magic
tech sky130l
timestamp 1731220306
<< checkpaint >>
rect -28 76 40 80
rect -28 12 68 76
rect -27 8 68 12
rect -24 -12 68 8
rect -24 -26 59 -12
rect -19 -28 54 -26
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 11 20 12
rect 15 8 16 11
rect 19 8 20 11
rect 15 6 20 8
rect 22 10 27 12
rect 22 7 23 10
rect 26 7 27 10
rect 22 6 27 7
<< ndc >>
rect 9 7 12 10
rect 16 8 19 11
rect 23 7 26 10
<< ntransistor >>
rect 13 6 15 12
rect 20 6 22 12
<< pdiffusion >>
rect 8 33 13 34
rect 8 30 9 33
rect 12 30 13 33
rect 8 19 13 30
rect 15 19 20 34
rect 22 23 27 34
rect 22 20 23 23
rect 26 20 27 23
rect 22 19 27 20
<< pdc >>
rect 9 30 12 33
rect 23 20 26 23
<< ptransistor >>
rect 13 19 15 34
rect 20 19 22 34
<< polysilicon >>
rect 10 43 15 44
rect 10 40 11 43
rect 14 40 15 43
rect 10 39 15 40
rect 13 34 15 39
rect 20 43 25 44
rect 20 40 21 43
rect 24 40 25 43
rect 20 39 25 40
rect 20 34 22 39
rect 13 12 15 19
rect 20 12 22 19
rect 13 4 15 6
rect 20 4 22 6
<< pc >>
rect 11 40 14 43
rect 21 40 24 43
<< m1 >>
rect 4 44 8 48
rect 5 43 8 44
rect 32 43 36 44
rect 5 40 11 43
rect 14 40 15 43
rect 20 40 21 43
rect 24 40 36 43
rect 9 33 12 34
rect 9 29 12 30
rect 32 23 36 24
rect 16 20 23 23
rect 26 20 36 23
rect 16 11 19 20
rect 9 10 12 11
rect 16 7 19 8
rect 23 10 26 11
rect 9 6 12 7
rect 23 6 26 7
<< m2c >>
rect 9 30 12 33
rect 9 7 12 10
rect 23 7 26 10
<< m2 >>
rect 8 33 13 34
rect 8 30 9 33
rect 12 30 13 33
rect 8 29 13 30
rect 8 10 27 11
rect 8 7 9 10
rect 12 7 23 10
rect 26 7 27 10
rect 8 6 27 7
<< labels >>
rlabel space 0 0 40 52 6 prboundary
rlabel ndiffusion 23 7 23 7 3 GND
rlabel ndiffusion 23 8 23 8 3 GND
rlabel ndiffusion 23 11 23 11 3 GND
rlabel ndiffusion 20 9 20 9 3 Y
rlabel pdiffusion 23 20 23 20 3 Y
rlabel pdiffusion 23 21 23 21 3 Y
rlabel pdiffusion 23 24 23 24 3 Y
rlabel polysilicon 21 35 21 35 3 B
rlabel polysilicon 21 40 21 40 3 B
rlabel polysilicon 21 44 21 44 3 B
rlabel polysilicon 21 5 21 5 3 B
rlabel ntransistor 21 7 21 7 3 B
rlabel polysilicon 21 13 21 13 3 B
rlabel ptransistor 21 20 21 20 3 B
rlabel ndiffusion 16 7 16 7 3 Y
rlabel ndiffusion 16 9 16 9 3 Y
rlabel ndiffusion 16 12 16 12 3 Y
rlabel polysilicon 14 35 14 35 3 A
rlabel polysilicon 14 5 14 5 3 A
rlabel ntransistor 14 7 14 7 3 A
rlabel polysilicon 14 13 14 13 3 A
rlabel ptransistor 14 20 14 20 3 A
rlabel polysilicon 11 40 11 40 3 A
rlabel polysilicon 11 41 11 41 3 A
rlabel polysilicon 11 44 11 44 3 A
rlabel pdiffusion 9 20 9 20 3 Vdd
rlabel m1 33 44 33 44 3 B
port 1 e
rlabel m1 33 24 33 24 3 Y
port 2 e
rlabel m1 24 11 24 11 3 GND
rlabel m1 25 41 25 41 3 B
port 1 e
rlabel pc 22 41 22 41 3 B
port 1 e
rlabel m1 27 21 27 21 3 Y
port 2 e
rlabel m1 21 41 21 41 3 B
port 1 e
rlabel pdc 24 21 24 21 3 Y
port 2 e
rlabel m1 24 7 24 7 3 GND
rlabel m1 17 8 17 8 3 Y
port 2 e
rlabel ndc 17 9 17 9 3 Y
port 2 e
rlabel m1 17 12 17 12 3 Y
port 2 e
rlabel m1 17 21 17 21 3 Y
port 2 e
rlabel m1 15 41 15 41 3 A
port 3 e
rlabel m1 10 7 10 7 3 GND
rlabel m1 10 11 10 11 3 GND
rlabel m1 10 30 10 30 3 Vdd
rlabel m1 10 34 10 34 3 Vdd
rlabel pc 12 41 12 41 3 A
port 3 e
rlabel m1 6 41 6 41 3 A
port 3 e
rlabel m1 6 44 6 44 3 A
port 3 e
rlabel m1 5 45 5 45 3 A
port 3 e
rlabel m2 27 8 27 8 3 GND
rlabel m2c 24 8 24 8 3 GND
rlabel m2 13 8 13 8 3 GND
rlabel m2 13 31 13 31 3 Vdd
rlabel m2c 10 8 10 8 3 GND
rlabel m2c 10 31 10 31 3 Vdd
rlabel m2 9 7 9 7 3 GND
rlabel m2 9 8 9 8 3 GND
rlabel m2 9 11 9 11 3 GND
rlabel m2 9 30 9 30 3 Vdd
rlabel m2 9 31 9 31 3 Vdd
rlabel m2 9 34 9 34 3 Vdd
<< end >>
