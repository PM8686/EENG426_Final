magic
tech sky130l
timestamp 1731220306
<< checkpaint >>
rect -24 103 76 104
rect -24 93 77 103
rect -24 92 79 93
rect -24 89 84 92
rect -24 87 97 89
rect -24 -14 102 87
rect -24 -16 97 -14
rect -16 -21 97 -16
rect -9 -27 60 -21
rect -8 -28 60 -27
<< ndiffusion >>
rect 8 26 13 28
rect 8 23 9 26
rect 12 23 13 26
rect 8 18 13 23
rect 15 18 20 28
rect 22 27 27 28
rect 22 24 23 27
rect 26 24 27 27
rect 22 18 27 24
rect 33 22 38 28
rect 33 19 34 22
rect 37 19 38 22
rect 33 18 38 19
rect 40 26 45 28
rect 40 23 41 26
rect 44 23 45 26
rect 40 18 45 23
rect 47 26 52 28
rect 47 23 48 26
rect 51 23 52 26
rect 47 18 52 23
rect 58 27 63 28
rect 58 24 59 27
rect 62 24 63 27
rect 58 18 63 24
rect 65 26 70 28
rect 65 23 66 26
rect 69 23 70 26
rect 65 18 70 23
<< ndc >>
rect 9 23 12 26
rect 23 24 26 27
rect 34 19 37 22
rect 41 23 44 26
rect 48 23 51 26
rect 59 24 62 27
rect 66 23 69 26
<< ntransistor >>
rect 13 18 15 28
rect 20 18 22 28
rect 38 18 40 28
rect 45 18 47 28
rect 63 18 65 28
<< pdiffusion >>
rect 8 47 13 55
rect 8 44 9 47
rect 12 44 13 47
rect 8 35 13 44
rect 15 50 19 55
rect 15 49 20 50
rect 15 46 16 49
rect 19 46 20 49
rect 15 35 20 46
rect 22 40 27 50
rect 58 47 63 55
rect 22 37 23 40
rect 26 37 27 40
rect 22 35 27 37
rect 33 39 38 45
rect 33 36 34 39
rect 37 36 38 39
rect 33 35 38 36
rect 40 35 45 45
rect 47 44 52 45
rect 47 41 48 44
rect 51 41 52 44
rect 47 35 52 41
rect 58 44 59 47
rect 62 44 63 47
rect 58 35 63 44
rect 65 39 70 55
rect 65 36 66 39
rect 69 36 70 39
rect 65 35 70 36
<< pdc >>
rect 9 44 12 47
rect 16 46 19 49
rect 23 37 26 40
rect 34 36 37 39
rect 48 41 51 44
rect 59 44 62 47
rect 66 36 69 39
<< ptransistor >>
rect 13 35 15 55
rect 20 35 22 50
rect 38 35 40 45
rect 45 35 47 45
rect 63 35 65 55
<< polysilicon >>
rect 8 62 15 63
rect 8 59 9 62
rect 12 59 15 62
rect 8 58 15 59
rect 41 60 47 61
rect 13 55 15 58
rect 20 57 28 58
rect 20 54 24 57
rect 27 54 28 57
rect 41 57 42 60
rect 45 57 47 60
rect 41 56 47 57
rect 20 53 28 54
rect 20 50 22 53
rect 35 52 40 53
rect 35 49 36 52
rect 39 49 40 52
rect 35 48 40 49
rect 38 45 40 48
rect 45 45 47 56
rect 63 55 65 57
rect 13 28 15 35
rect 20 28 22 35
rect 38 28 40 35
rect 45 28 47 35
rect 63 28 65 35
rect 13 16 15 18
rect 20 16 22 18
rect 38 16 40 18
rect 45 16 47 18
rect 63 16 65 18
rect 60 15 65 16
rect 60 12 61 15
rect 64 12 65 15
rect 60 11 65 12
<< pc >>
rect 9 59 12 62
rect 24 54 27 57
rect 42 57 45 60
rect 36 49 39 52
rect 61 12 64 15
<< m1 >>
rect 8 68 12 72
rect 9 62 12 68
rect 24 68 28 72
rect 40 71 44 72
rect 40 68 45 71
rect 9 58 12 59
rect 16 59 19 60
rect 16 49 19 56
rect 24 57 27 68
rect 42 60 45 68
rect 42 56 45 57
rect 48 59 51 60
rect 24 52 27 54
rect 24 49 36 52
rect 39 49 40 52
rect 9 47 12 48
rect 16 45 19 46
rect 9 43 12 44
rect 48 44 51 56
rect 59 47 62 48
rect 59 43 62 44
rect 48 40 51 41
rect 17 37 23 40
rect 26 37 27 40
rect 34 39 37 40
rect 8 26 12 27
rect 8 23 9 26
rect 8 16 12 23
rect 17 15 20 37
rect 17 11 20 12
rect 23 33 26 34
rect 23 27 26 30
rect 34 33 37 36
rect 65 36 66 39
rect 69 36 70 39
rect 34 29 37 30
rect 59 33 62 34
rect 65 33 70 36
rect 65 30 66 33
rect 69 30 70 33
rect 59 27 62 30
rect 23 8 26 24
rect 41 26 44 27
rect 34 22 37 23
rect 41 22 44 23
rect 48 26 51 27
rect 59 23 62 24
rect 66 26 69 27
rect 48 22 51 23
rect 66 22 69 23
rect 34 15 37 19
rect 34 11 37 12
rect 61 15 64 16
rect 61 11 64 12
rect 23 5 28 8
rect 24 4 28 5
<< m2c >>
rect 16 56 19 59
rect 48 56 51 59
rect 9 44 12 47
rect 59 44 62 47
rect 9 23 12 26
rect 17 12 20 15
rect 23 30 26 33
rect 34 30 37 33
rect 59 30 62 33
rect 66 30 69 33
rect 41 23 44 26
rect 48 23 51 26
rect 66 23 69 26
rect 34 12 37 15
rect 61 12 64 15
<< m2 >>
rect 15 59 52 60
rect 15 56 16 59
rect 19 56 48 59
rect 51 56 52 59
rect 15 55 52 56
rect 8 47 63 48
rect 8 44 9 47
rect 12 44 59 47
rect 62 44 63 47
rect 8 43 63 44
rect 22 33 70 34
rect 22 30 23 33
rect 26 30 34 33
rect 37 30 59 33
rect 62 30 66 33
rect 69 30 70 33
rect 22 29 70 30
rect 8 26 45 27
rect 8 23 9 26
rect 12 23 41 26
rect 44 23 45 26
rect 8 22 45 23
rect 47 26 70 27
rect 47 23 48 26
rect 51 23 66 26
rect 69 23 70 26
rect 47 22 70 23
rect 16 15 65 16
rect 16 12 17 15
rect 20 12 34 15
rect 37 12 61 15
rect 64 12 65 15
rect 16 11 65 12
<< labels >>
rlabel space 0 0 80 76 6 prboundary
rlabel ndiffusion 63 25 63 25 3 _q
rlabel ndiffusion 66 19 66 19 3 #10
rlabel ndiffusion 66 24 66 24 3 #10
rlabel ndiffusion 66 27 66 27 3 #10
rlabel ndiffusion 59 25 59 25 3 _q
rlabel pdiffusion 66 36 66 36 3 _q
rlabel pdiffusion 66 40 66 40 3 _q
rlabel ntransistor 64 19 64 19 3 _clk
rlabel polysilicon 64 29 64 29 3 _clk
rlabel ptransistor 64 36 64 36 3 _clk
rlabel polysilicon 64 56 64 56 3 _clk
rlabel ndiffusion 59 19 59 19 3 _q
rlabel ndiffusion 59 28 59 28 3 _q
rlabel pdiffusion 59 36 59 36 3 #7
rlabel pdiffusion 59 45 59 45 3 #7
rlabel pdiffusion 59 48 59 48 3 #7
rlabel pdiffusion 52 42 52 42 3 Vdd
rlabel polysilicon 46 58 46 58 3 q
rlabel polysilicon 46 46 46 46 3 q
rlabel ndiffusion 48 19 48 19 3 #10
rlabel pdiffusion 48 36 48 36 3 Vdd
rlabel pdiffusion 48 42 48 42 3 Vdd
rlabel pdiffusion 48 45 48 45 3 Vdd
rlabel polysilicon 42 57 42 57 3 q
rlabel polysilicon 42 58 42 58 3 q
rlabel polysilicon 42 61 42 61 3 q
rlabel polysilicon 64 17 64 17 3 _clk
rlabel ntransistor 46 19 46 19 3 q
rlabel polysilicon 46 29 46 29 3 q
rlabel ptransistor 46 36 46 36 3 q
rlabel ndiffusion 41 19 41 19 3 GND
rlabel ndiffusion 41 24 41 24 3 GND
rlabel ndiffusion 41 27 41 27 3 GND
rlabel ndiffusion 38 20 38 20 3 _clk
rlabel pdiffusion 38 37 38 37 3 _q
rlabel polysilicon 39 46 39 46 3 CLK
rlabel polysilicon 46 17 46 17 3 q
rlabel ntransistor 39 19 39 19 3 CLK
rlabel polysilicon 39 29 39 29 3 CLK
rlabel ptransistor 39 36 39 36 3 CLK
rlabel polysilicon 36 49 36 49 3 CLK
rlabel polysilicon 36 50 36 50 3 CLK
rlabel polysilicon 36 53 36 53 3 CLK
rlabel ndiffusion 34 19 34 19 3 _clk
rlabel ndiffusion 34 20 34 20 3 _clk
rlabel ndiffusion 34 23 34 23 3 _clk
rlabel ndiffusion 27 25 27 25 3 _q
rlabel pdiffusion 34 36 34 36 3 _q
rlabel pdiffusion 34 37 34 37 3 _q
rlabel pdiffusion 34 40 34 40 3 _q
rlabel polysilicon 28 55 28 55 3 CLK
rlabel polysilicon 39 17 39 17 3 CLK
rlabel ndiffusion 23 19 23 19 3 _q
rlabel ndiffusion 23 25 23 25 3 _q
rlabel ndiffusion 23 28 23 28 3 _q
rlabel pdiffusion 23 36 23 36 3 _clk
rlabel pdiffusion 23 38 23 38 3 _clk
rlabel pdiffusion 23 41 23 41 3 _clk
rlabel pdiffusion 20 47 20 47 3 Vdd
rlabel polysilicon 21 51 21 51 3 CLK
rlabel polysilicon 21 54 21 54 3 CLK
rlabel polysilicon 21 55 21 55 3 CLK
rlabel polysilicon 21 58 21 58 3 CLK
rlabel polysilicon 21 17 21 17 3 CLK
rlabel ntransistor 21 19 21 19 3 CLK
rlabel polysilicon 21 29 21 29 3 CLK
rlabel ptransistor 21 36 21 36 3 CLK
rlabel polysilicon 61 12 61 12 3 _clk
rlabel polysilicon 61 13 61 13 3 _clk
rlabel polysilicon 61 16 61 16 3 _clk
rlabel pdiffusion 16 36 16 36 3 Vdd
rlabel pdiffusion 16 47 16 47 3 Vdd
rlabel pdiffusion 16 50 16 50 3 Vdd
rlabel pdiffusion 16 51 16 51 3 Vdd
rlabel polysilicon 13 60 13 60 3 D
rlabel polysilicon 14 17 14 17 3 D
rlabel ntransistor 14 19 14 19 3 D
rlabel polysilicon 14 29 14 29 3 D
rlabel ptransistor 14 36 14 36 3 D
rlabel polysilicon 14 56 14 56 3 D
rlabel ndiffusion 9 19 9 19 3 GND
rlabel pdiffusion 9 36 9 36 3 #7
rlabel polysilicon 9 59 9 59 3 D
rlabel polysilicon 9 60 9 60 3 D
rlabel polysilicon 9 63 9 63 3 D
rlabel m1 70 37 70 37 3 _q
port 1 e
rlabel m1 67 27 67 27 3 #10
rlabel pdc 67 37 67 37 3 _q
port 1 e
rlabel m1 41 69 41 69 3 q
port 2 e
rlabel m1 41 72 41 72 3 q
port 2 e
rlabel m1 67 23 67 23 3 #10
rlabel m1 66 31 66 31 3 _q
port 1 e
rlabel m1 66 34 66 34 3 _q
port 1 e
rlabel m1 66 37 66 37 3 _q
port 1 e
rlabel m1 49 60 49 60 3 Vdd
rlabel m1 49 23 49 23 3 #10
rlabel m1 60 24 60 24 3 _q
port 1 e
rlabel ndc 60 25 60 25 3 _q
port 1 e
rlabel m1 60 28 60 28 3 _q
port 1 e
rlabel m1 60 34 60 34 3 _q
port 1 e
rlabel m1 60 44 60 44 3 #7
rlabel m1 60 48 60 48 3 #7
rlabel m1 43 57 43 57 3 q
port 2 e
rlabel pc 43 58 43 58 3 q
port 2 e
rlabel m1 43 61 43 61 3 q
port 2 e
rlabel m1 35 40 35 40 3 _q
port 1 e
rlabel m1 40 50 40 50 3 CLK
port 3 e
rlabel m1 62 12 62 12 3 _clk
rlabel m1 62 16 62 16 3 _clk
rlabel m1 42 23 42 23 3 GND
rlabel m1 49 27 49 27 3 #10
rlabel m1 49 41 49 41 3 Vdd
rlabel pdc 49 42 49 42 3 Vdd
rlabel m1 49 45 49 45 3 Vdd
rlabel m1 42 27 42 27 3 GND
rlabel pc 37 50 37 50 3 CLK
port 3 e
rlabel m1 35 30 35 30 3 _q
port 1 e
rlabel m1 35 34 35 34 3 _q
port 1 e
rlabel pdc 35 37 35 37 3 _q
port 1 e
rlabel m1 27 38 27 38 3 _clk
rlabel m1 25 50 25 50 3 CLK
port 3 e
rlabel m1 25 53 25 53 3 CLK
port 3 e
rlabel pc 25 55 25 55 3 CLK
port 3 e
rlabel m1 25 58 25 58 3 CLK
port 3 e
rlabel m1 25 69 25 69 3 CLK
port 3 e
rlabel m1 35 12 35 12 3 _clk
rlabel m1 35 16 35 16 3 _clk
rlabel ndc 35 20 35 20 3 _clk
rlabel m1 35 23 35 23 3 _clk
rlabel pdc 24 38 24 38 3 _clk
rlabel m1 25 5 25 5 3 _q
port 1 e
rlabel ndc 24 25 24 25 3 _q
port 1 e
rlabel m1 24 28 24 28 3 _q
port 1 e
rlabel m1 24 34 24 34 3 _q
port 1 e
rlabel m1 18 38 18 38 3 _clk
rlabel m1 24 6 24 6 3 _q
port 1 e
rlabel m1 24 9 24 9 3 _q
port 1 e
rlabel m1 17 46 17 46 3 Vdd
rlabel pdc 17 47 17 47 3 Vdd
rlabel m1 17 50 17 50 3 Vdd
rlabel m1 17 60 17 60 3 Vdd
rlabel m1 18 12 18 12 3 _clk
rlabel m1 18 16 18 16 3 _clk
rlabel m1 10 44 10 44 3 #7
rlabel m1 10 48 10 48 3 #7
rlabel m1 10 59 10 59 3 D
port 4 e
rlabel pc 10 60 10 60 3 D
port 4 e
rlabel m1 10 63 10 63 3 D
port 4 e
rlabel m1 9 17 9 17 3 GND
rlabel m1 9 69 9 69 3 D
port 4 e
rlabel m2 70 31 70 31 3 _q
port 1 e
rlabel m2c 67 31 67 31 3 _q
port 1 e
rlabel m2 63 31 63 31 3 _q
port 1 e
rlabel m2c 60 31 60 31 3 _q
port 1 e
rlabel m2 70 24 70 24 3 #10
rlabel m2 38 31 38 31 3 _q
port 1 e
rlabel m2c 67 24 67 24 3 #10
rlabel m2c 35 31 35 31 3 _q
port 1 e
rlabel m2 65 13 65 13 3 _clk
rlabel m2 52 24 52 24 3 #10
rlabel m2 27 31 27 31 3 _q
port 1 e
rlabel m2c 62 13 62 13 3 _clk
rlabel m2c 49 24 49 24 3 #10
rlabel m2c 24 31 24 31 3 _q
port 1 e
rlabel m2 52 57 52 57 3 Vdd
rlabel m2 38 13 38 13 3 _clk
rlabel m2 48 24 48 24 3 #10
rlabel m2 23 30 23 30 3 _q
port 1 e
rlabel m2 23 31 23 31 3 _q
port 1 e
rlabel m2 23 34 23 34 3 _q
port 1 e
rlabel m2c 49 57 49 57 3 Vdd
rlabel m2c 35 13 35 13 3 _clk
rlabel m2 20 57 20 57 3 Vdd
rlabel m2 21 13 21 13 3 _clk
rlabel m2 45 24 45 24 3 GND
rlabel m2 63 45 63 45 3 #7
rlabel m2c 17 57 17 57 3 Vdd
rlabel m2c 18 13 18 13 3 _clk
rlabel m2c 42 24 42 24 3 GND
rlabel m2c 60 45 60 45 3 #7
rlabel m2 16 56 16 56 3 Vdd
rlabel m2 16 57 16 57 3 Vdd
rlabel m2 16 60 16 60 3 Vdd
rlabel m2 17 12 17 12 3 _clk
rlabel m2 17 13 17 13 3 _clk
rlabel m2 17 16 17 16 3 _clk
rlabel m2 48 23 48 23 3 #10
rlabel m2 13 24 13 24 3 GND
rlabel m2 48 27 48 27 3 #10
rlabel m2 13 45 13 45 3 #7
rlabel m2c 10 24 10 24 3 GND
rlabel m2c 10 45 10 45 3 #7
rlabel m2 9 23 9 23 3 GND
rlabel m2 9 24 9 24 3 GND
rlabel m2 9 27 9 27 3 GND
rlabel m2 9 44 9 44 3 #7
rlabel m2 9 45 9 45 3 #7
rlabel m2 9 48 9 48 3 #7
<< end >>
