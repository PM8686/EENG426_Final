VERSION 5.6 ;

BUSBITCHARS "[]" ;

DIVIDERCHAR "/" ;

UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005000 ; 

CLEARANCEMEASURE EUCLIDEAN ; 

USEMINSPACING OBS ON ; 

SITE CoreSite
    CLASS CORE ;
    SIZE 0.540000 BY 0.900000 ;
END CoreSite

LAYER m1
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.270000 ;
   WIDTH 0.270000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.270000 ;
   PITCH 0.540000 0.540000 ;
END m1

LAYER v1
    TYPE CUT ;
    SPACING 0.270000 ;
    WIDTH 0.270000 ;
    ENCLOSURE ABOVE 0.090000 0.090000 ;
    ENCLOSURE BELOW 0.090000 0.090000 ;
END v1

LAYER m2
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.450000 ;
   WIDTH 0.450000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.450000 ;
   PITCH 0.900000 0.900000 ;
END m2

LAYER v2
    TYPE CUT ;
    SPACING 0.270000 ;
    WIDTH 0.270000 ;
    ENCLOSURE ABOVE 0.090000 0.090000 ;
    ENCLOSURE BELOW 0.090000 0.090000 ;
END v2

LAYER m3
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.450000 ;
   WIDTH 0.450000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.450000 ;
   PITCH 0.900000 0.900000 ;
END m3

LAYER v3
    TYPE CUT ;
    SPACING 0.270000 ;
    WIDTH 0.270000 ;
    ENCLOSURE ABOVE 0.090000 0.090000 ;
    ENCLOSURE BELOW 0.090000 0.090000 ;
END v3

LAYER m4
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.450000 ;
   WIDTH 0.450000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.450000 ;
   PITCH 0.900000 0.900000 ;
END m4

LAYER v4
    TYPE CUT ;
    SPACING 0.270000 ;
    WIDTH 0.270000 ;
    ENCLOSURE ABOVE 0.090000 0.090000 ;
    ENCLOSURE BELOW 0.090000 0.090000 ;
END v4

LAYER m5
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.450000 ;
   WIDTH 0.450000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.450000 ;
   PITCH 0.900000 0.900000 ;
END m5

LAYER v5
    TYPE CUT ;
    SPACING 0.270000 ;
    WIDTH 0.270000 ;
    ENCLOSURE ABOVE 0.090000 0.090000 ;
    ENCLOSURE BELOW 0.090000 0.090000 ;
END v5

LAYER m6
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.450000 ;
   WIDTH 0.450000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.450000 ;
   PITCH 0.900000 0.900000 ;
END m6

LAYER OVERLAP
   TYPE OVERLAP ;
END OVERLAP

VIA v1_C DEFAULT
   LAYER m1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v1 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v1_C

VIA v1_Ch
   LAYER m1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v1 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v1_Ch

VIA v1_Cv
   LAYER m1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v1 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v1_Cv

VIA v2_C DEFAULT
   LAYER m2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v2 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_C

VIA v2_Ch
   LAYER m2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v2 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_Ch

VIA v2_Cv
   LAYER m2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v2 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_Cv

VIA v3_C DEFAULT
   LAYER m3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v3 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m4 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v3_C

VIA v3_Ch
   LAYER m3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v3 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m4 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v3_Ch

VIA v3_Cv
   LAYER m3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v3 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m4 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v3_Cv

VIA v4_C DEFAULT
   LAYER m4 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v4 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m5 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v4_C

VIA v4_Ch
   LAYER m4 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v4 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m5 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v4_Ch

VIA v4_Cv
   LAYER m4 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v4 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m5 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v4_Cv

VIA v5_C DEFAULT
   LAYER m5 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v5 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m6 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v5_C

VIA v5_Ch
   LAYER m5 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v5 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m6 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v5_Ch

VIA v5_Cv
   LAYER m5 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v5 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m6 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v5_Cv

MACRO _0_0cell_0_0g0n_0x0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g0n_0x0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 3.240000 BY 9.900000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 8.730000 0.810000 9.000000 ;
        END
    END in_50_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 0.900000 0.810000 1.170000 ;
        END
        ANTENNADIFFAREA 3.888000 ;
    END out
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 1.620000 8.730000 1.890000 9.000000 ;
        END
        ANTENNADIFFAREA 3.888000 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 2.700000 8.730000 2.970000 9.000000 ;
        END
        ANTENNADIFFAREA 0.972000 ;
    END GND
    OBS
      LAYER m1 ;
         RECT 0.540000 1.620000 2.610000 8.190000 ;
    END
END _0_0cell_0_0g0n_0x0

MACRO _0_0std_0_0cells_0_0INVX1
    CLASS CORE ;
    FOREIGN _0_0std_0_0cells_0_0INVX1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.160000 BY 5.400000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 4.230000 0.810000 4.500000 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 0.900000 0.810000 1.170000 ;
        END
        ANTENNADIFFAREA 0.631800 ;
    END Y
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 1.080000 4.230000 1.350000 4.500000 ;
        END
        ANTENNADIFFAREA 0.388800 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 1.620000 4.230000 1.890000 4.500000 ;
        END
        ANTENNADIFFAREA 0.243000 ;
    END GND
    OBS
      LAYER m1 ;
         RECT 0.540000 1.620000 1.530000 3.690000 ;
    END
END _0_0std_0_0cells_0_0INVX1

MACRO _0_0std_0_0cells_0_0AND2X1
    CLASS CORE ;
    FOREIGN _0_0std_0_0cells_0_0AND2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 5.400000 BY 7.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 1.620000 6.030000 2.970000 6.300000 ;
        RECT 2.700000 5.760000 2.970000 6.030000 ;
        RECT 2.700000 5.670000 3.060000 5.760000 ;
        RECT 2.700000 5.490000 2.790000 5.670000 ;
        RECT 2.700000 5.400000 3.060000 5.490000 ;
        RECT 2.790000 5.490000 2.970000 5.670000 ;
        RECT 2.970000 5.490000 3.060000 5.670000 ;
        END
        ANTENNAGATEAREA 0.291600 ;
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 1.620000 1.710000 1.980000 1.800000 ;
        RECT 1.620000 1.530000 1.710000 1.710000 ;
        RECT 1.620000 1.440000 1.980000 1.530000 ;
        RECT 1.620000 0.990000 1.890000 1.440000 ;
        RECT 1.710000 1.530000 1.890000 1.710000 ;
        RECT 1.890000 1.530000 1.980000 1.710000 ;
        END
        ANTENNAGATEAREA 0.291600 ;
    END B
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 3.960000 4.320000 4.320000 4.410000 ;
        RECT 3.960000 2.520000 4.320000 2.610000 ;
        RECT 3.960000 2.790000 4.320000 2.880000 ;
        RECT 3.960000 2.610000 4.050000 2.790000 ;
        RECT 4.050000 6.030000 5.130000 6.300000 ;
        RECT 4.050000 4.680000 4.320000 6.030000 ;
        RECT 3.960000 4.590000 4.320000 4.680000 ;
        RECT 3.960000 4.410000 4.050000 4.590000 ;
        RECT 4.050000 2.880000 4.320000 4.320000 ;
        RECT 4.050000 2.610000 4.230000 2.790000 ;
        RECT 4.050000 4.410000 4.230000 4.590000 ;
        RECT 4.230000 2.610000 4.320000 2.790000 ;
        RECT 4.230000 4.410000 4.320000 4.590000 ;
        END
        ANTENNADIFFAREA 0.631800 ;
    END Y
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 1.620000 5.040000 2.070000 5.130000 ;
        RECT 1.620000 4.770000 1.710000 5.040000 ;
        RECT 1.620000 4.680000 2.070000 4.770000 ;
        RECT 1.710000 4.950000 1.980000 5.040000 ;
        RECT 1.710000 4.770000 1.890000 4.950000 ;
        RECT 1.890000 4.770000 1.980000 4.950000 ;
        RECT 1.980000 4.770000 2.070000 5.040000 ;
        RECT 2.970000 5.040000 3.420000 5.130000 ;
        RECT 2.970000 4.770000 3.060000 5.040000 ;
        RECT 2.970000 4.680000 3.420000 4.770000 ;
        RECT 3.060000 4.950000 3.330000 5.040000 ;
        RECT 3.060000 4.770000 3.150000 4.950000 ;
        RECT 3.150000 4.770000 3.330000 4.950000 ;
        RECT 3.330000 4.770000 3.420000 5.040000 ;
        LAYER v1 ;
        RECT 1.710000 4.950000 1.980000 5.040000 ;
        RECT 1.710000 4.770000 1.890000 4.950000 ;
        RECT 1.890000 4.770000 1.980000 4.950000 ;
        RECT 3.060000 4.950000 3.330000 5.040000 ;
        RECT 3.060000 4.770000 3.150000 4.950000 ;
        RECT 3.150000 4.770000 3.330000 4.950000 ;
        LAYER m2 ;
        RECT 0.630000 5.040000 3.420000 5.130000 ;
        RECT 0.630000 4.770000 1.710000 5.040000 ;
        RECT 0.630000 4.680000 3.420000 4.770000 ;
        RECT 1.710000 4.950000 1.980000 5.040000 ;
        RECT 1.710000 4.770000 1.890000 4.950000 ;
        RECT 1.890000 4.770000 1.980000 4.950000 ;
        RECT 1.980000 4.770000 3.060000 5.040000 ;
        RECT 3.060000 4.950000 3.330000 5.040000 ;
        RECT 3.060000 4.770000 3.150000 4.950000 ;
        RECT 3.150000 4.770000 3.330000 4.950000 ;
        RECT 3.330000 4.770000 3.420000 5.040000 ;
        END
        ANTENNADIFFAREA 0.777600 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 2.970000 2.250000 3.420000 2.340000 ;
        RECT 2.970000 1.980000 3.060000 2.250000 ;
        RECT 2.970000 1.890000 3.420000 1.980000 ;
        RECT 3.060000 2.070000 3.150000 2.250000 ;
        RECT 3.060000 1.980000 3.330000 2.070000 ;
        RECT 3.150000 2.070000 3.330000 2.250000 ;
        RECT 3.330000 1.980000 3.420000 2.250000 ;
        LAYER v1 ;
        RECT 3.060000 2.070000 3.150000 2.250000 ;
        RECT 3.060000 1.980000 3.330000 2.070000 ;
        RECT 3.150000 2.070000 3.330000 2.250000 ;
        LAYER m2 ;
        RECT 2.970000 2.250000 3.420000 2.340000 ;
        RECT 2.970000 1.980000 3.060000 2.250000 ;
        RECT 2.970000 0.900000 3.420000 1.980000 ;
        RECT 3.060000 2.070000 3.150000 2.250000 ;
        RECT 3.060000 1.980000 3.330000 2.070000 ;
        RECT 3.150000 2.070000 3.330000 2.250000 ;
        RECT 3.330000 1.980000 3.420000 2.250000 ;
        END
        ANTENNADIFFAREA 0.405000 ;
    END GND
    OBS
        LAYER m1 ;
        RECT 1.620000 3.690000 2.070000 3.780000 ;
        RECT 1.620000 3.420000 1.710000 3.690000 ;
        RECT 1.620000 3.330000 2.070000 3.420000 ;
        RECT 1.710000 3.420000 1.980000 3.690000 ;
        RECT 1.710000 2.790000 2.070000 2.880000 ;
        RECT 1.710000 2.610000 1.800000 2.790000 ;
        RECT 1.710000 2.520000 2.070000 2.610000 ;
        RECT 2.340000 4.590000 2.700000 4.680000 ;
        RECT 2.340000 4.410000 2.430000 4.590000 ;
        RECT 2.340000 4.320000 2.700000 4.410000 ;
        RECT 2.340000 3.780000 2.610000 4.320000 ;
        RECT 2.340000 3.690000 2.790000 3.780000 ;
        RECT 1.980000 3.420000 2.070000 3.690000 ;
        RECT 2.340000 3.330000 2.790000 3.420000 ;
        RECT 1.800000 2.880000 2.070000 3.330000 ;
        RECT 1.800000 2.610000 1.980000 2.790000 ;
        RECT 2.430000 4.410000 2.610000 4.590000 ;
        RECT 1.980000 2.610000 2.070000 2.790000 ;
        RECT 2.610000 4.410000 2.700000 4.590000 ;
        RECT 2.340000 3.420000 2.430000 3.690000 ;
        RECT 2.430000 3.420000 2.700000 3.690000 ;
        RECT 2.700000 3.420000 2.790000 3.690000 ;
        RECT 4.590000 3.690000 5.040000 3.780000 ;
        RECT 4.590000 3.420000 4.680000 3.690000 ;
        RECT 4.590000 3.330000 5.040000 3.420000 ;
        RECT 4.680000 3.600000 4.950000 3.690000 ;
        RECT 4.680000 3.420000 4.860000 3.600000 ;
        RECT 4.860000 3.420000 4.950000 3.600000 ;
        RECT 4.950000 3.420000 5.040000 3.690000 ;
        LAYER m2 ;
        RECT 1.620000 3.690000 5.040000 3.780000 ;
        RECT 1.620000 3.420000 1.710000 3.690000 ;
        RECT 1.620000 3.330000 5.040000 3.420000 ;
        RECT 1.710000 3.420000 1.980000 3.690000 ;
        RECT 1.980000 3.420000 2.430000 3.690000 ;
        RECT 2.430000 3.420000 2.700000 3.690000 ;
        RECT 2.700000 3.420000 4.680000 3.690000 ;
        RECT 4.680000 3.600000 4.950000 3.690000 ;
        RECT 4.680000 3.420000 4.860000 3.600000 ;
        RECT 4.860000 3.420000 4.950000 3.600000 ;
        RECT 4.950000 3.420000 5.040000 3.690000 ;
    END
END _0_0std_0_0cells_0_0AND2X1

MACRO _0_0std_0_0cells_0_0NOR2X1
    CLASS CORE ;
    FOREIGN _0_0std_0_0cells_0_0NOR2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 3.780000 BY 7.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.990000 2.070000 1.350000 2.160000 ;
        RECT 0.990000 1.890000 1.080000 2.070000 ;
        RECT 0.990000 1.800000 1.350000 1.890000 ;
        RECT 1.080000 1.890000 1.260000 2.070000 ;
        RECT 1.260000 1.890000 1.350000 2.070000 ;
        END
        ANTENNAGATEAREA 0.324000 ;
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 1.710000 6.210000 2.070000 6.300000 ;
        RECT 1.710000 6.030000 1.800000 6.210000 ;
        RECT 1.710000 5.940000 2.070000 6.030000 ;
        RECT 1.800000 6.030000 1.980000 6.210000 ;
        RECT 1.980000 6.030000 2.070000 6.210000 ;
        END
        ANTENNAGATEAREA 0.324000 ;
    END B
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 1.350000 2.790000 1.800000 2.880000 ;
        RECT 1.350000 5.220000 1.800000 5.310000 ;
        RECT 1.350000 4.860000 1.800000 4.950000 ;
        RECT 1.440000 2.880000 1.710000 4.860000 ;
        RECT 1.350000 2.520000 1.440000 2.790000 ;
        RECT 1.350000 4.950000 1.440000 5.220000 ;
        RECT 1.440000 2.520000 1.710000 2.790000 ;
        RECT 1.350000 2.430000 1.800000 2.520000 ;
        RECT 1.440000 4.950000 1.710000 5.220000 ;
        RECT 1.710000 2.520000 1.800000 2.790000 ;
        RECT 1.710000 4.950000 1.800000 5.220000 ;
        RECT 2.880000 4.950000 3.060000 5.130000 ;
        LAYER v1 ;
        RECT 1.440000 4.950000 1.710000 5.220000 ;
        LAYER m2 ;
        RECT 1.440000 4.950000 1.710000 5.220000 ;
        RECT 1.710000 4.950000 1.800000 5.220000 ;
        END
        ANTENNADIFFAREA 2.551500 ;
    END Y
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 0.540000 5.220000 0.990000 5.310000 ;
        RECT 0.540000 4.950000 0.630000 5.220000 ;
        RECT 0.540000 4.860000 0.990000 4.950000 ;
        RECT 0.630000 4.950000 0.900000 5.220000 ;
        RECT 0.900000 4.950000 0.990000 5.220000 ;
        RECT 2.790000 5.220000 3.060000 6.210000 ;
        RECT 2.790000 5.130000 3.150000 5.220000 ;
        RECT 2.790000 4.950000 2.880000 5.130000 ;
        RECT 2.790000 4.860000 3.150000 4.950000 ;
        RECT 3.060000 4.950000 3.150000 5.130000 ;
        LAYER v1 ;
        RECT 0.630000 4.950000 0.900000 5.220000 ;
        LAYER m2 ;
        RECT 0.540000 5.220000 1.800000 5.310000 ;
        RECT 0.540000 4.950000 0.630000 5.220000 ;
        RECT 0.540000 4.860000 1.800000 4.950000 ;
        RECT 0.630000 4.950000 0.900000 5.220000 ;
        RECT 0.900000 4.950000 1.440000 5.220000 ;
        END
        ANTENNADIFFAREA 0.850500 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 0.450000 2.700000 0.810000 2.790000 ;
        RECT 0.450000 2.520000 0.540000 2.700000 ;
        RECT 0.450000 2.430000 0.810000 2.520000 ;
        RECT 0.450000 1.530000 0.720000 2.430000 ;
        RECT 0.450000 1.440000 0.900000 1.530000 ;
        RECT 0.450000 1.170000 0.540000 1.440000 ;
        RECT 0.450000 1.080000 0.900000 1.170000 ;
        RECT 0.540000 2.520000 0.720000 2.700000 ;
        RECT 0.540000 1.170000 0.810000 1.440000 ;
        RECT 0.720000 2.520000 0.810000 2.700000 ;
        RECT 0.810000 1.170000 0.900000 1.440000 ;
        RECT 2.070000 1.440000 2.520000 1.530000 ;
        RECT 2.070000 1.170000 2.160000 1.440000 ;
        RECT 2.070000 1.080000 2.520000 1.170000 ;
        RECT 2.250000 1.530000 2.520000 2.430000 ;
        RECT 2.160000 1.170000 2.430000 1.440000 ;
        RECT 2.430000 1.170000 2.520000 1.440000 ;
        RECT 2.160000 2.430000 2.520000 2.520000 ;
        RECT 2.160000 2.700000 2.520000 2.790000 ;
        RECT 2.160000 2.520000 2.250000 2.700000 ;
        RECT 2.250000 2.520000 2.430000 2.700000 ;
        RECT 2.430000 2.520000 2.520000 2.700000 ;
        LAYER v1 ;
        RECT 0.540000 1.170000 0.810000 1.440000 ;
        RECT 2.160000 1.170000 2.430000 1.440000 ;
        LAYER m2 ;
        RECT 0.450000 1.440000 2.520000 1.530000 ;
        RECT 0.450000 1.170000 0.540000 1.440000 ;
        RECT 0.450000 1.080000 2.520000 1.170000 ;
        RECT 0.540000 1.170000 0.810000 1.440000 ;
        RECT 0.810000 1.170000 2.160000 1.440000 ;
        RECT 2.160000 1.170000 2.430000 1.440000 ;
        RECT 2.430000 1.170000 2.520000 1.440000 ;
        END
        ANTENNADIFFAREA 0.810000 ;
    END GND
END _0_0std_0_0cells_0_0NOR2X1

MACRO _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 6.480000 BY 10.800000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 9.630000 0.810000 9.900000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 1.620000 9.630000 1.890000 9.900000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 2.700000 9.630000 2.970000 9.900000 ;
        END
    END in_52_6
    PIN in_53_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 3.780000 9.630000 4.050000 9.900000 ;
        END
    END in_53_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 0.900000 0.810000 1.170000 ;
        END
        ANTENNADIFFAREA 2.138400 ;
    END out
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 4.860000 9.630000 5.130000 9.900000 ;
        END
        ANTENNADIFFAREA 5.054400 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 5.940000 9.630000 6.210000 9.900000 ;
        END
        ANTENNADIFFAREA 1.944000 ;
    END GND
    OBS
      LAYER m1 ;
         RECT 0.540000 1.620000 5.850000 9.090000 ;
    END
END _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0

MACRO _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 5.400000 BY 7.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 6.030000 0.810000 6.300000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 1.620000 6.030000 1.890000 6.300000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 2.700000 6.030000 2.970000 6.300000 ;
        END
    END in_52_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 0.900000 0.810000 1.170000 ;
        END
        ANTENNADIFFAREA 1.603800 ;
    END out
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 3.780000 6.030000 4.050000 6.300000 ;
        END
        ANTENNADIFFAREA 1.652400 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 4.860000 6.030000 5.130000 6.300000 ;
        END
        ANTENNADIFFAREA 0.972000 ;
    END GND
    OBS
      LAYER m1 ;
         RECT 0.540000 1.620000 4.770000 5.490000 ;
    END
END _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0

MACRO _0_0cell_0_0g0n_0x2
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g0n_0x2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.160000 BY 5.400000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 4.230000 0.810000 4.500000 ;
        END
    END in_50_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 0.900000 0.810000 1.170000 ;
        END
        ANTENNADIFFAREA 0.631800 ;
    END out
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 1.080000 4.230000 1.350000 4.500000 ;
        END
        ANTENNADIFFAREA 0.388800 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 1.620000 4.230000 1.890000 4.500000 ;
        END
        ANTENNADIFFAREA 0.243000 ;
    END GND
    OBS
      LAYER m1 ;
         RECT 0.540000 1.620000 1.530000 3.690000 ;
    END
END _0_0cell_0_0g0n_0x2

MACRO _0_0std_0_0cells_0_0OR2X1
    CLASS CORE ;
    FOREIGN _0_0std_0_0cells_0_0OR2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 4.860000 BY 6.300000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 1.710000 5.940000 2.070000 6.030000 ;
        RECT 1.710000 5.760000 1.800000 5.940000 ;
        RECT 1.710000 5.670000 2.070000 5.760000 ;
        RECT 1.800000 5.760000 1.980000 5.940000 ;
        RECT 1.980000 5.760000 2.070000 5.940000 ;
        END
        ANTENNAGATEAREA 0.324000 ;
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.990000 5.310000 1.350000 5.400000 ;
        RECT 0.990000 5.130000 1.080000 5.310000 ;
        RECT 0.990000 5.040000 1.350000 5.130000 ;
        RECT 1.080000 5.130000 1.260000 5.310000 ;
        RECT 1.260000 5.130000 1.350000 5.310000 ;
        END
        ANTENNAGATEAREA 0.324000 ;
    END B
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 3.150000 1.530000 3.510000 1.620000 ;
        RECT 3.240000 1.890000 3.510000 3.600000 ;
        RECT 3.150000 3.870000 3.510000 3.960000 ;
        RECT 3.150000 3.600000 3.510000 3.690000 ;
        RECT 3.150000 1.800000 3.510000 1.890000 ;
        RECT 3.150000 1.620000 3.240000 1.800000 ;
        RECT 3.150000 3.690000 3.240000 3.870000 ;
        RECT 3.240000 1.620000 3.420000 1.800000 ;
        RECT 3.240000 3.690000 3.420000 3.870000 ;
        RECT 3.420000 1.620000 3.510000 1.800000 ;
        RECT 3.420000 3.690000 3.510000 3.870000 ;
        END
        ANTENNADIFFAREA 2.211300 ;
    END Y
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 2.070000 3.870000 2.430000 3.960000 ;
        RECT 2.070000 3.690000 2.160000 3.870000 ;
        RECT 2.070000 3.600000 2.430000 3.690000 ;
        RECT 2.160000 3.960000 2.430000 5.400000 ;
        RECT 2.160000 3.690000 2.340000 3.870000 ;
        RECT 2.340000 3.690000 2.430000 3.870000 ;
        END
        ANTENNADIFFAREA 0.615600 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 0.450000 1.890000 0.900000 1.980000 ;
        RECT 0.450000 1.620000 0.540000 1.890000 ;
        RECT 0.450000 1.530000 0.900000 1.620000 ;
        RECT 0.540000 1.620000 0.810000 1.890000 ;
        RECT 0.810000 1.620000 0.900000 1.890000 ;
        RECT 1.980000 1.530000 2.430000 1.620000 ;
        RECT 1.980000 1.890000 2.430000 1.980000 ;
        RECT 1.980000 1.620000 2.070000 1.890000 ;
        RECT 2.070000 1.620000 2.340000 1.890000 ;
        RECT 2.340000 1.620000 2.430000 1.890000 ;
        LAYER v1 ;
        RECT 0.540000 1.620000 0.810000 1.890000 ;
        RECT 2.070000 1.620000 2.340000 1.890000 ;
        LAYER m2 ;
        RECT 0.450000 1.890000 2.430000 1.980000 ;
        RECT 0.450000 1.620000 0.540000 1.890000 ;
        RECT 0.450000 1.530000 2.430000 1.620000 ;
        RECT 0.540000 1.620000 0.810000 1.890000 ;
        RECT 0.810000 1.620000 2.070000 1.890000 ;
        RECT 2.070000 1.620000 2.340000 1.890000 ;
        RECT 2.340000 1.620000 2.430000 1.890000 ;
        END
        ANTENNADIFFAREA 0.607500 ;
    END GND
    OBS
        LAYER m1 ;
        RECT 0.360000 3.960000 0.810000 4.050000 ;
        RECT 0.360000 3.690000 0.450000 3.960000 ;
        RECT 0.360000 3.600000 0.810000 3.690000 ;
        RECT 0.360000 2.970000 0.810000 3.060000 ;
        RECT 0.360000 2.700000 0.450000 2.970000 ;
        RECT 0.360000 2.610000 0.810000 2.700000 ;
        RECT 0.450000 3.690000 0.720000 3.960000 ;
        RECT 0.450000 3.060000 0.720000 3.600000 ;
        RECT 0.450000 2.700000 0.720000 2.970000 ;
        RECT 0.720000 3.690000 0.810000 3.960000 ;
        RECT 0.720000 2.700000 0.810000 2.970000 ;
        RECT 1.260000 1.530000 1.710000 1.620000 ;
        RECT 1.350000 0.810000 1.620000 1.530000 ;
        RECT 1.350000 0.720000 1.800000 0.810000 ;
        RECT 1.350000 0.450000 1.440000 0.720000 ;
        RECT 1.350000 0.360000 1.800000 0.450000 ;
        RECT 1.440000 0.450000 1.710000 0.720000 ;
        RECT 2.340000 0.720000 2.790000 0.810000 ;
        RECT 1.710000 0.450000 1.800000 0.720000 ;
        RECT 2.340000 0.360000 2.790000 0.450000 ;
        RECT 1.260000 2.970000 1.710000 3.060000 ;
        RECT 1.260000 2.700000 1.350000 2.970000 ;
        RECT 1.260000 2.610000 1.710000 2.700000 ;
        RECT 1.260000 1.890000 1.710000 1.980000 ;
        RECT 1.260000 1.620000 1.350000 1.890000 ;
        RECT 2.340000 0.450000 2.430000 0.720000 ;
        RECT 1.350000 2.700000 1.620000 2.970000 ;
        RECT 1.350000 1.980000 1.620000 2.610000 ;
        RECT 1.350000 1.620000 1.620000 1.890000 ;
        RECT 2.430000 0.450000 2.700000 0.720000 ;
        RECT 1.620000 2.700000 1.710000 2.970000 ;
        RECT 1.620000 1.620000 1.710000 1.890000 ;
        RECT 2.700000 0.450000 2.790000 0.720000 ;
        LAYER m2 ;
        RECT 0.360000 2.970000 1.710000 3.060000 ;
        RECT 0.360000 2.700000 0.450000 2.970000 ;
        RECT 0.360000 2.610000 1.710000 2.700000 ;
        RECT 0.450000 2.700000 0.720000 2.970000 ;
        RECT 0.720000 2.700000 1.350000 2.970000 ;
        RECT 1.350000 2.700000 1.620000 2.970000 ;
        RECT 1.350000 0.720000 2.790000 0.810000 ;
        RECT 1.350000 0.450000 1.440000 0.720000 ;
        RECT 1.350000 0.360000 2.790000 0.450000 ;
        RECT 1.620000 2.700000 1.710000 2.970000 ;
        RECT 1.440000 0.450000 1.710000 0.720000 ;
        RECT 1.710000 0.450000 2.430000 0.720000 ;
        RECT 2.430000 0.450000 2.700000 0.720000 ;
        RECT 2.700000 0.450000 2.790000 0.720000 ;
    END
END _0_0std_0_0cells_0_0OR2X1

MACRO _0_0std_0_0cells_0_0LATCH
    CLASS CORE ;
    FOREIGN _0_0std_0_0cells_0_0LATCH 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 8.640000 BY 7.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 2.700000 5.220000 2.970000 6.300000 ;
        RECT 2.700000 5.130000 3.060000 5.220000 ;
        RECT 2.700000 4.950000 2.790000 5.130000 ;
        RECT 2.700000 4.860000 3.060000 4.950000 ;
        RECT 2.790000 4.950000 2.970000 5.130000 ;
        RECT 2.970000 4.950000 3.060000 5.130000 ;
        END
        ANTENNAGATEAREA 0.729000 ;
    END CLK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 6.750000 2.970000 8.370000 3.060000 ;
        RECT 6.750000 2.790000 6.840000 2.970000 ;
        RECT 6.750000 2.700000 7.110000 2.790000 ;
        RECT 6.840000 2.790000 7.020000 2.970000 ;
        RECT 7.020000 2.790000 8.370000 2.970000 ;
        END
        ANTENNAGATEAREA 0.486000 ;
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 4.770000 0.810000 6.300000 ;
        RECT 0.540000 4.680000 0.990000 4.770000 ;
        RECT 0.540000 4.410000 0.630000 4.680000 ;
        RECT 0.540000 4.320000 0.990000 4.410000 ;
        RECT 0.540000 1.980000 0.810000 4.320000 ;
        RECT 0.540000 1.890000 0.900000 1.980000 ;
        RECT 0.540000 1.710000 0.630000 1.890000 ;
        RECT 0.540000 1.620000 0.900000 1.710000 ;
        RECT 0.630000 4.500000 0.810000 4.680000 ;
        RECT 0.630000 4.410000 0.900000 4.500000 ;
        RECT 0.630000 1.710000 0.810000 1.890000 ;
        RECT 0.810000 4.500000 0.900000 4.680000 ;
        RECT 0.900000 4.410000 0.990000 4.680000 ;
        RECT 0.810000 1.710000 0.900000 1.890000 ;
        RECT 5.670000 4.770000 6.120000 4.860000 ;
        RECT 5.670000 4.680000 5.850000 4.770000 ;
        RECT 5.670000 4.410000 5.760000 4.680000 ;
        RECT 5.670000 4.320000 6.120000 4.410000 ;
        RECT 5.850000 4.680000 6.030000 4.770000 ;
        RECT 5.760000 4.590000 5.850000 4.680000 ;
        RECT 5.760000 4.410000 6.030000 4.590000 ;
        RECT 5.850000 4.590000 6.030000 4.680000 ;
        RECT 6.030000 4.410000 6.120000 4.770000 ;
        LAYER v1 ;
        RECT 0.630000 4.500000 0.810000 4.680000 ;
        RECT 0.630000 4.410000 0.900000 4.500000 ;
        RECT 0.810000 4.500000 0.900000 4.680000 ;
        RECT 5.760000 4.590000 5.850000 4.680000 ;
        RECT 5.760000 4.410000 6.030000 4.590000 ;
        RECT 5.850000 4.590000 6.030000 4.680000 ;
        LAYER m2 ;
        RECT 0.540000 4.680000 6.120000 4.770000 ;
        RECT 0.540000 4.410000 0.630000 4.680000 ;
        RECT 0.540000 4.320000 6.120000 4.410000 ;
        RECT 0.630000 4.500000 0.810000 4.680000 ;
        RECT 0.630000 4.410000 0.900000 4.500000 ;
        RECT 0.810000 4.500000 0.900000 4.680000 ;
        RECT 0.900000 4.410000 5.760000 4.680000 ;
        RECT 5.760000 4.590000 5.850000 4.680000 ;
        RECT 5.760000 4.410000 6.030000 4.590000 ;
        RECT 5.850000 4.590000 6.030000 4.680000 ;
        RECT 6.030000 4.410000 6.120000 4.680000 ;
        END
        ANTENNAGATEAREA 0.324000 ;
        ANTENNADIFFAREA 1.215000 ;
    END Q
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 1.260000 5.580000 1.710000 5.670000 ;
        RECT 1.260000 5.310000 1.350000 5.580000 ;
        RECT 1.260000 5.220000 1.710000 5.310000 ;
        RECT 1.350000 5.310000 1.620000 5.580000 ;
        RECT 1.620000 5.310000 1.710000 5.580000 ;
        RECT 1.440000 4.770000 1.710000 5.220000 ;
        RECT 1.440000 4.680000 1.800000 4.770000 ;
        RECT 1.440000 4.500000 1.530000 4.680000 ;
        RECT 1.440000 4.410000 1.800000 4.500000 ;
        RECT 1.530000 4.500000 1.710000 4.680000 ;
        RECT 1.710000 4.500000 1.800000 4.680000 ;
        RECT 6.390000 5.580000 6.840000 5.670000 ;
        RECT 6.390000 5.310000 6.480000 5.580000 ;
        RECT 6.390000 5.220000 6.840000 5.310000 ;
        RECT 6.480000 5.310000 6.750000 5.580000 ;
        RECT 6.750000 5.310000 6.840000 5.580000 ;
        RECT 6.480000 5.130000 6.840000 5.220000 ;
        RECT 6.480000 4.950000 6.570000 5.130000 ;
        RECT 6.480000 4.860000 6.840000 4.950000 ;
        RECT 6.570000 4.950000 6.750000 5.130000 ;
        RECT 6.750000 4.950000 6.840000 5.130000 ;
        LAYER v1 ;
        RECT 1.350000 5.310000 1.620000 5.580000 ;
        RECT 6.480000 5.310000 6.750000 5.580000 ;
        LAYER m2 ;
        RECT 1.260000 5.580000 6.840000 5.670000 ;
        RECT 1.260000 5.310000 1.350000 5.580000 ;
        RECT 1.260000 5.220000 6.840000 5.310000 ;
        RECT 1.350000 5.310000 1.620000 5.580000 ;
        RECT 1.620000 5.310000 6.480000 5.580000 ;
        RECT 6.480000 5.310000 6.750000 5.580000 ;
        RECT 6.750000 5.310000 6.840000 5.580000 ;
        END
        ANTENNADIFFAREA 1.701000 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 1.440000 1.350000 1.800000 1.440000 ;
        RECT 1.440000 1.170000 1.530000 1.350000 ;
        RECT 1.440000 1.080000 1.890000 1.170000 ;
        RECT 1.440000 0.810000 1.530000 1.080000 ;
        RECT 1.440000 0.720000 1.890000 0.810000 ;
        RECT 1.530000 1.170000 1.710000 1.350000 ;
        RECT 1.530000 0.810000 1.800000 1.080000 ;
        RECT 1.710000 1.170000 1.800000 1.350000 ;
        RECT 1.800000 0.810000 1.890000 1.080000 ;
        RECT 6.030000 1.080000 6.480000 1.170000 ;
        RECT 6.030000 0.810000 6.120000 1.080000 ;
        RECT 6.030000 0.720000 6.480000 0.810000 ;
        RECT 6.120000 0.810000 6.390000 1.080000 ;
        RECT 6.390000 0.810000 6.480000 1.080000 ;
        RECT 6.120000 1.350000 6.480000 1.440000 ;
        RECT 6.120000 1.170000 6.210000 1.350000 ;
        RECT 6.210000 1.170000 6.390000 1.350000 ;
        RECT 6.390000 1.170000 6.480000 1.350000 ;
        LAYER v1 ;
        RECT 1.530000 0.810000 1.800000 1.080000 ;
        RECT 6.120000 0.810000 6.390000 1.080000 ;
        LAYER m2 ;
        RECT 1.440000 1.080000 6.480000 1.170000 ;
        RECT 1.440000 0.810000 1.530000 1.080000 ;
        RECT 1.440000 0.720000 6.480000 0.810000 ;
        RECT 1.530000 0.810000 1.800000 1.080000 ;
        RECT 1.800000 0.810000 6.120000 1.080000 ;
        RECT 6.120000 0.810000 6.390000 1.080000 ;
        RECT 6.390000 0.810000 6.480000 1.080000 ;
        END
        ANTENNADIFFAREA 1.134000 ;
    END GND
    OBS
        LAYER m1 ;
        RECT 0.810000 0.450000 1.170000 0.540000 ;
        RECT 0.810000 0.270000 0.900000 0.450000 ;
        RECT 0.810000 0.180000 4.050000 0.270000 ;
        RECT 0.900000 0.270000 1.080000 0.450000 ;
        RECT 1.080000 0.270000 4.050000 0.450000 ;
        RECT 2.160000 1.620000 2.520000 1.710000 ;
        RECT 3.780000 1.080000 4.140000 1.170000 ;
        RECT 2.160000 3.690000 2.520000 3.780000 ;
        RECT 2.160000 3.510000 2.250000 3.690000 ;
        RECT 2.160000 3.420000 2.520000 3.510000 ;
        RECT 2.160000 1.890000 2.520000 1.980000 ;
        RECT 2.160000 1.710000 2.250000 1.890000 ;
        RECT 3.780000 0.450000 4.050000 1.080000 ;
        RECT 2.250000 3.510000 2.430000 3.690000 ;
        RECT 2.250000 2.970000 2.520000 3.420000 ;
        RECT 2.250000 2.880000 2.700000 2.970000 ;
        RECT 2.250000 2.610000 2.340000 2.880000 ;
        RECT 2.250000 2.520000 2.700000 2.610000 ;
        RECT 2.250000 1.980000 2.520000 2.520000 ;
        RECT 2.250000 1.710000 2.430000 1.890000 ;
        RECT 3.060000 1.620000 3.510000 1.710000 ;
        RECT 2.430000 3.510000 2.520000 3.690000 ;
        RECT 2.340000 2.610000 2.610000 2.880000 ;
        RECT 2.430000 1.710000 2.520000 1.890000 ;
        RECT 3.780000 1.440000 4.050000 3.420000 ;
        RECT 3.780000 1.350000 4.140000 1.440000 ;
        RECT 3.780000 1.170000 3.870000 1.350000 ;
        RECT 2.610000 2.610000 2.700000 2.880000 ;
        RECT 3.870000 1.170000 4.050000 1.350000 ;
        RECT 4.320000 2.880000 4.770000 2.970000 ;
        RECT 4.320000 2.610000 4.410000 2.880000 ;
        RECT 4.320000 2.520000 4.770000 2.610000 ;
        RECT 4.680000 1.620000 5.760000 1.710000 ;
        RECT 4.050000 1.170000 4.140000 1.350000 ;
        RECT 4.410000 2.790000 4.680000 2.880000 ;
        RECT 4.410000 2.610000 4.590000 2.790000 ;
        RECT 4.590000 2.610000 4.680000 2.790000 ;
        RECT 4.680000 1.890000 5.760000 1.980000 ;
        RECT 4.680000 1.710000 4.770000 1.890000 ;
        RECT 3.060000 3.780000 3.510000 3.870000 ;
        RECT 3.060000 3.510000 3.150000 3.780000 ;
        RECT 3.060000 3.420000 3.510000 3.510000 ;
        RECT 3.060000 1.980000 3.510000 2.070000 ;
        RECT 3.060000 1.710000 3.150000 1.980000 ;
        RECT 4.680000 2.610000 4.770000 2.880000 ;
        RECT 4.770000 1.710000 4.950000 1.890000 ;
        RECT 3.150000 3.690000 3.420000 3.780000 ;
        RECT 3.150000 3.510000 3.330000 3.690000 ;
        RECT 3.150000 1.890000 3.420000 1.980000 ;
        RECT 3.150000 1.710000 3.330000 1.890000 ;
        RECT 4.950000 1.710000 5.490000 1.890000 ;
        RECT 3.330000 3.510000 3.420000 3.690000 ;
        RECT 3.780000 3.420000 4.140000 3.510000 ;
        RECT 3.330000 1.710000 3.420000 1.890000 ;
        RECT 5.310000 3.780000 5.760000 3.870000 ;
        RECT 5.310000 3.510000 5.400000 3.780000 ;
        RECT 5.310000 3.420000 5.760000 3.510000 ;
        RECT 5.490000 1.710000 5.670000 1.890000 ;
        RECT 6.930000 1.620000 7.380000 1.710000 ;
        RECT 3.420000 3.510000 3.510000 3.780000 ;
        RECT 3.420000 1.710000 3.510000 1.980000 ;
        RECT 5.400000 3.690000 5.670000 3.780000 ;
        RECT 5.400000 3.510000 5.490000 3.690000 ;
        RECT 5.670000 1.710000 5.760000 1.890000 ;
        RECT 5.490000 3.510000 5.670000 3.690000 ;
        RECT 3.780000 3.690000 4.140000 3.780000 ;
        RECT 3.780000 3.510000 3.870000 3.690000 ;
        RECT 5.670000 3.510000 5.760000 3.780000 ;
        RECT 3.870000 3.510000 4.050000 3.690000 ;
        RECT 4.680000 5.130000 5.040000 5.220000 ;
        RECT 4.680000 4.950000 4.770000 5.130000 ;
        RECT 4.680000 4.860000 5.040000 4.950000 ;
        RECT 4.050000 3.510000 4.140000 3.690000 ;
        RECT 4.770000 5.940000 7.380000 6.210000 ;
        RECT 4.770000 5.220000 5.040000 5.940000 ;
        RECT 4.770000 4.950000 4.950000 5.130000 ;
        RECT 7.110000 5.220000 7.380000 5.940000 ;
        RECT 4.950000 4.950000 5.040000 5.130000 ;
        RECT 6.930000 1.980000 7.380000 2.070000 ;
        RECT 6.930000 1.710000 7.020000 1.980000 ;
        RECT 7.110000 5.130000 7.470000 5.220000 ;
        RECT 7.110000 4.860000 7.470000 4.950000 ;
        RECT 7.020000 1.890000 7.290000 1.980000 ;
        RECT 7.020000 1.710000 7.110000 1.890000 ;
        RECT 7.110000 1.710000 7.290000 1.890000 ;
        RECT 7.110000 4.950000 7.200000 5.130000 ;
        RECT 7.290000 1.710000 7.380000 1.980000 ;
        RECT 7.200000 4.950000 7.380000 5.130000 ;
        RECT 7.380000 4.950000 7.470000 5.130000 ;
        LAYER m2 ;
        RECT 2.250000 2.880000 4.770000 2.970000 ;
        RECT 2.250000 2.610000 2.340000 2.880000 ;
        RECT 2.250000 2.520000 4.770000 2.610000 ;
        RECT 2.340000 2.610000 2.610000 2.880000 ;
        RECT 2.610000 2.610000 4.410000 2.880000 ;
        RECT 3.060000 1.980000 7.380000 2.070000 ;
        RECT 3.060000 1.710000 3.150000 1.980000 ;
        RECT 3.060000 1.620000 7.380000 1.710000 ;
        RECT 3.060000 3.780000 5.760000 3.870000 ;
        RECT 3.060000 3.510000 3.150000 3.780000 ;
        RECT 3.060000 3.420000 5.760000 3.510000 ;
        RECT 4.410000 2.790000 4.680000 2.880000 ;
        RECT 4.410000 2.610000 4.590000 2.790000 ;
        RECT 3.150000 1.890000 3.420000 1.980000 ;
        RECT 3.150000 1.710000 3.330000 1.890000 ;
        RECT 3.150000 3.690000 3.420000 3.780000 ;
        RECT 3.150000 3.510000 3.330000 3.690000 ;
        RECT 4.590000 2.610000 4.680000 2.790000 ;
        RECT 3.330000 1.710000 3.420000 1.890000 ;
        RECT 3.330000 3.510000 3.420000 3.690000 ;
        RECT 4.680000 2.610000 4.770000 2.880000 ;
        RECT 3.420000 1.710000 7.020000 1.980000 ;
        RECT 3.420000 3.510000 5.400000 3.780000 ;
        RECT 7.020000 1.890000 7.290000 1.980000 ;
        RECT 7.020000 1.710000 7.110000 1.890000 ;
        RECT 5.400000 3.690000 5.670000 3.780000 ;
        RECT 5.400000 3.510000 5.490000 3.690000 ;
        RECT 7.110000 1.710000 7.290000 1.890000 ;
        RECT 5.490000 3.510000 5.670000 3.690000 ;
        RECT 7.290000 1.710000 7.380000 1.980000 ;
        RECT 5.670000 3.510000 5.760000 3.780000 ;
    END
END _0_0std_0_0cells_0_0LATCH

MACRO _0_0std_0_0cells_0_0TIELOX1
    CLASS CORE ;
    FOREIGN _0_0std_0_0cells_0_0TIELOX1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.700000 BY 4.500000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 1.440000 0.990000 2.430000 1.170000 ;
        RECT 1.440000 0.630000 1.800000 0.810000 ;
        RECT 1.440000 0.810000 1.530000 0.990000 ;
        RECT 1.530000 0.810000 1.710000 0.990000 ;
        RECT 1.710000 0.900000 2.430000 0.990000 ;
        RECT 1.710000 0.810000 1.800000 0.900000 ;
        END
        ANTENNADIFFAREA 0.178200 ;
    END Y
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 0.540000 2.880000 0.810000 3.600000 ;
        RECT 0.540000 2.790000 0.900000 2.880000 ;
        RECT 0.540000 2.610000 0.630000 2.790000 ;
        RECT 0.540000 2.520000 0.900000 2.610000 ;
        RECT 0.630000 2.610000 0.810000 2.790000 ;
        RECT 0.810000 2.610000 0.900000 2.790000 ;
        END
        ANTENNADIFFAREA 0.178200 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 0.540000 1.080000 0.810000 1.170000 ;
        RECT 0.540000 0.990000 0.900000 1.080000 ;
        RECT 0.540000 0.810000 0.630000 0.990000 ;
        RECT 0.540000 0.720000 0.900000 0.810000 ;
        RECT 0.540000 0.630000 0.810000 0.720000 ;
        RECT 0.630000 0.810000 0.810000 0.990000 ;
        RECT 0.810000 0.810000 0.900000 0.990000 ;
        END
        ANTENNADIFFAREA 0.178200 ;
    END GND
    OBS
        LAYER m1 ;
        RECT 1.440000 3.510000 1.800000 3.600000 ;
        RECT 1.440000 3.330000 1.530000 3.510000 ;
        RECT 1.440000 3.240000 1.800000 3.330000 ;
        RECT 1.440000 2.880000 1.710000 3.240000 ;
        RECT 1.440000 2.790000 1.800000 2.880000 ;
        RECT 1.440000 2.520000 1.800000 2.610000 ;
        RECT 1.530000 3.330000 1.710000 3.510000 ;
        RECT 1.710000 3.330000 1.800000 3.510000 ;
        RECT 1.440000 2.610000 1.530000 2.790000 ;
        RECT 1.530000 2.610000 1.710000 2.790000 ;
        RECT 1.710000 2.610000 1.800000 2.790000 ;
    END
END _0_0std_0_0cells_0_0TIELOX1

MACRO _0_0cell_0_0g0n1n2naa_012aax0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g0n1n2naa_012aax0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 6.480000 BY 7.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 6.030000 0.810000 6.300000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 1.620000 6.030000 1.890000 6.300000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 2.700000 6.030000 2.970000 6.300000 ;
        END
    END in_52_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 0.900000 0.810000 1.170000 ;
        END
        ANTENNADIFFAREA 0.194400 ;
    END out
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 3.780000 6.030000 4.050000 6.300000 ;
        END
        ANTENNADIFFAREA 0.729000 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 4.860000 6.030000 5.130000 6.300000 ;
        END
        ANTENNADIFFAREA 0.631800 ;
    END GND
    OBS
      LAYER m1 ;
         RECT 0.540000 1.620000 5.850000 5.490000 ;
    END
END _0_0cell_0_0g0n1n2naa_012aax0

MACRO _0_0std_0_0cells_0_0TIEHIX1
    CLASS CORE ;
    FOREIGN _0_0std_0_0cells_0_0TIEHIX1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.700000 BY 4.500000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 1.440000 2.790000 1.800000 2.880000 ;
        RECT 1.440000 2.520000 2.430000 2.610000 ;
        RECT 2.160000 2.790000 2.430000 3.600000 ;
        RECT 1.440000 2.610000 1.530000 2.790000 ;
        RECT 1.530000 2.610000 1.710000 2.790000 ;
        RECT 1.710000 2.610000 2.430000 2.790000 ;
        END
        ANTENNADIFFAREA 0.178200 ;
    END Y
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 0.540000 2.880000 0.810000 3.600000 ;
        RECT 0.540000 2.790000 0.900000 2.880000 ;
        RECT 0.540000 2.610000 0.630000 2.790000 ;
        RECT 0.540000 2.520000 0.900000 2.610000 ;
        RECT 0.630000 2.610000 0.810000 2.790000 ;
        RECT 0.810000 2.610000 0.900000 2.790000 ;
        END
        ANTENNADIFFAREA 0.178200 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 0.540000 1.080000 0.810000 1.170000 ;
        RECT 0.540000 0.990000 0.900000 1.080000 ;
        RECT 0.540000 0.810000 0.630000 0.990000 ;
        RECT 0.540000 0.720000 0.900000 0.810000 ;
        RECT 0.630000 0.810000 0.810000 0.990000 ;
        RECT 0.810000 0.810000 0.900000 0.990000 ;
        END
        ANTENNADIFFAREA 0.178200 ;
    END GND
    OBS
        LAYER m1 ;
        RECT 1.440000 0.990000 1.800000 1.080000 ;
        RECT 1.440000 0.450000 1.800000 0.810000 ;
        RECT 1.440000 0.270000 1.530000 0.450000 ;
        RECT 1.440000 0.180000 1.800000 0.270000 ;
        RECT 1.530000 0.270000 1.710000 0.450000 ;
        RECT 1.440000 0.810000 1.530000 0.990000 ;
        RECT 1.710000 0.270000 1.800000 0.450000 ;
        RECT 1.530000 0.810000 1.710000 0.990000 ;
        RECT 1.710000 0.810000 1.800000 0.990000 ;
    END
END _0_0std_0_0cells_0_0TIEHIX1

MACRO _0_0cell_0_0g0n_0x1
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g0n_0x1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.160000 BY 4.500000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 3.330000 0.810000 3.600000 ;
        END
    END in_50_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 0.900000 0.810000 1.170000 ;
        END
        ANTENNADIFFAREA 0.534600 ;
    END out
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 1.080000 3.330000 1.350000 3.600000 ;
        END
        ANTENNADIFFAREA 0.291600 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 1.620000 3.330000 1.890000 3.600000 ;
        END
        ANTENNADIFFAREA 0.243000 ;
    END GND
    OBS
      LAYER m1 ;
         RECT 0.540000 1.620000 1.530000 2.790000 ;
    END
END _0_0cell_0_0g0n_0x1

MACRO _0_0cell_0_0g0n1na_01ax0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g0n1na_01ax0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 5.940000 BY 6.300000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 5.130000 0.810000 5.400000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 2.160000 5.130000 2.430000 5.400000 ;
        END
    END in_51_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 0.900000 0.810000 1.170000 ;
        END
        ANTENNADIFFAREA 0.194400 ;
    END out
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 3.780000 5.130000 4.050000 5.400000 ;
        END
        ANTENNADIFFAREA 0.534600 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 5.400000 5.130000 5.670000 5.400000 ;
        END
        ANTENNADIFFAREA 0.469800 ;
    END GND
    OBS
      LAYER m1 ;
         RECT 0.540000 1.620000 5.310000 4.590000 ;
    END
END _0_0cell_0_0g0n1na_01ax0

MACRO _0_0std_0_0cells_0_0MUX2X1
    CLASS CORE ;
    FOREIGN _0_0std_0_0cells_0_0MUX2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 8.100000 BY 8.100000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 1.080000 6.210000 1.440000 7.740000 ;
        RECT 1.080000 6.030000 1.170000 6.210000 ;
        RECT 1.080000 5.940000 1.440000 6.030000 ;
        RECT 1.170000 6.030000 1.350000 6.210000 ;
        RECT 1.350000 6.030000 1.440000 6.210000 ;
        END
        ANTENNAGATEAREA 0.405000 ;
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 5.490000 6.300000 5.760000 7.740000 ;
        RECT 5.490000 6.210000 6.210000 6.300000 ;
        RECT 5.490000 6.030000 5.670000 6.210000 ;
        RECT 5.490000 5.940000 6.210000 6.030000 ;
        RECT 5.670000 6.030000 5.850000 6.210000 ;
        RECT 5.850000 6.030000 6.210000 6.210000 ;
        END
        ANTENNAGATEAREA 0.405000 ;
    END B
    PIN S
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 2.340000 0.450000 2.700000 0.540000 ;
        RECT 2.340000 0.270000 2.430000 0.450000 ;
        RECT 2.340000 0.180000 2.700000 0.270000 ;
        RECT 2.430000 0.270000 2.610000 0.450000 ;
        RECT 2.610000 0.270000 2.700000 0.450000 ;
        RECT 4.140000 6.210000 4.590000 6.300000 ;
        RECT 4.140000 6.030000 4.230000 6.210000 ;
        RECT 4.140000 5.940000 4.500000 6.030000 ;
        RECT 4.230000 6.030000 4.410000 6.210000 ;
        RECT 4.320000 6.300000 4.590000 7.740000 ;
        RECT 4.410000 6.030000 4.590000 6.210000 ;
        END
        ANTENNAGATEAREA 0.615600 ;
    END S
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 2.700000 1.980000 2.790000 2.250000 ;
        RECT 2.700000 1.890000 3.150000 1.980000 ;
        RECT 2.700000 2.250000 3.150000 2.340000 ;
        RECT 2.790000 2.070000 2.970000 2.250000 ;
        RECT 2.790000 1.980000 3.060000 2.070000 ;
        RECT 2.970000 2.070000 3.060000 2.250000 ;
        RECT 3.060000 1.980000 3.150000 2.250000 ;
        RECT 3.510000 4.770000 3.870000 4.860000 ;
        RECT 3.510000 4.590000 3.600000 4.770000 ;
        RECT 3.600000 4.590000 3.780000 4.770000 ;
        RECT 6.030000 2.250000 6.480000 2.340000 ;
        RECT 6.030000 1.980000 6.120000 2.250000 ;
        RECT 6.030000 1.890000 6.480000 1.980000 ;
        RECT 3.780000 4.590000 6.840000 4.770000 ;
        RECT 3.510000 4.500000 7.740000 4.590000 ;
        RECT 6.120000 2.070000 6.210000 2.250000 ;
        RECT 6.120000 1.980000 6.390000 2.070000 ;
        RECT 6.840000 4.590000 7.020000 4.770000 ;
        RECT 7.380000 2.250000 7.830000 2.340000 ;
        RECT 6.210000 2.070000 6.390000 2.250000 ;
        RECT 6.390000 1.980000 6.480000 2.250000 ;
        RECT 7.380000 1.890000 7.830000 1.980000 ;
        RECT 7.020000 4.590000 7.740000 4.770000 ;
        RECT 7.470000 2.340000 7.740000 4.500000 ;
        RECT 7.380000 1.980000 7.470000 2.250000 ;
        RECT 7.470000 1.980000 7.740000 2.250000 ;
        RECT 7.740000 1.980000 7.830000 2.250000 ;
        RECT 6.750000 4.770000 7.110000 4.860000 ;
        LAYER v1 ;
        RECT 2.790000 2.070000 2.970000 2.250000 ;
        RECT 2.790000 1.980000 3.060000 2.070000 ;
        RECT 2.970000 2.070000 3.060000 2.250000 ;
        RECT 6.120000 2.070000 6.210000 2.250000 ;
        RECT 6.120000 1.980000 6.390000 2.070000 ;
        RECT 6.210000 2.070000 6.390000 2.250000 ;
        RECT 7.470000 1.980000 7.740000 2.250000 ;
        LAYER m2 ;
        RECT 2.700000 2.250000 7.830000 2.340000 ;
        RECT 2.700000 1.980000 2.790000 2.250000 ;
        RECT 2.700000 1.890000 7.830000 1.980000 ;
        RECT 2.790000 2.070000 2.970000 2.250000 ;
        RECT 2.790000 1.980000 3.060000 2.070000 ;
        RECT 2.970000 2.070000 3.060000 2.250000 ;
        RECT 3.060000 1.980000 6.120000 2.250000 ;
        RECT 6.120000 2.070000 6.210000 2.250000 ;
        RECT 6.120000 1.980000 6.390000 2.070000 ;
        RECT 6.210000 2.070000 6.390000 2.250000 ;
        RECT 6.390000 1.980000 7.470000 2.250000 ;
        RECT 7.470000 1.980000 7.740000 2.250000 ;
        RECT 7.740000 1.980000 7.830000 2.250000 ;
        END
        ANTENNADIFFAREA 2.430000 ;
    END Y
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 1.800000 5.580000 2.250000 5.670000 ;
        RECT 1.800000 5.310000 1.890000 5.580000 ;
        RECT 1.800000 5.220000 2.250000 5.310000 ;
        RECT 1.890000 5.670000 2.160000 6.030000 ;
        RECT 1.890000 5.400000 2.070000 5.580000 ;
        RECT 1.890000 5.310000 2.160000 5.400000 ;
        RECT 2.700000 6.300000 2.970000 7.740000 ;
        RECT 1.890000 6.030000 2.970000 6.300000 ;
        RECT 2.070000 5.400000 2.160000 5.580000 ;
        RECT 2.160000 5.310000 2.250000 5.580000 ;
        RECT 5.130000 5.400000 5.580000 5.490000 ;
        RECT 5.130000 5.130000 5.220000 5.400000 ;
        RECT 5.130000 5.040000 5.580000 5.130000 ;
        RECT 5.220000 5.310000 5.490000 5.400000 ;
        RECT 5.220000 5.130000 5.400000 5.310000 ;
        RECT 5.400000 5.130000 5.490000 5.310000 ;
        RECT 5.490000 5.130000 5.580000 5.400000 ;
        LAYER v1 ;
        RECT 1.890000 5.400000 2.070000 5.580000 ;
        RECT 1.890000 5.310000 2.160000 5.400000 ;
        RECT 2.070000 5.400000 2.160000 5.580000 ;
        RECT 5.220000 5.310000 5.490000 5.400000 ;
        RECT 5.220000 5.130000 5.400000 5.310000 ;
        RECT 5.400000 5.130000 5.490000 5.310000 ;
        LAYER m2 ;
        RECT 1.800000 5.580000 5.580000 5.670000 ;
        RECT 1.800000 5.310000 1.890000 5.580000 ;
        RECT 1.800000 5.220000 5.220000 5.310000 ;
        RECT 1.890000 5.400000 2.070000 5.580000 ;
        RECT 1.890000 5.310000 2.160000 5.400000 ;
        RECT 2.070000 5.400000 2.160000 5.580000 ;
        RECT 2.160000 5.310000 5.220000 5.400000 ;
        RECT 2.160000 5.400000 5.580000 5.580000 ;
        RECT 5.220000 5.310000 5.490000 5.400000 ;
        RECT 5.130000 5.130000 5.220000 5.220000 ;
        RECT 5.130000 5.040000 5.580000 5.130000 ;
        RECT 5.220000 5.130000 5.400000 5.310000 ;
        RECT 5.400000 5.130000 5.490000 5.310000 ;
        RECT 5.490000 5.130000 5.580000 5.400000 ;
        END
        ANTENNADIFFAREA 1.344600 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 1.080000 2.250000 1.440000 2.340000 ;
        RECT 1.080000 2.070000 1.170000 2.250000 ;
        RECT 1.080000 1.980000 1.440000 2.070000 ;
        RECT 1.080000 1.350000 1.350000 1.980000 ;
        RECT 1.080000 1.260000 1.530000 1.350000 ;
        RECT 1.080000 0.990000 1.170000 1.260000 ;
        RECT 1.080000 0.900000 1.530000 0.990000 ;
        RECT 1.170000 2.070000 1.350000 2.250000 ;
        RECT 1.170000 0.990000 1.440000 1.260000 ;
        RECT 1.350000 2.070000 1.440000 2.250000 ;
        RECT 1.440000 0.990000 1.530000 1.260000 ;
        RECT 4.320000 1.260000 4.770000 1.350000 ;
        RECT 4.320000 0.990000 4.410000 1.260000 ;
        RECT 4.320000 0.900000 4.770000 0.990000 ;
        RECT 4.410000 1.350000 4.680000 2.430000 ;
        RECT 4.410000 0.990000 4.680000 1.260000 ;
        RECT 4.680000 0.990000 4.770000 1.260000 ;
        RECT 4.320000 2.520000 4.410000 2.700000 ;
        RECT 4.320000 2.430000 4.680000 2.520000 ;
        RECT 4.410000 2.520000 4.590000 2.700000 ;
        RECT 4.320000 2.700000 4.680000 2.790000 ;
        RECT 4.590000 2.520000 4.680000 2.700000 ;
        LAYER v1 ;
        RECT 1.170000 0.990000 1.440000 1.260000 ;
        RECT 4.410000 0.990000 4.680000 1.260000 ;
        LAYER m2 ;
        RECT 1.080000 1.260000 4.770000 1.350000 ;
        RECT 1.080000 0.990000 1.170000 1.260000 ;
        RECT 1.080000 0.900000 4.770000 0.990000 ;
        RECT 1.170000 0.990000 1.440000 1.260000 ;
        RECT 1.440000 0.990000 4.410000 1.260000 ;
        RECT 4.410000 0.990000 4.680000 1.260000 ;
        RECT 4.680000 0.990000 4.770000 1.260000 ;
        END
        ANTENNADIFFAREA 0.972000 ;
    END GND
    OBS
        LAYER m1 ;
        RECT 0.270000 6.930000 0.720000 7.020000 ;
        RECT 0.270000 6.660000 0.360000 6.930000 ;
        RECT 0.270000 6.570000 0.720000 6.660000 ;
        RECT 0.270000 4.680000 0.720000 4.770000 ;
        RECT 0.270000 4.410000 0.360000 4.680000 ;
        RECT 0.270000 4.320000 0.720000 4.410000 ;
        RECT 0.360000 6.660000 0.630000 6.930000 ;
        RECT 0.360000 4.410000 0.630000 4.680000 ;
        RECT 0.630000 6.660000 0.720000 6.930000 ;
        RECT 1.080000 4.680000 1.530000 4.770000 ;
        RECT 0.630000 4.410000 0.720000 4.680000 ;
        RECT 1.080000 4.320000 1.530000 4.410000 ;
        RECT 1.080000 4.410000 1.170000 4.680000 ;
        RECT 1.170000 4.590000 1.440000 4.680000 ;
        RECT 1.170000 4.410000 1.350000 4.590000 ;
        RECT 1.350000 4.410000 1.440000 4.590000 ;
        RECT 1.440000 4.410000 1.530000 4.680000 ;
        RECT 2.700000 4.590000 3.150000 4.770000 ;
        RECT 2.700000 4.410000 2.790000 4.590000 ;
        RECT 2.700000 4.140000 3.150000 4.410000 ;
        RECT 2.700000 3.870000 2.790000 4.140000 ;
        RECT 2.700000 3.780000 3.150000 3.870000 ;
        RECT 2.790000 4.410000 2.970000 4.590000 ;
        RECT 2.790000 3.870000 3.060000 4.140000 ;
        RECT 2.970000 4.410000 3.150000 4.590000 ;
        RECT 3.420000 4.140000 3.870000 4.230000 ;
        RECT 3.060000 3.870000 3.150000 4.140000 ;
        RECT 3.420000 2.790000 3.870000 3.870000 ;
        RECT 3.420000 2.610000 3.510000 2.790000 ;
        RECT 3.420000 2.430000 3.870000 2.610000 ;
        RECT 3.510000 2.610000 3.690000 2.790000 ;
        RECT 3.420000 3.870000 3.510000 4.140000 ;
        RECT 3.690000 2.610000 3.870000 2.790000 ;
        RECT 3.510000 3.870000 3.780000 4.140000 ;
        RECT 3.780000 3.870000 3.870000 4.140000 ;
        RECT 5.220000 2.520000 5.580000 2.610000 ;
        RECT 5.220000 3.240000 5.670000 3.330000 ;
        RECT 5.220000 2.970000 5.310000 3.240000 ;
        RECT 5.220000 2.880000 5.670000 2.970000 ;
        RECT 5.220000 2.790000 5.580000 2.880000 ;
        RECT 5.220000 2.610000 5.310000 2.790000 ;
        RECT 5.310000 2.970000 5.580000 3.240000 ;
        RECT 5.310000 2.610000 5.490000 2.790000 ;
        RECT 6.750000 2.520000 7.110000 2.610000 ;
        RECT 5.580000 2.970000 5.670000 3.240000 ;
        RECT 5.490000 2.610000 5.580000 2.790000 ;
        RECT 6.030000 5.580000 6.480000 5.670000 ;
        RECT 6.030000 5.310000 6.120000 5.580000 ;
        RECT 6.030000 5.220000 6.480000 5.310000 ;
        RECT 6.120000 5.310000 6.390000 5.580000 ;
        RECT 6.030000 6.930000 6.480000 7.020000 ;
        RECT 6.030000 6.660000 6.120000 6.930000 ;
        RECT 6.030000 6.570000 6.480000 6.660000 ;
        RECT 6.390000 5.310000 6.480000 5.580000 ;
        RECT 6.390000 4.140000 6.840000 4.230000 ;
        RECT 6.390000 3.870000 6.480000 4.140000 ;
        RECT 6.390000 3.780000 6.840000 3.870000 ;
        RECT 6.120000 6.660000 6.390000 6.930000 ;
        RECT 6.480000 4.050000 6.750000 4.140000 ;
        RECT 6.480000 3.870000 6.570000 4.050000 ;
        RECT 6.390000 6.660000 6.480000 6.930000 ;
        RECT 6.570000 3.870000 6.750000 4.050000 ;
        RECT 6.750000 3.240000 7.200000 3.330000 ;
        RECT 6.750000 2.970000 6.840000 3.240000 ;
        RECT 6.750000 2.880000 7.200000 2.970000 ;
        RECT 6.750000 2.790000 7.110000 2.880000 ;
        RECT 6.750000 2.610000 6.840000 2.790000 ;
        RECT 6.750000 3.870000 6.840000 4.140000 ;
        RECT 6.840000 2.970000 7.110000 3.240000 ;
        RECT 6.840000 2.610000 7.020000 2.790000 ;
        RECT 7.110000 2.970000 7.200000 3.240000 ;
        RECT 7.020000 2.610000 7.110000 2.790000 ;
        LAYER m2 ;
        RECT 0.270000 6.930000 6.480000 7.020000 ;
        RECT 0.270000 6.660000 0.360000 6.930000 ;
        RECT 0.270000 6.570000 6.480000 6.660000 ;
        RECT 0.270000 4.770000 0.720000 6.570000 ;
        RECT 0.270000 4.680000 1.530000 4.770000 ;
        RECT 0.270000 4.410000 0.360000 4.680000 ;
        RECT 0.270000 4.320000 1.530000 4.410000 ;
        RECT 0.360000 6.660000 0.630000 6.930000 ;
        RECT 0.360000 4.410000 0.630000 4.680000 ;
        RECT 0.630000 6.660000 6.120000 6.930000 ;
        RECT 0.630000 4.410000 1.170000 4.680000 ;
        RECT 6.120000 6.660000 6.390000 6.930000 ;
        RECT 1.170000 4.590000 1.440000 4.680000 ;
        RECT 1.170000 4.410000 1.350000 4.590000 ;
        RECT 6.390000 6.660000 6.480000 6.930000 ;
        RECT 6.030000 5.580000 6.480000 6.570000 ;
        RECT 1.350000 4.410000 1.440000 4.590000 ;
        RECT 1.440000 4.410000 1.530000 4.680000 ;
        RECT 2.700000 4.140000 6.840000 4.230000 ;
        RECT 2.700000 3.870000 2.790000 4.140000 ;
        RECT 2.700000 3.780000 6.840000 3.870000 ;
        RECT 2.790000 3.870000 3.060000 4.140000 ;
        RECT 3.060000 3.870000 3.510000 4.140000 ;
        RECT 3.510000 3.870000 3.780000 4.140000 ;
        RECT 3.780000 3.870000 6.480000 4.140000 ;
        RECT 5.220000 3.240000 7.200000 3.330000 ;
        RECT 5.220000 2.970000 5.310000 3.240000 ;
        RECT 5.220000 2.880000 7.200000 2.970000 ;
        RECT 6.480000 4.050000 6.750000 4.140000 ;
        RECT 6.480000 3.870000 6.570000 4.050000 ;
        RECT 5.310000 2.970000 5.580000 3.240000 ;
        RECT 6.570000 3.870000 6.750000 4.050000 ;
        RECT 5.580000 2.970000 6.840000 3.240000 ;
        RECT 6.750000 3.870000 6.840000 4.140000 ;
        RECT 6.840000 2.970000 7.110000 3.240000 ;
        RECT 7.110000 2.970000 7.200000 3.240000 ;
        RECT 6.030000 5.310000 6.120000 5.580000 ;
        RECT 6.030000 5.220000 6.480000 5.310000 ;
        RECT 6.120000 5.310000 6.390000 5.580000 ;
        RECT 6.390000 5.310000 6.480000 5.580000 ;
    END
END _0_0std_0_0cells_0_0MUX2X1

MACRO _0_0std_0_0cells_0_0NOR2X2
    CLASS CORE ;
    FOREIGN _0_0std_0_0cells_0_0NOR2X2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 4.320000 BY 9.000000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 1.440000 8.010000 1.800000 8.100000 ;
        RECT 1.440000 7.830000 1.530000 8.010000 ;
        RECT 1.440000 7.740000 1.800000 7.830000 ;
        RECT 1.530000 7.830000 1.710000 8.010000 ;
        RECT 1.710000 7.830000 1.800000 8.010000 ;
        END
        ANTENNAGATEAREA 0.648000 ;
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 2.250000 8.010000 2.610000 8.100000 ;
        RECT 2.250000 7.830000 2.340000 8.010000 ;
        RECT 2.250000 7.740000 2.610000 7.830000 ;
        RECT 2.340000 7.830000 2.520000 8.010000 ;
        RECT 2.520000 7.830000 2.610000 8.010000 ;
        END
        ANTENNAGATEAREA 0.648000 ;
    END B
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 1.890000 2.340000 1.980000 2.520000 ;
        RECT 1.890000 2.250000 2.250000 2.340000 ;
        RECT 1.800000 5.490000 2.250000 5.580000 ;
        RECT 1.980000 2.340000 2.160000 2.520000 ;
        RECT 1.890000 2.520000 2.250000 5.490000 ;
        RECT 2.160000 2.340000 2.250000 2.520000 ;
        RECT 1.800000 5.850000 2.250000 5.940000 ;
        RECT 1.800000 5.580000 1.890000 5.850000 ;
        RECT 3.150000 6.570000 3.240000 6.750000 ;
        RECT 3.150000 6.480000 3.510000 6.570000 ;
        RECT 1.890000 5.580000 2.160000 5.850000 ;
        RECT 3.240000 6.570000 3.420000 6.750000 ;
        RECT 2.160000 5.580000 2.250000 5.850000 ;
        RECT 3.420000 6.570000 3.510000 6.750000 ;
        LAYER v1 ;
        RECT 1.890000 5.580000 2.160000 5.850000 ;
        LAYER m2 ;
        RECT 1.890000 5.580000 2.160000 5.850000 ;
        RECT 2.160000 5.580000 2.250000 5.850000 ;
        END
        ANTENNADIFFAREA 5.103000 ;
    END Y
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 0.900000 5.850000 1.350000 5.940000 ;
        RECT 0.900000 5.580000 0.990000 5.850000 ;
        RECT 0.900000 5.490000 1.350000 5.580000 ;
        RECT 0.990000 5.580000 1.260000 5.850000 ;
        RECT 1.260000 5.580000 1.350000 5.850000 ;
        RECT 3.150000 6.750000 3.510000 6.840000 ;
        RECT 3.240000 6.840000 3.510000 8.010000 ;
        LAYER v1 ;
        RECT 0.990000 5.580000 1.260000 5.850000 ;
        LAYER m2 ;
        RECT 0.810000 5.850000 2.250000 5.940000 ;
        RECT 0.810000 5.580000 0.990000 5.850000 ;
        RECT 0.810000 5.400000 2.250000 5.580000 ;
        RECT 0.990000 5.580000 1.260000 5.850000 ;
        RECT 1.260000 5.580000 1.890000 5.850000 ;
        END
        ANTENNADIFFAREA 2.673000 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 0.810000 2.610000 1.170000 2.700000 ;
        RECT 0.810000 2.430000 0.900000 2.610000 ;
        RECT 0.810000 2.340000 1.170000 2.430000 ;
        RECT 0.810000 1.530000 1.080000 2.340000 ;
        RECT 0.810000 1.440000 1.260000 1.530000 ;
        RECT 0.810000 1.170000 0.900000 1.440000 ;
        RECT 0.810000 1.080000 1.260000 1.170000 ;
        RECT 0.900000 2.430000 1.080000 2.610000 ;
        RECT 0.900000 1.170000 1.170000 1.440000 ;
        RECT 1.080000 2.430000 1.170000 2.610000 ;
        RECT 1.170000 1.170000 1.260000 1.440000 ;
        RECT 3.060000 1.440000 3.510000 1.530000 ;
        RECT 3.060000 1.170000 3.150000 1.440000 ;
        RECT 3.060000 1.080000 3.510000 1.170000 ;
        RECT 3.240000 1.530000 3.510000 2.340000 ;
        RECT 3.150000 1.170000 3.420000 1.440000 ;
        RECT 3.150000 2.340000 3.510000 2.430000 ;
        RECT 3.420000 1.170000 3.510000 1.440000 ;
        RECT 3.150000 2.610000 3.510000 2.700000 ;
        RECT 3.150000 2.430000 3.240000 2.610000 ;
        RECT 3.240000 2.430000 3.420000 2.610000 ;
        RECT 3.420000 2.430000 3.510000 2.610000 ;
        LAYER v1 ;
        RECT 0.900000 1.170000 1.170000 1.440000 ;
        RECT 3.150000 1.170000 3.420000 1.440000 ;
        LAYER m2 ;
        RECT 0.810000 1.440000 3.510000 1.530000 ;
        RECT 0.810000 1.170000 0.900000 1.440000 ;
        RECT 0.810000 1.080000 3.510000 1.170000 ;
        RECT 0.900000 1.170000 1.170000 1.440000 ;
        RECT 1.170000 1.170000 3.150000 1.440000 ;
        RECT 3.150000 1.170000 3.420000 1.440000 ;
        RECT 3.420000 1.170000 3.510000 1.440000 ;
        END
        ANTENNADIFFAREA 1.944000 ;
    END GND
END _0_0std_0_0cells_0_0NOR2X2

MACRO _0_0std_0_0cells_0_0LATCHINV
    CLASS CORE ;
    FOREIGN _0_0std_0_0cells_0_0LATCHINV 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 7.560000 BY 9.000000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CLK
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 2.070000 7.110000 2.430000 8.190000 ;
        RECT 2.070000 6.930000 2.160000 7.110000 ;
        RECT 2.070000 6.840000 2.430000 6.930000 ;
        RECT 2.160000 6.930000 2.340000 7.110000 ;
        RECT 2.340000 6.930000 2.430000 7.110000 ;
        END
        ANTENNAGATEAREA 0.729000 ;
    END CLK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 7.110000 0.900000 8.190000 ;
        RECT 0.540000 6.930000 0.630000 7.110000 ;
        RECT 0.540000 6.840000 0.900000 6.930000 ;
        RECT 0.630000 6.930000 0.810000 7.110000 ;
        RECT 0.810000 6.930000 0.900000 7.110000 ;
        END
        ANTENNAGATEAREA 0.486000 ;
    END D
    PIN q
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 3.780000 7.110000 4.140000 8.190000 ;
        RECT 3.780000 6.930000 3.870000 7.110000 ;
        RECT 3.780000 6.840000 4.140000 6.930000 ;
        RECT 3.870000 6.930000 4.050000 7.110000 ;
        RECT 4.050000 6.930000 4.140000 7.110000 ;
        END
        ANTENNAGATEAREA 0.324000 ;
    END q
    PIN __q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 2.070000 3.240000 2.520000 3.330000 ;
        RECT 2.070000 2.970000 2.160000 3.240000 ;
        RECT 2.070000 2.880000 2.520000 2.970000 ;
        RECT 2.070000 2.790000 2.430000 2.880000 ;
        RECT 2.070000 2.610000 2.160000 2.790000 ;
        RECT 2.070000 2.520000 2.430000 2.610000 ;
        RECT 2.160000 2.970000 2.430000 3.240000 ;
        RECT 2.160000 2.610000 2.340000 2.790000 ;
        RECT 2.880000 5.130000 3.330000 5.220000 ;
        RECT 2.880000 4.860000 2.970000 5.130000 ;
        RECT 2.880000 4.770000 3.330000 4.860000 ;
        RECT 2.430000 2.970000 2.520000 3.240000 ;
        RECT 2.340000 2.610000 2.430000 2.790000 ;
        RECT 2.970000 4.950000 3.150000 5.130000 ;
        RECT 2.970000 4.860000 3.240000 4.950000 ;
        RECT 3.150000 4.950000 3.240000 5.130000 ;
        RECT 3.240000 4.860000 3.330000 5.130000 ;
        RECT 5.310000 2.520000 5.670000 2.610000 ;
        RECT 5.220000 3.240000 5.670000 3.330000 ;
        RECT 5.220000 2.970000 5.310000 3.240000 ;
        RECT 5.220000 2.880000 5.670000 2.970000 ;
        RECT 5.310000 2.970000 5.580000 3.240000 ;
        RECT 5.310000 2.790000 5.670000 2.880000 ;
        RECT 5.310000 2.610000 5.400000 2.790000 ;
        RECT 5.940000 3.240000 6.390000 3.330000 ;
        RECT 5.580000 2.970000 5.670000 3.240000 ;
        RECT 5.940000 2.880000 6.390000 2.970000 ;
        RECT 5.400000 2.610000 5.580000 2.790000 ;
        RECT 5.940000 5.130000 6.390000 5.220000 ;
        RECT 5.940000 4.860000 6.030000 5.130000 ;
        RECT 5.940000 4.770000 6.390000 4.860000 ;
        RECT 5.580000 2.610000 5.670000 2.790000 ;
        RECT 6.030000 4.950000 6.210000 5.130000 ;
        RECT 6.030000 4.860000 6.300000 4.950000 ;
        RECT 6.120000 4.050000 6.390000 4.770000 ;
        RECT 6.120000 3.780000 7.290000 4.050000 ;
        RECT 6.120000 3.330000 6.390000 3.780000 ;
        RECT 5.940000 2.970000 6.030000 3.240000 ;
        RECT 6.210000 4.950000 6.300000 5.130000 ;
        RECT 6.300000 4.860000 6.390000 5.130000 ;
        RECT 6.030000 2.970000 6.300000 3.240000 ;
        RECT 6.300000 2.970000 6.390000 3.240000 ;
        LAYER v1 ;
        RECT 2.160000 2.970000 2.430000 3.240000 ;
        RECT 2.970000 4.950000 3.150000 5.130000 ;
        RECT 2.970000 4.860000 3.240000 4.950000 ;
        RECT 3.150000 4.950000 3.240000 5.130000 ;
        RECT 6.030000 4.860000 6.300000 4.950000 ;
        RECT 6.030000 4.950000 6.210000 5.130000 ;
        RECT 5.310000 2.970000 5.580000 3.240000 ;
        RECT 6.210000 4.950000 6.300000 5.130000 ;
        RECT 6.030000 2.970000 6.300000 3.240000 ;
        LAYER m2 ;
        RECT 2.070000 3.240000 6.390000 3.330000 ;
        RECT 2.070000 2.970000 2.160000 3.240000 ;
        RECT 2.070000 2.880000 6.390000 2.970000 ;
        RECT 2.160000 2.970000 2.430000 3.240000 ;
        RECT 2.430000 2.970000 5.310000 3.240000 ;
        RECT 2.880000 5.130000 6.390000 5.220000 ;
        RECT 2.880000 4.860000 2.970000 5.130000 ;
        RECT 2.880000 4.770000 6.390000 4.860000 ;
        RECT 5.310000 2.970000 5.580000 3.240000 ;
        RECT 2.970000 4.950000 3.150000 5.130000 ;
        RECT 2.970000 4.860000 3.240000 4.950000 ;
        RECT 5.580000 2.970000 6.030000 3.240000 ;
        RECT 3.150000 4.950000 3.240000 5.130000 ;
        RECT 3.240000 4.860000 6.030000 5.130000 ;
        RECT 6.030000 2.970000 6.300000 3.240000 ;
        RECT 6.030000 4.950000 6.210000 5.130000 ;
        RECT 6.030000 4.860000 6.300000 4.950000 ;
        RECT 6.300000 2.970000 6.390000 3.240000 ;
        RECT 6.210000 4.950000 6.300000 5.130000 ;
        RECT 6.300000 4.860000 6.390000 5.130000 ;
        END
        ANTENNADIFFAREA 2.430000 ;
    END __q
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 1.260000 7.560000 1.710000 7.650000 ;
        RECT 1.260000 7.290000 1.350000 7.560000 ;
        RECT 1.260000 7.200000 1.710000 7.290000 ;
        RECT 1.350000 7.290000 1.620000 7.560000 ;
        RECT 1.620000 7.290000 1.710000 7.560000 ;
        RECT 1.260000 5.400000 1.620000 7.200000 ;
        RECT 1.260000 5.220000 1.350000 5.400000 ;
        RECT 1.260000 5.130000 1.620000 5.220000 ;
        RECT 1.350000 5.220000 1.530000 5.400000 ;
        RECT 1.530000 5.220000 1.620000 5.400000 ;
        RECT 4.410000 7.560000 4.860000 7.650000 ;
        RECT 4.410000 7.290000 4.500000 7.560000 ;
        RECT 4.410000 7.200000 4.860000 7.290000 ;
        RECT 4.500000 7.290000 4.770000 7.560000 ;
        RECT 5.220000 7.560000 5.670000 7.650000 ;
        RECT 4.770000 7.290000 4.860000 7.560000 ;
        RECT 5.220000 7.200000 5.670000 7.290000 ;
        RECT 5.220000 7.290000 5.310000 7.560000 ;
        RECT 5.310000 7.290000 5.580000 7.560000 ;
        RECT 4.410000 5.130000 4.770000 7.200000 ;
        RECT 4.410000 4.950000 4.500000 5.130000 ;
        RECT 4.410000 4.860000 4.770000 4.950000 ;
        RECT 5.580000 7.290000 5.670000 7.560000 ;
        RECT 4.500000 4.950000 4.680000 5.130000 ;
        RECT 4.680000 4.950000 4.770000 5.130000 ;
        RECT 5.400000 6.930000 5.670000 7.200000 ;
        LAYER v1 ;
        RECT 1.350000 7.290000 1.620000 7.560000 ;
        RECT 4.500000 7.290000 4.770000 7.560000 ;
        RECT 5.310000 7.290000 5.580000 7.560000 ;
        LAYER m2 ;
        RECT 1.260000 7.560000 5.670000 7.650000 ;
        RECT 1.260000 7.290000 1.350000 7.560000 ;
        RECT 1.260000 7.200000 5.670000 7.290000 ;
        RECT 1.350000 7.290000 1.620000 7.560000 ;
        RECT 1.620000 7.290000 4.500000 7.560000 ;
        RECT 4.500000 7.290000 4.770000 7.560000 ;
        RECT 4.770000 7.290000 5.310000 7.560000 ;
        RECT 5.310000 7.290000 5.580000 7.560000 ;
        RECT 5.580000 7.290000 5.670000 7.560000 ;
        END
        ANTENNADIFFAREA 1.377000 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 0.540000 2.250000 0.900000 2.340000 ;
        RECT 0.540000 2.070000 0.630000 2.250000 ;
        RECT 0.540000 1.530000 0.900000 2.070000 ;
        RECT 0.540000 1.440000 0.990000 1.530000 ;
        RECT 0.540000 1.170000 0.630000 1.440000 ;
        RECT 0.540000 1.080000 0.990000 1.170000 ;
        RECT 0.630000 2.070000 0.810000 2.250000 ;
        RECT 0.630000 1.170000 0.900000 1.440000 ;
        RECT 0.810000 2.070000 0.900000 2.250000 ;
        RECT 3.690000 1.530000 4.050000 2.070000 ;
        RECT 3.600000 1.440000 4.050000 1.530000 ;
        RECT 0.900000 1.170000 0.990000 1.440000 ;
        RECT 3.600000 1.080000 4.050000 1.170000 ;
        RECT 3.600000 1.170000 3.690000 1.440000 ;
        RECT 3.690000 1.170000 3.960000 1.440000 ;
        RECT 3.960000 1.170000 4.050000 1.440000 ;
        RECT 3.690000 2.250000 4.050000 2.340000 ;
        RECT 3.690000 2.070000 3.780000 2.250000 ;
        RECT 3.780000 2.070000 3.960000 2.250000 ;
        RECT 3.960000 2.070000 4.050000 2.250000 ;
        LAYER v1 ;
        RECT 0.630000 1.170000 0.900000 1.440000 ;
        RECT 3.690000 1.170000 3.960000 1.440000 ;
        LAYER m2 ;
        RECT 0.540000 1.440000 4.050000 1.530000 ;
        RECT 0.540000 1.170000 0.630000 1.440000 ;
        RECT 0.540000 1.080000 4.050000 1.170000 ;
        RECT 0.630000 1.170000 0.900000 1.440000 ;
        RECT 0.900000 1.170000 3.690000 1.440000 ;
        RECT 3.690000 1.170000 3.960000 1.440000 ;
        RECT 3.960000 1.170000 4.050000 1.440000 ;
        END
        ANTENNADIFFAREA 0.972000 ;
    END GND
    OBS
        LAYER m1 ;
        RECT 0.540000 6.030000 0.990000 6.120000 ;
        RECT 0.540000 5.760000 0.630000 6.030000 ;
        RECT 0.540000 5.670000 0.990000 5.760000 ;
        RECT 0.630000 5.850000 0.810000 6.030000 ;
        RECT 0.630000 5.760000 0.900000 5.850000 ;
        RECT 0.810000 5.850000 0.900000 6.030000 ;
        RECT 0.900000 5.760000 0.990000 6.030000 ;
        RECT 4.410000 1.980000 4.860000 2.070000 ;
        RECT 2.070000 4.590000 2.430000 4.680000 ;
        RECT 2.070000 4.410000 2.160000 4.590000 ;
        RECT 2.070000 4.230000 2.430000 4.410000 ;
        RECT 2.070000 4.140000 2.520000 4.230000 ;
        RECT 2.070000 3.870000 2.160000 4.140000 ;
        RECT 2.070000 3.780000 2.520000 3.870000 ;
        RECT 5.940000 1.980000 6.390000 2.070000 ;
        RECT 2.160000 4.410000 2.340000 4.590000 ;
        RECT 2.160000 3.870000 2.430000 4.140000 ;
        RECT 2.340000 4.410000 2.430000 4.590000 ;
        RECT 2.880000 4.140000 3.330000 4.230000 ;
        RECT 2.430000 3.870000 2.520000 4.140000 ;
        RECT 2.880000 3.780000 3.330000 3.870000 ;
        RECT 2.970000 2.520000 3.330000 2.610000 ;
        RECT 2.880000 3.870000 2.970000 4.140000 ;
        RECT 4.410000 2.340000 4.860000 2.430000 ;
        RECT 2.970000 3.870000 3.240000 4.140000 ;
        RECT 2.970000 2.790000 3.330000 3.780000 ;
        RECT 2.970000 2.610000 3.060000 2.790000 ;
        RECT 3.240000 3.870000 3.330000 4.140000 ;
        RECT 3.060000 2.610000 3.240000 2.790000 ;
        RECT 4.410000 2.070000 4.500000 2.340000 ;
        RECT 3.240000 2.610000 3.330000 2.790000 ;
        RECT 4.500000 2.250000 4.770000 2.340000 ;
        RECT 4.500000 2.070000 4.590000 2.250000 ;
        RECT 4.590000 2.070000 4.770000 2.250000 ;
        RECT 4.770000 2.070000 4.860000 2.340000 ;
        RECT 5.940000 2.340000 6.390000 2.430000 ;
        RECT 5.940000 2.070000 6.030000 2.340000 ;
        RECT 6.030000 2.250000 6.300000 2.340000 ;
        RECT 6.030000 2.070000 6.210000 2.250000 ;
        RECT 5.310000 4.140000 5.760000 4.230000 ;
        RECT 5.310000 3.870000 5.400000 4.140000 ;
        RECT 5.310000 3.780000 5.760000 3.870000 ;
        RECT 6.210000 2.070000 6.300000 2.250000 ;
        RECT 5.220000 6.030000 5.670000 6.120000 ;
        RECT 5.220000 5.760000 5.310000 6.030000 ;
        RECT 5.220000 5.670000 5.670000 5.760000 ;
        RECT 5.400000 4.050000 5.670000 4.140000 ;
        RECT 5.400000 3.870000 5.490000 4.050000 ;
        RECT 6.300000 2.070000 6.390000 2.340000 ;
        RECT 5.310000 5.850000 5.490000 6.030000 ;
        RECT 5.310000 5.760000 5.580000 5.850000 ;
        RECT 5.490000 3.870000 5.670000 4.050000 ;
        RECT 5.490000 5.850000 5.580000 6.030000 ;
        RECT 5.580000 5.760000 5.670000 6.030000 ;
        RECT 5.670000 3.870000 5.760000 4.140000 ;
        LAYER m2 ;
        RECT 0.540000 6.030000 5.670000 6.120000 ;
        RECT 0.540000 5.760000 0.630000 6.030000 ;
        RECT 0.540000 5.670000 5.670000 5.760000 ;
        RECT 0.630000 5.850000 0.810000 6.030000 ;
        RECT 0.630000 5.760000 0.900000 5.850000 ;
        RECT 0.810000 5.850000 0.900000 6.030000 ;
        RECT 0.900000 5.760000 5.310000 6.030000 ;
        RECT 4.410000 2.340000 6.390000 2.430000 ;
        RECT 4.410000 2.070000 4.500000 2.340000 ;
        RECT 4.410000 1.980000 6.390000 2.070000 ;
        RECT 5.310000 5.850000 5.490000 6.030000 ;
        RECT 5.310000 5.760000 5.580000 5.850000 ;
        RECT 4.500000 2.250000 4.770000 2.340000 ;
        RECT 4.500000 2.070000 4.590000 2.250000 ;
        RECT 5.490000 5.850000 5.580000 6.030000 ;
        RECT 5.580000 5.760000 5.670000 6.030000 ;
        RECT 2.070000 4.140000 5.760000 4.230000 ;
        RECT 2.070000 3.870000 2.160000 4.140000 ;
        RECT 2.070000 3.780000 5.760000 3.870000 ;
        RECT 4.590000 2.070000 4.770000 2.250000 ;
        RECT 2.160000 3.870000 2.430000 4.140000 ;
        RECT 4.770000 2.070000 6.030000 2.340000 ;
        RECT 2.430000 3.870000 2.970000 4.140000 ;
        RECT 6.030000 2.250000 6.300000 2.340000 ;
        RECT 6.030000 2.070000 6.210000 2.250000 ;
        RECT 2.970000 3.870000 3.240000 4.140000 ;
        RECT 6.210000 2.070000 6.300000 2.250000 ;
        RECT 3.240000 3.870000 5.400000 4.140000 ;
        RECT 6.300000 2.070000 6.390000 2.340000 ;
        RECT 5.400000 4.050000 5.670000 4.140000 ;
        RECT 5.400000 3.870000 5.490000 4.050000 ;
        RECT 5.490000 3.870000 5.670000 4.050000 ;
        RECT 5.670000 3.870000 5.760000 4.140000 ;
    END
END _0_0std_0_0cells_0_0LATCHINV

MACRO welltap_svt
    CLASS CORE WELLTAP ;
    FOREIGN welltap_svt 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.620000 BY 3.600000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 0.450000 2.430000 0.900000 2.520000 ;
        RECT 0.450000 2.160000 0.540000 2.430000 ;
        RECT 0.450000 2.070000 0.900000 2.160000 ;
        RECT 0.540000 2.340000 0.810000 2.430000 ;
        RECT 0.540000 2.160000 0.630000 2.340000 ;
        RECT 0.630000 2.160000 0.810000 2.340000 ;
        RECT 0.810000 2.160000 0.900000 2.430000 ;
        LAYER v1 ;
        RECT 0.540000 2.340000 0.810000 2.430000 ;
        RECT 0.540000 2.160000 0.630000 2.340000 ;
        RECT 0.630000 2.160000 0.810000 2.340000 ;
        LAYER m2 ;
        RECT 0.450000 2.430000 0.900000 2.970000 ;
        RECT 0.450000 2.160000 0.540000 2.430000 ;
        RECT 0.450000 2.070000 0.900000 2.160000 ;
        RECT 0.540000 2.340000 0.810000 2.430000 ;
        RECT 0.540000 2.160000 0.630000 2.340000 ;
        RECT 0.630000 2.160000 0.810000 2.340000 ;
        RECT 0.810000 2.160000 0.900000 2.430000 ;
        END
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 0.450000 1.440000 0.900000 1.530000 ;
        RECT 0.450000 1.170000 0.540000 1.440000 ;
        RECT 0.450000 1.080000 0.900000 1.170000 ;
        RECT 0.540000 1.260000 0.630000 1.440000 ;
        RECT 0.540000 1.170000 0.810000 1.260000 ;
        RECT 0.630000 1.260000 0.810000 1.440000 ;
        RECT 0.810000 1.170000 0.900000 1.440000 ;
        LAYER v1 ;
        RECT 0.540000 1.260000 0.630000 1.440000 ;
        RECT 0.540000 1.170000 0.810000 1.260000 ;
        RECT 0.630000 1.260000 0.810000 1.440000 ;
        LAYER m2 ;
        RECT 0.450000 1.440000 0.900000 1.530000 ;
        RECT 0.450000 1.170000 0.540000 1.440000 ;
        RECT 0.450000 0.630000 0.900000 1.170000 ;
        RECT 0.540000 1.260000 0.630000 1.440000 ;
        RECT 0.540000 1.170000 0.810000 1.260000 ;
        RECT 0.630000 1.260000 0.810000 1.440000 ;
        RECT 0.810000 1.170000 0.900000 1.440000 ;
        END
    END GND
END welltap_svt

MACRO circuitppnp
   CLASS CORE ;
   FOREIGN circuitppnp 0.000000 0.000000 ;
   ORIGIN 0.000000 0.000000 ; 
   SIZE 370.980000 BY 372.600000 ; 
   SYMMETRY X Y ;
   SITE CoreSite ;
END circuitppnp

MACRO circuitwell
   CLASS CORE ;
   FOREIGN circuitwell 0.000000 0.000000 ;
   ORIGIN 0.000000 0.000000 ; 
   SIZE 370.980000 BY 372.600000 ; 
   SYMMETRY X Y ;
   SITE CoreSite ;
END circuitwell

