magic
tech sky130l
timestamp 1731220337
<< m1 >>
rect 248 3335 252 3355
rect 2360 3231 2364 3263
rect 3088 3199 3092 3219
rect 3080 3063 3084 3095
rect 2024 2955 2028 2979
rect 1464 2911 1468 2931
rect 1176 2655 1180 2687
rect 2000 2515 2004 2539
rect 1216 2475 1220 2495
rect 2128 2479 2132 2499
rect 2472 2379 2476 2403
rect 1296 2343 1300 2363
rect 3184 2227 3192 2231
rect 2080 2207 2084 2227
rect 3184 2143 3188 2227
rect 928 2063 932 2099
rect 2072 2071 2076 2091
rect 2248 2071 2252 2091
rect 2880 2071 2884 2091
rect 3256 2071 3260 2111
rect 1952 1935 1956 1955
rect 2952 1823 2956 1863
rect 2448 1795 2452 1815
rect 2800 1795 2804 1815
rect 2840 1683 2844 1715
rect 944 1655 948 1675
rect 2888 1607 2892 1647
rect 392 1379 396 1399
rect 1224 1243 1228 1263
rect 1952 987 1956 1019
rect 2376 1003 2380 1019
rect 2544 963 2548 983
rect 448 827 452 847
rect 568 827 572 847
rect 1000 827 1004 863
rect 3120 719 3124 755
rect 2928 695 2932 715
rect 1240 551 1244 591
rect 1456 459 1460 539
rect 984 415 988 435
rect 792 279 796 315
rect 1160 311 1164 343
rect 896 279 900 299
rect 1080 151 1084 207
rect 1200 183 1204 207
rect 2720 155 2724 207
rect 2872 183 2876 207
<< m2c >>
rect 320 3495 324 3499
rect 488 3495 492 3499
rect 664 3495 668 3499
rect 840 3495 844 3499
rect 1008 3495 1012 3499
rect 1168 3495 1172 3499
rect 1312 3495 1316 3499
rect 1456 3495 1460 3499
rect 1600 3495 1604 3499
rect 1720 3495 1724 3499
rect 1880 3483 1884 3487
rect 2024 3483 2028 3487
rect 2192 3483 2196 3487
rect 2360 3483 2364 3487
rect 2528 3483 2532 3487
rect 2688 3483 2692 3487
rect 2848 3483 2852 3487
rect 3016 3483 3020 3487
rect 184 3375 188 3379
rect 304 3375 308 3379
rect 464 3375 468 3379
rect 624 3375 628 3379
rect 784 3375 788 3379
rect 944 3375 948 3379
rect 1112 3375 1116 3379
rect 1280 3375 1284 3379
rect 1448 3375 1452 3379
rect 2080 3367 2084 3371
rect 2200 3367 2204 3371
rect 2320 3367 2324 3371
rect 2440 3367 2444 3371
rect 2560 3367 2564 3371
rect 2672 3367 2676 3371
rect 2776 3367 2780 3371
rect 2880 3367 2884 3371
rect 2984 3367 2988 3371
rect 3088 3367 3092 3371
rect 3200 3367 3204 3371
rect 184 3355 188 3359
rect 248 3355 252 3359
rect 376 3355 380 3359
rect 584 3355 588 3359
rect 792 3355 796 3359
rect 984 3355 988 3359
rect 1168 3355 1172 3359
rect 1344 3355 1348 3359
rect 1512 3355 1516 3359
rect 1688 3355 1692 3359
rect 2208 3351 2212 3355
rect 2344 3351 2348 3355
rect 2480 3351 2484 3355
rect 2616 3351 2620 3355
rect 2752 3351 2756 3355
rect 2888 3351 2892 3355
rect 3024 3351 3028 3355
rect 3168 3351 3172 3355
rect 248 3331 252 3335
rect 2360 3263 2364 3267
rect 2136 3235 2140 3239
rect 2288 3235 2292 3239
rect 184 3231 188 3235
rect 328 3231 332 3235
rect 512 3231 516 3235
rect 696 3231 700 3235
rect 880 3231 884 3235
rect 1056 3231 1060 3235
rect 1224 3231 1228 3235
rect 1392 3231 1396 3235
rect 1552 3231 1556 3235
rect 1720 3231 1724 3235
rect 2448 3235 2452 3239
rect 2608 3235 2612 3239
rect 2768 3235 2772 3239
rect 2928 3235 2932 3239
rect 3088 3235 3092 3239
rect 3248 3235 3252 3239
rect 2360 3227 2364 3231
rect 1960 3219 1964 3223
rect 2096 3219 2100 3223
rect 2248 3219 2252 3223
rect 2408 3219 2412 3223
rect 2576 3219 2580 3223
rect 2736 3219 2740 3223
rect 2896 3219 2900 3223
rect 3056 3219 3060 3223
rect 3088 3219 3092 3223
rect 3216 3219 3220 3223
rect 3384 3219 3388 3223
rect 232 3211 236 3215
rect 376 3211 380 3215
rect 536 3211 540 3215
rect 696 3211 700 3215
rect 856 3211 860 3215
rect 1016 3211 1020 3215
rect 1184 3211 1188 3215
rect 1352 3211 1356 3215
rect 1520 3211 1524 3215
rect 3088 3195 3092 3199
rect 1880 3103 1884 3107
rect 2056 3103 2060 3107
rect 2256 3103 2260 3107
rect 2448 3103 2452 3107
rect 2632 3103 2636 3107
rect 2808 3103 2812 3107
rect 2968 3103 2972 3107
rect 3128 3103 3132 3107
rect 3280 3103 3284 3107
rect 3416 3103 3420 3107
rect 416 3095 420 3099
rect 536 3095 540 3099
rect 656 3095 660 3099
rect 776 3095 780 3099
rect 896 3095 900 3099
rect 1016 3095 1020 3099
rect 1128 3095 1132 3099
rect 1248 3095 1252 3099
rect 1368 3095 1372 3099
rect 3080 3095 3084 3099
rect 1880 3083 1884 3087
rect 2008 3083 2012 3087
rect 2168 3083 2172 3087
rect 2344 3083 2348 3087
rect 2536 3083 2540 3087
rect 2744 3083 2748 3087
rect 2968 3083 2972 3087
rect 488 3079 492 3083
rect 576 3079 580 3083
rect 664 3079 668 3083
rect 752 3079 756 3083
rect 840 3079 844 3083
rect 928 3079 932 3083
rect 1016 3079 1020 3083
rect 1104 3079 1108 3083
rect 1192 3079 1196 3083
rect 3200 3083 3204 3087
rect 3416 3083 3420 3087
rect 3080 3059 3084 3063
rect 2024 2979 2028 2983
rect 552 2955 556 2959
rect 640 2955 644 2959
rect 728 2955 732 2959
rect 816 2955 820 2959
rect 904 2955 908 2959
rect 992 2955 996 2959
rect 1080 2955 1084 2959
rect 1168 2955 1172 2959
rect 1256 2955 1260 2959
rect 1344 2955 1348 2959
rect 1880 2951 1884 2955
rect 1968 2951 1972 2955
rect 2024 2951 2028 2955
rect 2080 2951 2084 2955
rect 2192 2951 2196 2955
rect 2296 2951 2300 2955
rect 2408 2951 2412 2955
rect 2528 2951 2532 2955
rect 2672 2951 2676 2955
rect 2840 2951 2844 2955
rect 3032 2951 3036 2955
rect 3232 2951 3236 2955
rect 3416 2951 3420 2955
rect 376 2931 380 2935
rect 496 2931 500 2935
rect 624 2931 628 2935
rect 760 2931 764 2935
rect 896 2931 900 2935
rect 1024 2931 1028 2935
rect 1152 2931 1156 2935
rect 1280 2931 1284 2935
rect 1408 2931 1412 2935
rect 1464 2931 1468 2935
rect 1544 2931 1548 2935
rect 1880 2927 1884 2931
rect 2064 2927 2068 2931
rect 2264 2927 2268 2931
rect 2456 2927 2460 2931
rect 2640 2927 2644 2931
rect 2808 2927 2812 2931
rect 2960 2927 2964 2931
rect 3112 2927 3116 2931
rect 3256 2927 3260 2931
rect 3408 2927 3412 2931
rect 1464 2907 1468 2911
rect 1880 2811 1884 2815
rect 2048 2811 2052 2815
rect 2240 2811 2244 2815
rect 2432 2811 2436 2815
rect 2616 2811 2620 2815
rect 2784 2811 2788 2815
rect 2952 2811 2956 2815
rect 3112 2811 3116 2815
rect 3272 2811 3276 2815
rect 3416 2811 3420 2815
rect 184 2807 188 2811
rect 304 2807 308 2811
rect 464 2807 468 2811
rect 624 2807 628 2811
rect 784 2807 788 2811
rect 944 2807 948 2811
rect 1096 2807 1100 2811
rect 1240 2807 1244 2811
rect 1392 2807 1396 2811
rect 1544 2807 1548 2811
rect 1880 2795 1884 2799
rect 2064 2795 2068 2799
rect 2264 2795 2268 2799
rect 2456 2795 2460 2799
rect 2632 2795 2636 2799
rect 2800 2795 2804 2799
rect 2960 2795 2964 2799
rect 3120 2795 3124 2799
rect 3280 2795 3284 2799
rect 3416 2795 3420 2799
rect 184 2783 188 2787
rect 296 2783 300 2787
rect 440 2783 444 2787
rect 592 2783 596 2787
rect 744 2783 748 2787
rect 904 2783 908 2787
rect 1072 2783 1076 2787
rect 1240 2783 1244 2787
rect 1408 2783 1412 2787
rect 1576 2783 1580 2787
rect 1720 2783 1724 2787
rect 1176 2687 1180 2691
rect 296 2659 300 2663
rect 408 2659 412 2663
rect 528 2659 532 2663
rect 664 2659 668 2663
rect 808 2659 812 2663
rect 960 2659 964 2663
rect 1112 2659 1116 2663
rect 2088 2663 2092 2667
rect 2208 2663 2212 2667
rect 2328 2663 2332 2667
rect 2456 2663 2460 2667
rect 2592 2663 2596 2667
rect 2736 2663 2740 2667
rect 2896 2663 2900 2667
rect 3072 2663 3076 2667
rect 3256 2663 3260 2667
rect 3416 2663 3420 2667
rect 1264 2659 1268 2663
rect 1424 2659 1428 2663
rect 1584 2659 1588 2663
rect 1720 2659 1724 2663
rect 1176 2651 1180 2655
rect 512 2639 516 2643
rect 600 2639 604 2643
rect 688 2639 692 2643
rect 792 2639 796 2643
rect 904 2639 908 2643
rect 1032 2639 1036 2643
rect 1176 2639 1180 2643
rect 1328 2639 1332 2643
rect 1488 2639 1492 2643
rect 1656 2639 1660 2643
rect 1920 2639 1924 2643
rect 2016 2639 2020 2643
rect 2120 2639 2124 2643
rect 2232 2639 2236 2643
rect 2344 2639 2348 2643
rect 2480 2639 2484 2643
rect 2632 2639 2636 2643
rect 2808 2639 2812 2643
rect 3008 2639 3012 2643
rect 3216 2639 3220 2643
rect 3416 2639 3420 2643
rect 2000 2539 2004 2543
rect 552 2515 556 2519
rect 640 2515 644 2519
rect 728 2515 732 2519
rect 824 2515 828 2519
rect 928 2515 932 2519
rect 1040 2515 1044 2519
rect 1152 2515 1156 2519
rect 1272 2515 1276 2519
rect 1400 2515 1404 2519
rect 1528 2515 1532 2519
rect 1656 2515 1660 2519
rect 1880 2511 1884 2515
rect 1968 2511 1972 2515
rect 2000 2511 2004 2515
rect 2056 2511 2060 2515
rect 2160 2511 2164 2515
rect 2272 2511 2276 2515
rect 2392 2511 2396 2515
rect 2536 2511 2540 2515
rect 2696 2511 2700 2515
rect 2864 2511 2868 2515
rect 3048 2511 3052 2515
rect 3240 2511 3244 2515
rect 3416 2511 3420 2515
rect 2000 2499 2004 2503
rect 2088 2499 2092 2503
rect 2128 2499 2132 2503
rect 2184 2499 2188 2503
rect 2288 2499 2292 2503
rect 2416 2499 2420 2503
rect 2576 2499 2580 2503
rect 2760 2499 2764 2503
rect 2968 2499 2972 2503
rect 3192 2499 3196 2503
rect 3416 2499 3420 2503
rect 600 2495 604 2499
rect 784 2495 788 2499
rect 960 2495 964 2499
rect 1128 2495 1132 2499
rect 1216 2495 1220 2499
rect 1288 2495 1292 2499
rect 1448 2495 1452 2499
rect 1616 2495 1620 2499
rect 2128 2475 2132 2479
rect 1216 2471 1220 2475
rect 2472 2403 2476 2407
rect 464 2379 468 2383
rect 552 2379 556 2383
rect 648 2379 652 2383
rect 752 2379 756 2383
rect 856 2379 860 2383
rect 968 2379 972 2383
rect 1088 2379 1092 2383
rect 1216 2379 1220 2383
rect 1344 2379 1348 2383
rect 1472 2379 1476 2383
rect 2264 2377 2268 2381
rect 2912 2395 2916 2399
rect 2352 2375 2356 2379
rect 2440 2375 2444 2379
rect 2472 2375 2476 2379
rect 2528 2375 2532 2379
rect 2616 2375 2620 2379
rect 2704 2375 2708 2379
rect 2792 2375 2796 2379
rect 2888 2375 2892 2379
rect 2984 2375 2988 2379
rect 368 2363 372 2367
rect 480 2363 484 2367
rect 592 2363 596 2367
rect 704 2363 708 2367
rect 816 2363 820 2367
rect 928 2363 932 2367
rect 1040 2363 1044 2367
rect 1152 2363 1156 2367
rect 1264 2363 1268 2367
rect 1296 2363 1300 2367
rect 1384 2363 1388 2367
rect 2216 2363 2220 2367
rect 2312 2363 2316 2367
rect 2416 2363 2420 2367
rect 2520 2363 2524 2367
rect 2624 2363 2628 2367
rect 2736 2363 2740 2367
rect 2848 2363 2852 2367
rect 2960 2363 2964 2367
rect 3072 2363 3076 2367
rect 1296 2339 1300 2343
rect 200 2239 204 2243
rect 320 2239 324 2243
rect 440 2239 444 2243
rect 568 2239 572 2243
rect 696 2239 700 2243
rect 824 2239 828 2243
rect 944 2239 948 2243
rect 1064 2239 1068 2243
rect 1192 2239 1196 2243
rect 1320 2239 1324 2243
rect 1936 2239 1940 2243
rect 2088 2239 2092 2243
rect 2248 2239 2252 2243
rect 2424 2239 2428 2243
rect 2600 2239 2604 2243
rect 2768 2239 2772 2243
rect 2936 2239 2940 2243
rect 3104 2239 3108 2243
rect 3272 2239 3276 2243
rect 3416 2239 3420 2243
rect 1880 2227 1884 2231
rect 2016 2227 2020 2231
rect 2080 2227 2084 2231
rect 2184 2227 2188 2231
rect 2360 2227 2364 2231
rect 2536 2227 2540 2231
rect 2704 2227 2708 2231
rect 2864 2227 2868 2231
rect 3008 2227 3012 2231
rect 3152 2227 3156 2231
rect 3192 2227 3196 2231
rect 3296 2227 3300 2231
rect 3416 2227 3420 2231
rect 184 2223 188 2227
rect 296 2223 300 2227
rect 456 2223 460 2227
rect 632 2223 636 2227
rect 816 2223 820 2227
rect 1000 2223 1004 2227
rect 1184 2223 1188 2227
rect 1368 2223 1372 2227
rect 1552 2223 1556 2227
rect 1720 2223 1724 2227
rect 2080 2203 2084 2207
rect 3184 2139 3188 2143
rect 2976 2111 2980 2115
rect 3064 2111 3068 2115
rect 3152 2111 3156 2115
rect 3240 2111 3244 2115
rect 3256 2111 3260 2115
rect 3328 2111 3332 2115
rect 3416 2111 3420 2115
rect 184 2099 188 2103
rect 296 2099 300 2103
rect 440 2099 444 2103
rect 592 2099 596 2103
rect 744 2099 748 2103
rect 888 2099 892 2103
rect 928 2099 932 2103
rect 1024 2099 1028 2103
rect 1152 2099 1156 2103
rect 1280 2099 1284 2103
rect 1400 2099 1404 2103
rect 1512 2099 1516 2103
rect 1624 2099 1628 2103
rect 1720 2099 1724 2103
rect 184 2083 188 2087
rect 272 2083 276 2087
rect 392 2083 396 2087
rect 512 2083 516 2087
rect 632 2083 636 2087
rect 752 2083 756 2087
rect 872 2083 876 2087
rect 1880 2091 1884 2095
rect 2040 2091 2044 2095
rect 2072 2091 2076 2095
rect 2216 2091 2220 2095
rect 2248 2091 2252 2095
rect 2392 2091 2396 2095
rect 2552 2091 2556 2095
rect 2704 2091 2708 2095
rect 2840 2091 2844 2095
rect 2880 2091 2884 2095
rect 2968 2091 2972 2095
rect 3088 2091 3092 2095
rect 3208 2091 3212 2095
rect 984 2083 988 2087
rect 1096 2083 1100 2087
rect 1208 2083 1212 2087
rect 1328 2083 1332 2087
rect 2072 2067 2076 2071
rect 2248 2067 2252 2071
rect 2880 2067 2884 2071
rect 3320 2091 3324 2095
rect 3416 2091 3420 2095
rect 3256 2067 3260 2071
rect 928 2059 932 2063
rect 1880 1971 1884 1975
rect 2064 1971 2068 1975
rect 2272 1971 2276 1975
rect 2480 1971 2484 1975
rect 2680 1971 2684 1975
rect 2872 1971 2876 1975
rect 3056 1971 3060 1975
rect 3248 1971 3252 1975
rect 3416 1971 3420 1975
rect 184 1959 188 1963
rect 288 1959 292 1963
rect 416 1959 420 1963
rect 552 1959 556 1963
rect 688 1959 692 1963
rect 824 1959 828 1963
rect 960 1959 964 1963
rect 1096 1959 1100 1963
rect 1232 1959 1236 1963
rect 1376 1959 1380 1963
rect 1912 1955 1916 1959
rect 1952 1955 1956 1959
rect 2048 1955 2052 1959
rect 2192 1955 2196 1959
rect 2336 1955 2340 1959
rect 2480 1955 2484 1959
rect 2624 1955 2628 1959
rect 2760 1955 2764 1959
rect 2880 1955 2884 1959
rect 3000 1955 3004 1959
rect 3112 1955 3116 1959
rect 3216 1955 3220 1959
rect 3328 1955 3332 1959
rect 3416 1955 3420 1959
rect 344 1943 348 1947
rect 472 1943 476 1947
rect 608 1943 612 1947
rect 752 1943 756 1947
rect 904 1943 908 1947
rect 1056 1943 1060 1947
rect 1208 1943 1212 1947
rect 1360 1943 1364 1947
rect 1520 1943 1524 1947
rect 1952 1931 1956 1935
rect 2952 1863 2956 1867
rect 2616 1855 2620 1859
rect 2064 1835 2068 1839
rect 2160 1835 2164 1839
rect 2264 1835 2268 1839
rect 2376 1835 2380 1839
rect 2488 1835 2492 1839
rect 2592 1835 2596 1839
rect 2696 1835 2700 1839
rect 2808 1835 2812 1839
rect 2920 1835 2924 1839
rect 480 1827 484 1831
rect 624 1827 628 1831
rect 776 1827 780 1831
rect 936 1827 940 1831
rect 1096 1827 1100 1831
rect 1248 1827 1252 1831
rect 1400 1827 1404 1831
rect 1560 1827 1564 1831
rect 1720 1827 1724 1831
rect 3032 1835 3036 1839
rect 2152 1815 2156 1819
rect 2240 1815 2244 1819
rect 2328 1815 2332 1819
rect 2416 1815 2420 1819
rect 2448 1815 2452 1819
rect 2504 1815 2508 1819
rect 2592 1815 2596 1819
rect 2680 1815 2684 1819
rect 2768 1815 2772 1819
rect 2800 1815 2804 1819
rect 2856 1815 2860 1819
rect 2944 1817 2948 1821
rect 2952 1819 2956 1823
rect 560 1811 564 1815
rect 680 1811 684 1815
rect 808 1811 812 1815
rect 936 1811 940 1815
rect 1072 1811 1076 1815
rect 1200 1811 1204 1815
rect 1328 1811 1332 1815
rect 1456 1811 1460 1815
rect 1584 1811 1588 1815
rect 1720 1811 1724 1815
rect 2448 1791 2452 1795
rect 2800 1791 2804 1795
rect 2840 1715 2844 1719
rect 1024 1711 1028 1715
rect 488 1691 492 1695
rect 584 1691 588 1695
rect 688 1691 692 1695
rect 792 1691 796 1695
rect 896 1691 900 1695
rect 1000 1691 1004 1695
rect 1104 1691 1108 1695
rect 1208 1691 1212 1695
rect 1320 1691 1324 1695
rect 1432 1691 1436 1695
rect 2192 1687 2196 1691
rect 2280 1687 2284 1691
rect 2368 1687 2372 1691
rect 2456 1687 2460 1691
rect 2544 1687 2548 1691
rect 2632 1687 2636 1691
rect 2720 1687 2724 1691
rect 2808 1687 2812 1691
rect 2896 1687 2900 1691
rect 2840 1679 2844 1683
rect 448 1675 452 1679
rect 536 1675 540 1679
rect 624 1675 628 1679
rect 712 1675 716 1679
rect 808 1675 812 1679
rect 904 1675 908 1679
rect 944 1675 948 1679
rect 1000 1675 1004 1679
rect 1096 1675 1100 1679
rect 1192 1675 1196 1679
rect 2152 1671 2156 1675
rect 2240 1671 2244 1675
rect 2328 1671 2332 1675
rect 2416 1671 2420 1675
rect 2504 1671 2508 1675
rect 2592 1671 2596 1675
rect 2680 1671 2684 1675
rect 2768 1671 2772 1675
rect 2856 1671 2860 1675
rect 2944 1671 2948 1675
rect 944 1651 948 1655
rect 2888 1647 2892 1651
rect 2888 1603 2892 1607
rect 328 1555 332 1559
rect 432 1555 436 1559
rect 544 1555 548 1559
rect 656 1555 660 1559
rect 768 1555 772 1559
rect 880 1555 884 1559
rect 992 1555 996 1559
rect 1104 1555 1108 1559
rect 1216 1555 1220 1559
rect 1328 1555 1332 1559
rect 2112 1551 2116 1555
rect 2208 1551 2212 1555
rect 2304 1551 2308 1555
rect 2408 1551 2412 1555
rect 2512 1551 2516 1555
rect 2616 1551 2620 1555
rect 2720 1551 2724 1555
rect 2824 1551 2828 1555
rect 2936 1551 2940 1555
rect 1968 1539 1972 1543
rect 2088 1539 2092 1543
rect 2216 1539 2220 1543
rect 2344 1539 2348 1543
rect 2472 1539 2476 1543
rect 2600 1539 2604 1543
rect 2728 1539 2732 1543
rect 2848 1539 2852 1543
rect 2976 1539 2980 1543
rect 3104 1539 3108 1543
rect 232 1535 236 1539
rect 376 1535 380 1539
rect 520 1535 524 1539
rect 672 1535 676 1539
rect 816 1535 820 1539
rect 960 1535 964 1539
rect 1096 1535 1100 1539
rect 1224 1535 1228 1539
rect 1360 1535 1364 1539
rect 1496 1535 1500 1539
rect 1904 1435 1908 1439
rect 2664 1435 2668 1439
rect 208 1415 212 1419
rect 424 1415 428 1419
rect 632 1415 636 1419
rect 832 1415 836 1419
rect 1008 1415 1012 1419
rect 1176 1415 1180 1419
rect 1328 1415 1332 1419
rect 1480 1415 1484 1419
rect 1640 1415 1644 1419
rect 1880 1415 1884 1419
rect 2000 1415 2004 1419
rect 2160 1415 2164 1419
rect 2320 1415 2324 1419
rect 2480 1415 2484 1419
rect 2640 1415 2644 1419
rect 2784 1415 2788 1419
rect 2920 1415 2924 1419
rect 3056 1415 3060 1419
rect 3184 1415 3188 1419
rect 3312 1415 3316 1419
rect 3416 1415 3420 1419
rect 184 1399 188 1403
rect 352 1399 356 1403
rect 392 1399 396 1403
rect 544 1399 548 1403
rect 728 1399 732 1403
rect 904 1399 908 1403
rect 1064 1399 1068 1403
rect 1216 1399 1220 1403
rect 1352 1399 1356 1403
rect 1480 1399 1484 1403
rect 1608 1399 1612 1403
rect 1720 1399 1724 1403
rect 1880 1399 1884 1403
rect 2056 1399 2060 1403
rect 2248 1399 2252 1403
rect 2432 1399 2436 1403
rect 2608 1399 2612 1403
rect 2768 1399 2772 1403
rect 2912 1399 2916 1403
rect 3048 1399 3052 1403
rect 3176 1399 3180 1403
rect 3304 1399 3308 1403
rect 3416 1399 3420 1403
rect 392 1375 396 1379
rect 184 1279 188 1283
rect 296 1279 300 1283
rect 448 1279 452 1283
rect 608 1279 612 1283
rect 776 1279 780 1283
rect 944 1279 948 1283
rect 1112 1279 1116 1283
rect 1272 1279 1276 1283
rect 1424 1279 1428 1283
rect 1584 1279 1588 1283
rect 1720 1279 1724 1283
rect 1880 1275 1884 1279
rect 2016 1275 2020 1279
rect 2192 1275 2196 1279
rect 2376 1275 2380 1279
rect 2560 1275 2564 1279
rect 2736 1275 2740 1279
rect 2912 1275 2916 1279
rect 3088 1275 3092 1279
rect 3264 1275 3268 1279
rect 3416 1275 3420 1279
rect 184 1263 188 1267
rect 272 1263 276 1267
rect 368 1263 372 1267
rect 480 1263 484 1267
rect 600 1263 604 1267
rect 728 1263 732 1267
rect 872 1263 876 1267
rect 1024 1263 1028 1267
rect 1192 1263 1196 1267
rect 1224 1263 1228 1267
rect 1368 1263 1372 1267
rect 1552 1263 1556 1267
rect 1720 1263 1724 1267
rect 1880 1263 1884 1267
rect 2144 1263 2148 1267
rect 2408 1263 2412 1267
rect 2648 1263 2652 1267
rect 2856 1263 2860 1267
rect 3056 1263 3060 1267
rect 3248 1263 3252 1267
rect 3416 1263 3420 1267
rect 1224 1239 1228 1243
rect 184 1139 188 1143
rect 280 1139 284 1143
rect 408 1139 412 1143
rect 536 1139 540 1143
rect 664 1139 668 1143
rect 792 1139 796 1143
rect 920 1139 924 1143
rect 1040 1139 1044 1143
rect 1168 1139 1172 1143
rect 1296 1139 1300 1143
rect 1984 1139 1988 1143
rect 2088 1139 2092 1143
rect 2208 1139 2212 1143
rect 2336 1139 2340 1143
rect 2472 1139 2476 1143
rect 2616 1139 2620 1143
rect 2752 1139 2756 1143
rect 2888 1139 2892 1143
rect 3024 1139 3028 1143
rect 3160 1139 3164 1143
rect 3296 1139 3300 1143
rect 3416 1139 3420 1143
rect 296 1123 300 1127
rect 416 1123 420 1127
rect 544 1123 548 1127
rect 672 1123 676 1127
rect 808 1123 812 1127
rect 936 1123 940 1127
rect 1064 1123 1068 1127
rect 1192 1123 1196 1127
rect 1320 1123 1324 1127
rect 1448 1123 1452 1127
rect 1992 1121 1996 1125
rect 2112 1119 2116 1123
rect 2240 1119 2244 1123
rect 2368 1119 2372 1123
rect 2504 1119 2508 1123
rect 2648 1119 2652 1123
rect 2800 1119 2804 1123
rect 2952 1119 2956 1123
rect 3112 1119 3116 1123
rect 3272 1119 3276 1123
rect 3416 1119 3420 1123
rect 1920 1019 1924 1023
rect 1952 1019 1956 1023
rect 2328 1019 2332 1023
rect 2376 1019 2380 1023
rect 480 1003 484 1007
rect 592 1003 596 1007
rect 712 1003 716 1007
rect 840 1003 844 1007
rect 968 1003 972 1007
rect 1088 1003 1092 1007
rect 1208 1003 1212 1007
rect 1328 1003 1332 1007
rect 1456 1003 1460 1007
rect 1584 1003 1588 1007
rect 1896 999 1900 1003
rect 2032 999 2036 1003
rect 2168 999 2172 1003
rect 2304 999 2308 1003
rect 2376 999 2380 1003
rect 2440 999 2444 1003
rect 2592 999 2596 1003
rect 2752 999 2756 1003
rect 2912 999 2916 1003
rect 3080 999 3084 1003
rect 3256 999 3260 1003
rect 3416 999 3420 1003
rect 616 983 620 987
rect 728 983 732 987
rect 840 983 844 987
rect 960 983 964 987
rect 1080 983 1084 987
rect 1192 983 1196 987
rect 1304 983 1308 987
rect 1408 983 1412 987
rect 1520 983 1524 987
rect 1632 983 1636 987
rect 1720 983 1724 987
rect 1880 983 1884 987
rect 1952 983 1956 987
rect 2024 983 2028 987
rect 2184 983 2188 987
rect 2344 983 2348 987
rect 2512 983 2516 987
rect 2544 983 2548 987
rect 2680 983 2684 987
rect 2856 983 2860 987
rect 3040 983 3044 987
rect 3232 983 3236 987
rect 3416 983 3420 987
rect 2544 959 2548 963
rect 2200 887 2204 891
rect 2176 867 2180 871
rect 2264 867 2268 871
rect 2352 867 2356 871
rect 2440 867 2444 871
rect 2528 867 2532 871
rect 2616 867 2620 871
rect 2704 867 2708 871
rect 2792 867 2796 871
rect 2880 867 2884 871
rect 464 863 468 867
rect 608 863 612 867
rect 776 863 780 867
rect 960 863 964 867
rect 1000 863 1004 867
rect 1168 863 1172 867
rect 1384 863 1388 867
rect 1608 863 1612 867
rect 184 847 188 851
rect 280 847 284 851
rect 408 847 412 851
rect 448 847 452 851
rect 536 847 540 851
rect 568 847 572 851
rect 672 847 676 851
rect 800 847 804 851
rect 928 847 932 851
rect 448 823 452 827
rect 568 823 572 827
rect 1056 847 1060 851
rect 1184 847 1188 851
rect 1320 847 1324 851
rect 2208 847 2212 851
rect 2296 847 2300 851
rect 2384 847 2388 851
rect 2472 847 2476 851
rect 2576 847 2580 851
rect 2688 847 2692 851
rect 2816 847 2820 851
rect 2960 847 2964 851
rect 3112 847 3116 851
rect 3272 847 3276 851
rect 3416 847 3420 851
rect 1000 823 1004 827
rect 3120 755 3124 759
rect 184 727 188 731
rect 272 727 276 731
rect 392 727 396 731
rect 520 727 524 731
rect 656 727 660 731
rect 792 727 796 731
rect 936 727 940 731
rect 1088 727 1092 731
rect 1240 727 1244 731
rect 1400 727 1404 731
rect 2112 727 2116 731
rect 2224 727 2228 731
rect 2344 727 2348 731
rect 2472 727 2476 731
rect 2608 727 2612 731
rect 2760 727 2764 731
rect 2920 727 2924 731
rect 3088 727 3092 731
rect 3264 727 3268 731
rect 3416 727 3420 731
rect 1976 715 1980 719
rect 2120 715 2124 719
rect 2280 715 2284 719
rect 2440 715 2444 719
rect 2600 715 2604 719
rect 2752 715 2756 719
rect 2896 715 2900 719
rect 2928 715 2932 719
rect 3032 715 3036 719
rect 3120 715 3124 719
rect 3168 715 3172 719
rect 3304 715 3308 719
rect 3416 715 3420 719
rect 216 711 220 715
rect 344 711 348 715
rect 480 711 484 715
rect 624 711 628 715
rect 776 711 780 715
rect 928 711 932 715
rect 1080 711 1084 715
rect 1232 711 1236 715
rect 1392 711 1396 715
rect 1552 711 1556 715
rect 2928 691 2932 695
rect 504 591 508 595
rect 608 591 612 595
rect 728 591 732 595
rect 848 591 852 595
rect 976 591 980 595
rect 1104 591 1108 595
rect 1232 591 1236 595
rect 1240 591 1244 595
rect 1360 591 1364 595
rect 1496 591 1500 595
rect 1632 591 1636 595
rect 1880 591 1884 595
rect 2016 591 2020 595
rect 2184 591 2188 595
rect 2360 591 2364 595
rect 2536 591 2540 595
rect 2704 591 2708 595
rect 2864 591 2868 595
rect 3008 591 3012 595
rect 3152 591 3156 595
rect 3296 591 3300 595
rect 3416 591 3420 595
rect 648 571 652 575
rect 752 571 756 575
rect 864 571 868 575
rect 976 571 980 575
rect 1088 571 1092 575
rect 1200 571 1204 575
rect 1880 579 1884 583
rect 2016 579 2020 583
rect 2176 579 2180 583
rect 2336 579 2340 583
rect 2504 579 2508 583
rect 2672 579 2676 583
rect 2848 579 2852 583
rect 3032 579 3036 583
rect 3216 579 3220 583
rect 3408 579 3412 583
rect 1304 571 1308 575
rect 1408 571 1412 575
rect 1520 571 1524 575
rect 1632 571 1636 575
rect 1720 571 1724 575
rect 1240 547 1244 551
rect 1456 539 1460 543
rect 1648 475 1652 479
rect 352 455 356 459
rect 480 455 484 459
rect 616 455 620 459
rect 752 455 756 459
rect 896 455 900 459
rect 1032 455 1036 459
rect 1160 455 1164 459
rect 1280 455 1284 459
rect 1400 455 1404 459
rect 1456 455 1460 459
rect 1512 455 1516 459
rect 1624 455 1628 459
rect 1720 455 1724 459
rect 1880 447 1884 451
rect 2016 447 2020 451
rect 2176 447 2180 451
rect 2344 447 2348 451
rect 2528 447 2532 451
rect 2728 447 2732 451
rect 2936 447 2940 451
rect 3160 447 3164 451
rect 3384 447 3388 451
rect 184 435 188 439
rect 304 435 308 439
rect 464 435 468 439
rect 632 435 636 439
rect 792 435 796 439
rect 952 435 956 439
rect 984 435 988 439
rect 1096 435 1100 439
rect 1232 435 1236 439
rect 1360 435 1364 439
rect 1488 435 1492 439
rect 1616 435 1620 439
rect 1720 435 1724 439
rect 1880 435 1884 439
rect 2008 435 2012 439
rect 2160 435 2164 439
rect 2320 435 2324 439
rect 2504 435 2508 439
rect 2704 435 2708 439
rect 2920 435 2924 439
rect 3152 435 3156 439
rect 3384 435 3388 439
rect 984 411 988 415
rect 1160 343 1164 347
rect 184 315 188 319
rect 272 315 276 319
rect 392 315 396 319
rect 520 315 524 319
rect 648 315 652 319
rect 768 315 772 319
rect 792 315 796 319
rect 888 315 892 319
rect 1008 315 1012 319
rect 1128 315 1132 319
rect 312 299 316 303
rect 424 299 428 303
rect 536 299 540 303
rect 648 299 652 303
rect 760 299 764 303
rect 1256 315 1260 319
rect 1976 315 1980 319
rect 2088 315 2092 319
rect 2208 315 2212 319
rect 2336 315 2340 319
rect 2472 315 2476 319
rect 2632 315 2636 319
rect 2808 315 2812 319
rect 3000 315 3004 319
rect 3200 315 3204 319
rect 3408 315 3412 319
rect 1160 307 1164 311
rect 2272 303 2276 307
rect 2360 303 2364 307
rect 2448 303 2452 307
rect 2536 303 2540 307
rect 2624 303 2628 307
rect 2728 303 2732 307
rect 2848 303 2852 307
rect 2976 303 2980 307
rect 3120 303 3124 307
rect 3272 303 3276 307
rect 3416 303 3420 307
rect 864 299 868 303
rect 896 299 900 303
rect 968 299 972 303
rect 1072 299 1076 303
rect 1176 299 1180 303
rect 1288 299 1292 303
rect 792 275 796 279
rect 896 275 900 279
rect 1080 207 1084 211
rect 496 179 500 183
rect 584 179 588 183
rect 672 179 676 183
rect 760 179 764 183
rect 856 179 860 183
rect 952 179 956 183
rect 1048 179 1052 183
rect 1200 207 1204 211
rect 2720 207 2724 211
rect 1152 179 1156 183
rect 1200 179 1204 183
rect 1256 179 1260 183
rect 1360 179 1364 183
rect 2192 179 2196 183
rect 2312 179 2316 183
rect 2432 179 2436 183
rect 2560 179 2564 183
rect 2688 179 2692 183
rect 2872 207 2876 211
rect 2816 179 2820 183
rect 2872 179 2876 183
rect 2944 179 2948 183
rect 3064 179 3068 183
rect 3184 179 3188 183
rect 3312 179 3316 183
rect 3416 179 3420 183
rect 2720 151 2724 155
rect 1080 147 1084 151
rect 1880 143 1884 147
rect 1968 143 1972 147
rect 2056 143 2060 147
rect 2144 143 2148 147
rect 2232 143 2236 147
rect 2344 143 2348 147
rect 2456 143 2460 147
rect 2560 143 2564 147
rect 2664 143 2668 147
rect 2768 143 2772 147
rect 2864 143 2868 147
rect 2960 143 2964 147
rect 3056 143 3060 147
rect 3152 143 3156 147
rect 3240 143 3244 147
rect 3328 143 3332 147
rect 3416 143 3420 147
rect 312 139 316 143
rect 400 139 404 143
rect 488 139 492 143
rect 576 139 580 143
rect 664 139 668 143
rect 752 139 756 143
rect 840 139 844 143
rect 928 139 932 143
rect 1016 139 1020 143
rect 1104 139 1108 143
rect 1192 139 1196 143
rect 1280 139 1284 143
rect 1368 139 1372 143
rect 1456 139 1460 143
rect 1544 139 1548 143
rect 1632 139 1636 143
rect 1720 139 1724 143
<< m2 >>
rect 1342 3507 1348 3508
rect 1342 3506 1343 3507
rect 1159 3504 1343 3506
rect 1159 3502 1161 3504
rect 1342 3503 1343 3504
rect 1347 3503 1348 3507
rect 1342 3502 1348 3503
rect 1084 3500 1161 3502
rect 206 3499 212 3500
rect 206 3495 207 3499
rect 211 3498 212 3499
rect 319 3499 325 3500
rect 319 3498 320 3499
rect 211 3496 320 3498
rect 211 3495 212 3496
rect 206 3494 212 3495
rect 319 3495 320 3496
rect 324 3495 325 3499
rect 319 3494 325 3495
rect 342 3499 348 3500
rect 342 3495 343 3499
rect 347 3498 348 3499
rect 487 3499 493 3500
rect 487 3498 488 3499
rect 347 3496 488 3498
rect 347 3495 348 3496
rect 342 3494 348 3495
rect 487 3495 488 3496
rect 492 3495 493 3499
rect 487 3494 493 3495
rect 510 3499 516 3500
rect 510 3495 511 3499
rect 515 3498 516 3499
rect 663 3499 669 3500
rect 663 3498 664 3499
rect 515 3496 664 3498
rect 515 3495 516 3496
rect 510 3494 516 3495
rect 663 3495 664 3496
rect 668 3495 669 3499
rect 663 3494 669 3495
rect 686 3499 692 3500
rect 686 3495 687 3499
rect 691 3498 692 3499
rect 839 3499 845 3500
rect 839 3498 840 3499
rect 691 3496 840 3498
rect 691 3495 692 3496
rect 686 3494 692 3495
rect 839 3495 840 3496
rect 844 3495 845 3499
rect 839 3494 845 3495
rect 1007 3499 1013 3500
rect 1007 3495 1008 3499
rect 1012 3498 1013 3499
rect 1084 3498 1086 3500
rect 1167 3499 1173 3500
rect 1167 3498 1168 3499
rect 1012 3496 1086 3498
rect 1159 3496 1168 3498
rect 1012 3495 1013 3496
rect 1007 3494 1013 3495
rect 1090 3495 1096 3496
rect 1090 3491 1091 3495
rect 1095 3494 1096 3495
rect 1159 3494 1161 3496
rect 1167 3495 1168 3496
rect 1172 3495 1173 3499
rect 1167 3494 1173 3495
rect 1190 3499 1196 3500
rect 1190 3495 1191 3499
rect 1195 3498 1196 3499
rect 1311 3499 1317 3500
rect 1311 3498 1312 3499
rect 1195 3496 1312 3498
rect 1195 3495 1196 3496
rect 1190 3494 1196 3495
rect 1311 3495 1312 3496
rect 1316 3495 1317 3499
rect 1311 3494 1317 3495
rect 1334 3499 1340 3500
rect 1334 3495 1335 3499
rect 1339 3498 1340 3499
rect 1455 3499 1461 3500
rect 1455 3498 1456 3499
rect 1339 3496 1456 3498
rect 1339 3495 1340 3496
rect 1334 3494 1340 3495
rect 1455 3495 1456 3496
rect 1460 3495 1461 3499
rect 1455 3494 1461 3495
rect 1478 3499 1484 3500
rect 1478 3495 1479 3499
rect 1483 3498 1484 3499
rect 1599 3499 1605 3500
rect 1599 3498 1600 3499
rect 1483 3496 1600 3498
rect 1483 3495 1484 3496
rect 1478 3494 1484 3495
rect 1599 3495 1600 3496
rect 1604 3495 1605 3499
rect 1599 3494 1605 3495
rect 1622 3499 1628 3500
rect 1622 3495 1623 3499
rect 1627 3498 1628 3499
rect 1719 3499 1725 3500
rect 1719 3498 1720 3499
rect 1627 3496 1720 3498
rect 1627 3495 1628 3496
rect 1622 3494 1628 3495
rect 1719 3495 1720 3496
rect 1724 3495 1725 3499
rect 1719 3494 1725 3495
rect 1095 3492 1161 3494
rect 1095 3491 1096 3492
rect 1090 3490 1096 3491
rect 1879 3487 1885 3488
rect 1879 3486 1880 3487
rect 110 3484 116 3485
rect 1766 3484 1772 3485
rect 110 3480 111 3484
rect 115 3480 116 3484
rect 110 3479 116 3480
rect 134 3483 140 3484
rect 134 3479 135 3483
rect 139 3479 140 3483
rect 134 3478 140 3479
rect 270 3483 276 3484
rect 270 3479 271 3483
rect 275 3479 276 3483
rect 270 3478 276 3479
rect 438 3483 444 3484
rect 438 3479 439 3483
rect 443 3479 444 3483
rect 438 3478 444 3479
rect 614 3483 620 3484
rect 614 3479 615 3483
rect 619 3479 620 3483
rect 614 3478 620 3479
rect 790 3483 796 3484
rect 790 3479 791 3483
rect 795 3479 796 3483
rect 790 3478 796 3479
rect 958 3483 964 3484
rect 958 3479 959 3483
rect 963 3479 964 3483
rect 958 3478 964 3479
rect 1118 3483 1124 3484
rect 1118 3479 1119 3483
rect 1123 3479 1124 3483
rect 1118 3478 1124 3479
rect 1262 3483 1268 3484
rect 1262 3479 1263 3483
rect 1267 3479 1268 3483
rect 1262 3478 1268 3479
rect 1406 3483 1412 3484
rect 1406 3479 1407 3483
rect 1411 3479 1412 3483
rect 1406 3478 1412 3479
rect 1550 3483 1556 3484
rect 1550 3479 1551 3483
rect 1555 3479 1556 3483
rect 1550 3478 1556 3479
rect 1670 3483 1676 3484
rect 1670 3479 1671 3483
rect 1675 3479 1676 3483
rect 1766 3480 1767 3484
rect 1771 3480 1772 3484
rect 1766 3479 1772 3480
rect 1796 3484 1880 3486
rect 1670 3478 1676 3479
rect 206 3475 212 3476
rect 206 3471 207 3475
rect 211 3471 212 3475
rect 206 3470 212 3471
rect 342 3475 348 3476
rect 342 3471 343 3475
rect 347 3471 348 3475
rect 342 3470 348 3471
rect 510 3475 516 3476
rect 510 3471 511 3475
rect 515 3471 516 3475
rect 510 3470 516 3471
rect 686 3475 692 3476
rect 686 3471 687 3475
rect 691 3471 692 3475
rect 686 3470 692 3471
rect 782 3475 788 3476
rect 782 3471 783 3475
rect 787 3474 788 3475
rect 1090 3475 1096 3476
rect 1090 3474 1091 3475
rect 787 3472 833 3474
rect 1033 3472 1091 3474
rect 787 3471 788 3472
rect 782 3470 788 3471
rect 1090 3471 1091 3472
rect 1095 3471 1096 3475
rect 1090 3470 1096 3471
rect 1190 3475 1196 3476
rect 1190 3471 1191 3475
rect 1195 3471 1196 3475
rect 1190 3470 1196 3471
rect 1334 3475 1340 3476
rect 1334 3471 1335 3475
rect 1339 3471 1340 3475
rect 1334 3470 1340 3471
rect 1478 3475 1484 3476
rect 1478 3471 1479 3475
rect 1483 3471 1484 3475
rect 1478 3470 1484 3471
rect 1622 3475 1628 3476
rect 1622 3471 1623 3475
rect 1627 3471 1628 3475
rect 1796 3474 1798 3484
rect 1879 3483 1880 3484
rect 1884 3483 1885 3487
rect 1879 3482 1885 3483
rect 1902 3487 1908 3488
rect 1902 3483 1903 3487
rect 1907 3486 1908 3487
rect 2023 3487 2029 3488
rect 2023 3486 2024 3487
rect 1907 3484 2024 3486
rect 1907 3483 1908 3484
rect 1902 3482 1908 3483
rect 2023 3483 2024 3484
rect 2028 3483 2029 3487
rect 2023 3482 2029 3483
rect 2046 3487 2052 3488
rect 2046 3483 2047 3487
rect 2051 3486 2052 3487
rect 2191 3487 2197 3488
rect 2191 3486 2192 3487
rect 2051 3484 2192 3486
rect 2051 3483 2052 3484
rect 2046 3482 2052 3483
rect 2191 3483 2192 3484
rect 2196 3483 2197 3487
rect 2191 3482 2197 3483
rect 2214 3487 2220 3488
rect 2214 3483 2215 3487
rect 2219 3486 2220 3487
rect 2359 3487 2365 3488
rect 2359 3486 2360 3487
rect 2219 3484 2360 3486
rect 2219 3483 2220 3484
rect 2214 3482 2220 3483
rect 2359 3483 2360 3484
rect 2364 3483 2365 3487
rect 2359 3482 2365 3483
rect 2527 3487 2533 3488
rect 2527 3483 2528 3487
rect 2532 3486 2533 3487
rect 2574 3487 2580 3488
rect 2574 3486 2575 3487
rect 2532 3484 2575 3486
rect 2532 3483 2533 3484
rect 2527 3482 2533 3483
rect 2574 3483 2575 3484
rect 2579 3483 2580 3487
rect 2574 3482 2580 3483
rect 2586 3487 2592 3488
rect 2586 3483 2587 3487
rect 2591 3486 2592 3487
rect 2687 3487 2693 3488
rect 2687 3486 2688 3487
rect 2591 3484 2688 3486
rect 2591 3483 2592 3484
rect 2586 3482 2592 3483
rect 2687 3483 2688 3484
rect 2692 3483 2693 3487
rect 2687 3482 2693 3483
rect 2710 3487 2716 3488
rect 2710 3483 2711 3487
rect 2715 3486 2716 3487
rect 2847 3487 2853 3488
rect 2847 3486 2848 3487
rect 2715 3484 2848 3486
rect 2715 3483 2716 3484
rect 2710 3482 2716 3483
rect 2847 3483 2848 3484
rect 2852 3483 2853 3487
rect 2847 3482 2853 3483
rect 2870 3487 2876 3488
rect 2870 3483 2871 3487
rect 2875 3486 2876 3487
rect 3015 3487 3021 3488
rect 3015 3486 3016 3487
rect 2875 3484 3016 3486
rect 2875 3483 2876 3484
rect 2870 3482 2876 3483
rect 3015 3483 3016 3484
rect 3020 3483 3021 3487
rect 3015 3482 3021 3483
rect 1745 3472 1798 3474
rect 1806 3472 1812 3473
rect 3462 3472 3468 3473
rect 1622 3470 1628 3471
rect 1806 3468 1807 3472
rect 1811 3468 1812 3472
rect 110 3467 116 3468
rect 110 3463 111 3467
rect 115 3463 116 3467
rect 1766 3467 1772 3468
rect 1806 3467 1812 3468
rect 1830 3471 1836 3472
rect 1830 3467 1831 3471
rect 1835 3467 1836 3471
rect 110 3462 116 3463
rect 134 3464 140 3465
rect 134 3460 135 3464
rect 139 3460 140 3464
rect 134 3459 140 3460
rect 270 3464 276 3465
rect 270 3460 271 3464
rect 275 3460 276 3464
rect 270 3459 276 3460
rect 438 3464 444 3465
rect 438 3460 439 3464
rect 443 3460 444 3464
rect 438 3459 444 3460
rect 614 3464 620 3465
rect 614 3460 615 3464
rect 619 3460 620 3464
rect 614 3459 620 3460
rect 790 3464 796 3465
rect 790 3460 791 3464
rect 795 3460 796 3464
rect 790 3459 796 3460
rect 958 3464 964 3465
rect 958 3460 959 3464
rect 963 3460 964 3464
rect 958 3459 964 3460
rect 1118 3464 1124 3465
rect 1118 3460 1119 3464
rect 1123 3460 1124 3464
rect 1118 3459 1124 3460
rect 1262 3464 1268 3465
rect 1262 3460 1263 3464
rect 1267 3460 1268 3464
rect 1262 3459 1268 3460
rect 1406 3464 1412 3465
rect 1406 3460 1407 3464
rect 1411 3460 1412 3464
rect 1406 3459 1412 3460
rect 1550 3464 1556 3465
rect 1550 3460 1551 3464
rect 1555 3460 1556 3464
rect 1550 3459 1556 3460
rect 1670 3464 1676 3465
rect 1670 3460 1671 3464
rect 1675 3460 1676 3464
rect 1766 3463 1767 3467
rect 1771 3463 1772 3467
rect 1830 3466 1836 3467
rect 1974 3471 1980 3472
rect 1974 3467 1975 3471
rect 1979 3467 1980 3471
rect 1974 3466 1980 3467
rect 2142 3471 2148 3472
rect 2142 3467 2143 3471
rect 2147 3467 2148 3471
rect 2142 3466 2148 3467
rect 2310 3471 2316 3472
rect 2310 3467 2311 3471
rect 2315 3467 2316 3471
rect 2310 3466 2316 3467
rect 2478 3471 2484 3472
rect 2478 3467 2479 3471
rect 2483 3467 2484 3471
rect 2478 3466 2484 3467
rect 2638 3471 2644 3472
rect 2638 3467 2639 3471
rect 2643 3467 2644 3471
rect 2638 3466 2644 3467
rect 2798 3471 2804 3472
rect 2798 3467 2799 3471
rect 2803 3467 2804 3471
rect 2798 3466 2804 3467
rect 2966 3471 2972 3472
rect 2966 3467 2967 3471
rect 2971 3467 2972 3471
rect 3462 3468 3463 3472
rect 3467 3468 3468 3472
rect 3462 3467 3468 3468
rect 2966 3466 2972 3467
rect 1766 3462 1772 3463
rect 1902 3463 1908 3464
rect 1670 3459 1676 3460
rect 1902 3459 1903 3463
rect 1907 3459 1908 3463
rect 1902 3458 1908 3459
rect 2046 3463 2052 3464
rect 2046 3459 2047 3463
rect 2051 3459 2052 3463
rect 2046 3458 2052 3459
rect 2214 3463 2220 3464
rect 2214 3459 2215 3463
rect 2219 3459 2220 3463
rect 2214 3458 2220 3459
rect 2222 3463 2228 3464
rect 2222 3459 2223 3463
rect 2227 3462 2228 3463
rect 2586 3463 2592 3464
rect 2586 3462 2587 3463
rect 2227 3460 2353 3462
rect 2553 3460 2587 3462
rect 2227 3459 2228 3460
rect 2222 3458 2228 3459
rect 2586 3459 2587 3460
rect 2591 3459 2592 3463
rect 2586 3458 2592 3459
rect 2710 3463 2716 3464
rect 2710 3459 2711 3463
rect 2715 3459 2716 3463
rect 2710 3458 2716 3459
rect 2870 3463 2876 3464
rect 2870 3459 2871 3463
rect 2875 3459 2876 3463
rect 2870 3458 2876 3459
rect 2882 3463 2888 3464
rect 2882 3459 2883 3463
rect 2887 3462 2888 3463
rect 2887 3460 3009 3462
rect 2887 3459 2888 3460
rect 2882 3458 2888 3459
rect 1806 3455 1812 3456
rect 1806 3451 1807 3455
rect 1811 3451 1812 3455
rect 3462 3455 3468 3456
rect 1806 3450 1812 3451
rect 1830 3452 1836 3453
rect 1830 3448 1831 3452
rect 1835 3448 1836 3452
rect 1830 3447 1836 3448
rect 1974 3452 1980 3453
rect 1974 3448 1975 3452
rect 1979 3448 1980 3452
rect 1974 3447 1980 3448
rect 2142 3452 2148 3453
rect 2142 3448 2143 3452
rect 2147 3448 2148 3452
rect 2142 3447 2148 3448
rect 2310 3452 2316 3453
rect 2310 3448 2311 3452
rect 2315 3448 2316 3452
rect 2310 3447 2316 3448
rect 2478 3452 2484 3453
rect 2478 3448 2479 3452
rect 2483 3448 2484 3452
rect 2478 3447 2484 3448
rect 2638 3452 2644 3453
rect 2638 3448 2639 3452
rect 2643 3448 2644 3452
rect 2638 3447 2644 3448
rect 2798 3452 2804 3453
rect 2798 3448 2799 3452
rect 2803 3448 2804 3452
rect 2798 3447 2804 3448
rect 2966 3452 2972 3453
rect 2966 3448 2967 3452
rect 2971 3448 2972 3452
rect 3462 3451 3463 3455
rect 3467 3451 3468 3455
rect 3462 3450 3468 3451
rect 2966 3447 2972 3448
rect 186 3423 192 3424
rect 186 3419 187 3423
rect 191 3422 192 3423
rect 191 3420 498 3422
rect 191 3419 192 3420
rect 186 3418 192 3419
rect 134 3416 140 3417
rect 110 3413 116 3414
rect 110 3409 111 3413
rect 115 3409 116 3413
rect 134 3412 135 3416
rect 139 3412 140 3416
rect 134 3411 140 3412
rect 254 3416 260 3417
rect 254 3412 255 3416
rect 259 3412 260 3416
rect 254 3411 260 3412
rect 414 3416 420 3417
rect 414 3412 415 3416
rect 419 3412 420 3416
rect 414 3411 420 3412
rect 110 3408 116 3409
rect 206 3407 212 3408
rect 206 3403 207 3407
rect 211 3403 212 3407
rect 206 3402 212 3403
rect 326 3407 332 3408
rect 326 3403 327 3407
rect 331 3403 332 3407
rect 326 3402 332 3403
rect 486 3407 492 3408
rect 486 3403 487 3407
rect 491 3403 492 3407
rect 496 3406 498 3420
rect 2082 3419 2088 3420
rect 574 3416 580 3417
rect 574 3412 575 3416
rect 579 3412 580 3416
rect 574 3411 580 3412
rect 734 3416 740 3417
rect 734 3412 735 3416
rect 739 3412 740 3416
rect 734 3411 740 3412
rect 894 3416 900 3417
rect 894 3412 895 3416
rect 899 3412 900 3416
rect 894 3411 900 3412
rect 1062 3416 1068 3417
rect 1062 3412 1063 3416
rect 1067 3412 1068 3416
rect 1062 3411 1068 3412
rect 1230 3416 1236 3417
rect 1230 3412 1231 3416
rect 1235 3412 1236 3416
rect 1230 3411 1236 3412
rect 1398 3416 1404 3417
rect 1398 3412 1399 3416
rect 1403 3412 1404 3416
rect 2082 3415 2083 3419
rect 2087 3418 2088 3419
rect 2222 3419 2228 3420
rect 2222 3418 2223 3419
rect 2087 3416 2223 3418
rect 2087 3415 2088 3416
rect 2082 3414 2088 3415
rect 2222 3415 2223 3416
rect 2227 3415 2228 3419
rect 2222 3414 2228 3415
rect 1398 3411 1404 3412
rect 1766 3413 1772 3414
rect 1766 3409 1767 3413
rect 1771 3409 1772 3413
rect 1766 3408 1772 3409
rect 2030 3408 2036 3409
rect 654 3407 660 3408
rect 496 3404 617 3406
rect 486 3402 492 3403
rect 654 3403 655 3407
rect 659 3406 660 3407
rect 1022 3407 1028 3408
rect 1022 3406 1023 3407
rect 659 3404 777 3406
rect 969 3404 1023 3406
rect 659 3403 660 3404
rect 654 3402 660 3403
rect 1022 3403 1023 3404
rect 1027 3403 1028 3407
rect 1022 3402 1028 3403
rect 1134 3407 1140 3408
rect 1134 3403 1135 3407
rect 1139 3403 1140 3407
rect 1134 3402 1140 3403
rect 1302 3407 1308 3408
rect 1302 3403 1303 3407
rect 1307 3403 1308 3407
rect 1302 3402 1308 3403
rect 1342 3407 1348 3408
rect 1342 3403 1343 3407
rect 1347 3406 1348 3407
rect 1347 3404 1441 3406
rect 1806 3405 1812 3406
rect 1347 3403 1348 3404
rect 1342 3402 1348 3403
rect 1806 3401 1807 3405
rect 1811 3401 1812 3405
rect 2030 3404 2031 3408
rect 2035 3404 2036 3408
rect 2030 3403 2036 3404
rect 2150 3408 2156 3409
rect 2150 3404 2151 3408
rect 2155 3404 2156 3408
rect 2150 3403 2156 3404
rect 2270 3408 2276 3409
rect 2270 3404 2271 3408
rect 2275 3404 2276 3408
rect 2270 3403 2276 3404
rect 2390 3408 2396 3409
rect 2390 3404 2391 3408
rect 2395 3404 2396 3408
rect 2390 3403 2396 3404
rect 2510 3408 2516 3409
rect 2510 3404 2511 3408
rect 2515 3404 2516 3408
rect 2510 3403 2516 3404
rect 2622 3408 2628 3409
rect 2622 3404 2623 3408
rect 2627 3404 2628 3408
rect 2622 3403 2628 3404
rect 2726 3408 2732 3409
rect 2726 3404 2727 3408
rect 2731 3404 2732 3408
rect 2726 3403 2732 3404
rect 2830 3408 2836 3409
rect 2830 3404 2831 3408
rect 2835 3404 2836 3408
rect 2830 3403 2836 3404
rect 2934 3408 2940 3409
rect 2934 3404 2935 3408
rect 2939 3404 2940 3408
rect 2934 3403 2940 3404
rect 3038 3408 3044 3409
rect 3038 3404 3039 3408
rect 3043 3404 3044 3408
rect 3038 3403 3044 3404
rect 3150 3408 3156 3409
rect 3150 3404 3151 3408
rect 3155 3404 3156 3408
rect 3150 3403 3156 3404
rect 3462 3405 3468 3406
rect 1806 3400 1812 3401
rect 3462 3401 3463 3405
rect 3467 3401 3468 3405
rect 3462 3400 3468 3401
rect 2102 3399 2108 3400
rect 134 3397 140 3398
rect 110 3396 116 3397
rect 110 3392 111 3396
rect 115 3392 116 3396
rect 134 3393 135 3397
rect 139 3393 140 3397
rect 134 3392 140 3393
rect 254 3397 260 3398
rect 254 3393 255 3397
rect 259 3393 260 3397
rect 254 3392 260 3393
rect 414 3397 420 3398
rect 414 3393 415 3397
rect 419 3393 420 3397
rect 414 3392 420 3393
rect 574 3397 580 3398
rect 574 3393 575 3397
rect 579 3393 580 3397
rect 574 3392 580 3393
rect 734 3397 740 3398
rect 734 3393 735 3397
rect 739 3393 740 3397
rect 734 3392 740 3393
rect 894 3397 900 3398
rect 894 3393 895 3397
rect 899 3393 900 3397
rect 894 3392 900 3393
rect 1062 3397 1068 3398
rect 1062 3393 1063 3397
rect 1067 3393 1068 3397
rect 1062 3392 1068 3393
rect 1230 3397 1236 3398
rect 1230 3393 1231 3397
rect 1235 3393 1236 3397
rect 1230 3392 1236 3393
rect 1398 3397 1404 3398
rect 1398 3393 1399 3397
rect 1403 3393 1404 3397
rect 1398 3392 1404 3393
rect 1766 3396 1772 3397
rect 1766 3392 1767 3396
rect 1771 3392 1772 3396
rect 2102 3395 2103 3399
rect 2107 3395 2108 3399
rect 2102 3394 2108 3395
rect 2222 3399 2228 3400
rect 2222 3395 2223 3399
rect 2227 3395 2228 3399
rect 2222 3394 2228 3395
rect 2342 3399 2348 3400
rect 2342 3395 2343 3399
rect 2347 3395 2348 3399
rect 2342 3394 2348 3395
rect 2350 3399 2356 3400
rect 2350 3395 2351 3399
rect 2355 3398 2356 3399
rect 2574 3399 2580 3400
rect 2355 3396 2433 3398
rect 2355 3395 2356 3396
rect 2350 3394 2356 3395
rect 2574 3395 2575 3399
rect 2579 3395 2580 3399
rect 2574 3394 2580 3395
rect 2590 3399 2596 3400
rect 2590 3395 2591 3399
rect 2595 3398 2596 3399
rect 2702 3399 2708 3400
rect 2595 3396 2665 3398
rect 2595 3395 2596 3396
rect 2590 3394 2596 3395
rect 2702 3395 2703 3399
rect 2707 3398 2708 3399
rect 2902 3399 2908 3400
rect 2707 3396 2769 3398
rect 2707 3395 2708 3396
rect 2702 3394 2708 3395
rect 2902 3395 2903 3399
rect 2907 3395 2908 3399
rect 2902 3394 2908 3395
rect 3006 3399 3012 3400
rect 3006 3395 3007 3399
rect 3011 3395 3012 3399
rect 3006 3394 3012 3395
rect 3110 3399 3116 3400
rect 3110 3395 3111 3399
rect 3115 3395 3116 3399
rect 3110 3394 3116 3395
rect 3214 3399 3220 3400
rect 3214 3395 3215 3399
rect 3219 3395 3220 3399
rect 3214 3394 3220 3395
rect 110 3391 116 3392
rect 1766 3391 1772 3392
rect 2030 3389 2036 3390
rect 1806 3388 1812 3389
rect 1806 3384 1807 3388
rect 1811 3384 1812 3388
rect 2030 3385 2031 3389
rect 2035 3385 2036 3389
rect 2030 3384 2036 3385
rect 2150 3389 2156 3390
rect 2150 3385 2151 3389
rect 2155 3385 2156 3389
rect 2150 3384 2156 3385
rect 2270 3389 2276 3390
rect 2270 3385 2271 3389
rect 2275 3385 2276 3389
rect 2270 3384 2276 3385
rect 2390 3389 2396 3390
rect 2390 3385 2391 3389
rect 2395 3385 2396 3389
rect 2390 3384 2396 3385
rect 2510 3389 2516 3390
rect 2510 3385 2511 3389
rect 2515 3385 2516 3389
rect 2510 3384 2516 3385
rect 2622 3389 2628 3390
rect 2622 3385 2623 3389
rect 2627 3385 2628 3389
rect 2622 3384 2628 3385
rect 2726 3389 2732 3390
rect 2726 3385 2727 3389
rect 2731 3385 2732 3389
rect 2726 3384 2732 3385
rect 2830 3389 2836 3390
rect 2830 3385 2831 3389
rect 2835 3385 2836 3389
rect 2830 3384 2836 3385
rect 2934 3389 2940 3390
rect 2934 3385 2935 3389
rect 2939 3385 2940 3389
rect 2934 3384 2940 3385
rect 3038 3389 3044 3390
rect 3038 3385 3039 3389
rect 3043 3385 3044 3389
rect 3038 3384 3044 3385
rect 3150 3389 3156 3390
rect 3150 3385 3151 3389
rect 3155 3385 3156 3389
rect 3150 3384 3156 3385
rect 3462 3388 3468 3389
rect 3462 3384 3463 3388
rect 3467 3384 3468 3388
rect 1806 3383 1812 3384
rect 3462 3383 3468 3384
rect 183 3379 192 3380
rect 183 3375 184 3379
rect 191 3375 192 3379
rect 183 3374 192 3375
rect 206 3379 212 3380
rect 206 3375 207 3379
rect 211 3378 212 3379
rect 303 3379 309 3380
rect 303 3378 304 3379
rect 211 3376 304 3378
rect 211 3375 212 3376
rect 206 3374 212 3375
rect 303 3375 304 3376
rect 308 3375 309 3379
rect 303 3374 309 3375
rect 326 3379 332 3380
rect 326 3375 327 3379
rect 331 3378 332 3379
rect 463 3379 469 3380
rect 463 3378 464 3379
rect 331 3376 464 3378
rect 331 3375 332 3376
rect 326 3374 332 3375
rect 463 3375 464 3376
rect 468 3375 469 3379
rect 463 3374 469 3375
rect 623 3379 629 3380
rect 623 3375 624 3379
rect 628 3378 629 3379
rect 654 3379 660 3380
rect 654 3378 655 3379
rect 628 3376 655 3378
rect 628 3375 629 3376
rect 623 3374 629 3375
rect 654 3375 655 3376
rect 659 3375 660 3379
rect 654 3374 660 3375
rect 782 3379 789 3380
rect 782 3375 783 3379
rect 788 3375 789 3379
rect 782 3374 789 3375
rect 943 3379 949 3380
rect 943 3375 944 3379
rect 948 3378 949 3379
rect 1006 3379 1012 3380
rect 1006 3378 1007 3379
rect 948 3376 1007 3378
rect 948 3375 949 3376
rect 943 3374 949 3375
rect 1006 3375 1007 3376
rect 1011 3375 1012 3379
rect 1006 3374 1012 3375
rect 1022 3379 1028 3380
rect 1022 3375 1023 3379
rect 1027 3378 1028 3379
rect 1111 3379 1117 3380
rect 1111 3378 1112 3379
rect 1027 3376 1112 3378
rect 1027 3375 1028 3376
rect 1022 3374 1028 3375
rect 1111 3375 1112 3376
rect 1116 3375 1117 3379
rect 1111 3374 1117 3375
rect 1134 3379 1140 3380
rect 1134 3375 1135 3379
rect 1139 3378 1140 3379
rect 1279 3379 1285 3380
rect 1279 3378 1280 3379
rect 1139 3376 1280 3378
rect 1139 3375 1140 3376
rect 1134 3374 1140 3375
rect 1279 3375 1280 3376
rect 1284 3375 1285 3379
rect 1279 3374 1285 3375
rect 1302 3379 1308 3380
rect 1302 3375 1303 3379
rect 1307 3378 1308 3379
rect 1447 3379 1453 3380
rect 1447 3378 1448 3379
rect 1307 3376 1448 3378
rect 1307 3375 1308 3376
rect 1302 3374 1308 3375
rect 1447 3375 1448 3376
rect 1452 3375 1453 3379
rect 1447 3374 1453 3375
rect 2079 3371 2088 3372
rect 614 3367 620 3368
rect 614 3366 615 3367
rect 480 3364 615 3366
rect 183 3359 189 3360
rect 183 3355 184 3359
rect 188 3358 189 3359
rect 247 3359 253 3360
rect 247 3358 248 3359
rect 188 3356 248 3358
rect 188 3355 189 3356
rect 183 3354 189 3355
rect 247 3355 248 3356
rect 252 3355 253 3359
rect 247 3354 253 3355
rect 375 3359 381 3360
rect 375 3355 376 3359
rect 380 3358 381 3359
rect 480 3358 482 3364
rect 614 3363 615 3364
rect 619 3363 620 3367
rect 2079 3367 2080 3371
rect 2087 3367 2088 3371
rect 2079 3366 2088 3367
rect 2102 3371 2108 3372
rect 2102 3367 2103 3371
rect 2107 3370 2108 3371
rect 2199 3371 2205 3372
rect 2199 3370 2200 3371
rect 2107 3368 2200 3370
rect 2107 3367 2108 3368
rect 2102 3366 2108 3367
rect 2199 3367 2200 3368
rect 2204 3367 2205 3371
rect 2199 3366 2205 3367
rect 2222 3371 2228 3372
rect 2222 3367 2223 3371
rect 2227 3370 2228 3371
rect 2319 3371 2325 3372
rect 2319 3370 2320 3371
rect 2227 3368 2320 3370
rect 2227 3367 2228 3368
rect 2222 3366 2228 3367
rect 2319 3367 2320 3368
rect 2324 3367 2325 3371
rect 2319 3366 2325 3367
rect 2342 3371 2348 3372
rect 2342 3367 2343 3371
rect 2347 3370 2348 3371
rect 2439 3371 2445 3372
rect 2439 3370 2440 3371
rect 2347 3368 2440 3370
rect 2347 3367 2348 3368
rect 2342 3366 2348 3367
rect 2439 3367 2440 3368
rect 2444 3367 2445 3371
rect 2439 3366 2445 3367
rect 2559 3371 2565 3372
rect 2559 3367 2560 3371
rect 2564 3370 2565 3371
rect 2590 3371 2596 3372
rect 2590 3370 2591 3371
rect 2564 3368 2591 3370
rect 2564 3367 2565 3368
rect 2559 3366 2565 3367
rect 2590 3367 2591 3368
rect 2595 3367 2596 3371
rect 2590 3366 2596 3367
rect 2671 3371 2677 3372
rect 2671 3367 2672 3371
rect 2676 3370 2677 3371
rect 2702 3371 2708 3372
rect 2702 3370 2703 3371
rect 2676 3368 2703 3370
rect 2676 3367 2677 3368
rect 2671 3366 2677 3367
rect 2702 3367 2703 3368
rect 2707 3367 2708 3371
rect 2702 3366 2708 3367
rect 2774 3371 2781 3372
rect 2774 3367 2775 3371
rect 2780 3367 2781 3371
rect 2774 3366 2781 3367
rect 2879 3371 2888 3372
rect 2879 3367 2880 3371
rect 2887 3367 2888 3371
rect 2879 3366 2888 3367
rect 2902 3371 2908 3372
rect 2902 3367 2903 3371
rect 2907 3370 2908 3371
rect 2983 3371 2989 3372
rect 2983 3370 2984 3371
rect 2907 3368 2984 3370
rect 2907 3367 2908 3368
rect 2902 3366 2908 3367
rect 2983 3367 2984 3368
rect 2988 3367 2989 3371
rect 2983 3366 2989 3367
rect 3006 3371 3012 3372
rect 3006 3367 3007 3371
rect 3011 3370 3012 3371
rect 3087 3371 3093 3372
rect 3087 3370 3088 3371
rect 3011 3368 3088 3370
rect 3011 3367 3012 3368
rect 3006 3366 3012 3367
rect 3087 3367 3088 3368
rect 3092 3367 3093 3371
rect 3087 3366 3093 3367
rect 3110 3371 3116 3372
rect 3110 3367 3111 3371
rect 3115 3370 3116 3371
rect 3199 3371 3205 3372
rect 3199 3370 3200 3371
rect 3115 3368 3200 3370
rect 3115 3367 3116 3368
rect 3110 3366 3116 3367
rect 3199 3367 3200 3368
rect 3204 3367 3205 3371
rect 3199 3366 3205 3367
rect 614 3362 620 3363
rect 2350 3363 2356 3364
rect 2350 3362 2351 3363
rect 2224 3360 2351 3362
rect 380 3356 482 3358
rect 486 3359 492 3360
rect 380 3355 381 3356
rect 375 3354 381 3355
rect 486 3355 487 3359
rect 491 3358 492 3359
rect 583 3359 589 3360
rect 583 3358 584 3359
rect 491 3356 584 3358
rect 491 3355 492 3356
rect 486 3354 492 3355
rect 583 3355 584 3356
rect 588 3355 589 3359
rect 583 3354 589 3355
rect 606 3359 612 3360
rect 606 3355 607 3359
rect 611 3358 612 3359
rect 791 3359 797 3360
rect 791 3358 792 3359
rect 611 3356 792 3358
rect 611 3355 612 3356
rect 606 3354 612 3355
rect 791 3355 792 3356
rect 796 3355 797 3359
rect 791 3354 797 3355
rect 983 3359 989 3360
rect 983 3355 984 3359
rect 988 3358 989 3359
rect 1070 3359 1076 3360
rect 1070 3358 1071 3359
rect 988 3356 1071 3358
rect 988 3355 989 3356
rect 983 3354 989 3355
rect 1070 3355 1071 3356
rect 1075 3355 1076 3359
rect 1070 3354 1076 3355
rect 1167 3359 1173 3360
rect 1167 3355 1168 3359
rect 1172 3358 1173 3359
rect 1198 3359 1204 3360
rect 1198 3358 1199 3359
rect 1172 3356 1199 3358
rect 1172 3355 1173 3356
rect 1167 3354 1173 3355
rect 1198 3355 1199 3356
rect 1203 3355 1204 3359
rect 1198 3354 1204 3355
rect 1343 3359 1349 3360
rect 1343 3355 1344 3359
rect 1348 3358 1349 3359
rect 1374 3359 1380 3360
rect 1374 3358 1375 3359
rect 1348 3356 1375 3358
rect 1348 3355 1349 3356
rect 1343 3354 1349 3355
rect 1374 3355 1375 3356
rect 1379 3355 1380 3359
rect 1374 3354 1380 3355
rect 1511 3359 1517 3360
rect 1511 3355 1512 3359
rect 1516 3358 1517 3359
rect 1598 3359 1604 3360
rect 1598 3358 1599 3359
rect 1516 3356 1599 3358
rect 1516 3355 1517 3356
rect 1511 3354 1517 3355
rect 1598 3355 1599 3356
rect 1603 3355 1604 3359
rect 1598 3354 1604 3355
rect 1687 3359 1693 3360
rect 1687 3355 1688 3359
rect 1692 3358 1693 3359
rect 1734 3359 1740 3360
rect 1734 3358 1735 3359
rect 1692 3356 1735 3358
rect 1692 3355 1693 3356
rect 1687 3354 1693 3355
rect 1734 3355 1735 3356
rect 1739 3355 1740 3359
rect 1734 3354 1740 3355
rect 2207 3355 2213 3356
rect 2207 3351 2208 3355
rect 2212 3354 2213 3355
rect 2224 3354 2226 3360
rect 2350 3359 2351 3360
rect 2355 3359 2356 3363
rect 2350 3358 2356 3359
rect 2212 3352 2226 3354
rect 2230 3355 2236 3356
rect 2212 3351 2213 3352
rect 2207 3350 2213 3351
rect 2230 3351 2231 3355
rect 2235 3354 2236 3355
rect 2343 3355 2349 3356
rect 2343 3354 2344 3355
rect 2235 3352 2344 3354
rect 2235 3351 2236 3352
rect 2230 3350 2236 3351
rect 2343 3351 2344 3352
rect 2348 3351 2349 3355
rect 2343 3350 2349 3351
rect 2366 3355 2372 3356
rect 2366 3351 2367 3355
rect 2371 3354 2372 3355
rect 2479 3355 2485 3356
rect 2479 3354 2480 3355
rect 2371 3352 2480 3354
rect 2371 3351 2372 3352
rect 2366 3350 2372 3351
rect 2479 3351 2480 3352
rect 2484 3351 2485 3355
rect 2479 3350 2485 3351
rect 2502 3355 2508 3356
rect 2502 3351 2503 3355
rect 2507 3354 2508 3355
rect 2615 3355 2621 3356
rect 2615 3354 2616 3355
rect 2507 3352 2616 3354
rect 2507 3351 2508 3352
rect 2502 3350 2508 3351
rect 2615 3351 2616 3352
rect 2620 3351 2621 3355
rect 2615 3350 2621 3351
rect 2751 3355 2757 3356
rect 2751 3351 2752 3355
rect 2756 3354 2757 3355
rect 2782 3355 2788 3356
rect 2782 3354 2783 3355
rect 2756 3352 2783 3354
rect 2756 3351 2757 3352
rect 2751 3350 2757 3351
rect 2782 3351 2783 3352
rect 2787 3351 2788 3355
rect 2782 3350 2788 3351
rect 2887 3355 2893 3356
rect 2887 3351 2888 3355
rect 2892 3354 2893 3355
rect 2918 3355 2924 3356
rect 2918 3354 2919 3355
rect 2892 3352 2919 3354
rect 2892 3351 2893 3352
rect 2887 3350 2893 3351
rect 2918 3351 2919 3352
rect 2923 3351 2924 3355
rect 2918 3350 2924 3351
rect 3023 3355 3029 3356
rect 3023 3351 3024 3355
rect 3028 3354 3029 3355
rect 3054 3355 3060 3356
rect 3054 3354 3055 3355
rect 3028 3352 3055 3354
rect 3028 3351 3029 3352
rect 3023 3350 3029 3351
rect 3054 3351 3055 3352
rect 3059 3351 3060 3355
rect 3054 3350 3060 3351
rect 3167 3355 3173 3356
rect 3167 3351 3168 3355
rect 3172 3354 3173 3355
rect 3214 3355 3220 3356
rect 3214 3354 3215 3355
rect 3172 3352 3215 3354
rect 3172 3351 3173 3352
rect 3167 3350 3173 3351
rect 3214 3351 3215 3352
rect 3219 3351 3220 3355
rect 3214 3350 3220 3351
rect 110 3344 116 3345
rect 1766 3344 1772 3345
rect 110 3340 111 3344
rect 115 3340 116 3344
rect 110 3339 116 3340
rect 134 3343 140 3344
rect 134 3339 135 3343
rect 139 3339 140 3343
rect 134 3338 140 3339
rect 326 3343 332 3344
rect 326 3339 327 3343
rect 331 3339 332 3343
rect 326 3338 332 3339
rect 534 3343 540 3344
rect 534 3339 535 3343
rect 539 3339 540 3343
rect 534 3338 540 3339
rect 742 3343 748 3344
rect 742 3339 743 3343
rect 747 3339 748 3343
rect 742 3338 748 3339
rect 934 3343 940 3344
rect 934 3339 935 3343
rect 939 3339 940 3343
rect 934 3338 940 3339
rect 1118 3343 1124 3344
rect 1118 3339 1119 3343
rect 1123 3339 1124 3343
rect 1118 3338 1124 3339
rect 1294 3343 1300 3344
rect 1294 3339 1295 3343
rect 1299 3339 1300 3343
rect 1294 3338 1300 3339
rect 1462 3343 1468 3344
rect 1462 3339 1463 3343
rect 1467 3339 1468 3343
rect 1462 3338 1468 3339
rect 1638 3343 1644 3344
rect 1638 3339 1639 3343
rect 1643 3339 1644 3343
rect 1766 3340 1767 3344
rect 1771 3340 1772 3344
rect 1766 3339 1772 3340
rect 1806 3340 1812 3341
rect 3462 3340 3468 3341
rect 1638 3338 1644 3339
rect 1806 3336 1807 3340
rect 1811 3336 1812 3340
rect 247 3335 253 3336
rect 247 3331 248 3335
rect 252 3334 253 3335
rect 606 3335 612 3336
rect 252 3332 369 3334
rect 252 3331 253 3332
rect 247 3330 253 3331
rect 606 3331 607 3335
rect 611 3331 612 3335
rect 606 3330 612 3331
rect 614 3335 620 3336
rect 614 3331 615 3335
rect 619 3334 620 3335
rect 1006 3335 1012 3336
rect 619 3332 785 3334
rect 619 3331 620 3332
rect 614 3330 620 3331
rect 1006 3331 1007 3335
rect 1011 3331 1012 3335
rect 1006 3330 1012 3331
rect 1070 3335 1076 3336
rect 1070 3331 1071 3335
rect 1075 3334 1076 3335
rect 1198 3335 1204 3336
rect 1075 3332 1161 3334
rect 1075 3331 1076 3332
rect 1070 3330 1076 3331
rect 1198 3331 1199 3335
rect 1203 3334 1204 3335
rect 1374 3335 1380 3336
rect 1203 3332 1337 3334
rect 1203 3331 1204 3332
rect 1198 3330 1204 3331
rect 1374 3331 1375 3335
rect 1379 3334 1380 3335
rect 1598 3335 1604 3336
rect 1806 3335 1812 3336
rect 2158 3339 2164 3340
rect 2158 3335 2159 3339
rect 2163 3335 2164 3339
rect 1379 3332 1505 3334
rect 1379 3331 1380 3332
rect 1374 3330 1380 3331
rect 1598 3331 1599 3335
rect 1603 3334 1604 3335
rect 2158 3334 2164 3335
rect 2294 3339 2300 3340
rect 2294 3335 2295 3339
rect 2299 3335 2300 3339
rect 2294 3334 2300 3335
rect 2430 3339 2436 3340
rect 2430 3335 2431 3339
rect 2435 3335 2436 3339
rect 2430 3334 2436 3335
rect 2566 3339 2572 3340
rect 2566 3335 2567 3339
rect 2571 3335 2572 3339
rect 2566 3334 2572 3335
rect 2702 3339 2708 3340
rect 2702 3335 2703 3339
rect 2707 3335 2708 3339
rect 2702 3334 2708 3335
rect 2838 3339 2844 3340
rect 2838 3335 2839 3339
rect 2843 3335 2844 3339
rect 2838 3334 2844 3335
rect 2974 3339 2980 3340
rect 2974 3335 2975 3339
rect 2979 3335 2980 3339
rect 2974 3334 2980 3335
rect 3118 3339 3124 3340
rect 3118 3335 3119 3339
rect 3123 3335 3124 3339
rect 3462 3336 3463 3340
rect 3467 3336 3468 3340
rect 3462 3335 3468 3336
rect 3118 3334 3124 3335
rect 1603 3332 1681 3334
rect 1603 3331 1604 3332
rect 1598 3330 1604 3331
rect 2230 3331 2236 3332
rect 110 3327 116 3328
rect 110 3323 111 3327
rect 115 3323 116 3327
rect 198 3327 204 3328
rect 110 3322 116 3323
rect 134 3324 140 3325
rect 134 3320 135 3324
rect 139 3320 140 3324
rect 198 3323 199 3327
rect 203 3326 204 3327
rect 208 3326 210 3329
rect 203 3324 210 3326
rect 1766 3327 1772 3328
rect 326 3324 332 3325
rect 203 3323 204 3324
rect 198 3322 204 3323
rect 134 3319 140 3320
rect 326 3320 327 3324
rect 331 3320 332 3324
rect 326 3319 332 3320
rect 534 3324 540 3325
rect 534 3320 535 3324
rect 539 3320 540 3324
rect 534 3319 540 3320
rect 742 3324 748 3325
rect 742 3320 743 3324
rect 747 3320 748 3324
rect 742 3319 748 3320
rect 934 3324 940 3325
rect 934 3320 935 3324
rect 939 3320 940 3324
rect 934 3319 940 3320
rect 1118 3324 1124 3325
rect 1118 3320 1119 3324
rect 1123 3320 1124 3324
rect 1118 3319 1124 3320
rect 1294 3324 1300 3325
rect 1294 3320 1295 3324
rect 1299 3320 1300 3324
rect 1294 3319 1300 3320
rect 1462 3324 1468 3325
rect 1462 3320 1463 3324
rect 1467 3320 1468 3324
rect 1462 3319 1468 3320
rect 1638 3324 1644 3325
rect 1638 3320 1639 3324
rect 1643 3320 1644 3324
rect 1766 3323 1767 3327
rect 1771 3323 1772 3327
rect 2230 3327 2231 3331
rect 2235 3327 2236 3331
rect 2230 3326 2236 3327
rect 2366 3331 2372 3332
rect 2366 3327 2367 3331
rect 2371 3327 2372 3331
rect 2366 3326 2372 3327
rect 2502 3331 2508 3332
rect 2502 3327 2503 3331
rect 2507 3327 2508 3331
rect 2774 3331 2780 3332
rect 2502 3326 2508 3327
rect 2638 3327 2644 3328
rect 1766 3322 1772 3323
rect 1806 3323 1812 3324
rect 1638 3319 1644 3320
rect 1806 3319 1807 3323
rect 1811 3319 1812 3323
rect 2638 3323 2639 3327
rect 2643 3323 2644 3327
rect 2774 3327 2775 3331
rect 2779 3327 2780 3331
rect 2918 3331 2924 3332
rect 2774 3326 2780 3327
rect 2910 3327 2916 3328
rect 2638 3322 2644 3323
rect 2910 3323 2911 3327
rect 2915 3323 2916 3327
rect 2918 3327 2919 3331
rect 2923 3330 2924 3331
rect 3054 3331 3060 3332
rect 2923 3328 3017 3330
rect 2923 3327 2924 3328
rect 2918 3326 2924 3327
rect 3054 3327 3055 3331
rect 3059 3330 3060 3331
rect 3059 3328 3161 3330
rect 3059 3327 3060 3328
rect 3054 3326 3060 3327
rect 2910 3322 2916 3323
rect 3462 3323 3468 3324
rect 1806 3318 1812 3319
rect 2158 3320 2164 3321
rect 2158 3316 2159 3320
rect 2163 3316 2164 3320
rect 2158 3315 2164 3316
rect 2294 3320 2300 3321
rect 2294 3316 2295 3320
rect 2299 3316 2300 3320
rect 2294 3315 2300 3316
rect 2430 3320 2436 3321
rect 2430 3316 2431 3320
rect 2435 3316 2436 3320
rect 2430 3315 2436 3316
rect 2566 3320 2572 3321
rect 2566 3316 2567 3320
rect 2571 3316 2572 3320
rect 2566 3315 2572 3316
rect 2702 3320 2708 3321
rect 2702 3316 2703 3320
rect 2707 3316 2708 3320
rect 2702 3315 2708 3316
rect 2838 3320 2844 3321
rect 2838 3316 2839 3320
rect 2843 3316 2844 3320
rect 2838 3315 2844 3316
rect 2974 3320 2980 3321
rect 2974 3316 2975 3320
rect 2979 3316 2980 3320
rect 2974 3315 2980 3316
rect 3118 3320 3124 3321
rect 3118 3316 3119 3320
rect 3123 3316 3124 3320
rect 3462 3319 3463 3323
rect 3467 3319 3468 3323
rect 3462 3318 3468 3319
rect 3118 3315 3124 3316
rect 234 3279 240 3280
rect 234 3275 235 3279
rect 239 3278 240 3279
rect 239 3276 730 3278
rect 239 3275 240 3276
rect 234 3274 240 3275
rect 134 3272 140 3273
rect 110 3269 116 3270
rect 110 3265 111 3269
rect 115 3265 116 3269
rect 134 3268 135 3272
rect 139 3268 140 3272
rect 134 3267 140 3268
rect 278 3272 284 3273
rect 278 3268 279 3272
rect 283 3268 284 3272
rect 278 3267 284 3268
rect 462 3272 468 3273
rect 462 3268 463 3272
rect 467 3268 468 3272
rect 462 3267 468 3268
rect 646 3272 652 3273
rect 646 3268 647 3272
rect 651 3268 652 3272
rect 646 3267 652 3268
rect 110 3264 116 3265
rect 206 3263 212 3264
rect 206 3259 207 3263
rect 211 3259 212 3263
rect 206 3258 212 3259
rect 350 3263 356 3264
rect 350 3259 351 3263
rect 355 3259 356 3263
rect 350 3258 356 3259
rect 534 3263 540 3264
rect 534 3259 535 3263
rect 539 3259 540 3263
rect 534 3258 540 3259
rect 718 3263 724 3264
rect 718 3259 719 3263
rect 723 3259 724 3263
rect 728 3262 730 3276
rect 2086 3276 2092 3277
rect 1806 3273 1812 3274
rect 830 3272 836 3273
rect 830 3268 831 3272
rect 835 3268 836 3272
rect 830 3267 836 3268
rect 1006 3272 1012 3273
rect 1006 3268 1007 3272
rect 1011 3268 1012 3272
rect 1006 3267 1012 3268
rect 1174 3272 1180 3273
rect 1174 3268 1175 3272
rect 1179 3268 1180 3272
rect 1174 3267 1180 3268
rect 1342 3272 1348 3273
rect 1342 3268 1343 3272
rect 1347 3268 1348 3272
rect 1342 3267 1348 3268
rect 1502 3272 1508 3273
rect 1502 3268 1503 3272
rect 1507 3268 1508 3272
rect 1502 3267 1508 3268
rect 1670 3272 1676 3273
rect 1670 3268 1671 3272
rect 1675 3268 1676 3272
rect 1670 3267 1676 3268
rect 1766 3269 1772 3270
rect 1766 3265 1767 3269
rect 1771 3265 1772 3269
rect 1806 3269 1807 3273
rect 1811 3269 1812 3273
rect 2086 3272 2087 3276
rect 2091 3272 2092 3276
rect 2086 3271 2092 3272
rect 2238 3276 2244 3277
rect 2238 3272 2239 3276
rect 2243 3272 2244 3276
rect 2238 3271 2244 3272
rect 2398 3276 2404 3277
rect 2398 3272 2399 3276
rect 2403 3272 2404 3276
rect 2398 3271 2404 3272
rect 2558 3276 2564 3277
rect 2558 3272 2559 3276
rect 2563 3272 2564 3276
rect 2558 3271 2564 3272
rect 2718 3276 2724 3277
rect 2718 3272 2719 3276
rect 2723 3272 2724 3276
rect 2718 3271 2724 3272
rect 2878 3276 2884 3277
rect 2878 3272 2879 3276
rect 2883 3272 2884 3276
rect 2878 3271 2884 3272
rect 3038 3276 3044 3277
rect 3038 3272 3039 3276
rect 3043 3272 3044 3276
rect 3038 3271 3044 3272
rect 3198 3276 3204 3277
rect 3198 3272 3199 3276
rect 3203 3272 3204 3276
rect 3198 3271 3204 3272
rect 3462 3273 3468 3274
rect 1806 3268 1812 3269
rect 3462 3269 3463 3273
rect 3467 3269 3468 3273
rect 3462 3268 3468 3269
rect 1766 3264 1772 3265
rect 2158 3267 2164 3268
rect 1114 3263 1120 3264
rect 1114 3262 1115 3263
rect 728 3260 873 3262
rect 1081 3260 1115 3262
rect 718 3258 724 3259
rect 1114 3259 1115 3260
rect 1119 3259 1120 3263
rect 1114 3258 1120 3259
rect 1246 3263 1252 3264
rect 1246 3259 1247 3263
rect 1251 3259 1252 3263
rect 1246 3258 1252 3259
rect 1414 3263 1420 3264
rect 1414 3259 1415 3263
rect 1419 3259 1420 3263
rect 1414 3258 1420 3259
rect 1574 3263 1580 3264
rect 1574 3259 1575 3263
rect 1579 3259 1580 3263
rect 1574 3258 1580 3259
rect 1734 3263 1740 3264
rect 1734 3259 1735 3263
rect 1739 3259 1740 3263
rect 2158 3263 2159 3267
rect 2163 3263 2164 3267
rect 2158 3262 2164 3263
rect 2310 3267 2316 3268
rect 2310 3263 2311 3267
rect 2315 3263 2316 3267
rect 2310 3262 2316 3263
rect 2359 3267 2365 3268
rect 2359 3263 2360 3267
rect 2364 3266 2365 3267
rect 2478 3267 2484 3268
rect 2364 3264 2441 3266
rect 2364 3263 2365 3264
rect 2359 3262 2365 3263
rect 2478 3263 2479 3267
rect 2483 3266 2484 3267
rect 2782 3267 2788 3268
rect 2483 3264 2601 3266
rect 2483 3263 2484 3264
rect 2478 3262 2484 3263
rect 2782 3263 2783 3267
rect 2787 3263 2788 3267
rect 2782 3262 2788 3263
rect 2950 3267 2956 3268
rect 2950 3263 2951 3267
rect 2955 3263 2956 3267
rect 2950 3262 2956 3263
rect 3110 3267 3116 3268
rect 3110 3263 3111 3267
rect 3115 3263 3116 3267
rect 3110 3262 3116 3263
rect 3262 3267 3268 3268
rect 3262 3263 3263 3267
rect 3267 3263 3268 3267
rect 3262 3262 3268 3263
rect 1734 3258 1740 3259
rect 2086 3257 2092 3258
rect 1806 3256 1812 3257
rect 134 3253 140 3254
rect 110 3252 116 3253
rect 110 3248 111 3252
rect 115 3248 116 3252
rect 134 3249 135 3253
rect 139 3249 140 3253
rect 134 3248 140 3249
rect 278 3253 284 3254
rect 278 3249 279 3253
rect 283 3249 284 3253
rect 278 3248 284 3249
rect 462 3253 468 3254
rect 462 3249 463 3253
rect 467 3249 468 3253
rect 462 3248 468 3249
rect 646 3253 652 3254
rect 646 3249 647 3253
rect 651 3249 652 3253
rect 646 3248 652 3249
rect 830 3253 836 3254
rect 830 3249 831 3253
rect 835 3249 836 3253
rect 830 3248 836 3249
rect 1006 3253 1012 3254
rect 1006 3249 1007 3253
rect 1011 3249 1012 3253
rect 1006 3248 1012 3249
rect 1174 3253 1180 3254
rect 1174 3249 1175 3253
rect 1179 3249 1180 3253
rect 1174 3248 1180 3249
rect 1342 3253 1348 3254
rect 1342 3249 1343 3253
rect 1347 3249 1348 3253
rect 1342 3248 1348 3249
rect 1502 3253 1508 3254
rect 1502 3249 1503 3253
rect 1507 3249 1508 3253
rect 1502 3248 1508 3249
rect 1670 3253 1676 3254
rect 1670 3249 1671 3253
rect 1675 3249 1676 3253
rect 1670 3248 1676 3249
rect 1766 3252 1772 3253
rect 1766 3248 1767 3252
rect 1771 3248 1772 3252
rect 1806 3252 1807 3256
rect 1811 3252 1812 3256
rect 2086 3253 2087 3257
rect 2091 3253 2092 3257
rect 2086 3252 2092 3253
rect 2238 3257 2244 3258
rect 2238 3253 2239 3257
rect 2243 3253 2244 3257
rect 2238 3252 2244 3253
rect 2398 3257 2404 3258
rect 2398 3253 2399 3257
rect 2403 3253 2404 3257
rect 2398 3252 2404 3253
rect 2558 3257 2564 3258
rect 2558 3253 2559 3257
rect 2563 3253 2564 3257
rect 2558 3252 2564 3253
rect 2718 3257 2724 3258
rect 2718 3253 2719 3257
rect 2723 3253 2724 3257
rect 2718 3252 2724 3253
rect 2878 3257 2884 3258
rect 2878 3253 2879 3257
rect 2883 3253 2884 3257
rect 2878 3252 2884 3253
rect 3038 3257 3044 3258
rect 3038 3253 3039 3257
rect 3043 3253 3044 3257
rect 3038 3252 3044 3253
rect 3198 3257 3204 3258
rect 3198 3253 3199 3257
rect 3203 3253 3204 3257
rect 3198 3252 3204 3253
rect 3462 3256 3468 3257
rect 3462 3252 3463 3256
rect 3467 3252 3468 3256
rect 1806 3251 1812 3252
rect 3462 3251 3468 3252
rect 110 3247 116 3248
rect 1766 3247 1772 3248
rect 2135 3239 2141 3240
rect 183 3235 189 3236
rect 183 3231 184 3235
rect 188 3234 189 3235
rect 198 3235 204 3236
rect 198 3234 199 3235
rect 188 3232 199 3234
rect 188 3231 189 3232
rect 183 3230 189 3231
rect 198 3231 199 3232
rect 203 3231 204 3235
rect 198 3230 204 3231
rect 206 3235 212 3236
rect 206 3231 207 3235
rect 211 3234 212 3235
rect 327 3235 333 3236
rect 327 3234 328 3235
rect 211 3232 328 3234
rect 211 3231 212 3232
rect 206 3230 212 3231
rect 327 3231 328 3232
rect 332 3231 333 3235
rect 327 3230 333 3231
rect 350 3235 356 3236
rect 350 3231 351 3235
rect 355 3234 356 3235
rect 511 3235 517 3236
rect 511 3234 512 3235
rect 355 3232 512 3234
rect 355 3231 356 3232
rect 350 3230 356 3231
rect 511 3231 512 3232
rect 516 3231 517 3235
rect 511 3230 517 3231
rect 534 3235 540 3236
rect 534 3231 535 3235
rect 539 3234 540 3235
rect 695 3235 701 3236
rect 695 3234 696 3235
rect 539 3232 696 3234
rect 539 3231 540 3232
rect 534 3230 540 3231
rect 695 3231 696 3232
rect 700 3231 701 3235
rect 695 3230 701 3231
rect 718 3235 724 3236
rect 718 3231 719 3235
rect 723 3234 724 3235
rect 879 3235 885 3236
rect 879 3234 880 3235
rect 723 3232 880 3234
rect 723 3231 724 3232
rect 718 3230 724 3231
rect 879 3231 880 3232
rect 884 3231 885 3235
rect 879 3230 885 3231
rect 1055 3235 1061 3236
rect 1055 3231 1056 3235
rect 1060 3234 1061 3235
rect 1114 3235 1120 3236
rect 1060 3232 1110 3234
rect 1060 3231 1061 3232
rect 1055 3230 1061 3231
rect 1108 3226 1110 3232
rect 1114 3231 1115 3235
rect 1119 3234 1120 3235
rect 1223 3235 1229 3236
rect 1223 3234 1224 3235
rect 1119 3232 1224 3234
rect 1119 3231 1120 3232
rect 1114 3230 1120 3231
rect 1223 3231 1224 3232
rect 1228 3231 1229 3235
rect 1223 3230 1229 3231
rect 1246 3235 1252 3236
rect 1246 3231 1247 3235
rect 1251 3234 1252 3235
rect 1391 3235 1397 3236
rect 1391 3234 1392 3235
rect 1251 3232 1392 3234
rect 1251 3231 1252 3232
rect 1246 3230 1252 3231
rect 1391 3231 1392 3232
rect 1396 3231 1397 3235
rect 1391 3230 1397 3231
rect 1414 3235 1420 3236
rect 1414 3231 1415 3235
rect 1419 3234 1420 3235
rect 1551 3235 1557 3236
rect 1551 3234 1552 3235
rect 1419 3232 1552 3234
rect 1419 3231 1420 3232
rect 1414 3230 1420 3231
rect 1551 3231 1552 3232
rect 1556 3231 1557 3235
rect 1551 3230 1557 3231
rect 1574 3235 1580 3236
rect 1574 3231 1575 3235
rect 1579 3234 1580 3235
rect 1719 3235 1725 3236
rect 1719 3234 1720 3235
rect 1579 3232 1720 3234
rect 1579 3231 1580 3232
rect 1574 3230 1580 3231
rect 1719 3231 1720 3232
rect 1724 3231 1725 3235
rect 2135 3235 2136 3239
rect 2140 3238 2141 3239
rect 2158 3239 2164 3240
rect 2140 3236 2154 3238
rect 2140 3235 2141 3236
rect 2135 3234 2141 3235
rect 1719 3230 1725 3231
rect 2152 3230 2154 3236
rect 2158 3235 2159 3239
rect 2163 3238 2164 3239
rect 2287 3239 2293 3240
rect 2287 3238 2288 3239
rect 2163 3236 2288 3238
rect 2163 3235 2164 3236
rect 2158 3234 2164 3235
rect 2287 3235 2288 3236
rect 2292 3235 2293 3239
rect 2287 3234 2293 3235
rect 2447 3239 2453 3240
rect 2447 3235 2448 3239
rect 2452 3238 2453 3239
rect 2478 3239 2484 3240
rect 2478 3238 2479 3239
rect 2452 3236 2479 3238
rect 2452 3235 2453 3236
rect 2447 3234 2453 3235
rect 2478 3235 2479 3236
rect 2483 3235 2484 3239
rect 2478 3234 2484 3235
rect 2607 3239 2613 3240
rect 2607 3235 2608 3239
rect 2612 3238 2613 3239
rect 2638 3239 2644 3240
rect 2638 3238 2639 3239
rect 2612 3236 2639 3238
rect 2612 3235 2613 3236
rect 2607 3234 2613 3235
rect 2638 3235 2639 3236
rect 2643 3235 2644 3239
rect 2638 3234 2644 3235
rect 2758 3239 2764 3240
rect 2758 3235 2759 3239
rect 2763 3238 2764 3239
rect 2767 3239 2773 3240
rect 2767 3238 2768 3239
rect 2763 3236 2768 3238
rect 2763 3235 2764 3236
rect 2758 3234 2764 3235
rect 2767 3235 2768 3236
rect 2772 3235 2773 3239
rect 2767 3234 2773 3235
rect 2910 3239 2916 3240
rect 2910 3235 2911 3239
rect 2915 3238 2916 3239
rect 2927 3239 2933 3240
rect 2927 3238 2928 3239
rect 2915 3236 2928 3238
rect 2915 3235 2916 3236
rect 2910 3234 2916 3235
rect 2927 3235 2928 3236
rect 2932 3235 2933 3239
rect 2927 3234 2933 3235
rect 2950 3239 2956 3240
rect 2950 3235 2951 3239
rect 2955 3238 2956 3239
rect 3087 3239 3093 3240
rect 3087 3238 3088 3239
rect 2955 3236 3088 3238
rect 2955 3235 2956 3236
rect 2950 3234 2956 3235
rect 3087 3235 3088 3236
rect 3092 3235 3093 3239
rect 3087 3234 3093 3235
rect 3110 3239 3116 3240
rect 3110 3235 3111 3239
rect 3115 3238 3116 3239
rect 3247 3239 3253 3240
rect 3247 3238 3248 3239
rect 3115 3236 3248 3238
rect 3115 3235 3116 3236
rect 3110 3234 3116 3235
rect 3247 3235 3248 3236
rect 3252 3235 3253 3239
rect 3247 3234 3253 3235
rect 2359 3231 2365 3232
rect 2359 3230 2360 3231
rect 1256 3228 1386 3230
rect 2152 3228 2360 3230
rect 1256 3226 1258 3228
rect 1108 3224 1258 3226
rect 1384 3226 1386 3228
rect 1398 3227 1404 3228
rect 1398 3226 1399 3227
rect 1384 3224 1399 3226
rect 1278 3223 1284 3224
rect 1278 3222 1279 3223
rect 1159 3220 1279 3222
rect 1159 3218 1161 3220
rect 1278 3219 1279 3220
rect 1283 3219 1284 3223
rect 1398 3223 1399 3224
rect 1403 3223 1404 3227
rect 2359 3227 2360 3228
rect 2364 3227 2365 3231
rect 2359 3226 2365 3227
rect 1398 3222 1404 3223
rect 1959 3223 1968 3224
rect 1278 3218 1284 3219
rect 1959 3219 1960 3223
rect 1967 3219 1968 3223
rect 1959 3218 1968 3219
rect 1982 3223 1988 3224
rect 1982 3219 1983 3223
rect 1987 3222 1988 3223
rect 2095 3223 2101 3224
rect 2095 3222 2096 3223
rect 1987 3220 2096 3222
rect 1987 3219 1988 3220
rect 1982 3218 1988 3219
rect 2095 3219 2096 3220
rect 2100 3219 2101 3223
rect 2095 3218 2101 3219
rect 2118 3223 2124 3224
rect 2118 3219 2119 3223
rect 2123 3222 2124 3223
rect 2247 3223 2253 3224
rect 2247 3222 2248 3223
rect 2123 3220 2248 3222
rect 2123 3219 2124 3220
rect 2118 3218 2124 3219
rect 2247 3219 2248 3220
rect 2252 3219 2253 3223
rect 2247 3218 2253 3219
rect 2310 3223 2316 3224
rect 2310 3219 2311 3223
rect 2315 3222 2316 3223
rect 2407 3223 2413 3224
rect 2407 3222 2408 3223
rect 2315 3220 2408 3222
rect 2315 3219 2316 3220
rect 2310 3218 2316 3219
rect 2407 3219 2408 3220
rect 2412 3219 2413 3223
rect 2407 3218 2413 3219
rect 2430 3223 2436 3224
rect 2430 3219 2431 3223
rect 2435 3222 2436 3223
rect 2575 3223 2581 3224
rect 2575 3222 2576 3223
rect 2435 3220 2576 3222
rect 2435 3219 2436 3220
rect 2430 3218 2436 3219
rect 2575 3219 2576 3220
rect 2580 3219 2581 3223
rect 2575 3218 2581 3219
rect 2735 3223 2741 3224
rect 2735 3219 2736 3223
rect 2740 3222 2741 3223
rect 2806 3223 2812 3224
rect 2806 3222 2807 3223
rect 2740 3220 2807 3222
rect 2740 3219 2741 3220
rect 2735 3218 2741 3219
rect 2806 3219 2807 3220
rect 2811 3219 2812 3223
rect 2806 3218 2812 3219
rect 2830 3223 2836 3224
rect 2830 3219 2831 3223
rect 2835 3222 2836 3223
rect 2895 3223 2901 3224
rect 2895 3222 2896 3223
rect 2835 3220 2896 3222
rect 2835 3219 2836 3220
rect 2830 3218 2836 3219
rect 2895 3219 2896 3220
rect 2900 3219 2901 3223
rect 2895 3218 2901 3219
rect 3055 3223 3061 3224
rect 3055 3219 3056 3223
rect 3060 3222 3061 3223
rect 3087 3223 3093 3224
rect 3087 3222 3088 3223
rect 3060 3220 3088 3222
rect 3060 3219 3061 3220
rect 3055 3218 3061 3219
rect 3087 3219 3088 3220
rect 3092 3219 3093 3223
rect 3087 3218 3093 3219
rect 3215 3223 3221 3224
rect 3215 3219 3216 3223
rect 3220 3222 3221 3223
rect 3262 3223 3268 3224
rect 3262 3222 3263 3223
rect 3220 3220 3263 3222
rect 3220 3219 3221 3220
rect 3215 3218 3221 3219
rect 3262 3219 3263 3220
rect 3267 3219 3268 3223
rect 3262 3218 3268 3219
rect 3302 3223 3308 3224
rect 3302 3219 3303 3223
rect 3307 3222 3308 3223
rect 3383 3223 3389 3224
rect 3383 3222 3384 3223
rect 3307 3220 3384 3222
rect 3307 3219 3308 3220
rect 3302 3218 3308 3219
rect 3383 3219 3384 3220
rect 3388 3219 3389 3223
rect 3383 3218 3389 3219
rect 1088 3216 1161 3218
rect 231 3215 240 3216
rect 231 3211 232 3215
rect 239 3211 240 3215
rect 231 3210 240 3211
rect 254 3215 260 3216
rect 254 3211 255 3215
rect 259 3214 260 3215
rect 375 3215 381 3216
rect 375 3214 376 3215
rect 259 3212 376 3214
rect 259 3211 260 3212
rect 254 3210 260 3211
rect 375 3211 376 3212
rect 380 3211 381 3215
rect 375 3210 381 3211
rect 398 3215 404 3216
rect 398 3211 399 3215
rect 403 3214 404 3215
rect 535 3215 541 3216
rect 535 3214 536 3215
rect 403 3212 536 3214
rect 403 3211 404 3212
rect 398 3210 404 3211
rect 535 3211 536 3212
rect 540 3211 541 3215
rect 535 3210 541 3211
rect 558 3215 564 3216
rect 558 3211 559 3215
rect 563 3214 564 3215
rect 695 3215 701 3216
rect 695 3214 696 3215
rect 563 3212 696 3214
rect 563 3211 564 3212
rect 558 3210 564 3211
rect 695 3211 696 3212
rect 700 3211 701 3215
rect 695 3210 701 3211
rect 718 3215 724 3216
rect 718 3211 719 3215
rect 723 3214 724 3215
rect 855 3215 861 3216
rect 855 3214 856 3215
rect 723 3212 856 3214
rect 723 3211 724 3212
rect 718 3210 724 3211
rect 855 3211 856 3212
rect 860 3211 861 3215
rect 855 3210 861 3211
rect 1015 3215 1021 3216
rect 1015 3211 1016 3215
rect 1020 3214 1021 3215
rect 1088 3214 1090 3216
rect 1183 3215 1189 3216
rect 1183 3214 1184 3215
rect 1020 3212 1090 3214
rect 1159 3212 1184 3214
rect 1020 3211 1021 3212
rect 1015 3210 1021 3211
rect 1094 3211 1100 3212
rect 1094 3207 1095 3211
rect 1099 3210 1100 3211
rect 1159 3210 1161 3212
rect 1183 3211 1184 3212
rect 1188 3211 1189 3215
rect 1183 3210 1189 3211
rect 1250 3215 1256 3216
rect 1250 3211 1251 3215
rect 1255 3214 1256 3215
rect 1351 3215 1357 3216
rect 1351 3214 1352 3215
rect 1255 3212 1352 3214
rect 1255 3211 1256 3212
rect 1250 3210 1256 3211
rect 1351 3211 1352 3212
rect 1356 3211 1357 3215
rect 1351 3210 1357 3211
rect 1374 3215 1380 3216
rect 1374 3211 1375 3215
rect 1379 3214 1380 3215
rect 1519 3215 1525 3216
rect 1519 3214 1520 3215
rect 1379 3212 1520 3214
rect 1379 3211 1380 3212
rect 1374 3210 1380 3211
rect 1519 3211 1520 3212
rect 1524 3211 1525 3215
rect 1519 3210 1525 3211
rect 1099 3208 1161 3210
rect 1806 3208 1812 3209
rect 3462 3208 3468 3209
rect 1099 3207 1100 3208
rect 1094 3206 1100 3207
rect 1806 3204 1807 3208
rect 1811 3204 1812 3208
rect 1806 3203 1812 3204
rect 1910 3207 1916 3208
rect 1910 3203 1911 3207
rect 1915 3203 1916 3207
rect 1910 3202 1916 3203
rect 2046 3207 2052 3208
rect 2046 3203 2047 3207
rect 2051 3203 2052 3207
rect 2046 3202 2052 3203
rect 2198 3207 2204 3208
rect 2198 3203 2199 3207
rect 2203 3203 2204 3207
rect 2198 3202 2204 3203
rect 2358 3207 2364 3208
rect 2358 3203 2359 3207
rect 2363 3203 2364 3207
rect 2358 3202 2364 3203
rect 2526 3207 2532 3208
rect 2526 3203 2527 3207
rect 2531 3203 2532 3207
rect 2526 3202 2532 3203
rect 2686 3207 2692 3208
rect 2686 3203 2687 3207
rect 2691 3203 2692 3207
rect 2686 3202 2692 3203
rect 2846 3207 2852 3208
rect 2846 3203 2847 3207
rect 2851 3203 2852 3207
rect 2846 3202 2852 3203
rect 3006 3207 3012 3208
rect 3006 3203 3007 3207
rect 3011 3203 3012 3207
rect 3006 3202 3012 3203
rect 3166 3207 3172 3208
rect 3166 3203 3167 3207
rect 3171 3203 3172 3207
rect 3166 3202 3172 3203
rect 3334 3207 3340 3208
rect 3334 3203 3335 3207
rect 3339 3203 3340 3207
rect 3462 3204 3463 3208
rect 3467 3204 3468 3208
rect 3462 3203 3468 3204
rect 3334 3202 3340 3203
rect 110 3200 116 3201
rect 1766 3200 1772 3201
rect 110 3196 111 3200
rect 115 3196 116 3200
rect 110 3195 116 3196
rect 182 3199 188 3200
rect 182 3195 183 3199
rect 187 3195 188 3199
rect 182 3194 188 3195
rect 326 3199 332 3200
rect 326 3195 327 3199
rect 331 3195 332 3199
rect 326 3194 332 3195
rect 486 3199 492 3200
rect 486 3195 487 3199
rect 491 3195 492 3199
rect 486 3194 492 3195
rect 646 3199 652 3200
rect 646 3195 647 3199
rect 651 3195 652 3199
rect 646 3194 652 3195
rect 806 3199 812 3200
rect 806 3195 807 3199
rect 811 3195 812 3199
rect 806 3194 812 3195
rect 966 3199 972 3200
rect 966 3195 967 3199
rect 971 3195 972 3199
rect 966 3194 972 3195
rect 1134 3199 1140 3200
rect 1134 3195 1135 3199
rect 1139 3195 1140 3199
rect 1134 3194 1140 3195
rect 1302 3199 1308 3200
rect 1302 3195 1303 3199
rect 1307 3195 1308 3199
rect 1302 3194 1308 3195
rect 1470 3199 1476 3200
rect 1470 3195 1471 3199
rect 1475 3195 1476 3199
rect 1766 3196 1767 3200
rect 1771 3196 1772 3200
rect 1766 3195 1772 3196
rect 1982 3199 1988 3200
rect 1982 3195 1983 3199
rect 1987 3195 1988 3199
rect 1470 3194 1476 3195
rect 1982 3194 1988 3195
rect 2118 3199 2124 3200
rect 2118 3195 2119 3199
rect 2123 3195 2124 3199
rect 2430 3199 2436 3200
rect 2118 3194 2124 3195
rect 2270 3195 2276 3196
rect 254 3191 260 3192
rect 254 3187 255 3191
rect 259 3187 260 3191
rect 254 3186 260 3187
rect 398 3191 404 3192
rect 398 3187 399 3191
rect 403 3187 404 3191
rect 398 3186 404 3187
rect 558 3191 564 3192
rect 558 3187 559 3191
rect 563 3187 564 3191
rect 558 3186 564 3187
rect 718 3191 724 3192
rect 718 3187 719 3191
rect 723 3187 724 3191
rect 718 3186 724 3187
rect 734 3191 740 3192
rect 734 3187 735 3191
rect 739 3190 740 3191
rect 1094 3191 1100 3192
rect 1094 3190 1095 3191
rect 739 3188 849 3190
rect 1041 3188 1095 3190
rect 739 3187 740 3188
rect 734 3186 740 3187
rect 1094 3187 1095 3188
rect 1099 3187 1100 3191
rect 1250 3191 1256 3192
rect 1250 3190 1251 3191
rect 1209 3188 1251 3190
rect 1094 3186 1100 3187
rect 1250 3187 1251 3188
rect 1255 3187 1256 3191
rect 1250 3186 1256 3187
rect 1374 3191 1380 3192
rect 1374 3187 1375 3191
rect 1379 3187 1380 3191
rect 1374 3186 1380 3187
rect 1398 3191 1404 3192
rect 1398 3187 1399 3191
rect 1403 3190 1404 3191
rect 1806 3191 1812 3192
rect 1403 3188 1513 3190
rect 1403 3187 1404 3188
rect 1398 3186 1404 3187
rect 1806 3187 1807 3191
rect 1811 3187 1812 3191
rect 2270 3191 2271 3195
rect 2275 3191 2276 3195
rect 2430 3195 2431 3199
rect 2435 3195 2436 3199
rect 2430 3194 2436 3195
rect 2478 3199 2484 3200
rect 2478 3195 2479 3199
rect 2483 3198 2484 3199
rect 2758 3199 2764 3200
rect 2483 3196 2569 3198
rect 2483 3195 2484 3196
rect 2478 3194 2484 3195
rect 2758 3195 2759 3199
rect 2763 3195 2764 3199
rect 2758 3194 2764 3195
rect 2806 3199 2812 3200
rect 2806 3195 2807 3199
rect 2811 3198 2812 3199
rect 2966 3199 2972 3200
rect 2811 3196 2889 3198
rect 2811 3195 2812 3196
rect 2806 3194 2812 3195
rect 2966 3195 2967 3199
rect 2971 3198 2972 3199
rect 3087 3199 3093 3200
rect 2971 3196 3049 3198
rect 2971 3195 2972 3196
rect 2966 3194 2972 3195
rect 3087 3195 3088 3199
rect 3092 3198 3093 3199
rect 3092 3196 3209 3198
rect 3092 3195 3093 3196
rect 3087 3194 3093 3195
rect 3406 3195 3412 3196
rect 2270 3190 2276 3191
rect 3406 3191 3407 3195
rect 3411 3191 3412 3195
rect 3406 3190 3412 3191
rect 3462 3191 3468 3192
rect 1806 3186 1812 3187
rect 1910 3188 1916 3189
rect 1910 3184 1911 3188
rect 1915 3184 1916 3188
rect 110 3183 116 3184
rect 110 3179 111 3183
rect 115 3179 116 3183
rect 1766 3183 1772 3184
rect 1910 3183 1916 3184
rect 2046 3188 2052 3189
rect 2046 3184 2047 3188
rect 2051 3184 2052 3188
rect 2046 3183 2052 3184
rect 2198 3188 2204 3189
rect 2198 3184 2199 3188
rect 2203 3184 2204 3188
rect 2198 3183 2204 3184
rect 2358 3188 2364 3189
rect 2358 3184 2359 3188
rect 2363 3184 2364 3188
rect 2358 3183 2364 3184
rect 2526 3188 2532 3189
rect 2526 3184 2527 3188
rect 2531 3184 2532 3188
rect 2526 3183 2532 3184
rect 2686 3188 2692 3189
rect 2686 3184 2687 3188
rect 2691 3184 2692 3188
rect 2686 3183 2692 3184
rect 2846 3188 2852 3189
rect 2846 3184 2847 3188
rect 2851 3184 2852 3188
rect 2846 3183 2852 3184
rect 3006 3188 3012 3189
rect 3006 3184 3007 3188
rect 3011 3184 3012 3188
rect 3006 3183 3012 3184
rect 3166 3188 3172 3189
rect 3166 3184 3167 3188
rect 3171 3184 3172 3188
rect 3166 3183 3172 3184
rect 3334 3188 3340 3189
rect 3334 3184 3335 3188
rect 3339 3184 3340 3188
rect 3462 3187 3463 3191
rect 3467 3187 3468 3191
rect 3462 3186 3468 3187
rect 3334 3183 3340 3184
rect 110 3178 116 3179
rect 182 3180 188 3181
rect 182 3176 183 3180
rect 187 3176 188 3180
rect 182 3175 188 3176
rect 326 3180 332 3181
rect 326 3176 327 3180
rect 331 3176 332 3180
rect 326 3175 332 3176
rect 486 3180 492 3181
rect 486 3176 487 3180
rect 491 3176 492 3180
rect 486 3175 492 3176
rect 646 3180 652 3181
rect 646 3176 647 3180
rect 651 3176 652 3180
rect 646 3175 652 3176
rect 806 3180 812 3181
rect 806 3176 807 3180
rect 811 3176 812 3180
rect 806 3175 812 3176
rect 966 3180 972 3181
rect 966 3176 967 3180
rect 971 3176 972 3180
rect 966 3175 972 3176
rect 1134 3180 1140 3181
rect 1134 3176 1135 3180
rect 1139 3176 1140 3180
rect 1134 3175 1140 3176
rect 1302 3180 1308 3181
rect 1302 3176 1303 3180
rect 1307 3176 1308 3180
rect 1302 3175 1308 3176
rect 1470 3180 1476 3181
rect 1470 3176 1471 3180
rect 1475 3176 1476 3180
rect 1766 3179 1767 3183
rect 1771 3179 1772 3183
rect 1766 3178 1772 3179
rect 1962 3179 1968 3180
rect 1470 3175 1476 3176
rect 1962 3175 1963 3179
rect 1967 3178 1968 3179
rect 2478 3179 2484 3180
rect 2478 3178 2479 3179
rect 1967 3176 2479 3178
rect 1967 3175 1968 3176
rect 1962 3174 1968 3175
rect 2478 3175 2479 3176
rect 2483 3175 2484 3179
rect 2478 3174 2484 3175
rect 418 3147 424 3148
rect 418 3143 419 3147
rect 423 3146 424 3147
rect 734 3147 740 3148
rect 734 3146 735 3147
rect 423 3144 735 3146
rect 423 3143 424 3144
rect 418 3142 424 3143
rect 734 3143 735 3144
rect 739 3143 740 3147
rect 734 3142 740 3143
rect 1830 3144 1836 3145
rect 1806 3141 1812 3142
rect 1806 3137 1807 3141
rect 1811 3137 1812 3141
rect 1830 3140 1831 3144
rect 1835 3140 1836 3144
rect 1830 3139 1836 3140
rect 2006 3144 2012 3145
rect 2006 3140 2007 3144
rect 2011 3140 2012 3144
rect 2006 3139 2012 3140
rect 2206 3144 2212 3145
rect 2206 3140 2207 3144
rect 2211 3140 2212 3144
rect 2206 3139 2212 3140
rect 2398 3144 2404 3145
rect 2398 3140 2399 3144
rect 2403 3140 2404 3144
rect 2398 3139 2404 3140
rect 2582 3144 2588 3145
rect 2582 3140 2583 3144
rect 2587 3140 2588 3144
rect 2582 3139 2588 3140
rect 2758 3144 2764 3145
rect 2758 3140 2759 3144
rect 2763 3140 2764 3144
rect 2758 3139 2764 3140
rect 2918 3144 2924 3145
rect 2918 3140 2919 3144
rect 2923 3140 2924 3144
rect 2918 3139 2924 3140
rect 3078 3144 3084 3145
rect 3078 3140 3079 3144
rect 3083 3140 3084 3144
rect 3078 3139 3084 3140
rect 3230 3144 3236 3145
rect 3230 3140 3231 3144
rect 3235 3140 3236 3144
rect 3230 3139 3236 3140
rect 3366 3144 3372 3145
rect 3366 3140 3367 3144
rect 3371 3140 3372 3144
rect 3366 3139 3372 3140
rect 3462 3141 3468 3142
rect 366 3136 372 3137
rect 110 3133 116 3134
rect 110 3129 111 3133
rect 115 3129 116 3133
rect 366 3132 367 3136
rect 371 3132 372 3136
rect 366 3131 372 3132
rect 486 3136 492 3137
rect 486 3132 487 3136
rect 491 3132 492 3136
rect 486 3131 492 3132
rect 606 3136 612 3137
rect 606 3132 607 3136
rect 611 3132 612 3136
rect 606 3131 612 3132
rect 726 3136 732 3137
rect 726 3132 727 3136
rect 731 3132 732 3136
rect 726 3131 732 3132
rect 846 3136 852 3137
rect 846 3132 847 3136
rect 851 3132 852 3136
rect 846 3131 852 3132
rect 966 3136 972 3137
rect 966 3132 967 3136
rect 971 3132 972 3136
rect 966 3131 972 3132
rect 1078 3136 1084 3137
rect 1078 3132 1079 3136
rect 1083 3132 1084 3136
rect 1078 3131 1084 3132
rect 1198 3136 1204 3137
rect 1198 3132 1199 3136
rect 1203 3132 1204 3136
rect 1198 3131 1204 3132
rect 1318 3136 1324 3137
rect 1806 3136 1812 3137
rect 3462 3137 3463 3141
rect 3467 3137 3468 3141
rect 3462 3136 3468 3137
rect 1318 3132 1319 3136
rect 1323 3132 1324 3136
rect 1894 3135 1900 3136
rect 1318 3131 1324 3132
rect 1766 3133 1772 3134
rect 110 3128 116 3129
rect 1766 3129 1767 3133
rect 1771 3129 1772 3133
rect 1894 3131 1895 3135
rect 1899 3131 1900 3135
rect 1894 3130 1900 3131
rect 1910 3135 1916 3136
rect 1910 3131 1911 3135
rect 1915 3134 1916 3135
rect 2278 3135 2284 3136
rect 1915 3132 2049 3134
rect 1915 3131 1916 3132
rect 1910 3130 1916 3131
rect 2278 3131 2279 3135
rect 2283 3131 2284 3135
rect 2278 3130 2284 3131
rect 2286 3135 2292 3136
rect 2286 3131 2287 3135
rect 2291 3134 2292 3135
rect 2742 3135 2748 3136
rect 2742 3134 2743 3135
rect 2291 3132 2441 3134
rect 2657 3132 2743 3134
rect 2291 3131 2292 3132
rect 2286 3130 2292 3131
rect 2742 3131 2743 3132
rect 2747 3131 2748 3135
rect 2742 3130 2748 3131
rect 2830 3135 2836 3136
rect 2830 3131 2831 3135
rect 2835 3131 2836 3135
rect 2830 3130 2836 3131
rect 2990 3135 2996 3136
rect 2990 3131 2991 3135
rect 2995 3131 2996 3135
rect 2990 3130 2996 3131
rect 3150 3135 3156 3136
rect 3150 3131 3151 3135
rect 3155 3131 3156 3135
rect 3150 3130 3156 3131
rect 3302 3135 3308 3136
rect 3302 3131 3303 3135
rect 3307 3131 3308 3135
rect 3302 3130 3308 3131
rect 3430 3135 3436 3136
rect 3430 3131 3431 3135
rect 3435 3131 3436 3135
rect 3430 3130 3436 3131
rect 1766 3128 1772 3129
rect 438 3127 444 3128
rect 438 3123 439 3127
rect 443 3123 444 3127
rect 438 3122 444 3123
rect 558 3127 564 3128
rect 558 3123 559 3127
rect 563 3123 564 3127
rect 558 3122 564 3123
rect 678 3127 684 3128
rect 678 3123 679 3127
rect 683 3123 684 3127
rect 678 3122 684 3123
rect 686 3127 692 3128
rect 686 3123 687 3127
rect 691 3126 692 3127
rect 918 3127 924 3128
rect 691 3124 769 3126
rect 691 3123 692 3124
rect 686 3122 692 3123
rect 918 3123 919 3127
rect 923 3123 924 3127
rect 918 3122 924 3123
rect 1038 3127 1044 3128
rect 1038 3123 1039 3127
rect 1043 3123 1044 3127
rect 1038 3122 1044 3123
rect 1150 3127 1156 3128
rect 1150 3123 1151 3127
rect 1155 3123 1156 3127
rect 1150 3122 1156 3123
rect 1270 3127 1276 3128
rect 1270 3123 1271 3127
rect 1275 3123 1276 3127
rect 1270 3122 1276 3123
rect 1278 3127 1284 3128
rect 1278 3123 1279 3127
rect 1283 3126 1284 3127
rect 1283 3124 1361 3126
rect 1830 3125 1836 3126
rect 1806 3124 1812 3125
rect 1283 3123 1284 3124
rect 1278 3122 1284 3123
rect 1806 3120 1807 3124
rect 1811 3120 1812 3124
rect 1830 3121 1831 3125
rect 1835 3121 1836 3125
rect 1830 3120 1836 3121
rect 2006 3125 2012 3126
rect 2006 3121 2007 3125
rect 2011 3121 2012 3125
rect 2006 3120 2012 3121
rect 2206 3125 2212 3126
rect 2206 3121 2207 3125
rect 2211 3121 2212 3125
rect 2206 3120 2212 3121
rect 2398 3125 2404 3126
rect 2398 3121 2399 3125
rect 2403 3121 2404 3125
rect 2398 3120 2404 3121
rect 2582 3125 2588 3126
rect 2582 3121 2583 3125
rect 2587 3121 2588 3125
rect 2582 3120 2588 3121
rect 2758 3125 2764 3126
rect 2758 3121 2759 3125
rect 2763 3121 2764 3125
rect 2758 3120 2764 3121
rect 2918 3125 2924 3126
rect 2918 3121 2919 3125
rect 2923 3121 2924 3125
rect 2918 3120 2924 3121
rect 3078 3125 3084 3126
rect 3078 3121 3079 3125
rect 3083 3121 3084 3125
rect 3078 3120 3084 3121
rect 3230 3125 3236 3126
rect 3230 3121 3231 3125
rect 3235 3121 3236 3125
rect 3230 3120 3236 3121
rect 3366 3125 3372 3126
rect 3366 3121 3367 3125
rect 3371 3121 3372 3125
rect 3366 3120 3372 3121
rect 3462 3124 3468 3125
rect 3462 3120 3463 3124
rect 3467 3120 3468 3124
rect 1806 3119 1812 3120
rect 3462 3119 3468 3120
rect 366 3117 372 3118
rect 110 3116 116 3117
rect 110 3112 111 3116
rect 115 3112 116 3116
rect 366 3113 367 3117
rect 371 3113 372 3117
rect 366 3112 372 3113
rect 486 3117 492 3118
rect 486 3113 487 3117
rect 491 3113 492 3117
rect 486 3112 492 3113
rect 606 3117 612 3118
rect 606 3113 607 3117
rect 611 3113 612 3117
rect 606 3112 612 3113
rect 726 3117 732 3118
rect 726 3113 727 3117
rect 731 3113 732 3117
rect 726 3112 732 3113
rect 846 3117 852 3118
rect 846 3113 847 3117
rect 851 3113 852 3117
rect 846 3112 852 3113
rect 966 3117 972 3118
rect 966 3113 967 3117
rect 971 3113 972 3117
rect 966 3112 972 3113
rect 1078 3117 1084 3118
rect 1078 3113 1079 3117
rect 1083 3113 1084 3117
rect 1078 3112 1084 3113
rect 1198 3117 1204 3118
rect 1198 3113 1199 3117
rect 1203 3113 1204 3117
rect 1198 3112 1204 3113
rect 1318 3117 1324 3118
rect 1318 3113 1319 3117
rect 1323 3113 1324 3117
rect 1318 3112 1324 3113
rect 1766 3116 1772 3117
rect 1766 3112 1767 3116
rect 1771 3112 1772 3116
rect 110 3111 116 3112
rect 1766 3111 1772 3112
rect 1879 3107 1885 3108
rect 1879 3103 1880 3107
rect 1884 3106 1885 3107
rect 1910 3107 1916 3108
rect 1910 3106 1911 3107
rect 1884 3104 1911 3106
rect 1884 3103 1885 3104
rect 1879 3102 1885 3103
rect 1910 3103 1911 3104
rect 1915 3103 1916 3107
rect 1910 3102 1916 3103
rect 2055 3107 2061 3108
rect 2055 3103 2056 3107
rect 2060 3106 2061 3107
rect 2255 3107 2261 3108
rect 2060 3104 2250 3106
rect 2060 3103 2061 3104
rect 2055 3102 2061 3103
rect 415 3099 424 3100
rect 415 3095 416 3099
rect 423 3095 424 3099
rect 415 3094 424 3095
rect 438 3099 444 3100
rect 438 3095 439 3099
rect 443 3098 444 3099
rect 535 3099 541 3100
rect 535 3098 536 3099
rect 443 3096 536 3098
rect 443 3095 444 3096
rect 438 3094 444 3095
rect 535 3095 536 3096
rect 540 3095 541 3099
rect 535 3094 541 3095
rect 558 3099 564 3100
rect 558 3095 559 3099
rect 563 3098 564 3099
rect 655 3099 661 3100
rect 655 3098 656 3099
rect 563 3096 656 3098
rect 563 3095 564 3096
rect 558 3094 564 3095
rect 655 3095 656 3096
rect 660 3095 661 3099
rect 655 3094 661 3095
rect 678 3099 684 3100
rect 678 3095 679 3099
rect 683 3098 684 3099
rect 775 3099 781 3100
rect 775 3098 776 3099
rect 683 3096 776 3098
rect 683 3095 684 3096
rect 678 3094 684 3095
rect 775 3095 776 3096
rect 780 3095 781 3099
rect 775 3094 781 3095
rect 895 3099 901 3100
rect 895 3095 896 3099
rect 900 3098 901 3099
rect 918 3099 924 3100
rect 900 3096 914 3098
rect 900 3095 901 3096
rect 895 3094 901 3095
rect 686 3091 692 3092
rect 686 3090 687 3091
rect 504 3088 687 3090
rect 487 3083 493 3084
rect 487 3079 488 3083
rect 492 3082 493 3083
rect 504 3082 506 3088
rect 686 3087 687 3088
rect 691 3087 692 3091
rect 912 3090 914 3096
rect 918 3095 919 3099
rect 923 3098 924 3099
rect 1015 3099 1021 3100
rect 1015 3098 1016 3099
rect 923 3096 1016 3098
rect 923 3095 924 3096
rect 918 3094 924 3095
rect 1015 3095 1016 3096
rect 1020 3095 1021 3099
rect 1015 3094 1021 3095
rect 1038 3099 1044 3100
rect 1038 3095 1039 3099
rect 1043 3098 1044 3099
rect 1127 3099 1133 3100
rect 1127 3098 1128 3099
rect 1043 3096 1128 3098
rect 1043 3095 1044 3096
rect 1038 3094 1044 3095
rect 1127 3095 1128 3096
rect 1132 3095 1133 3099
rect 1127 3094 1133 3095
rect 1150 3099 1156 3100
rect 1150 3095 1151 3099
rect 1155 3098 1156 3099
rect 1247 3099 1253 3100
rect 1247 3098 1248 3099
rect 1155 3096 1248 3098
rect 1155 3095 1156 3096
rect 1150 3094 1156 3095
rect 1247 3095 1248 3096
rect 1252 3095 1253 3099
rect 1247 3094 1253 3095
rect 1270 3099 1276 3100
rect 1270 3095 1271 3099
rect 1275 3098 1276 3099
rect 1367 3099 1373 3100
rect 1367 3098 1368 3099
rect 1275 3096 1368 3098
rect 1275 3095 1276 3096
rect 1270 3094 1276 3095
rect 1367 3095 1368 3096
rect 1372 3095 1373 3099
rect 2248 3098 2250 3104
rect 2255 3103 2256 3107
rect 2260 3106 2261 3107
rect 2270 3107 2276 3108
rect 2270 3106 2271 3107
rect 2260 3104 2271 3106
rect 2260 3103 2261 3104
rect 2255 3102 2261 3103
rect 2270 3103 2271 3104
rect 2275 3103 2276 3107
rect 2270 3102 2276 3103
rect 2278 3107 2284 3108
rect 2278 3103 2279 3107
rect 2283 3106 2284 3107
rect 2447 3107 2453 3108
rect 2447 3106 2448 3107
rect 2283 3104 2448 3106
rect 2283 3103 2284 3104
rect 2278 3102 2284 3103
rect 2447 3103 2448 3104
rect 2452 3103 2453 3107
rect 2447 3102 2453 3103
rect 2631 3107 2637 3108
rect 2631 3103 2632 3107
rect 2636 3106 2637 3107
rect 2742 3107 2748 3108
rect 2636 3104 2738 3106
rect 2636 3103 2637 3104
rect 2631 3102 2637 3103
rect 2286 3099 2292 3100
rect 2286 3098 2287 3099
rect 2248 3096 2287 3098
rect 1367 3094 1373 3095
rect 2286 3095 2287 3096
rect 2291 3095 2292 3099
rect 2736 3098 2738 3104
rect 2742 3103 2743 3107
rect 2747 3106 2748 3107
rect 2807 3107 2813 3108
rect 2807 3106 2808 3107
rect 2747 3104 2808 3106
rect 2747 3103 2748 3104
rect 2742 3102 2748 3103
rect 2807 3103 2808 3104
rect 2812 3103 2813 3107
rect 2807 3102 2813 3103
rect 2966 3107 2973 3108
rect 2966 3103 2967 3107
rect 2972 3103 2973 3107
rect 2966 3102 2973 3103
rect 2990 3107 2996 3108
rect 2990 3103 2991 3107
rect 2995 3106 2996 3107
rect 3127 3107 3133 3108
rect 3127 3106 3128 3107
rect 2995 3104 3128 3106
rect 2995 3103 2996 3104
rect 2990 3102 2996 3103
rect 3127 3103 3128 3104
rect 3132 3103 3133 3107
rect 3127 3102 3133 3103
rect 3150 3107 3156 3108
rect 3150 3103 3151 3107
rect 3155 3106 3156 3107
rect 3279 3107 3285 3108
rect 3279 3106 3280 3107
rect 3155 3104 3280 3106
rect 3155 3103 3156 3104
rect 3150 3102 3156 3103
rect 3279 3103 3280 3104
rect 3284 3103 3285 3107
rect 3279 3102 3285 3103
rect 3406 3107 3412 3108
rect 3406 3103 3407 3107
rect 3411 3106 3412 3107
rect 3415 3107 3421 3108
rect 3415 3106 3416 3107
rect 3411 3104 3416 3106
rect 3411 3103 3412 3104
rect 3406 3102 3412 3103
rect 3415 3103 3416 3104
rect 3420 3103 3421 3107
rect 3415 3102 3421 3103
rect 3079 3099 3085 3100
rect 3079 3098 3080 3099
rect 2736 3096 3080 3098
rect 2286 3094 2292 3095
rect 3079 3095 3080 3096
rect 3084 3095 3085 3099
rect 3079 3094 3085 3095
rect 1134 3091 1140 3092
rect 1134 3090 1135 3091
rect 912 3088 1135 3090
rect 686 3086 692 3087
rect 1134 3087 1135 3088
rect 1139 3087 1140 3091
rect 1134 3086 1140 3087
rect 1879 3087 1885 3088
rect 492 3080 506 3082
rect 510 3083 516 3084
rect 492 3079 493 3080
rect 487 3078 493 3079
rect 510 3079 511 3083
rect 515 3082 516 3083
rect 575 3083 581 3084
rect 575 3082 576 3083
rect 515 3080 576 3082
rect 515 3079 516 3080
rect 510 3078 516 3079
rect 575 3079 576 3080
rect 580 3079 581 3083
rect 575 3078 581 3079
rect 598 3083 604 3084
rect 598 3079 599 3083
rect 603 3082 604 3083
rect 663 3083 669 3084
rect 663 3082 664 3083
rect 603 3080 664 3082
rect 603 3079 604 3080
rect 598 3078 604 3079
rect 663 3079 664 3080
rect 668 3079 669 3083
rect 663 3078 669 3079
rect 686 3083 692 3084
rect 686 3079 687 3083
rect 691 3082 692 3083
rect 751 3083 757 3084
rect 751 3082 752 3083
rect 691 3080 752 3082
rect 691 3079 692 3080
rect 686 3078 692 3079
rect 751 3079 752 3080
rect 756 3079 757 3083
rect 751 3078 757 3079
rect 774 3083 780 3084
rect 774 3079 775 3083
rect 779 3082 780 3083
rect 839 3083 845 3084
rect 839 3082 840 3083
rect 779 3080 840 3082
rect 779 3079 780 3080
rect 774 3078 780 3079
rect 839 3079 840 3080
rect 844 3079 845 3083
rect 839 3078 845 3079
rect 926 3083 933 3084
rect 926 3079 927 3083
rect 932 3079 933 3083
rect 926 3078 933 3079
rect 950 3083 956 3084
rect 950 3079 951 3083
rect 955 3082 956 3083
rect 1015 3083 1021 3084
rect 1015 3082 1016 3083
rect 955 3080 1016 3082
rect 955 3079 956 3080
rect 950 3078 956 3079
rect 1015 3079 1016 3080
rect 1020 3079 1021 3083
rect 1015 3078 1021 3079
rect 1038 3083 1044 3084
rect 1038 3079 1039 3083
rect 1043 3082 1044 3083
rect 1103 3083 1109 3084
rect 1103 3082 1104 3083
rect 1043 3080 1104 3082
rect 1043 3079 1044 3080
rect 1038 3078 1044 3079
rect 1103 3079 1104 3080
rect 1108 3079 1109 3083
rect 1103 3078 1109 3079
rect 1126 3083 1132 3084
rect 1126 3079 1127 3083
rect 1131 3082 1132 3083
rect 1191 3083 1197 3084
rect 1191 3082 1192 3083
rect 1131 3080 1192 3082
rect 1131 3079 1132 3080
rect 1126 3078 1132 3079
rect 1191 3079 1192 3080
rect 1196 3079 1197 3083
rect 1879 3083 1880 3087
rect 1884 3086 1885 3087
rect 1894 3087 1900 3088
rect 1894 3086 1895 3087
rect 1884 3084 1895 3086
rect 1884 3083 1885 3084
rect 1879 3082 1885 3083
rect 1894 3083 1895 3084
rect 1899 3083 1900 3087
rect 1894 3082 1900 3083
rect 1902 3087 1908 3088
rect 1902 3083 1903 3087
rect 1907 3086 1908 3087
rect 2007 3087 2013 3088
rect 2007 3086 2008 3087
rect 1907 3084 2008 3086
rect 1907 3083 1908 3084
rect 1902 3082 1908 3083
rect 2007 3083 2008 3084
rect 2012 3083 2013 3087
rect 2007 3082 2013 3083
rect 2030 3087 2036 3088
rect 2030 3083 2031 3087
rect 2035 3086 2036 3087
rect 2167 3087 2173 3088
rect 2167 3086 2168 3087
rect 2035 3084 2168 3086
rect 2035 3083 2036 3084
rect 2030 3082 2036 3083
rect 2167 3083 2168 3084
rect 2172 3083 2173 3087
rect 2167 3082 2173 3083
rect 2190 3087 2196 3088
rect 2190 3083 2191 3087
rect 2195 3086 2196 3087
rect 2343 3087 2349 3088
rect 2343 3086 2344 3087
rect 2195 3084 2344 3086
rect 2195 3083 2196 3084
rect 2190 3082 2196 3083
rect 2343 3083 2344 3084
rect 2348 3083 2349 3087
rect 2343 3082 2349 3083
rect 2535 3087 2541 3088
rect 2535 3083 2536 3087
rect 2540 3086 2541 3087
rect 2550 3087 2556 3088
rect 2550 3086 2551 3087
rect 2540 3084 2551 3086
rect 2540 3083 2541 3084
rect 2535 3082 2541 3083
rect 2550 3083 2551 3084
rect 2555 3083 2556 3087
rect 2550 3082 2556 3083
rect 2558 3087 2564 3088
rect 2558 3083 2559 3087
rect 2563 3086 2564 3087
rect 2743 3087 2749 3088
rect 2743 3086 2744 3087
rect 2563 3084 2744 3086
rect 2563 3083 2564 3084
rect 2558 3082 2564 3083
rect 2743 3083 2744 3084
rect 2748 3083 2749 3087
rect 2743 3082 2749 3083
rect 2766 3087 2772 3088
rect 2766 3083 2767 3087
rect 2771 3086 2772 3087
rect 2967 3087 2973 3088
rect 2967 3086 2968 3087
rect 2771 3084 2968 3086
rect 2771 3083 2772 3084
rect 2766 3082 2772 3083
rect 2967 3083 2968 3084
rect 2972 3083 2973 3087
rect 2967 3082 2973 3083
rect 2990 3087 2996 3088
rect 2990 3083 2991 3087
rect 2995 3086 2996 3087
rect 3199 3087 3205 3088
rect 3199 3086 3200 3087
rect 2995 3084 3200 3086
rect 2995 3083 2996 3084
rect 2990 3082 2996 3083
rect 3199 3083 3200 3084
rect 3204 3083 3205 3087
rect 3199 3082 3205 3083
rect 3415 3087 3421 3088
rect 3415 3083 3416 3087
rect 3420 3086 3421 3087
rect 3430 3087 3436 3088
rect 3430 3086 3431 3087
rect 3420 3084 3431 3086
rect 3420 3083 3421 3084
rect 3415 3082 3421 3083
rect 3430 3083 3431 3084
rect 3435 3083 3436 3087
rect 3430 3082 3436 3083
rect 1191 3078 1197 3079
rect 1806 3072 1812 3073
rect 3462 3072 3468 3073
rect 110 3068 116 3069
rect 1766 3068 1772 3069
rect 110 3064 111 3068
rect 115 3064 116 3068
rect 110 3063 116 3064
rect 438 3067 444 3068
rect 438 3063 439 3067
rect 443 3063 444 3067
rect 438 3062 444 3063
rect 526 3067 532 3068
rect 526 3063 527 3067
rect 531 3063 532 3067
rect 526 3062 532 3063
rect 614 3067 620 3068
rect 614 3063 615 3067
rect 619 3063 620 3067
rect 614 3062 620 3063
rect 702 3067 708 3068
rect 702 3063 703 3067
rect 707 3063 708 3067
rect 702 3062 708 3063
rect 790 3067 796 3068
rect 790 3063 791 3067
rect 795 3063 796 3067
rect 790 3062 796 3063
rect 878 3067 884 3068
rect 878 3063 879 3067
rect 883 3063 884 3067
rect 878 3062 884 3063
rect 966 3067 972 3068
rect 966 3063 967 3067
rect 971 3063 972 3067
rect 966 3062 972 3063
rect 1054 3067 1060 3068
rect 1054 3063 1055 3067
rect 1059 3063 1060 3067
rect 1054 3062 1060 3063
rect 1142 3067 1148 3068
rect 1142 3063 1143 3067
rect 1147 3063 1148 3067
rect 1766 3064 1767 3068
rect 1771 3064 1772 3068
rect 1806 3068 1807 3072
rect 1811 3068 1812 3072
rect 1806 3067 1812 3068
rect 1830 3071 1836 3072
rect 1830 3067 1831 3071
rect 1835 3067 1836 3071
rect 1830 3066 1836 3067
rect 1958 3071 1964 3072
rect 1958 3067 1959 3071
rect 1963 3067 1964 3071
rect 1958 3066 1964 3067
rect 2118 3071 2124 3072
rect 2118 3067 2119 3071
rect 2123 3067 2124 3071
rect 2118 3066 2124 3067
rect 2294 3071 2300 3072
rect 2294 3067 2295 3071
rect 2299 3067 2300 3071
rect 2294 3066 2300 3067
rect 2486 3071 2492 3072
rect 2486 3067 2487 3071
rect 2491 3067 2492 3071
rect 2486 3066 2492 3067
rect 2694 3071 2700 3072
rect 2694 3067 2695 3071
rect 2699 3067 2700 3071
rect 2694 3066 2700 3067
rect 2918 3071 2924 3072
rect 2918 3067 2919 3071
rect 2923 3067 2924 3071
rect 2918 3066 2924 3067
rect 3150 3071 3156 3072
rect 3150 3067 3151 3071
rect 3155 3067 3156 3071
rect 3150 3066 3156 3067
rect 3366 3071 3372 3072
rect 3366 3067 3367 3071
rect 3371 3067 3372 3071
rect 3462 3068 3463 3072
rect 3467 3068 3468 3072
rect 3462 3067 3468 3068
rect 3366 3066 3372 3067
rect 1766 3063 1772 3064
rect 1902 3063 1908 3064
rect 1142 3062 1148 3063
rect 510 3059 516 3060
rect 510 3055 511 3059
rect 515 3055 516 3059
rect 510 3054 516 3055
rect 598 3059 604 3060
rect 598 3055 599 3059
rect 603 3055 604 3059
rect 598 3054 604 3055
rect 686 3059 692 3060
rect 686 3055 687 3059
rect 691 3055 692 3059
rect 686 3054 692 3055
rect 774 3059 780 3060
rect 774 3055 775 3059
rect 779 3055 780 3059
rect 950 3059 956 3060
rect 774 3054 780 3055
rect 862 3055 868 3056
rect 110 3051 116 3052
rect 110 3047 111 3051
rect 115 3047 116 3051
rect 862 3051 863 3055
rect 867 3051 868 3055
rect 950 3055 951 3059
rect 955 3055 956 3059
rect 950 3054 956 3055
rect 1038 3059 1044 3060
rect 1038 3055 1039 3059
rect 1043 3055 1044 3059
rect 1038 3054 1044 3055
rect 1126 3059 1132 3060
rect 1126 3055 1127 3059
rect 1131 3055 1132 3059
rect 1126 3054 1132 3055
rect 1134 3059 1140 3060
rect 1134 3055 1135 3059
rect 1139 3058 1140 3059
rect 1902 3059 1903 3063
rect 1907 3059 1908 3063
rect 1902 3058 1908 3059
rect 2030 3063 2036 3064
rect 2030 3059 2031 3063
rect 2035 3059 2036 3063
rect 2030 3058 2036 3059
rect 2190 3063 2196 3064
rect 2190 3059 2191 3063
rect 2195 3059 2196 3063
rect 2558 3063 2564 3064
rect 2190 3058 2196 3059
rect 2200 3060 2337 3062
rect 1139 3056 1185 3058
rect 1139 3055 1140 3056
rect 1134 3054 1140 3055
rect 1806 3055 1812 3056
rect 862 3050 868 3051
rect 1766 3051 1772 3052
rect 110 3046 116 3047
rect 438 3048 444 3049
rect 438 3044 439 3048
rect 443 3044 444 3048
rect 438 3043 444 3044
rect 526 3048 532 3049
rect 526 3044 527 3048
rect 531 3044 532 3048
rect 526 3043 532 3044
rect 614 3048 620 3049
rect 614 3044 615 3048
rect 619 3044 620 3048
rect 614 3043 620 3044
rect 702 3048 708 3049
rect 702 3044 703 3048
rect 707 3044 708 3048
rect 702 3043 708 3044
rect 790 3048 796 3049
rect 790 3044 791 3048
rect 795 3044 796 3048
rect 790 3043 796 3044
rect 878 3048 884 3049
rect 878 3044 879 3048
rect 883 3044 884 3048
rect 878 3043 884 3044
rect 966 3048 972 3049
rect 966 3044 967 3048
rect 971 3044 972 3048
rect 966 3043 972 3044
rect 1054 3048 1060 3049
rect 1054 3044 1055 3048
rect 1059 3044 1060 3048
rect 1054 3043 1060 3044
rect 1142 3048 1148 3049
rect 1142 3044 1143 3048
rect 1147 3044 1148 3048
rect 1766 3047 1767 3051
rect 1771 3047 1772 3051
rect 1806 3051 1807 3055
rect 1811 3051 1812 3055
rect 2182 3055 2188 3056
rect 1806 3050 1812 3051
rect 1830 3052 1836 3053
rect 1830 3048 1831 3052
rect 1835 3048 1836 3052
rect 1830 3047 1836 3048
rect 1958 3052 1964 3053
rect 1958 3048 1959 3052
rect 1963 3048 1964 3052
rect 1958 3047 1964 3048
rect 2118 3052 2124 3053
rect 2118 3048 2119 3052
rect 2123 3048 2124 3052
rect 2182 3051 2183 3055
rect 2187 3054 2188 3055
rect 2200 3054 2202 3060
rect 2558 3059 2559 3063
rect 2563 3059 2564 3063
rect 2558 3058 2564 3059
rect 2766 3063 2772 3064
rect 2766 3059 2767 3063
rect 2771 3059 2772 3063
rect 2766 3058 2772 3059
rect 2990 3063 2996 3064
rect 2990 3059 2991 3063
rect 2995 3059 2996 3063
rect 2990 3058 2996 3059
rect 3079 3063 3085 3064
rect 3079 3059 3080 3063
rect 3084 3062 3085 3063
rect 3084 3060 3193 3062
rect 3084 3059 3085 3060
rect 3079 3058 3085 3059
rect 2187 3052 2202 3054
rect 3430 3055 3436 3056
rect 2294 3052 2300 3053
rect 2187 3051 2188 3052
rect 2182 3050 2188 3051
rect 2118 3047 2124 3048
rect 2294 3048 2295 3052
rect 2299 3048 2300 3052
rect 2294 3047 2300 3048
rect 2486 3052 2492 3053
rect 2486 3048 2487 3052
rect 2491 3048 2492 3052
rect 2486 3047 2492 3048
rect 2694 3052 2700 3053
rect 2694 3048 2695 3052
rect 2699 3048 2700 3052
rect 2694 3047 2700 3048
rect 2918 3052 2924 3053
rect 2918 3048 2919 3052
rect 2923 3048 2924 3052
rect 2918 3047 2924 3048
rect 3150 3052 3156 3053
rect 3150 3048 3151 3052
rect 3155 3048 3156 3052
rect 3150 3047 3156 3048
rect 3366 3052 3372 3053
rect 3366 3048 3367 3052
rect 3371 3048 3372 3052
rect 3430 3051 3431 3055
rect 3435 3054 3436 3055
rect 3440 3054 3442 3057
rect 3435 3052 3442 3054
rect 3462 3055 3468 3056
rect 3435 3051 3436 3052
rect 3430 3050 3436 3051
rect 3462 3051 3463 3055
rect 3467 3051 3468 3055
rect 3462 3050 3468 3051
rect 3366 3047 3372 3048
rect 1766 3046 1772 3047
rect 1142 3043 1148 3044
rect 2550 2999 2556 3000
rect 502 2996 508 2997
rect 110 2993 116 2994
rect 110 2989 111 2993
rect 115 2989 116 2993
rect 502 2992 503 2996
rect 507 2992 508 2996
rect 502 2991 508 2992
rect 590 2996 596 2997
rect 590 2992 591 2996
rect 595 2992 596 2996
rect 590 2991 596 2992
rect 678 2996 684 2997
rect 678 2992 679 2996
rect 683 2992 684 2996
rect 678 2991 684 2992
rect 766 2996 772 2997
rect 766 2992 767 2996
rect 771 2992 772 2996
rect 766 2991 772 2992
rect 854 2996 860 2997
rect 854 2992 855 2996
rect 859 2992 860 2996
rect 854 2991 860 2992
rect 942 2996 948 2997
rect 942 2992 943 2996
rect 947 2992 948 2996
rect 942 2991 948 2992
rect 1030 2996 1036 2997
rect 1030 2992 1031 2996
rect 1035 2992 1036 2996
rect 1030 2991 1036 2992
rect 1118 2996 1124 2997
rect 1118 2992 1119 2996
rect 1123 2992 1124 2996
rect 1118 2991 1124 2992
rect 1206 2996 1212 2997
rect 1206 2992 1207 2996
rect 1211 2992 1212 2996
rect 1206 2991 1212 2992
rect 1294 2996 1300 2997
rect 1294 2992 1295 2996
rect 1299 2992 1300 2996
rect 2550 2995 2551 2999
rect 2555 2998 2556 2999
rect 2555 2996 3066 2998
rect 2555 2995 2556 2996
rect 2550 2994 2556 2995
rect 1294 2991 1300 2992
rect 1766 2993 1772 2994
rect 110 2988 116 2989
rect 1766 2989 1767 2993
rect 1771 2989 1772 2993
rect 1830 2992 1836 2993
rect 1766 2988 1772 2989
rect 1806 2989 1812 2990
rect 574 2987 580 2988
rect 574 2983 575 2987
rect 579 2983 580 2987
rect 574 2982 580 2983
rect 662 2987 668 2988
rect 662 2983 663 2987
rect 667 2983 668 2987
rect 662 2982 668 2983
rect 750 2987 756 2988
rect 750 2983 751 2987
rect 755 2983 756 2987
rect 750 2982 756 2983
rect 758 2987 764 2988
rect 758 2983 759 2987
rect 763 2986 764 2987
rect 846 2987 852 2988
rect 763 2984 809 2986
rect 763 2983 764 2984
rect 758 2982 764 2983
rect 846 2983 847 2987
rect 851 2986 852 2987
rect 934 2987 940 2988
rect 851 2984 897 2986
rect 851 2983 852 2984
rect 846 2982 852 2983
rect 934 2983 935 2987
rect 939 2986 940 2987
rect 1022 2987 1028 2988
rect 939 2984 985 2986
rect 939 2983 940 2984
rect 934 2982 940 2983
rect 1022 2983 1023 2987
rect 1027 2986 1028 2987
rect 1190 2987 1196 2988
rect 1027 2984 1073 2986
rect 1027 2983 1028 2984
rect 1022 2982 1028 2983
rect 1190 2983 1191 2987
rect 1195 2983 1196 2987
rect 1190 2982 1196 2983
rect 1278 2987 1284 2988
rect 1278 2983 1279 2987
rect 1283 2983 1284 2987
rect 1278 2982 1284 2983
rect 1286 2987 1292 2988
rect 1286 2983 1287 2987
rect 1291 2986 1292 2987
rect 1291 2984 1337 2986
rect 1806 2985 1807 2989
rect 1811 2985 1812 2989
rect 1830 2988 1831 2992
rect 1835 2988 1836 2992
rect 1830 2987 1836 2988
rect 1918 2992 1924 2993
rect 1918 2988 1919 2992
rect 1923 2988 1924 2992
rect 1918 2987 1924 2988
rect 2030 2992 2036 2993
rect 2030 2988 2031 2992
rect 2035 2988 2036 2992
rect 2030 2987 2036 2988
rect 2142 2992 2148 2993
rect 2142 2988 2143 2992
rect 2147 2988 2148 2992
rect 2142 2987 2148 2988
rect 2246 2992 2252 2993
rect 2246 2988 2247 2992
rect 2251 2988 2252 2992
rect 2246 2987 2252 2988
rect 2358 2992 2364 2993
rect 2358 2988 2359 2992
rect 2363 2988 2364 2992
rect 2358 2987 2364 2988
rect 2478 2992 2484 2993
rect 2478 2988 2479 2992
rect 2483 2988 2484 2992
rect 2478 2987 2484 2988
rect 2622 2992 2628 2993
rect 2622 2988 2623 2992
rect 2627 2988 2628 2992
rect 2622 2987 2628 2988
rect 2790 2992 2796 2993
rect 2790 2988 2791 2992
rect 2795 2988 2796 2992
rect 2790 2987 2796 2988
rect 2982 2992 2988 2993
rect 2982 2988 2983 2992
rect 2987 2988 2988 2992
rect 2982 2987 2988 2988
rect 1806 2984 1812 2985
rect 1291 2983 1292 2984
rect 1286 2982 1292 2983
rect 1894 2983 1900 2984
rect 1894 2979 1895 2983
rect 1899 2979 1900 2983
rect 1894 2978 1900 2979
rect 1910 2983 1916 2984
rect 1910 2979 1911 2983
rect 1915 2982 1916 2983
rect 2023 2983 2029 2984
rect 1915 2980 1961 2982
rect 1915 2979 1916 2980
rect 1910 2978 1916 2979
rect 2023 2979 2024 2983
rect 2028 2982 2029 2983
rect 2214 2983 2220 2984
rect 2028 2980 2073 2982
rect 2028 2979 2029 2980
rect 2023 2978 2029 2979
rect 2214 2979 2215 2983
rect 2219 2979 2220 2983
rect 2214 2978 2220 2979
rect 2318 2983 2324 2984
rect 2318 2979 2319 2983
rect 2323 2979 2324 2983
rect 2318 2978 2324 2979
rect 2430 2983 2436 2984
rect 2430 2979 2431 2983
rect 2435 2979 2436 2983
rect 2430 2978 2436 2979
rect 2550 2983 2556 2984
rect 2550 2979 2551 2983
rect 2555 2979 2556 2983
rect 2550 2978 2556 2979
rect 2694 2983 2700 2984
rect 2694 2979 2695 2983
rect 2699 2979 2700 2983
rect 2694 2978 2700 2979
rect 2862 2983 2868 2984
rect 2862 2979 2863 2983
rect 2867 2979 2868 2983
rect 2862 2978 2868 2979
rect 3054 2983 3060 2984
rect 3054 2979 3055 2983
rect 3059 2979 3060 2983
rect 3064 2982 3066 2996
rect 3182 2992 3188 2993
rect 3182 2988 3183 2992
rect 3187 2988 3188 2992
rect 3182 2987 3188 2988
rect 3366 2992 3372 2993
rect 3366 2988 3367 2992
rect 3371 2988 3372 2992
rect 3366 2987 3372 2988
rect 3462 2989 3468 2990
rect 3462 2985 3463 2989
rect 3467 2985 3468 2989
rect 3462 2984 3468 2985
rect 3438 2983 3444 2984
rect 3064 2980 3225 2982
rect 3054 2978 3060 2979
rect 3438 2979 3439 2983
rect 3443 2979 3444 2983
rect 3438 2978 3444 2979
rect 502 2977 508 2978
rect 110 2976 116 2977
rect 110 2972 111 2976
rect 115 2972 116 2976
rect 502 2973 503 2977
rect 507 2973 508 2977
rect 502 2972 508 2973
rect 590 2977 596 2978
rect 590 2973 591 2977
rect 595 2973 596 2977
rect 590 2972 596 2973
rect 678 2977 684 2978
rect 678 2973 679 2977
rect 683 2973 684 2977
rect 678 2972 684 2973
rect 766 2977 772 2978
rect 766 2973 767 2977
rect 771 2973 772 2977
rect 766 2972 772 2973
rect 854 2977 860 2978
rect 854 2973 855 2977
rect 859 2973 860 2977
rect 854 2972 860 2973
rect 942 2977 948 2978
rect 942 2973 943 2977
rect 947 2973 948 2977
rect 942 2972 948 2973
rect 1030 2977 1036 2978
rect 1030 2973 1031 2977
rect 1035 2973 1036 2977
rect 1030 2972 1036 2973
rect 1118 2977 1124 2978
rect 1118 2973 1119 2977
rect 1123 2973 1124 2977
rect 1118 2972 1124 2973
rect 1206 2977 1212 2978
rect 1206 2973 1207 2977
rect 1211 2973 1212 2977
rect 1206 2972 1212 2973
rect 1294 2977 1300 2978
rect 1294 2973 1295 2977
rect 1299 2973 1300 2977
rect 1294 2972 1300 2973
rect 1766 2976 1772 2977
rect 1766 2972 1767 2976
rect 1771 2972 1772 2976
rect 1830 2973 1836 2974
rect 110 2971 116 2972
rect 1766 2971 1772 2972
rect 1806 2972 1812 2973
rect 1806 2968 1807 2972
rect 1811 2968 1812 2972
rect 1830 2969 1831 2973
rect 1835 2969 1836 2973
rect 1830 2968 1836 2969
rect 1918 2973 1924 2974
rect 1918 2969 1919 2973
rect 1923 2969 1924 2973
rect 1918 2968 1924 2969
rect 2030 2973 2036 2974
rect 2030 2969 2031 2973
rect 2035 2969 2036 2973
rect 2030 2968 2036 2969
rect 2142 2973 2148 2974
rect 2142 2969 2143 2973
rect 2147 2969 2148 2973
rect 2142 2968 2148 2969
rect 2246 2973 2252 2974
rect 2246 2969 2247 2973
rect 2251 2969 2252 2973
rect 2246 2968 2252 2969
rect 2358 2973 2364 2974
rect 2358 2969 2359 2973
rect 2363 2969 2364 2973
rect 2358 2968 2364 2969
rect 2478 2973 2484 2974
rect 2478 2969 2479 2973
rect 2483 2969 2484 2973
rect 2478 2968 2484 2969
rect 2622 2973 2628 2974
rect 2622 2969 2623 2973
rect 2627 2969 2628 2973
rect 2622 2968 2628 2969
rect 2790 2973 2796 2974
rect 2790 2969 2791 2973
rect 2795 2969 2796 2973
rect 2790 2968 2796 2969
rect 2982 2973 2988 2974
rect 2982 2969 2983 2973
rect 2987 2969 2988 2973
rect 2982 2968 2988 2969
rect 3182 2973 3188 2974
rect 3182 2969 3183 2973
rect 3187 2969 3188 2973
rect 3182 2968 3188 2969
rect 3366 2973 3372 2974
rect 3366 2969 3367 2973
rect 3371 2969 3372 2973
rect 3366 2968 3372 2969
rect 3462 2972 3468 2973
rect 3462 2968 3463 2972
rect 3467 2968 3468 2972
rect 1806 2967 1812 2968
rect 3462 2967 3468 2968
rect 551 2959 557 2960
rect 551 2955 552 2959
rect 556 2958 557 2959
rect 574 2959 580 2960
rect 556 2956 570 2958
rect 556 2955 557 2956
rect 551 2954 557 2955
rect 568 2950 570 2956
rect 574 2955 575 2959
rect 579 2958 580 2959
rect 639 2959 645 2960
rect 639 2958 640 2959
rect 579 2956 640 2958
rect 579 2955 580 2956
rect 574 2954 580 2955
rect 639 2955 640 2956
rect 644 2955 645 2959
rect 639 2954 645 2955
rect 662 2959 668 2960
rect 662 2955 663 2959
rect 667 2958 668 2959
rect 727 2959 733 2960
rect 727 2958 728 2959
rect 667 2956 728 2958
rect 667 2955 668 2956
rect 662 2954 668 2955
rect 727 2955 728 2956
rect 732 2955 733 2959
rect 727 2954 733 2955
rect 815 2959 821 2960
rect 815 2955 816 2959
rect 820 2958 821 2959
rect 846 2959 852 2960
rect 846 2958 847 2959
rect 820 2956 847 2958
rect 820 2955 821 2956
rect 815 2954 821 2955
rect 846 2955 847 2956
rect 851 2955 852 2959
rect 846 2954 852 2955
rect 862 2959 868 2960
rect 862 2955 863 2959
rect 867 2958 868 2959
rect 903 2959 909 2960
rect 903 2958 904 2959
rect 867 2956 904 2958
rect 867 2955 868 2956
rect 862 2954 868 2955
rect 903 2955 904 2956
rect 908 2955 909 2959
rect 903 2954 909 2955
rect 991 2959 997 2960
rect 991 2955 992 2959
rect 996 2958 997 2959
rect 1022 2959 1028 2960
rect 1022 2958 1023 2959
rect 996 2956 1023 2958
rect 996 2955 997 2956
rect 991 2954 997 2955
rect 1022 2955 1023 2956
rect 1027 2955 1028 2959
rect 1022 2954 1028 2955
rect 1079 2959 1085 2960
rect 1079 2955 1080 2959
rect 1084 2958 1085 2959
rect 1166 2959 1173 2960
rect 1084 2956 1162 2958
rect 1084 2955 1085 2956
rect 1079 2954 1085 2955
rect 758 2951 764 2952
rect 758 2950 759 2951
rect 568 2948 759 2950
rect 758 2947 759 2948
rect 763 2947 764 2951
rect 1160 2950 1162 2956
rect 1166 2955 1167 2959
rect 1172 2955 1173 2959
rect 1166 2954 1173 2955
rect 1190 2959 1196 2960
rect 1190 2955 1191 2959
rect 1195 2958 1196 2959
rect 1255 2959 1261 2960
rect 1255 2958 1256 2959
rect 1195 2956 1256 2958
rect 1195 2955 1196 2956
rect 1190 2954 1196 2955
rect 1255 2955 1256 2956
rect 1260 2955 1261 2959
rect 1255 2954 1261 2955
rect 1278 2959 1284 2960
rect 1278 2955 1279 2959
rect 1283 2958 1284 2959
rect 1343 2959 1349 2960
rect 1343 2958 1344 2959
rect 1283 2956 1344 2958
rect 1283 2955 1284 2956
rect 1278 2954 1284 2955
rect 1343 2955 1344 2956
rect 1348 2955 1349 2959
rect 1343 2954 1349 2955
rect 1879 2955 1885 2956
rect 1286 2951 1292 2952
rect 1286 2950 1287 2951
rect 1160 2948 1287 2950
rect 758 2946 764 2947
rect 1286 2947 1287 2948
rect 1291 2947 1292 2951
rect 1879 2951 1880 2955
rect 1884 2954 1885 2955
rect 1910 2955 1916 2956
rect 1910 2954 1911 2955
rect 1884 2952 1911 2954
rect 1884 2951 1885 2952
rect 1879 2950 1885 2951
rect 1910 2951 1911 2952
rect 1915 2951 1916 2955
rect 1910 2950 1916 2951
rect 1967 2955 1973 2956
rect 1967 2951 1968 2955
rect 1972 2954 1973 2955
rect 2023 2955 2029 2956
rect 2023 2954 2024 2955
rect 1972 2952 2024 2954
rect 1972 2951 1973 2952
rect 1967 2950 1973 2951
rect 2023 2951 2024 2952
rect 2028 2951 2029 2955
rect 2023 2950 2029 2951
rect 2079 2955 2085 2956
rect 2079 2951 2080 2955
rect 2084 2954 2085 2955
rect 2182 2955 2188 2956
rect 2182 2954 2183 2955
rect 2084 2952 2183 2954
rect 2084 2951 2085 2952
rect 2079 2950 2085 2951
rect 2182 2951 2183 2952
rect 2187 2951 2188 2955
rect 2182 2950 2188 2951
rect 2191 2955 2200 2956
rect 2191 2951 2192 2955
rect 2199 2951 2200 2955
rect 2191 2950 2200 2951
rect 2214 2955 2220 2956
rect 2214 2951 2215 2955
rect 2219 2954 2220 2955
rect 2295 2955 2301 2956
rect 2295 2954 2296 2955
rect 2219 2952 2296 2954
rect 2219 2951 2220 2952
rect 2214 2950 2220 2951
rect 2295 2951 2296 2952
rect 2300 2951 2301 2955
rect 2295 2950 2301 2951
rect 2318 2955 2324 2956
rect 2318 2951 2319 2955
rect 2323 2954 2324 2955
rect 2407 2955 2413 2956
rect 2407 2954 2408 2955
rect 2323 2952 2408 2954
rect 2323 2951 2324 2952
rect 2318 2950 2324 2951
rect 2407 2951 2408 2952
rect 2412 2951 2413 2955
rect 2407 2950 2413 2951
rect 2430 2955 2436 2956
rect 2430 2951 2431 2955
rect 2435 2954 2436 2955
rect 2527 2955 2533 2956
rect 2527 2954 2528 2955
rect 2435 2952 2528 2954
rect 2435 2951 2436 2952
rect 2430 2950 2436 2951
rect 2527 2951 2528 2952
rect 2532 2951 2533 2955
rect 2527 2950 2533 2951
rect 2550 2955 2556 2956
rect 2550 2951 2551 2955
rect 2555 2954 2556 2955
rect 2671 2955 2677 2956
rect 2671 2954 2672 2955
rect 2555 2952 2672 2954
rect 2555 2951 2556 2952
rect 2550 2950 2556 2951
rect 2671 2951 2672 2952
rect 2676 2951 2677 2955
rect 2671 2950 2677 2951
rect 2694 2955 2700 2956
rect 2694 2951 2695 2955
rect 2699 2954 2700 2955
rect 2839 2955 2845 2956
rect 2839 2954 2840 2955
rect 2699 2952 2840 2954
rect 2699 2951 2700 2952
rect 2694 2950 2700 2951
rect 2839 2951 2840 2952
rect 2844 2951 2845 2955
rect 2839 2950 2845 2951
rect 2862 2955 2868 2956
rect 2862 2951 2863 2955
rect 2867 2954 2868 2955
rect 3031 2955 3037 2956
rect 3031 2954 3032 2955
rect 2867 2952 3032 2954
rect 2867 2951 2868 2952
rect 2862 2950 2868 2951
rect 3031 2951 3032 2952
rect 3036 2951 3037 2955
rect 3031 2950 3037 2951
rect 3054 2955 3060 2956
rect 3054 2951 3055 2955
rect 3059 2954 3060 2955
rect 3231 2955 3237 2956
rect 3231 2954 3232 2955
rect 3059 2952 3232 2954
rect 3059 2951 3060 2952
rect 3054 2950 3060 2951
rect 3231 2951 3232 2952
rect 3236 2951 3237 2955
rect 3231 2950 3237 2951
rect 3415 2955 3421 2956
rect 3415 2951 3416 2955
rect 3420 2954 3421 2955
rect 3430 2955 3436 2956
rect 3430 2954 3431 2955
rect 3420 2952 3431 2954
rect 3420 2951 3421 2952
rect 3415 2950 3421 2951
rect 3430 2951 3431 2952
rect 3435 2951 3436 2955
rect 3430 2950 3436 2951
rect 1286 2946 1292 2947
rect 798 2943 804 2944
rect 798 2942 799 2943
rect 392 2940 799 2942
rect 375 2935 381 2936
rect 375 2931 376 2935
rect 380 2934 381 2935
rect 392 2934 394 2940
rect 798 2939 799 2940
rect 803 2939 804 2943
rect 1182 2943 1188 2944
rect 1182 2942 1183 2943
rect 798 2938 804 2939
rect 1092 2940 1183 2942
rect 380 2932 394 2934
rect 398 2935 404 2936
rect 380 2931 381 2932
rect 375 2930 381 2931
rect 398 2931 399 2935
rect 403 2934 404 2935
rect 495 2935 501 2936
rect 495 2934 496 2935
rect 403 2932 496 2934
rect 403 2931 404 2932
rect 398 2930 404 2931
rect 495 2931 496 2932
rect 500 2931 501 2935
rect 495 2930 501 2931
rect 518 2935 524 2936
rect 518 2931 519 2935
rect 523 2934 524 2935
rect 623 2935 629 2936
rect 623 2934 624 2935
rect 523 2932 624 2934
rect 523 2931 524 2932
rect 518 2930 524 2931
rect 623 2931 624 2932
rect 628 2931 629 2935
rect 623 2930 629 2931
rect 750 2935 756 2936
rect 750 2931 751 2935
rect 755 2934 756 2935
rect 759 2935 765 2936
rect 759 2934 760 2935
rect 755 2932 760 2934
rect 755 2931 756 2932
rect 750 2930 756 2931
rect 759 2931 760 2932
rect 764 2931 765 2935
rect 759 2930 765 2931
rect 782 2935 788 2936
rect 782 2931 783 2935
rect 787 2934 788 2935
rect 895 2935 901 2936
rect 895 2934 896 2935
rect 787 2932 896 2934
rect 787 2931 788 2932
rect 782 2930 788 2931
rect 895 2931 896 2932
rect 900 2931 901 2935
rect 895 2930 901 2931
rect 1023 2935 1029 2936
rect 1023 2931 1024 2935
rect 1028 2934 1029 2935
rect 1092 2934 1094 2940
rect 1182 2939 1183 2940
rect 1187 2939 1188 2943
rect 1182 2938 1188 2939
rect 1151 2935 1157 2936
rect 1151 2934 1152 2935
rect 1028 2932 1094 2934
rect 1096 2932 1152 2934
rect 1028 2931 1029 2932
rect 1023 2930 1029 2931
rect 110 2920 116 2921
rect 110 2916 111 2920
rect 115 2916 116 2920
rect 110 2915 116 2916
rect 326 2919 332 2920
rect 326 2915 327 2919
rect 331 2915 332 2919
rect 326 2914 332 2915
rect 446 2919 452 2920
rect 446 2915 447 2919
rect 451 2915 452 2919
rect 446 2914 452 2915
rect 574 2919 580 2920
rect 574 2915 575 2919
rect 579 2915 580 2919
rect 574 2914 580 2915
rect 710 2919 716 2920
rect 710 2915 711 2919
rect 715 2915 716 2919
rect 710 2914 716 2915
rect 846 2919 852 2920
rect 846 2915 847 2919
rect 851 2915 852 2919
rect 846 2914 852 2915
rect 974 2919 980 2920
rect 974 2915 975 2919
rect 979 2915 980 2919
rect 974 2914 980 2915
rect 398 2911 404 2912
rect 398 2907 399 2911
rect 403 2907 404 2911
rect 398 2906 404 2907
rect 518 2911 524 2912
rect 518 2907 519 2911
rect 523 2907 524 2911
rect 518 2906 524 2907
rect 782 2911 788 2912
rect 782 2907 783 2911
rect 787 2907 788 2911
rect 782 2906 788 2907
rect 798 2911 804 2912
rect 798 2907 799 2911
rect 803 2910 804 2911
rect 1096 2910 1098 2932
rect 1151 2931 1152 2932
rect 1156 2931 1157 2935
rect 1151 2930 1157 2931
rect 1279 2935 1285 2936
rect 1279 2931 1280 2935
rect 1284 2934 1285 2935
rect 1310 2935 1316 2936
rect 1310 2934 1311 2935
rect 1284 2932 1311 2934
rect 1284 2931 1285 2932
rect 1279 2930 1285 2931
rect 1310 2931 1311 2932
rect 1315 2931 1316 2935
rect 1310 2930 1316 2931
rect 1407 2935 1413 2936
rect 1407 2931 1408 2935
rect 1412 2934 1413 2935
rect 1463 2935 1469 2936
rect 1463 2934 1464 2935
rect 1412 2932 1464 2934
rect 1412 2931 1413 2932
rect 1407 2930 1413 2931
rect 1463 2931 1464 2932
rect 1468 2931 1469 2935
rect 1463 2930 1469 2931
rect 1543 2935 1549 2936
rect 1543 2931 1544 2935
rect 1548 2934 1549 2935
rect 1558 2935 1564 2936
rect 1558 2934 1559 2935
rect 1548 2932 1559 2934
rect 1548 2931 1549 2932
rect 1543 2930 1549 2931
rect 1558 2931 1559 2932
rect 1563 2931 1564 2935
rect 1558 2930 1564 2931
rect 1879 2931 1885 2932
rect 1879 2927 1880 2931
rect 1884 2930 1885 2931
rect 1894 2931 1900 2932
rect 1894 2930 1895 2931
rect 1884 2928 1895 2930
rect 1884 2927 1885 2928
rect 1879 2926 1885 2927
rect 1894 2927 1895 2928
rect 1899 2927 1900 2931
rect 1894 2926 1900 2927
rect 1902 2931 1908 2932
rect 1902 2927 1903 2931
rect 1907 2930 1908 2931
rect 2063 2931 2069 2932
rect 2063 2930 2064 2931
rect 1907 2928 2064 2930
rect 1907 2927 1908 2928
rect 1902 2926 1908 2927
rect 2063 2927 2064 2928
rect 2068 2927 2069 2931
rect 2063 2926 2069 2927
rect 2263 2931 2269 2932
rect 2263 2927 2264 2931
rect 2268 2930 2269 2931
rect 2294 2931 2300 2932
rect 2294 2930 2295 2931
rect 2268 2928 2295 2930
rect 2268 2927 2269 2928
rect 2263 2926 2269 2927
rect 2294 2927 2295 2928
rect 2299 2927 2300 2931
rect 2294 2926 2300 2927
rect 2455 2931 2461 2932
rect 2455 2927 2456 2931
rect 2460 2930 2461 2931
rect 2486 2931 2492 2932
rect 2486 2930 2487 2931
rect 2460 2928 2487 2930
rect 2460 2927 2461 2928
rect 2455 2926 2461 2927
rect 2486 2927 2487 2928
rect 2491 2927 2492 2931
rect 2486 2926 2492 2927
rect 2638 2931 2645 2932
rect 2638 2927 2639 2931
rect 2644 2927 2645 2931
rect 2638 2926 2645 2927
rect 2807 2931 2813 2932
rect 2807 2927 2808 2931
rect 2812 2930 2813 2931
rect 2894 2931 2900 2932
rect 2894 2930 2895 2931
rect 2812 2928 2895 2930
rect 2812 2927 2813 2928
rect 2807 2926 2813 2927
rect 2894 2927 2895 2928
rect 2899 2927 2900 2931
rect 2894 2926 2900 2927
rect 2959 2931 2965 2932
rect 2959 2927 2960 2931
rect 2964 2930 2965 2931
rect 2990 2931 2996 2932
rect 2990 2930 2991 2931
rect 2964 2928 2991 2930
rect 2964 2927 2965 2928
rect 2959 2926 2965 2927
rect 2990 2927 2991 2928
rect 2995 2927 2996 2931
rect 2990 2926 2996 2927
rect 3111 2931 3117 2932
rect 3111 2927 3112 2931
rect 3116 2930 3117 2931
rect 3142 2931 3148 2932
rect 3142 2930 3143 2931
rect 3116 2928 3143 2930
rect 3116 2927 3117 2928
rect 3111 2926 3117 2927
rect 3142 2927 3143 2928
rect 3147 2927 3148 2931
rect 3142 2926 3148 2927
rect 3255 2931 3261 2932
rect 3255 2927 3256 2931
rect 3260 2930 3261 2931
rect 3286 2931 3292 2932
rect 3286 2930 3287 2931
rect 3260 2928 3287 2930
rect 3260 2927 3261 2928
rect 3255 2926 3261 2927
rect 3286 2927 3287 2928
rect 3291 2927 3292 2931
rect 3286 2926 3292 2927
rect 3294 2931 3300 2932
rect 3294 2927 3295 2931
rect 3299 2930 3300 2931
rect 3407 2931 3413 2932
rect 3407 2930 3408 2931
rect 3299 2928 3408 2930
rect 3299 2927 3300 2928
rect 3294 2926 3300 2927
rect 3407 2927 3408 2928
rect 3412 2927 3413 2931
rect 3407 2926 3413 2927
rect 1766 2920 1772 2921
rect 1102 2919 1108 2920
rect 1102 2915 1103 2919
rect 1107 2915 1108 2919
rect 1230 2919 1236 2920
rect 1102 2914 1108 2915
rect 1166 2915 1172 2916
rect 1166 2911 1167 2915
rect 1171 2911 1172 2915
rect 1230 2915 1231 2919
rect 1235 2915 1236 2919
rect 1230 2914 1236 2915
rect 1358 2919 1364 2920
rect 1358 2915 1359 2919
rect 1363 2915 1364 2919
rect 1358 2914 1364 2915
rect 1494 2919 1500 2920
rect 1494 2915 1495 2919
rect 1499 2915 1500 2919
rect 1766 2916 1767 2920
rect 1771 2916 1772 2920
rect 1766 2915 1772 2916
rect 1806 2916 1812 2917
rect 3462 2916 3468 2917
rect 1494 2914 1500 2915
rect 1806 2912 1807 2916
rect 1811 2912 1812 2916
rect 1166 2910 1172 2911
rect 1182 2911 1188 2912
rect 803 2908 889 2910
rect 1049 2908 1098 2910
rect 1168 2908 1177 2910
rect 803 2907 804 2908
rect 798 2906 804 2907
rect 1182 2907 1183 2911
rect 1187 2910 1188 2911
rect 1310 2911 1316 2912
rect 1187 2908 1273 2910
rect 1187 2907 1188 2908
rect 1182 2906 1188 2907
rect 1310 2907 1311 2911
rect 1315 2910 1316 2911
rect 1463 2911 1469 2912
rect 1806 2911 1812 2912
rect 1830 2915 1836 2916
rect 1830 2911 1831 2915
rect 1835 2911 1836 2915
rect 1315 2908 1401 2910
rect 1315 2907 1316 2908
rect 1310 2906 1316 2907
rect 1463 2907 1464 2911
rect 1468 2910 1469 2911
rect 1830 2910 1836 2911
rect 2014 2915 2020 2916
rect 2014 2911 2015 2915
rect 2019 2911 2020 2915
rect 2014 2910 2020 2911
rect 2214 2915 2220 2916
rect 2214 2911 2215 2915
rect 2219 2911 2220 2915
rect 2214 2910 2220 2911
rect 2406 2915 2412 2916
rect 2406 2911 2407 2915
rect 2411 2911 2412 2915
rect 2406 2910 2412 2911
rect 2590 2915 2596 2916
rect 2590 2911 2591 2915
rect 2595 2911 2596 2915
rect 2590 2910 2596 2911
rect 2758 2915 2764 2916
rect 2758 2911 2759 2915
rect 2763 2911 2764 2915
rect 2758 2910 2764 2911
rect 2910 2915 2916 2916
rect 2910 2911 2911 2915
rect 2915 2911 2916 2915
rect 2910 2910 2916 2911
rect 3062 2915 3068 2916
rect 3062 2911 3063 2915
rect 3067 2911 3068 2915
rect 3062 2910 3068 2911
rect 3206 2915 3212 2916
rect 3206 2911 3207 2915
rect 3211 2911 3212 2915
rect 3206 2910 3212 2911
rect 3358 2915 3364 2916
rect 3358 2911 3359 2915
rect 3363 2911 3364 2915
rect 3462 2912 3463 2916
rect 3467 2912 3468 2916
rect 3462 2911 3468 2912
rect 3358 2910 3364 2911
rect 1468 2908 1537 2910
rect 1468 2907 1469 2908
rect 1463 2906 1469 2907
rect 1902 2907 1908 2908
rect 640 2904 649 2906
rect 110 2903 116 2904
rect 110 2899 111 2903
rect 115 2899 116 2903
rect 638 2903 644 2904
rect 110 2898 116 2899
rect 326 2900 332 2901
rect 326 2896 327 2900
rect 331 2896 332 2900
rect 326 2895 332 2896
rect 446 2900 452 2901
rect 446 2896 447 2900
rect 451 2896 452 2900
rect 446 2895 452 2896
rect 574 2900 580 2901
rect 574 2896 575 2900
rect 579 2896 580 2900
rect 638 2899 639 2903
rect 643 2899 644 2903
rect 1766 2903 1772 2904
rect 638 2898 644 2899
rect 710 2900 716 2901
rect 574 2895 580 2896
rect 710 2896 711 2900
rect 715 2896 716 2900
rect 710 2895 716 2896
rect 846 2900 852 2901
rect 846 2896 847 2900
rect 851 2896 852 2900
rect 846 2895 852 2896
rect 974 2900 980 2901
rect 974 2896 975 2900
rect 979 2896 980 2900
rect 974 2895 980 2896
rect 1102 2900 1108 2901
rect 1102 2896 1103 2900
rect 1107 2896 1108 2900
rect 1102 2895 1108 2896
rect 1230 2900 1236 2901
rect 1230 2896 1231 2900
rect 1235 2896 1236 2900
rect 1230 2895 1236 2896
rect 1358 2900 1364 2901
rect 1358 2896 1359 2900
rect 1363 2896 1364 2900
rect 1358 2895 1364 2896
rect 1494 2900 1500 2901
rect 1494 2896 1495 2900
rect 1499 2896 1500 2900
rect 1766 2899 1767 2903
rect 1771 2899 1772 2903
rect 1902 2903 1903 2907
rect 1907 2903 1908 2907
rect 2194 2907 2200 2908
rect 1902 2902 1908 2903
rect 2086 2903 2092 2904
rect 1766 2898 1772 2899
rect 1806 2899 1812 2900
rect 1494 2895 1500 2896
rect 1806 2895 1807 2899
rect 1811 2895 1812 2899
rect 2086 2899 2087 2903
rect 2091 2899 2092 2903
rect 2194 2903 2195 2907
rect 2199 2906 2200 2907
rect 2294 2907 2300 2908
rect 2199 2904 2257 2906
rect 2199 2903 2200 2904
rect 2194 2902 2200 2903
rect 2294 2903 2295 2907
rect 2299 2906 2300 2907
rect 2486 2907 2492 2908
rect 2299 2904 2449 2906
rect 2299 2903 2300 2904
rect 2294 2902 2300 2903
rect 2486 2903 2487 2907
rect 2491 2906 2492 2907
rect 2894 2907 2900 2908
rect 2491 2904 2633 2906
rect 2491 2903 2492 2904
rect 2486 2902 2492 2903
rect 2830 2903 2836 2904
rect 2086 2898 2092 2899
rect 2830 2899 2831 2903
rect 2835 2899 2836 2903
rect 2894 2903 2895 2907
rect 2899 2906 2900 2907
rect 2990 2907 2996 2908
rect 2899 2904 2953 2906
rect 2899 2903 2900 2904
rect 2894 2902 2900 2903
rect 2990 2903 2991 2907
rect 2995 2906 2996 2907
rect 3142 2907 3148 2908
rect 2995 2904 3105 2906
rect 2995 2903 2996 2904
rect 2990 2902 2996 2903
rect 3142 2903 3143 2907
rect 3147 2906 3148 2907
rect 3286 2907 3292 2908
rect 3147 2904 3249 2906
rect 3147 2903 3148 2904
rect 3142 2902 3148 2903
rect 3286 2903 3287 2907
rect 3291 2906 3292 2907
rect 3291 2904 3401 2906
rect 3291 2903 3292 2904
rect 3286 2902 3292 2903
rect 2830 2898 2836 2899
rect 3462 2899 3468 2900
rect 1806 2894 1812 2895
rect 1830 2896 1836 2897
rect 1830 2892 1831 2896
rect 1835 2892 1836 2896
rect 1830 2891 1836 2892
rect 2014 2896 2020 2897
rect 2014 2892 2015 2896
rect 2019 2892 2020 2896
rect 2014 2891 2020 2892
rect 2214 2896 2220 2897
rect 2214 2892 2215 2896
rect 2219 2892 2220 2896
rect 2214 2891 2220 2892
rect 2406 2896 2412 2897
rect 2406 2892 2407 2896
rect 2411 2892 2412 2896
rect 2406 2891 2412 2892
rect 2590 2896 2596 2897
rect 2590 2892 2591 2896
rect 2595 2892 2596 2896
rect 2590 2891 2596 2892
rect 2758 2896 2764 2897
rect 2758 2892 2759 2896
rect 2763 2892 2764 2896
rect 2758 2891 2764 2892
rect 2910 2896 2916 2897
rect 2910 2892 2911 2896
rect 2915 2892 2916 2896
rect 2910 2891 2916 2892
rect 3062 2896 3068 2897
rect 3062 2892 3063 2896
rect 3067 2892 3068 2896
rect 3062 2891 3068 2892
rect 3206 2896 3212 2897
rect 3206 2892 3207 2896
rect 3211 2892 3212 2896
rect 3206 2891 3212 2892
rect 3358 2896 3364 2897
rect 3358 2892 3359 2896
rect 3363 2892 3364 2896
rect 3462 2895 3463 2899
rect 3467 2895 3468 2899
rect 3462 2894 3468 2895
rect 3358 2891 3364 2892
rect 1830 2852 1836 2853
rect 1806 2849 1812 2850
rect 134 2848 140 2849
rect 110 2845 116 2846
rect 110 2841 111 2845
rect 115 2841 116 2845
rect 134 2844 135 2848
rect 139 2844 140 2848
rect 134 2843 140 2844
rect 254 2848 260 2849
rect 254 2844 255 2848
rect 259 2844 260 2848
rect 254 2843 260 2844
rect 414 2848 420 2849
rect 414 2844 415 2848
rect 419 2844 420 2848
rect 414 2843 420 2844
rect 574 2848 580 2849
rect 574 2844 575 2848
rect 579 2844 580 2848
rect 574 2843 580 2844
rect 734 2848 740 2849
rect 734 2844 735 2848
rect 739 2844 740 2848
rect 734 2843 740 2844
rect 894 2848 900 2849
rect 894 2844 895 2848
rect 899 2844 900 2848
rect 894 2843 900 2844
rect 1046 2848 1052 2849
rect 1046 2844 1047 2848
rect 1051 2844 1052 2848
rect 1046 2843 1052 2844
rect 1190 2848 1196 2849
rect 1190 2844 1191 2848
rect 1195 2844 1196 2848
rect 1190 2843 1196 2844
rect 1342 2848 1348 2849
rect 1342 2844 1343 2848
rect 1347 2844 1348 2848
rect 1342 2843 1348 2844
rect 1494 2848 1500 2849
rect 1494 2844 1495 2848
rect 1499 2844 1500 2848
rect 1494 2843 1500 2844
rect 1766 2845 1772 2846
rect 110 2840 116 2841
rect 1766 2841 1767 2845
rect 1771 2841 1772 2845
rect 1806 2845 1807 2849
rect 1811 2845 1812 2849
rect 1830 2848 1831 2852
rect 1835 2848 1836 2852
rect 1830 2847 1836 2848
rect 1998 2852 2004 2853
rect 1998 2848 1999 2852
rect 2003 2848 2004 2852
rect 1998 2847 2004 2848
rect 2190 2852 2196 2853
rect 2190 2848 2191 2852
rect 2195 2848 2196 2852
rect 2190 2847 2196 2848
rect 2382 2852 2388 2853
rect 2382 2848 2383 2852
rect 2387 2848 2388 2852
rect 2382 2847 2388 2848
rect 2566 2852 2572 2853
rect 2566 2848 2567 2852
rect 2571 2848 2572 2852
rect 2566 2847 2572 2848
rect 2734 2852 2740 2853
rect 2734 2848 2735 2852
rect 2739 2848 2740 2852
rect 2734 2847 2740 2848
rect 2902 2852 2908 2853
rect 2902 2848 2903 2852
rect 2907 2848 2908 2852
rect 2902 2847 2908 2848
rect 3062 2852 3068 2853
rect 3062 2848 3063 2852
rect 3067 2848 3068 2852
rect 3062 2847 3068 2848
rect 3222 2852 3228 2853
rect 3222 2848 3223 2852
rect 3227 2848 3228 2852
rect 3222 2847 3228 2848
rect 3366 2852 3372 2853
rect 3366 2848 3367 2852
rect 3371 2848 3372 2852
rect 3366 2847 3372 2848
rect 3462 2849 3468 2850
rect 1806 2844 1812 2845
rect 3462 2845 3463 2849
rect 3467 2845 3468 2849
rect 3462 2844 3468 2845
rect 1766 2840 1772 2841
rect 1894 2843 1900 2844
rect 198 2839 204 2840
rect 198 2835 199 2839
rect 203 2835 204 2839
rect 198 2834 204 2835
rect 214 2839 220 2840
rect 214 2835 215 2839
rect 219 2838 220 2839
rect 334 2839 340 2840
rect 219 2836 297 2838
rect 219 2835 220 2836
rect 214 2834 220 2835
rect 334 2835 335 2839
rect 339 2838 340 2839
rect 646 2839 652 2840
rect 339 2836 457 2838
rect 339 2835 340 2836
rect 334 2834 340 2835
rect 646 2835 647 2839
rect 651 2835 652 2839
rect 646 2834 652 2835
rect 726 2839 732 2840
rect 726 2835 727 2839
rect 731 2838 732 2839
rect 966 2839 972 2840
rect 731 2836 777 2838
rect 731 2835 732 2836
rect 726 2834 732 2835
rect 966 2835 967 2839
rect 971 2835 972 2839
rect 966 2834 972 2835
rect 1118 2839 1124 2840
rect 1118 2835 1119 2839
rect 1123 2835 1124 2839
rect 1118 2834 1124 2835
rect 1262 2839 1268 2840
rect 1262 2835 1263 2839
rect 1267 2835 1268 2839
rect 1262 2834 1268 2835
rect 1414 2839 1420 2840
rect 1414 2835 1415 2839
rect 1419 2835 1420 2839
rect 1414 2834 1420 2835
rect 1558 2839 1564 2840
rect 1558 2835 1559 2839
rect 1563 2835 1564 2839
rect 1894 2839 1895 2843
rect 1899 2839 1900 2843
rect 1894 2838 1900 2839
rect 1910 2843 1916 2844
rect 1910 2839 1911 2843
rect 1915 2842 1916 2843
rect 2262 2843 2268 2844
rect 1915 2840 2041 2842
rect 1915 2839 1916 2840
rect 1910 2838 1916 2839
rect 2262 2839 2263 2843
rect 2267 2839 2268 2843
rect 2262 2838 2268 2839
rect 2454 2843 2460 2844
rect 2454 2839 2455 2843
rect 2459 2839 2460 2843
rect 2454 2838 2460 2839
rect 2638 2843 2644 2844
rect 2638 2839 2639 2843
rect 2643 2839 2644 2843
rect 2862 2843 2868 2844
rect 2862 2842 2863 2843
rect 2809 2840 2863 2842
rect 2638 2838 2644 2839
rect 2862 2839 2863 2840
rect 2867 2839 2868 2843
rect 2862 2838 2868 2839
rect 2974 2843 2980 2844
rect 2974 2839 2975 2843
rect 2979 2839 2980 2843
rect 2974 2838 2980 2839
rect 3126 2843 3132 2844
rect 3126 2839 3127 2843
rect 3131 2839 3132 2843
rect 3126 2838 3132 2839
rect 3294 2843 3300 2844
rect 3294 2839 3295 2843
rect 3299 2839 3300 2843
rect 3294 2838 3300 2839
rect 3430 2843 3436 2844
rect 3430 2839 3431 2843
rect 3435 2839 3436 2843
rect 3430 2838 3436 2839
rect 1558 2834 1564 2835
rect 1830 2833 1836 2834
rect 1806 2832 1812 2833
rect 134 2829 140 2830
rect 110 2828 116 2829
rect 110 2824 111 2828
rect 115 2824 116 2828
rect 134 2825 135 2829
rect 139 2825 140 2829
rect 134 2824 140 2825
rect 254 2829 260 2830
rect 254 2825 255 2829
rect 259 2825 260 2829
rect 254 2824 260 2825
rect 414 2829 420 2830
rect 414 2825 415 2829
rect 419 2825 420 2829
rect 414 2824 420 2825
rect 574 2829 580 2830
rect 574 2825 575 2829
rect 579 2825 580 2829
rect 574 2824 580 2825
rect 734 2829 740 2830
rect 734 2825 735 2829
rect 739 2825 740 2829
rect 734 2824 740 2825
rect 894 2829 900 2830
rect 894 2825 895 2829
rect 899 2825 900 2829
rect 894 2824 900 2825
rect 1046 2829 1052 2830
rect 1046 2825 1047 2829
rect 1051 2825 1052 2829
rect 1046 2824 1052 2825
rect 1190 2829 1196 2830
rect 1190 2825 1191 2829
rect 1195 2825 1196 2829
rect 1190 2824 1196 2825
rect 1342 2829 1348 2830
rect 1342 2825 1343 2829
rect 1347 2825 1348 2829
rect 1342 2824 1348 2825
rect 1494 2829 1500 2830
rect 1494 2825 1495 2829
rect 1499 2825 1500 2829
rect 1494 2824 1500 2825
rect 1766 2828 1772 2829
rect 1766 2824 1767 2828
rect 1771 2824 1772 2828
rect 1806 2828 1807 2832
rect 1811 2828 1812 2832
rect 1830 2829 1831 2833
rect 1835 2829 1836 2833
rect 1830 2828 1836 2829
rect 1998 2833 2004 2834
rect 1998 2829 1999 2833
rect 2003 2829 2004 2833
rect 1998 2828 2004 2829
rect 2190 2833 2196 2834
rect 2190 2829 2191 2833
rect 2195 2829 2196 2833
rect 2190 2828 2196 2829
rect 2382 2833 2388 2834
rect 2382 2829 2383 2833
rect 2387 2829 2388 2833
rect 2382 2828 2388 2829
rect 2566 2833 2572 2834
rect 2566 2829 2567 2833
rect 2571 2829 2572 2833
rect 2566 2828 2572 2829
rect 2734 2833 2740 2834
rect 2734 2829 2735 2833
rect 2739 2829 2740 2833
rect 2734 2828 2740 2829
rect 2902 2833 2908 2834
rect 2902 2829 2903 2833
rect 2907 2829 2908 2833
rect 2902 2828 2908 2829
rect 3062 2833 3068 2834
rect 3062 2829 3063 2833
rect 3067 2829 3068 2833
rect 3062 2828 3068 2829
rect 3222 2833 3228 2834
rect 3222 2829 3223 2833
rect 3227 2829 3228 2833
rect 3222 2828 3228 2829
rect 3366 2833 3372 2834
rect 3366 2829 3367 2833
rect 3371 2829 3372 2833
rect 3366 2828 3372 2829
rect 3462 2832 3468 2833
rect 3462 2828 3463 2832
rect 3467 2828 3468 2832
rect 1806 2827 1812 2828
rect 3462 2827 3468 2828
rect 110 2823 116 2824
rect 1766 2823 1772 2824
rect 1879 2815 1885 2816
rect 183 2811 189 2812
rect 183 2807 184 2811
rect 188 2810 189 2811
rect 214 2811 220 2812
rect 214 2810 215 2811
rect 188 2808 215 2810
rect 188 2807 189 2808
rect 183 2806 189 2807
rect 214 2807 215 2808
rect 219 2807 220 2811
rect 214 2806 220 2807
rect 303 2811 309 2812
rect 303 2807 304 2811
rect 308 2810 309 2811
rect 334 2811 340 2812
rect 334 2810 335 2811
rect 308 2808 335 2810
rect 308 2807 309 2808
rect 303 2806 309 2807
rect 334 2807 335 2808
rect 339 2807 340 2811
rect 334 2806 340 2807
rect 463 2811 469 2812
rect 463 2807 464 2811
rect 468 2810 469 2811
rect 623 2811 629 2812
rect 468 2808 598 2810
rect 468 2807 469 2808
rect 463 2806 469 2807
rect 596 2802 598 2808
rect 623 2807 624 2811
rect 628 2810 629 2811
rect 638 2811 644 2812
rect 638 2810 639 2811
rect 628 2808 639 2810
rect 628 2807 629 2808
rect 623 2806 629 2807
rect 638 2807 639 2808
rect 643 2807 644 2811
rect 638 2806 644 2807
rect 646 2811 652 2812
rect 646 2807 647 2811
rect 651 2810 652 2811
rect 783 2811 789 2812
rect 783 2810 784 2811
rect 651 2808 784 2810
rect 651 2807 652 2808
rect 646 2806 652 2807
rect 783 2807 784 2808
rect 788 2807 789 2811
rect 783 2806 789 2807
rect 943 2811 949 2812
rect 943 2807 944 2811
rect 948 2810 949 2811
rect 966 2811 972 2812
rect 948 2808 962 2810
rect 948 2807 949 2808
rect 943 2806 949 2807
rect 726 2803 732 2804
rect 726 2802 727 2803
rect 596 2800 727 2802
rect 726 2799 727 2800
rect 731 2799 732 2803
rect 960 2802 962 2808
rect 966 2807 967 2811
rect 971 2810 972 2811
rect 1095 2811 1101 2812
rect 1095 2810 1096 2811
rect 971 2808 1096 2810
rect 971 2807 972 2808
rect 966 2806 972 2807
rect 1095 2807 1096 2808
rect 1100 2807 1101 2811
rect 1095 2806 1101 2807
rect 1118 2811 1124 2812
rect 1118 2807 1119 2811
rect 1123 2810 1124 2811
rect 1239 2811 1245 2812
rect 1239 2810 1240 2811
rect 1123 2808 1240 2810
rect 1123 2807 1124 2808
rect 1118 2806 1124 2807
rect 1239 2807 1240 2808
rect 1244 2807 1245 2811
rect 1239 2806 1245 2807
rect 1262 2811 1268 2812
rect 1262 2807 1263 2811
rect 1267 2810 1268 2811
rect 1391 2811 1397 2812
rect 1391 2810 1392 2811
rect 1267 2808 1392 2810
rect 1267 2807 1268 2808
rect 1262 2806 1268 2807
rect 1391 2807 1392 2808
rect 1396 2807 1397 2811
rect 1391 2806 1397 2807
rect 1414 2811 1420 2812
rect 1414 2807 1415 2811
rect 1419 2810 1420 2811
rect 1543 2811 1549 2812
rect 1543 2810 1544 2811
rect 1419 2808 1544 2810
rect 1419 2807 1420 2808
rect 1414 2806 1420 2807
rect 1543 2807 1544 2808
rect 1548 2807 1549 2811
rect 1879 2811 1880 2815
rect 1884 2814 1885 2815
rect 1910 2815 1916 2816
rect 1910 2814 1911 2815
rect 1884 2812 1911 2814
rect 1884 2811 1885 2812
rect 1879 2810 1885 2811
rect 1910 2811 1911 2812
rect 1915 2811 1916 2815
rect 1910 2810 1916 2811
rect 2047 2815 2053 2816
rect 2047 2811 2048 2815
rect 2052 2814 2053 2815
rect 2086 2815 2092 2816
rect 2086 2814 2087 2815
rect 2052 2812 2087 2814
rect 2052 2811 2053 2812
rect 2047 2810 2053 2811
rect 2086 2811 2087 2812
rect 2091 2811 2092 2815
rect 2086 2810 2092 2811
rect 2146 2815 2152 2816
rect 2146 2811 2147 2815
rect 2151 2814 2152 2815
rect 2239 2815 2245 2816
rect 2239 2814 2240 2815
rect 2151 2812 2240 2814
rect 2151 2811 2152 2812
rect 2146 2810 2152 2811
rect 2239 2811 2240 2812
rect 2244 2811 2245 2815
rect 2239 2810 2245 2811
rect 2262 2815 2268 2816
rect 2262 2811 2263 2815
rect 2267 2814 2268 2815
rect 2431 2815 2437 2816
rect 2431 2814 2432 2815
rect 2267 2812 2432 2814
rect 2267 2811 2268 2812
rect 2262 2810 2268 2811
rect 2431 2811 2432 2812
rect 2436 2811 2437 2815
rect 2431 2810 2437 2811
rect 2454 2815 2460 2816
rect 2454 2811 2455 2815
rect 2459 2814 2460 2815
rect 2615 2815 2621 2816
rect 2615 2814 2616 2815
rect 2459 2812 2616 2814
rect 2459 2811 2460 2812
rect 2454 2810 2460 2811
rect 2615 2811 2616 2812
rect 2620 2811 2621 2815
rect 2615 2810 2621 2811
rect 2783 2815 2789 2816
rect 2783 2811 2784 2815
rect 2788 2814 2789 2815
rect 2830 2815 2836 2816
rect 2830 2814 2831 2815
rect 2788 2812 2831 2814
rect 2788 2811 2789 2812
rect 2783 2810 2789 2811
rect 2830 2811 2831 2812
rect 2835 2811 2836 2815
rect 2830 2810 2836 2811
rect 2862 2815 2868 2816
rect 2862 2811 2863 2815
rect 2867 2814 2868 2815
rect 2951 2815 2957 2816
rect 2951 2814 2952 2815
rect 2867 2812 2952 2814
rect 2867 2811 2868 2812
rect 2862 2810 2868 2811
rect 2951 2811 2952 2812
rect 2956 2811 2957 2815
rect 2951 2810 2957 2811
rect 2974 2815 2980 2816
rect 2974 2811 2975 2815
rect 2979 2814 2980 2815
rect 3111 2815 3117 2816
rect 3111 2814 3112 2815
rect 2979 2812 3112 2814
rect 2979 2811 2980 2812
rect 2974 2810 2980 2811
rect 3111 2811 3112 2812
rect 3116 2811 3117 2815
rect 3111 2810 3117 2811
rect 3271 2815 3277 2816
rect 3271 2811 3272 2815
rect 3276 2814 3277 2815
rect 3302 2815 3308 2816
rect 3302 2814 3303 2815
rect 3276 2812 3303 2814
rect 3276 2811 3277 2812
rect 3271 2810 3277 2811
rect 3302 2811 3303 2812
rect 3307 2811 3308 2815
rect 3302 2810 3308 2811
rect 3415 2815 3421 2816
rect 3415 2811 3416 2815
rect 3420 2814 3421 2815
rect 3438 2815 3444 2816
rect 3438 2814 3439 2815
rect 3420 2812 3439 2814
rect 3420 2811 3421 2812
rect 3415 2810 3421 2811
rect 3438 2811 3439 2812
rect 3443 2811 3444 2815
rect 3438 2810 3444 2811
rect 1543 2806 1549 2807
rect 2990 2807 2996 2808
rect 2990 2806 2991 2807
rect 2736 2804 2991 2806
rect 1278 2803 1284 2804
rect 1278 2802 1279 2803
rect 960 2800 1279 2802
rect 726 2798 732 2799
rect 1278 2799 1279 2800
rect 1283 2799 1284 2803
rect 1278 2798 1284 2799
rect 1879 2799 1885 2800
rect 1879 2795 1880 2799
rect 1884 2798 1885 2799
rect 1894 2799 1900 2800
rect 1894 2798 1895 2799
rect 1884 2796 1895 2798
rect 1884 2795 1885 2796
rect 1879 2794 1885 2795
rect 1894 2795 1895 2796
rect 1899 2795 1900 2799
rect 1894 2794 1900 2795
rect 2063 2799 2069 2800
rect 2063 2795 2064 2799
rect 2068 2798 2069 2799
rect 2094 2799 2100 2800
rect 2094 2798 2095 2799
rect 2068 2796 2095 2798
rect 2068 2795 2069 2796
rect 2063 2794 2069 2795
rect 2094 2795 2095 2796
rect 2099 2795 2100 2799
rect 2094 2794 2100 2795
rect 2263 2799 2269 2800
rect 2263 2795 2264 2799
rect 2268 2798 2269 2799
rect 2294 2799 2300 2800
rect 2294 2798 2295 2799
rect 2268 2796 2295 2798
rect 2268 2795 2269 2796
rect 2263 2794 2269 2795
rect 2294 2795 2295 2796
rect 2299 2795 2300 2799
rect 2294 2794 2300 2795
rect 2455 2799 2461 2800
rect 2455 2795 2456 2799
rect 2460 2798 2461 2799
rect 2470 2799 2476 2800
rect 2470 2798 2471 2799
rect 2460 2796 2471 2798
rect 2460 2795 2461 2796
rect 2455 2794 2461 2795
rect 2470 2795 2471 2796
rect 2475 2795 2476 2799
rect 2470 2794 2476 2795
rect 2631 2799 2637 2800
rect 2631 2795 2632 2799
rect 2636 2798 2637 2799
rect 2736 2798 2738 2804
rect 2990 2803 2991 2804
rect 2995 2803 2996 2807
rect 2990 2802 2996 2803
rect 2636 2796 2738 2798
rect 2742 2799 2748 2800
rect 2636 2795 2637 2796
rect 2631 2794 2637 2795
rect 2742 2795 2743 2799
rect 2747 2798 2748 2799
rect 2799 2799 2805 2800
rect 2799 2798 2800 2799
rect 2747 2796 2800 2798
rect 2747 2795 2748 2796
rect 2742 2794 2748 2795
rect 2799 2795 2800 2796
rect 2804 2795 2805 2799
rect 2799 2794 2805 2795
rect 2822 2799 2828 2800
rect 2822 2795 2823 2799
rect 2827 2798 2828 2799
rect 2959 2799 2965 2800
rect 2959 2798 2960 2799
rect 2827 2796 2960 2798
rect 2827 2795 2828 2796
rect 2822 2794 2828 2795
rect 2959 2795 2960 2796
rect 2964 2795 2965 2799
rect 2959 2794 2965 2795
rect 3119 2799 3125 2800
rect 3119 2795 3120 2799
rect 3124 2795 3125 2799
rect 3119 2794 3125 2795
rect 3262 2799 3268 2800
rect 3262 2795 3263 2799
rect 3267 2798 3268 2799
rect 3279 2799 3285 2800
rect 3279 2798 3280 2799
rect 3267 2796 3280 2798
rect 3267 2795 3268 2796
rect 3262 2794 3268 2795
rect 3279 2795 3280 2796
rect 3284 2795 3285 2799
rect 3279 2794 3285 2795
rect 3415 2799 3421 2800
rect 3415 2795 3416 2799
rect 3420 2798 3421 2799
rect 3430 2799 3436 2800
rect 3430 2798 3431 2799
rect 3420 2796 3431 2798
rect 3420 2795 3421 2796
rect 3415 2794 3421 2795
rect 3430 2795 3431 2796
rect 3435 2795 3436 2799
rect 3430 2794 3436 2795
rect 183 2787 189 2788
rect 183 2783 184 2787
rect 188 2786 189 2787
rect 198 2787 204 2788
rect 198 2786 199 2787
rect 188 2784 199 2786
rect 188 2783 189 2784
rect 183 2782 189 2783
rect 198 2783 199 2784
rect 203 2783 204 2787
rect 198 2782 204 2783
rect 206 2787 212 2788
rect 206 2783 207 2787
rect 211 2786 212 2787
rect 295 2787 301 2788
rect 295 2786 296 2787
rect 211 2784 296 2786
rect 211 2783 212 2784
rect 206 2782 212 2783
rect 295 2783 296 2784
rect 300 2783 301 2787
rect 295 2782 301 2783
rect 318 2787 324 2788
rect 318 2783 319 2787
rect 323 2786 324 2787
rect 439 2787 445 2788
rect 439 2786 440 2787
rect 323 2784 440 2786
rect 323 2783 324 2784
rect 318 2782 324 2783
rect 439 2783 440 2784
rect 444 2783 445 2787
rect 439 2782 445 2783
rect 462 2787 468 2788
rect 462 2783 463 2787
rect 467 2786 468 2787
rect 591 2787 597 2788
rect 591 2786 592 2787
rect 467 2784 592 2786
rect 467 2783 468 2784
rect 462 2782 468 2783
rect 591 2783 592 2784
rect 596 2783 597 2787
rect 591 2782 597 2783
rect 614 2787 620 2788
rect 614 2783 615 2787
rect 619 2786 620 2787
rect 743 2787 749 2788
rect 743 2786 744 2787
rect 619 2784 744 2786
rect 619 2783 620 2784
rect 614 2782 620 2783
rect 743 2783 744 2784
rect 748 2783 749 2787
rect 743 2782 749 2783
rect 902 2787 909 2788
rect 902 2783 903 2787
rect 908 2783 909 2787
rect 902 2782 909 2783
rect 926 2787 932 2788
rect 926 2783 927 2787
rect 931 2786 932 2787
rect 1071 2787 1077 2788
rect 1071 2786 1072 2787
rect 931 2784 1072 2786
rect 931 2783 932 2784
rect 926 2782 932 2783
rect 1071 2783 1072 2784
rect 1076 2783 1077 2787
rect 1071 2782 1077 2783
rect 1094 2787 1100 2788
rect 1094 2783 1095 2787
rect 1099 2786 1100 2787
rect 1239 2787 1245 2788
rect 1239 2786 1240 2787
rect 1099 2784 1240 2786
rect 1099 2783 1100 2784
rect 1094 2782 1100 2783
rect 1239 2783 1240 2784
rect 1244 2783 1245 2787
rect 1239 2782 1245 2783
rect 1262 2787 1268 2788
rect 1262 2783 1263 2787
rect 1267 2786 1268 2787
rect 1407 2787 1413 2788
rect 1407 2786 1408 2787
rect 1267 2784 1408 2786
rect 1267 2783 1268 2784
rect 1262 2782 1268 2783
rect 1407 2783 1408 2784
rect 1412 2783 1413 2787
rect 1407 2782 1413 2783
rect 1575 2787 1581 2788
rect 1575 2783 1576 2787
rect 1580 2786 1581 2787
rect 1606 2787 1612 2788
rect 1606 2786 1607 2787
rect 1580 2784 1607 2786
rect 1580 2783 1581 2784
rect 1575 2782 1581 2783
rect 1606 2783 1607 2784
rect 1611 2783 1612 2787
rect 1606 2782 1612 2783
rect 1719 2787 1725 2788
rect 1719 2783 1720 2787
rect 1724 2786 1725 2787
rect 1724 2784 1798 2786
rect 1724 2783 1725 2784
rect 1719 2782 1725 2783
rect 1796 2774 1798 2784
rect 1806 2784 1812 2785
rect 3462 2784 3468 2785
rect 1806 2780 1807 2784
rect 1811 2780 1812 2784
rect 1806 2779 1812 2780
rect 1830 2783 1836 2784
rect 1830 2779 1831 2783
rect 1835 2779 1836 2783
rect 1830 2778 1836 2779
rect 2014 2783 2020 2784
rect 2014 2779 2015 2783
rect 2019 2779 2020 2783
rect 2146 2783 2152 2784
rect 2146 2782 2147 2783
rect 2014 2778 2020 2779
rect 2088 2780 2147 2782
rect 110 2772 116 2773
rect 1766 2772 1772 2773
rect 1796 2772 1873 2774
rect 2088 2773 2090 2780
rect 2146 2779 2147 2780
rect 2151 2779 2152 2783
rect 2146 2778 2152 2779
rect 2214 2783 2220 2784
rect 2214 2779 2215 2783
rect 2219 2779 2220 2783
rect 2214 2778 2220 2779
rect 2406 2783 2412 2784
rect 2406 2779 2407 2783
rect 2411 2779 2412 2783
rect 2406 2778 2412 2779
rect 2582 2783 2588 2784
rect 2582 2779 2583 2783
rect 2587 2779 2588 2783
rect 2582 2778 2588 2779
rect 2750 2783 2756 2784
rect 2750 2779 2751 2783
rect 2755 2779 2756 2783
rect 2750 2778 2756 2779
rect 2910 2783 2916 2784
rect 2910 2779 2911 2783
rect 2915 2779 2916 2783
rect 2910 2778 2916 2779
rect 3070 2783 3076 2784
rect 3070 2779 3071 2783
rect 3075 2779 3076 2783
rect 3070 2778 3076 2779
rect 3230 2783 3236 2784
rect 3230 2779 3231 2783
rect 3235 2779 3236 2783
rect 3230 2778 3236 2779
rect 3366 2783 3372 2784
rect 3366 2779 3367 2783
rect 3371 2779 3372 2783
rect 3462 2780 3463 2784
rect 3467 2780 3468 2784
rect 3462 2779 3468 2780
rect 3366 2778 3372 2779
rect 2094 2775 2100 2776
rect 110 2768 111 2772
rect 115 2768 116 2772
rect 110 2767 116 2768
rect 134 2771 140 2772
rect 134 2767 135 2771
rect 139 2767 140 2771
rect 134 2766 140 2767
rect 246 2771 252 2772
rect 246 2767 247 2771
rect 251 2767 252 2771
rect 246 2766 252 2767
rect 390 2771 396 2772
rect 390 2767 391 2771
rect 395 2767 396 2771
rect 390 2766 396 2767
rect 542 2771 548 2772
rect 542 2767 543 2771
rect 547 2767 548 2771
rect 542 2766 548 2767
rect 694 2771 700 2772
rect 694 2767 695 2771
rect 699 2767 700 2771
rect 694 2766 700 2767
rect 854 2771 860 2772
rect 854 2767 855 2771
rect 859 2767 860 2771
rect 854 2766 860 2767
rect 1022 2771 1028 2772
rect 1022 2767 1023 2771
rect 1027 2767 1028 2771
rect 1022 2766 1028 2767
rect 1190 2771 1196 2772
rect 1190 2767 1191 2771
rect 1195 2767 1196 2771
rect 1190 2766 1196 2767
rect 1358 2771 1364 2772
rect 1358 2767 1359 2771
rect 1363 2767 1364 2771
rect 1358 2766 1364 2767
rect 1526 2771 1532 2772
rect 1526 2767 1527 2771
rect 1531 2767 1532 2771
rect 1526 2766 1532 2767
rect 1670 2771 1676 2772
rect 1670 2767 1671 2771
rect 1675 2767 1676 2771
rect 1766 2768 1767 2772
rect 1771 2768 1772 2772
rect 2094 2771 2095 2775
rect 2099 2774 2100 2775
rect 2294 2775 2300 2776
rect 2099 2772 2257 2774
rect 2099 2771 2100 2772
rect 2094 2770 2100 2771
rect 2294 2771 2295 2775
rect 2299 2774 2300 2775
rect 2742 2775 2748 2776
rect 2742 2774 2743 2775
rect 2299 2772 2449 2774
rect 2657 2772 2743 2774
rect 2299 2771 2300 2772
rect 2294 2770 2300 2771
rect 2742 2771 2743 2772
rect 2747 2771 2748 2775
rect 2742 2770 2748 2771
rect 2822 2775 2828 2776
rect 2822 2771 2823 2775
rect 2827 2771 2828 2775
rect 2990 2775 2996 2776
rect 2822 2770 2828 2771
rect 2982 2771 2988 2772
rect 1766 2767 1772 2768
rect 1806 2767 1812 2768
rect 1670 2766 1676 2767
rect 206 2763 212 2764
rect 206 2759 207 2763
rect 211 2759 212 2763
rect 206 2758 212 2759
rect 318 2763 324 2764
rect 318 2759 319 2763
rect 323 2759 324 2763
rect 318 2758 324 2759
rect 462 2763 468 2764
rect 462 2759 463 2763
rect 467 2759 468 2763
rect 462 2758 468 2759
rect 614 2763 620 2764
rect 614 2759 615 2763
rect 619 2759 620 2763
rect 614 2758 620 2759
rect 622 2763 628 2764
rect 622 2759 623 2763
rect 627 2762 628 2763
rect 926 2763 932 2764
rect 627 2760 737 2762
rect 627 2759 628 2760
rect 622 2758 628 2759
rect 926 2759 927 2763
rect 931 2759 932 2763
rect 926 2758 932 2759
rect 1094 2763 1100 2764
rect 1094 2759 1095 2763
rect 1099 2759 1100 2763
rect 1094 2758 1100 2759
rect 1262 2763 1268 2764
rect 1262 2759 1263 2763
rect 1267 2759 1268 2763
rect 1262 2758 1268 2759
rect 1278 2763 1284 2764
rect 1278 2759 1279 2763
rect 1283 2762 1284 2763
rect 1606 2763 1612 2764
rect 1283 2760 1401 2762
rect 1283 2759 1284 2760
rect 1278 2758 1284 2759
rect 1598 2759 1604 2760
rect 110 2755 116 2756
rect 110 2751 111 2755
rect 115 2751 116 2755
rect 1598 2755 1599 2759
rect 1603 2755 1604 2759
rect 1606 2759 1607 2763
rect 1611 2762 1612 2763
rect 1806 2763 1807 2767
rect 1811 2763 1812 2767
rect 2982 2767 2983 2771
rect 2987 2767 2988 2771
rect 2990 2771 2991 2775
rect 2995 2774 2996 2775
rect 3302 2775 3308 2776
rect 2995 2772 3113 2774
rect 2995 2771 2996 2772
rect 2990 2770 2996 2771
rect 3302 2771 3303 2775
rect 3307 2771 3308 2775
rect 3302 2770 3308 2771
rect 3438 2771 3444 2772
rect 2982 2766 2988 2767
rect 3438 2767 3439 2771
rect 3443 2767 3444 2771
rect 3438 2766 3444 2767
rect 3462 2767 3468 2768
rect 1806 2762 1812 2763
rect 1830 2764 1836 2765
rect 1611 2760 1713 2762
rect 1830 2760 1831 2764
rect 1835 2760 1836 2764
rect 1611 2759 1612 2760
rect 1830 2759 1836 2760
rect 2014 2764 2020 2765
rect 2014 2760 2015 2764
rect 2019 2760 2020 2764
rect 2014 2759 2020 2760
rect 2214 2764 2220 2765
rect 2214 2760 2215 2764
rect 2219 2760 2220 2764
rect 2214 2759 2220 2760
rect 2406 2764 2412 2765
rect 2406 2760 2407 2764
rect 2411 2760 2412 2764
rect 2406 2759 2412 2760
rect 2582 2764 2588 2765
rect 2582 2760 2583 2764
rect 2587 2760 2588 2764
rect 2582 2759 2588 2760
rect 2750 2764 2756 2765
rect 2750 2760 2751 2764
rect 2755 2760 2756 2764
rect 2750 2759 2756 2760
rect 2910 2764 2916 2765
rect 2910 2760 2911 2764
rect 2915 2760 2916 2764
rect 2910 2759 2916 2760
rect 3070 2764 3076 2765
rect 3070 2760 3071 2764
rect 3075 2760 3076 2764
rect 3070 2759 3076 2760
rect 3230 2764 3236 2765
rect 3230 2760 3231 2764
rect 3235 2760 3236 2764
rect 3230 2759 3236 2760
rect 3366 2764 3372 2765
rect 3366 2760 3367 2764
rect 3371 2760 3372 2764
rect 3462 2763 3463 2767
rect 3467 2763 3468 2767
rect 3462 2762 3468 2763
rect 3366 2759 3372 2760
rect 1606 2758 1612 2759
rect 1598 2754 1604 2755
rect 1766 2755 1772 2756
rect 110 2750 116 2751
rect 134 2752 140 2753
rect 134 2748 135 2752
rect 139 2748 140 2752
rect 134 2747 140 2748
rect 246 2752 252 2753
rect 246 2748 247 2752
rect 251 2748 252 2752
rect 246 2747 252 2748
rect 390 2752 396 2753
rect 390 2748 391 2752
rect 395 2748 396 2752
rect 390 2747 396 2748
rect 542 2752 548 2753
rect 542 2748 543 2752
rect 547 2748 548 2752
rect 542 2747 548 2748
rect 694 2752 700 2753
rect 694 2748 695 2752
rect 699 2748 700 2752
rect 694 2747 700 2748
rect 854 2752 860 2753
rect 854 2748 855 2752
rect 859 2748 860 2752
rect 854 2747 860 2748
rect 1022 2752 1028 2753
rect 1022 2748 1023 2752
rect 1027 2748 1028 2752
rect 1022 2747 1028 2748
rect 1190 2752 1196 2753
rect 1190 2748 1191 2752
rect 1195 2748 1196 2752
rect 1190 2747 1196 2748
rect 1358 2752 1364 2753
rect 1358 2748 1359 2752
rect 1363 2748 1364 2752
rect 1358 2747 1364 2748
rect 1526 2752 1532 2753
rect 1526 2748 1527 2752
rect 1531 2748 1532 2752
rect 1526 2747 1532 2748
rect 1670 2752 1676 2753
rect 1670 2748 1671 2752
rect 1675 2748 1676 2752
rect 1766 2751 1767 2755
rect 1771 2751 1772 2755
rect 1766 2750 1772 2751
rect 1670 2747 1676 2748
rect 298 2715 304 2716
rect 298 2711 299 2715
rect 303 2714 304 2715
rect 622 2715 628 2716
rect 622 2714 623 2715
rect 303 2712 623 2714
rect 303 2711 304 2712
rect 298 2710 304 2711
rect 622 2711 623 2712
rect 627 2711 628 2715
rect 622 2710 628 2711
rect 2038 2704 2044 2705
rect 1806 2701 1812 2702
rect 246 2700 252 2701
rect 110 2697 116 2698
rect 110 2693 111 2697
rect 115 2693 116 2697
rect 246 2696 247 2700
rect 251 2696 252 2700
rect 246 2695 252 2696
rect 358 2700 364 2701
rect 358 2696 359 2700
rect 363 2696 364 2700
rect 358 2695 364 2696
rect 478 2700 484 2701
rect 478 2696 479 2700
rect 483 2696 484 2700
rect 478 2695 484 2696
rect 614 2700 620 2701
rect 614 2696 615 2700
rect 619 2696 620 2700
rect 614 2695 620 2696
rect 758 2700 764 2701
rect 758 2696 759 2700
rect 763 2696 764 2700
rect 758 2695 764 2696
rect 910 2700 916 2701
rect 910 2696 911 2700
rect 915 2696 916 2700
rect 910 2695 916 2696
rect 1062 2700 1068 2701
rect 1062 2696 1063 2700
rect 1067 2696 1068 2700
rect 1062 2695 1068 2696
rect 1214 2700 1220 2701
rect 1214 2696 1215 2700
rect 1219 2696 1220 2700
rect 1214 2695 1220 2696
rect 1374 2700 1380 2701
rect 1374 2696 1375 2700
rect 1379 2696 1380 2700
rect 1374 2695 1380 2696
rect 1534 2700 1540 2701
rect 1534 2696 1535 2700
rect 1539 2696 1540 2700
rect 1534 2695 1540 2696
rect 1670 2700 1676 2701
rect 1670 2696 1671 2700
rect 1675 2696 1676 2700
rect 1670 2695 1676 2696
rect 1766 2697 1772 2698
rect 110 2692 116 2693
rect 1766 2693 1767 2697
rect 1771 2693 1772 2697
rect 1806 2697 1807 2701
rect 1811 2697 1812 2701
rect 2038 2700 2039 2704
rect 2043 2700 2044 2704
rect 2038 2699 2044 2700
rect 2158 2704 2164 2705
rect 2158 2700 2159 2704
rect 2163 2700 2164 2704
rect 2158 2699 2164 2700
rect 2278 2704 2284 2705
rect 2278 2700 2279 2704
rect 2283 2700 2284 2704
rect 2278 2699 2284 2700
rect 2406 2704 2412 2705
rect 2406 2700 2407 2704
rect 2411 2700 2412 2704
rect 2406 2699 2412 2700
rect 2542 2704 2548 2705
rect 2542 2700 2543 2704
rect 2547 2700 2548 2704
rect 2542 2699 2548 2700
rect 2686 2704 2692 2705
rect 2686 2700 2687 2704
rect 2691 2700 2692 2704
rect 2686 2699 2692 2700
rect 2846 2704 2852 2705
rect 2846 2700 2847 2704
rect 2851 2700 2852 2704
rect 2846 2699 2852 2700
rect 3022 2704 3028 2705
rect 3022 2700 3023 2704
rect 3027 2700 3028 2704
rect 3022 2699 3028 2700
rect 3206 2704 3212 2705
rect 3206 2700 3207 2704
rect 3211 2700 3212 2704
rect 3206 2699 3212 2700
rect 3366 2704 3372 2705
rect 3366 2700 3367 2704
rect 3371 2700 3372 2704
rect 3366 2699 3372 2700
rect 3462 2701 3468 2702
rect 1806 2696 1812 2697
rect 3462 2697 3463 2701
rect 3467 2697 3468 2701
rect 3462 2696 3468 2697
rect 1766 2692 1772 2693
rect 2110 2695 2116 2696
rect 318 2691 324 2692
rect 318 2687 319 2691
rect 323 2687 324 2691
rect 318 2686 324 2687
rect 430 2691 436 2692
rect 430 2687 431 2691
rect 435 2687 436 2691
rect 430 2686 436 2687
rect 550 2691 556 2692
rect 550 2687 551 2691
rect 555 2687 556 2691
rect 550 2686 556 2687
rect 686 2691 692 2692
rect 686 2687 687 2691
rect 691 2687 692 2691
rect 686 2686 692 2687
rect 694 2691 700 2692
rect 694 2687 695 2691
rect 699 2690 700 2691
rect 902 2691 908 2692
rect 699 2688 801 2690
rect 699 2687 700 2688
rect 694 2686 700 2687
rect 902 2687 903 2691
rect 907 2690 908 2691
rect 1134 2691 1140 2692
rect 907 2688 953 2690
rect 907 2687 908 2688
rect 902 2686 908 2687
rect 1134 2687 1135 2691
rect 1139 2687 1140 2691
rect 1134 2686 1140 2687
rect 1175 2691 1181 2692
rect 1175 2687 1176 2691
rect 1180 2690 1181 2691
rect 1446 2691 1452 2692
rect 1180 2688 1257 2690
rect 1180 2687 1181 2688
rect 1175 2686 1181 2687
rect 1446 2687 1447 2691
rect 1451 2687 1452 2691
rect 1446 2686 1452 2687
rect 1606 2691 1612 2692
rect 1606 2687 1607 2691
rect 1611 2687 1612 2691
rect 1606 2686 1612 2687
rect 1638 2691 1644 2692
rect 1638 2687 1639 2691
rect 1643 2690 1644 2691
rect 2110 2691 2111 2695
rect 2115 2691 2116 2695
rect 2110 2690 2116 2691
rect 2230 2695 2236 2696
rect 2230 2691 2231 2695
rect 2235 2691 2236 2695
rect 2230 2690 2236 2691
rect 2350 2695 2356 2696
rect 2350 2691 2351 2695
rect 2355 2691 2356 2695
rect 2350 2690 2356 2691
rect 2470 2695 2476 2696
rect 2470 2691 2471 2695
rect 2475 2691 2476 2695
rect 2470 2690 2476 2691
rect 2614 2695 2620 2696
rect 2614 2691 2615 2695
rect 2619 2691 2620 2695
rect 2766 2695 2772 2696
rect 2766 2694 2767 2695
rect 2761 2692 2767 2694
rect 2614 2690 2620 2691
rect 2766 2691 2767 2692
rect 2771 2691 2772 2695
rect 2766 2690 2772 2691
rect 2774 2695 2780 2696
rect 2774 2691 2775 2695
rect 2779 2694 2780 2695
rect 3094 2695 3100 2696
rect 2779 2692 2889 2694
rect 2779 2691 2780 2692
rect 2774 2690 2780 2691
rect 3094 2691 3095 2695
rect 3099 2691 3100 2695
rect 3094 2690 3100 2691
rect 3102 2695 3108 2696
rect 3102 2691 3103 2695
rect 3107 2694 3108 2695
rect 3430 2695 3436 2696
rect 3107 2692 3249 2694
rect 3107 2691 3108 2692
rect 3102 2690 3108 2691
rect 3430 2691 3431 2695
rect 3435 2691 3436 2695
rect 3430 2690 3436 2691
rect 1643 2688 1713 2690
rect 1643 2687 1644 2688
rect 1638 2686 1644 2687
rect 2038 2685 2044 2686
rect 1806 2684 1812 2685
rect 246 2681 252 2682
rect 110 2680 116 2681
rect 110 2676 111 2680
rect 115 2676 116 2680
rect 246 2677 247 2681
rect 251 2677 252 2681
rect 246 2676 252 2677
rect 358 2681 364 2682
rect 358 2677 359 2681
rect 363 2677 364 2681
rect 358 2676 364 2677
rect 478 2681 484 2682
rect 478 2677 479 2681
rect 483 2677 484 2681
rect 478 2676 484 2677
rect 614 2681 620 2682
rect 614 2677 615 2681
rect 619 2677 620 2681
rect 614 2676 620 2677
rect 758 2681 764 2682
rect 758 2677 759 2681
rect 763 2677 764 2681
rect 758 2676 764 2677
rect 910 2681 916 2682
rect 910 2677 911 2681
rect 915 2677 916 2681
rect 910 2676 916 2677
rect 1062 2681 1068 2682
rect 1062 2677 1063 2681
rect 1067 2677 1068 2681
rect 1062 2676 1068 2677
rect 1214 2681 1220 2682
rect 1214 2677 1215 2681
rect 1219 2677 1220 2681
rect 1214 2676 1220 2677
rect 1374 2681 1380 2682
rect 1374 2677 1375 2681
rect 1379 2677 1380 2681
rect 1374 2676 1380 2677
rect 1534 2681 1540 2682
rect 1534 2677 1535 2681
rect 1539 2677 1540 2681
rect 1534 2676 1540 2677
rect 1670 2681 1676 2682
rect 1670 2677 1671 2681
rect 1675 2677 1676 2681
rect 1670 2676 1676 2677
rect 1766 2680 1772 2681
rect 1766 2676 1767 2680
rect 1771 2676 1772 2680
rect 1806 2680 1807 2684
rect 1811 2680 1812 2684
rect 2038 2681 2039 2685
rect 2043 2681 2044 2685
rect 2038 2680 2044 2681
rect 2158 2685 2164 2686
rect 2158 2681 2159 2685
rect 2163 2681 2164 2685
rect 2158 2680 2164 2681
rect 2278 2685 2284 2686
rect 2278 2681 2279 2685
rect 2283 2681 2284 2685
rect 2278 2680 2284 2681
rect 2406 2685 2412 2686
rect 2406 2681 2407 2685
rect 2411 2681 2412 2685
rect 2406 2680 2412 2681
rect 2542 2685 2548 2686
rect 2542 2681 2543 2685
rect 2547 2681 2548 2685
rect 2542 2680 2548 2681
rect 2686 2685 2692 2686
rect 2686 2681 2687 2685
rect 2691 2681 2692 2685
rect 2686 2680 2692 2681
rect 2846 2685 2852 2686
rect 2846 2681 2847 2685
rect 2851 2681 2852 2685
rect 2846 2680 2852 2681
rect 3022 2685 3028 2686
rect 3022 2681 3023 2685
rect 3027 2681 3028 2685
rect 3022 2680 3028 2681
rect 3206 2685 3212 2686
rect 3206 2681 3207 2685
rect 3211 2681 3212 2685
rect 3206 2680 3212 2681
rect 3366 2685 3372 2686
rect 3366 2681 3367 2685
rect 3371 2681 3372 2685
rect 3366 2680 3372 2681
rect 3462 2684 3468 2685
rect 3462 2680 3463 2684
rect 3467 2680 3468 2684
rect 1806 2679 1812 2680
rect 3462 2679 3468 2680
rect 110 2675 116 2676
rect 1766 2675 1772 2676
rect 2087 2667 2093 2668
rect 295 2663 304 2664
rect 295 2659 296 2663
rect 303 2659 304 2663
rect 295 2658 304 2659
rect 318 2663 324 2664
rect 318 2659 319 2663
rect 323 2662 324 2663
rect 407 2663 413 2664
rect 407 2662 408 2663
rect 323 2660 408 2662
rect 323 2659 324 2660
rect 318 2658 324 2659
rect 407 2659 408 2660
rect 412 2659 413 2663
rect 407 2658 413 2659
rect 430 2663 436 2664
rect 430 2659 431 2663
rect 435 2662 436 2663
rect 527 2663 533 2664
rect 527 2662 528 2663
rect 435 2660 528 2662
rect 435 2659 436 2660
rect 430 2658 436 2659
rect 527 2659 528 2660
rect 532 2659 533 2663
rect 527 2658 533 2659
rect 550 2663 556 2664
rect 550 2659 551 2663
rect 555 2662 556 2663
rect 663 2663 669 2664
rect 663 2662 664 2663
rect 555 2660 664 2662
rect 555 2659 556 2660
rect 550 2658 556 2659
rect 663 2659 664 2660
rect 668 2659 669 2663
rect 663 2658 669 2659
rect 686 2663 692 2664
rect 686 2659 687 2663
rect 691 2662 692 2663
rect 807 2663 813 2664
rect 807 2662 808 2663
rect 691 2660 808 2662
rect 691 2659 692 2660
rect 686 2658 692 2659
rect 807 2659 808 2660
rect 812 2659 813 2663
rect 807 2658 813 2659
rect 959 2663 965 2664
rect 959 2659 960 2663
rect 964 2662 965 2663
rect 1054 2663 1060 2664
rect 964 2660 1050 2662
rect 964 2659 965 2660
rect 959 2658 965 2659
rect 1048 2654 1050 2660
rect 1054 2659 1055 2663
rect 1059 2662 1060 2663
rect 1111 2663 1117 2664
rect 1111 2662 1112 2663
rect 1059 2660 1112 2662
rect 1059 2659 1060 2660
rect 1054 2658 1060 2659
rect 1111 2659 1112 2660
rect 1116 2659 1117 2663
rect 1111 2658 1117 2659
rect 1134 2663 1140 2664
rect 1134 2659 1135 2663
rect 1139 2662 1140 2663
rect 1263 2663 1269 2664
rect 1263 2662 1264 2663
rect 1139 2660 1264 2662
rect 1139 2659 1140 2660
rect 1134 2658 1140 2659
rect 1263 2659 1264 2660
rect 1268 2659 1269 2663
rect 1263 2658 1269 2659
rect 1423 2663 1429 2664
rect 1423 2659 1424 2663
rect 1428 2662 1429 2663
rect 1583 2663 1589 2664
rect 1428 2660 1570 2662
rect 1428 2659 1429 2660
rect 1423 2658 1429 2659
rect 1175 2655 1181 2656
rect 1175 2654 1176 2655
rect 1048 2652 1176 2654
rect 694 2651 700 2652
rect 694 2650 695 2651
rect 528 2648 695 2650
rect 511 2643 517 2644
rect 511 2639 512 2643
rect 516 2642 517 2643
rect 528 2642 530 2648
rect 694 2647 695 2648
rect 699 2647 700 2651
rect 1175 2651 1176 2652
rect 1180 2651 1181 2655
rect 1568 2654 1570 2660
rect 1583 2659 1584 2663
rect 1588 2662 1589 2663
rect 1598 2663 1604 2664
rect 1598 2662 1599 2663
rect 1588 2660 1599 2662
rect 1588 2659 1589 2660
rect 1583 2658 1589 2659
rect 1598 2659 1599 2660
rect 1603 2659 1604 2663
rect 1598 2658 1604 2659
rect 1606 2663 1612 2664
rect 1606 2659 1607 2663
rect 1611 2662 1612 2663
rect 1719 2663 1725 2664
rect 1719 2662 1720 2663
rect 1611 2660 1720 2662
rect 1611 2659 1612 2660
rect 1606 2658 1612 2659
rect 1719 2659 1720 2660
rect 1724 2659 1725 2663
rect 2087 2663 2088 2667
rect 2092 2666 2093 2667
rect 2110 2667 2116 2668
rect 2092 2664 2106 2666
rect 2092 2663 2093 2664
rect 2087 2662 2093 2663
rect 1719 2658 1725 2659
rect 2104 2658 2106 2664
rect 2110 2663 2111 2667
rect 2115 2666 2116 2667
rect 2207 2667 2213 2668
rect 2207 2666 2208 2667
rect 2115 2664 2208 2666
rect 2115 2663 2116 2664
rect 2110 2662 2116 2663
rect 2207 2663 2208 2664
rect 2212 2663 2213 2667
rect 2207 2662 2213 2663
rect 2230 2667 2236 2668
rect 2230 2663 2231 2667
rect 2235 2666 2236 2667
rect 2327 2667 2333 2668
rect 2327 2666 2328 2667
rect 2235 2664 2328 2666
rect 2235 2663 2236 2664
rect 2230 2662 2236 2663
rect 2327 2663 2328 2664
rect 2332 2663 2333 2667
rect 2327 2662 2333 2663
rect 2350 2667 2356 2668
rect 2350 2663 2351 2667
rect 2355 2666 2356 2667
rect 2455 2667 2461 2668
rect 2455 2666 2456 2667
rect 2355 2664 2456 2666
rect 2355 2663 2356 2664
rect 2350 2662 2356 2663
rect 2455 2663 2456 2664
rect 2460 2663 2461 2667
rect 2455 2662 2461 2663
rect 2591 2667 2597 2668
rect 2591 2663 2592 2667
rect 2596 2666 2597 2667
rect 2614 2667 2620 2668
rect 2596 2664 2610 2666
rect 2596 2663 2597 2664
rect 2591 2662 2597 2663
rect 2262 2659 2268 2660
rect 2262 2658 2263 2659
rect 2104 2656 2263 2658
rect 1638 2655 1644 2656
rect 1638 2654 1639 2655
rect 1568 2652 1639 2654
rect 1175 2650 1181 2651
rect 1638 2651 1639 2652
rect 1643 2651 1644 2655
rect 2262 2655 2263 2656
rect 2267 2655 2268 2659
rect 2608 2658 2610 2664
rect 2614 2663 2615 2667
rect 2619 2666 2620 2667
rect 2735 2667 2741 2668
rect 2735 2666 2736 2667
rect 2619 2664 2736 2666
rect 2619 2663 2620 2664
rect 2614 2662 2620 2663
rect 2735 2663 2736 2664
rect 2740 2663 2741 2667
rect 2735 2662 2741 2663
rect 2895 2667 2901 2668
rect 2895 2663 2896 2667
rect 2900 2666 2901 2667
rect 2982 2667 2988 2668
rect 2900 2664 2978 2666
rect 2900 2663 2901 2664
rect 2895 2662 2901 2663
rect 2774 2659 2780 2660
rect 2774 2658 2775 2659
rect 2608 2656 2775 2658
rect 2262 2654 2268 2655
rect 2774 2655 2775 2656
rect 2779 2655 2780 2659
rect 2976 2658 2978 2664
rect 2982 2663 2983 2667
rect 2987 2666 2988 2667
rect 3071 2667 3077 2668
rect 3071 2666 3072 2667
rect 2987 2664 3072 2666
rect 2987 2663 2988 2664
rect 2982 2662 2988 2663
rect 3071 2663 3072 2664
rect 3076 2663 3077 2667
rect 3071 2662 3077 2663
rect 3094 2667 3100 2668
rect 3094 2663 3095 2667
rect 3099 2666 3100 2667
rect 3255 2667 3261 2668
rect 3255 2666 3256 2667
rect 3099 2664 3256 2666
rect 3099 2663 3100 2664
rect 3094 2662 3100 2663
rect 3255 2663 3256 2664
rect 3260 2663 3261 2667
rect 3255 2662 3261 2663
rect 3415 2667 3421 2668
rect 3415 2663 3416 2667
rect 3420 2666 3421 2667
rect 3438 2667 3444 2668
rect 3438 2666 3439 2667
rect 3420 2664 3439 2666
rect 3420 2663 3421 2664
rect 3415 2662 3421 2663
rect 3438 2663 3439 2664
rect 3443 2663 3444 2667
rect 3438 2662 3444 2663
rect 3102 2659 3108 2660
rect 3102 2658 3103 2659
rect 2976 2656 3103 2658
rect 2774 2654 2780 2655
rect 3102 2655 3103 2656
rect 3107 2655 3108 2659
rect 3102 2654 3108 2655
rect 1638 2650 1644 2651
rect 3138 2651 3144 2652
rect 3138 2650 3139 2651
rect 694 2646 700 2647
rect 2736 2648 3139 2650
rect 516 2640 530 2642
rect 534 2643 540 2644
rect 516 2639 517 2640
rect 511 2638 517 2639
rect 534 2639 535 2643
rect 539 2642 540 2643
rect 599 2643 605 2644
rect 599 2642 600 2643
rect 539 2640 600 2642
rect 539 2639 540 2640
rect 534 2638 540 2639
rect 599 2639 600 2640
rect 604 2639 605 2643
rect 599 2638 605 2639
rect 622 2643 628 2644
rect 622 2639 623 2643
rect 627 2642 628 2643
rect 687 2643 693 2644
rect 687 2642 688 2643
rect 627 2640 688 2642
rect 627 2639 628 2640
rect 622 2638 628 2639
rect 687 2639 688 2640
rect 692 2639 693 2643
rect 687 2638 693 2639
rect 710 2643 716 2644
rect 710 2639 711 2643
rect 715 2642 716 2643
rect 791 2643 797 2644
rect 791 2642 792 2643
rect 715 2640 792 2642
rect 715 2639 716 2640
rect 710 2638 716 2639
rect 791 2639 792 2640
rect 796 2639 797 2643
rect 791 2638 797 2639
rect 814 2643 820 2644
rect 814 2639 815 2643
rect 819 2642 820 2643
rect 903 2643 909 2644
rect 903 2642 904 2643
rect 819 2640 904 2642
rect 819 2639 820 2640
rect 814 2638 820 2639
rect 903 2639 904 2640
rect 908 2639 909 2643
rect 903 2638 909 2639
rect 1031 2643 1037 2644
rect 1031 2639 1032 2643
rect 1036 2642 1037 2643
rect 1106 2643 1112 2644
rect 1106 2642 1107 2643
rect 1036 2640 1107 2642
rect 1036 2639 1037 2640
rect 1031 2638 1037 2639
rect 1106 2639 1107 2640
rect 1111 2639 1112 2643
rect 1106 2638 1112 2639
rect 1175 2643 1181 2644
rect 1175 2639 1176 2643
rect 1180 2642 1181 2643
rect 1206 2643 1212 2644
rect 1206 2642 1207 2643
rect 1180 2640 1207 2642
rect 1180 2639 1181 2640
rect 1175 2638 1181 2639
rect 1206 2639 1207 2640
rect 1211 2639 1212 2643
rect 1206 2638 1212 2639
rect 1294 2643 1300 2644
rect 1294 2639 1295 2643
rect 1299 2642 1300 2643
rect 1327 2643 1333 2644
rect 1327 2642 1328 2643
rect 1299 2640 1328 2642
rect 1299 2639 1300 2640
rect 1294 2638 1300 2639
rect 1327 2639 1328 2640
rect 1332 2639 1333 2643
rect 1327 2638 1333 2639
rect 1446 2643 1452 2644
rect 1446 2639 1447 2643
rect 1451 2642 1452 2643
rect 1487 2643 1493 2644
rect 1487 2642 1488 2643
rect 1451 2640 1488 2642
rect 1451 2639 1452 2640
rect 1446 2638 1452 2639
rect 1487 2639 1488 2640
rect 1492 2639 1493 2643
rect 1487 2638 1493 2639
rect 1510 2643 1516 2644
rect 1510 2639 1511 2643
rect 1515 2642 1516 2643
rect 1655 2643 1661 2644
rect 1655 2642 1656 2643
rect 1515 2640 1656 2642
rect 1515 2639 1516 2640
rect 1510 2638 1516 2639
rect 1655 2639 1656 2640
rect 1660 2639 1661 2643
rect 1655 2638 1661 2639
rect 1902 2643 1908 2644
rect 1902 2639 1903 2643
rect 1907 2642 1908 2643
rect 1919 2643 1925 2644
rect 1919 2642 1920 2643
rect 1907 2640 1920 2642
rect 1907 2639 1908 2640
rect 1902 2638 1908 2639
rect 1919 2639 1920 2640
rect 1924 2639 1925 2643
rect 1919 2638 1925 2639
rect 1942 2643 1948 2644
rect 1942 2639 1943 2643
rect 1947 2642 1948 2643
rect 2015 2643 2021 2644
rect 2015 2642 2016 2643
rect 1947 2640 2016 2642
rect 1947 2639 1948 2640
rect 1942 2638 1948 2639
rect 2015 2639 2016 2640
rect 2020 2639 2021 2643
rect 2015 2638 2021 2639
rect 2062 2643 2068 2644
rect 2062 2639 2063 2643
rect 2067 2642 2068 2643
rect 2119 2643 2125 2644
rect 2119 2642 2120 2643
rect 2067 2640 2120 2642
rect 2067 2639 2068 2640
rect 2062 2638 2068 2639
rect 2119 2639 2120 2640
rect 2124 2639 2125 2643
rect 2119 2638 2125 2639
rect 2142 2643 2148 2644
rect 2142 2639 2143 2643
rect 2147 2642 2148 2643
rect 2231 2643 2237 2644
rect 2231 2642 2232 2643
rect 2147 2640 2232 2642
rect 2147 2639 2148 2640
rect 2142 2638 2148 2639
rect 2231 2639 2232 2640
rect 2236 2639 2237 2643
rect 2231 2638 2237 2639
rect 2254 2643 2260 2644
rect 2254 2639 2255 2643
rect 2259 2642 2260 2643
rect 2343 2643 2349 2644
rect 2343 2642 2344 2643
rect 2259 2640 2344 2642
rect 2259 2639 2260 2640
rect 2254 2638 2260 2639
rect 2343 2639 2344 2640
rect 2348 2639 2349 2643
rect 2343 2638 2349 2639
rect 2479 2643 2485 2644
rect 2479 2639 2480 2643
rect 2484 2642 2485 2643
rect 2510 2643 2516 2644
rect 2510 2642 2511 2643
rect 2484 2640 2511 2642
rect 2484 2639 2485 2640
rect 2479 2638 2485 2639
rect 2510 2639 2511 2640
rect 2515 2639 2516 2643
rect 2510 2638 2516 2639
rect 2631 2643 2637 2644
rect 2631 2639 2632 2643
rect 2636 2642 2637 2643
rect 2736 2642 2738 2648
rect 3138 2647 3139 2648
rect 3143 2647 3144 2651
rect 3138 2646 3144 2647
rect 2636 2640 2738 2642
rect 2766 2643 2772 2644
rect 2636 2639 2637 2640
rect 2631 2638 2637 2639
rect 2766 2639 2767 2643
rect 2771 2642 2772 2643
rect 2807 2643 2813 2644
rect 2807 2642 2808 2643
rect 2771 2640 2808 2642
rect 2771 2639 2772 2640
rect 2766 2638 2772 2639
rect 2807 2639 2808 2640
rect 2812 2639 2813 2643
rect 2807 2638 2813 2639
rect 2830 2643 2836 2644
rect 2830 2639 2831 2643
rect 2835 2642 2836 2643
rect 3007 2643 3013 2644
rect 3007 2642 3008 2643
rect 2835 2640 3008 2642
rect 2835 2639 2836 2640
rect 2830 2638 2836 2639
rect 3007 2639 3008 2640
rect 3012 2639 3013 2643
rect 3007 2638 3013 2639
rect 3030 2643 3036 2644
rect 3030 2639 3031 2643
rect 3035 2642 3036 2643
rect 3215 2643 3221 2644
rect 3215 2642 3216 2643
rect 3035 2640 3216 2642
rect 3035 2639 3036 2640
rect 3030 2638 3036 2639
rect 3215 2639 3216 2640
rect 3220 2639 3221 2643
rect 3215 2638 3221 2639
rect 3415 2643 3421 2644
rect 3415 2639 3416 2643
rect 3420 2642 3421 2643
rect 3430 2643 3436 2644
rect 3430 2642 3431 2643
rect 3420 2640 3431 2642
rect 3420 2639 3421 2640
rect 3415 2638 3421 2639
rect 3430 2639 3431 2640
rect 3435 2639 3436 2643
rect 3430 2638 3436 2639
rect 110 2628 116 2629
rect 1766 2628 1772 2629
rect 110 2624 111 2628
rect 115 2624 116 2628
rect 110 2623 116 2624
rect 462 2627 468 2628
rect 462 2623 463 2627
rect 467 2623 468 2627
rect 462 2622 468 2623
rect 550 2627 556 2628
rect 550 2623 551 2627
rect 555 2623 556 2627
rect 550 2622 556 2623
rect 638 2627 644 2628
rect 638 2623 639 2627
rect 643 2623 644 2627
rect 638 2622 644 2623
rect 742 2627 748 2628
rect 742 2623 743 2627
rect 747 2623 748 2627
rect 742 2622 748 2623
rect 854 2627 860 2628
rect 854 2623 855 2627
rect 859 2623 860 2627
rect 854 2622 860 2623
rect 982 2627 988 2628
rect 982 2623 983 2627
rect 987 2623 988 2627
rect 982 2622 988 2623
rect 1126 2627 1132 2628
rect 1126 2623 1127 2627
rect 1131 2623 1132 2627
rect 1126 2622 1132 2623
rect 1278 2627 1284 2628
rect 1278 2623 1279 2627
rect 1283 2623 1284 2627
rect 1278 2622 1284 2623
rect 1438 2627 1444 2628
rect 1438 2623 1439 2627
rect 1443 2623 1444 2627
rect 1438 2622 1444 2623
rect 1606 2627 1612 2628
rect 1606 2623 1607 2627
rect 1611 2623 1612 2627
rect 1766 2624 1767 2628
rect 1771 2624 1772 2628
rect 1766 2623 1772 2624
rect 1806 2628 1812 2629
rect 3462 2628 3468 2629
rect 1806 2624 1807 2628
rect 1811 2624 1812 2628
rect 1806 2623 1812 2624
rect 1870 2627 1876 2628
rect 1870 2623 1871 2627
rect 1875 2623 1876 2627
rect 1606 2622 1612 2623
rect 1870 2622 1876 2623
rect 1966 2627 1972 2628
rect 1966 2623 1967 2627
rect 1971 2623 1972 2627
rect 1966 2622 1972 2623
rect 2070 2627 2076 2628
rect 2070 2623 2071 2627
rect 2075 2623 2076 2627
rect 2070 2622 2076 2623
rect 2182 2627 2188 2628
rect 2182 2623 2183 2627
rect 2187 2623 2188 2627
rect 2182 2622 2188 2623
rect 2294 2627 2300 2628
rect 2294 2623 2295 2627
rect 2299 2623 2300 2627
rect 2294 2622 2300 2623
rect 2430 2627 2436 2628
rect 2430 2623 2431 2627
rect 2435 2623 2436 2627
rect 2430 2622 2436 2623
rect 2582 2627 2588 2628
rect 2582 2623 2583 2627
rect 2587 2623 2588 2627
rect 2582 2622 2588 2623
rect 2758 2627 2764 2628
rect 2758 2623 2759 2627
rect 2763 2623 2764 2627
rect 2758 2622 2764 2623
rect 2958 2627 2964 2628
rect 2958 2623 2959 2627
rect 2963 2623 2964 2627
rect 2958 2622 2964 2623
rect 3166 2627 3172 2628
rect 3166 2623 3167 2627
rect 3171 2623 3172 2627
rect 3166 2622 3172 2623
rect 3366 2627 3372 2628
rect 3366 2623 3367 2627
rect 3371 2623 3372 2627
rect 3462 2624 3463 2628
rect 3467 2624 3468 2628
rect 3462 2623 3468 2624
rect 3366 2622 3372 2623
rect 534 2619 540 2620
rect 534 2615 535 2619
rect 539 2615 540 2619
rect 534 2614 540 2615
rect 622 2619 628 2620
rect 622 2615 623 2619
rect 627 2615 628 2619
rect 622 2614 628 2615
rect 710 2619 716 2620
rect 710 2615 711 2619
rect 715 2615 716 2619
rect 710 2614 716 2615
rect 814 2619 820 2620
rect 814 2615 815 2619
rect 819 2615 820 2619
rect 814 2614 820 2615
rect 822 2619 828 2620
rect 822 2615 823 2619
rect 827 2618 828 2619
rect 1054 2619 1060 2620
rect 827 2616 897 2618
rect 827 2615 828 2616
rect 822 2614 828 2615
rect 1054 2615 1055 2619
rect 1059 2615 1060 2619
rect 1054 2614 1060 2615
rect 1106 2619 1112 2620
rect 1106 2615 1107 2619
rect 1111 2618 1112 2619
rect 1206 2619 1212 2620
rect 1111 2616 1169 2618
rect 1111 2615 1112 2616
rect 1106 2614 1112 2615
rect 1206 2615 1207 2619
rect 1211 2618 1212 2619
rect 1510 2619 1516 2620
rect 1211 2616 1321 2618
rect 1211 2615 1212 2616
rect 1206 2614 1212 2615
rect 1510 2615 1511 2619
rect 1515 2615 1516 2619
rect 1942 2619 1948 2620
rect 1510 2614 1516 2615
rect 1678 2615 1684 2616
rect 110 2611 116 2612
rect 110 2607 111 2611
rect 115 2607 116 2611
rect 1678 2611 1679 2615
rect 1683 2611 1684 2615
rect 1942 2615 1943 2619
rect 1947 2615 1948 2619
rect 2062 2619 2068 2620
rect 2062 2618 2063 2619
rect 2041 2616 2063 2618
rect 1942 2614 1948 2615
rect 2062 2615 2063 2616
rect 2067 2615 2068 2619
rect 2062 2614 2068 2615
rect 2142 2619 2148 2620
rect 2142 2615 2143 2619
rect 2147 2615 2148 2619
rect 2142 2614 2148 2615
rect 2254 2619 2260 2620
rect 2254 2615 2255 2619
rect 2259 2615 2260 2619
rect 2254 2614 2260 2615
rect 2262 2619 2268 2620
rect 2262 2615 2263 2619
rect 2267 2618 2268 2619
rect 2394 2619 2400 2620
rect 2267 2616 2337 2618
rect 2267 2615 2268 2616
rect 2262 2614 2268 2615
rect 2394 2615 2395 2619
rect 2399 2618 2400 2619
rect 2510 2619 2516 2620
rect 2399 2616 2473 2618
rect 2399 2615 2400 2616
rect 2394 2614 2400 2615
rect 2510 2615 2511 2619
rect 2515 2618 2516 2619
rect 2830 2619 2836 2620
rect 2515 2616 2625 2618
rect 2515 2615 2516 2616
rect 2510 2614 2516 2615
rect 2830 2615 2831 2619
rect 2835 2615 2836 2619
rect 2830 2614 2836 2615
rect 3030 2619 3036 2620
rect 3030 2615 3031 2619
rect 3035 2615 3036 2619
rect 3030 2614 3036 2615
rect 3138 2619 3144 2620
rect 3138 2615 3139 2619
rect 3143 2618 3144 2619
rect 3143 2616 3209 2618
rect 3143 2615 3144 2616
rect 3138 2614 3144 2615
rect 3438 2615 3444 2616
rect 1678 2610 1684 2611
rect 1766 2611 1772 2612
rect 110 2606 116 2607
rect 462 2608 468 2609
rect 462 2604 463 2608
rect 467 2604 468 2608
rect 462 2603 468 2604
rect 550 2608 556 2609
rect 550 2604 551 2608
rect 555 2604 556 2608
rect 550 2603 556 2604
rect 638 2608 644 2609
rect 638 2604 639 2608
rect 643 2604 644 2608
rect 638 2603 644 2604
rect 742 2608 748 2609
rect 742 2604 743 2608
rect 747 2604 748 2608
rect 742 2603 748 2604
rect 854 2608 860 2609
rect 854 2604 855 2608
rect 859 2604 860 2608
rect 854 2603 860 2604
rect 982 2608 988 2609
rect 982 2604 983 2608
rect 987 2604 988 2608
rect 982 2603 988 2604
rect 1126 2608 1132 2609
rect 1126 2604 1127 2608
rect 1131 2604 1132 2608
rect 1126 2603 1132 2604
rect 1278 2608 1284 2609
rect 1278 2604 1279 2608
rect 1283 2604 1284 2608
rect 1278 2603 1284 2604
rect 1438 2608 1444 2609
rect 1438 2604 1439 2608
rect 1443 2604 1444 2608
rect 1438 2603 1444 2604
rect 1606 2608 1612 2609
rect 1606 2604 1607 2608
rect 1611 2604 1612 2608
rect 1766 2607 1767 2611
rect 1771 2607 1772 2611
rect 1766 2606 1772 2607
rect 1806 2611 1812 2612
rect 1806 2607 1807 2611
rect 1811 2607 1812 2611
rect 3438 2611 3439 2615
rect 3443 2611 3444 2615
rect 3438 2610 3444 2611
rect 3462 2611 3468 2612
rect 1806 2606 1812 2607
rect 1870 2608 1876 2609
rect 1606 2603 1612 2604
rect 1870 2604 1871 2608
rect 1875 2604 1876 2608
rect 1870 2603 1876 2604
rect 1966 2608 1972 2609
rect 1966 2604 1967 2608
rect 1971 2604 1972 2608
rect 1966 2603 1972 2604
rect 2070 2608 2076 2609
rect 2070 2604 2071 2608
rect 2075 2604 2076 2608
rect 2070 2603 2076 2604
rect 2182 2608 2188 2609
rect 2182 2604 2183 2608
rect 2187 2604 2188 2608
rect 2182 2603 2188 2604
rect 2294 2608 2300 2609
rect 2294 2604 2295 2608
rect 2299 2604 2300 2608
rect 2294 2603 2300 2604
rect 2430 2608 2436 2609
rect 2430 2604 2431 2608
rect 2435 2604 2436 2608
rect 2430 2603 2436 2604
rect 2582 2608 2588 2609
rect 2582 2604 2583 2608
rect 2587 2604 2588 2608
rect 2582 2603 2588 2604
rect 2758 2608 2764 2609
rect 2758 2604 2759 2608
rect 2763 2604 2764 2608
rect 2758 2603 2764 2604
rect 2958 2608 2964 2609
rect 2958 2604 2959 2608
rect 2963 2604 2964 2608
rect 2958 2603 2964 2604
rect 3166 2608 3172 2609
rect 3166 2604 3167 2608
rect 3171 2604 3172 2608
rect 3166 2603 3172 2604
rect 3366 2608 3372 2609
rect 3366 2604 3367 2608
rect 3371 2604 3372 2608
rect 3462 2607 3463 2611
rect 3467 2607 3468 2611
rect 3462 2606 3468 2607
rect 3366 2603 3372 2604
rect 2578 2559 2584 2560
rect 502 2556 508 2557
rect 110 2553 116 2554
rect 110 2549 111 2553
rect 115 2549 116 2553
rect 502 2552 503 2556
rect 507 2552 508 2556
rect 502 2551 508 2552
rect 590 2556 596 2557
rect 590 2552 591 2556
rect 595 2552 596 2556
rect 590 2551 596 2552
rect 678 2556 684 2557
rect 678 2552 679 2556
rect 683 2552 684 2556
rect 678 2551 684 2552
rect 774 2556 780 2557
rect 774 2552 775 2556
rect 779 2552 780 2556
rect 774 2551 780 2552
rect 878 2556 884 2557
rect 878 2552 879 2556
rect 883 2552 884 2556
rect 878 2551 884 2552
rect 990 2556 996 2557
rect 990 2552 991 2556
rect 995 2552 996 2556
rect 990 2551 996 2552
rect 1102 2556 1108 2557
rect 1102 2552 1103 2556
rect 1107 2552 1108 2556
rect 1102 2551 1108 2552
rect 1222 2556 1228 2557
rect 1222 2552 1223 2556
rect 1227 2552 1228 2556
rect 1222 2551 1228 2552
rect 1350 2556 1356 2557
rect 1350 2552 1351 2556
rect 1355 2552 1356 2556
rect 1350 2551 1356 2552
rect 1478 2556 1484 2557
rect 1478 2552 1479 2556
rect 1483 2552 1484 2556
rect 1478 2551 1484 2552
rect 1606 2556 1612 2557
rect 1606 2552 1607 2556
rect 1611 2552 1612 2556
rect 2578 2555 2579 2559
rect 2583 2558 2584 2559
rect 2583 2556 2946 2558
rect 2583 2555 2584 2556
rect 2578 2554 2584 2555
rect 1606 2551 1612 2552
rect 1766 2553 1772 2554
rect 110 2548 116 2549
rect 1766 2549 1767 2553
rect 1771 2549 1772 2553
rect 1830 2552 1836 2553
rect 1766 2548 1772 2549
rect 1806 2549 1812 2550
rect 574 2547 580 2548
rect 574 2543 575 2547
rect 579 2543 580 2547
rect 574 2542 580 2543
rect 662 2547 668 2548
rect 662 2543 663 2547
rect 667 2543 668 2547
rect 662 2542 668 2543
rect 750 2547 756 2548
rect 750 2543 751 2547
rect 755 2543 756 2547
rect 750 2542 756 2543
rect 846 2547 852 2548
rect 846 2543 847 2547
rect 851 2543 852 2547
rect 846 2542 852 2543
rect 950 2547 956 2548
rect 950 2543 951 2547
rect 955 2543 956 2547
rect 950 2542 956 2543
rect 1062 2547 1068 2548
rect 1062 2543 1063 2547
rect 1067 2543 1068 2547
rect 1062 2542 1068 2543
rect 1174 2547 1180 2548
rect 1174 2543 1175 2547
rect 1179 2543 1180 2547
rect 1174 2542 1180 2543
rect 1294 2547 1300 2548
rect 1294 2543 1295 2547
rect 1299 2543 1300 2547
rect 1294 2542 1300 2543
rect 1422 2547 1428 2548
rect 1422 2543 1423 2547
rect 1427 2543 1428 2547
rect 1422 2542 1428 2543
rect 1430 2547 1436 2548
rect 1430 2543 1431 2547
rect 1435 2546 1436 2547
rect 1558 2547 1564 2548
rect 1435 2544 1521 2546
rect 1435 2543 1436 2544
rect 1430 2542 1436 2543
rect 1558 2543 1559 2547
rect 1563 2546 1564 2547
rect 1563 2544 1649 2546
rect 1806 2545 1807 2549
rect 1811 2545 1812 2549
rect 1830 2548 1831 2552
rect 1835 2548 1836 2552
rect 1830 2547 1836 2548
rect 1918 2552 1924 2553
rect 1918 2548 1919 2552
rect 1923 2548 1924 2552
rect 1918 2547 1924 2548
rect 2006 2552 2012 2553
rect 2006 2548 2007 2552
rect 2011 2548 2012 2552
rect 2006 2547 2012 2548
rect 2110 2552 2116 2553
rect 2110 2548 2111 2552
rect 2115 2548 2116 2552
rect 2110 2547 2116 2548
rect 2222 2552 2228 2553
rect 2222 2548 2223 2552
rect 2227 2548 2228 2552
rect 2222 2547 2228 2548
rect 2342 2552 2348 2553
rect 2342 2548 2343 2552
rect 2347 2548 2348 2552
rect 2342 2547 2348 2548
rect 2486 2552 2492 2553
rect 2486 2548 2487 2552
rect 2491 2548 2492 2552
rect 2486 2547 2492 2548
rect 2646 2552 2652 2553
rect 2646 2548 2647 2552
rect 2651 2548 2652 2552
rect 2646 2547 2652 2548
rect 2814 2552 2820 2553
rect 2814 2548 2815 2552
rect 2819 2548 2820 2552
rect 2814 2547 2820 2548
rect 1806 2544 1812 2545
rect 1563 2543 1564 2544
rect 1558 2542 1564 2543
rect 1902 2543 1908 2544
rect 1902 2539 1903 2543
rect 1907 2539 1908 2543
rect 1902 2538 1908 2539
rect 1910 2543 1916 2544
rect 1910 2539 1911 2543
rect 1915 2542 1916 2543
rect 1999 2543 2005 2544
rect 1915 2540 1961 2542
rect 1915 2539 1916 2540
rect 1910 2538 1916 2539
rect 1999 2539 2000 2543
rect 2004 2542 2005 2543
rect 2086 2543 2092 2544
rect 2004 2540 2049 2542
rect 2004 2539 2005 2540
rect 1999 2538 2005 2539
rect 2086 2539 2087 2543
rect 2091 2542 2092 2543
rect 2190 2543 2196 2544
rect 2091 2540 2153 2542
rect 2091 2539 2092 2540
rect 2086 2538 2092 2539
rect 2190 2539 2191 2543
rect 2195 2542 2196 2543
rect 2414 2543 2420 2544
rect 2195 2540 2265 2542
rect 2195 2539 2196 2540
rect 2190 2538 2196 2539
rect 2414 2539 2415 2543
rect 2419 2539 2420 2543
rect 2414 2538 2420 2539
rect 2558 2543 2564 2544
rect 2558 2539 2559 2543
rect 2563 2539 2564 2543
rect 2558 2538 2564 2539
rect 2718 2543 2724 2544
rect 2718 2539 2719 2543
rect 2723 2539 2724 2543
rect 2718 2538 2724 2539
rect 2886 2543 2892 2544
rect 2886 2539 2887 2543
rect 2891 2539 2892 2543
rect 2944 2542 2946 2556
rect 2998 2552 3004 2553
rect 2998 2548 2999 2552
rect 3003 2548 3004 2552
rect 2998 2547 3004 2548
rect 3190 2552 3196 2553
rect 3190 2548 3191 2552
rect 3195 2548 3196 2552
rect 3190 2547 3196 2548
rect 3366 2552 3372 2553
rect 3366 2548 3367 2552
rect 3371 2548 3372 2552
rect 3366 2547 3372 2548
rect 3462 2549 3468 2550
rect 3462 2545 3463 2549
rect 3467 2545 3468 2549
rect 3462 2544 3468 2545
rect 3262 2543 3268 2544
rect 2944 2540 3041 2542
rect 2886 2538 2892 2539
rect 3262 2539 3263 2543
rect 3267 2539 3268 2543
rect 3262 2538 3268 2539
rect 3430 2543 3436 2544
rect 3430 2539 3431 2543
rect 3435 2539 3436 2543
rect 3430 2538 3436 2539
rect 502 2537 508 2538
rect 110 2536 116 2537
rect 110 2532 111 2536
rect 115 2532 116 2536
rect 502 2533 503 2537
rect 507 2533 508 2537
rect 502 2532 508 2533
rect 590 2537 596 2538
rect 590 2533 591 2537
rect 595 2533 596 2537
rect 590 2532 596 2533
rect 678 2537 684 2538
rect 678 2533 679 2537
rect 683 2533 684 2537
rect 678 2532 684 2533
rect 774 2537 780 2538
rect 774 2533 775 2537
rect 779 2533 780 2537
rect 774 2532 780 2533
rect 878 2537 884 2538
rect 878 2533 879 2537
rect 883 2533 884 2537
rect 878 2532 884 2533
rect 990 2537 996 2538
rect 990 2533 991 2537
rect 995 2533 996 2537
rect 990 2532 996 2533
rect 1102 2537 1108 2538
rect 1102 2533 1103 2537
rect 1107 2533 1108 2537
rect 1102 2532 1108 2533
rect 1222 2537 1228 2538
rect 1222 2533 1223 2537
rect 1227 2533 1228 2537
rect 1222 2532 1228 2533
rect 1350 2537 1356 2538
rect 1350 2533 1351 2537
rect 1355 2533 1356 2537
rect 1350 2532 1356 2533
rect 1478 2537 1484 2538
rect 1478 2533 1479 2537
rect 1483 2533 1484 2537
rect 1478 2532 1484 2533
rect 1606 2537 1612 2538
rect 1606 2533 1607 2537
rect 1611 2533 1612 2537
rect 1606 2532 1612 2533
rect 1766 2536 1772 2537
rect 1766 2532 1767 2536
rect 1771 2532 1772 2536
rect 1830 2533 1836 2534
rect 110 2531 116 2532
rect 1766 2531 1772 2532
rect 1806 2532 1812 2533
rect 1806 2528 1807 2532
rect 1811 2528 1812 2532
rect 1830 2529 1831 2533
rect 1835 2529 1836 2533
rect 1830 2528 1836 2529
rect 1918 2533 1924 2534
rect 1918 2529 1919 2533
rect 1923 2529 1924 2533
rect 1918 2528 1924 2529
rect 2006 2533 2012 2534
rect 2006 2529 2007 2533
rect 2011 2529 2012 2533
rect 2006 2528 2012 2529
rect 2110 2533 2116 2534
rect 2110 2529 2111 2533
rect 2115 2529 2116 2533
rect 2110 2528 2116 2529
rect 2222 2533 2228 2534
rect 2222 2529 2223 2533
rect 2227 2529 2228 2533
rect 2222 2528 2228 2529
rect 2342 2533 2348 2534
rect 2342 2529 2343 2533
rect 2347 2529 2348 2533
rect 2342 2528 2348 2529
rect 2486 2533 2492 2534
rect 2486 2529 2487 2533
rect 2491 2529 2492 2533
rect 2486 2528 2492 2529
rect 2646 2533 2652 2534
rect 2646 2529 2647 2533
rect 2651 2529 2652 2533
rect 2646 2528 2652 2529
rect 2814 2533 2820 2534
rect 2814 2529 2815 2533
rect 2819 2529 2820 2533
rect 2814 2528 2820 2529
rect 2998 2533 3004 2534
rect 2998 2529 2999 2533
rect 3003 2529 3004 2533
rect 2998 2528 3004 2529
rect 3190 2533 3196 2534
rect 3190 2529 3191 2533
rect 3195 2529 3196 2533
rect 3190 2528 3196 2529
rect 3366 2533 3372 2534
rect 3366 2529 3367 2533
rect 3371 2529 3372 2533
rect 3366 2528 3372 2529
rect 3462 2532 3468 2533
rect 3462 2528 3463 2532
rect 3467 2528 3468 2532
rect 1806 2527 1812 2528
rect 3462 2527 3468 2528
rect 551 2519 557 2520
rect 551 2515 552 2519
rect 556 2518 557 2519
rect 574 2519 580 2520
rect 556 2516 570 2518
rect 556 2515 557 2516
rect 551 2514 557 2515
rect 568 2510 570 2516
rect 574 2515 575 2519
rect 579 2518 580 2519
rect 639 2519 645 2520
rect 639 2518 640 2519
rect 579 2516 640 2518
rect 579 2515 580 2516
rect 574 2514 580 2515
rect 639 2515 640 2516
rect 644 2515 645 2519
rect 639 2514 645 2515
rect 662 2519 668 2520
rect 662 2515 663 2519
rect 667 2518 668 2519
rect 727 2519 733 2520
rect 727 2518 728 2519
rect 667 2516 728 2518
rect 667 2515 668 2516
rect 662 2514 668 2515
rect 727 2515 728 2516
rect 732 2515 733 2519
rect 727 2514 733 2515
rect 750 2519 756 2520
rect 750 2515 751 2519
rect 755 2518 756 2519
rect 823 2519 829 2520
rect 823 2518 824 2519
rect 755 2516 824 2518
rect 755 2515 756 2516
rect 750 2514 756 2515
rect 823 2515 824 2516
rect 828 2515 829 2519
rect 823 2514 829 2515
rect 846 2519 852 2520
rect 846 2515 847 2519
rect 851 2518 852 2519
rect 927 2519 933 2520
rect 927 2518 928 2519
rect 851 2516 928 2518
rect 851 2515 852 2516
rect 846 2514 852 2515
rect 927 2515 928 2516
rect 932 2515 933 2519
rect 927 2514 933 2515
rect 950 2519 956 2520
rect 950 2515 951 2519
rect 955 2518 956 2519
rect 1039 2519 1045 2520
rect 1039 2518 1040 2519
rect 955 2516 1040 2518
rect 955 2515 956 2516
rect 950 2514 956 2515
rect 1039 2515 1040 2516
rect 1044 2515 1045 2519
rect 1039 2514 1045 2515
rect 1062 2519 1068 2520
rect 1062 2515 1063 2519
rect 1067 2518 1068 2519
rect 1151 2519 1157 2520
rect 1151 2518 1152 2519
rect 1067 2516 1152 2518
rect 1067 2515 1068 2516
rect 1062 2514 1068 2515
rect 1151 2515 1152 2516
rect 1156 2515 1157 2519
rect 1151 2514 1157 2515
rect 1174 2519 1180 2520
rect 1174 2515 1175 2519
rect 1179 2518 1180 2519
rect 1271 2519 1277 2520
rect 1271 2518 1272 2519
rect 1179 2516 1272 2518
rect 1179 2515 1180 2516
rect 1174 2514 1180 2515
rect 1271 2515 1272 2516
rect 1276 2515 1277 2519
rect 1271 2514 1277 2515
rect 1399 2519 1405 2520
rect 1399 2515 1400 2519
rect 1404 2518 1405 2519
rect 1430 2519 1436 2520
rect 1430 2518 1431 2519
rect 1404 2516 1431 2518
rect 1404 2515 1405 2516
rect 1399 2514 1405 2515
rect 1430 2515 1431 2516
rect 1435 2515 1436 2519
rect 1430 2514 1436 2515
rect 1527 2519 1533 2520
rect 1527 2515 1528 2519
rect 1532 2518 1533 2519
rect 1558 2519 1564 2520
rect 1558 2518 1559 2519
rect 1532 2516 1559 2518
rect 1532 2515 1533 2516
rect 1527 2514 1533 2515
rect 1558 2515 1559 2516
rect 1563 2515 1564 2519
rect 1558 2514 1564 2515
rect 1655 2519 1661 2520
rect 1655 2515 1656 2519
rect 1660 2518 1661 2519
rect 1678 2519 1684 2520
rect 1678 2518 1679 2519
rect 1660 2516 1679 2518
rect 1660 2515 1661 2516
rect 1655 2514 1661 2515
rect 1678 2515 1679 2516
rect 1683 2515 1684 2519
rect 1678 2514 1684 2515
rect 1879 2515 1885 2516
rect 822 2511 828 2512
rect 822 2510 823 2511
rect 568 2508 823 2510
rect 822 2507 823 2508
rect 827 2507 828 2511
rect 1879 2511 1880 2515
rect 1884 2514 1885 2515
rect 1910 2515 1916 2516
rect 1910 2514 1911 2515
rect 1884 2512 1911 2514
rect 1884 2511 1885 2512
rect 1879 2510 1885 2511
rect 1910 2511 1911 2512
rect 1915 2511 1916 2515
rect 1910 2510 1916 2511
rect 1967 2515 1973 2516
rect 1967 2511 1968 2515
rect 1972 2514 1973 2515
rect 1999 2515 2005 2516
rect 1999 2514 2000 2515
rect 1972 2512 2000 2514
rect 1972 2511 1973 2512
rect 1967 2510 1973 2511
rect 1999 2511 2000 2512
rect 2004 2511 2005 2515
rect 1999 2510 2005 2511
rect 2055 2515 2061 2516
rect 2055 2511 2056 2515
rect 2060 2514 2061 2515
rect 2086 2515 2092 2516
rect 2086 2514 2087 2515
rect 2060 2512 2087 2514
rect 2060 2511 2061 2512
rect 2055 2510 2061 2511
rect 2086 2511 2087 2512
rect 2091 2511 2092 2515
rect 2086 2510 2092 2511
rect 2159 2515 2165 2516
rect 2159 2511 2160 2515
rect 2164 2514 2165 2515
rect 2190 2515 2196 2516
rect 2190 2514 2191 2515
rect 2164 2512 2191 2514
rect 2164 2511 2165 2512
rect 2159 2510 2165 2511
rect 2190 2511 2191 2512
rect 2195 2511 2196 2515
rect 2190 2510 2196 2511
rect 2206 2515 2212 2516
rect 2206 2511 2207 2515
rect 2211 2514 2212 2515
rect 2271 2515 2277 2516
rect 2271 2514 2272 2515
rect 2211 2512 2272 2514
rect 2211 2511 2212 2512
rect 2206 2510 2212 2511
rect 2271 2511 2272 2512
rect 2276 2511 2277 2515
rect 2271 2510 2277 2511
rect 2391 2515 2400 2516
rect 2391 2511 2392 2515
rect 2399 2511 2400 2515
rect 2391 2510 2400 2511
rect 2414 2515 2420 2516
rect 2414 2511 2415 2515
rect 2419 2514 2420 2515
rect 2535 2515 2541 2516
rect 2535 2514 2536 2515
rect 2419 2512 2536 2514
rect 2419 2511 2420 2512
rect 2414 2510 2420 2511
rect 2535 2511 2536 2512
rect 2540 2511 2541 2515
rect 2535 2510 2541 2511
rect 2558 2515 2564 2516
rect 2558 2511 2559 2515
rect 2563 2514 2564 2515
rect 2695 2515 2701 2516
rect 2695 2514 2696 2515
rect 2563 2512 2696 2514
rect 2563 2511 2564 2512
rect 2558 2510 2564 2511
rect 2695 2511 2696 2512
rect 2700 2511 2701 2515
rect 2695 2510 2701 2511
rect 2718 2515 2724 2516
rect 2718 2511 2719 2515
rect 2723 2514 2724 2515
rect 2863 2515 2869 2516
rect 2863 2514 2864 2515
rect 2723 2512 2864 2514
rect 2723 2511 2724 2512
rect 2718 2510 2724 2511
rect 2863 2511 2864 2512
rect 2868 2511 2869 2515
rect 2863 2510 2869 2511
rect 2886 2515 2892 2516
rect 2886 2511 2887 2515
rect 2891 2514 2892 2515
rect 3047 2515 3053 2516
rect 3047 2514 3048 2515
rect 2891 2512 3048 2514
rect 2891 2511 2892 2512
rect 2886 2510 2892 2511
rect 3047 2511 3048 2512
rect 3052 2511 3053 2515
rect 3047 2510 3053 2511
rect 3239 2515 3248 2516
rect 3239 2511 3240 2515
rect 3247 2511 3248 2515
rect 3239 2510 3248 2511
rect 3415 2515 3421 2516
rect 3415 2511 3416 2515
rect 3420 2514 3421 2515
rect 3438 2515 3444 2516
rect 3438 2514 3439 2515
rect 3420 2512 3439 2514
rect 3420 2511 3421 2512
rect 3415 2510 3421 2511
rect 3438 2511 3439 2512
rect 3443 2511 3444 2515
rect 3438 2510 3444 2511
rect 822 2506 828 2507
rect 1518 2507 1524 2508
rect 1518 2506 1519 2507
rect 1416 2504 1519 2506
rect 599 2499 605 2500
rect 599 2495 600 2499
rect 604 2498 605 2499
rect 630 2499 636 2500
rect 630 2498 631 2499
rect 604 2496 631 2498
rect 604 2495 605 2496
rect 599 2494 605 2495
rect 630 2495 631 2496
rect 635 2495 636 2499
rect 630 2494 636 2495
rect 783 2499 789 2500
rect 783 2495 784 2499
rect 788 2498 789 2499
rect 814 2499 820 2500
rect 814 2498 815 2499
rect 788 2496 815 2498
rect 788 2495 789 2496
rect 783 2494 789 2495
rect 814 2495 815 2496
rect 819 2495 820 2499
rect 814 2494 820 2495
rect 959 2499 965 2500
rect 959 2495 960 2499
rect 964 2498 965 2499
rect 1127 2499 1133 2500
rect 964 2496 994 2498
rect 964 2495 965 2496
rect 959 2494 965 2495
rect 990 2495 996 2496
rect 990 2491 991 2495
rect 995 2491 996 2495
rect 1127 2495 1128 2499
rect 1132 2498 1133 2499
rect 1215 2499 1221 2500
rect 1215 2498 1216 2499
rect 1132 2496 1216 2498
rect 1132 2495 1133 2496
rect 1127 2494 1133 2495
rect 1215 2495 1216 2496
rect 1220 2495 1221 2499
rect 1215 2494 1221 2495
rect 1287 2499 1293 2500
rect 1287 2495 1288 2499
rect 1292 2498 1293 2499
rect 1416 2498 1418 2504
rect 1518 2503 1519 2504
rect 1523 2503 1524 2507
rect 1518 2502 1524 2503
rect 1999 2503 2005 2504
rect 1292 2496 1418 2498
rect 1422 2499 1428 2500
rect 1292 2495 1293 2496
rect 1287 2494 1293 2495
rect 1422 2495 1423 2499
rect 1427 2498 1428 2499
rect 1447 2499 1453 2500
rect 1447 2498 1448 2499
rect 1427 2496 1448 2498
rect 1427 2495 1428 2496
rect 1422 2494 1428 2495
rect 1447 2495 1448 2496
rect 1452 2495 1453 2499
rect 1447 2494 1453 2495
rect 1470 2499 1476 2500
rect 1470 2495 1471 2499
rect 1475 2498 1476 2499
rect 1615 2499 1621 2500
rect 1615 2498 1616 2499
rect 1475 2496 1616 2498
rect 1475 2495 1476 2496
rect 1470 2494 1476 2495
rect 1615 2495 1616 2496
rect 1620 2495 1621 2499
rect 1999 2499 2000 2503
rect 2004 2502 2005 2503
rect 2014 2503 2020 2504
rect 2014 2502 2015 2503
rect 2004 2500 2015 2502
rect 2004 2499 2005 2500
rect 1999 2498 2005 2499
rect 2014 2499 2015 2500
rect 2019 2499 2020 2503
rect 2014 2498 2020 2499
rect 2022 2503 2028 2504
rect 2022 2499 2023 2503
rect 2027 2502 2028 2503
rect 2087 2503 2093 2504
rect 2087 2502 2088 2503
rect 2027 2500 2088 2502
rect 2027 2499 2028 2500
rect 2022 2498 2028 2499
rect 2087 2499 2088 2500
rect 2092 2499 2093 2503
rect 2087 2498 2093 2499
rect 2127 2503 2133 2504
rect 2127 2499 2128 2503
rect 2132 2502 2133 2503
rect 2183 2503 2189 2504
rect 2183 2502 2184 2503
rect 2132 2500 2184 2502
rect 2132 2499 2133 2500
rect 2127 2498 2133 2499
rect 2183 2499 2184 2500
rect 2188 2499 2189 2503
rect 2183 2498 2189 2499
rect 2287 2503 2293 2504
rect 2287 2499 2288 2503
rect 2292 2502 2293 2503
rect 2318 2503 2324 2504
rect 2318 2502 2319 2503
rect 2292 2500 2319 2502
rect 2292 2499 2293 2500
rect 2287 2498 2293 2499
rect 2318 2499 2319 2500
rect 2323 2499 2324 2503
rect 2318 2498 2324 2499
rect 2374 2503 2380 2504
rect 2374 2499 2375 2503
rect 2379 2502 2380 2503
rect 2415 2503 2421 2504
rect 2415 2502 2416 2503
rect 2379 2500 2416 2502
rect 2379 2499 2380 2500
rect 2374 2498 2380 2499
rect 2415 2499 2416 2500
rect 2420 2499 2421 2503
rect 2415 2498 2421 2499
rect 2575 2503 2584 2504
rect 2575 2499 2576 2503
rect 2583 2499 2584 2503
rect 2575 2498 2584 2499
rect 2598 2503 2604 2504
rect 2598 2499 2599 2503
rect 2603 2502 2604 2503
rect 2759 2503 2765 2504
rect 2759 2502 2760 2503
rect 2603 2500 2760 2502
rect 2603 2499 2604 2500
rect 2598 2498 2604 2499
rect 2759 2499 2760 2500
rect 2764 2499 2765 2503
rect 2759 2498 2765 2499
rect 2782 2503 2788 2504
rect 2782 2499 2783 2503
rect 2787 2502 2788 2503
rect 2967 2503 2973 2504
rect 2967 2502 2968 2503
rect 2787 2500 2968 2502
rect 2787 2499 2788 2500
rect 2782 2498 2788 2499
rect 2967 2499 2968 2500
rect 2972 2499 2973 2503
rect 2967 2498 2973 2499
rect 2990 2503 2996 2504
rect 2990 2499 2991 2503
rect 2995 2502 2996 2503
rect 3191 2503 3197 2504
rect 3191 2502 3192 2503
rect 2995 2500 3192 2502
rect 2995 2499 2996 2500
rect 2990 2498 2996 2499
rect 3191 2499 3192 2500
rect 3196 2499 3197 2503
rect 3191 2498 3197 2499
rect 3415 2503 3421 2504
rect 3415 2499 3416 2503
rect 3420 2502 3421 2503
rect 3430 2503 3436 2504
rect 3430 2502 3431 2503
rect 3420 2500 3431 2502
rect 3420 2499 3421 2500
rect 3415 2498 3421 2499
rect 3430 2499 3431 2500
rect 3435 2499 3436 2503
rect 3430 2498 3436 2499
rect 1615 2494 1621 2495
rect 990 2490 996 2491
rect 1806 2488 1812 2489
rect 3462 2488 3468 2489
rect 110 2484 116 2485
rect 1766 2484 1772 2485
rect 110 2480 111 2484
rect 115 2480 116 2484
rect 110 2479 116 2480
rect 550 2483 556 2484
rect 550 2479 551 2483
rect 555 2479 556 2483
rect 550 2478 556 2479
rect 734 2483 740 2484
rect 734 2479 735 2483
rect 739 2479 740 2483
rect 734 2478 740 2479
rect 910 2483 916 2484
rect 910 2479 911 2483
rect 915 2479 916 2483
rect 910 2478 916 2479
rect 1078 2483 1084 2484
rect 1078 2479 1079 2483
rect 1083 2479 1084 2483
rect 1078 2478 1084 2479
rect 1238 2483 1244 2484
rect 1238 2479 1239 2483
rect 1243 2479 1244 2483
rect 1238 2478 1244 2479
rect 1398 2483 1404 2484
rect 1398 2479 1399 2483
rect 1403 2479 1404 2483
rect 1398 2478 1404 2479
rect 1566 2483 1572 2484
rect 1566 2479 1567 2483
rect 1571 2479 1572 2483
rect 1766 2480 1767 2484
rect 1771 2480 1772 2484
rect 1806 2484 1807 2488
rect 1811 2484 1812 2488
rect 1806 2483 1812 2484
rect 1950 2487 1956 2488
rect 1950 2483 1951 2487
rect 1955 2483 1956 2487
rect 1950 2482 1956 2483
rect 2038 2487 2044 2488
rect 2038 2483 2039 2487
rect 2043 2483 2044 2487
rect 2038 2482 2044 2483
rect 2134 2487 2140 2488
rect 2134 2483 2135 2487
rect 2139 2483 2140 2487
rect 2134 2482 2140 2483
rect 2238 2487 2244 2488
rect 2238 2483 2239 2487
rect 2243 2483 2244 2487
rect 2238 2482 2244 2483
rect 2366 2487 2372 2488
rect 2366 2483 2367 2487
rect 2371 2483 2372 2487
rect 2366 2482 2372 2483
rect 2526 2487 2532 2488
rect 2526 2483 2527 2487
rect 2531 2483 2532 2487
rect 2526 2482 2532 2483
rect 2710 2487 2716 2488
rect 2710 2483 2711 2487
rect 2715 2483 2716 2487
rect 2710 2482 2716 2483
rect 2918 2487 2924 2488
rect 2918 2483 2919 2487
rect 2923 2483 2924 2487
rect 2918 2482 2924 2483
rect 3142 2487 3148 2488
rect 3142 2483 3143 2487
rect 3147 2483 3148 2487
rect 3142 2482 3148 2483
rect 3366 2487 3372 2488
rect 3366 2483 3367 2487
rect 3371 2483 3372 2487
rect 3462 2484 3463 2488
rect 3467 2484 3468 2488
rect 3462 2483 3468 2484
rect 3366 2482 3372 2483
rect 1766 2479 1772 2480
rect 2022 2479 2028 2480
rect 1566 2478 1572 2479
rect 630 2475 636 2476
rect 622 2471 628 2472
rect 110 2467 116 2468
rect 110 2463 111 2467
rect 115 2463 116 2467
rect 622 2467 623 2471
rect 627 2467 628 2471
rect 630 2471 631 2475
rect 635 2474 636 2475
rect 814 2475 820 2476
rect 635 2472 777 2474
rect 635 2471 636 2472
rect 630 2470 636 2471
rect 814 2471 815 2475
rect 819 2474 820 2475
rect 1215 2475 1221 2476
rect 819 2472 953 2474
rect 819 2471 820 2472
rect 814 2470 820 2471
rect 1150 2471 1156 2472
rect 622 2466 628 2467
rect 1150 2467 1151 2471
rect 1155 2467 1156 2471
rect 1215 2471 1216 2475
rect 1220 2474 1221 2475
rect 1470 2475 1476 2476
rect 1220 2472 1281 2474
rect 1220 2471 1221 2472
rect 1215 2470 1221 2471
rect 1470 2471 1471 2475
rect 1475 2471 1476 2475
rect 1470 2470 1476 2471
rect 1518 2475 1524 2476
rect 1518 2471 1519 2475
rect 1523 2474 1524 2475
rect 2022 2475 2023 2479
rect 2027 2475 2028 2479
rect 2127 2479 2133 2480
rect 2127 2478 2128 2479
rect 2113 2476 2128 2478
rect 2022 2474 2028 2475
rect 2127 2475 2128 2476
rect 2132 2475 2133 2479
rect 2127 2474 2133 2475
rect 2206 2479 2212 2480
rect 2206 2475 2207 2479
rect 2211 2475 2212 2479
rect 2206 2474 2212 2475
rect 2214 2479 2220 2480
rect 2214 2475 2215 2479
rect 2219 2478 2220 2479
rect 2318 2479 2324 2480
rect 2219 2476 2281 2478
rect 2219 2475 2220 2476
rect 2214 2474 2220 2475
rect 2318 2475 2319 2479
rect 2323 2478 2324 2479
rect 2598 2479 2604 2480
rect 2323 2476 2409 2478
rect 2323 2475 2324 2476
rect 2318 2474 2324 2475
rect 2598 2475 2599 2479
rect 2603 2475 2604 2479
rect 2598 2474 2604 2475
rect 2782 2479 2788 2480
rect 2782 2475 2783 2479
rect 2787 2475 2788 2479
rect 2782 2474 2788 2475
rect 2990 2479 2996 2480
rect 2990 2475 2991 2479
rect 2995 2475 2996 2479
rect 2990 2474 2996 2475
rect 3078 2479 3084 2480
rect 3078 2475 3079 2479
rect 3083 2478 3084 2479
rect 3242 2479 3248 2480
rect 3083 2476 3185 2478
rect 3083 2475 3084 2476
rect 3078 2474 3084 2475
rect 3242 2475 3243 2479
rect 3247 2478 3248 2479
rect 3247 2476 3409 2478
rect 3247 2475 3248 2476
rect 3242 2474 3248 2475
rect 1523 2472 1609 2474
rect 1523 2471 1524 2472
rect 1518 2470 1524 2471
rect 1806 2471 1812 2472
rect 1150 2466 1156 2467
rect 1766 2467 1772 2468
rect 110 2462 116 2463
rect 550 2464 556 2465
rect 550 2460 551 2464
rect 555 2460 556 2464
rect 550 2459 556 2460
rect 734 2464 740 2465
rect 734 2460 735 2464
rect 739 2460 740 2464
rect 734 2459 740 2460
rect 910 2464 916 2465
rect 910 2460 911 2464
rect 915 2460 916 2464
rect 910 2459 916 2460
rect 1078 2464 1084 2465
rect 1078 2460 1079 2464
rect 1083 2460 1084 2464
rect 1078 2459 1084 2460
rect 1238 2464 1244 2465
rect 1238 2460 1239 2464
rect 1243 2460 1244 2464
rect 1238 2459 1244 2460
rect 1398 2464 1404 2465
rect 1398 2460 1399 2464
rect 1403 2460 1404 2464
rect 1398 2459 1404 2460
rect 1566 2464 1572 2465
rect 1566 2460 1567 2464
rect 1571 2460 1572 2464
rect 1766 2463 1767 2467
rect 1771 2463 1772 2467
rect 1806 2467 1807 2471
rect 1811 2467 1812 2471
rect 3462 2471 3468 2472
rect 1806 2466 1812 2467
rect 1950 2468 1956 2469
rect 1950 2464 1951 2468
rect 1955 2464 1956 2468
rect 1950 2463 1956 2464
rect 2038 2468 2044 2469
rect 2038 2464 2039 2468
rect 2043 2464 2044 2468
rect 2038 2463 2044 2464
rect 2134 2468 2140 2469
rect 2134 2464 2135 2468
rect 2139 2464 2140 2468
rect 2134 2463 2140 2464
rect 2238 2468 2244 2469
rect 2238 2464 2239 2468
rect 2243 2464 2244 2468
rect 2238 2463 2244 2464
rect 2366 2468 2372 2469
rect 2366 2464 2367 2468
rect 2371 2464 2372 2468
rect 2366 2463 2372 2464
rect 2526 2468 2532 2469
rect 2526 2464 2527 2468
rect 2531 2464 2532 2468
rect 2526 2463 2532 2464
rect 2710 2468 2716 2469
rect 2710 2464 2711 2468
rect 2715 2464 2716 2468
rect 2710 2463 2716 2464
rect 2918 2468 2924 2469
rect 2918 2464 2919 2468
rect 2923 2464 2924 2468
rect 2918 2463 2924 2464
rect 3142 2468 3148 2469
rect 3142 2464 3143 2468
rect 3147 2464 3148 2468
rect 3142 2463 3148 2464
rect 3366 2468 3372 2469
rect 3366 2464 3367 2468
rect 3371 2464 3372 2468
rect 3462 2467 3463 2471
rect 3467 2467 3468 2471
rect 3462 2466 3468 2467
rect 3366 2463 3372 2464
rect 1766 2462 1772 2463
rect 1566 2459 1572 2460
rect 2618 2431 2624 2432
rect 2618 2427 2619 2431
rect 2623 2430 2624 2431
rect 3078 2431 3084 2432
rect 3078 2430 3079 2431
rect 2623 2428 3079 2430
rect 2623 2427 2624 2428
rect 2618 2426 2624 2427
rect 3078 2427 3079 2428
rect 3083 2427 3084 2431
rect 3078 2426 3084 2427
rect 2262 2423 2268 2424
rect 414 2420 420 2421
rect 110 2417 116 2418
rect 110 2413 111 2417
rect 115 2413 116 2417
rect 414 2416 415 2420
rect 419 2416 420 2420
rect 414 2415 420 2416
rect 502 2420 508 2421
rect 502 2416 503 2420
rect 507 2416 508 2420
rect 502 2415 508 2416
rect 598 2420 604 2421
rect 598 2416 599 2420
rect 603 2416 604 2420
rect 598 2415 604 2416
rect 702 2420 708 2421
rect 702 2416 703 2420
rect 707 2416 708 2420
rect 702 2415 708 2416
rect 806 2420 812 2421
rect 806 2416 807 2420
rect 811 2416 812 2420
rect 806 2415 812 2416
rect 918 2420 924 2421
rect 918 2416 919 2420
rect 923 2416 924 2420
rect 918 2415 924 2416
rect 1038 2420 1044 2421
rect 1038 2416 1039 2420
rect 1043 2416 1044 2420
rect 1038 2415 1044 2416
rect 1166 2420 1172 2421
rect 1166 2416 1167 2420
rect 1171 2416 1172 2420
rect 1166 2415 1172 2416
rect 1294 2420 1300 2421
rect 1294 2416 1295 2420
rect 1299 2416 1300 2420
rect 1294 2415 1300 2416
rect 1422 2420 1428 2421
rect 1422 2416 1423 2420
rect 1427 2416 1428 2420
rect 2262 2419 2263 2423
rect 2267 2422 2268 2423
rect 2750 2423 2756 2424
rect 2267 2420 2386 2422
rect 2267 2419 2268 2420
rect 2262 2418 2268 2419
rect 1422 2415 1428 2416
rect 1766 2417 1772 2418
rect 110 2412 116 2413
rect 1766 2413 1767 2417
rect 1771 2413 1772 2417
rect 2214 2416 2220 2417
rect 1766 2412 1772 2413
rect 1806 2413 1812 2414
rect 486 2411 492 2412
rect 486 2407 487 2411
rect 491 2407 492 2411
rect 486 2406 492 2407
rect 574 2411 580 2412
rect 574 2407 575 2411
rect 579 2407 580 2411
rect 574 2406 580 2407
rect 582 2411 588 2412
rect 582 2407 583 2411
rect 587 2410 588 2411
rect 774 2411 780 2412
rect 587 2408 641 2410
rect 587 2407 588 2408
rect 582 2406 588 2407
rect 774 2407 775 2411
rect 779 2407 780 2411
rect 774 2406 780 2407
rect 878 2411 884 2412
rect 878 2407 879 2411
rect 883 2407 884 2411
rect 878 2406 884 2407
rect 990 2411 996 2412
rect 990 2407 991 2411
rect 995 2407 996 2411
rect 990 2406 996 2407
rect 998 2411 1004 2412
rect 998 2407 999 2411
rect 1003 2410 1004 2411
rect 1238 2411 1244 2412
rect 1003 2408 1081 2410
rect 1003 2407 1004 2408
rect 998 2406 1004 2407
rect 1238 2407 1239 2411
rect 1243 2407 1244 2411
rect 1238 2406 1244 2407
rect 1366 2411 1372 2412
rect 1366 2407 1367 2411
rect 1371 2407 1372 2411
rect 1366 2406 1372 2407
rect 1386 2411 1392 2412
rect 1386 2407 1387 2411
rect 1391 2410 1392 2411
rect 1391 2408 1465 2410
rect 1806 2409 1807 2413
rect 1811 2409 1812 2413
rect 2214 2412 2215 2416
rect 2219 2412 2220 2416
rect 2214 2411 2220 2412
rect 2302 2416 2308 2417
rect 2302 2412 2303 2416
rect 2307 2412 2308 2416
rect 2302 2411 2308 2412
rect 1806 2408 1812 2409
rect 1391 2407 1392 2408
rect 1386 2406 1392 2407
rect 2286 2407 2292 2408
rect 2286 2403 2287 2407
rect 2291 2403 2292 2407
rect 2286 2402 2292 2403
rect 2374 2407 2380 2408
rect 2374 2403 2375 2407
rect 2379 2403 2380 2407
rect 2384 2406 2386 2420
rect 2750 2419 2751 2423
rect 2755 2422 2756 2423
rect 2755 2420 2922 2422
rect 2755 2419 2756 2420
rect 2750 2418 2756 2419
rect 2390 2416 2396 2417
rect 2390 2412 2391 2416
rect 2395 2412 2396 2416
rect 2390 2411 2396 2412
rect 2478 2416 2484 2417
rect 2478 2412 2479 2416
rect 2483 2412 2484 2416
rect 2478 2411 2484 2412
rect 2566 2416 2572 2417
rect 2566 2412 2567 2416
rect 2571 2412 2572 2416
rect 2566 2411 2572 2412
rect 2654 2416 2660 2417
rect 2654 2412 2655 2416
rect 2659 2412 2660 2416
rect 2654 2411 2660 2412
rect 2742 2416 2748 2417
rect 2742 2412 2743 2416
rect 2747 2412 2748 2416
rect 2742 2411 2748 2412
rect 2838 2416 2844 2417
rect 2838 2412 2839 2416
rect 2843 2412 2844 2416
rect 2838 2411 2844 2412
rect 2471 2407 2477 2408
rect 2384 2404 2433 2406
rect 2374 2402 2380 2403
rect 2471 2403 2472 2407
rect 2476 2406 2477 2407
rect 2638 2407 2644 2408
rect 2476 2404 2521 2406
rect 2476 2403 2477 2404
rect 2471 2402 2477 2403
rect 2638 2403 2639 2407
rect 2643 2403 2644 2407
rect 2638 2402 2644 2403
rect 2726 2407 2732 2408
rect 2726 2403 2727 2407
rect 2731 2403 2732 2407
rect 2726 2402 2732 2403
rect 2814 2407 2820 2408
rect 2814 2403 2815 2407
rect 2819 2403 2820 2407
rect 2920 2406 2922 2420
rect 2934 2416 2940 2417
rect 2934 2412 2935 2416
rect 2939 2412 2940 2416
rect 2934 2411 2940 2412
rect 3462 2413 3468 2414
rect 3462 2409 3463 2413
rect 3467 2409 3468 2413
rect 3462 2408 3468 2409
rect 2920 2404 2977 2406
rect 2814 2402 2820 2403
rect 414 2401 420 2402
rect 110 2400 116 2401
rect 110 2396 111 2400
rect 115 2396 116 2400
rect 414 2397 415 2401
rect 419 2397 420 2401
rect 414 2396 420 2397
rect 502 2401 508 2402
rect 502 2397 503 2401
rect 507 2397 508 2401
rect 502 2396 508 2397
rect 598 2401 604 2402
rect 598 2397 599 2401
rect 603 2397 604 2401
rect 598 2396 604 2397
rect 702 2401 708 2402
rect 702 2397 703 2401
rect 707 2397 708 2401
rect 702 2396 708 2397
rect 806 2401 812 2402
rect 806 2397 807 2401
rect 811 2397 812 2401
rect 806 2396 812 2397
rect 918 2401 924 2402
rect 918 2397 919 2401
rect 923 2397 924 2401
rect 918 2396 924 2397
rect 1038 2401 1044 2402
rect 1038 2397 1039 2401
rect 1043 2397 1044 2401
rect 1038 2396 1044 2397
rect 1166 2401 1172 2402
rect 1166 2397 1167 2401
rect 1171 2397 1172 2401
rect 1166 2396 1172 2397
rect 1294 2401 1300 2402
rect 1294 2397 1295 2401
rect 1299 2397 1300 2401
rect 1294 2396 1300 2397
rect 1422 2401 1428 2402
rect 1422 2397 1423 2401
rect 1427 2397 1428 2401
rect 1422 2396 1428 2397
rect 1766 2400 1772 2401
rect 1766 2396 1767 2400
rect 1771 2396 1772 2400
rect 2911 2399 2917 2400
rect 2214 2397 2220 2398
rect 110 2395 116 2396
rect 1766 2395 1772 2396
rect 1806 2396 1812 2397
rect 1806 2392 1807 2396
rect 1811 2392 1812 2396
rect 2214 2393 2215 2397
rect 2219 2393 2220 2397
rect 2214 2392 2220 2393
rect 2302 2397 2308 2398
rect 2302 2393 2303 2397
rect 2307 2393 2308 2397
rect 2302 2392 2308 2393
rect 2390 2397 2396 2398
rect 2390 2393 2391 2397
rect 2395 2393 2396 2397
rect 2390 2392 2396 2393
rect 2478 2397 2484 2398
rect 2478 2393 2479 2397
rect 2483 2393 2484 2397
rect 2478 2392 2484 2393
rect 2566 2397 2572 2398
rect 2566 2393 2567 2397
rect 2571 2393 2572 2397
rect 2566 2392 2572 2393
rect 2654 2397 2660 2398
rect 2654 2393 2655 2397
rect 2659 2393 2660 2397
rect 2654 2392 2660 2393
rect 2742 2397 2748 2398
rect 2742 2393 2743 2397
rect 2747 2393 2748 2397
rect 2742 2392 2748 2393
rect 2838 2397 2844 2398
rect 2838 2393 2839 2397
rect 2843 2393 2844 2397
rect 2911 2395 2912 2399
rect 2916 2398 2917 2399
rect 2926 2399 2932 2400
rect 2926 2398 2927 2399
rect 2916 2396 2927 2398
rect 2916 2395 2917 2396
rect 2911 2394 2917 2395
rect 2926 2395 2927 2396
rect 2931 2395 2932 2399
rect 2926 2394 2932 2395
rect 2934 2397 2940 2398
rect 2838 2392 2844 2393
rect 2934 2393 2935 2397
rect 2939 2393 2940 2397
rect 2934 2392 2940 2393
rect 3462 2396 3468 2397
rect 3462 2392 3463 2396
rect 3467 2392 3468 2396
rect 1806 2391 1812 2392
rect 3462 2391 3468 2392
rect 463 2383 469 2384
rect 463 2379 464 2383
rect 468 2382 469 2383
rect 486 2383 492 2384
rect 468 2380 482 2382
rect 468 2379 469 2380
rect 463 2378 469 2379
rect 480 2374 482 2380
rect 486 2379 487 2383
rect 491 2382 492 2383
rect 551 2383 557 2384
rect 551 2382 552 2383
rect 491 2380 552 2382
rect 491 2379 492 2380
rect 486 2378 492 2379
rect 551 2379 552 2380
rect 556 2379 557 2383
rect 551 2378 557 2379
rect 622 2383 628 2384
rect 622 2379 623 2383
rect 627 2382 628 2383
rect 647 2383 653 2384
rect 647 2382 648 2383
rect 627 2380 648 2382
rect 627 2379 628 2380
rect 622 2378 628 2379
rect 647 2379 648 2380
rect 652 2379 653 2383
rect 647 2378 653 2379
rect 751 2383 757 2384
rect 751 2379 752 2383
rect 756 2382 757 2383
rect 774 2383 780 2384
rect 756 2380 770 2382
rect 756 2379 757 2380
rect 751 2378 757 2379
rect 582 2375 588 2376
rect 582 2374 583 2375
rect 480 2372 583 2374
rect 582 2371 583 2372
rect 587 2371 588 2375
rect 768 2374 770 2380
rect 774 2379 775 2383
rect 779 2382 780 2383
rect 855 2383 861 2384
rect 855 2382 856 2383
rect 779 2380 856 2382
rect 779 2379 780 2380
rect 774 2378 780 2379
rect 855 2379 856 2380
rect 860 2379 861 2383
rect 855 2378 861 2379
rect 878 2383 884 2384
rect 878 2379 879 2383
rect 883 2382 884 2383
rect 967 2383 973 2384
rect 967 2382 968 2383
rect 883 2380 968 2382
rect 883 2379 884 2380
rect 878 2378 884 2379
rect 967 2379 968 2380
rect 972 2379 973 2383
rect 967 2378 973 2379
rect 1062 2383 1068 2384
rect 1062 2379 1063 2383
rect 1067 2382 1068 2383
rect 1087 2383 1093 2384
rect 1087 2382 1088 2383
rect 1067 2380 1088 2382
rect 1067 2379 1068 2380
rect 1062 2378 1068 2379
rect 1087 2379 1088 2380
rect 1092 2379 1093 2383
rect 1087 2378 1093 2379
rect 1150 2383 1156 2384
rect 1150 2379 1151 2383
rect 1155 2382 1156 2383
rect 1215 2383 1221 2384
rect 1215 2382 1216 2383
rect 1155 2380 1216 2382
rect 1155 2379 1156 2380
rect 1150 2378 1156 2379
rect 1215 2379 1216 2380
rect 1220 2379 1221 2383
rect 1215 2378 1221 2379
rect 1238 2383 1244 2384
rect 1238 2379 1239 2383
rect 1243 2382 1244 2383
rect 1343 2383 1349 2384
rect 1343 2382 1344 2383
rect 1243 2380 1344 2382
rect 1243 2379 1244 2380
rect 1238 2378 1244 2379
rect 1343 2379 1344 2380
rect 1348 2379 1349 2383
rect 1343 2378 1349 2379
rect 1366 2383 1372 2384
rect 1366 2379 1367 2383
rect 1371 2382 1372 2383
rect 1471 2383 1477 2384
rect 1471 2382 1472 2383
rect 1371 2380 1472 2382
rect 1371 2379 1372 2380
rect 1366 2378 1372 2379
rect 1471 2379 1472 2380
rect 1476 2379 1477 2383
rect 1471 2378 1477 2379
rect 2262 2383 2268 2384
rect 2262 2379 2263 2383
rect 2267 2382 2268 2383
rect 2267 2381 2269 2382
rect 2262 2378 2264 2379
rect 2263 2377 2264 2378
rect 2268 2377 2269 2381
rect 2263 2376 2269 2377
rect 2286 2379 2292 2380
rect 998 2375 1004 2376
rect 998 2374 999 2375
rect 768 2372 999 2374
rect 582 2370 588 2371
rect 998 2371 999 2372
rect 1003 2371 1004 2375
rect 2286 2375 2287 2379
rect 2291 2378 2292 2379
rect 2351 2379 2357 2380
rect 2351 2378 2352 2379
rect 2291 2376 2352 2378
rect 2291 2375 2292 2376
rect 2286 2374 2292 2375
rect 2351 2375 2352 2376
rect 2356 2375 2357 2379
rect 2351 2374 2357 2375
rect 2439 2379 2445 2380
rect 2439 2375 2440 2379
rect 2444 2378 2445 2379
rect 2471 2379 2477 2380
rect 2471 2378 2472 2379
rect 2444 2376 2472 2378
rect 2444 2375 2445 2376
rect 2439 2374 2445 2375
rect 2471 2375 2472 2376
rect 2476 2375 2477 2379
rect 2471 2374 2477 2375
rect 2527 2379 2533 2380
rect 2527 2375 2528 2379
rect 2532 2378 2533 2379
rect 2550 2379 2556 2380
rect 2550 2378 2551 2379
rect 2532 2376 2551 2378
rect 2532 2375 2533 2376
rect 2527 2374 2533 2375
rect 2550 2375 2551 2376
rect 2555 2375 2556 2379
rect 2550 2374 2556 2375
rect 2615 2379 2624 2380
rect 2615 2375 2616 2379
rect 2623 2375 2624 2379
rect 2615 2374 2624 2375
rect 2638 2379 2644 2380
rect 2638 2375 2639 2379
rect 2643 2378 2644 2379
rect 2703 2379 2709 2380
rect 2703 2378 2704 2379
rect 2643 2376 2704 2378
rect 2643 2375 2644 2376
rect 2638 2374 2644 2375
rect 2703 2375 2704 2376
rect 2708 2375 2709 2379
rect 2703 2374 2709 2375
rect 2726 2379 2732 2380
rect 2726 2375 2727 2379
rect 2731 2378 2732 2379
rect 2791 2379 2797 2380
rect 2791 2378 2792 2379
rect 2731 2376 2792 2378
rect 2731 2375 2732 2376
rect 2726 2374 2732 2375
rect 2791 2375 2792 2376
rect 2796 2375 2797 2379
rect 2791 2374 2797 2375
rect 2814 2379 2820 2380
rect 2814 2375 2815 2379
rect 2819 2378 2820 2379
rect 2887 2379 2893 2380
rect 2887 2378 2888 2379
rect 2819 2376 2888 2378
rect 2819 2375 2820 2376
rect 2814 2374 2820 2375
rect 2887 2375 2888 2376
rect 2892 2375 2893 2379
rect 2887 2374 2893 2375
rect 2926 2379 2932 2380
rect 2926 2375 2927 2379
rect 2931 2378 2932 2379
rect 2983 2379 2989 2380
rect 2983 2378 2984 2379
rect 2931 2376 2984 2378
rect 2931 2375 2932 2376
rect 2926 2374 2932 2375
rect 2983 2375 2984 2376
rect 2988 2375 2989 2379
rect 2983 2374 2989 2375
rect 998 2370 1004 2371
rect 367 2367 373 2368
rect 367 2363 368 2367
rect 372 2366 373 2367
rect 398 2367 404 2368
rect 398 2366 399 2367
rect 372 2364 399 2366
rect 372 2363 373 2364
rect 367 2362 373 2363
rect 398 2363 399 2364
rect 403 2363 404 2367
rect 398 2362 404 2363
rect 479 2367 485 2368
rect 479 2363 480 2367
rect 484 2366 485 2367
rect 550 2367 556 2368
rect 550 2366 551 2367
rect 484 2364 551 2366
rect 484 2363 485 2364
rect 479 2362 485 2363
rect 550 2363 551 2364
rect 555 2363 556 2367
rect 550 2362 556 2363
rect 574 2367 580 2368
rect 574 2363 575 2367
rect 579 2366 580 2367
rect 591 2367 597 2368
rect 591 2366 592 2367
rect 579 2364 592 2366
rect 579 2363 580 2364
rect 574 2362 580 2363
rect 591 2363 592 2364
rect 596 2363 597 2367
rect 591 2362 597 2363
rect 614 2367 620 2368
rect 614 2363 615 2367
rect 619 2366 620 2367
rect 703 2367 709 2368
rect 703 2366 704 2367
rect 619 2364 704 2366
rect 619 2363 620 2364
rect 614 2362 620 2363
rect 703 2363 704 2364
rect 708 2363 709 2367
rect 703 2362 709 2363
rect 815 2367 821 2368
rect 815 2363 816 2367
rect 820 2366 821 2367
rect 846 2367 852 2368
rect 846 2366 847 2367
rect 820 2364 847 2366
rect 820 2363 821 2364
rect 815 2362 821 2363
rect 846 2363 847 2364
rect 851 2363 852 2367
rect 846 2362 852 2363
rect 866 2367 872 2368
rect 866 2363 867 2367
rect 871 2366 872 2367
rect 927 2367 933 2368
rect 927 2366 928 2367
rect 871 2364 928 2366
rect 871 2363 872 2364
rect 866 2362 872 2363
rect 927 2363 928 2364
rect 932 2363 933 2367
rect 927 2362 933 2363
rect 950 2367 956 2368
rect 950 2363 951 2367
rect 955 2366 956 2367
rect 1039 2367 1045 2368
rect 1039 2366 1040 2367
rect 955 2364 1040 2366
rect 955 2363 956 2364
rect 950 2362 956 2363
rect 1039 2363 1040 2364
rect 1044 2363 1045 2367
rect 1039 2362 1045 2363
rect 1151 2367 1157 2368
rect 1151 2363 1152 2367
rect 1156 2366 1157 2367
rect 1206 2367 1212 2368
rect 1206 2366 1207 2367
rect 1156 2364 1207 2366
rect 1156 2363 1157 2364
rect 1151 2362 1157 2363
rect 1206 2363 1207 2364
rect 1211 2363 1212 2367
rect 1206 2362 1212 2363
rect 1263 2367 1269 2368
rect 1263 2363 1264 2367
rect 1268 2366 1269 2367
rect 1295 2367 1301 2368
rect 1295 2366 1296 2367
rect 1268 2364 1296 2366
rect 1268 2363 1269 2364
rect 1263 2362 1269 2363
rect 1295 2363 1296 2364
rect 1300 2363 1301 2367
rect 1295 2362 1301 2363
rect 1383 2367 1392 2368
rect 1383 2363 1384 2367
rect 1391 2363 1392 2367
rect 1383 2362 1392 2363
rect 2215 2367 2221 2368
rect 2215 2363 2216 2367
rect 2220 2366 2221 2367
rect 2230 2367 2236 2368
rect 2230 2366 2231 2367
rect 2220 2364 2231 2366
rect 2220 2363 2221 2364
rect 2215 2362 2221 2363
rect 2230 2363 2231 2364
rect 2235 2363 2236 2367
rect 2230 2362 2236 2363
rect 2238 2367 2244 2368
rect 2238 2363 2239 2367
rect 2243 2366 2244 2367
rect 2311 2367 2317 2368
rect 2311 2366 2312 2367
rect 2243 2364 2312 2366
rect 2243 2363 2244 2364
rect 2238 2362 2244 2363
rect 2311 2363 2312 2364
rect 2316 2363 2317 2367
rect 2311 2362 2317 2363
rect 2334 2367 2340 2368
rect 2334 2363 2335 2367
rect 2339 2366 2340 2367
rect 2415 2367 2421 2368
rect 2415 2366 2416 2367
rect 2339 2364 2416 2366
rect 2339 2363 2340 2364
rect 2334 2362 2340 2363
rect 2415 2363 2416 2364
rect 2420 2363 2421 2367
rect 2415 2362 2421 2363
rect 2438 2367 2444 2368
rect 2438 2363 2439 2367
rect 2443 2366 2444 2367
rect 2519 2367 2525 2368
rect 2519 2366 2520 2367
rect 2443 2364 2520 2366
rect 2443 2363 2444 2364
rect 2438 2362 2444 2363
rect 2519 2363 2520 2364
rect 2524 2363 2525 2367
rect 2519 2362 2525 2363
rect 2542 2367 2548 2368
rect 2542 2363 2543 2367
rect 2547 2366 2548 2367
rect 2623 2367 2629 2368
rect 2623 2366 2624 2367
rect 2547 2364 2624 2366
rect 2547 2363 2548 2364
rect 2542 2362 2548 2363
rect 2623 2363 2624 2364
rect 2628 2363 2629 2367
rect 2623 2362 2629 2363
rect 2735 2367 2741 2368
rect 2735 2363 2736 2367
rect 2740 2366 2741 2367
rect 2750 2367 2756 2368
rect 2750 2366 2751 2367
rect 2740 2364 2751 2366
rect 2740 2363 2741 2364
rect 2735 2362 2741 2363
rect 2750 2363 2751 2364
rect 2755 2363 2756 2367
rect 2750 2362 2756 2363
rect 2758 2367 2764 2368
rect 2758 2363 2759 2367
rect 2763 2366 2764 2367
rect 2847 2367 2853 2368
rect 2847 2366 2848 2367
rect 2763 2364 2848 2366
rect 2763 2363 2764 2364
rect 2758 2362 2764 2363
rect 2847 2363 2848 2364
rect 2852 2363 2853 2367
rect 2847 2362 2853 2363
rect 2870 2367 2876 2368
rect 2870 2363 2871 2367
rect 2875 2366 2876 2367
rect 2959 2367 2965 2368
rect 2959 2366 2960 2367
rect 2875 2364 2960 2366
rect 2875 2363 2876 2364
rect 2870 2362 2876 2363
rect 2959 2363 2960 2364
rect 2964 2363 2965 2367
rect 2959 2362 2965 2363
rect 2982 2367 2988 2368
rect 2982 2363 2983 2367
rect 2987 2366 2988 2367
rect 3071 2367 3077 2368
rect 3071 2366 3072 2367
rect 2987 2364 3072 2366
rect 2987 2363 2988 2364
rect 2982 2362 2988 2363
rect 3071 2363 3072 2364
rect 3076 2363 3077 2367
rect 3071 2362 3077 2363
rect 110 2352 116 2353
rect 1766 2352 1772 2353
rect 110 2348 111 2352
rect 115 2348 116 2352
rect 110 2347 116 2348
rect 318 2351 324 2352
rect 318 2347 319 2351
rect 323 2347 324 2351
rect 318 2346 324 2347
rect 430 2351 436 2352
rect 430 2347 431 2351
rect 435 2347 436 2351
rect 430 2346 436 2347
rect 542 2351 548 2352
rect 542 2347 543 2351
rect 547 2347 548 2351
rect 542 2346 548 2347
rect 654 2351 660 2352
rect 654 2347 655 2351
rect 659 2347 660 2351
rect 654 2346 660 2347
rect 766 2351 772 2352
rect 766 2347 767 2351
rect 771 2347 772 2351
rect 766 2346 772 2347
rect 878 2351 884 2352
rect 878 2347 879 2351
rect 883 2347 884 2351
rect 878 2346 884 2347
rect 990 2351 996 2352
rect 990 2347 991 2351
rect 995 2347 996 2351
rect 990 2346 996 2347
rect 1102 2351 1108 2352
rect 1102 2347 1103 2351
rect 1107 2347 1108 2351
rect 1102 2346 1108 2347
rect 1214 2351 1220 2352
rect 1214 2347 1215 2351
rect 1219 2347 1220 2351
rect 1214 2346 1220 2347
rect 1334 2351 1340 2352
rect 1334 2347 1335 2351
rect 1339 2347 1340 2351
rect 1766 2348 1767 2352
rect 1771 2348 1772 2352
rect 1766 2347 1772 2348
rect 1806 2352 1812 2353
rect 3462 2352 3468 2353
rect 1806 2348 1807 2352
rect 1811 2348 1812 2352
rect 1806 2347 1812 2348
rect 2166 2351 2172 2352
rect 2166 2347 2167 2351
rect 2171 2347 2172 2351
rect 1334 2346 1340 2347
rect 2166 2346 2172 2347
rect 2262 2351 2268 2352
rect 2262 2347 2263 2351
rect 2267 2347 2268 2351
rect 2262 2346 2268 2347
rect 2366 2351 2372 2352
rect 2366 2347 2367 2351
rect 2371 2347 2372 2351
rect 2366 2346 2372 2347
rect 2470 2351 2476 2352
rect 2470 2347 2471 2351
rect 2475 2347 2476 2351
rect 2470 2346 2476 2347
rect 2574 2351 2580 2352
rect 2574 2347 2575 2351
rect 2579 2347 2580 2351
rect 2574 2346 2580 2347
rect 2686 2351 2692 2352
rect 2686 2347 2687 2351
rect 2691 2347 2692 2351
rect 2686 2346 2692 2347
rect 2798 2351 2804 2352
rect 2798 2347 2799 2351
rect 2803 2347 2804 2351
rect 2798 2346 2804 2347
rect 2910 2351 2916 2352
rect 2910 2347 2911 2351
rect 2915 2347 2916 2351
rect 2910 2346 2916 2347
rect 3022 2351 3028 2352
rect 3022 2347 3023 2351
rect 3027 2347 3028 2351
rect 3462 2348 3463 2352
rect 3467 2348 3468 2352
rect 3462 2347 3468 2348
rect 3022 2346 3028 2347
rect 398 2343 404 2344
rect 398 2339 399 2343
rect 403 2342 404 2343
rect 614 2343 620 2344
rect 403 2340 473 2342
rect 403 2339 404 2340
rect 398 2338 404 2339
rect 614 2339 615 2343
rect 619 2339 620 2343
rect 866 2343 872 2344
rect 866 2342 867 2343
rect 614 2338 620 2339
rect 624 2340 697 2342
rect 841 2340 867 2342
rect 110 2335 116 2336
rect 110 2331 111 2335
rect 115 2331 116 2335
rect 392 2334 394 2337
rect 398 2335 404 2336
rect 398 2334 399 2335
rect 110 2330 116 2331
rect 318 2332 324 2333
rect 392 2332 399 2334
rect 318 2328 319 2332
rect 323 2328 324 2332
rect 398 2331 399 2332
rect 403 2331 404 2335
rect 398 2330 404 2331
rect 430 2332 436 2333
rect 318 2327 324 2328
rect 430 2328 431 2332
rect 435 2328 436 2332
rect 430 2327 436 2328
rect 542 2332 548 2333
rect 542 2328 543 2332
rect 547 2328 548 2332
rect 542 2327 548 2328
rect 550 2327 556 2328
rect 550 2323 551 2327
rect 555 2326 556 2327
rect 624 2326 626 2340
rect 866 2339 867 2340
rect 871 2339 872 2343
rect 866 2338 872 2339
rect 950 2343 956 2344
rect 950 2339 951 2343
rect 955 2339 956 2343
rect 950 2338 956 2339
rect 1062 2343 1068 2344
rect 1062 2339 1063 2343
rect 1067 2339 1068 2343
rect 1062 2338 1068 2339
rect 1070 2343 1076 2344
rect 1070 2339 1071 2343
rect 1075 2342 1076 2343
rect 1206 2343 1212 2344
rect 1075 2340 1145 2342
rect 1075 2339 1076 2340
rect 1070 2338 1076 2339
rect 1206 2339 1207 2343
rect 1211 2342 1212 2343
rect 1295 2343 1301 2344
rect 1211 2340 1257 2342
rect 1211 2339 1212 2340
rect 1206 2338 1212 2339
rect 1295 2339 1296 2343
rect 1300 2342 1301 2343
rect 2238 2343 2244 2344
rect 1300 2340 1377 2342
rect 1300 2339 1301 2340
rect 1295 2338 1301 2339
rect 2238 2339 2239 2343
rect 2243 2339 2244 2343
rect 2238 2338 2244 2339
rect 2334 2343 2340 2344
rect 2334 2339 2335 2343
rect 2339 2339 2340 2343
rect 2334 2338 2340 2339
rect 2438 2343 2444 2344
rect 2438 2339 2439 2343
rect 2443 2339 2444 2343
rect 2438 2338 2444 2339
rect 2542 2343 2548 2344
rect 2542 2339 2543 2343
rect 2547 2339 2548 2343
rect 2542 2338 2548 2339
rect 2550 2343 2556 2344
rect 2550 2339 2551 2343
rect 2555 2342 2556 2343
rect 2758 2343 2764 2344
rect 2555 2340 2617 2342
rect 2555 2339 2556 2340
rect 2550 2338 2556 2339
rect 2758 2339 2759 2343
rect 2763 2339 2764 2343
rect 2758 2338 2764 2339
rect 2870 2343 2876 2344
rect 2870 2339 2871 2343
rect 2875 2339 2876 2343
rect 2870 2338 2876 2339
rect 2982 2343 2988 2344
rect 2982 2339 2983 2343
rect 2987 2339 2988 2343
rect 2982 2338 2988 2339
rect 2990 2343 2996 2344
rect 2990 2339 2991 2343
rect 2995 2342 2996 2343
rect 2995 2340 3065 2342
rect 2995 2339 2996 2340
rect 2990 2338 2996 2339
rect 1766 2335 1772 2336
rect 654 2332 660 2333
rect 654 2328 655 2332
rect 659 2328 660 2332
rect 654 2327 660 2328
rect 766 2332 772 2333
rect 766 2328 767 2332
rect 771 2328 772 2332
rect 766 2327 772 2328
rect 878 2332 884 2333
rect 878 2328 879 2332
rect 883 2328 884 2332
rect 878 2327 884 2328
rect 990 2332 996 2333
rect 990 2328 991 2332
rect 995 2328 996 2332
rect 990 2327 996 2328
rect 1102 2332 1108 2333
rect 1102 2328 1103 2332
rect 1107 2328 1108 2332
rect 1102 2327 1108 2328
rect 1214 2332 1220 2333
rect 1214 2328 1215 2332
rect 1219 2328 1220 2332
rect 1214 2327 1220 2328
rect 1334 2332 1340 2333
rect 1334 2328 1335 2332
rect 1339 2328 1340 2332
rect 1766 2331 1767 2335
rect 1771 2331 1772 2335
rect 1766 2330 1772 2331
rect 1806 2335 1812 2336
rect 1806 2331 1807 2335
rect 1811 2331 1812 2335
rect 3462 2335 3468 2336
rect 1806 2330 1812 2331
rect 2166 2332 2172 2333
rect 1334 2327 1340 2328
rect 2166 2328 2167 2332
rect 2171 2328 2172 2332
rect 2166 2327 2172 2328
rect 2262 2332 2268 2333
rect 2262 2328 2263 2332
rect 2267 2328 2268 2332
rect 2262 2327 2268 2328
rect 2366 2332 2372 2333
rect 2366 2328 2367 2332
rect 2371 2328 2372 2332
rect 2366 2327 2372 2328
rect 2470 2332 2476 2333
rect 2470 2328 2471 2332
rect 2475 2328 2476 2332
rect 2470 2327 2476 2328
rect 2574 2332 2580 2333
rect 2574 2328 2575 2332
rect 2579 2328 2580 2332
rect 2574 2327 2580 2328
rect 2686 2332 2692 2333
rect 2686 2328 2687 2332
rect 2691 2328 2692 2332
rect 2686 2327 2692 2328
rect 2798 2332 2804 2333
rect 2798 2328 2799 2332
rect 2803 2328 2804 2332
rect 2798 2327 2804 2328
rect 2910 2332 2916 2333
rect 2910 2328 2911 2332
rect 2915 2328 2916 2332
rect 2910 2327 2916 2328
rect 3022 2332 3028 2333
rect 3022 2328 3023 2332
rect 3027 2328 3028 2332
rect 3462 2331 3463 2335
rect 3467 2331 3468 2335
rect 3462 2330 3468 2331
rect 3022 2327 3028 2328
rect 555 2324 626 2326
rect 555 2323 556 2324
rect 550 2322 556 2323
rect 202 2287 208 2288
rect 202 2283 203 2287
rect 207 2286 208 2287
rect 2230 2287 2236 2288
rect 207 2284 602 2286
rect 207 2283 208 2284
rect 202 2282 208 2283
rect 150 2280 156 2281
rect 110 2277 116 2278
rect 110 2273 111 2277
rect 115 2273 116 2277
rect 150 2276 151 2280
rect 155 2276 156 2280
rect 150 2275 156 2276
rect 270 2280 276 2281
rect 270 2276 271 2280
rect 275 2276 276 2280
rect 270 2275 276 2276
rect 390 2280 396 2281
rect 390 2276 391 2280
rect 395 2276 396 2280
rect 390 2275 396 2276
rect 518 2280 524 2281
rect 518 2276 519 2280
rect 523 2276 524 2280
rect 518 2275 524 2276
rect 110 2272 116 2273
rect 222 2271 228 2272
rect 222 2267 223 2271
rect 227 2267 228 2271
rect 222 2266 228 2267
rect 342 2271 348 2272
rect 342 2267 343 2271
rect 347 2267 348 2271
rect 342 2266 348 2267
rect 462 2271 468 2272
rect 462 2267 463 2271
rect 467 2267 468 2271
rect 462 2266 468 2267
rect 590 2271 596 2272
rect 590 2267 591 2271
rect 595 2267 596 2271
rect 600 2270 602 2284
rect 2230 2283 2231 2287
rect 2235 2286 2236 2287
rect 2235 2284 2458 2286
rect 2235 2283 2236 2284
rect 2230 2282 2236 2283
rect 646 2280 652 2281
rect 646 2276 647 2280
rect 651 2276 652 2280
rect 646 2275 652 2276
rect 774 2280 780 2281
rect 774 2276 775 2280
rect 779 2276 780 2280
rect 774 2275 780 2276
rect 894 2280 900 2281
rect 894 2276 895 2280
rect 899 2276 900 2280
rect 894 2275 900 2276
rect 1014 2280 1020 2281
rect 1014 2276 1015 2280
rect 1019 2276 1020 2280
rect 1014 2275 1020 2276
rect 1142 2280 1148 2281
rect 1142 2276 1143 2280
rect 1147 2276 1148 2280
rect 1142 2275 1148 2276
rect 1270 2280 1276 2281
rect 1270 2276 1271 2280
rect 1275 2276 1276 2280
rect 1886 2280 1892 2281
rect 1270 2275 1276 2276
rect 1766 2277 1772 2278
rect 1766 2273 1767 2277
rect 1771 2273 1772 2277
rect 1766 2272 1772 2273
rect 1806 2277 1812 2278
rect 1806 2273 1807 2277
rect 1811 2273 1812 2277
rect 1886 2276 1887 2280
rect 1891 2276 1892 2280
rect 1886 2275 1892 2276
rect 2038 2280 2044 2281
rect 2038 2276 2039 2280
rect 2043 2276 2044 2280
rect 2038 2275 2044 2276
rect 2198 2280 2204 2281
rect 2198 2276 2199 2280
rect 2203 2276 2204 2280
rect 2198 2275 2204 2276
rect 2374 2280 2380 2281
rect 2374 2276 2375 2280
rect 2379 2276 2380 2280
rect 2374 2275 2380 2276
rect 1806 2272 1812 2273
rect 846 2271 852 2272
rect 600 2268 689 2270
rect 590 2266 596 2267
rect 846 2267 847 2271
rect 851 2267 852 2271
rect 846 2266 852 2267
rect 854 2271 860 2272
rect 854 2267 855 2271
rect 859 2270 860 2271
rect 1086 2271 1092 2272
rect 859 2268 937 2270
rect 859 2267 860 2268
rect 854 2266 860 2267
rect 1086 2267 1087 2271
rect 1091 2267 1092 2271
rect 1086 2266 1092 2267
rect 1214 2271 1220 2272
rect 1214 2267 1215 2271
rect 1219 2267 1220 2271
rect 1214 2266 1220 2267
rect 1222 2271 1228 2272
rect 1222 2267 1223 2271
rect 1227 2270 1228 2271
rect 1958 2271 1964 2272
rect 1227 2268 1313 2270
rect 1227 2267 1228 2268
rect 1222 2266 1228 2267
rect 1958 2267 1959 2271
rect 1963 2267 1964 2271
rect 1958 2266 1964 2267
rect 2110 2271 2116 2272
rect 2110 2267 2111 2271
rect 2115 2267 2116 2271
rect 2110 2266 2116 2267
rect 2270 2271 2276 2272
rect 2270 2267 2271 2271
rect 2275 2267 2276 2271
rect 2270 2266 2276 2267
rect 2446 2271 2452 2272
rect 2446 2267 2447 2271
rect 2451 2267 2452 2271
rect 2456 2270 2458 2284
rect 2550 2280 2556 2281
rect 2550 2276 2551 2280
rect 2555 2276 2556 2280
rect 2550 2275 2556 2276
rect 2718 2280 2724 2281
rect 2718 2276 2719 2280
rect 2723 2276 2724 2280
rect 2718 2275 2724 2276
rect 2886 2280 2892 2281
rect 2886 2276 2887 2280
rect 2891 2276 2892 2280
rect 2886 2275 2892 2276
rect 3054 2280 3060 2281
rect 3054 2276 3055 2280
rect 3059 2276 3060 2280
rect 3054 2275 3060 2276
rect 3222 2280 3228 2281
rect 3222 2276 3223 2280
rect 3227 2276 3228 2280
rect 3222 2275 3228 2276
rect 3366 2280 3372 2281
rect 3366 2276 3367 2280
rect 3371 2276 3372 2280
rect 3366 2275 3372 2276
rect 3462 2277 3468 2278
rect 3462 2273 3463 2277
rect 3467 2273 3468 2277
rect 3462 2272 3468 2273
rect 2706 2271 2712 2272
rect 2456 2268 2593 2270
rect 2446 2266 2452 2267
rect 2706 2267 2707 2271
rect 2711 2270 2712 2271
rect 2798 2271 2804 2272
rect 2711 2268 2761 2270
rect 2711 2267 2712 2268
rect 2706 2266 2712 2267
rect 2798 2267 2799 2271
rect 2803 2270 2804 2271
rect 3126 2271 3132 2272
rect 2803 2268 2929 2270
rect 2803 2267 2804 2268
rect 2798 2266 2804 2267
rect 3126 2267 3127 2271
rect 3131 2267 3132 2271
rect 3126 2266 3132 2267
rect 3294 2271 3300 2272
rect 3294 2267 3295 2271
rect 3299 2267 3300 2271
rect 3294 2266 3300 2267
rect 3430 2271 3436 2272
rect 3430 2267 3431 2271
rect 3435 2267 3436 2271
rect 3430 2266 3436 2267
rect 150 2261 156 2262
rect 110 2260 116 2261
rect 110 2256 111 2260
rect 115 2256 116 2260
rect 150 2257 151 2261
rect 155 2257 156 2261
rect 150 2256 156 2257
rect 270 2261 276 2262
rect 270 2257 271 2261
rect 275 2257 276 2261
rect 270 2256 276 2257
rect 390 2261 396 2262
rect 390 2257 391 2261
rect 395 2257 396 2261
rect 390 2256 396 2257
rect 518 2261 524 2262
rect 518 2257 519 2261
rect 523 2257 524 2261
rect 518 2256 524 2257
rect 646 2261 652 2262
rect 646 2257 647 2261
rect 651 2257 652 2261
rect 646 2256 652 2257
rect 774 2261 780 2262
rect 774 2257 775 2261
rect 779 2257 780 2261
rect 774 2256 780 2257
rect 894 2261 900 2262
rect 894 2257 895 2261
rect 899 2257 900 2261
rect 894 2256 900 2257
rect 1014 2261 1020 2262
rect 1014 2257 1015 2261
rect 1019 2257 1020 2261
rect 1014 2256 1020 2257
rect 1142 2261 1148 2262
rect 1142 2257 1143 2261
rect 1147 2257 1148 2261
rect 1142 2256 1148 2257
rect 1270 2261 1276 2262
rect 1886 2261 1892 2262
rect 1270 2257 1271 2261
rect 1275 2257 1276 2261
rect 1270 2256 1276 2257
rect 1766 2260 1772 2261
rect 1766 2256 1767 2260
rect 1771 2256 1772 2260
rect 110 2255 116 2256
rect 1766 2255 1772 2256
rect 1806 2260 1812 2261
rect 1806 2256 1807 2260
rect 1811 2256 1812 2260
rect 1886 2257 1887 2261
rect 1891 2257 1892 2261
rect 1886 2256 1892 2257
rect 2038 2261 2044 2262
rect 2038 2257 2039 2261
rect 2043 2257 2044 2261
rect 2038 2256 2044 2257
rect 2198 2261 2204 2262
rect 2198 2257 2199 2261
rect 2203 2257 2204 2261
rect 2198 2256 2204 2257
rect 2374 2261 2380 2262
rect 2374 2257 2375 2261
rect 2379 2257 2380 2261
rect 2374 2256 2380 2257
rect 2550 2261 2556 2262
rect 2550 2257 2551 2261
rect 2555 2257 2556 2261
rect 2550 2256 2556 2257
rect 2718 2261 2724 2262
rect 2718 2257 2719 2261
rect 2723 2257 2724 2261
rect 2718 2256 2724 2257
rect 2886 2261 2892 2262
rect 2886 2257 2887 2261
rect 2891 2257 2892 2261
rect 2886 2256 2892 2257
rect 3054 2261 3060 2262
rect 3054 2257 3055 2261
rect 3059 2257 3060 2261
rect 3054 2256 3060 2257
rect 3222 2261 3228 2262
rect 3222 2257 3223 2261
rect 3227 2257 3228 2261
rect 3222 2256 3228 2257
rect 3366 2261 3372 2262
rect 3366 2257 3367 2261
rect 3371 2257 3372 2261
rect 3366 2256 3372 2257
rect 3462 2260 3468 2261
rect 3462 2256 3463 2260
rect 3467 2256 3468 2260
rect 1806 2255 1812 2256
rect 3462 2255 3468 2256
rect 199 2243 208 2244
rect 199 2239 200 2243
rect 207 2239 208 2243
rect 199 2238 208 2239
rect 222 2243 228 2244
rect 222 2239 223 2243
rect 227 2242 228 2243
rect 319 2243 325 2244
rect 319 2242 320 2243
rect 227 2240 320 2242
rect 227 2239 228 2240
rect 222 2238 228 2239
rect 319 2239 320 2240
rect 324 2239 325 2243
rect 319 2238 325 2239
rect 398 2243 404 2244
rect 398 2239 399 2243
rect 403 2242 404 2243
rect 439 2243 445 2244
rect 439 2242 440 2243
rect 403 2240 440 2242
rect 403 2239 404 2240
rect 398 2238 404 2239
rect 439 2239 440 2240
rect 444 2239 445 2243
rect 439 2238 445 2239
rect 462 2243 468 2244
rect 462 2239 463 2243
rect 467 2242 468 2243
rect 567 2243 573 2244
rect 567 2242 568 2243
rect 467 2240 568 2242
rect 467 2239 468 2240
rect 462 2238 468 2239
rect 567 2239 568 2240
rect 572 2239 573 2243
rect 567 2238 573 2239
rect 590 2243 596 2244
rect 590 2239 591 2243
rect 595 2242 596 2243
rect 695 2243 701 2244
rect 695 2242 696 2243
rect 595 2240 696 2242
rect 595 2239 596 2240
rect 590 2238 596 2239
rect 695 2239 696 2240
rect 700 2239 701 2243
rect 695 2238 701 2239
rect 823 2243 829 2244
rect 823 2239 824 2243
rect 828 2242 829 2243
rect 854 2243 860 2244
rect 854 2242 855 2243
rect 828 2240 855 2242
rect 828 2239 829 2240
rect 823 2238 829 2239
rect 854 2239 855 2240
rect 859 2239 860 2243
rect 854 2238 860 2239
rect 942 2243 949 2244
rect 942 2239 943 2243
rect 948 2239 949 2243
rect 942 2238 949 2239
rect 1063 2243 1069 2244
rect 1063 2239 1064 2243
rect 1068 2239 1069 2243
rect 1063 2238 1069 2239
rect 1086 2243 1092 2244
rect 1086 2239 1087 2243
rect 1091 2242 1092 2243
rect 1191 2243 1197 2244
rect 1191 2242 1192 2243
rect 1091 2240 1192 2242
rect 1091 2239 1092 2240
rect 1086 2238 1092 2239
rect 1191 2239 1192 2240
rect 1196 2239 1197 2243
rect 1191 2238 1197 2239
rect 1214 2243 1220 2244
rect 1214 2239 1215 2243
rect 1219 2242 1220 2243
rect 1319 2243 1325 2244
rect 1319 2242 1320 2243
rect 1219 2240 1320 2242
rect 1219 2239 1220 2240
rect 1214 2238 1220 2239
rect 1319 2239 1320 2240
rect 1324 2239 1325 2243
rect 1319 2238 1325 2239
rect 1935 2243 1941 2244
rect 1935 2239 1936 2243
rect 1940 2242 1941 2243
rect 1950 2243 1956 2244
rect 1950 2242 1951 2243
rect 1940 2240 1951 2242
rect 1940 2239 1941 2240
rect 1935 2238 1941 2239
rect 1950 2239 1951 2240
rect 1955 2239 1956 2243
rect 1950 2238 1956 2239
rect 1958 2243 1964 2244
rect 1958 2239 1959 2243
rect 1963 2242 1964 2243
rect 2087 2243 2093 2244
rect 2087 2242 2088 2243
rect 1963 2240 2088 2242
rect 1963 2239 1964 2240
rect 1958 2238 1964 2239
rect 2087 2239 2088 2240
rect 2092 2239 2093 2243
rect 2087 2238 2093 2239
rect 2110 2243 2116 2244
rect 2110 2239 2111 2243
rect 2115 2242 2116 2243
rect 2247 2243 2253 2244
rect 2247 2242 2248 2243
rect 2115 2240 2248 2242
rect 2115 2239 2116 2240
rect 2110 2238 2116 2239
rect 2247 2239 2248 2240
rect 2252 2239 2253 2243
rect 2247 2238 2253 2239
rect 2270 2243 2276 2244
rect 2270 2239 2271 2243
rect 2275 2242 2276 2243
rect 2423 2243 2429 2244
rect 2423 2242 2424 2243
rect 2275 2240 2424 2242
rect 2275 2239 2276 2240
rect 2270 2238 2276 2239
rect 2423 2239 2424 2240
rect 2428 2239 2429 2243
rect 2423 2238 2429 2239
rect 2446 2243 2452 2244
rect 2446 2239 2447 2243
rect 2451 2242 2452 2243
rect 2599 2243 2605 2244
rect 2599 2242 2600 2243
rect 2451 2240 2600 2242
rect 2451 2239 2452 2240
rect 2446 2238 2452 2239
rect 2599 2239 2600 2240
rect 2604 2239 2605 2243
rect 2599 2238 2605 2239
rect 2767 2243 2773 2244
rect 2767 2239 2768 2243
rect 2772 2242 2773 2243
rect 2798 2243 2804 2244
rect 2798 2242 2799 2243
rect 2772 2240 2799 2242
rect 2772 2239 2773 2240
rect 2767 2238 2773 2239
rect 2798 2239 2799 2240
rect 2803 2239 2804 2243
rect 2798 2238 2804 2239
rect 2935 2243 2941 2244
rect 2935 2239 2936 2243
rect 2940 2242 2941 2243
rect 2990 2243 2996 2244
rect 2990 2242 2991 2243
rect 2940 2240 2991 2242
rect 2940 2239 2941 2240
rect 2935 2238 2941 2239
rect 2990 2239 2991 2240
rect 2995 2239 2996 2243
rect 2990 2238 2996 2239
rect 3030 2243 3036 2244
rect 3030 2239 3031 2243
rect 3035 2242 3036 2243
rect 3103 2243 3109 2244
rect 3103 2242 3104 2243
rect 3035 2240 3104 2242
rect 3035 2239 3036 2240
rect 3030 2238 3036 2239
rect 3103 2239 3104 2240
rect 3108 2239 3109 2243
rect 3103 2238 3109 2239
rect 3126 2243 3132 2244
rect 3126 2239 3127 2243
rect 3131 2242 3132 2243
rect 3271 2243 3277 2244
rect 3271 2242 3272 2243
rect 3131 2240 3272 2242
rect 3131 2239 3132 2240
rect 3126 2238 3132 2239
rect 3271 2239 3272 2240
rect 3276 2239 3277 2243
rect 3271 2238 3277 2239
rect 3294 2243 3300 2244
rect 3294 2239 3295 2243
rect 3299 2242 3300 2243
rect 3415 2243 3421 2244
rect 3415 2242 3416 2243
rect 3299 2240 3416 2242
rect 3299 2239 3300 2240
rect 3294 2238 3300 2239
rect 3415 2239 3416 2240
rect 3420 2239 3421 2243
rect 3415 2238 3421 2239
rect 738 2235 744 2236
rect 738 2234 739 2235
rect 319 2232 739 2234
rect 183 2227 189 2228
rect 183 2223 184 2227
rect 188 2226 189 2227
rect 214 2227 220 2228
rect 214 2226 215 2227
rect 188 2224 215 2226
rect 188 2223 189 2224
rect 183 2222 189 2223
rect 214 2223 215 2224
rect 219 2223 220 2227
rect 214 2222 220 2223
rect 295 2227 301 2228
rect 295 2223 296 2227
rect 300 2226 301 2227
rect 319 2226 321 2232
rect 738 2231 739 2232
rect 743 2231 744 2235
rect 738 2230 744 2231
rect 1742 2231 1748 2232
rect 300 2224 321 2226
rect 342 2227 348 2228
rect 300 2223 301 2224
rect 295 2222 301 2223
rect 342 2223 343 2227
rect 347 2226 348 2227
rect 455 2227 461 2228
rect 455 2226 456 2227
rect 347 2224 456 2226
rect 347 2223 348 2224
rect 342 2222 348 2223
rect 455 2223 456 2224
rect 460 2223 461 2227
rect 455 2222 461 2223
rect 478 2227 484 2228
rect 478 2223 479 2227
rect 483 2226 484 2227
rect 631 2227 637 2228
rect 631 2226 632 2227
rect 483 2224 632 2226
rect 483 2223 484 2224
rect 478 2222 484 2223
rect 631 2223 632 2224
rect 636 2223 637 2227
rect 631 2222 637 2223
rect 654 2227 660 2228
rect 654 2223 655 2227
rect 659 2226 660 2227
rect 815 2227 821 2228
rect 815 2226 816 2227
rect 659 2224 816 2226
rect 659 2223 660 2224
rect 654 2222 660 2223
rect 815 2223 816 2224
rect 820 2223 821 2227
rect 815 2222 821 2223
rect 999 2227 1005 2228
rect 999 2223 1000 2227
rect 1004 2226 1005 2227
rect 1078 2227 1084 2228
rect 1078 2226 1079 2227
rect 1004 2224 1079 2226
rect 1004 2223 1005 2224
rect 999 2222 1005 2223
rect 1078 2223 1079 2224
rect 1083 2223 1084 2227
rect 1078 2222 1084 2223
rect 1183 2227 1189 2228
rect 1183 2223 1184 2227
rect 1188 2226 1189 2227
rect 1222 2227 1228 2228
rect 1222 2226 1223 2227
rect 1188 2224 1223 2226
rect 1188 2223 1189 2224
rect 1183 2222 1189 2223
rect 1222 2223 1223 2224
rect 1227 2223 1228 2227
rect 1222 2222 1228 2223
rect 1302 2227 1308 2228
rect 1302 2223 1303 2227
rect 1307 2226 1308 2227
rect 1367 2227 1373 2228
rect 1367 2226 1368 2227
rect 1307 2224 1368 2226
rect 1307 2223 1308 2224
rect 1302 2222 1308 2223
rect 1367 2223 1368 2224
rect 1372 2223 1373 2227
rect 1367 2222 1373 2223
rect 1390 2227 1396 2228
rect 1390 2223 1391 2227
rect 1395 2226 1396 2227
rect 1551 2227 1557 2228
rect 1551 2226 1552 2227
rect 1395 2224 1552 2226
rect 1395 2223 1396 2224
rect 1390 2222 1396 2223
rect 1551 2223 1552 2224
rect 1556 2223 1557 2227
rect 1551 2222 1557 2223
rect 1574 2227 1580 2228
rect 1574 2223 1575 2227
rect 1579 2226 1580 2227
rect 1719 2227 1725 2228
rect 1719 2226 1720 2227
rect 1579 2224 1720 2226
rect 1579 2223 1580 2224
rect 1574 2222 1580 2223
rect 1719 2223 1720 2224
rect 1724 2223 1725 2227
rect 1742 2227 1743 2231
rect 1747 2230 1748 2231
rect 1879 2231 1885 2232
rect 1879 2230 1880 2231
rect 1747 2228 1880 2230
rect 1747 2227 1748 2228
rect 1742 2226 1748 2227
rect 1879 2227 1880 2228
rect 1884 2227 1885 2231
rect 1879 2226 1885 2227
rect 1902 2231 1908 2232
rect 1902 2227 1903 2231
rect 1907 2230 1908 2231
rect 2015 2231 2021 2232
rect 2015 2230 2016 2231
rect 1907 2228 2016 2230
rect 1907 2227 1908 2228
rect 1902 2226 1908 2227
rect 2015 2227 2016 2228
rect 2020 2227 2021 2231
rect 2015 2226 2021 2227
rect 2079 2231 2085 2232
rect 2079 2227 2080 2231
rect 2084 2230 2085 2231
rect 2183 2231 2189 2232
rect 2183 2230 2184 2231
rect 2084 2228 2184 2230
rect 2084 2227 2085 2228
rect 2079 2226 2085 2227
rect 2183 2227 2184 2228
rect 2188 2227 2189 2231
rect 2183 2226 2189 2227
rect 2206 2231 2212 2232
rect 2206 2227 2207 2231
rect 2211 2230 2212 2231
rect 2359 2231 2365 2232
rect 2359 2230 2360 2231
rect 2211 2228 2360 2230
rect 2211 2227 2212 2228
rect 2206 2226 2212 2227
rect 2359 2227 2360 2228
rect 2364 2227 2365 2231
rect 2359 2226 2365 2227
rect 2382 2231 2388 2232
rect 2382 2227 2383 2231
rect 2387 2230 2388 2231
rect 2535 2231 2541 2232
rect 2535 2230 2536 2231
rect 2387 2228 2536 2230
rect 2387 2227 2388 2228
rect 2382 2226 2388 2227
rect 2535 2227 2536 2228
rect 2540 2227 2541 2231
rect 2535 2226 2541 2227
rect 2703 2231 2712 2232
rect 2703 2227 2704 2231
rect 2711 2227 2712 2231
rect 2703 2226 2712 2227
rect 2726 2231 2732 2232
rect 2726 2227 2727 2231
rect 2731 2230 2732 2231
rect 2863 2231 2869 2232
rect 2863 2230 2864 2231
rect 2731 2228 2864 2230
rect 2731 2227 2732 2228
rect 2726 2226 2732 2227
rect 2863 2227 2864 2228
rect 2868 2227 2869 2231
rect 2863 2226 2869 2227
rect 3007 2231 3013 2232
rect 3007 2227 3008 2231
rect 3012 2230 3013 2231
rect 3038 2231 3044 2232
rect 3038 2230 3039 2231
rect 3012 2228 3039 2230
rect 3012 2227 3013 2228
rect 3007 2226 3013 2227
rect 3038 2227 3039 2228
rect 3043 2227 3044 2231
rect 3038 2226 3044 2227
rect 3151 2231 3157 2232
rect 3151 2227 3152 2231
rect 3156 2230 3157 2231
rect 3182 2231 3188 2232
rect 3182 2230 3183 2231
rect 3156 2228 3183 2230
rect 3156 2227 3157 2228
rect 3151 2226 3157 2227
rect 3182 2227 3183 2228
rect 3187 2227 3188 2231
rect 3182 2226 3188 2227
rect 3191 2231 3197 2232
rect 3191 2227 3192 2231
rect 3196 2230 3197 2231
rect 3295 2231 3301 2232
rect 3295 2230 3296 2231
rect 3196 2228 3296 2230
rect 3196 2227 3197 2228
rect 3191 2226 3197 2227
rect 3295 2227 3296 2228
rect 3300 2227 3301 2231
rect 3295 2226 3301 2227
rect 3415 2231 3421 2232
rect 3415 2227 3416 2231
rect 3420 2230 3421 2231
rect 3430 2231 3436 2232
rect 3430 2230 3431 2231
rect 3420 2228 3431 2230
rect 3420 2227 3421 2228
rect 3415 2226 3421 2227
rect 3430 2227 3431 2228
rect 3435 2227 3436 2231
rect 3430 2226 3436 2227
rect 1719 2222 1725 2223
rect 1806 2216 1812 2217
rect 3462 2216 3468 2217
rect 110 2212 116 2213
rect 1766 2212 1772 2213
rect 110 2208 111 2212
rect 115 2208 116 2212
rect 110 2207 116 2208
rect 134 2211 140 2212
rect 134 2207 135 2211
rect 139 2207 140 2211
rect 134 2206 140 2207
rect 246 2211 252 2212
rect 246 2207 247 2211
rect 251 2207 252 2211
rect 246 2206 252 2207
rect 406 2211 412 2212
rect 406 2207 407 2211
rect 411 2207 412 2211
rect 406 2206 412 2207
rect 582 2211 588 2212
rect 582 2207 583 2211
rect 587 2207 588 2211
rect 582 2206 588 2207
rect 766 2211 772 2212
rect 766 2207 767 2211
rect 771 2207 772 2211
rect 766 2206 772 2207
rect 950 2211 956 2212
rect 950 2207 951 2211
rect 955 2207 956 2211
rect 950 2206 956 2207
rect 1134 2211 1140 2212
rect 1134 2207 1135 2211
rect 1139 2207 1140 2211
rect 1134 2206 1140 2207
rect 1318 2211 1324 2212
rect 1318 2207 1319 2211
rect 1323 2207 1324 2211
rect 1318 2206 1324 2207
rect 1502 2211 1508 2212
rect 1502 2207 1503 2211
rect 1507 2207 1508 2211
rect 1502 2206 1508 2207
rect 1670 2211 1676 2212
rect 1670 2207 1671 2211
rect 1675 2207 1676 2211
rect 1766 2208 1767 2212
rect 1771 2208 1772 2212
rect 1806 2212 1807 2216
rect 1811 2212 1812 2216
rect 1806 2211 1812 2212
rect 1830 2215 1836 2216
rect 1830 2211 1831 2215
rect 1835 2211 1836 2215
rect 1830 2210 1836 2211
rect 1966 2215 1972 2216
rect 1966 2211 1967 2215
rect 1971 2211 1972 2215
rect 1966 2210 1972 2211
rect 2134 2215 2140 2216
rect 2134 2211 2135 2215
rect 2139 2211 2140 2215
rect 2134 2210 2140 2211
rect 2310 2215 2316 2216
rect 2310 2211 2311 2215
rect 2315 2211 2316 2215
rect 2310 2210 2316 2211
rect 2486 2215 2492 2216
rect 2486 2211 2487 2215
rect 2491 2211 2492 2215
rect 2486 2210 2492 2211
rect 2654 2215 2660 2216
rect 2654 2211 2655 2215
rect 2659 2211 2660 2215
rect 2654 2210 2660 2211
rect 2814 2215 2820 2216
rect 2814 2211 2815 2215
rect 2819 2211 2820 2215
rect 2814 2210 2820 2211
rect 2958 2215 2964 2216
rect 2958 2211 2959 2215
rect 2963 2211 2964 2215
rect 2958 2210 2964 2211
rect 3102 2215 3108 2216
rect 3102 2211 3103 2215
rect 3107 2211 3108 2215
rect 3102 2210 3108 2211
rect 3246 2215 3252 2216
rect 3246 2211 3247 2215
rect 3251 2211 3252 2215
rect 3246 2210 3252 2211
rect 3366 2215 3372 2216
rect 3366 2211 3367 2215
rect 3371 2211 3372 2215
rect 3462 2212 3463 2216
rect 3467 2212 3468 2216
rect 3462 2211 3468 2212
rect 3366 2210 3372 2211
rect 1766 2207 1772 2208
rect 1902 2207 1908 2208
rect 1670 2206 1676 2207
rect 214 2203 220 2204
rect 214 2199 215 2203
rect 219 2202 220 2203
rect 478 2203 484 2204
rect 219 2200 289 2202
rect 219 2199 220 2200
rect 214 2198 220 2199
rect 478 2199 479 2203
rect 483 2199 484 2203
rect 478 2198 484 2199
rect 654 2203 660 2204
rect 654 2199 655 2203
rect 659 2199 660 2203
rect 654 2198 660 2199
rect 738 2203 744 2204
rect 738 2199 739 2203
rect 743 2202 744 2203
rect 942 2203 948 2204
rect 743 2200 809 2202
rect 743 2199 744 2200
rect 738 2198 744 2199
rect 942 2199 943 2203
rect 947 2202 948 2203
rect 1078 2203 1084 2204
rect 947 2200 993 2202
rect 947 2199 948 2200
rect 942 2198 948 2199
rect 1078 2199 1079 2203
rect 1083 2202 1084 2203
rect 1390 2203 1396 2204
rect 1083 2200 1177 2202
rect 1083 2199 1084 2200
rect 1078 2198 1084 2199
rect 1390 2199 1391 2203
rect 1395 2199 1396 2203
rect 1390 2198 1396 2199
rect 1574 2203 1580 2204
rect 1574 2199 1575 2203
rect 1579 2199 1580 2203
rect 1574 2198 1580 2199
rect 1742 2203 1748 2204
rect 1742 2199 1743 2203
rect 1747 2199 1748 2203
rect 1902 2203 1903 2207
rect 1907 2203 1908 2207
rect 2079 2207 2085 2208
rect 2079 2206 2080 2207
rect 2041 2204 2080 2206
rect 1902 2202 1908 2203
rect 2079 2203 2080 2204
rect 2084 2203 2085 2207
rect 2079 2202 2085 2203
rect 2206 2207 2212 2208
rect 2206 2203 2207 2207
rect 2211 2203 2212 2207
rect 2206 2202 2212 2203
rect 2382 2207 2388 2208
rect 2382 2203 2383 2207
rect 2387 2203 2388 2207
rect 2382 2202 2388 2203
rect 2418 2207 2424 2208
rect 2418 2203 2419 2207
rect 2423 2206 2424 2207
rect 2726 2207 2732 2208
rect 2423 2204 2529 2206
rect 2423 2203 2424 2204
rect 2418 2202 2424 2203
rect 2726 2203 2727 2207
rect 2731 2203 2732 2207
rect 3030 2207 3036 2208
rect 2726 2202 2732 2203
rect 2886 2203 2892 2204
rect 1742 2198 1748 2199
rect 1806 2199 1812 2200
rect 110 2195 116 2196
rect 110 2191 111 2195
rect 115 2191 116 2195
rect 198 2195 204 2196
rect 110 2190 116 2191
rect 134 2192 140 2193
rect 134 2188 135 2192
rect 139 2188 140 2192
rect 198 2191 199 2195
rect 203 2194 204 2195
rect 208 2194 210 2197
rect 203 2192 210 2194
rect 1766 2195 1772 2196
rect 246 2192 252 2193
rect 203 2191 204 2192
rect 198 2190 204 2191
rect 134 2187 140 2188
rect 246 2188 247 2192
rect 251 2188 252 2192
rect 246 2187 252 2188
rect 406 2192 412 2193
rect 406 2188 407 2192
rect 411 2188 412 2192
rect 406 2187 412 2188
rect 582 2192 588 2193
rect 582 2188 583 2192
rect 587 2188 588 2192
rect 582 2187 588 2188
rect 766 2192 772 2193
rect 766 2188 767 2192
rect 771 2188 772 2192
rect 766 2187 772 2188
rect 950 2192 956 2193
rect 950 2188 951 2192
rect 955 2188 956 2192
rect 950 2187 956 2188
rect 1134 2192 1140 2193
rect 1134 2188 1135 2192
rect 1139 2188 1140 2192
rect 1134 2187 1140 2188
rect 1318 2192 1324 2193
rect 1318 2188 1319 2192
rect 1323 2188 1324 2192
rect 1318 2187 1324 2188
rect 1502 2192 1508 2193
rect 1502 2188 1503 2192
rect 1507 2188 1508 2192
rect 1502 2187 1508 2188
rect 1670 2192 1676 2193
rect 1670 2188 1671 2192
rect 1675 2188 1676 2192
rect 1766 2191 1767 2195
rect 1771 2191 1772 2195
rect 1806 2195 1807 2199
rect 1811 2195 1812 2199
rect 2886 2199 2887 2203
rect 2891 2199 2892 2203
rect 3030 2203 3031 2207
rect 3035 2203 3036 2207
rect 3030 2202 3036 2203
rect 3038 2207 3044 2208
rect 3038 2203 3039 2207
rect 3043 2206 3044 2207
rect 3182 2207 3188 2208
rect 3043 2204 3145 2206
rect 3043 2203 3044 2204
rect 3038 2202 3044 2203
rect 3182 2203 3183 2207
rect 3187 2206 3188 2207
rect 3187 2204 3289 2206
rect 3187 2203 3188 2204
rect 3182 2202 3188 2203
rect 3438 2203 3444 2204
rect 2886 2198 2892 2199
rect 3438 2199 3439 2203
rect 3443 2199 3444 2203
rect 3438 2198 3444 2199
rect 3462 2199 3468 2200
rect 1806 2194 1812 2195
rect 1830 2196 1836 2197
rect 1830 2192 1831 2196
rect 1835 2192 1836 2196
rect 1830 2191 1836 2192
rect 1966 2196 1972 2197
rect 1966 2192 1967 2196
rect 1971 2192 1972 2196
rect 1966 2191 1972 2192
rect 2134 2196 2140 2197
rect 2134 2192 2135 2196
rect 2139 2192 2140 2196
rect 2134 2191 2140 2192
rect 2310 2196 2316 2197
rect 2310 2192 2311 2196
rect 2315 2192 2316 2196
rect 2310 2191 2316 2192
rect 2486 2196 2492 2197
rect 2486 2192 2487 2196
rect 2491 2192 2492 2196
rect 2486 2191 2492 2192
rect 2654 2196 2660 2197
rect 2654 2192 2655 2196
rect 2659 2192 2660 2196
rect 2654 2191 2660 2192
rect 2814 2196 2820 2197
rect 2814 2192 2815 2196
rect 2819 2192 2820 2196
rect 2814 2191 2820 2192
rect 2958 2196 2964 2197
rect 2958 2192 2959 2196
rect 2963 2192 2964 2196
rect 2958 2191 2964 2192
rect 3102 2196 3108 2197
rect 3102 2192 3103 2196
rect 3107 2192 3108 2196
rect 3102 2191 3108 2192
rect 3246 2196 3252 2197
rect 3246 2192 3247 2196
rect 3251 2192 3252 2196
rect 3246 2191 3252 2192
rect 3366 2196 3372 2197
rect 3366 2192 3367 2196
rect 3371 2192 3372 2196
rect 3462 2195 3463 2199
rect 3467 2195 3468 2199
rect 3462 2194 3468 2195
rect 3366 2191 3372 2192
rect 1766 2190 1772 2191
rect 1670 2187 1676 2188
rect 1950 2187 1956 2188
rect 1950 2183 1951 2187
rect 1955 2186 1956 2187
rect 2418 2187 2424 2188
rect 2418 2186 2419 2187
rect 1955 2184 2419 2186
rect 1955 2183 1956 2184
rect 1950 2182 1956 2183
rect 2418 2183 2419 2184
rect 2423 2183 2424 2187
rect 2418 2182 2424 2183
rect 2926 2152 2932 2153
rect 1806 2149 1812 2150
rect 1806 2145 1807 2149
rect 1811 2145 1812 2149
rect 2926 2148 2927 2152
rect 2931 2148 2932 2152
rect 2926 2147 2932 2148
rect 3014 2152 3020 2153
rect 3014 2148 3015 2152
rect 3019 2148 3020 2152
rect 3014 2147 3020 2148
rect 3102 2152 3108 2153
rect 3102 2148 3103 2152
rect 3107 2148 3108 2152
rect 3102 2147 3108 2148
rect 3190 2152 3196 2153
rect 3190 2148 3191 2152
rect 3195 2148 3196 2152
rect 3190 2147 3196 2148
rect 3278 2152 3284 2153
rect 3278 2148 3279 2152
rect 3283 2148 3284 2152
rect 3278 2147 3284 2148
rect 3366 2152 3372 2153
rect 3366 2148 3367 2152
rect 3371 2148 3372 2152
rect 3366 2147 3372 2148
rect 3462 2149 3468 2150
rect 1806 2144 1812 2145
rect 3462 2145 3463 2149
rect 3467 2145 3468 2149
rect 3462 2144 3468 2145
rect 2998 2143 3004 2144
rect 134 2140 140 2141
rect 110 2137 116 2138
rect 110 2133 111 2137
rect 115 2133 116 2137
rect 134 2136 135 2140
rect 139 2136 140 2140
rect 134 2135 140 2136
rect 246 2140 252 2141
rect 246 2136 247 2140
rect 251 2136 252 2140
rect 246 2135 252 2136
rect 390 2140 396 2141
rect 390 2136 391 2140
rect 395 2136 396 2140
rect 390 2135 396 2136
rect 542 2140 548 2141
rect 542 2136 543 2140
rect 547 2136 548 2140
rect 542 2135 548 2136
rect 694 2140 700 2141
rect 694 2136 695 2140
rect 699 2136 700 2140
rect 694 2135 700 2136
rect 838 2140 844 2141
rect 838 2136 839 2140
rect 843 2136 844 2140
rect 838 2135 844 2136
rect 974 2140 980 2141
rect 974 2136 975 2140
rect 979 2136 980 2140
rect 974 2135 980 2136
rect 1102 2140 1108 2141
rect 1102 2136 1103 2140
rect 1107 2136 1108 2140
rect 1102 2135 1108 2136
rect 1230 2140 1236 2141
rect 1230 2136 1231 2140
rect 1235 2136 1236 2140
rect 1230 2135 1236 2136
rect 1350 2140 1356 2141
rect 1350 2136 1351 2140
rect 1355 2136 1356 2140
rect 1350 2135 1356 2136
rect 1462 2140 1468 2141
rect 1462 2136 1463 2140
rect 1467 2136 1468 2140
rect 1462 2135 1468 2136
rect 1574 2140 1580 2141
rect 1574 2136 1575 2140
rect 1579 2136 1580 2140
rect 1574 2135 1580 2136
rect 1670 2140 1676 2141
rect 1670 2136 1671 2140
rect 1675 2136 1676 2140
rect 2998 2139 2999 2143
rect 3003 2139 3004 2143
rect 2998 2138 3004 2139
rect 3086 2143 3092 2144
rect 3086 2139 3087 2143
rect 3091 2139 3092 2143
rect 3183 2143 3189 2144
rect 3183 2142 3184 2143
rect 3177 2140 3184 2142
rect 3086 2138 3092 2139
rect 3183 2139 3184 2140
rect 3188 2139 3189 2143
rect 3183 2138 3189 2139
rect 3254 2143 3260 2144
rect 3254 2139 3255 2143
rect 3259 2139 3260 2143
rect 3254 2138 3260 2139
rect 3350 2143 3356 2144
rect 3350 2139 3351 2143
rect 3355 2139 3356 2143
rect 3350 2138 3356 2139
rect 3358 2143 3364 2144
rect 3358 2139 3359 2143
rect 3363 2142 3364 2143
rect 3363 2140 3409 2142
rect 3363 2139 3364 2140
rect 3358 2138 3364 2139
rect 1670 2135 1676 2136
rect 1766 2137 1772 2138
rect 110 2132 116 2133
rect 1766 2133 1767 2137
rect 1771 2133 1772 2137
rect 2926 2133 2932 2134
rect 1766 2132 1772 2133
rect 1806 2132 1812 2133
rect 206 2131 212 2132
rect 206 2127 207 2131
rect 211 2127 212 2131
rect 206 2126 212 2127
rect 318 2131 324 2132
rect 318 2127 319 2131
rect 323 2127 324 2131
rect 318 2126 324 2127
rect 462 2131 468 2132
rect 462 2127 463 2131
rect 467 2127 468 2131
rect 462 2126 468 2127
rect 614 2131 620 2132
rect 614 2127 615 2131
rect 619 2127 620 2131
rect 614 2126 620 2127
rect 622 2131 628 2132
rect 622 2127 623 2131
rect 627 2130 628 2131
rect 950 2131 956 2132
rect 950 2130 951 2131
rect 627 2128 737 2130
rect 913 2128 951 2130
rect 627 2127 628 2128
rect 622 2126 628 2127
rect 950 2127 951 2128
rect 955 2127 956 2131
rect 1054 2131 1060 2132
rect 1054 2130 1055 2131
rect 1049 2128 1055 2130
rect 950 2126 956 2127
rect 1054 2127 1055 2128
rect 1059 2127 1060 2131
rect 1054 2126 1060 2127
rect 1174 2131 1180 2132
rect 1174 2127 1175 2131
rect 1179 2127 1180 2131
rect 1174 2126 1180 2127
rect 1302 2131 1308 2132
rect 1302 2127 1303 2131
rect 1307 2127 1308 2131
rect 1302 2126 1308 2127
rect 1310 2131 1316 2132
rect 1310 2127 1311 2131
rect 1315 2130 1316 2131
rect 1430 2131 1436 2132
rect 1315 2128 1393 2130
rect 1315 2127 1316 2128
rect 1310 2126 1316 2127
rect 1430 2127 1431 2131
rect 1435 2130 1436 2131
rect 1542 2131 1548 2132
rect 1435 2128 1505 2130
rect 1435 2127 1436 2128
rect 1430 2126 1436 2127
rect 1542 2127 1543 2131
rect 1547 2130 1548 2131
rect 1654 2131 1660 2132
rect 1547 2128 1617 2130
rect 1547 2127 1548 2128
rect 1542 2126 1548 2127
rect 1654 2127 1655 2131
rect 1659 2130 1660 2131
rect 1659 2128 1713 2130
rect 1806 2128 1807 2132
rect 1811 2128 1812 2132
rect 2926 2129 2927 2133
rect 2931 2129 2932 2133
rect 2926 2128 2932 2129
rect 3014 2133 3020 2134
rect 3014 2129 3015 2133
rect 3019 2129 3020 2133
rect 3014 2128 3020 2129
rect 3102 2133 3108 2134
rect 3102 2129 3103 2133
rect 3107 2129 3108 2133
rect 3102 2128 3108 2129
rect 3190 2133 3196 2134
rect 3190 2129 3191 2133
rect 3195 2129 3196 2133
rect 3190 2128 3196 2129
rect 3278 2133 3284 2134
rect 3278 2129 3279 2133
rect 3283 2129 3284 2133
rect 3278 2128 3284 2129
rect 3366 2133 3372 2134
rect 3366 2129 3367 2133
rect 3371 2129 3372 2133
rect 3366 2128 3372 2129
rect 3462 2132 3468 2133
rect 3462 2128 3463 2132
rect 3467 2128 3468 2132
rect 1659 2127 1660 2128
rect 1806 2127 1812 2128
rect 3462 2127 3468 2128
rect 1654 2126 1660 2127
rect 134 2121 140 2122
rect 110 2120 116 2121
rect 110 2116 111 2120
rect 115 2116 116 2120
rect 134 2117 135 2121
rect 139 2117 140 2121
rect 134 2116 140 2117
rect 246 2121 252 2122
rect 246 2117 247 2121
rect 251 2117 252 2121
rect 246 2116 252 2117
rect 390 2121 396 2122
rect 390 2117 391 2121
rect 395 2117 396 2121
rect 390 2116 396 2117
rect 542 2121 548 2122
rect 542 2117 543 2121
rect 547 2117 548 2121
rect 542 2116 548 2117
rect 694 2121 700 2122
rect 694 2117 695 2121
rect 699 2117 700 2121
rect 694 2116 700 2117
rect 838 2121 844 2122
rect 838 2117 839 2121
rect 843 2117 844 2121
rect 838 2116 844 2117
rect 974 2121 980 2122
rect 974 2117 975 2121
rect 979 2117 980 2121
rect 974 2116 980 2117
rect 1102 2121 1108 2122
rect 1102 2117 1103 2121
rect 1107 2117 1108 2121
rect 1102 2116 1108 2117
rect 1230 2121 1236 2122
rect 1230 2117 1231 2121
rect 1235 2117 1236 2121
rect 1230 2116 1236 2117
rect 1350 2121 1356 2122
rect 1350 2117 1351 2121
rect 1355 2117 1356 2121
rect 1350 2116 1356 2117
rect 1462 2121 1468 2122
rect 1462 2117 1463 2121
rect 1467 2117 1468 2121
rect 1462 2116 1468 2117
rect 1574 2121 1580 2122
rect 1574 2117 1575 2121
rect 1579 2117 1580 2121
rect 1574 2116 1580 2117
rect 1670 2121 1676 2122
rect 1670 2117 1671 2121
rect 1675 2117 1676 2121
rect 1670 2116 1676 2117
rect 1766 2120 1772 2121
rect 1766 2116 1767 2120
rect 1771 2116 1772 2120
rect 110 2115 116 2116
rect 1766 2115 1772 2116
rect 2886 2115 2892 2116
rect 2886 2111 2887 2115
rect 2891 2114 2892 2115
rect 2975 2115 2981 2116
rect 2975 2114 2976 2115
rect 2891 2112 2976 2114
rect 2891 2111 2892 2112
rect 2886 2110 2892 2111
rect 2975 2111 2976 2112
rect 2980 2111 2981 2115
rect 2975 2110 2981 2111
rect 2998 2115 3004 2116
rect 2998 2111 2999 2115
rect 3003 2114 3004 2115
rect 3063 2115 3069 2116
rect 3063 2114 3064 2115
rect 3003 2112 3064 2114
rect 3003 2111 3004 2112
rect 2998 2110 3004 2111
rect 3063 2111 3064 2112
rect 3068 2111 3069 2115
rect 3063 2110 3069 2111
rect 3086 2115 3092 2116
rect 3086 2111 3087 2115
rect 3091 2114 3092 2115
rect 3151 2115 3157 2116
rect 3151 2114 3152 2115
rect 3091 2112 3152 2114
rect 3091 2111 3092 2112
rect 3086 2110 3092 2111
rect 3151 2111 3152 2112
rect 3156 2111 3157 2115
rect 3151 2110 3157 2111
rect 3239 2115 3245 2116
rect 3239 2111 3240 2115
rect 3244 2114 3245 2115
rect 3255 2115 3261 2116
rect 3255 2114 3256 2115
rect 3244 2112 3256 2114
rect 3244 2111 3245 2112
rect 3239 2110 3245 2111
rect 3255 2111 3256 2112
rect 3260 2111 3261 2115
rect 3255 2110 3261 2111
rect 3327 2115 3333 2116
rect 3327 2111 3328 2115
rect 3332 2114 3333 2115
rect 3358 2115 3364 2116
rect 3358 2114 3359 2115
rect 3332 2112 3359 2114
rect 3332 2111 3333 2112
rect 3327 2110 3333 2111
rect 3358 2111 3359 2112
rect 3363 2111 3364 2115
rect 3358 2110 3364 2111
rect 3415 2115 3421 2116
rect 3415 2111 3416 2115
rect 3420 2114 3421 2115
rect 3438 2115 3444 2116
rect 3438 2114 3439 2115
rect 3420 2112 3439 2114
rect 3420 2111 3421 2112
rect 3415 2110 3421 2111
rect 3438 2111 3439 2112
rect 3443 2111 3444 2115
rect 3438 2110 3444 2111
rect 183 2103 189 2104
rect 183 2099 184 2103
rect 188 2102 189 2103
rect 198 2103 204 2104
rect 198 2102 199 2103
rect 188 2100 199 2102
rect 188 2099 189 2100
rect 183 2098 189 2099
rect 198 2099 199 2100
rect 203 2099 204 2103
rect 198 2098 204 2099
rect 206 2103 212 2104
rect 206 2099 207 2103
rect 211 2102 212 2103
rect 295 2103 301 2104
rect 295 2102 296 2103
rect 211 2100 296 2102
rect 211 2099 212 2100
rect 206 2098 212 2099
rect 295 2099 296 2100
rect 300 2099 301 2103
rect 295 2098 301 2099
rect 318 2103 324 2104
rect 318 2099 319 2103
rect 323 2102 324 2103
rect 439 2103 445 2104
rect 439 2102 440 2103
rect 323 2100 440 2102
rect 323 2099 324 2100
rect 318 2098 324 2099
rect 439 2099 440 2100
rect 444 2099 445 2103
rect 439 2098 445 2099
rect 462 2103 468 2104
rect 462 2099 463 2103
rect 467 2102 468 2103
rect 591 2103 597 2104
rect 591 2102 592 2103
rect 467 2100 592 2102
rect 467 2099 468 2100
rect 462 2098 468 2099
rect 591 2099 592 2100
rect 596 2099 597 2103
rect 591 2098 597 2099
rect 614 2103 620 2104
rect 614 2099 615 2103
rect 619 2102 620 2103
rect 743 2103 749 2104
rect 743 2102 744 2103
rect 619 2100 744 2102
rect 619 2099 620 2100
rect 614 2098 620 2099
rect 743 2099 744 2100
rect 748 2099 749 2103
rect 743 2098 749 2099
rect 887 2103 893 2104
rect 887 2099 888 2103
rect 892 2102 893 2103
rect 927 2103 933 2104
rect 927 2102 928 2103
rect 892 2100 928 2102
rect 892 2099 893 2100
rect 887 2098 893 2099
rect 927 2099 928 2100
rect 932 2099 933 2103
rect 927 2098 933 2099
rect 950 2103 956 2104
rect 950 2099 951 2103
rect 955 2102 956 2103
rect 1023 2103 1029 2104
rect 1023 2102 1024 2103
rect 955 2100 1024 2102
rect 955 2099 956 2100
rect 950 2098 956 2099
rect 1023 2099 1024 2100
rect 1028 2099 1029 2103
rect 1023 2098 1029 2099
rect 1151 2103 1157 2104
rect 1151 2099 1152 2103
rect 1156 2102 1157 2103
rect 1174 2103 1180 2104
rect 1156 2100 1161 2102
rect 1156 2099 1157 2100
rect 1151 2098 1157 2099
rect 622 2095 628 2096
rect 622 2094 623 2095
rect 216 2092 623 2094
rect 183 2087 189 2088
rect 183 2083 184 2087
rect 188 2086 189 2087
rect 216 2086 218 2092
rect 622 2091 623 2092
rect 627 2091 628 2095
rect 1159 2094 1161 2100
rect 1174 2099 1175 2103
rect 1179 2102 1180 2103
rect 1279 2103 1285 2104
rect 1279 2102 1280 2103
rect 1179 2100 1280 2102
rect 1179 2099 1180 2100
rect 1174 2098 1180 2099
rect 1279 2099 1280 2100
rect 1284 2099 1285 2103
rect 1279 2098 1285 2099
rect 1399 2103 1405 2104
rect 1399 2099 1400 2103
rect 1404 2102 1405 2103
rect 1430 2103 1436 2104
rect 1430 2102 1431 2103
rect 1404 2100 1431 2102
rect 1404 2099 1405 2100
rect 1399 2098 1405 2099
rect 1430 2099 1431 2100
rect 1435 2099 1436 2103
rect 1430 2098 1436 2099
rect 1511 2103 1517 2104
rect 1511 2099 1512 2103
rect 1516 2102 1517 2103
rect 1542 2103 1548 2104
rect 1542 2102 1543 2103
rect 1516 2100 1543 2102
rect 1516 2099 1517 2100
rect 1511 2098 1517 2099
rect 1542 2099 1543 2100
rect 1547 2099 1548 2103
rect 1542 2098 1548 2099
rect 1623 2103 1629 2104
rect 1623 2099 1624 2103
rect 1628 2102 1629 2103
rect 1654 2103 1660 2104
rect 1654 2102 1655 2103
rect 1628 2100 1655 2102
rect 1628 2099 1629 2100
rect 1623 2098 1629 2099
rect 1654 2099 1655 2100
rect 1659 2099 1660 2103
rect 1654 2098 1660 2099
rect 1719 2103 1725 2104
rect 1719 2099 1720 2103
rect 1724 2102 1725 2103
rect 1786 2103 1792 2104
rect 1786 2102 1787 2103
rect 1724 2100 1787 2102
rect 1724 2099 1725 2100
rect 1719 2098 1725 2099
rect 1786 2099 1787 2100
rect 1791 2099 1792 2103
rect 3254 2103 3260 2104
rect 3254 2102 3255 2103
rect 1786 2098 1792 2099
rect 3080 2100 3255 2102
rect 1310 2095 1316 2096
rect 1310 2094 1311 2095
rect 1159 2092 1311 2094
rect 622 2090 628 2091
rect 1310 2091 1311 2092
rect 1315 2091 1316 2095
rect 1310 2090 1316 2091
rect 1879 2095 1885 2096
rect 1879 2091 1880 2095
rect 1884 2094 1885 2095
rect 1938 2095 1944 2096
rect 1938 2094 1939 2095
rect 1884 2092 1939 2094
rect 1884 2091 1885 2092
rect 1879 2090 1885 2091
rect 1938 2091 1939 2092
rect 1943 2091 1944 2095
rect 1938 2090 1944 2091
rect 2039 2095 2045 2096
rect 2039 2091 2040 2095
rect 2044 2094 2045 2095
rect 2071 2095 2077 2096
rect 2071 2094 2072 2095
rect 2044 2092 2072 2094
rect 2044 2091 2045 2092
rect 2039 2090 2045 2091
rect 2071 2091 2072 2092
rect 2076 2091 2077 2095
rect 2071 2090 2077 2091
rect 2215 2095 2221 2096
rect 2215 2091 2216 2095
rect 2220 2094 2221 2095
rect 2247 2095 2253 2096
rect 2247 2094 2248 2095
rect 2220 2092 2248 2094
rect 2220 2091 2221 2092
rect 2215 2090 2221 2091
rect 2247 2091 2248 2092
rect 2252 2091 2253 2095
rect 2247 2090 2253 2091
rect 2391 2095 2400 2096
rect 2391 2091 2392 2095
rect 2399 2091 2400 2095
rect 2391 2090 2400 2091
rect 2551 2095 2557 2096
rect 2551 2091 2552 2095
rect 2556 2094 2557 2095
rect 2582 2095 2588 2096
rect 2582 2094 2583 2095
rect 2556 2092 2583 2094
rect 2556 2091 2557 2092
rect 2551 2090 2557 2091
rect 2582 2091 2583 2092
rect 2587 2091 2588 2095
rect 2582 2090 2588 2091
rect 2703 2095 2709 2096
rect 2703 2091 2704 2095
rect 2708 2094 2709 2095
rect 2734 2095 2740 2096
rect 2734 2094 2735 2095
rect 2708 2092 2735 2094
rect 2708 2091 2709 2092
rect 2703 2090 2709 2091
rect 2734 2091 2735 2092
rect 2739 2091 2740 2095
rect 2734 2090 2740 2091
rect 2839 2095 2845 2096
rect 2839 2091 2840 2095
rect 2844 2094 2845 2095
rect 2879 2095 2885 2096
rect 2879 2094 2880 2095
rect 2844 2092 2880 2094
rect 2844 2091 2845 2092
rect 2839 2090 2845 2091
rect 2879 2091 2880 2092
rect 2884 2091 2885 2095
rect 2879 2090 2885 2091
rect 2967 2095 2973 2096
rect 2967 2091 2968 2095
rect 2972 2094 2973 2095
rect 3080 2094 3082 2100
rect 3254 2099 3255 2100
rect 3259 2099 3260 2103
rect 3254 2098 3260 2099
rect 2972 2092 3082 2094
rect 3086 2095 3093 2096
rect 2972 2091 2973 2092
rect 2967 2090 2973 2091
rect 3086 2091 3087 2095
rect 3092 2091 3093 2095
rect 3086 2090 3093 2091
rect 3110 2095 3116 2096
rect 3110 2091 3111 2095
rect 3115 2094 3116 2095
rect 3207 2095 3213 2096
rect 3207 2094 3208 2095
rect 3115 2092 3208 2094
rect 3115 2091 3116 2092
rect 3110 2090 3116 2091
rect 3207 2091 3208 2092
rect 3212 2091 3213 2095
rect 3207 2090 3213 2091
rect 3230 2095 3236 2096
rect 3230 2091 3231 2095
rect 3235 2094 3236 2095
rect 3319 2095 3325 2096
rect 3319 2094 3320 2095
rect 3235 2092 3320 2094
rect 3235 2091 3236 2092
rect 3230 2090 3236 2091
rect 3319 2091 3320 2092
rect 3324 2091 3325 2095
rect 3319 2090 3325 2091
rect 3350 2095 3356 2096
rect 3350 2091 3351 2095
rect 3355 2094 3356 2095
rect 3415 2095 3421 2096
rect 3415 2094 3416 2095
rect 3355 2092 3416 2094
rect 3355 2091 3356 2092
rect 3350 2090 3356 2091
rect 3415 2091 3416 2092
rect 3420 2091 3421 2095
rect 3415 2090 3421 2091
rect 271 2087 277 2088
rect 271 2086 272 2087
rect 188 2084 218 2086
rect 220 2084 272 2086
rect 188 2083 189 2084
rect 183 2082 189 2083
rect 220 2078 222 2084
rect 271 2083 272 2084
rect 276 2083 277 2087
rect 271 2082 277 2083
rect 294 2087 300 2088
rect 294 2083 295 2087
rect 299 2086 300 2087
rect 391 2087 397 2088
rect 391 2086 392 2087
rect 299 2084 392 2086
rect 299 2083 300 2084
rect 294 2082 300 2083
rect 391 2083 392 2084
rect 396 2083 397 2087
rect 391 2082 397 2083
rect 414 2087 420 2088
rect 414 2083 415 2087
rect 419 2086 420 2087
rect 511 2087 517 2088
rect 511 2086 512 2087
rect 419 2084 512 2086
rect 419 2083 420 2084
rect 414 2082 420 2083
rect 511 2083 512 2084
rect 516 2083 517 2087
rect 511 2082 517 2083
rect 534 2087 540 2088
rect 534 2083 535 2087
rect 539 2086 540 2087
rect 631 2087 637 2088
rect 631 2086 632 2087
rect 539 2084 632 2086
rect 539 2083 540 2084
rect 534 2082 540 2083
rect 631 2083 632 2084
rect 636 2083 637 2087
rect 631 2082 637 2083
rect 751 2087 760 2088
rect 751 2083 752 2087
rect 759 2083 760 2087
rect 751 2082 760 2083
rect 774 2087 780 2088
rect 774 2083 775 2087
rect 779 2086 780 2087
rect 871 2087 877 2088
rect 871 2086 872 2087
rect 779 2084 872 2086
rect 779 2083 780 2084
rect 774 2082 780 2083
rect 871 2083 872 2084
rect 876 2083 877 2087
rect 871 2082 877 2083
rect 894 2087 900 2088
rect 894 2083 895 2087
rect 899 2086 900 2087
rect 983 2087 989 2088
rect 983 2086 984 2087
rect 899 2084 984 2086
rect 899 2083 900 2084
rect 894 2082 900 2083
rect 983 2083 984 2084
rect 988 2083 989 2087
rect 983 2082 989 2083
rect 1054 2087 1060 2088
rect 1054 2083 1055 2087
rect 1059 2086 1060 2087
rect 1095 2087 1101 2088
rect 1095 2086 1096 2087
rect 1059 2084 1096 2086
rect 1059 2083 1060 2084
rect 1054 2082 1060 2083
rect 1095 2083 1096 2084
rect 1100 2083 1101 2087
rect 1095 2082 1101 2083
rect 1118 2087 1124 2088
rect 1118 2083 1119 2087
rect 1123 2086 1124 2087
rect 1207 2087 1213 2088
rect 1207 2086 1208 2087
rect 1123 2084 1208 2086
rect 1123 2083 1124 2084
rect 1118 2082 1124 2083
rect 1207 2083 1208 2084
rect 1212 2083 1213 2087
rect 1207 2082 1213 2083
rect 1258 2087 1264 2088
rect 1258 2083 1259 2087
rect 1263 2086 1264 2087
rect 1327 2087 1333 2088
rect 1327 2086 1328 2087
rect 1263 2084 1328 2086
rect 1263 2083 1264 2084
rect 1258 2082 1264 2083
rect 1327 2083 1328 2084
rect 1332 2083 1333 2087
rect 1327 2082 1333 2083
rect 208 2076 222 2078
rect 1806 2080 1812 2081
rect 3462 2080 3468 2081
rect 1806 2076 1807 2080
rect 1811 2076 1812 2080
rect 110 2072 116 2073
rect 110 2068 111 2072
rect 115 2068 116 2072
rect 110 2067 116 2068
rect 134 2071 140 2072
rect 134 2067 135 2071
rect 139 2067 140 2071
rect 134 2066 140 2067
rect 208 2061 210 2076
rect 1806 2075 1812 2076
rect 1830 2079 1836 2080
rect 1830 2075 1831 2079
rect 1835 2075 1836 2079
rect 1830 2074 1836 2075
rect 1990 2079 1996 2080
rect 1990 2075 1991 2079
rect 1995 2075 1996 2079
rect 1990 2074 1996 2075
rect 2166 2079 2172 2080
rect 2166 2075 2167 2079
rect 2171 2075 2172 2079
rect 2166 2074 2172 2075
rect 2342 2079 2348 2080
rect 2342 2075 2343 2079
rect 2347 2075 2348 2079
rect 2342 2074 2348 2075
rect 2502 2079 2508 2080
rect 2502 2075 2503 2079
rect 2507 2075 2508 2079
rect 2502 2074 2508 2075
rect 2654 2079 2660 2080
rect 2654 2075 2655 2079
rect 2659 2075 2660 2079
rect 2654 2074 2660 2075
rect 2790 2079 2796 2080
rect 2790 2075 2791 2079
rect 2795 2075 2796 2079
rect 2790 2074 2796 2075
rect 2918 2079 2924 2080
rect 2918 2075 2919 2079
rect 2923 2075 2924 2079
rect 2918 2074 2924 2075
rect 3038 2079 3044 2080
rect 3038 2075 3039 2079
rect 3043 2075 3044 2079
rect 3038 2074 3044 2075
rect 3158 2079 3164 2080
rect 3158 2075 3159 2079
rect 3163 2075 3164 2079
rect 3158 2074 3164 2075
rect 3270 2079 3276 2080
rect 3270 2075 3271 2079
rect 3275 2075 3276 2079
rect 3270 2074 3276 2075
rect 3366 2079 3372 2080
rect 3366 2075 3367 2079
rect 3371 2075 3372 2079
rect 3462 2076 3463 2080
rect 3467 2076 3468 2080
rect 3462 2075 3468 2076
rect 3366 2074 3372 2075
rect 1766 2072 1772 2073
rect 222 2071 228 2072
rect 222 2067 223 2071
rect 227 2067 228 2071
rect 222 2066 228 2067
rect 342 2071 348 2072
rect 342 2067 343 2071
rect 347 2067 348 2071
rect 342 2066 348 2067
rect 462 2071 468 2072
rect 462 2067 463 2071
rect 467 2067 468 2071
rect 462 2066 468 2067
rect 582 2071 588 2072
rect 582 2067 583 2071
rect 587 2067 588 2071
rect 582 2066 588 2067
rect 702 2071 708 2072
rect 702 2067 703 2071
rect 707 2067 708 2071
rect 702 2066 708 2067
rect 822 2071 828 2072
rect 822 2067 823 2071
rect 827 2067 828 2071
rect 822 2066 828 2067
rect 934 2071 940 2072
rect 934 2067 935 2071
rect 939 2067 940 2071
rect 934 2066 940 2067
rect 1046 2071 1052 2072
rect 1046 2067 1047 2071
rect 1051 2067 1052 2071
rect 1046 2066 1052 2067
rect 1158 2071 1164 2072
rect 1158 2067 1159 2071
rect 1163 2067 1164 2071
rect 1158 2066 1164 2067
rect 1278 2071 1284 2072
rect 1278 2067 1279 2071
rect 1283 2067 1284 2071
rect 1766 2068 1767 2072
rect 1771 2068 1772 2072
rect 1766 2067 1772 2068
rect 1786 2071 1792 2072
rect 1786 2067 1787 2071
rect 1791 2070 1792 2071
rect 1938 2071 1944 2072
rect 1791 2068 1873 2070
rect 1791 2067 1792 2068
rect 1278 2066 1284 2067
rect 1786 2066 1792 2067
rect 1938 2067 1939 2071
rect 1943 2070 1944 2071
rect 2071 2071 2077 2072
rect 1943 2068 2033 2070
rect 1943 2067 1944 2068
rect 1938 2066 1944 2067
rect 2071 2067 2072 2071
rect 2076 2070 2077 2071
rect 2247 2071 2253 2072
rect 2076 2068 2209 2070
rect 2076 2067 2077 2068
rect 2071 2066 2077 2067
rect 2247 2067 2248 2071
rect 2252 2070 2253 2071
rect 2582 2071 2588 2072
rect 2252 2068 2385 2070
rect 2252 2067 2253 2068
rect 2247 2066 2253 2067
rect 2574 2067 2580 2068
rect 294 2063 300 2064
rect 294 2059 295 2063
rect 299 2059 300 2063
rect 294 2058 300 2059
rect 414 2063 420 2064
rect 414 2059 415 2063
rect 419 2059 420 2063
rect 414 2058 420 2059
rect 534 2063 540 2064
rect 534 2059 535 2063
rect 539 2059 540 2063
rect 534 2058 540 2059
rect 542 2063 548 2064
rect 542 2059 543 2063
rect 547 2062 548 2063
rect 774 2063 780 2064
rect 547 2060 625 2062
rect 547 2059 548 2060
rect 542 2058 548 2059
rect 774 2059 775 2063
rect 779 2059 780 2063
rect 774 2058 780 2059
rect 894 2063 900 2064
rect 894 2059 895 2063
rect 899 2059 900 2063
rect 894 2058 900 2059
rect 927 2063 933 2064
rect 927 2059 928 2063
rect 932 2062 933 2063
rect 1118 2063 1124 2064
rect 932 2060 977 2062
rect 932 2059 933 2060
rect 927 2058 933 2059
rect 1118 2059 1119 2063
rect 1123 2059 1124 2063
rect 1258 2063 1264 2064
rect 1258 2062 1259 2063
rect 1233 2060 1259 2062
rect 1118 2058 1124 2059
rect 1258 2059 1259 2060
rect 1263 2059 1264 2063
rect 1258 2058 1264 2059
rect 1270 2063 1276 2064
rect 1270 2059 1271 2063
rect 1275 2062 1276 2063
rect 1806 2063 1812 2064
rect 1275 2060 1321 2062
rect 1275 2059 1276 2060
rect 1270 2058 1276 2059
rect 1806 2059 1807 2063
rect 1811 2059 1812 2063
rect 2574 2063 2575 2067
rect 2579 2063 2580 2067
rect 2582 2067 2583 2071
rect 2587 2070 2588 2071
rect 2734 2071 2740 2072
rect 2587 2068 2697 2070
rect 2587 2067 2588 2068
rect 2582 2066 2588 2067
rect 2734 2067 2735 2071
rect 2739 2070 2740 2071
rect 2879 2071 2885 2072
rect 2739 2068 2833 2070
rect 2739 2067 2740 2068
rect 2734 2066 2740 2067
rect 2879 2067 2880 2071
rect 2884 2070 2885 2071
rect 3110 2071 3116 2072
rect 2884 2068 2961 2070
rect 2884 2067 2885 2068
rect 2879 2066 2885 2067
rect 3110 2067 3111 2071
rect 3115 2067 3116 2071
rect 3110 2066 3116 2067
rect 3230 2071 3236 2072
rect 3230 2067 3231 2071
rect 3235 2067 3236 2071
rect 3230 2066 3236 2067
rect 3255 2071 3261 2072
rect 3255 2067 3256 2071
rect 3260 2070 3261 2071
rect 3260 2068 3313 2070
rect 3260 2067 3261 2068
rect 3255 2066 3261 2067
rect 3438 2067 3444 2068
rect 2574 2062 2580 2063
rect 3438 2063 3439 2067
rect 3443 2063 3444 2067
rect 3438 2062 3444 2063
rect 3462 2063 3468 2064
rect 1806 2058 1812 2059
rect 1830 2060 1836 2061
rect 1830 2056 1831 2060
rect 1835 2056 1836 2060
rect 110 2055 116 2056
rect 110 2051 111 2055
rect 115 2051 116 2055
rect 1766 2055 1772 2056
rect 1830 2055 1836 2056
rect 1990 2060 1996 2061
rect 1990 2056 1991 2060
rect 1995 2056 1996 2060
rect 1990 2055 1996 2056
rect 2166 2060 2172 2061
rect 2166 2056 2167 2060
rect 2171 2056 2172 2060
rect 2166 2055 2172 2056
rect 2342 2060 2348 2061
rect 2342 2056 2343 2060
rect 2347 2056 2348 2060
rect 2342 2055 2348 2056
rect 2502 2060 2508 2061
rect 2502 2056 2503 2060
rect 2507 2056 2508 2060
rect 2502 2055 2508 2056
rect 2654 2060 2660 2061
rect 2654 2056 2655 2060
rect 2659 2056 2660 2060
rect 2654 2055 2660 2056
rect 2790 2060 2796 2061
rect 2790 2056 2791 2060
rect 2795 2056 2796 2060
rect 2790 2055 2796 2056
rect 2918 2060 2924 2061
rect 2918 2056 2919 2060
rect 2923 2056 2924 2060
rect 2918 2055 2924 2056
rect 3038 2060 3044 2061
rect 3038 2056 3039 2060
rect 3043 2056 3044 2060
rect 3038 2055 3044 2056
rect 3158 2060 3164 2061
rect 3158 2056 3159 2060
rect 3163 2056 3164 2060
rect 3158 2055 3164 2056
rect 3270 2060 3276 2061
rect 3270 2056 3271 2060
rect 3275 2056 3276 2060
rect 3270 2055 3276 2056
rect 3366 2060 3372 2061
rect 3366 2056 3367 2060
rect 3371 2056 3372 2060
rect 3462 2059 3463 2063
rect 3467 2059 3468 2063
rect 3462 2058 3468 2059
rect 3366 2055 3372 2056
rect 110 2050 116 2051
rect 134 2052 140 2053
rect 134 2048 135 2052
rect 139 2048 140 2052
rect 134 2047 140 2048
rect 222 2052 228 2053
rect 222 2048 223 2052
rect 227 2048 228 2052
rect 222 2047 228 2048
rect 342 2052 348 2053
rect 342 2048 343 2052
rect 347 2048 348 2052
rect 342 2047 348 2048
rect 462 2052 468 2053
rect 462 2048 463 2052
rect 467 2048 468 2052
rect 462 2047 468 2048
rect 582 2052 588 2053
rect 582 2048 583 2052
rect 587 2048 588 2052
rect 582 2047 588 2048
rect 702 2052 708 2053
rect 702 2048 703 2052
rect 707 2048 708 2052
rect 702 2047 708 2048
rect 822 2052 828 2053
rect 822 2048 823 2052
rect 827 2048 828 2052
rect 822 2047 828 2048
rect 934 2052 940 2053
rect 934 2048 935 2052
rect 939 2048 940 2052
rect 934 2047 940 2048
rect 1046 2052 1052 2053
rect 1046 2048 1047 2052
rect 1051 2048 1052 2052
rect 1046 2047 1052 2048
rect 1158 2052 1164 2053
rect 1158 2048 1159 2052
rect 1163 2048 1164 2052
rect 1158 2047 1164 2048
rect 1278 2052 1284 2053
rect 1278 2048 1279 2052
rect 1283 2048 1284 2052
rect 1766 2051 1767 2055
rect 1771 2051 1772 2055
rect 1766 2050 1772 2051
rect 1278 2047 1284 2048
rect 186 2015 192 2016
rect 186 2011 187 2015
rect 191 2014 192 2015
rect 542 2015 548 2016
rect 542 2014 543 2015
rect 191 2012 543 2014
rect 191 2011 192 2012
rect 186 2010 192 2011
rect 542 2011 543 2012
rect 547 2011 548 2015
rect 542 2010 548 2011
rect 1830 2012 1836 2013
rect 1806 2009 1812 2010
rect 1806 2005 1807 2009
rect 1811 2005 1812 2009
rect 1830 2008 1831 2012
rect 1835 2008 1836 2012
rect 1830 2007 1836 2008
rect 2014 2012 2020 2013
rect 2014 2008 2015 2012
rect 2019 2008 2020 2012
rect 2014 2007 2020 2008
rect 2222 2012 2228 2013
rect 2222 2008 2223 2012
rect 2227 2008 2228 2012
rect 2222 2007 2228 2008
rect 2430 2012 2436 2013
rect 2430 2008 2431 2012
rect 2435 2008 2436 2012
rect 2430 2007 2436 2008
rect 2630 2012 2636 2013
rect 2630 2008 2631 2012
rect 2635 2008 2636 2012
rect 2630 2007 2636 2008
rect 2822 2012 2828 2013
rect 2822 2008 2823 2012
rect 2827 2008 2828 2012
rect 2822 2007 2828 2008
rect 3006 2012 3012 2013
rect 3006 2008 3007 2012
rect 3011 2008 3012 2012
rect 3006 2007 3012 2008
rect 3198 2012 3204 2013
rect 3198 2008 3199 2012
rect 3203 2008 3204 2012
rect 3198 2007 3204 2008
rect 3366 2012 3372 2013
rect 3366 2008 3367 2012
rect 3371 2008 3372 2012
rect 3366 2007 3372 2008
rect 3462 2009 3468 2010
rect 1806 2004 1812 2005
rect 3462 2005 3463 2009
rect 3467 2005 3468 2009
rect 3462 2004 3468 2005
rect 1966 2003 1972 2004
rect 1966 2002 1967 2003
rect 134 2000 140 2001
rect 110 1997 116 1998
rect 110 1993 111 1997
rect 115 1993 116 1997
rect 134 1996 135 2000
rect 139 1996 140 2000
rect 134 1995 140 1996
rect 238 2000 244 2001
rect 238 1996 239 2000
rect 243 1996 244 2000
rect 238 1995 244 1996
rect 366 2000 372 2001
rect 366 1996 367 2000
rect 371 1996 372 2000
rect 366 1995 372 1996
rect 502 2000 508 2001
rect 502 1996 503 2000
rect 507 1996 508 2000
rect 502 1995 508 1996
rect 638 2000 644 2001
rect 638 1996 639 2000
rect 643 1996 644 2000
rect 638 1995 644 1996
rect 774 2000 780 2001
rect 774 1996 775 2000
rect 779 1996 780 2000
rect 774 1995 780 1996
rect 910 2000 916 2001
rect 910 1996 911 2000
rect 915 1996 916 2000
rect 910 1995 916 1996
rect 1046 2000 1052 2001
rect 1046 1996 1047 2000
rect 1051 1996 1052 2000
rect 1046 1995 1052 1996
rect 1182 2000 1188 2001
rect 1182 1996 1183 2000
rect 1187 1996 1188 2000
rect 1182 1995 1188 1996
rect 1326 2000 1332 2001
rect 1905 2000 1967 2002
rect 1326 1996 1327 2000
rect 1331 1996 1332 2000
rect 1966 1999 1967 2000
rect 1971 1999 1972 2003
rect 1966 1998 1972 1999
rect 2086 2003 2092 2004
rect 2086 1999 2087 2003
rect 2091 1999 2092 2003
rect 2086 1998 2092 1999
rect 2294 2003 2300 2004
rect 2294 1999 2295 2003
rect 2299 1999 2300 2003
rect 2294 1998 2300 1999
rect 2394 2003 2400 2004
rect 2394 1999 2395 2003
rect 2399 2002 2400 2003
rect 2702 2003 2708 2004
rect 2399 2000 2473 2002
rect 2399 1999 2400 2000
rect 2394 1998 2400 1999
rect 2702 1999 2703 2003
rect 2707 1999 2708 2003
rect 2702 1998 2708 1999
rect 2894 2003 2900 2004
rect 2894 1999 2895 2003
rect 2899 1999 2900 2003
rect 2894 1998 2900 1999
rect 2998 2003 3004 2004
rect 2998 1999 2999 2003
rect 3003 2002 3004 2003
rect 3086 2003 3092 2004
rect 3003 2000 3049 2002
rect 3003 1999 3004 2000
rect 2998 1998 3004 1999
rect 3086 1999 3087 2003
rect 3091 2002 3092 2003
rect 3430 2003 3436 2004
rect 3091 2000 3241 2002
rect 3091 1999 3092 2000
rect 3086 1998 3092 1999
rect 3430 1999 3431 2003
rect 3435 1999 3436 2003
rect 3430 1998 3436 1999
rect 1326 1995 1332 1996
rect 1766 1997 1772 1998
rect 110 1992 116 1993
rect 1766 1993 1767 1997
rect 1771 1993 1772 1997
rect 1830 1993 1836 1994
rect 1766 1992 1772 1993
rect 1806 1992 1812 1993
rect 206 1991 212 1992
rect 206 1987 207 1991
rect 211 1987 212 1991
rect 206 1986 212 1987
rect 310 1991 316 1992
rect 310 1987 311 1991
rect 315 1987 316 1991
rect 310 1986 316 1987
rect 438 1991 444 1992
rect 438 1987 439 1991
rect 443 1987 444 1991
rect 438 1986 444 1987
rect 574 1991 580 1992
rect 574 1987 575 1991
rect 579 1987 580 1991
rect 574 1986 580 1987
rect 582 1991 588 1992
rect 582 1987 583 1991
rect 587 1990 588 1991
rect 754 1991 760 1992
rect 587 1988 681 1990
rect 587 1987 588 1988
rect 582 1986 588 1987
rect 754 1987 755 1991
rect 759 1990 760 1991
rect 854 1991 860 1992
rect 759 1988 817 1990
rect 759 1987 760 1988
rect 754 1986 760 1987
rect 854 1987 855 1991
rect 859 1990 860 1991
rect 1134 1991 1140 1992
rect 1134 1990 1135 1991
rect 859 1988 953 1990
rect 1121 1988 1135 1990
rect 859 1987 860 1988
rect 854 1986 860 1987
rect 1134 1987 1135 1988
rect 1139 1987 1140 1991
rect 1134 1986 1140 1987
rect 1254 1991 1260 1992
rect 1254 1987 1255 1991
rect 1259 1987 1260 1991
rect 1254 1986 1260 1987
rect 1398 1991 1404 1992
rect 1398 1987 1399 1991
rect 1403 1987 1404 1991
rect 1806 1988 1807 1992
rect 1811 1988 1812 1992
rect 1830 1989 1831 1993
rect 1835 1989 1836 1993
rect 1830 1988 1836 1989
rect 2014 1993 2020 1994
rect 2014 1989 2015 1993
rect 2019 1989 2020 1993
rect 2014 1988 2020 1989
rect 2222 1993 2228 1994
rect 2222 1989 2223 1993
rect 2227 1989 2228 1993
rect 2222 1988 2228 1989
rect 2430 1993 2436 1994
rect 2430 1989 2431 1993
rect 2435 1989 2436 1993
rect 2430 1988 2436 1989
rect 2630 1993 2636 1994
rect 2630 1989 2631 1993
rect 2635 1989 2636 1993
rect 2630 1988 2636 1989
rect 2822 1993 2828 1994
rect 2822 1989 2823 1993
rect 2827 1989 2828 1993
rect 2822 1988 2828 1989
rect 3006 1993 3012 1994
rect 3006 1989 3007 1993
rect 3011 1989 3012 1993
rect 3006 1988 3012 1989
rect 3198 1993 3204 1994
rect 3198 1989 3199 1993
rect 3203 1989 3204 1993
rect 3198 1988 3204 1989
rect 3366 1993 3372 1994
rect 3366 1989 3367 1993
rect 3371 1989 3372 1993
rect 3366 1988 3372 1989
rect 3462 1992 3468 1993
rect 3462 1988 3463 1992
rect 3467 1988 3468 1992
rect 1806 1987 1812 1988
rect 3462 1987 3468 1988
rect 1398 1986 1404 1987
rect 134 1981 140 1982
rect 110 1980 116 1981
rect 110 1976 111 1980
rect 115 1976 116 1980
rect 134 1977 135 1981
rect 139 1977 140 1981
rect 134 1976 140 1977
rect 238 1981 244 1982
rect 238 1977 239 1981
rect 243 1977 244 1981
rect 238 1976 244 1977
rect 366 1981 372 1982
rect 366 1977 367 1981
rect 371 1977 372 1981
rect 366 1976 372 1977
rect 502 1981 508 1982
rect 502 1977 503 1981
rect 507 1977 508 1981
rect 502 1976 508 1977
rect 638 1981 644 1982
rect 638 1977 639 1981
rect 643 1977 644 1981
rect 638 1976 644 1977
rect 774 1981 780 1982
rect 774 1977 775 1981
rect 779 1977 780 1981
rect 774 1976 780 1977
rect 910 1981 916 1982
rect 910 1977 911 1981
rect 915 1977 916 1981
rect 910 1976 916 1977
rect 1046 1981 1052 1982
rect 1046 1977 1047 1981
rect 1051 1977 1052 1981
rect 1046 1976 1052 1977
rect 1182 1981 1188 1982
rect 1182 1977 1183 1981
rect 1187 1977 1188 1981
rect 1182 1976 1188 1977
rect 1326 1981 1332 1982
rect 1326 1977 1327 1981
rect 1331 1977 1332 1981
rect 1326 1976 1332 1977
rect 1766 1980 1772 1981
rect 1766 1976 1767 1980
rect 1771 1976 1772 1980
rect 110 1975 116 1976
rect 1766 1975 1772 1976
rect 1879 1975 1885 1976
rect 1879 1971 1880 1975
rect 1884 1974 1885 1975
rect 1934 1975 1940 1976
rect 1934 1974 1935 1975
rect 1884 1972 1935 1974
rect 1884 1971 1885 1972
rect 1879 1970 1885 1971
rect 1934 1971 1935 1972
rect 1939 1971 1940 1975
rect 1934 1970 1940 1971
rect 1966 1975 1972 1976
rect 1966 1971 1967 1975
rect 1971 1974 1972 1975
rect 2063 1975 2069 1976
rect 2063 1974 2064 1975
rect 1971 1972 2064 1974
rect 1971 1971 1972 1972
rect 1966 1970 1972 1971
rect 2063 1971 2064 1972
rect 2068 1971 2069 1975
rect 2063 1970 2069 1971
rect 2086 1975 2092 1976
rect 2086 1971 2087 1975
rect 2091 1974 2092 1975
rect 2271 1975 2277 1976
rect 2271 1974 2272 1975
rect 2091 1972 2272 1974
rect 2091 1971 2092 1972
rect 2086 1970 2092 1971
rect 2271 1971 2272 1972
rect 2276 1971 2277 1975
rect 2271 1970 2277 1971
rect 2294 1975 2300 1976
rect 2294 1971 2295 1975
rect 2299 1974 2300 1975
rect 2479 1975 2485 1976
rect 2479 1974 2480 1975
rect 2299 1972 2480 1974
rect 2299 1971 2300 1972
rect 2294 1970 2300 1971
rect 2479 1971 2480 1972
rect 2484 1971 2485 1975
rect 2479 1970 2485 1971
rect 2574 1975 2580 1976
rect 2574 1971 2575 1975
rect 2579 1974 2580 1975
rect 2679 1975 2685 1976
rect 2679 1974 2680 1975
rect 2579 1972 2680 1974
rect 2579 1971 2580 1972
rect 2574 1970 2580 1971
rect 2679 1971 2680 1972
rect 2684 1971 2685 1975
rect 2679 1970 2685 1971
rect 2702 1975 2708 1976
rect 2702 1971 2703 1975
rect 2707 1974 2708 1975
rect 2871 1975 2877 1976
rect 2871 1974 2872 1975
rect 2707 1972 2872 1974
rect 2707 1971 2708 1972
rect 2702 1970 2708 1971
rect 2871 1971 2872 1972
rect 2876 1971 2877 1975
rect 2871 1970 2877 1971
rect 2894 1975 2900 1976
rect 2894 1971 2895 1975
rect 2899 1974 2900 1975
rect 3055 1975 3061 1976
rect 3055 1974 3056 1975
rect 2899 1972 3056 1974
rect 2899 1971 2900 1972
rect 2894 1970 2900 1971
rect 3055 1971 3056 1972
rect 3060 1971 3061 1975
rect 3055 1970 3061 1971
rect 3238 1975 3244 1976
rect 3238 1971 3239 1975
rect 3243 1974 3244 1975
rect 3247 1975 3253 1976
rect 3247 1974 3248 1975
rect 3243 1972 3248 1974
rect 3243 1971 3244 1972
rect 3238 1970 3244 1971
rect 3247 1971 3248 1972
rect 3252 1971 3253 1975
rect 3247 1970 3253 1971
rect 3415 1975 3421 1976
rect 3415 1971 3416 1975
rect 3420 1974 3421 1975
rect 3438 1975 3444 1976
rect 3438 1974 3439 1975
rect 3420 1972 3439 1974
rect 3420 1971 3421 1972
rect 3415 1970 3421 1971
rect 3438 1971 3439 1972
rect 3443 1971 3444 1975
rect 3438 1970 3444 1971
rect 2366 1967 2372 1968
rect 2366 1966 2367 1967
rect 2292 1964 2367 1966
rect 183 1963 192 1964
rect 183 1959 184 1963
rect 191 1959 192 1963
rect 183 1958 192 1959
rect 206 1963 212 1964
rect 206 1959 207 1963
rect 211 1962 212 1963
rect 287 1963 293 1964
rect 287 1962 288 1963
rect 211 1960 288 1962
rect 211 1959 212 1960
rect 206 1958 212 1959
rect 287 1959 288 1960
rect 292 1959 293 1963
rect 287 1958 293 1959
rect 310 1963 316 1964
rect 310 1959 311 1963
rect 315 1962 316 1963
rect 415 1963 421 1964
rect 415 1962 416 1963
rect 315 1960 416 1962
rect 315 1959 316 1960
rect 310 1958 316 1959
rect 415 1959 416 1960
rect 420 1959 421 1963
rect 415 1958 421 1959
rect 438 1963 444 1964
rect 438 1959 439 1963
rect 443 1962 444 1963
rect 551 1963 557 1964
rect 551 1962 552 1963
rect 443 1960 552 1962
rect 443 1959 444 1960
rect 438 1958 444 1959
rect 551 1959 552 1960
rect 556 1959 557 1963
rect 551 1958 557 1959
rect 574 1963 580 1964
rect 574 1959 575 1963
rect 579 1962 580 1963
rect 687 1963 693 1964
rect 687 1962 688 1963
rect 579 1960 688 1962
rect 579 1959 580 1960
rect 574 1958 580 1959
rect 687 1959 688 1960
rect 692 1959 693 1963
rect 687 1958 693 1959
rect 823 1963 829 1964
rect 823 1959 824 1963
rect 828 1962 829 1963
rect 854 1963 860 1964
rect 854 1962 855 1963
rect 828 1960 855 1962
rect 828 1959 829 1960
rect 823 1958 829 1959
rect 854 1959 855 1960
rect 859 1959 860 1963
rect 854 1958 860 1959
rect 959 1963 968 1964
rect 959 1959 960 1963
rect 967 1959 968 1963
rect 959 1958 968 1959
rect 1095 1963 1101 1964
rect 1095 1959 1096 1963
rect 1100 1962 1101 1963
rect 1134 1963 1140 1964
rect 1100 1960 1130 1962
rect 1100 1959 1101 1960
rect 1095 1958 1101 1959
rect 582 1955 588 1956
rect 582 1954 583 1955
rect 396 1952 583 1954
rect 343 1947 349 1948
rect 343 1943 344 1947
rect 348 1946 349 1947
rect 396 1946 398 1952
rect 582 1951 583 1952
rect 587 1951 588 1955
rect 1128 1954 1130 1960
rect 1134 1959 1135 1963
rect 1139 1962 1140 1963
rect 1231 1963 1237 1964
rect 1231 1962 1232 1963
rect 1139 1960 1232 1962
rect 1139 1959 1140 1960
rect 1134 1958 1140 1959
rect 1231 1959 1232 1960
rect 1236 1959 1237 1963
rect 1231 1958 1237 1959
rect 1254 1963 1260 1964
rect 1254 1959 1255 1963
rect 1259 1962 1260 1963
rect 1375 1963 1381 1964
rect 1375 1962 1376 1963
rect 1259 1960 1376 1962
rect 1259 1959 1260 1960
rect 1254 1958 1260 1959
rect 1375 1959 1376 1960
rect 1380 1959 1381 1963
rect 1375 1958 1381 1959
rect 1911 1959 1917 1960
rect 1270 1955 1276 1956
rect 1270 1954 1271 1955
rect 1128 1952 1271 1954
rect 582 1950 588 1951
rect 1270 1951 1271 1952
rect 1275 1951 1276 1955
rect 1911 1955 1912 1959
rect 1916 1958 1917 1959
rect 1951 1959 1957 1960
rect 1951 1958 1952 1959
rect 1916 1956 1952 1958
rect 1916 1955 1917 1956
rect 1911 1954 1917 1955
rect 1951 1955 1952 1956
rect 1956 1955 1957 1959
rect 1951 1954 1957 1955
rect 2047 1959 2053 1960
rect 2047 1955 2048 1959
rect 2052 1958 2053 1959
rect 2078 1959 2084 1960
rect 2078 1958 2079 1959
rect 2052 1956 2079 1958
rect 2052 1955 2053 1956
rect 2047 1954 2053 1955
rect 2078 1955 2079 1956
rect 2083 1955 2084 1959
rect 2078 1954 2084 1955
rect 2191 1959 2197 1960
rect 2191 1955 2192 1959
rect 2196 1958 2197 1959
rect 2292 1958 2294 1964
rect 2366 1963 2367 1964
rect 2371 1963 2372 1967
rect 3246 1967 3252 1968
rect 3246 1966 3247 1967
rect 2366 1962 2372 1963
rect 3128 1964 3247 1966
rect 2196 1956 2294 1958
rect 2298 1959 2304 1960
rect 2196 1955 2197 1956
rect 2191 1954 2197 1955
rect 2298 1955 2299 1959
rect 2303 1958 2304 1959
rect 2335 1959 2341 1960
rect 2335 1958 2336 1959
rect 2303 1956 2336 1958
rect 2303 1955 2304 1956
rect 2298 1954 2304 1955
rect 2335 1955 2336 1956
rect 2340 1955 2341 1959
rect 2335 1954 2341 1955
rect 2358 1959 2364 1960
rect 2358 1955 2359 1959
rect 2363 1958 2364 1959
rect 2479 1959 2485 1960
rect 2479 1958 2480 1959
rect 2363 1956 2480 1958
rect 2363 1955 2364 1956
rect 2358 1954 2364 1955
rect 2479 1955 2480 1956
rect 2484 1955 2485 1959
rect 2479 1954 2485 1955
rect 2623 1959 2629 1960
rect 2623 1955 2624 1959
rect 2628 1958 2629 1959
rect 2654 1959 2660 1960
rect 2654 1958 2655 1959
rect 2628 1956 2655 1958
rect 2628 1955 2629 1956
rect 2623 1954 2629 1955
rect 2654 1955 2655 1956
rect 2659 1955 2660 1959
rect 2654 1954 2660 1955
rect 2759 1959 2765 1960
rect 2759 1955 2760 1959
rect 2764 1958 2765 1959
rect 2798 1959 2804 1960
rect 2798 1958 2799 1959
rect 2764 1956 2799 1958
rect 2764 1955 2765 1956
rect 2759 1954 2765 1955
rect 2798 1955 2799 1956
rect 2803 1955 2804 1959
rect 2798 1954 2804 1955
rect 2879 1959 2885 1960
rect 2879 1955 2880 1959
rect 2884 1958 2885 1959
rect 2910 1959 2916 1960
rect 2910 1958 2911 1959
rect 2884 1956 2911 1958
rect 2884 1955 2885 1956
rect 2879 1954 2885 1955
rect 2910 1955 2911 1956
rect 2915 1955 2916 1959
rect 2910 1954 2916 1955
rect 2998 1959 3005 1960
rect 2998 1955 2999 1959
rect 3004 1955 3005 1959
rect 2998 1954 3005 1955
rect 3111 1959 3117 1960
rect 3111 1955 3112 1959
rect 3116 1958 3117 1959
rect 3128 1958 3130 1964
rect 3246 1963 3247 1964
rect 3251 1963 3252 1967
rect 3246 1962 3252 1963
rect 3116 1956 3130 1958
rect 3134 1959 3140 1960
rect 3116 1955 3117 1956
rect 3111 1954 3117 1955
rect 3134 1955 3135 1959
rect 3139 1958 3140 1959
rect 3215 1959 3221 1960
rect 3215 1958 3216 1959
rect 3139 1956 3216 1958
rect 3139 1955 3140 1956
rect 3134 1954 3140 1955
rect 3215 1955 3216 1956
rect 3220 1955 3221 1959
rect 3215 1954 3221 1955
rect 3327 1959 3333 1960
rect 3327 1955 3328 1959
rect 3332 1958 3333 1959
rect 3358 1959 3364 1960
rect 3358 1958 3359 1959
rect 3332 1956 3359 1958
rect 3332 1955 3333 1956
rect 3327 1954 3333 1955
rect 3358 1955 3359 1956
rect 3363 1955 3364 1959
rect 3358 1954 3364 1955
rect 3415 1959 3421 1960
rect 3415 1955 3416 1959
rect 3420 1958 3421 1959
rect 3430 1959 3436 1960
rect 3430 1958 3431 1959
rect 3420 1956 3431 1958
rect 3420 1955 3421 1956
rect 3415 1954 3421 1955
rect 3430 1955 3431 1956
rect 3435 1955 3436 1959
rect 3430 1954 3436 1955
rect 1270 1950 1276 1951
rect 348 1944 398 1946
rect 402 1947 408 1948
rect 348 1943 349 1944
rect 343 1942 349 1943
rect 402 1943 403 1947
rect 407 1946 408 1947
rect 471 1947 477 1948
rect 471 1946 472 1947
rect 407 1944 472 1946
rect 407 1943 408 1944
rect 402 1942 408 1943
rect 471 1943 472 1944
rect 476 1943 477 1947
rect 471 1942 477 1943
rect 494 1947 500 1948
rect 494 1943 495 1947
rect 499 1946 500 1947
rect 607 1947 613 1948
rect 607 1946 608 1947
rect 499 1944 608 1946
rect 499 1943 500 1944
rect 494 1942 500 1943
rect 607 1943 608 1944
rect 612 1943 613 1947
rect 607 1942 613 1943
rect 630 1947 636 1948
rect 630 1943 631 1947
rect 635 1946 636 1947
rect 751 1947 757 1948
rect 751 1946 752 1947
rect 635 1944 752 1946
rect 635 1943 636 1944
rect 630 1942 636 1943
rect 751 1943 752 1944
rect 756 1943 757 1947
rect 751 1942 757 1943
rect 903 1947 909 1948
rect 903 1943 904 1947
rect 908 1946 909 1947
rect 950 1947 956 1948
rect 950 1946 951 1947
rect 908 1944 951 1946
rect 908 1943 909 1944
rect 903 1942 909 1943
rect 950 1943 951 1944
rect 955 1943 956 1947
rect 1055 1947 1061 1948
rect 1055 1946 1056 1947
rect 950 1942 956 1943
rect 980 1944 1056 1946
rect 110 1932 116 1933
rect 110 1928 111 1932
rect 115 1928 116 1932
rect 110 1927 116 1928
rect 294 1931 300 1932
rect 294 1927 295 1931
rect 299 1927 300 1931
rect 294 1926 300 1927
rect 422 1931 428 1932
rect 422 1927 423 1931
rect 427 1927 428 1931
rect 422 1926 428 1927
rect 558 1931 564 1932
rect 558 1927 559 1931
rect 563 1927 564 1931
rect 558 1926 564 1927
rect 702 1931 708 1932
rect 702 1927 703 1931
rect 707 1927 708 1931
rect 702 1926 708 1927
rect 854 1931 860 1932
rect 854 1927 855 1931
rect 859 1927 860 1931
rect 980 1930 982 1944
rect 1055 1943 1056 1944
rect 1060 1943 1061 1947
rect 1055 1942 1061 1943
rect 1207 1947 1213 1948
rect 1207 1943 1208 1947
rect 1212 1946 1213 1947
rect 1238 1947 1244 1948
rect 1238 1946 1239 1947
rect 1212 1944 1239 1946
rect 1212 1943 1213 1944
rect 1207 1942 1213 1943
rect 1238 1943 1239 1944
rect 1243 1943 1244 1947
rect 1238 1942 1244 1943
rect 1359 1947 1365 1948
rect 1359 1943 1360 1947
rect 1364 1946 1365 1947
rect 1390 1947 1396 1948
rect 1390 1946 1391 1947
rect 1364 1944 1391 1946
rect 1364 1943 1365 1944
rect 1359 1942 1365 1943
rect 1390 1943 1391 1944
rect 1395 1943 1396 1947
rect 1390 1942 1396 1943
rect 1398 1947 1404 1948
rect 1398 1943 1399 1947
rect 1403 1946 1404 1947
rect 1519 1947 1525 1948
rect 1519 1946 1520 1947
rect 1403 1944 1520 1946
rect 1403 1943 1404 1944
rect 1398 1942 1404 1943
rect 1519 1943 1520 1944
rect 1524 1943 1525 1947
rect 1519 1942 1525 1943
rect 1806 1944 1812 1945
rect 3462 1944 3468 1945
rect 1806 1940 1807 1944
rect 1811 1940 1812 1944
rect 1806 1939 1812 1940
rect 1862 1943 1868 1944
rect 1862 1939 1863 1943
rect 1867 1939 1868 1943
rect 1862 1938 1868 1939
rect 1998 1943 2004 1944
rect 1998 1939 1999 1943
rect 2003 1939 2004 1943
rect 1998 1938 2004 1939
rect 2142 1943 2148 1944
rect 2142 1939 2143 1943
rect 2147 1939 2148 1943
rect 2142 1938 2148 1939
rect 2286 1943 2292 1944
rect 2286 1939 2287 1943
rect 2291 1939 2292 1943
rect 2286 1938 2292 1939
rect 2430 1943 2436 1944
rect 2430 1939 2431 1943
rect 2435 1939 2436 1943
rect 2430 1938 2436 1939
rect 2574 1943 2580 1944
rect 2574 1939 2575 1943
rect 2579 1939 2580 1943
rect 2574 1938 2580 1939
rect 2710 1943 2716 1944
rect 2710 1939 2711 1943
rect 2715 1939 2716 1943
rect 2710 1938 2716 1939
rect 2830 1943 2836 1944
rect 2830 1939 2831 1943
rect 2835 1939 2836 1943
rect 2830 1938 2836 1939
rect 2950 1943 2956 1944
rect 2950 1939 2951 1943
rect 2955 1939 2956 1943
rect 2950 1938 2956 1939
rect 3062 1943 3068 1944
rect 3062 1939 3063 1943
rect 3067 1939 3068 1943
rect 3062 1938 3068 1939
rect 3166 1943 3172 1944
rect 3166 1939 3167 1943
rect 3171 1939 3172 1943
rect 3166 1938 3172 1939
rect 3278 1943 3284 1944
rect 3278 1939 3279 1943
rect 3283 1939 3284 1943
rect 3278 1938 3284 1939
rect 3366 1943 3372 1944
rect 3366 1939 3367 1943
rect 3371 1939 3372 1943
rect 3462 1940 3463 1944
rect 3467 1940 3468 1944
rect 3462 1939 3468 1940
rect 3366 1938 3372 1939
rect 1934 1935 1940 1936
rect 1766 1932 1772 1933
rect 854 1926 860 1927
rect 928 1928 982 1930
rect 1006 1931 1012 1932
rect 402 1923 408 1924
rect 402 1922 403 1923
rect 369 1920 403 1922
rect 402 1919 403 1920
rect 407 1919 408 1923
rect 402 1918 408 1919
rect 494 1923 500 1924
rect 494 1919 495 1923
rect 499 1919 500 1923
rect 494 1918 500 1919
rect 630 1923 636 1924
rect 630 1919 631 1923
rect 635 1919 636 1923
rect 928 1921 930 1928
rect 1006 1927 1007 1931
rect 1011 1927 1012 1931
rect 1006 1926 1012 1927
rect 1158 1931 1164 1932
rect 1158 1927 1159 1931
rect 1163 1927 1164 1931
rect 1158 1926 1164 1927
rect 1310 1931 1316 1932
rect 1310 1927 1311 1931
rect 1315 1927 1316 1931
rect 1310 1926 1316 1927
rect 1470 1931 1476 1932
rect 1470 1927 1471 1931
rect 1475 1927 1476 1931
rect 1766 1928 1767 1932
rect 1771 1928 1772 1932
rect 1934 1931 1935 1935
rect 1939 1931 1940 1935
rect 1934 1930 1940 1931
rect 1951 1935 1957 1936
rect 1951 1931 1952 1935
rect 1956 1934 1957 1935
rect 2078 1935 2084 1936
rect 1956 1932 2041 1934
rect 1956 1931 1957 1932
rect 1951 1930 1957 1931
rect 2078 1931 2079 1935
rect 2083 1934 2084 1935
rect 2358 1935 2364 1936
rect 2083 1932 2185 1934
rect 2083 1931 2084 1932
rect 2078 1930 2084 1931
rect 2358 1931 2359 1935
rect 2363 1931 2364 1935
rect 2358 1930 2364 1931
rect 2366 1935 2372 1936
rect 2366 1931 2367 1935
rect 2371 1934 2372 1935
rect 2654 1935 2660 1936
rect 2371 1932 2473 1934
rect 2371 1931 2372 1932
rect 2366 1930 2372 1931
rect 2654 1931 2655 1935
rect 2659 1934 2660 1935
rect 2798 1935 2804 1936
rect 2659 1932 2753 1934
rect 2659 1931 2660 1932
rect 2654 1930 2660 1931
rect 2798 1931 2799 1935
rect 2803 1934 2804 1935
rect 2910 1935 2916 1936
rect 2803 1932 2873 1934
rect 2803 1931 2804 1932
rect 2798 1930 2804 1931
rect 2910 1931 2911 1935
rect 2915 1934 2916 1935
rect 3134 1935 3140 1936
rect 2915 1932 2993 1934
rect 2915 1931 2916 1932
rect 2910 1930 2916 1931
rect 3134 1931 3135 1935
rect 3139 1931 3140 1935
rect 3134 1930 3140 1931
rect 3238 1935 3244 1936
rect 3238 1931 3239 1935
rect 3243 1931 3244 1935
rect 3238 1930 3244 1931
rect 3246 1935 3252 1936
rect 3246 1931 3247 1935
rect 3251 1934 3252 1935
rect 3358 1935 3364 1936
rect 3251 1932 3321 1934
rect 3251 1931 3252 1932
rect 3246 1930 3252 1931
rect 3358 1931 3359 1935
rect 3363 1934 3364 1935
rect 3363 1932 3409 1934
rect 3363 1931 3364 1932
rect 3358 1930 3364 1931
rect 1766 1927 1772 1928
rect 1806 1927 1812 1928
rect 1470 1926 1476 1927
rect 962 1923 968 1924
rect 630 1918 636 1919
rect 774 1919 780 1920
rect 110 1915 116 1916
rect 110 1911 111 1915
rect 115 1911 116 1915
rect 774 1915 775 1919
rect 779 1915 780 1919
rect 962 1919 963 1923
rect 967 1922 968 1923
rect 1238 1923 1244 1924
rect 967 1920 1049 1922
rect 967 1919 968 1920
rect 962 1918 968 1919
rect 1230 1919 1236 1920
rect 774 1914 780 1915
rect 1230 1915 1231 1919
rect 1235 1915 1236 1919
rect 1238 1919 1239 1923
rect 1243 1922 1244 1923
rect 1390 1923 1396 1924
rect 1243 1920 1353 1922
rect 1243 1919 1244 1920
rect 1238 1918 1244 1919
rect 1390 1919 1391 1923
rect 1395 1922 1396 1923
rect 1806 1923 1807 1927
rect 1811 1923 1812 1927
rect 2638 1927 2644 1928
rect 1806 1922 1812 1923
rect 1862 1924 1868 1925
rect 1395 1920 1513 1922
rect 1862 1920 1863 1924
rect 1867 1920 1868 1924
rect 1395 1919 1396 1920
rect 1862 1919 1868 1920
rect 1998 1924 2004 1925
rect 1998 1920 1999 1924
rect 2003 1920 2004 1924
rect 1998 1919 2004 1920
rect 2142 1924 2148 1925
rect 2142 1920 2143 1924
rect 2147 1920 2148 1924
rect 2142 1919 2148 1920
rect 2286 1924 2292 1925
rect 2286 1920 2287 1924
rect 2291 1920 2292 1924
rect 2286 1919 2292 1920
rect 2430 1924 2436 1925
rect 2430 1920 2431 1924
rect 2435 1920 2436 1924
rect 2430 1919 2436 1920
rect 2574 1924 2580 1925
rect 2574 1920 2575 1924
rect 2579 1920 2580 1924
rect 2638 1923 2639 1927
rect 2643 1926 2644 1927
rect 2648 1926 2650 1929
rect 2643 1924 2650 1926
rect 3462 1927 3468 1928
rect 2710 1924 2716 1925
rect 2643 1923 2644 1924
rect 2638 1922 2644 1923
rect 2574 1919 2580 1920
rect 2710 1920 2711 1924
rect 2715 1920 2716 1924
rect 2710 1919 2716 1920
rect 2830 1924 2836 1925
rect 2830 1920 2831 1924
rect 2835 1920 2836 1924
rect 2830 1919 2836 1920
rect 2950 1924 2956 1925
rect 2950 1920 2951 1924
rect 2955 1920 2956 1924
rect 2950 1919 2956 1920
rect 3062 1924 3068 1925
rect 3062 1920 3063 1924
rect 3067 1920 3068 1924
rect 3062 1919 3068 1920
rect 3166 1924 3172 1925
rect 3166 1920 3167 1924
rect 3171 1920 3172 1924
rect 3166 1919 3172 1920
rect 3278 1924 3284 1925
rect 3278 1920 3279 1924
rect 3283 1920 3284 1924
rect 3278 1919 3284 1920
rect 3366 1924 3372 1925
rect 3366 1920 3367 1924
rect 3371 1920 3372 1924
rect 3462 1923 3463 1927
rect 3467 1923 3468 1927
rect 3462 1922 3468 1923
rect 3366 1919 3372 1920
rect 1390 1918 1396 1919
rect 1230 1914 1236 1915
rect 1766 1915 1772 1916
rect 110 1910 116 1911
rect 294 1912 300 1913
rect 294 1908 295 1912
rect 299 1908 300 1912
rect 294 1907 300 1908
rect 422 1912 428 1913
rect 422 1908 423 1912
rect 427 1908 428 1912
rect 422 1907 428 1908
rect 558 1912 564 1913
rect 558 1908 559 1912
rect 563 1908 564 1912
rect 558 1907 564 1908
rect 702 1912 708 1913
rect 702 1908 703 1912
rect 707 1908 708 1912
rect 702 1907 708 1908
rect 854 1912 860 1913
rect 854 1908 855 1912
rect 859 1908 860 1912
rect 854 1907 860 1908
rect 1006 1912 1012 1913
rect 1006 1908 1007 1912
rect 1011 1908 1012 1912
rect 1006 1907 1012 1908
rect 1158 1912 1164 1913
rect 1158 1908 1159 1912
rect 1163 1908 1164 1912
rect 1158 1907 1164 1908
rect 1310 1912 1316 1913
rect 1310 1908 1311 1912
rect 1315 1908 1316 1912
rect 1310 1907 1316 1908
rect 1470 1912 1476 1913
rect 1470 1908 1471 1912
rect 1475 1908 1476 1912
rect 1766 1911 1767 1915
rect 1771 1911 1772 1915
rect 1766 1910 1772 1911
rect 1470 1907 1476 1908
rect 2014 1876 2020 1877
rect 1806 1873 1812 1874
rect 1806 1869 1807 1873
rect 1811 1869 1812 1873
rect 2014 1872 2015 1876
rect 2019 1872 2020 1876
rect 2014 1871 2020 1872
rect 2110 1876 2116 1877
rect 2110 1872 2111 1876
rect 2115 1872 2116 1876
rect 2110 1871 2116 1872
rect 2214 1876 2220 1877
rect 2214 1872 2215 1876
rect 2219 1872 2220 1876
rect 2214 1871 2220 1872
rect 2326 1876 2332 1877
rect 2326 1872 2327 1876
rect 2331 1872 2332 1876
rect 2326 1871 2332 1872
rect 2438 1876 2444 1877
rect 2438 1872 2439 1876
rect 2443 1872 2444 1876
rect 2438 1871 2444 1872
rect 2542 1876 2548 1877
rect 2542 1872 2543 1876
rect 2547 1872 2548 1876
rect 2542 1871 2548 1872
rect 2646 1876 2652 1877
rect 2646 1872 2647 1876
rect 2651 1872 2652 1876
rect 2646 1871 2652 1872
rect 2758 1876 2764 1877
rect 2758 1872 2759 1876
rect 2763 1872 2764 1876
rect 2758 1871 2764 1872
rect 2870 1876 2876 1877
rect 2870 1872 2871 1876
rect 2875 1872 2876 1876
rect 2870 1871 2876 1872
rect 2982 1876 2988 1877
rect 2982 1872 2983 1876
rect 2987 1872 2988 1876
rect 2982 1871 2988 1872
rect 3462 1873 3468 1874
rect 430 1868 436 1869
rect 110 1865 116 1866
rect 110 1861 111 1865
rect 115 1861 116 1865
rect 430 1864 431 1868
rect 435 1864 436 1868
rect 430 1863 436 1864
rect 574 1868 580 1869
rect 574 1864 575 1868
rect 579 1864 580 1868
rect 574 1863 580 1864
rect 726 1868 732 1869
rect 726 1864 727 1868
rect 731 1864 732 1868
rect 726 1863 732 1864
rect 886 1868 892 1869
rect 886 1864 887 1868
rect 891 1864 892 1868
rect 886 1863 892 1864
rect 1046 1868 1052 1869
rect 1046 1864 1047 1868
rect 1051 1864 1052 1868
rect 1046 1863 1052 1864
rect 1198 1868 1204 1869
rect 1198 1864 1199 1868
rect 1203 1864 1204 1868
rect 1198 1863 1204 1864
rect 1350 1868 1356 1869
rect 1350 1864 1351 1868
rect 1355 1864 1356 1868
rect 1350 1863 1356 1864
rect 1510 1868 1516 1869
rect 1510 1864 1511 1868
rect 1515 1864 1516 1868
rect 1510 1863 1516 1864
rect 1670 1868 1676 1869
rect 1806 1868 1812 1869
rect 3462 1869 3463 1873
rect 3467 1869 3468 1873
rect 3462 1868 3468 1869
rect 1670 1864 1671 1868
rect 1675 1864 1676 1868
rect 2086 1867 2092 1868
rect 1670 1863 1676 1864
rect 1766 1865 1772 1866
rect 110 1860 116 1861
rect 1766 1861 1767 1865
rect 1771 1861 1772 1865
rect 2086 1863 2087 1867
rect 2091 1863 2092 1867
rect 2086 1862 2092 1863
rect 2182 1867 2188 1868
rect 2182 1863 2183 1867
rect 2187 1863 2188 1867
rect 2298 1867 2304 1868
rect 2298 1866 2299 1867
rect 2289 1864 2299 1866
rect 2182 1862 2188 1863
rect 2298 1863 2299 1864
rect 2303 1863 2304 1867
rect 2298 1862 2304 1863
rect 2306 1867 2312 1868
rect 2306 1863 2307 1867
rect 2311 1866 2312 1867
rect 2406 1867 2412 1868
rect 2311 1864 2369 1866
rect 2311 1863 2312 1864
rect 2306 1862 2312 1863
rect 2406 1863 2407 1867
rect 2411 1866 2412 1867
rect 2718 1867 2724 1868
rect 2411 1864 2481 1866
rect 2411 1863 2412 1864
rect 2406 1862 2412 1863
rect 2718 1863 2719 1867
rect 2723 1863 2724 1867
rect 2718 1862 2724 1863
rect 2830 1867 2836 1868
rect 2830 1863 2831 1867
rect 2835 1863 2836 1867
rect 2830 1862 2836 1863
rect 2942 1867 2948 1868
rect 2942 1863 2943 1867
rect 2947 1863 2948 1867
rect 2942 1862 2948 1863
rect 2951 1867 2957 1868
rect 2951 1863 2952 1867
rect 2956 1866 2957 1867
rect 2956 1864 3025 1866
rect 2956 1863 2957 1864
rect 2951 1862 2957 1863
rect 1766 1860 1772 1861
rect 502 1859 508 1860
rect 502 1855 503 1859
rect 507 1855 508 1859
rect 502 1854 508 1855
rect 510 1859 516 1860
rect 510 1855 511 1859
rect 515 1858 516 1859
rect 654 1859 660 1860
rect 515 1856 617 1858
rect 515 1855 516 1856
rect 510 1854 516 1855
rect 654 1855 655 1859
rect 659 1858 660 1859
rect 950 1859 956 1860
rect 659 1856 769 1858
rect 659 1855 660 1856
rect 654 1854 660 1855
rect 950 1855 951 1859
rect 955 1855 956 1859
rect 950 1854 956 1855
rect 966 1859 972 1860
rect 966 1855 967 1859
rect 971 1858 972 1859
rect 1270 1859 1276 1860
rect 971 1856 1089 1858
rect 971 1855 972 1856
rect 966 1854 972 1855
rect 1270 1855 1271 1859
rect 1275 1855 1276 1859
rect 1270 1854 1276 1855
rect 1422 1859 1428 1860
rect 1422 1855 1423 1859
rect 1427 1855 1428 1859
rect 1422 1854 1428 1855
rect 1582 1859 1588 1860
rect 1582 1855 1583 1859
rect 1587 1855 1588 1859
rect 1582 1854 1588 1855
rect 1734 1859 1740 1860
rect 1734 1855 1735 1859
rect 1739 1855 1740 1859
rect 2615 1859 2621 1860
rect 2014 1857 2020 1858
rect 1734 1854 1740 1855
rect 1806 1856 1812 1857
rect 1806 1852 1807 1856
rect 1811 1852 1812 1856
rect 2014 1853 2015 1857
rect 2019 1853 2020 1857
rect 2014 1852 2020 1853
rect 2110 1857 2116 1858
rect 2110 1853 2111 1857
rect 2115 1853 2116 1857
rect 2110 1852 2116 1853
rect 2214 1857 2220 1858
rect 2214 1853 2215 1857
rect 2219 1853 2220 1857
rect 2214 1852 2220 1853
rect 2326 1857 2332 1858
rect 2326 1853 2327 1857
rect 2331 1853 2332 1857
rect 2326 1852 2332 1853
rect 2438 1857 2444 1858
rect 2438 1853 2439 1857
rect 2443 1853 2444 1857
rect 2438 1852 2444 1853
rect 2542 1857 2548 1858
rect 2542 1853 2543 1857
rect 2547 1853 2548 1857
rect 2615 1855 2616 1859
rect 2620 1855 2621 1859
rect 2615 1854 2621 1855
rect 2646 1857 2652 1858
rect 2542 1852 2548 1853
rect 1806 1851 1812 1852
rect 2617 1850 2619 1854
rect 2646 1853 2647 1857
rect 2651 1853 2652 1857
rect 2646 1852 2652 1853
rect 2758 1857 2764 1858
rect 2758 1853 2759 1857
rect 2763 1853 2764 1857
rect 2758 1852 2764 1853
rect 2870 1857 2876 1858
rect 2870 1853 2871 1857
rect 2875 1853 2876 1857
rect 2870 1852 2876 1853
rect 2982 1857 2988 1858
rect 2982 1853 2983 1857
rect 2987 1853 2988 1857
rect 2982 1852 2988 1853
rect 3462 1856 3468 1857
rect 3462 1852 3463 1856
rect 3467 1852 3468 1856
rect 3462 1851 3468 1852
rect 430 1849 436 1850
rect 110 1848 116 1849
rect 110 1844 111 1848
rect 115 1844 116 1848
rect 430 1845 431 1849
rect 435 1845 436 1849
rect 430 1844 436 1845
rect 574 1849 580 1850
rect 574 1845 575 1849
rect 579 1845 580 1849
rect 574 1844 580 1845
rect 726 1849 732 1850
rect 726 1845 727 1849
rect 731 1845 732 1849
rect 726 1844 732 1845
rect 886 1849 892 1850
rect 886 1845 887 1849
rect 891 1845 892 1849
rect 886 1844 892 1845
rect 1046 1849 1052 1850
rect 1046 1845 1047 1849
rect 1051 1845 1052 1849
rect 1046 1844 1052 1845
rect 1198 1849 1204 1850
rect 1198 1845 1199 1849
rect 1203 1845 1204 1849
rect 1198 1844 1204 1845
rect 1350 1849 1356 1850
rect 1350 1845 1351 1849
rect 1355 1845 1356 1849
rect 1350 1844 1356 1845
rect 1510 1849 1516 1850
rect 1510 1845 1511 1849
rect 1515 1845 1516 1849
rect 1510 1844 1516 1845
rect 1670 1849 1676 1850
rect 1670 1845 1671 1849
rect 1675 1845 1676 1849
rect 1670 1844 1676 1845
rect 1766 1848 1772 1849
rect 2617 1848 2650 1850
rect 1766 1844 1767 1848
rect 1771 1844 1772 1848
rect 110 1843 116 1844
rect 1766 1843 1772 1844
rect 2063 1839 2069 1840
rect 2063 1835 2064 1839
rect 2068 1838 2069 1839
rect 2086 1839 2092 1840
rect 2068 1836 2082 1838
rect 2068 1835 2069 1836
rect 2063 1834 2069 1835
rect 479 1831 485 1832
rect 479 1827 480 1831
rect 484 1830 485 1831
rect 510 1831 516 1832
rect 510 1830 511 1831
rect 484 1828 511 1830
rect 484 1827 485 1828
rect 479 1826 485 1827
rect 510 1827 511 1828
rect 515 1827 516 1831
rect 510 1826 516 1827
rect 623 1831 629 1832
rect 623 1827 624 1831
rect 628 1830 629 1831
rect 654 1831 660 1832
rect 654 1830 655 1831
rect 628 1828 655 1830
rect 628 1827 629 1828
rect 623 1826 629 1827
rect 654 1827 655 1828
rect 659 1827 660 1831
rect 654 1826 660 1827
rect 774 1831 781 1832
rect 774 1827 775 1831
rect 780 1827 781 1831
rect 774 1826 781 1827
rect 935 1831 941 1832
rect 935 1827 936 1831
rect 940 1830 941 1831
rect 966 1831 972 1832
rect 966 1830 967 1831
rect 940 1828 967 1830
rect 940 1827 941 1828
rect 935 1826 941 1827
rect 966 1827 967 1828
rect 971 1827 972 1831
rect 966 1826 972 1827
rect 1094 1831 1101 1832
rect 1094 1827 1095 1831
rect 1100 1827 1101 1831
rect 1094 1826 1101 1827
rect 1230 1831 1236 1832
rect 1230 1827 1231 1831
rect 1235 1830 1236 1831
rect 1247 1831 1253 1832
rect 1247 1830 1248 1831
rect 1235 1828 1248 1830
rect 1235 1827 1236 1828
rect 1230 1826 1236 1827
rect 1247 1827 1248 1828
rect 1252 1827 1253 1831
rect 1247 1826 1253 1827
rect 1270 1831 1276 1832
rect 1270 1827 1271 1831
rect 1275 1830 1276 1831
rect 1399 1831 1405 1832
rect 1399 1830 1400 1831
rect 1275 1828 1400 1830
rect 1275 1827 1276 1828
rect 1270 1826 1276 1827
rect 1399 1827 1400 1828
rect 1404 1827 1405 1831
rect 1399 1826 1405 1827
rect 1422 1831 1428 1832
rect 1422 1827 1423 1831
rect 1427 1830 1428 1831
rect 1559 1831 1565 1832
rect 1559 1830 1560 1831
rect 1427 1828 1560 1830
rect 1427 1827 1428 1828
rect 1422 1826 1428 1827
rect 1559 1827 1560 1828
rect 1564 1827 1565 1831
rect 1559 1826 1565 1827
rect 1582 1831 1588 1832
rect 1582 1827 1583 1831
rect 1587 1830 1588 1831
rect 1719 1831 1725 1832
rect 1719 1830 1720 1831
rect 1587 1828 1720 1830
rect 1587 1827 1588 1828
rect 1582 1826 1588 1827
rect 1719 1827 1720 1828
rect 1724 1827 1725 1831
rect 2080 1830 2082 1836
rect 2086 1835 2087 1839
rect 2091 1838 2092 1839
rect 2159 1839 2165 1840
rect 2159 1838 2160 1839
rect 2091 1836 2160 1838
rect 2091 1835 2092 1836
rect 2086 1834 2092 1835
rect 2159 1835 2160 1836
rect 2164 1835 2165 1839
rect 2159 1834 2165 1835
rect 2182 1839 2188 1840
rect 2182 1835 2183 1839
rect 2187 1838 2188 1839
rect 2263 1839 2269 1840
rect 2263 1838 2264 1839
rect 2187 1836 2264 1838
rect 2187 1835 2188 1836
rect 2182 1834 2188 1835
rect 2263 1835 2264 1836
rect 2268 1835 2269 1839
rect 2263 1834 2269 1835
rect 2375 1839 2381 1840
rect 2375 1835 2376 1839
rect 2380 1838 2381 1839
rect 2406 1839 2412 1840
rect 2406 1838 2407 1839
rect 2380 1836 2407 1838
rect 2380 1835 2381 1836
rect 2375 1834 2381 1835
rect 2406 1835 2407 1836
rect 2411 1835 2412 1839
rect 2406 1834 2412 1835
rect 2487 1839 2493 1840
rect 2487 1835 2488 1839
rect 2492 1838 2493 1839
rect 2526 1839 2532 1840
rect 2526 1838 2527 1839
rect 2492 1836 2527 1838
rect 2492 1835 2493 1836
rect 2487 1834 2493 1835
rect 2526 1835 2527 1836
rect 2531 1835 2532 1839
rect 2526 1834 2532 1835
rect 2591 1839 2597 1840
rect 2591 1835 2592 1839
rect 2596 1838 2597 1839
rect 2638 1839 2644 1840
rect 2638 1838 2639 1839
rect 2596 1836 2639 1838
rect 2596 1835 2597 1836
rect 2591 1834 2597 1835
rect 2638 1835 2639 1836
rect 2643 1835 2644 1839
rect 2648 1838 2650 1848
rect 2695 1839 2701 1840
rect 2695 1838 2696 1839
rect 2648 1836 2696 1838
rect 2638 1834 2644 1835
rect 2695 1835 2696 1836
rect 2700 1835 2701 1839
rect 2695 1834 2701 1835
rect 2718 1839 2724 1840
rect 2718 1835 2719 1839
rect 2723 1838 2724 1839
rect 2807 1839 2813 1840
rect 2807 1838 2808 1839
rect 2723 1836 2808 1838
rect 2723 1835 2724 1836
rect 2718 1834 2724 1835
rect 2807 1835 2808 1836
rect 2812 1835 2813 1839
rect 2807 1834 2813 1835
rect 2830 1839 2836 1840
rect 2830 1835 2831 1839
rect 2835 1838 2836 1839
rect 2919 1839 2925 1840
rect 2919 1838 2920 1839
rect 2835 1836 2920 1838
rect 2835 1835 2836 1836
rect 2830 1834 2836 1835
rect 2919 1835 2920 1836
rect 2924 1835 2925 1839
rect 2919 1834 2925 1835
rect 2942 1839 2948 1840
rect 2942 1835 2943 1839
rect 2947 1838 2948 1839
rect 3031 1839 3037 1840
rect 3031 1838 3032 1839
rect 2947 1836 3032 1838
rect 2947 1835 2948 1836
rect 2942 1834 2948 1835
rect 3031 1835 3032 1836
rect 3036 1835 3037 1839
rect 3031 1834 3037 1835
rect 2306 1831 2312 1832
rect 2306 1830 2307 1831
rect 2080 1828 2307 1830
rect 1719 1826 1725 1827
rect 2306 1827 2307 1828
rect 2311 1827 2312 1831
rect 2306 1826 2312 1827
rect 2710 1827 2716 1828
rect 2710 1826 2711 1827
rect 2608 1824 2711 1826
rect 1358 1823 1364 1824
rect 1358 1822 1359 1823
rect 1216 1820 1359 1822
rect 502 1815 508 1816
rect 502 1811 503 1815
rect 507 1814 508 1815
rect 559 1815 565 1816
rect 559 1814 560 1815
rect 507 1812 560 1814
rect 507 1811 508 1812
rect 502 1810 508 1811
rect 559 1811 560 1812
rect 564 1811 565 1815
rect 559 1810 565 1811
rect 582 1815 588 1816
rect 582 1811 583 1815
rect 587 1814 588 1815
rect 679 1815 685 1816
rect 679 1814 680 1815
rect 587 1812 680 1814
rect 587 1811 588 1812
rect 582 1810 588 1811
rect 679 1811 680 1812
rect 684 1811 685 1815
rect 679 1810 685 1811
rect 807 1815 813 1816
rect 807 1811 808 1815
rect 812 1814 813 1815
rect 822 1815 828 1816
rect 822 1814 823 1815
rect 812 1812 823 1814
rect 812 1811 813 1812
rect 807 1810 813 1811
rect 822 1811 823 1812
rect 827 1811 828 1815
rect 822 1810 828 1811
rect 830 1815 836 1816
rect 830 1811 831 1815
rect 835 1814 836 1815
rect 935 1815 941 1816
rect 935 1814 936 1815
rect 835 1812 936 1814
rect 835 1811 836 1812
rect 830 1810 836 1811
rect 935 1811 936 1812
rect 940 1811 941 1815
rect 935 1810 941 1811
rect 958 1815 964 1816
rect 958 1811 959 1815
rect 963 1814 964 1815
rect 1071 1815 1077 1816
rect 1071 1814 1072 1815
rect 963 1812 1072 1814
rect 963 1811 964 1812
rect 958 1810 964 1811
rect 1071 1811 1072 1812
rect 1076 1811 1077 1815
rect 1071 1810 1077 1811
rect 1199 1815 1205 1816
rect 1199 1811 1200 1815
rect 1204 1814 1205 1815
rect 1216 1814 1218 1820
rect 1358 1819 1359 1820
rect 1363 1819 1364 1823
rect 1358 1818 1364 1819
rect 2151 1819 2157 1820
rect 1204 1812 1218 1814
rect 1222 1815 1228 1816
rect 1204 1811 1205 1812
rect 1199 1810 1205 1811
rect 1222 1811 1223 1815
rect 1227 1814 1228 1815
rect 1327 1815 1333 1816
rect 1327 1814 1328 1815
rect 1227 1812 1328 1814
rect 1227 1811 1228 1812
rect 1222 1810 1228 1811
rect 1327 1811 1328 1812
rect 1332 1811 1333 1815
rect 1327 1810 1333 1811
rect 1455 1815 1461 1816
rect 1455 1811 1456 1815
rect 1460 1814 1461 1815
rect 1486 1815 1492 1816
rect 1486 1814 1487 1815
rect 1460 1812 1487 1814
rect 1460 1811 1461 1812
rect 1455 1810 1461 1811
rect 1486 1811 1487 1812
rect 1491 1811 1492 1815
rect 1486 1810 1492 1811
rect 1583 1815 1589 1816
rect 1583 1811 1584 1815
rect 1588 1814 1589 1815
rect 1614 1815 1620 1816
rect 1614 1814 1615 1815
rect 1588 1812 1615 1814
rect 1588 1811 1589 1812
rect 1583 1810 1589 1811
rect 1614 1811 1615 1812
rect 1619 1811 1620 1815
rect 1614 1810 1620 1811
rect 1719 1815 1725 1816
rect 1719 1811 1720 1815
rect 1724 1814 1725 1815
rect 1734 1815 1740 1816
rect 1734 1814 1735 1815
rect 1724 1812 1735 1814
rect 1724 1811 1725 1812
rect 1719 1810 1725 1811
rect 1734 1811 1735 1812
rect 1739 1811 1740 1815
rect 2151 1815 2152 1819
rect 2156 1818 2157 1819
rect 2206 1819 2212 1820
rect 2206 1818 2207 1819
rect 2156 1816 2207 1818
rect 2156 1815 2157 1816
rect 2151 1814 2157 1815
rect 2206 1815 2207 1816
rect 2211 1815 2212 1819
rect 2239 1819 2245 1820
rect 2239 1818 2240 1819
rect 2206 1814 2212 1815
rect 2216 1816 2240 1818
rect 1734 1810 1740 1811
rect 2216 1810 2218 1816
rect 2239 1815 2240 1816
rect 2244 1815 2245 1819
rect 2239 1814 2245 1815
rect 2262 1819 2268 1820
rect 2262 1815 2263 1819
rect 2267 1818 2268 1819
rect 2327 1819 2333 1820
rect 2327 1818 2328 1819
rect 2267 1816 2328 1818
rect 2267 1815 2268 1816
rect 2262 1814 2268 1815
rect 2327 1815 2328 1816
rect 2332 1815 2333 1819
rect 2327 1814 2333 1815
rect 2350 1819 2356 1820
rect 2350 1815 2351 1819
rect 2355 1818 2356 1819
rect 2415 1819 2421 1820
rect 2415 1818 2416 1819
rect 2355 1816 2416 1818
rect 2355 1815 2356 1816
rect 2350 1814 2356 1815
rect 2415 1815 2416 1816
rect 2420 1815 2421 1819
rect 2415 1814 2421 1815
rect 2447 1819 2453 1820
rect 2447 1815 2448 1819
rect 2452 1818 2453 1819
rect 2503 1819 2509 1820
rect 2503 1818 2504 1819
rect 2452 1816 2504 1818
rect 2452 1815 2453 1816
rect 2447 1814 2453 1815
rect 2503 1815 2504 1816
rect 2508 1815 2509 1819
rect 2503 1814 2509 1815
rect 2591 1819 2597 1820
rect 2591 1815 2592 1819
rect 2596 1818 2597 1819
rect 2608 1818 2610 1824
rect 2710 1823 2711 1824
rect 2715 1823 2716 1827
rect 2710 1822 2716 1823
rect 2951 1823 2957 1824
rect 2951 1822 2952 1823
rect 2943 1821 2952 1822
rect 2596 1816 2610 1818
rect 2614 1819 2620 1820
rect 2596 1815 2597 1816
rect 2591 1814 2597 1815
rect 2614 1815 2615 1819
rect 2619 1818 2620 1819
rect 2679 1819 2685 1820
rect 2679 1818 2680 1819
rect 2619 1816 2680 1818
rect 2619 1815 2620 1816
rect 2614 1814 2620 1815
rect 2679 1815 2680 1816
rect 2684 1815 2685 1819
rect 2679 1814 2685 1815
rect 2767 1819 2773 1820
rect 2767 1815 2768 1819
rect 2772 1818 2773 1819
rect 2799 1819 2805 1820
rect 2799 1818 2800 1819
rect 2772 1816 2800 1818
rect 2772 1815 2773 1816
rect 2767 1814 2773 1815
rect 2799 1815 2800 1816
rect 2804 1815 2805 1819
rect 2799 1814 2805 1815
rect 2855 1819 2861 1820
rect 2855 1815 2856 1819
rect 2860 1818 2861 1819
rect 2886 1819 2892 1820
rect 2886 1818 2887 1819
rect 2860 1816 2887 1818
rect 2860 1815 2861 1816
rect 2855 1814 2861 1815
rect 2886 1815 2887 1816
rect 2891 1815 2892 1819
rect 2943 1817 2944 1821
rect 2948 1820 2952 1821
rect 2948 1817 2949 1820
rect 2951 1819 2952 1820
rect 2956 1819 2957 1823
rect 2951 1818 2957 1819
rect 2943 1816 2949 1817
rect 2886 1814 2892 1815
rect 2184 1808 2218 1810
rect 1806 1804 1812 1805
rect 110 1800 116 1801
rect 1766 1800 1772 1801
rect 110 1796 111 1800
rect 115 1796 116 1800
rect 110 1795 116 1796
rect 510 1799 516 1800
rect 510 1795 511 1799
rect 515 1795 516 1799
rect 510 1794 516 1795
rect 630 1799 636 1800
rect 630 1795 631 1799
rect 635 1795 636 1799
rect 630 1794 636 1795
rect 758 1799 764 1800
rect 758 1795 759 1799
rect 763 1795 764 1799
rect 758 1794 764 1795
rect 886 1799 892 1800
rect 886 1795 887 1799
rect 891 1795 892 1799
rect 886 1794 892 1795
rect 1022 1799 1028 1800
rect 1022 1795 1023 1799
rect 1027 1795 1028 1799
rect 1022 1794 1028 1795
rect 1150 1799 1156 1800
rect 1150 1795 1151 1799
rect 1155 1795 1156 1799
rect 1150 1794 1156 1795
rect 1278 1799 1284 1800
rect 1278 1795 1279 1799
rect 1283 1795 1284 1799
rect 1278 1794 1284 1795
rect 1406 1799 1412 1800
rect 1406 1795 1407 1799
rect 1411 1795 1412 1799
rect 1406 1794 1412 1795
rect 1534 1799 1540 1800
rect 1534 1795 1535 1799
rect 1539 1795 1540 1799
rect 1534 1794 1540 1795
rect 1670 1799 1676 1800
rect 1670 1795 1671 1799
rect 1675 1795 1676 1799
rect 1766 1796 1767 1800
rect 1771 1796 1772 1800
rect 1806 1800 1807 1804
rect 1811 1800 1812 1804
rect 1806 1799 1812 1800
rect 2102 1803 2108 1804
rect 2102 1799 2103 1803
rect 2107 1799 2108 1803
rect 2102 1798 2108 1799
rect 1766 1795 1772 1796
rect 1670 1794 1676 1795
rect 2184 1794 2186 1808
rect 3462 1804 3468 1805
rect 2190 1803 2196 1804
rect 2190 1799 2191 1803
rect 2195 1799 2196 1803
rect 2190 1798 2196 1799
rect 2278 1803 2284 1804
rect 2278 1799 2279 1803
rect 2283 1799 2284 1803
rect 2278 1798 2284 1799
rect 2366 1803 2372 1804
rect 2366 1799 2367 1803
rect 2371 1799 2372 1803
rect 2366 1798 2372 1799
rect 2454 1803 2460 1804
rect 2454 1799 2455 1803
rect 2459 1799 2460 1803
rect 2454 1798 2460 1799
rect 2542 1803 2548 1804
rect 2542 1799 2543 1803
rect 2547 1799 2548 1803
rect 2542 1798 2548 1799
rect 2630 1803 2636 1804
rect 2630 1799 2631 1803
rect 2635 1799 2636 1803
rect 2630 1798 2636 1799
rect 2718 1803 2724 1804
rect 2718 1799 2719 1803
rect 2723 1799 2724 1803
rect 2718 1798 2724 1799
rect 2806 1803 2812 1804
rect 2806 1799 2807 1803
rect 2811 1799 2812 1803
rect 2806 1798 2812 1799
rect 2894 1803 2900 1804
rect 2894 1799 2895 1803
rect 2899 1799 2900 1803
rect 3462 1800 3463 1804
rect 3467 1800 3468 1804
rect 3462 1799 3468 1800
rect 2894 1798 2900 1799
rect 2177 1792 2186 1794
rect 2262 1795 2268 1796
rect 582 1791 588 1792
rect 582 1787 583 1791
rect 587 1787 588 1791
rect 830 1791 836 1792
rect 582 1786 588 1787
rect 702 1787 708 1788
rect 110 1783 116 1784
rect 110 1779 111 1783
rect 115 1779 116 1783
rect 702 1783 703 1787
rect 707 1783 708 1787
rect 830 1787 831 1791
rect 835 1787 836 1791
rect 830 1786 836 1787
rect 958 1791 964 1792
rect 958 1787 959 1791
rect 963 1787 964 1791
rect 958 1786 964 1787
rect 1094 1791 1100 1792
rect 1094 1787 1095 1791
rect 1099 1787 1100 1791
rect 1094 1786 1100 1787
rect 1222 1791 1228 1792
rect 1222 1787 1223 1791
rect 1227 1787 1228 1791
rect 1222 1786 1228 1787
rect 1358 1791 1364 1792
rect 1358 1787 1359 1791
rect 1363 1790 1364 1791
rect 1486 1791 1492 1792
rect 1363 1788 1449 1790
rect 1363 1787 1364 1788
rect 1358 1786 1364 1787
rect 1486 1787 1487 1791
rect 1491 1790 1492 1791
rect 1614 1791 1620 1792
rect 1491 1788 1577 1790
rect 1491 1787 1492 1788
rect 1486 1786 1492 1787
rect 1614 1787 1615 1791
rect 1619 1790 1620 1791
rect 2262 1791 2263 1795
rect 2267 1791 2268 1795
rect 2262 1790 2268 1791
rect 2350 1795 2356 1796
rect 2350 1791 2351 1795
rect 2355 1791 2356 1795
rect 2447 1795 2453 1796
rect 2447 1794 2448 1795
rect 2441 1792 2448 1794
rect 2350 1790 2356 1791
rect 2447 1791 2448 1792
rect 2452 1791 2453 1795
rect 2447 1790 2453 1791
rect 2526 1795 2532 1796
rect 2526 1791 2527 1795
rect 2531 1791 2532 1795
rect 2526 1790 2532 1791
rect 2614 1795 2620 1796
rect 2614 1791 2615 1795
rect 2619 1791 2620 1795
rect 2710 1795 2716 1796
rect 2614 1790 2620 1791
rect 2702 1791 2708 1792
rect 1619 1788 1713 1790
rect 1619 1787 1620 1788
rect 1614 1786 1620 1787
rect 1806 1787 1812 1788
rect 702 1782 708 1783
rect 1352 1782 1354 1785
rect 1362 1783 1368 1784
rect 1362 1782 1363 1783
rect 110 1778 116 1779
rect 510 1780 516 1781
rect 510 1776 511 1780
rect 515 1776 516 1780
rect 510 1775 516 1776
rect 630 1780 636 1781
rect 630 1776 631 1780
rect 635 1776 636 1780
rect 630 1775 636 1776
rect 758 1780 764 1781
rect 758 1776 759 1780
rect 763 1776 764 1780
rect 758 1775 764 1776
rect 886 1780 892 1781
rect 886 1776 887 1780
rect 891 1776 892 1780
rect 886 1775 892 1776
rect 1022 1780 1028 1781
rect 1022 1776 1023 1780
rect 1027 1776 1028 1780
rect 1022 1775 1028 1776
rect 1150 1780 1156 1781
rect 1150 1776 1151 1780
rect 1155 1776 1156 1780
rect 1150 1775 1156 1776
rect 1278 1780 1284 1781
rect 1352 1780 1363 1782
rect 1278 1776 1279 1780
rect 1283 1776 1284 1780
rect 1362 1779 1363 1780
rect 1367 1779 1368 1783
rect 1766 1783 1772 1784
rect 1362 1778 1368 1779
rect 1406 1780 1412 1781
rect 1278 1775 1284 1776
rect 1406 1776 1407 1780
rect 1411 1776 1412 1780
rect 1406 1775 1412 1776
rect 1534 1780 1540 1781
rect 1534 1776 1535 1780
rect 1539 1776 1540 1780
rect 1534 1775 1540 1776
rect 1670 1780 1676 1781
rect 1670 1776 1671 1780
rect 1675 1776 1676 1780
rect 1766 1779 1767 1783
rect 1771 1779 1772 1783
rect 1806 1783 1807 1787
rect 1811 1783 1812 1787
rect 2702 1787 2703 1791
rect 2707 1787 2708 1791
rect 2710 1791 2711 1795
rect 2715 1794 2716 1795
rect 2799 1795 2805 1796
rect 2715 1792 2761 1794
rect 2715 1791 2716 1792
rect 2710 1790 2716 1791
rect 2799 1791 2800 1795
rect 2804 1794 2805 1795
rect 2886 1795 2892 1796
rect 2804 1792 2849 1794
rect 2804 1791 2805 1792
rect 2799 1790 2805 1791
rect 2886 1791 2887 1795
rect 2891 1794 2892 1795
rect 2891 1792 2937 1794
rect 2891 1791 2892 1792
rect 2886 1790 2892 1791
rect 2702 1786 2708 1787
rect 3462 1787 3468 1788
rect 1806 1782 1812 1783
rect 2102 1784 2108 1785
rect 2102 1780 2103 1784
rect 2107 1780 2108 1784
rect 2102 1779 2108 1780
rect 2190 1784 2196 1785
rect 2190 1780 2191 1784
rect 2195 1780 2196 1784
rect 2190 1779 2196 1780
rect 2278 1784 2284 1785
rect 2278 1780 2279 1784
rect 2283 1780 2284 1784
rect 2278 1779 2284 1780
rect 2366 1784 2372 1785
rect 2366 1780 2367 1784
rect 2371 1780 2372 1784
rect 2366 1779 2372 1780
rect 2454 1784 2460 1785
rect 2454 1780 2455 1784
rect 2459 1780 2460 1784
rect 2454 1779 2460 1780
rect 2542 1784 2548 1785
rect 2542 1780 2543 1784
rect 2547 1780 2548 1784
rect 2542 1779 2548 1780
rect 2630 1784 2636 1785
rect 2630 1780 2631 1784
rect 2635 1780 2636 1784
rect 2630 1779 2636 1780
rect 2718 1784 2724 1785
rect 2718 1780 2719 1784
rect 2723 1780 2724 1784
rect 2718 1779 2724 1780
rect 2806 1784 2812 1785
rect 2806 1780 2807 1784
rect 2811 1780 2812 1784
rect 2806 1779 2812 1780
rect 2894 1784 2900 1785
rect 2894 1780 2895 1784
rect 2899 1780 2900 1784
rect 3462 1783 3463 1787
rect 3467 1783 3468 1787
rect 3462 1782 3468 1783
rect 2894 1779 2900 1780
rect 1766 1778 1772 1779
rect 1670 1775 1676 1776
rect 438 1732 444 1733
rect 110 1729 116 1730
rect 110 1725 111 1729
rect 115 1725 116 1729
rect 438 1728 439 1732
rect 443 1728 444 1732
rect 438 1727 444 1728
rect 534 1732 540 1733
rect 534 1728 535 1732
rect 539 1728 540 1732
rect 534 1727 540 1728
rect 638 1732 644 1733
rect 638 1728 639 1732
rect 643 1728 644 1732
rect 638 1727 644 1728
rect 742 1732 748 1733
rect 742 1728 743 1732
rect 747 1728 748 1732
rect 742 1727 748 1728
rect 846 1732 852 1733
rect 846 1728 847 1732
rect 851 1728 852 1732
rect 846 1727 852 1728
rect 950 1732 956 1733
rect 950 1728 951 1732
rect 955 1728 956 1732
rect 950 1727 956 1728
rect 1054 1732 1060 1733
rect 1054 1728 1055 1732
rect 1059 1728 1060 1732
rect 1054 1727 1060 1728
rect 1158 1732 1164 1733
rect 1158 1728 1159 1732
rect 1163 1728 1164 1732
rect 1158 1727 1164 1728
rect 1270 1732 1276 1733
rect 1270 1728 1271 1732
rect 1275 1728 1276 1732
rect 1270 1727 1276 1728
rect 1382 1732 1388 1733
rect 1382 1728 1383 1732
rect 1387 1728 1388 1732
rect 1382 1727 1388 1728
rect 1766 1729 1772 1730
rect 110 1724 116 1725
rect 1766 1725 1767 1729
rect 1771 1725 1772 1729
rect 2142 1728 2148 1729
rect 1766 1724 1772 1725
rect 1806 1725 1812 1726
rect 502 1723 508 1724
rect 502 1719 503 1723
rect 507 1719 508 1723
rect 502 1718 508 1719
rect 518 1723 524 1724
rect 518 1719 519 1723
rect 523 1722 524 1723
rect 614 1723 620 1724
rect 523 1720 577 1722
rect 523 1719 524 1720
rect 518 1718 524 1719
rect 614 1719 615 1723
rect 619 1722 620 1723
rect 814 1723 820 1724
rect 619 1720 681 1722
rect 619 1719 620 1720
rect 614 1718 620 1719
rect 814 1719 815 1723
rect 819 1719 820 1723
rect 814 1718 820 1719
rect 822 1723 828 1724
rect 822 1719 823 1723
rect 827 1722 828 1723
rect 1030 1723 1036 1724
rect 827 1720 889 1722
rect 827 1719 828 1720
rect 822 1718 828 1719
rect 1030 1719 1031 1723
rect 1035 1722 1036 1723
rect 1134 1723 1140 1724
rect 1035 1720 1097 1722
rect 1035 1719 1036 1720
rect 1030 1718 1036 1719
rect 1134 1719 1135 1723
rect 1139 1722 1140 1723
rect 1238 1723 1244 1724
rect 1139 1720 1201 1722
rect 1139 1719 1140 1720
rect 1134 1718 1140 1719
rect 1238 1719 1239 1723
rect 1243 1722 1244 1723
rect 1350 1723 1356 1724
rect 1243 1720 1313 1722
rect 1243 1719 1244 1720
rect 1238 1718 1244 1719
rect 1350 1719 1351 1723
rect 1355 1722 1356 1723
rect 1355 1720 1425 1722
rect 1806 1721 1807 1725
rect 1811 1721 1812 1725
rect 2142 1724 2143 1728
rect 2147 1724 2148 1728
rect 2142 1723 2148 1724
rect 2230 1728 2236 1729
rect 2230 1724 2231 1728
rect 2235 1724 2236 1728
rect 2230 1723 2236 1724
rect 2318 1728 2324 1729
rect 2318 1724 2319 1728
rect 2323 1724 2324 1728
rect 2318 1723 2324 1724
rect 2406 1728 2412 1729
rect 2406 1724 2407 1728
rect 2411 1724 2412 1728
rect 2406 1723 2412 1724
rect 2494 1728 2500 1729
rect 2494 1724 2495 1728
rect 2499 1724 2500 1728
rect 2494 1723 2500 1724
rect 2582 1728 2588 1729
rect 2582 1724 2583 1728
rect 2587 1724 2588 1728
rect 2582 1723 2588 1724
rect 2670 1728 2676 1729
rect 2670 1724 2671 1728
rect 2675 1724 2676 1728
rect 2670 1723 2676 1724
rect 2758 1728 2764 1729
rect 2758 1724 2759 1728
rect 2763 1724 2764 1728
rect 2758 1723 2764 1724
rect 2846 1728 2852 1729
rect 2846 1724 2847 1728
rect 2851 1724 2852 1728
rect 2846 1723 2852 1724
rect 3462 1725 3468 1726
rect 1806 1720 1812 1721
rect 3462 1721 3463 1725
rect 3467 1721 3468 1725
rect 3462 1720 3468 1721
rect 1355 1719 1356 1720
rect 1350 1718 1356 1719
rect 2206 1719 2212 1720
rect 1023 1715 1029 1716
rect 438 1713 444 1714
rect 110 1712 116 1713
rect 110 1708 111 1712
rect 115 1708 116 1712
rect 438 1709 439 1713
rect 443 1709 444 1713
rect 438 1708 444 1709
rect 534 1713 540 1714
rect 534 1709 535 1713
rect 539 1709 540 1713
rect 534 1708 540 1709
rect 638 1713 644 1714
rect 638 1709 639 1713
rect 643 1709 644 1713
rect 638 1708 644 1709
rect 742 1713 748 1714
rect 742 1709 743 1713
rect 747 1709 748 1713
rect 742 1708 748 1709
rect 846 1713 852 1714
rect 846 1709 847 1713
rect 851 1709 852 1713
rect 846 1708 852 1709
rect 950 1713 956 1714
rect 950 1709 951 1713
rect 955 1709 956 1713
rect 1023 1711 1024 1715
rect 1028 1714 1029 1715
rect 2206 1715 2207 1719
rect 2211 1715 2212 1719
rect 2206 1714 2212 1715
rect 2222 1719 2228 1720
rect 2222 1715 2223 1719
rect 2227 1718 2228 1719
rect 2310 1719 2316 1720
rect 2227 1716 2273 1718
rect 2227 1715 2228 1716
rect 2222 1714 2228 1715
rect 2310 1715 2311 1719
rect 2315 1718 2316 1719
rect 2398 1719 2404 1720
rect 2315 1716 2361 1718
rect 2315 1715 2316 1716
rect 2310 1714 2316 1715
rect 2398 1715 2399 1719
rect 2403 1718 2404 1719
rect 2486 1719 2492 1720
rect 2403 1716 2449 1718
rect 2403 1715 2404 1716
rect 2398 1714 2404 1715
rect 2486 1715 2487 1719
rect 2491 1718 2492 1719
rect 2646 1719 2652 1720
rect 2491 1716 2537 1718
rect 2491 1715 2492 1716
rect 2486 1714 2492 1715
rect 2646 1715 2647 1719
rect 2651 1715 2652 1719
rect 2646 1714 2652 1715
rect 2742 1719 2748 1720
rect 2742 1715 2743 1719
rect 2747 1715 2748 1719
rect 2742 1714 2748 1715
rect 2830 1719 2836 1720
rect 2830 1715 2831 1719
rect 2835 1715 2836 1719
rect 2830 1714 2836 1715
rect 2839 1719 2845 1720
rect 2839 1715 2840 1719
rect 2844 1718 2845 1719
rect 2844 1716 2889 1718
rect 2844 1715 2845 1716
rect 2839 1714 2845 1715
rect 1028 1712 1046 1714
rect 1028 1711 1029 1712
rect 1023 1710 1029 1711
rect 950 1708 956 1709
rect 110 1707 116 1708
rect 1044 1706 1046 1712
rect 1054 1713 1060 1714
rect 1054 1709 1055 1713
rect 1059 1709 1060 1713
rect 1054 1708 1060 1709
rect 1158 1713 1164 1714
rect 1158 1709 1159 1713
rect 1163 1709 1164 1713
rect 1158 1708 1164 1709
rect 1270 1713 1276 1714
rect 1270 1709 1271 1713
rect 1275 1709 1276 1713
rect 1270 1708 1276 1709
rect 1382 1713 1388 1714
rect 1382 1709 1383 1713
rect 1387 1709 1388 1713
rect 1382 1708 1388 1709
rect 1766 1712 1772 1713
rect 1766 1708 1767 1712
rect 1771 1708 1772 1712
rect 2142 1709 2148 1710
rect 1078 1707 1084 1708
rect 1766 1707 1772 1708
rect 1806 1708 1812 1709
rect 1078 1706 1079 1707
rect 1044 1704 1079 1706
rect 1078 1703 1079 1704
rect 1083 1703 1084 1707
rect 1806 1704 1807 1708
rect 1811 1704 1812 1708
rect 2142 1705 2143 1709
rect 2147 1705 2148 1709
rect 2142 1704 2148 1705
rect 2230 1709 2236 1710
rect 2230 1705 2231 1709
rect 2235 1705 2236 1709
rect 2230 1704 2236 1705
rect 2318 1709 2324 1710
rect 2318 1705 2319 1709
rect 2323 1705 2324 1709
rect 2318 1704 2324 1705
rect 2406 1709 2412 1710
rect 2406 1705 2407 1709
rect 2411 1705 2412 1709
rect 2406 1704 2412 1705
rect 2494 1709 2500 1710
rect 2494 1705 2495 1709
rect 2499 1705 2500 1709
rect 2494 1704 2500 1705
rect 2582 1709 2588 1710
rect 2582 1705 2583 1709
rect 2587 1705 2588 1709
rect 2582 1704 2588 1705
rect 2670 1709 2676 1710
rect 2670 1705 2671 1709
rect 2675 1705 2676 1709
rect 2670 1704 2676 1705
rect 2758 1709 2764 1710
rect 2758 1705 2759 1709
rect 2763 1705 2764 1709
rect 2758 1704 2764 1705
rect 2846 1709 2852 1710
rect 2846 1705 2847 1709
rect 2851 1705 2852 1709
rect 2846 1704 2852 1705
rect 3462 1708 3468 1709
rect 3462 1704 3463 1708
rect 3467 1704 3468 1708
rect 1806 1703 1812 1704
rect 3462 1703 3468 1704
rect 1078 1702 1084 1703
rect 487 1695 493 1696
rect 487 1691 488 1695
rect 492 1694 493 1695
rect 518 1695 524 1696
rect 518 1694 519 1695
rect 492 1692 519 1694
rect 492 1691 493 1692
rect 487 1690 493 1691
rect 518 1691 519 1692
rect 523 1691 524 1695
rect 518 1690 524 1691
rect 583 1695 589 1696
rect 583 1691 584 1695
rect 588 1694 589 1695
rect 614 1695 620 1696
rect 614 1694 615 1695
rect 588 1692 615 1694
rect 588 1691 589 1692
rect 583 1690 589 1691
rect 614 1691 615 1692
rect 619 1691 620 1695
rect 614 1690 620 1691
rect 687 1695 693 1696
rect 687 1691 688 1695
rect 692 1694 693 1695
rect 702 1695 708 1696
rect 702 1694 703 1695
rect 692 1692 703 1694
rect 692 1691 693 1692
rect 687 1690 693 1691
rect 702 1691 703 1692
rect 707 1691 708 1695
rect 702 1690 708 1691
rect 734 1695 740 1696
rect 734 1691 735 1695
rect 739 1694 740 1695
rect 791 1695 797 1696
rect 791 1694 792 1695
rect 739 1692 792 1694
rect 739 1691 740 1692
rect 734 1690 740 1691
rect 791 1691 792 1692
rect 796 1691 797 1695
rect 791 1690 797 1691
rect 814 1695 820 1696
rect 814 1691 815 1695
rect 819 1694 820 1695
rect 895 1695 901 1696
rect 895 1694 896 1695
rect 819 1692 896 1694
rect 819 1691 820 1692
rect 814 1690 820 1691
rect 895 1691 896 1692
rect 900 1691 901 1695
rect 895 1690 901 1691
rect 999 1695 1005 1696
rect 999 1691 1000 1695
rect 1004 1694 1005 1695
rect 1030 1695 1036 1696
rect 1030 1694 1031 1695
rect 1004 1692 1031 1694
rect 1004 1691 1005 1692
rect 999 1690 1005 1691
rect 1030 1691 1031 1692
rect 1035 1691 1036 1695
rect 1030 1690 1036 1691
rect 1103 1695 1109 1696
rect 1103 1691 1104 1695
rect 1108 1694 1109 1695
rect 1134 1695 1140 1696
rect 1134 1694 1135 1695
rect 1108 1692 1135 1694
rect 1108 1691 1109 1692
rect 1103 1690 1109 1691
rect 1134 1691 1135 1692
rect 1139 1691 1140 1695
rect 1134 1690 1140 1691
rect 1207 1695 1213 1696
rect 1207 1691 1208 1695
rect 1212 1694 1213 1695
rect 1238 1695 1244 1696
rect 1238 1694 1239 1695
rect 1212 1692 1239 1694
rect 1212 1691 1213 1692
rect 1207 1690 1213 1691
rect 1238 1691 1239 1692
rect 1243 1691 1244 1695
rect 1238 1690 1244 1691
rect 1319 1695 1325 1696
rect 1319 1691 1320 1695
rect 1324 1694 1325 1695
rect 1350 1695 1356 1696
rect 1350 1694 1351 1695
rect 1324 1692 1351 1694
rect 1324 1691 1325 1692
rect 1319 1690 1325 1691
rect 1350 1691 1351 1692
rect 1355 1691 1356 1695
rect 1350 1690 1356 1691
rect 1362 1695 1368 1696
rect 1362 1691 1363 1695
rect 1367 1694 1368 1695
rect 1431 1695 1437 1696
rect 1431 1694 1432 1695
rect 1367 1692 1432 1694
rect 1367 1691 1368 1692
rect 1362 1690 1368 1691
rect 1431 1691 1432 1692
rect 1436 1691 1437 1695
rect 1431 1690 1437 1691
rect 2191 1691 2197 1692
rect 1126 1687 1132 1688
rect 1126 1686 1127 1687
rect 1076 1684 1127 1686
rect 447 1679 453 1680
rect 447 1675 448 1679
rect 452 1678 453 1679
rect 502 1679 508 1680
rect 502 1678 503 1679
rect 452 1676 503 1678
rect 452 1675 453 1676
rect 447 1674 453 1675
rect 502 1675 503 1676
rect 507 1675 508 1679
rect 535 1679 541 1680
rect 535 1678 536 1679
rect 502 1674 508 1675
rect 512 1676 536 1678
rect 512 1670 514 1676
rect 535 1675 536 1676
rect 540 1675 541 1679
rect 535 1674 541 1675
rect 623 1679 629 1680
rect 623 1675 624 1679
rect 628 1678 629 1679
rect 670 1679 676 1680
rect 670 1678 671 1679
rect 628 1676 671 1678
rect 628 1675 629 1676
rect 623 1674 629 1675
rect 670 1675 671 1676
rect 675 1675 676 1679
rect 711 1679 717 1680
rect 711 1678 712 1679
rect 670 1674 676 1675
rect 680 1676 712 1678
rect 680 1670 682 1676
rect 711 1675 712 1676
rect 716 1675 717 1679
rect 711 1674 717 1675
rect 807 1679 813 1680
rect 807 1675 808 1679
rect 812 1678 813 1679
rect 838 1679 844 1680
rect 838 1678 839 1679
rect 812 1676 839 1678
rect 812 1675 813 1676
rect 807 1674 813 1675
rect 838 1675 839 1676
rect 843 1675 844 1679
rect 838 1674 844 1675
rect 903 1679 909 1680
rect 903 1675 904 1679
rect 908 1678 909 1679
rect 943 1679 949 1680
rect 943 1678 944 1679
rect 908 1676 944 1678
rect 908 1675 909 1676
rect 903 1674 909 1675
rect 943 1675 944 1676
rect 948 1675 949 1679
rect 943 1674 949 1675
rect 999 1679 1005 1680
rect 999 1675 1000 1679
rect 1004 1678 1005 1679
rect 1076 1678 1078 1684
rect 1126 1683 1127 1684
rect 1131 1683 1132 1687
rect 2191 1687 2192 1691
rect 2196 1690 2197 1691
rect 2222 1691 2228 1692
rect 2222 1690 2223 1691
rect 2196 1688 2223 1690
rect 2196 1687 2197 1688
rect 2191 1686 2197 1687
rect 2222 1687 2223 1688
rect 2227 1687 2228 1691
rect 2222 1686 2228 1687
rect 2279 1691 2285 1692
rect 2279 1687 2280 1691
rect 2284 1690 2285 1691
rect 2310 1691 2316 1692
rect 2310 1690 2311 1691
rect 2284 1688 2311 1690
rect 2284 1687 2285 1688
rect 2279 1686 2285 1687
rect 2310 1687 2311 1688
rect 2315 1687 2316 1691
rect 2310 1686 2316 1687
rect 2367 1691 2373 1692
rect 2367 1687 2368 1691
rect 2372 1690 2373 1691
rect 2398 1691 2404 1692
rect 2398 1690 2399 1691
rect 2372 1688 2399 1690
rect 2372 1687 2373 1688
rect 2367 1686 2373 1687
rect 2398 1687 2399 1688
rect 2403 1687 2404 1691
rect 2398 1686 2404 1687
rect 2455 1691 2461 1692
rect 2455 1687 2456 1691
rect 2460 1690 2461 1691
rect 2486 1691 2492 1692
rect 2486 1690 2487 1691
rect 2460 1688 2487 1690
rect 2460 1687 2461 1688
rect 2455 1686 2461 1687
rect 2486 1687 2487 1688
rect 2491 1687 2492 1691
rect 2486 1686 2492 1687
rect 2526 1691 2532 1692
rect 2526 1687 2527 1691
rect 2531 1690 2532 1691
rect 2543 1691 2549 1692
rect 2543 1690 2544 1691
rect 2531 1688 2544 1690
rect 2531 1687 2532 1688
rect 2526 1686 2532 1687
rect 2543 1687 2544 1688
rect 2548 1687 2549 1691
rect 2543 1686 2549 1687
rect 2631 1691 2637 1692
rect 2631 1687 2632 1691
rect 2636 1690 2637 1691
rect 2702 1691 2708 1692
rect 2636 1688 2698 1690
rect 2636 1687 2637 1688
rect 2631 1686 2637 1687
rect 1126 1682 1132 1683
rect 2446 1683 2452 1684
rect 2446 1682 2447 1683
rect 2168 1680 2447 1682
rect 1004 1676 1078 1678
rect 1082 1679 1088 1680
rect 1004 1675 1005 1676
rect 999 1674 1005 1675
rect 1082 1675 1083 1679
rect 1087 1678 1088 1679
rect 1095 1679 1101 1680
rect 1095 1678 1096 1679
rect 1087 1676 1096 1678
rect 1087 1675 1088 1676
rect 1082 1674 1088 1675
rect 1095 1675 1096 1676
rect 1100 1675 1101 1679
rect 1095 1674 1101 1675
rect 1118 1679 1124 1680
rect 1118 1675 1119 1679
rect 1123 1678 1124 1679
rect 1191 1679 1197 1680
rect 1191 1678 1192 1679
rect 1123 1676 1192 1678
rect 1123 1675 1124 1676
rect 1118 1674 1124 1675
rect 1191 1675 1192 1676
rect 1196 1675 1197 1679
rect 1191 1674 1197 1675
rect 2151 1675 2157 1676
rect 2151 1671 2152 1675
rect 2156 1674 2157 1675
rect 2168 1674 2170 1680
rect 2446 1679 2447 1680
rect 2451 1679 2452 1683
rect 2696 1682 2698 1688
rect 2702 1687 2703 1691
rect 2707 1690 2708 1691
rect 2719 1691 2725 1692
rect 2719 1690 2720 1691
rect 2707 1688 2720 1690
rect 2707 1687 2708 1688
rect 2702 1686 2708 1687
rect 2719 1687 2720 1688
rect 2724 1687 2725 1691
rect 2719 1686 2725 1687
rect 2742 1691 2748 1692
rect 2742 1687 2743 1691
rect 2747 1690 2748 1691
rect 2807 1691 2813 1692
rect 2807 1690 2808 1691
rect 2747 1688 2808 1690
rect 2747 1687 2748 1688
rect 2742 1686 2748 1687
rect 2807 1687 2808 1688
rect 2812 1687 2813 1691
rect 2807 1686 2813 1687
rect 2830 1691 2836 1692
rect 2830 1687 2831 1691
rect 2835 1690 2836 1691
rect 2895 1691 2901 1692
rect 2895 1690 2896 1691
rect 2835 1688 2896 1690
rect 2835 1687 2836 1688
rect 2830 1686 2836 1687
rect 2895 1687 2896 1688
rect 2900 1687 2901 1691
rect 2895 1686 2901 1687
rect 2839 1683 2845 1684
rect 2839 1682 2840 1683
rect 2696 1680 2840 1682
rect 2446 1678 2452 1679
rect 2839 1679 2840 1680
rect 2844 1679 2845 1683
rect 2839 1678 2845 1679
rect 2156 1672 2170 1674
rect 2174 1675 2180 1676
rect 2156 1671 2157 1672
rect 2151 1670 2157 1671
rect 2174 1671 2175 1675
rect 2179 1674 2180 1675
rect 2239 1675 2245 1676
rect 2239 1674 2240 1675
rect 2179 1672 2240 1674
rect 2179 1671 2180 1672
rect 2174 1670 2180 1671
rect 2239 1671 2240 1672
rect 2244 1671 2245 1675
rect 2239 1670 2245 1671
rect 2262 1675 2268 1676
rect 2262 1671 2263 1675
rect 2267 1674 2268 1675
rect 2327 1675 2333 1676
rect 2327 1674 2328 1675
rect 2267 1672 2328 1674
rect 2267 1671 2268 1672
rect 2262 1670 2268 1671
rect 2327 1671 2328 1672
rect 2332 1671 2333 1675
rect 2327 1670 2333 1671
rect 2350 1675 2356 1676
rect 2350 1671 2351 1675
rect 2355 1674 2356 1675
rect 2415 1675 2421 1676
rect 2415 1674 2416 1675
rect 2355 1672 2416 1674
rect 2355 1671 2356 1672
rect 2350 1670 2356 1671
rect 2415 1671 2416 1672
rect 2420 1671 2421 1675
rect 2415 1670 2421 1671
rect 2438 1675 2444 1676
rect 2438 1671 2439 1675
rect 2443 1674 2444 1675
rect 2503 1675 2509 1676
rect 2503 1674 2504 1675
rect 2443 1672 2504 1674
rect 2443 1671 2444 1672
rect 2438 1670 2444 1671
rect 2503 1671 2504 1672
rect 2508 1671 2509 1675
rect 2503 1670 2509 1671
rect 2591 1675 2597 1676
rect 2591 1671 2592 1675
rect 2596 1674 2597 1675
rect 2646 1675 2652 1676
rect 2646 1674 2647 1675
rect 2596 1672 2647 1674
rect 2596 1671 2597 1672
rect 2591 1670 2597 1671
rect 2646 1671 2647 1672
rect 2651 1671 2652 1675
rect 2679 1675 2685 1676
rect 2679 1674 2680 1675
rect 2646 1670 2652 1671
rect 2656 1672 2680 1674
rect 480 1668 514 1670
rect 656 1668 682 1670
rect 110 1664 116 1665
rect 110 1660 111 1664
rect 115 1660 116 1664
rect 110 1659 116 1660
rect 398 1663 404 1664
rect 398 1659 399 1663
rect 403 1659 404 1663
rect 398 1658 404 1659
rect 480 1654 482 1668
rect 486 1663 492 1664
rect 486 1659 487 1663
rect 491 1659 492 1663
rect 486 1658 492 1659
rect 574 1663 580 1664
rect 574 1659 575 1663
rect 579 1659 580 1663
rect 574 1658 580 1659
rect 656 1654 658 1668
rect 2656 1666 2658 1672
rect 2679 1671 2680 1672
rect 2684 1671 2685 1675
rect 2679 1670 2685 1671
rect 2702 1675 2708 1676
rect 2702 1671 2703 1675
rect 2707 1674 2708 1675
rect 2767 1675 2773 1676
rect 2767 1674 2768 1675
rect 2707 1672 2768 1674
rect 2707 1671 2708 1672
rect 2702 1670 2708 1671
rect 2767 1671 2768 1672
rect 2772 1671 2773 1675
rect 2767 1670 2773 1671
rect 2790 1675 2796 1676
rect 2790 1671 2791 1675
rect 2795 1674 2796 1675
rect 2855 1675 2861 1676
rect 2855 1674 2856 1675
rect 2795 1672 2856 1674
rect 2795 1671 2796 1672
rect 2790 1670 2796 1671
rect 2855 1671 2856 1672
rect 2860 1671 2861 1675
rect 2855 1670 2861 1671
rect 2878 1675 2884 1676
rect 2878 1671 2879 1675
rect 2883 1674 2884 1675
rect 2943 1675 2949 1676
rect 2943 1674 2944 1675
rect 2883 1672 2944 1674
rect 2883 1671 2884 1672
rect 2878 1670 2884 1671
rect 2943 1671 2944 1672
rect 2948 1671 2949 1675
rect 2943 1670 2949 1671
rect 1766 1664 1772 1665
rect 662 1663 668 1664
rect 662 1659 663 1663
rect 667 1659 668 1663
rect 662 1658 668 1659
rect 758 1663 764 1664
rect 758 1659 759 1663
rect 763 1659 764 1663
rect 758 1658 764 1659
rect 854 1663 860 1664
rect 854 1659 855 1663
rect 859 1659 860 1663
rect 854 1658 860 1659
rect 950 1663 956 1664
rect 950 1659 951 1663
rect 955 1659 956 1663
rect 950 1658 956 1659
rect 1046 1663 1052 1664
rect 1046 1659 1047 1663
rect 1051 1659 1052 1663
rect 1046 1658 1052 1659
rect 1142 1663 1148 1664
rect 1142 1659 1143 1663
rect 1147 1659 1148 1663
rect 1766 1660 1767 1664
rect 1771 1660 1772 1664
rect 2624 1664 2658 1666
rect 1766 1659 1772 1660
rect 1806 1660 1812 1661
rect 1142 1658 1148 1659
rect 1806 1656 1807 1660
rect 1811 1656 1812 1660
rect 473 1652 482 1654
rect 649 1652 658 1654
rect 734 1655 740 1656
rect 558 1651 564 1652
rect 110 1647 116 1648
rect 110 1643 111 1647
rect 115 1643 116 1647
rect 558 1647 559 1651
rect 563 1647 564 1651
rect 734 1651 735 1655
rect 739 1651 740 1655
rect 734 1650 740 1651
rect 838 1655 844 1656
rect 838 1651 839 1655
rect 843 1654 844 1655
rect 943 1655 949 1656
rect 843 1652 897 1654
rect 843 1651 844 1652
rect 838 1650 844 1651
rect 943 1651 944 1655
rect 948 1654 949 1655
rect 1118 1655 1124 1656
rect 948 1652 993 1654
rect 948 1651 949 1652
rect 943 1650 949 1651
rect 1118 1651 1119 1655
rect 1123 1651 1124 1655
rect 1118 1650 1124 1651
rect 1126 1655 1132 1656
rect 1806 1655 1812 1656
rect 2102 1659 2108 1660
rect 2102 1655 2103 1659
rect 2107 1655 2108 1659
rect 1126 1651 1127 1655
rect 1131 1654 1132 1655
rect 2102 1654 2108 1655
rect 2190 1659 2196 1660
rect 2190 1655 2191 1659
rect 2195 1655 2196 1659
rect 2190 1654 2196 1655
rect 2278 1659 2284 1660
rect 2278 1655 2279 1659
rect 2283 1655 2284 1659
rect 2278 1654 2284 1655
rect 2366 1659 2372 1660
rect 2366 1655 2367 1659
rect 2371 1655 2372 1659
rect 2366 1654 2372 1655
rect 2454 1659 2460 1660
rect 2454 1655 2455 1659
rect 2459 1655 2460 1659
rect 2454 1654 2460 1655
rect 2542 1659 2548 1660
rect 2542 1655 2543 1659
rect 2547 1655 2548 1659
rect 2542 1654 2548 1655
rect 1131 1652 1185 1654
rect 1131 1651 1132 1652
rect 1126 1650 1132 1651
rect 2174 1651 2180 1652
rect 558 1646 564 1647
rect 832 1646 834 1649
rect 838 1647 844 1648
rect 838 1646 839 1647
rect 110 1642 116 1643
rect 398 1644 404 1645
rect 398 1640 399 1644
rect 403 1640 404 1644
rect 398 1639 404 1640
rect 486 1644 492 1645
rect 486 1640 487 1644
rect 491 1640 492 1644
rect 486 1639 492 1640
rect 574 1644 580 1645
rect 574 1640 575 1644
rect 579 1640 580 1644
rect 574 1639 580 1640
rect 662 1644 668 1645
rect 662 1640 663 1644
rect 667 1640 668 1644
rect 662 1639 668 1640
rect 758 1644 764 1645
rect 832 1644 839 1646
rect 758 1640 759 1644
rect 763 1640 764 1644
rect 838 1643 839 1644
rect 843 1643 844 1647
rect 1766 1647 1772 1648
rect 838 1642 844 1643
rect 854 1644 860 1645
rect 758 1639 764 1640
rect 854 1640 855 1644
rect 859 1640 860 1644
rect 854 1639 860 1640
rect 950 1644 956 1645
rect 950 1640 951 1644
rect 955 1640 956 1644
rect 950 1639 956 1640
rect 1046 1644 1052 1645
rect 1046 1640 1047 1644
rect 1051 1640 1052 1644
rect 1046 1639 1052 1640
rect 1142 1644 1148 1645
rect 1142 1640 1143 1644
rect 1147 1640 1148 1644
rect 1766 1643 1767 1647
rect 1771 1643 1772 1647
rect 2174 1647 2175 1651
rect 2179 1647 2180 1651
rect 2174 1646 2180 1647
rect 2262 1651 2268 1652
rect 2262 1647 2263 1651
rect 2267 1647 2268 1651
rect 2262 1646 2268 1647
rect 2350 1651 2356 1652
rect 2350 1647 2351 1651
rect 2355 1647 2356 1651
rect 2350 1646 2356 1647
rect 2438 1651 2444 1652
rect 2438 1647 2439 1651
rect 2443 1647 2444 1651
rect 2438 1646 2444 1647
rect 2526 1651 2532 1652
rect 2526 1647 2527 1651
rect 2531 1647 2532 1651
rect 2624 1650 2626 1664
rect 3462 1660 3468 1661
rect 2630 1659 2636 1660
rect 2630 1655 2631 1659
rect 2635 1655 2636 1659
rect 2630 1654 2636 1655
rect 2718 1659 2724 1660
rect 2718 1655 2719 1659
rect 2723 1655 2724 1659
rect 2718 1654 2724 1655
rect 2806 1659 2812 1660
rect 2806 1655 2807 1659
rect 2811 1655 2812 1659
rect 2806 1654 2812 1655
rect 2894 1659 2900 1660
rect 2894 1655 2895 1659
rect 2899 1655 2900 1659
rect 3462 1656 3463 1660
rect 3467 1656 3468 1660
rect 3462 1655 3468 1656
rect 2894 1654 2900 1655
rect 2617 1648 2626 1650
rect 2702 1651 2708 1652
rect 2526 1646 2532 1647
rect 2702 1647 2703 1651
rect 2707 1647 2708 1651
rect 2702 1646 2708 1647
rect 2790 1651 2796 1652
rect 2790 1647 2791 1651
rect 2795 1647 2796 1651
rect 2790 1646 2796 1647
rect 2878 1651 2884 1652
rect 2878 1647 2879 1651
rect 2883 1647 2884 1651
rect 2878 1646 2884 1647
rect 2887 1651 2893 1652
rect 2887 1647 2888 1651
rect 2892 1650 2893 1651
rect 2892 1648 2937 1650
rect 2892 1647 2893 1648
rect 2887 1646 2893 1647
rect 1766 1642 1772 1643
rect 1806 1643 1812 1644
rect 1142 1639 1148 1640
rect 1806 1639 1807 1643
rect 1811 1639 1812 1643
rect 3462 1643 3468 1644
rect 1806 1638 1812 1639
rect 2102 1640 2108 1641
rect 2102 1636 2103 1640
rect 2107 1636 2108 1640
rect 2102 1635 2108 1636
rect 2190 1640 2196 1641
rect 2190 1636 2191 1640
rect 2195 1636 2196 1640
rect 2190 1635 2196 1636
rect 2278 1640 2284 1641
rect 2278 1636 2279 1640
rect 2283 1636 2284 1640
rect 2278 1635 2284 1636
rect 2366 1640 2372 1641
rect 2366 1636 2367 1640
rect 2371 1636 2372 1640
rect 2366 1635 2372 1636
rect 2454 1640 2460 1641
rect 2454 1636 2455 1640
rect 2459 1636 2460 1640
rect 2454 1635 2460 1636
rect 2542 1640 2548 1641
rect 2542 1636 2543 1640
rect 2547 1636 2548 1640
rect 2542 1635 2548 1636
rect 2630 1640 2636 1641
rect 2630 1636 2631 1640
rect 2635 1636 2636 1640
rect 2630 1635 2636 1636
rect 2718 1640 2724 1641
rect 2718 1636 2719 1640
rect 2723 1636 2724 1640
rect 2718 1635 2724 1636
rect 2806 1640 2812 1641
rect 2806 1636 2807 1640
rect 2811 1636 2812 1640
rect 2806 1635 2812 1636
rect 2894 1640 2900 1641
rect 2894 1636 2895 1640
rect 2899 1636 2900 1640
rect 3462 1639 3463 1643
rect 3467 1639 3468 1643
rect 3462 1638 3468 1639
rect 2894 1635 2900 1636
rect 2618 1607 2624 1608
rect 2618 1603 2619 1607
rect 2623 1606 2624 1607
rect 2887 1607 2893 1608
rect 2887 1606 2888 1607
rect 2623 1604 2888 1606
rect 2623 1603 2624 1604
rect 2618 1602 2624 1603
rect 2887 1603 2888 1604
rect 2892 1603 2893 1607
rect 2887 1602 2893 1603
rect 2602 1599 2608 1600
rect 278 1596 284 1597
rect 110 1593 116 1594
rect 110 1589 111 1593
rect 115 1589 116 1593
rect 278 1592 279 1596
rect 283 1592 284 1596
rect 278 1591 284 1592
rect 382 1596 388 1597
rect 382 1592 383 1596
rect 387 1592 388 1596
rect 382 1591 388 1592
rect 494 1596 500 1597
rect 494 1592 495 1596
rect 499 1592 500 1596
rect 494 1591 500 1592
rect 606 1596 612 1597
rect 606 1592 607 1596
rect 611 1592 612 1596
rect 606 1591 612 1592
rect 718 1596 724 1597
rect 718 1592 719 1596
rect 723 1592 724 1596
rect 718 1591 724 1592
rect 830 1596 836 1597
rect 830 1592 831 1596
rect 835 1592 836 1596
rect 830 1591 836 1592
rect 942 1596 948 1597
rect 942 1592 943 1596
rect 947 1592 948 1596
rect 942 1591 948 1592
rect 1054 1596 1060 1597
rect 1054 1592 1055 1596
rect 1059 1592 1060 1596
rect 1054 1591 1060 1592
rect 1166 1596 1172 1597
rect 1166 1592 1167 1596
rect 1171 1592 1172 1596
rect 1166 1591 1172 1592
rect 1278 1596 1284 1597
rect 1278 1592 1279 1596
rect 1283 1592 1284 1596
rect 2602 1595 2603 1599
rect 2607 1598 2608 1599
rect 2607 1596 2882 1598
rect 2607 1595 2608 1596
rect 2602 1594 2608 1595
rect 1278 1591 1284 1592
rect 1766 1593 1772 1594
rect 110 1588 116 1589
rect 1766 1589 1767 1593
rect 1771 1589 1772 1593
rect 2062 1592 2068 1593
rect 1766 1588 1772 1589
rect 1806 1589 1812 1590
rect 350 1587 356 1588
rect 350 1583 351 1587
rect 355 1583 356 1587
rect 350 1582 356 1583
rect 454 1587 460 1588
rect 454 1583 455 1587
rect 459 1583 460 1587
rect 454 1582 460 1583
rect 462 1587 468 1588
rect 462 1583 463 1587
rect 467 1586 468 1587
rect 670 1587 676 1588
rect 467 1584 537 1586
rect 467 1583 468 1584
rect 462 1582 468 1583
rect 670 1583 671 1587
rect 675 1583 676 1587
rect 670 1582 676 1583
rect 686 1587 692 1588
rect 686 1583 687 1587
rect 691 1586 692 1587
rect 902 1587 908 1588
rect 691 1584 761 1586
rect 691 1583 692 1584
rect 686 1582 692 1583
rect 902 1583 903 1587
rect 907 1583 908 1587
rect 902 1582 908 1583
rect 1014 1587 1020 1588
rect 1014 1583 1015 1587
rect 1019 1583 1020 1587
rect 1014 1582 1020 1583
rect 1126 1587 1132 1588
rect 1126 1583 1127 1587
rect 1131 1583 1132 1587
rect 1126 1582 1132 1583
rect 1238 1587 1244 1588
rect 1238 1583 1239 1587
rect 1243 1583 1244 1587
rect 1238 1582 1244 1583
rect 1246 1587 1252 1588
rect 1246 1583 1247 1587
rect 1251 1586 1252 1587
rect 1251 1584 1321 1586
rect 1806 1585 1807 1589
rect 1811 1585 1812 1589
rect 2062 1588 2063 1592
rect 2067 1588 2068 1592
rect 2062 1587 2068 1588
rect 2158 1592 2164 1593
rect 2158 1588 2159 1592
rect 2163 1588 2164 1592
rect 2158 1587 2164 1588
rect 2254 1592 2260 1593
rect 2254 1588 2255 1592
rect 2259 1588 2260 1592
rect 2254 1587 2260 1588
rect 2358 1592 2364 1593
rect 2358 1588 2359 1592
rect 2363 1588 2364 1592
rect 2358 1587 2364 1588
rect 2462 1592 2468 1593
rect 2462 1588 2463 1592
rect 2467 1588 2468 1592
rect 2462 1587 2468 1588
rect 2566 1592 2572 1593
rect 2566 1588 2567 1592
rect 2571 1588 2572 1592
rect 2566 1587 2572 1588
rect 2670 1592 2676 1593
rect 2670 1588 2671 1592
rect 2675 1588 2676 1592
rect 2670 1587 2676 1588
rect 2774 1592 2780 1593
rect 2774 1588 2775 1592
rect 2779 1588 2780 1592
rect 2774 1587 2780 1588
rect 1806 1584 1812 1585
rect 1251 1583 1252 1584
rect 1246 1582 1252 1583
rect 2134 1583 2140 1584
rect 2134 1579 2135 1583
rect 2139 1579 2140 1583
rect 2134 1578 2140 1579
rect 2230 1583 2236 1584
rect 2230 1579 2231 1583
rect 2235 1579 2236 1583
rect 2230 1578 2236 1579
rect 2326 1583 2332 1584
rect 2326 1579 2327 1583
rect 2331 1579 2332 1583
rect 2326 1578 2332 1579
rect 2430 1583 2436 1584
rect 2430 1579 2431 1583
rect 2435 1579 2436 1583
rect 2430 1578 2436 1579
rect 2446 1583 2452 1584
rect 2446 1579 2447 1583
rect 2451 1582 2452 1583
rect 2638 1583 2644 1584
rect 2451 1580 2505 1582
rect 2451 1579 2452 1580
rect 2446 1578 2452 1579
rect 2638 1579 2639 1583
rect 2643 1579 2644 1583
rect 2638 1578 2644 1579
rect 2742 1583 2748 1584
rect 2742 1579 2743 1583
rect 2747 1579 2748 1583
rect 2742 1578 2748 1579
rect 2846 1583 2852 1584
rect 2846 1579 2847 1583
rect 2851 1579 2852 1583
rect 2880 1582 2882 1596
rect 2886 1592 2892 1593
rect 2886 1588 2887 1592
rect 2891 1588 2892 1592
rect 2886 1587 2892 1588
rect 3462 1589 3468 1590
rect 3462 1585 3463 1589
rect 3467 1585 3468 1589
rect 3462 1584 3468 1585
rect 2880 1580 2929 1582
rect 2846 1578 2852 1579
rect 278 1577 284 1578
rect 110 1576 116 1577
rect 110 1572 111 1576
rect 115 1572 116 1576
rect 278 1573 279 1577
rect 283 1573 284 1577
rect 278 1572 284 1573
rect 382 1577 388 1578
rect 382 1573 383 1577
rect 387 1573 388 1577
rect 382 1572 388 1573
rect 494 1577 500 1578
rect 494 1573 495 1577
rect 499 1573 500 1577
rect 494 1572 500 1573
rect 606 1577 612 1578
rect 606 1573 607 1577
rect 611 1573 612 1577
rect 606 1572 612 1573
rect 718 1577 724 1578
rect 718 1573 719 1577
rect 723 1573 724 1577
rect 718 1572 724 1573
rect 830 1577 836 1578
rect 830 1573 831 1577
rect 835 1573 836 1577
rect 830 1572 836 1573
rect 942 1577 948 1578
rect 942 1573 943 1577
rect 947 1573 948 1577
rect 942 1572 948 1573
rect 1054 1577 1060 1578
rect 1054 1573 1055 1577
rect 1059 1573 1060 1577
rect 1054 1572 1060 1573
rect 1166 1577 1172 1578
rect 1166 1573 1167 1577
rect 1171 1573 1172 1577
rect 1166 1572 1172 1573
rect 1278 1577 1284 1578
rect 1278 1573 1279 1577
rect 1283 1573 1284 1577
rect 1278 1572 1284 1573
rect 1766 1576 1772 1577
rect 1766 1572 1767 1576
rect 1771 1572 1772 1576
rect 2062 1573 2068 1574
rect 110 1571 116 1572
rect 1766 1571 1772 1572
rect 1806 1572 1812 1573
rect 1806 1568 1807 1572
rect 1811 1568 1812 1572
rect 2062 1569 2063 1573
rect 2067 1569 2068 1573
rect 2062 1568 2068 1569
rect 2158 1573 2164 1574
rect 2158 1569 2159 1573
rect 2163 1569 2164 1573
rect 2158 1568 2164 1569
rect 2254 1573 2260 1574
rect 2254 1569 2255 1573
rect 2259 1569 2260 1573
rect 2254 1568 2260 1569
rect 2358 1573 2364 1574
rect 2358 1569 2359 1573
rect 2363 1569 2364 1573
rect 2358 1568 2364 1569
rect 2462 1573 2468 1574
rect 2462 1569 2463 1573
rect 2467 1569 2468 1573
rect 2462 1568 2468 1569
rect 2566 1573 2572 1574
rect 2566 1569 2567 1573
rect 2571 1569 2572 1573
rect 2566 1568 2572 1569
rect 2670 1573 2676 1574
rect 2670 1569 2671 1573
rect 2675 1569 2676 1573
rect 2670 1568 2676 1569
rect 2774 1573 2780 1574
rect 2774 1569 2775 1573
rect 2779 1569 2780 1573
rect 2774 1568 2780 1569
rect 2886 1573 2892 1574
rect 2886 1569 2887 1573
rect 2891 1569 2892 1573
rect 2886 1568 2892 1569
rect 3462 1572 3468 1573
rect 3462 1568 3463 1572
rect 3467 1568 3468 1572
rect 1806 1567 1812 1568
rect 3462 1567 3468 1568
rect 327 1559 333 1560
rect 327 1555 328 1559
rect 332 1558 333 1559
rect 350 1559 356 1560
rect 332 1556 346 1558
rect 332 1555 333 1556
rect 327 1554 333 1555
rect 344 1550 346 1556
rect 350 1555 351 1559
rect 355 1558 356 1559
rect 431 1559 437 1560
rect 431 1558 432 1559
rect 355 1556 432 1558
rect 355 1555 356 1556
rect 350 1554 356 1555
rect 431 1555 432 1556
rect 436 1555 437 1559
rect 431 1554 437 1555
rect 543 1559 549 1560
rect 543 1555 544 1559
rect 548 1558 549 1559
rect 558 1559 564 1560
rect 558 1558 559 1559
rect 548 1556 559 1558
rect 548 1555 549 1556
rect 543 1554 549 1555
rect 558 1555 559 1556
rect 563 1555 564 1559
rect 558 1554 564 1555
rect 655 1559 661 1560
rect 655 1555 656 1559
rect 660 1558 661 1559
rect 686 1559 692 1560
rect 686 1558 687 1559
rect 660 1556 687 1558
rect 660 1555 661 1556
rect 655 1554 661 1555
rect 686 1555 687 1556
rect 691 1555 692 1559
rect 686 1554 692 1555
rect 694 1559 700 1560
rect 694 1555 695 1559
rect 699 1558 700 1559
rect 767 1559 773 1560
rect 767 1558 768 1559
rect 699 1556 768 1558
rect 699 1555 700 1556
rect 694 1554 700 1555
rect 767 1555 768 1556
rect 772 1555 773 1559
rect 767 1554 773 1555
rect 838 1559 844 1560
rect 838 1555 839 1559
rect 843 1558 844 1559
rect 879 1559 885 1560
rect 879 1558 880 1559
rect 843 1556 880 1558
rect 843 1555 844 1556
rect 838 1554 844 1555
rect 879 1555 880 1556
rect 884 1555 885 1559
rect 879 1554 885 1555
rect 902 1559 908 1560
rect 902 1555 903 1559
rect 907 1558 908 1559
rect 991 1559 997 1560
rect 991 1558 992 1559
rect 907 1556 992 1558
rect 907 1555 908 1556
rect 902 1554 908 1555
rect 991 1555 992 1556
rect 996 1555 997 1559
rect 991 1554 997 1555
rect 1014 1559 1020 1560
rect 1014 1555 1015 1559
rect 1019 1558 1020 1559
rect 1103 1559 1109 1560
rect 1103 1558 1104 1559
rect 1019 1556 1104 1558
rect 1019 1555 1020 1556
rect 1014 1554 1020 1555
rect 1103 1555 1104 1556
rect 1108 1555 1109 1559
rect 1103 1554 1109 1555
rect 1126 1559 1132 1560
rect 1126 1555 1127 1559
rect 1131 1558 1132 1559
rect 1215 1559 1221 1560
rect 1215 1558 1216 1559
rect 1131 1556 1216 1558
rect 1131 1555 1132 1556
rect 1126 1554 1132 1555
rect 1215 1555 1216 1556
rect 1220 1555 1221 1559
rect 1215 1554 1221 1555
rect 1238 1559 1244 1560
rect 1238 1555 1239 1559
rect 1243 1558 1244 1559
rect 1327 1559 1333 1560
rect 1327 1558 1328 1559
rect 1243 1556 1328 1558
rect 1243 1555 1244 1556
rect 1238 1554 1244 1555
rect 1327 1555 1328 1556
rect 1332 1555 1333 1559
rect 1327 1554 1333 1555
rect 2110 1555 2117 1556
rect 462 1551 468 1552
rect 462 1550 463 1551
rect 344 1548 463 1550
rect 462 1547 463 1548
rect 467 1547 468 1551
rect 2110 1551 2111 1555
rect 2116 1551 2117 1555
rect 2110 1550 2117 1551
rect 2134 1555 2140 1556
rect 2134 1551 2135 1555
rect 2139 1554 2140 1555
rect 2207 1555 2213 1556
rect 2207 1554 2208 1555
rect 2139 1552 2208 1554
rect 2139 1551 2140 1552
rect 2134 1550 2140 1551
rect 2207 1551 2208 1552
rect 2212 1551 2213 1555
rect 2207 1550 2213 1551
rect 2230 1555 2236 1556
rect 2230 1551 2231 1555
rect 2235 1554 2236 1555
rect 2303 1555 2309 1556
rect 2303 1554 2304 1555
rect 2235 1552 2304 1554
rect 2235 1551 2236 1552
rect 2230 1550 2236 1551
rect 2303 1551 2304 1552
rect 2308 1551 2309 1555
rect 2303 1550 2309 1551
rect 2326 1555 2332 1556
rect 2326 1551 2327 1555
rect 2331 1554 2332 1555
rect 2407 1555 2413 1556
rect 2407 1554 2408 1555
rect 2331 1552 2408 1554
rect 2331 1551 2332 1552
rect 2326 1550 2332 1551
rect 2407 1551 2408 1552
rect 2412 1551 2413 1555
rect 2407 1550 2413 1551
rect 2430 1555 2436 1556
rect 2430 1551 2431 1555
rect 2435 1554 2436 1555
rect 2511 1555 2517 1556
rect 2511 1554 2512 1555
rect 2435 1552 2512 1554
rect 2435 1551 2436 1552
rect 2430 1550 2436 1551
rect 2511 1551 2512 1552
rect 2516 1551 2517 1555
rect 2511 1550 2517 1551
rect 2615 1555 2624 1556
rect 2615 1551 2616 1555
rect 2623 1551 2624 1555
rect 2615 1550 2624 1551
rect 2638 1555 2644 1556
rect 2638 1551 2639 1555
rect 2643 1554 2644 1555
rect 2719 1555 2725 1556
rect 2719 1554 2720 1555
rect 2643 1552 2720 1554
rect 2643 1551 2644 1552
rect 2638 1550 2644 1551
rect 2719 1551 2720 1552
rect 2724 1551 2725 1555
rect 2719 1550 2725 1551
rect 2742 1555 2748 1556
rect 2742 1551 2743 1555
rect 2747 1554 2748 1555
rect 2823 1555 2829 1556
rect 2823 1554 2824 1555
rect 2747 1552 2824 1554
rect 2747 1551 2748 1552
rect 2742 1550 2748 1551
rect 2823 1551 2824 1552
rect 2828 1551 2829 1555
rect 2823 1550 2829 1551
rect 2846 1555 2852 1556
rect 2846 1551 2847 1555
rect 2851 1554 2852 1555
rect 2935 1555 2941 1556
rect 2935 1554 2936 1555
rect 2851 1552 2936 1554
rect 2851 1551 2852 1552
rect 2846 1550 2852 1551
rect 2935 1551 2936 1552
rect 2940 1551 2941 1555
rect 2935 1550 2941 1551
rect 462 1546 468 1547
rect 1246 1547 1252 1548
rect 1246 1546 1247 1547
rect 1060 1544 1247 1546
rect 231 1539 237 1540
rect 231 1535 232 1539
rect 236 1538 237 1539
rect 290 1539 296 1540
rect 290 1538 291 1539
rect 236 1536 291 1538
rect 236 1535 237 1536
rect 231 1534 237 1535
rect 290 1535 291 1536
rect 295 1535 296 1539
rect 290 1534 296 1535
rect 375 1539 381 1540
rect 375 1535 376 1539
rect 380 1538 381 1539
rect 406 1539 412 1540
rect 406 1538 407 1539
rect 380 1536 407 1538
rect 380 1535 381 1536
rect 375 1534 381 1535
rect 406 1535 407 1536
rect 411 1535 412 1539
rect 406 1534 412 1535
rect 454 1539 460 1540
rect 454 1535 455 1539
rect 459 1538 460 1539
rect 519 1539 525 1540
rect 519 1538 520 1539
rect 459 1536 520 1538
rect 459 1535 460 1536
rect 454 1534 460 1535
rect 519 1535 520 1536
rect 524 1535 525 1539
rect 519 1534 525 1535
rect 671 1539 677 1540
rect 671 1535 672 1539
rect 676 1538 677 1539
rect 702 1539 708 1540
rect 702 1538 703 1539
rect 676 1536 703 1538
rect 676 1535 677 1536
rect 671 1534 677 1535
rect 702 1535 703 1536
rect 707 1535 708 1539
rect 702 1534 708 1535
rect 815 1539 821 1540
rect 815 1535 816 1539
rect 820 1538 821 1539
rect 846 1539 852 1540
rect 846 1538 847 1539
rect 820 1536 847 1538
rect 820 1535 821 1536
rect 815 1534 821 1535
rect 846 1535 847 1536
rect 851 1535 852 1539
rect 846 1534 852 1535
rect 959 1539 965 1540
rect 959 1535 960 1539
rect 964 1538 965 1539
rect 1060 1538 1062 1544
rect 1246 1543 1247 1544
rect 1251 1543 1252 1547
rect 1246 1542 1252 1543
rect 1967 1543 1973 1544
rect 1095 1539 1101 1540
rect 1095 1538 1096 1539
rect 964 1536 1062 1538
rect 1064 1536 1096 1538
rect 964 1535 965 1536
rect 959 1534 965 1535
rect 1064 1530 1066 1536
rect 1095 1535 1096 1536
rect 1100 1535 1101 1539
rect 1095 1534 1101 1535
rect 1118 1539 1124 1540
rect 1118 1535 1119 1539
rect 1123 1538 1124 1539
rect 1223 1539 1229 1540
rect 1223 1538 1224 1539
rect 1123 1536 1224 1538
rect 1123 1535 1124 1536
rect 1118 1534 1124 1535
rect 1223 1535 1224 1536
rect 1228 1535 1229 1539
rect 1223 1534 1229 1535
rect 1246 1539 1252 1540
rect 1246 1535 1247 1539
rect 1251 1538 1252 1539
rect 1359 1539 1365 1540
rect 1359 1538 1360 1539
rect 1251 1536 1360 1538
rect 1251 1535 1252 1536
rect 1246 1534 1252 1535
rect 1359 1535 1360 1536
rect 1364 1535 1365 1539
rect 1359 1534 1365 1535
rect 1382 1539 1388 1540
rect 1382 1535 1383 1539
rect 1387 1538 1388 1539
rect 1495 1539 1501 1540
rect 1495 1538 1496 1539
rect 1387 1536 1496 1538
rect 1387 1535 1388 1536
rect 1382 1534 1388 1535
rect 1495 1535 1496 1536
rect 1500 1535 1501 1539
rect 1967 1539 1968 1543
rect 1972 1542 1973 1543
rect 1982 1543 1988 1544
rect 1982 1542 1983 1543
rect 1972 1540 1983 1542
rect 1972 1539 1973 1540
rect 1967 1538 1973 1539
rect 1982 1539 1983 1540
rect 1987 1539 1988 1543
rect 1982 1538 1988 1539
rect 1990 1543 1996 1544
rect 1990 1539 1991 1543
rect 1995 1542 1996 1543
rect 2087 1543 2093 1544
rect 2087 1542 2088 1543
rect 1995 1540 2088 1542
rect 1995 1539 1996 1540
rect 1990 1538 1996 1539
rect 2087 1539 2088 1540
rect 2092 1539 2093 1543
rect 2087 1538 2093 1539
rect 2110 1543 2116 1544
rect 2110 1539 2111 1543
rect 2115 1542 2116 1543
rect 2215 1543 2221 1544
rect 2215 1542 2216 1543
rect 2115 1540 2216 1542
rect 2115 1539 2116 1540
rect 2110 1538 2116 1539
rect 2215 1539 2216 1540
rect 2220 1539 2221 1543
rect 2215 1538 2221 1539
rect 2238 1543 2244 1544
rect 2238 1539 2239 1543
rect 2243 1542 2244 1543
rect 2343 1543 2349 1544
rect 2343 1542 2344 1543
rect 2243 1540 2344 1542
rect 2243 1539 2244 1540
rect 2238 1538 2244 1539
rect 2343 1539 2344 1540
rect 2348 1539 2349 1543
rect 2343 1538 2349 1539
rect 2366 1543 2372 1544
rect 2366 1539 2367 1543
rect 2371 1542 2372 1543
rect 2471 1543 2477 1544
rect 2471 1542 2472 1543
rect 2371 1540 2472 1542
rect 2371 1539 2372 1540
rect 2366 1538 2372 1539
rect 2471 1539 2472 1540
rect 2476 1539 2477 1543
rect 2471 1538 2477 1539
rect 2599 1543 2608 1544
rect 2599 1539 2600 1543
rect 2607 1539 2608 1543
rect 2599 1538 2608 1539
rect 2622 1543 2628 1544
rect 2622 1539 2623 1543
rect 2627 1542 2628 1543
rect 2727 1543 2733 1544
rect 2727 1542 2728 1543
rect 2627 1540 2728 1542
rect 2627 1539 2628 1540
rect 2622 1538 2628 1539
rect 2727 1539 2728 1540
rect 2732 1539 2733 1543
rect 2727 1538 2733 1539
rect 2750 1543 2756 1544
rect 2750 1539 2751 1543
rect 2755 1542 2756 1543
rect 2847 1543 2853 1544
rect 2847 1542 2848 1543
rect 2755 1540 2848 1542
rect 2755 1539 2756 1540
rect 2750 1538 2756 1539
rect 2847 1539 2848 1540
rect 2852 1539 2853 1543
rect 2847 1538 2853 1539
rect 2870 1543 2876 1544
rect 2870 1539 2871 1543
rect 2875 1542 2876 1543
rect 2975 1543 2981 1544
rect 2975 1542 2976 1543
rect 2875 1540 2976 1542
rect 2875 1539 2876 1540
rect 2870 1538 2876 1539
rect 2975 1539 2976 1540
rect 2980 1539 2981 1543
rect 2975 1538 2981 1539
rect 2998 1543 3004 1544
rect 2998 1539 2999 1543
rect 3003 1542 3004 1543
rect 3103 1543 3109 1544
rect 3103 1542 3104 1543
rect 3003 1540 3104 1542
rect 3003 1539 3004 1540
rect 2998 1538 3004 1539
rect 3103 1539 3104 1540
rect 3108 1539 3109 1543
rect 3103 1538 3109 1539
rect 1495 1534 1501 1535
rect 1028 1528 1066 1530
rect 1806 1528 1812 1529
rect 3462 1528 3468 1529
rect 110 1524 116 1525
rect 110 1520 111 1524
rect 115 1520 116 1524
rect 110 1519 116 1520
rect 182 1523 188 1524
rect 182 1519 183 1523
rect 187 1519 188 1523
rect 182 1518 188 1519
rect 326 1523 332 1524
rect 326 1519 327 1523
rect 331 1519 332 1523
rect 326 1518 332 1519
rect 470 1523 476 1524
rect 470 1519 471 1523
rect 475 1519 476 1523
rect 470 1518 476 1519
rect 622 1523 628 1524
rect 622 1519 623 1523
rect 627 1519 628 1523
rect 622 1518 628 1519
rect 766 1523 772 1524
rect 766 1519 767 1523
rect 771 1519 772 1523
rect 766 1518 772 1519
rect 910 1523 916 1524
rect 910 1519 911 1523
rect 915 1519 916 1523
rect 910 1518 916 1519
rect 290 1515 296 1516
rect 254 1511 260 1512
rect 110 1507 116 1508
rect 110 1503 111 1507
rect 115 1503 116 1507
rect 254 1507 255 1511
rect 259 1507 260 1511
rect 290 1511 291 1515
rect 295 1514 296 1515
rect 406 1515 412 1516
rect 295 1512 369 1514
rect 295 1511 296 1512
rect 290 1510 296 1511
rect 406 1511 407 1515
rect 411 1514 412 1515
rect 694 1515 700 1516
rect 411 1512 513 1514
rect 411 1511 412 1512
rect 406 1510 412 1511
rect 694 1511 695 1515
rect 699 1511 700 1515
rect 694 1510 700 1511
rect 702 1515 708 1516
rect 702 1511 703 1515
rect 707 1514 708 1515
rect 1028 1514 1030 1528
rect 1766 1524 1772 1525
rect 1046 1523 1052 1524
rect 1046 1519 1047 1523
rect 1051 1519 1052 1523
rect 1046 1518 1052 1519
rect 1174 1523 1180 1524
rect 1174 1519 1175 1523
rect 1179 1519 1180 1523
rect 1174 1518 1180 1519
rect 1310 1523 1316 1524
rect 1310 1519 1311 1523
rect 1315 1519 1316 1523
rect 1310 1518 1316 1519
rect 1446 1523 1452 1524
rect 1446 1519 1447 1523
rect 1451 1519 1452 1523
rect 1766 1520 1767 1524
rect 1771 1520 1772 1524
rect 1806 1524 1807 1528
rect 1811 1524 1812 1528
rect 1806 1523 1812 1524
rect 1918 1527 1924 1528
rect 1918 1523 1919 1527
rect 1923 1523 1924 1527
rect 1918 1522 1924 1523
rect 2038 1527 2044 1528
rect 2038 1523 2039 1527
rect 2043 1523 2044 1527
rect 2038 1522 2044 1523
rect 2166 1527 2172 1528
rect 2166 1523 2167 1527
rect 2171 1523 2172 1527
rect 2166 1522 2172 1523
rect 2294 1527 2300 1528
rect 2294 1523 2295 1527
rect 2299 1523 2300 1527
rect 2294 1522 2300 1523
rect 2422 1527 2428 1528
rect 2422 1523 2423 1527
rect 2427 1523 2428 1527
rect 2422 1522 2428 1523
rect 2550 1527 2556 1528
rect 2550 1523 2551 1527
rect 2555 1523 2556 1527
rect 2550 1522 2556 1523
rect 2678 1527 2684 1528
rect 2678 1523 2679 1527
rect 2683 1523 2684 1527
rect 2678 1522 2684 1523
rect 2798 1527 2804 1528
rect 2798 1523 2799 1527
rect 2803 1523 2804 1527
rect 2798 1522 2804 1523
rect 2926 1527 2932 1528
rect 2926 1523 2927 1527
rect 2931 1523 2932 1527
rect 2926 1522 2932 1523
rect 3054 1527 3060 1528
rect 3054 1523 3055 1527
rect 3059 1523 3060 1527
rect 3462 1524 3463 1528
rect 3467 1524 3468 1528
rect 3462 1523 3468 1524
rect 3054 1522 3060 1523
rect 1766 1519 1772 1520
rect 1990 1519 1996 1520
rect 1446 1518 1452 1519
rect 707 1512 809 1514
rect 985 1512 1030 1514
rect 1118 1515 1124 1516
rect 707 1511 708 1512
rect 702 1510 708 1511
rect 1118 1511 1119 1515
rect 1123 1511 1124 1515
rect 1118 1510 1124 1511
rect 1246 1515 1252 1516
rect 1246 1511 1247 1515
rect 1251 1511 1252 1515
rect 1246 1510 1252 1511
rect 1382 1515 1388 1516
rect 1382 1511 1383 1515
rect 1387 1511 1388 1515
rect 1382 1510 1388 1511
rect 1398 1515 1404 1516
rect 1398 1511 1399 1515
rect 1403 1514 1404 1515
rect 1990 1515 1991 1519
rect 1995 1515 1996 1519
rect 1990 1514 1996 1515
rect 2110 1519 2116 1520
rect 2110 1515 2111 1519
rect 2115 1515 2116 1519
rect 2110 1514 2116 1515
rect 2238 1519 2244 1520
rect 2238 1515 2239 1519
rect 2243 1515 2244 1519
rect 2238 1514 2244 1515
rect 2366 1519 2372 1520
rect 2366 1515 2367 1519
rect 2371 1515 2372 1519
rect 2366 1514 2372 1515
rect 2374 1519 2380 1520
rect 2374 1515 2375 1519
rect 2379 1518 2380 1519
rect 2622 1519 2628 1520
rect 2379 1516 2465 1518
rect 2379 1515 2380 1516
rect 2374 1514 2380 1515
rect 2622 1515 2623 1519
rect 2627 1515 2628 1519
rect 2622 1514 2628 1515
rect 2750 1519 2756 1520
rect 2750 1515 2751 1519
rect 2755 1515 2756 1519
rect 2750 1514 2756 1515
rect 2870 1519 2876 1520
rect 2870 1515 2871 1519
rect 2875 1515 2876 1519
rect 2870 1514 2876 1515
rect 2998 1519 3004 1520
rect 2998 1515 2999 1519
rect 3003 1515 3004 1519
rect 2998 1514 3004 1515
rect 3018 1519 3024 1520
rect 3018 1515 3019 1519
rect 3023 1518 3024 1519
rect 3023 1516 3097 1518
rect 3023 1515 3024 1516
rect 3018 1514 3024 1515
rect 1403 1512 1489 1514
rect 1403 1511 1404 1512
rect 1398 1510 1404 1511
rect 1806 1511 1812 1512
rect 254 1506 260 1507
rect 1766 1507 1772 1508
rect 110 1502 116 1503
rect 182 1504 188 1505
rect 182 1500 183 1504
rect 187 1500 188 1504
rect 182 1499 188 1500
rect 326 1504 332 1505
rect 326 1500 327 1504
rect 331 1500 332 1504
rect 326 1499 332 1500
rect 470 1504 476 1505
rect 470 1500 471 1504
rect 475 1500 476 1504
rect 470 1499 476 1500
rect 622 1504 628 1505
rect 622 1500 623 1504
rect 627 1500 628 1504
rect 622 1499 628 1500
rect 766 1504 772 1505
rect 766 1500 767 1504
rect 771 1500 772 1504
rect 766 1499 772 1500
rect 910 1504 916 1505
rect 910 1500 911 1504
rect 915 1500 916 1504
rect 910 1499 916 1500
rect 1046 1504 1052 1505
rect 1046 1500 1047 1504
rect 1051 1500 1052 1504
rect 1046 1499 1052 1500
rect 1174 1504 1180 1505
rect 1174 1500 1175 1504
rect 1179 1500 1180 1504
rect 1174 1499 1180 1500
rect 1310 1504 1316 1505
rect 1310 1500 1311 1504
rect 1315 1500 1316 1504
rect 1310 1499 1316 1500
rect 1446 1504 1452 1505
rect 1446 1500 1447 1504
rect 1451 1500 1452 1504
rect 1766 1503 1767 1507
rect 1771 1503 1772 1507
rect 1806 1507 1807 1511
rect 1811 1507 1812 1511
rect 3462 1511 3468 1512
rect 1806 1506 1812 1507
rect 1918 1508 1924 1509
rect 1918 1504 1919 1508
rect 1923 1504 1924 1508
rect 1918 1503 1924 1504
rect 2038 1508 2044 1509
rect 2038 1504 2039 1508
rect 2043 1504 2044 1508
rect 2038 1503 2044 1504
rect 2166 1508 2172 1509
rect 2166 1504 2167 1508
rect 2171 1504 2172 1508
rect 2166 1503 2172 1504
rect 2294 1508 2300 1509
rect 2294 1504 2295 1508
rect 2299 1504 2300 1508
rect 2294 1503 2300 1504
rect 2422 1508 2428 1509
rect 2422 1504 2423 1508
rect 2427 1504 2428 1508
rect 2422 1503 2428 1504
rect 2550 1508 2556 1509
rect 2550 1504 2551 1508
rect 2555 1504 2556 1508
rect 2550 1503 2556 1504
rect 2678 1508 2684 1509
rect 2678 1504 2679 1508
rect 2683 1504 2684 1508
rect 2678 1503 2684 1504
rect 2798 1508 2804 1509
rect 2798 1504 2799 1508
rect 2803 1504 2804 1508
rect 2798 1503 2804 1504
rect 2926 1508 2932 1509
rect 2926 1504 2927 1508
rect 2931 1504 2932 1508
rect 2926 1503 2932 1504
rect 3054 1508 3060 1509
rect 3054 1504 3055 1508
rect 3059 1504 3060 1508
rect 3462 1507 3463 1511
rect 3467 1507 3468 1511
rect 3462 1506 3468 1507
rect 3054 1503 3060 1504
rect 1766 1502 1772 1503
rect 1446 1499 1452 1500
rect 2118 1499 2124 1500
rect 2118 1495 2119 1499
rect 2123 1498 2124 1499
rect 2374 1499 2380 1500
rect 2374 1498 2375 1499
rect 2123 1496 2375 1498
rect 2123 1495 2124 1496
rect 2118 1494 2124 1495
rect 2374 1495 2375 1496
rect 2379 1495 2380 1499
rect 2374 1494 2380 1495
rect 1066 1463 1072 1464
rect 1066 1459 1067 1463
rect 1071 1462 1072 1463
rect 1982 1463 1988 1464
rect 1071 1460 1514 1462
rect 1071 1459 1072 1460
rect 1066 1458 1072 1459
rect 158 1456 164 1457
rect 110 1453 116 1454
rect 110 1449 111 1453
rect 115 1449 116 1453
rect 158 1452 159 1456
rect 163 1452 164 1456
rect 158 1451 164 1452
rect 374 1456 380 1457
rect 374 1452 375 1456
rect 379 1452 380 1456
rect 374 1451 380 1452
rect 582 1456 588 1457
rect 582 1452 583 1456
rect 587 1452 588 1456
rect 582 1451 588 1452
rect 782 1456 788 1457
rect 782 1452 783 1456
rect 787 1452 788 1456
rect 782 1451 788 1452
rect 958 1456 964 1457
rect 958 1452 959 1456
rect 963 1452 964 1456
rect 958 1451 964 1452
rect 1126 1456 1132 1457
rect 1126 1452 1127 1456
rect 1131 1452 1132 1456
rect 1126 1451 1132 1452
rect 1278 1456 1284 1457
rect 1278 1452 1279 1456
rect 1283 1452 1284 1456
rect 1278 1451 1284 1452
rect 1430 1456 1436 1457
rect 1430 1452 1431 1456
rect 1435 1452 1436 1456
rect 1430 1451 1436 1452
rect 110 1448 116 1449
rect 262 1447 268 1448
rect 262 1446 263 1447
rect 233 1444 263 1446
rect 262 1443 263 1444
rect 267 1443 268 1447
rect 262 1442 268 1443
rect 446 1447 452 1448
rect 446 1443 447 1447
rect 451 1443 452 1447
rect 446 1442 452 1443
rect 654 1447 660 1448
rect 654 1443 655 1447
rect 659 1443 660 1447
rect 654 1442 660 1443
rect 846 1447 852 1448
rect 846 1443 847 1447
rect 851 1443 852 1447
rect 1090 1447 1096 1448
rect 1090 1446 1091 1447
rect 1033 1444 1091 1446
rect 846 1442 852 1443
rect 1090 1443 1091 1444
rect 1095 1443 1096 1447
rect 1090 1442 1096 1443
rect 1198 1447 1204 1448
rect 1198 1443 1199 1447
rect 1203 1443 1204 1447
rect 1198 1442 1204 1443
rect 1350 1447 1356 1448
rect 1350 1443 1351 1447
rect 1355 1443 1356 1447
rect 1350 1442 1356 1443
rect 1502 1447 1508 1448
rect 1502 1443 1503 1447
rect 1507 1443 1508 1447
rect 1512 1446 1514 1460
rect 1982 1459 1983 1463
rect 1987 1462 1988 1463
rect 2610 1463 2616 1464
rect 1987 1460 2354 1462
rect 1987 1459 1988 1460
rect 1982 1458 1988 1459
rect 1590 1456 1596 1457
rect 1590 1452 1591 1456
rect 1595 1452 1596 1456
rect 1830 1456 1836 1457
rect 1590 1451 1596 1452
rect 1766 1453 1772 1454
rect 1766 1449 1767 1453
rect 1771 1449 1772 1453
rect 1766 1448 1772 1449
rect 1806 1453 1812 1454
rect 1806 1449 1807 1453
rect 1811 1449 1812 1453
rect 1830 1452 1831 1456
rect 1835 1452 1836 1456
rect 1830 1451 1836 1452
rect 1950 1456 1956 1457
rect 1950 1452 1951 1456
rect 1955 1452 1956 1456
rect 1950 1451 1956 1452
rect 2110 1456 2116 1457
rect 2110 1452 2111 1456
rect 2115 1452 2116 1456
rect 2110 1451 2116 1452
rect 2270 1456 2276 1457
rect 2270 1452 2271 1456
rect 2275 1452 2276 1456
rect 2270 1451 2276 1452
rect 1806 1448 1812 1449
rect 2022 1447 2028 1448
rect 1512 1444 1633 1446
rect 1502 1442 1508 1443
rect 2022 1443 2023 1447
rect 2027 1443 2028 1447
rect 2022 1442 2028 1443
rect 2182 1447 2188 1448
rect 2182 1443 2183 1447
rect 2187 1443 2188 1447
rect 2182 1442 2188 1443
rect 2342 1447 2348 1448
rect 2342 1443 2343 1447
rect 2347 1443 2348 1447
rect 2352 1446 2354 1460
rect 2610 1459 2611 1463
rect 2615 1462 2616 1463
rect 2615 1460 3090 1462
rect 2615 1459 2616 1460
rect 2610 1458 2616 1459
rect 2430 1456 2436 1457
rect 2430 1452 2431 1456
rect 2435 1452 2436 1456
rect 2430 1451 2436 1452
rect 2590 1456 2596 1457
rect 2590 1452 2591 1456
rect 2595 1452 2596 1456
rect 2590 1451 2596 1452
rect 2734 1456 2740 1457
rect 2734 1452 2735 1456
rect 2739 1452 2740 1456
rect 2734 1451 2740 1452
rect 2870 1456 2876 1457
rect 2870 1452 2871 1456
rect 2875 1452 2876 1456
rect 2870 1451 2876 1452
rect 3006 1456 3012 1457
rect 3006 1452 3007 1456
rect 3011 1452 3012 1456
rect 3006 1451 3012 1452
rect 2806 1447 2812 1448
rect 2352 1444 2473 1446
rect 2342 1442 2348 1443
rect 2806 1443 2807 1447
rect 2811 1443 2812 1447
rect 2806 1442 2812 1443
rect 2942 1447 2948 1448
rect 2942 1443 2943 1447
rect 2947 1443 2948 1447
rect 2942 1442 2948 1443
rect 3078 1447 3084 1448
rect 3078 1443 3079 1447
rect 3083 1443 3084 1447
rect 3088 1446 3090 1460
rect 3134 1456 3140 1457
rect 3134 1452 3135 1456
rect 3139 1452 3140 1456
rect 3134 1451 3140 1452
rect 3262 1456 3268 1457
rect 3262 1452 3263 1456
rect 3267 1452 3268 1456
rect 3262 1451 3268 1452
rect 3366 1456 3372 1457
rect 3366 1452 3367 1456
rect 3371 1452 3372 1456
rect 3366 1451 3372 1452
rect 3462 1453 3468 1454
rect 3462 1449 3463 1453
rect 3467 1449 3468 1453
rect 3462 1448 3468 1449
rect 3334 1447 3340 1448
rect 3088 1444 3177 1446
rect 3078 1442 3084 1443
rect 3334 1443 3335 1447
rect 3339 1443 3340 1447
rect 3334 1442 3340 1443
rect 3430 1447 3436 1448
rect 3430 1443 3431 1447
rect 3435 1443 3436 1447
rect 3430 1442 3436 1443
rect 1903 1439 1909 1440
rect 158 1437 164 1438
rect 110 1436 116 1437
rect 110 1432 111 1436
rect 115 1432 116 1436
rect 158 1433 159 1437
rect 163 1433 164 1437
rect 158 1432 164 1433
rect 374 1437 380 1438
rect 374 1433 375 1437
rect 379 1433 380 1437
rect 374 1432 380 1433
rect 582 1437 588 1438
rect 582 1433 583 1437
rect 587 1433 588 1437
rect 582 1432 588 1433
rect 782 1437 788 1438
rect 782 1433 783 1437
rect 787 1433 788 1437
rect 782 1432 788 1433
rect 958 1437 964 1438
rect 958 1433 959 1437
rect 963 1433 964 1437
rect 958 1432 964 1433
rect 1126 1437 1132 1438
rect 1126 1433 1127 1437
rect 1131 1433 1132 1437
rect 1126 1432 1132 1433
rect 1278 1437 1284 1438
rect 1278 1433 1279 1437
rect 1283 1433 1284 1437
rect 1278 1432 1284 1433
rect 1430 1437 1436 1438
rect 1430 1433 1431 1437
rect 1435 1433 1436 1437
rect 1430 1432 1436 1433
rect 1590 1437 1596 1438
rect 1830 1437 1836 1438
rect 1590 1433 1591 1437
rect 1595 1433 1596 1437
rect 1590 1432 1596 1433
rect 1766 1436 1772 1437
rect 1766 1432 1767 1436
rect 1771 1432 1772 1436
rect 110 1431 116 1432
rect 1766 1431 1772 1432
rect 1806 1436 1812 1437
rect 1806 1432 1807 1436
rect 1811 1432 1812 1436
rect 1830 1433 1831 1437
rect 1835 1433 1836 1437
rect 1903 1435 1904 1439
rect 1908 1438 1909 1439
rect 2663 1439 2669 1440
rect 1908 1436 1938 1438
rect 1908 1435 1909 1436
rect 1903 1434 1909 1435
rect 1830 1432 1836 1433
rect 1806 1431 1812 1432
rect 1936 1422 1938 1436
rect 1950 1437 1956 1438
rect 1950 1433 1951 1437
rect 1955 1433 1956 1437
rect 1950 1432 1956 1433
rect 2110 1437 2116 1438
rect 2110 1433 2111 1437
rect 2115 1433 2116 1437
rect 2110 1432 2116 1433
rect 2270 1437 2276 1438
rect 2270 1433 2271 1437
rect 2275 1433 2276 1437
rect 2270 1432 2276 1433
rect 2430 1437 2436 1438
rect 2430 1433 2431 1437
rect 2435 1433 2436 1437
rect 2430 1432 2436 1433
rect 2590 1437 2596 1438
rect 2590 1433 2591 1437
rect 2595 1433 2596 1437
rect 2663 1435 2664 1439
rect 2668 1438 2669 1439
rect 2668 1436 2710 1438
rect 2668 1435 2669 1436
rect 2663 1434 2669 1435
rect 2590 1432 2596 1433
rect 2708 1430 2710 1436
rect 2734 1437 2740 1438
rect 2734 1433 2735 1437
rect 2739 1433 2740 1437
rect 2734 1432 2740 1433
rect 2870 1437 2876 1438
rect 2870 1433 2871 1437
rect 2875 1433 2876 1437
rect 2870 1432 2876 1433
rect 3006 1437 3012 1438
rect 3006 1433 3007 1437
rect 3011 1433 3012 1437
rect 3006 1432 3012 1433
rect 3134 1437 3140 1438
rect 3134 1433 3135 1437
rect 3139 1433 3140 1437
rect 3134 1432 3140 1433
rect 3262 1437 3268 1438
rect 3262 1433 3263 1437
rect 3267 1433 3268 1437
rect 3262 1432 3268 1433
rect 3366 1437 3372 1438
rect 3366 1433 3367 1437
rect 3371 1433 3372 1437
rect 3366 1432 3372 1433
rect 3462 1436 3468 1437
rect 3462 1432 3463 1436
rect 3467 1432 3468 1436
rect 3462 1431 3468 1432
rect 2708 1428 2746 1430
rect 1936 1420 2001 1422
rect 207 1419 213 1420
rect 207 1415 208 1419
rect 212 1418 213 1419
rect 254 1419 260 1420
rect 254 1418 255 1419
rect 212 1416 255 1418
rect 212 1415 213 1416
rect 207 1414 213 1415
rect 254 1415 255 1416
rect 259 1415 260 1419
rect 254 1414 260 1415
rect 262 1419 268 1420
rect 262 1415 263 1419
rect 267 1418 268 1419
rect 423 1419 429 1420
rect 423 1418 424 1419
rect 267 1416 424 1418
rect 267 1415 268 1416
rect 262 1414 268 1415
rect 423 1415 424 1416
rect 428 1415 429 1419
rect 423 1414 429 1415
rect 631 1419 640 1420
rect 631 1415 632 1419
rect 639 1415 640 1419
rect 631 1414 640 1415
rect 654 1419 660 1420
rect 654 1415 655 1419
rect 659 1418 660 1419
rect 831 1419 837 1420
rect 831 1418 832 1419
rect 659 1416 832 1418
rect 659 1415 660 1416
rect 654 1414 660 1415
rect 831 1415 832 1416
rect 836 1415 837 1419
rect 831 1414 837 1415
rect 1007 1419 1013 1420
rect 1007 1415 1008 1419
rect 1012 1418 1013 1419
rect 1090 1419 1096 1420
rect 1012 1416 1086 1418
rect 1012 1415 1013 1416
rect 1007 1414 1013 1415
rect 1084 1410 1086 1416
rect 1090 1415 1091 1419
rect 1095 1418 1096 1419
rect 1175 1419 1181 1420
rect 1175 1418 1176 1419
rect 1095 1416 1176 1418
rect 1095 1415 1096 1416
rect 1090 1414 1096 1415
rect 1175 1415 1176 1416
rect 1180 1415 1181 1419
rect 1175 1414 1181 1415
rect 1198 1419 1204 1420
rect 1198 1415 1199 1419
rect 1203 1418 1204 1419
rect 1327 1419 1333 1420
rect 1327 1418 1328 1419
rect 1203 1416 1328 1418
rect 1203 1415 1204 1416
rect 1198 1414 1204 1415
rect 1327 1415 1328 1416
rect 1332 1415 1333 1419
rect 1327 1414 1333 1415
rect 1350 1419 1356 1420
rect 1350 1415 1351 1419
rect 1355 1418 1356 1419
rect 1479 1419 1485 1420
rect 1479 1418 1480 1419
rect 1355 1416 1480 1418
rect 1355 1415 1356 1416
rect 1350 1414 1356 1415
rect 1479 1415 1480 1416
rect 1484 1415 1485 1419
rect 1479 1414 1485 1415
rect 1502 1419 1508 1420
rect 1502 1415 1503 1419
rect 1507 1418 1508 1419
rect 1639 1419 1645 1420
rect 1639 1418 1640 1419
rect 1507 1416 1640 1418
rect 1507 1415 1508 1416
rect 1502 1414 1508 1415
rect 1639 1415 1640 1416
rect 1644 1415 1645 1419
rect 1639 1414 1645 1415
rect 1879 1419 1885 1420
rect 1879 1415 1880 1419
rect 1884 1418 1885 1419
rect 1999 1419 2005 1420
rect 1884 1416 1942 1418
rect 1884 1415 1885 1416
rect 1879 1414 1885 1415
rect 1398 1411 1404 1412
rect 1398 1410 1399 1411
rect 1084 1408 1399 1410
rect 1398 1407 1399 1408
rect 1403 1407 1404 1411
rect 1398 1406 1404 1407
rect 1742 1411 1748 1412
rect 1742 1407 1743 1411
rect 1747 1410 1748 1411
rect 1940 1410 1942 1416
rect 1999 1415 2000 1419
rect 2004 1415 2005 1419
rect 1999 1414 2005 1415
rect 2022 1419 2028 1420
rect 2022 1415 2023 1419
rect 2027 1418 2028 1419
rect 2159 1419 2165 1420
rect 2159 1418 2160 1419
rect 2027 1416 2160 1418
rect 2027 1415 2028 1416
rect 2022 1414 2028 1415
rect 2159 1415 2160 1416
rect 2164 1415 2165 1419
rect 2159 1414 2165 1415
rect 2182 1419 2188 1420
rect 2182 1415 2183 1419
rect 2187 1418 2188 1419
rect 2319 1419 2325 1420
rect 2319 1418 2320 1419
rect 2187 1416 2320 1418
rect 2187 1415 2188 1416
rect 2182 1414 2188 1415
rect 2319 1415 2320 1416
rect 2324 1415 2325 1419
rect 2319 1414 2325 1415
rect 2342 1419 2348 1420
rect 2342 1415 2343 1419
rect 2347 1418 2348 1419
rect 2479 1419 2485 1420
rect 2479 1418 2480 1419
rect 2347 1416 2480 1418
rect 2347 1415 2348 1416
rect 2342 1414 2348 1415
rect 2479 1415 2480 1416
rect 2484 1415 2485 1419
rect 2479 1414 2485 1415
rect 2639 1419 2645 1420
rect 2639 1415 2640 1419
rect 2644 1418 2645 1419
rect 2744 1418 2746 1428
rect 2783 1419 2789 1420
rect 2783 1418 2784 1419
rect 2644 1416 2742 1418
rect 2744 1416 2784 1418
rect 2644 1415 2645 1416
rect 2639 1414 2645 1415
rect 2342 1411 2348 1412
rect 2342 1410 2343 1411
rect 1747 1408 1906 1410
rect 1940 1408 2343 1410
rect 1747 1407 1748 1408
rect 1742 1406 1748 1407
rect 183 1403 189 1404
rect 183 1399 184 1403
rect 188 1402 189 1403
rect 282 1403 288 1404
rect 282 1402 283 1403
rect 188 1400 283 1402
rect 188 1399 189 1400
rect 183 1398 189 1399
rect 282 1399 283 1400
rect 287 1399 288 1403
rect 282 1398 288 1399
rect 351 1403 357 1404
rect 351 1399 352 1403
rect 356 1402 357 1403
rect 391 1403 397 1404
rect 391 1402 392 1403
rect 356 1400 392 1402
rect 356 1399 357 1400
rect 351 1398 357 1399
rect 391 1399 392 1400
rect 396 1399 397 1403
rect 391 1398 397 1399
rect 446 1403 452 1404
rect 446 1399 447 1403
rect 451 1402 452 1403
rect 543 1403 549 1404
rect 543 1402 544 1403
rect 451 1400 544 1402
rect 451 1399 452 1400
rect 446 1398 452 1399
rect 543 1399 544 1400
rect 548 1399 549 1403
rect 543 1398 549 1399
rect 727 1403 733 1404
rect 727 1399 728 1403
rect 732 1402 733 1403
rect 758 1403 764 1404
rect 758 1402 759 1403
rect 732 1400 759 1402
rect 732 1399 733 1400
rect 727 1398 733 1399
rect 758 1399 759 1400
rect 763 1399 764 1403
rect 758 1398 764 1399
rect 903 1403 909 1404
rect 903 1399 904 1403
rect 908 1402 909 1403
rect 974 1403 980 1404
rect 974 1402 975 1403
rect 908 1400 975 1402
rect 908 1399 909 1400
rect 903 1398 909 1399
rect 974 1399 975 1400
rect 979 1399 980 1403
rect 974 1398 980 1399
rect 1063 1403 1072 1404
rect 1063 1399 1064 1403
rect 1071 1399 1072 1403
rect 1063 1398 1072 1399
rect 1086 1403 1092 1404
rect 1086 1399 1087 1403
rect 1091 1402 1092 1403
rect 1215 1403 1221 1404
rect 1215 1402 1216 1403
rect 1091 1400 1216 1402
rect 1091 1399 1092 1400
rect 1086 1398 1092 1399
rect 1215 1399 1216 1400
rect 1220 1399 1221 1403
rect 1215 1398 1221 1399
rect 1238 1403 1244 1404
rect 1238 1399 1239 1403
rect 1243 1402 1244 1403
rect 1351 1403 1357 1404
rect 1351 1402 1352 1403
rect 1243 1400 1352 1402
rect 1243 1399 1244 1400
rect 1238 1398 1244 1399
rect 1351 1399 1352 1400
rect 1356 1399 1357 1403
rect 1351 1398 1357 1399
rect 1374 1403 1380 1404
rect 1374 1399 1375 1403
rect 1379 1402 1380 1403
rect 1479 1403 1485 1404
rect 1479 1402 1480 1403
rect 1379 1400 1480 1402
rect 1379 1399 1380 1400
rect 1374 1398 1380 1399
rect 1479 1399 1480 1400
rect 1484 1399 1485 1403
rect 1479 1398 1485 1399
rect 1502 1403 1508 1404
rect 1502 1399 1503 1403
rect 1507 1402 1508 1403
rect 1607 1403 1613 1404
rect 1607 1402 1608 1403
rect 1507 1400 1608 1402
rect 1507 1399 1508 1400
rect 1502 1398 1508 1399
rect 1607 1399 1608 1400
rect 1612 1399 1613 1403
rect 1607 1398 1613 1399
rect 1719 1403 1725 1404
rect 1719 1399 1720 1403
rect 1724 1402 1725 1403
rect 1750 1403 1756 1404
rect 1750 1402 1751 1403
rect 1724 1400 1751 1402
rect 1724 1399 1725 1400
rect 1719 1398 1725 1399
rect 1750 1399 1751 1400
rect 1755 1399 1756 1403
rect 1750 1398 1756 1399
rect 1879 1403 1885 1404
rect 1879 1399 1880 1403
rect 1884 1402 1885 1403
rect 1894 1403 1900 1404
rect 1894 1402 1895 1403
rect 1884 1400 1895 1402
rect 1884 1399 1885 1400
rect 1879 1398 1885 1399
rect 1894 1399 1895 1400
rect 1899 1399 1900 1403
rect 1904 1402 1906 1408
rect 2342 1407 2343 1408
rect 2347 1407 2348 1411
rect 2740 1410 2742 1416
rect 2783 1415 2784 1416
rect 2788 1415 2789 1419
rect 2783 1414 2789 1415
rect 2806 1419 2812 1420
rect 2806 1415 2807 1419
rect 2811 1418 2812 1419
rect 2919 1419 2925 1420
rect 2919 1418 2920 1419
rect 2811 1416 2920 1418
rect 2811 1415 2812 1416
rect 2806 1414 2812 1415
rect 2919 1415 2920 1416
rect 2924 1415 2925 1419
rect 2919 1414 2925 1415
rect 2942 1419 2948 1420
rect 2942 1415 2943 1419
rect 2947 1418 2948 1419
rect 3055 1419 3061 1420
rect 3055 1418 3056 1419
rect 2947 1416 3056 1418
rect 2947 1415 2948 1416
rect 2942 1414 2948 1415
rect 3055 1415 3056 1416
rect 3060 1415 3061 1419
rect 3055 1414 3061 1415
rect 3078 1419 3084 1420
rect 3078 1415 3079 1419
rect 3083 1418 3084 1419
rect 3183 1419 3189 1420
rect 3183 1418 3184 1419
rect 3083 1416 3184 1418
rect 3083 1415 3084 1416
rect 3078 1414 3084 1415
rect 3183 1415 3184 1416
rect 3188 1415 3189 1419
rect 3183 1414 3189 1415
rect 3311 1419 3317 1420
rect 3311 1415 3312 1419
rect 3316 1418 3317 1419
rect 3326 1419 3332 1420
rect 3326 1418 3327 1419
rect 3316 1416 3327 1418
rect 3316 1415 3317 1416
rect 3311 1414 3317 1415
rect 3326 1415 3327 1416
rect 3331 1415 3332 1419
rect 3326 1414 3332 1415
rect 3334 1419 3340 1420
rect 3334 1415 3335 1419
rect 3339 1418 3340 1419
rect 3415 1419 3421 1420
rect 3415 1418 3416 1419
rect 3339 1416 3416 1418
rect 3339 1415 3340 1416
rect 3334 1414 3340 1415
rect 3415 1415 3416 1416
rect 3420 1415 3421 1419
rect 3415 1414 3421 1415
rect 3018 1411 3024 1412
rect 3018 1410 3019 1411
rect 2740 1408 3019 1410
rect 2342 1406 2348 1407
rect 3018 1407 3019 1408
rect 3023 1407 3024 1411
rect 3018 1406 3024 1407
rect 2055 1403 2061 1404
rect 2055 1402 2056 1403
rect 1904 1400 2056 1402
rect 1894 1398 1900 1399
rect 2055 1399 2056 1400
rect 2060 1399 2061 1403
rect 2055 1398 2061 1399
rect 2078 1403 2084 1404
rect 2078 1399 2079 1403
rect 2083 1402 2084 1403
rect 2247 1403 2253 1404
rect 2247 1402 2248 1403
rect 2083 1400 2248 1402
rect 2083 1399 2084 1400
rect 2078 1398 2084 1399
rect 2247 1399 2248 1400
rect 2252 1399 2253 1403
rect 2247 1398 2253 1399
rect 2334 1403 2340 1404
rect 2334 1399 2335 1403
rect 2339 1402 2340 1403
rect 2431 1403 2437 1404
rect 2431 1402 2432 1403
rect 2339 1400 2432 1402
rect 2339 1399 2340 1400
rect 2334 1398 2340 1399
rect 2431 1399 2432 1400
rect 2436 1399 2437 1403
rect 2431 1398 2437 1399
rect 2607 1403 2616 1404
rect 2607 1399 2608 1403
rect 2615 1399 2616 1403
rect 2607 1398 2616 1399
rect 2630 1403 2636 1404
rect 2630 1399 2631 1403
rect 2635 1402 2636 1403
rect 2767 1403 2773 1404
rect 2767 1402 2768 1403
rect 2635 1400 2768 1402
rect 2635 1399 2636 1400
rect 2630 1398 2636 1399
rect 2767 1399 2768 1400
rect 2772 1399 2773 1403
rect 2767 1398 2773 1399
rect 2790 1403 2796 1404
rect 2790 1399 2791 1403
rect 2795 1402 2796 1403
rect 2911 1403 2917 1404
rect 2911 1402 2912 1403
rect 2795 1400 2912 1402
rect 2795 1399 2796 1400
rect 2790 1398 2796 1399
rect 2911 1399 2912 1400
rect 2916 1399 2917 1403
rect 2911 1398 2917 1399
rect 2934 1403 2940 1404
rect 2934 1399 2935 1403
rect 2939 1402 2940 1403
rect 3047 1403 3053 1404
rect 3047 1402 3048 1403
rect 2939 1400 3048 1402
rect 2939 1399 2940 1400
rect 2934 1398 2940 1399
rect 3047 1399 3048 1400
rect 3052 1399 3053 1403
rect 3047 1398 3053 1399
rect 3070 1403 3076 1404
rect 3070 1399 3071 1403
rect 3075 1402 3076 1403
rect 3175 1403 3181 1404
rect 3175 1402 3176 1403
rect 3075 1400 3176 1402
rect 3075 1399 3076 1400
rect 3070 1398 3076 1399
rect 3175 1399 3176 1400
rect 3180 1399 3181 1403
rect 3175 1398 3181 1399
rect 3198 1403 3204 1404
rect 3198 1399 3199 1403
rect 3203 1402 3204 1403
rect 3303 1403 3309 1404
rect 3303 1402 3304 1403
rect 3203 1400 3304 1402
rect 3203 1399 3204 1400
rect 3198 1398 3204 1399
rect 3303 1399 3304 1400
rect 3308 1399 3309 1403
rect 3303 1398 3309 1399
rect 3415 1403 3421 1404
rect 3415 1399 3416 1403
rect 3420 1402 3421 1403
rect 3430 1403 3436 1404
rect 3430 1402 3431 1403
rect 3420 1400 3431 1402
rect 3420 1399 3421 1400
rect 3415 1398 3421 1399
rect 3430 1399 3431 1400
rect 3435 1399 3436 1403
rect 3430 1398 3436 1399
rect 110 1388 116 1389
rect 1766 1388 1772 1389
rect 110 1384 111 1388
rect 115 1384 116 1388
rect 110 1383 116 1384
rect 134 1387 140 1388
rect 134 1383 135 1387
rect 139 1383 140 1387
rect 134 1382 140 1383
rect 302 1387 308 1388
rect 302 1383 303 1387
rect 307 1383 308 1387
rect 302 1382 308 1383
rect 494 1387 500 1388
rect 494 1383 495 1387
rect 499 1383 500 1387
rect 494 1382 500 1383
rect 678 1387 684 1388
rect 678 1383 679 1387
rect 683 1383 684 1387
rect 678 1382 684 1383
rect 854 1387 860 1388
rect 854 1383 855 1387
rect 859 1383 860 1387
rect 854 1382 860 1383
rect 1014 1387 1020 1388
rect 1014 1383 1015 1387
rect 1019 1383 1020 1387
rect 1014 1382 1020 1383
rect 1166 1387 1172 1388
rect 1166 1383 1167 1387
rect 1171 1383 1172 1387
rect 1166 1382 1172 1383
rect 1302 1387 1308 1388
rect 1302 1383 1303 1387
rect 1307 1383 1308 1387
rect 1302 1382 1308 1383
rect 1430 1387 1436 1388
rect 1430 1383 1431 1387
rect 1435 1383 1436 1387
rect 1430 1382 1436 1383
rect 1558 1387 1564 1388
rect 1558 1383 1559 1387
rect 1563 1383 1564 1387
rect 1558 1382 1564 1383
rect 1670 1387 1676 1388
rect 1670 1383 1671 1387
rect 1675 1383 1676 1387
rect 1766 1384 1767 1388
rect 1771 1384 1772 1388
rect 1766 1383 1772 1384
rect 1806 1388 1812 1389
rect 3462 1388 3468 1389
rect 1806 1384 1807 1388
rect 1811 1384 1812 1388
rect 1806 1383 1812 1384
rect 1830 1387 1836 1388
rect 1830 1383 1831 1387
rect 1835 1383 1836 1387
rect 1670 1382 1676 1383
rect 1830 1382 1836 1383
rect 2006 1387 2012 1388
rect 2006 1383 2007 1387
rect 2011 1383 2012 1387
rect 2006 1382 2012 1383
rect 2198 1387 2204 1388
rect 2198 1383 2199 1387
rect 2203 1383 2204 1387
rect 2198 1382 2204 1383
rect 2382 1387 2388 1388
rect 2382 1383 2383 1387
rect 2387 1383 2388 1387
rect 2382 1382 2388 1383
rect 2558 1387 2564 1388
rect 2558 1383 2559 1387
rect 2563 1383 2564 1387
rect 2558 1382 2564 1383
rect 2718 1387 2724 1388
rect 2718 1383 2719 1387
rect 2723 1383 2724 1387
rect 2718 1382 2724 1383
rect 2862 1387 2868 1388
rect 2862 1383 2863 1387
rect 2867 1383 2868 1387
rect 2862 1382 2868 1383
rect 2998 1387 3004 1388
rect 2998 1383 2999 1387
rect 3003 1383 3004 1387
rect 2998 1382 3004 1383
rect 3126 1387 3132 1388
rect 3126 1383 3127 1387
rect 3131 1383 3132 1387
rect 3126 1382 3132 1383
rect 3254 1387 3260 1388
rect 3254 1383 3255 1387
rect 3259 1383 3260 1387
rect 3254 1382 3260 1383
rect 3366 1387 3372 1388
rect 3366 1383 3367 1387
rect 3371 1383 3372 1387
rect 3462 1384 3463 1388
rect 3467 1384 3468 1388
rect 3462 1383 3468 1384
rect 3366 1382 3372 1383
rect 282 1379 288 1380
rect 282 1375 283 1379
rect 287 1378 288 1379
rect 391 1379 397 1380
rect 287 1376 345 1378
rect 287 1375 288 1376
rect 282 1374 288 1375
rect 391 1375 392 1379
rect 396 1378 397 1379
rect 634 1379 640 1380
rect 396 1376 537 1378
rect 396 1375 397 1376
rect 391 1374 397 1375
rect 634 1375 635 1379
rect 639 1378 640 1379
rect 758 1379 764 1380
rect 639 1376 721 1378
rect 639 1375 640 1376
rect 634 1374 640 1375
rect 758 1375 759 1379
rect 763 1378 764 1379
rect 1086 1379 1092 1380
rect 763 1376 897 1378
rect 763 1375 764 1376
rect 758 1374 764 1375
rect 1086 1375 1087 1379
rect 1091 1375 1092 1379
rect 1086 1374 1092 1375
rect 1238 1379 1244 1380
rect 1238 1375 1239 1379
rect 1243 1375 1244 1379
rect 1238 1374 1244 1375
rect 1374 1379 1380 1380
rect 1374 1375 1375 1379
rect 1379 1375 1380 1379
rect 1374 1374 1380 1375
rect 1502 1379 1508 1380
rect 1502 1375 1503 1379
rect 1507 1375 1508 1379
rect 1502 1374 1508 1375
rect 1510 1379 1516 1380
rect 1510 1375 1511 1379
rect 1515 1378 1516 1379
rect 1742 1379 1748 1380
rect 1515 1376 1601 1378
rect 1515 1375 1516 1376
rect 1510 1374 1516 1375
rect 1742 1375 1743 1379
rect 1747 1375 1748 1379
rect 1742 1374 1748 1375
rect 1750 1379 1756 1380
rect 1750 1375 1751 1379
rect 1755 1378 1756 1379
rect 2078 1379 2084 1380
rect 1755 1376 1873 1378
rect 1755 1375 1756 1376
rect 1750 1374 1756 1375
rect 2078 1375 2079 1379
rect 2083 1375 2084 1379
rect 2334 1379 2340 1380
rect 2334 1378 2335 1379
rect 2273 1376 2335 1378
rect 2078 1374 2084 1375
rect 2334 1375 2335 1376
rect 2339 1375 2340 1379
rect 2334 1374 2340 1375
rect 2342 1379 2348 1380
rect 2342 1375 2343 1379
rect 2347 1378 2348 1379
rect 2630 1379 2636 1380
rect 2347 1376 2425 1378
rect 2347 1375 2348 1376
rect 2342 1374 2348 1375
rect 2630 1375 2631 1379
rect 2635 1375 2636 1379
rect 2630 1374 2636 1375
rect 2790 1379 2796 1380
rect 2790 1375 2791 1379
rect 2795 1375 2796 1379
rect 2790 1374 2796 1375
rect 2934 1379 2940 1380
rect 2934 1375 2935 1379
rect 2939 1375 2940 1379
rect 2934 1374 2940 1375
rect 3070 1379 3076 1380
rect 3070 1375 3071 1379
rect 3075 1375 3076 1379
rect 3070 1374 3076 1375
rect 3198 1379 3204 1380
rect 3198 1375 3199 1379
rect 3203 1375 3204 1379
rect 3198 1374 3204 1375
rect 3326 1379 3332 1380
rect 3326 1375 3327 1379
rect 3331 1375 3332 1379
rect 3326 1374 3332 1375
rect 3438 1375 3444 1376
rect 110 1371 116 1372
rect 110 1367 111 1371
rect 115 1367 116 1371
rect 198 1371 204 1372
rect 110 1366 116 1367
rect 134 1368 140 1369
rect 134 1364 135 1368
rect 139 1364 140 1368
rect 198 1367 199 1371
rect 203 1370 204 1371
rect 208 1370 210 1373
rect 203 1368 210 1370
rect 1766 1371 1772 1372
rect 302 1368 308 1369
rect 203 1367 204 1368
rect 198 1366 204 1367
rect 134 1363 140 1364
rect 302 1364 303 1368
rect 307 1364 308 1368
rect 302 1363 308 1364
rect 494 1368 500 1369
rect 494 1364 495 1368
rect 499 1364 500 1368
rect 494 1363 500 1364
rect 678 1368 684 1369
rect 678 1364 679 1368
rect 683 1364 684 1368
rect 678 1363 684 1364
rect 854 1368 860 1369
rect 854 1364 855 1368
rect 859 1364 860 1368
rect 854 1363 860 1364
rect 1014 1368 1020 1369
rect 1014 1364 1015 1368
rect 1019 1364 1020 1368
rect 1014 1363 1020 1364
rect 1166 1368 1172 1369
rect 1166 1364 1167 1368
rect 1171 1364 1172 1368
rect 1166 1363 1172 1364
rect 1302 1368 1308 1369
rect 1302 1364 1303 1368
rect 1307 1364 1308 1368
rect 1302 1363 1308 1364
rect 1430 1368 1436 1369
rect 1430 1364 1431 1368
rect 1435 1364 1436 1368
rect 1430 1363 1436 1364
rect 1558 1368 1564 1369
rect 1558 1364 1559 1368
rect 1563 1364 1564 1368
rect 1558 1363 1564 1364
rect 1670 1368 1676 1369
rect 1670 1364 1671 1368
rect 1675 1364 1676 1368
rect 1766 1367 1767 1371
rect 1771 1367 1772 1371
rect 1766 1366 1772 1367
rect 1806 1371 1812 1372
rect 1806 1367 1807 1371
rect 1811 1367 1812 1371
rect 3438 1371 3439 1375
rect 3443 1371 3444 1375
rect 3438 1370 3444 1371
rect 3462 1371 3468 1372
rect 1806 1366 1812 1367
rect 1830 1368 1836 1369
rect 1670 1363 1676 1364
rect 1830 1364 1831 1368
rect 1835 1364 1836 1368
rect 1830 1363 1836 1364
rect 2006 1368 2012 1369
rect 2006 1364 2007 1368
rect 2011 1364 2012 1368
rect 2006 1363 2012 1364
rect 2198 1368 2204 1369
rect 2198 1364 2199 1368
rect 2203 1364 2204 1368
rect 2198 1363 2204 1364
rect 2382 1368 2388 1369
rect 2382 1364 2383 1368
rect 2387 1364 2388 1368
rect 2382 1363 2388 1364
rect 2558 1368 2564 1369
rect 2558 1364 2559 1368
rect 2563 1364 2564 1368
rect 2558 1363 2564 1364
rect 2718 1368 2724 1369
rect 2718 1364 2719 1368
rect 2723 1364 2724 1368
rect 2718 1363 2724 1364
rect 2862 1368 2868 1369
rect 2862 1364 2863 1368
rect 2867 1364 2868 1368
rect 2862 1363 2868 1364
rect 2998 1368 3004 1369
rect 2998 1364 2999 1368
rect 3003 1364 3004 1368
rect 2998 1363 3004 1364
rect 3126 1368 3132 1369
rect 3126 1364 3127 1368
rect 3131 1364 3132 1368
rect 3126 1363 3132 1364
rect 3254 1368 3260 1369
rect 3254 1364 3255 1368
rect 3259 1364 3260 1368
rect 3254 1363 3260 1364
rect 3366 1368 3372 1369
rect 3366 1364 3367 1368
rect 3371 1364 3372 1368
rect 3462 1367 3463 1371
rect 3467 1367 3468 1371
rect 3462 1366 3468 1367
rect 3366 1363 3372 1364
rect 2018 1323 2024 1324
rect 134 1320 140 1321
rect 110 1317 116 1318
rect 110 1313 111 1317
rect 115 1313 116 1317
rect 134 1316 135 1320
rect 139 1316 140 1320
rect 134 1315 140 1316
rect 246 1320 252 1321
rect 246 1316 247 1320
rect 251 1316 252 1320
rect 246 1315 252 1316
rect 398 1320 404 1321
rect 398 1316 399 1320
rect 403 1316 404 1320
rect 398 1315 404 1316
rect 558 1320 564 1321
rect 558 1316 559 1320
rect 563 1316 564 1320
rect 558 1315 564 1316
rect 726 1320 732 1321
rect 726 1316 727 1320
rect 731 1316 732 1320
rect 726 1315 732 1316
rect 894 1320 900 1321
rect 894 1316 895 1320
rect 899 1316 900 1320
rect 894 1315 900 1316
rect 1062 1320 1068 1321
rect 1062 1316 1063 1320
rect 1067 1316 1068 1320
rect 1062 1315 1068 1316
rect 1222 1320 1228 1321
rect 1222 1316 1223 1320
rect 1227 1316 1228 1320
rect 1222 1315 1228 1316
rect 1374 1320 1380 1321
rect 1374 1316 1375 1320
rect 1379 1316 1380 1320
rect 1374 1315 1380 1316
rect 1534 1320 1540 1321
rect 1534 1316 1535 1320
rect 1539 1316 1540 1320
rect 1534 1315 1540 1316
rect 1670 1320 1676 1321
rect 1670 1316 1671 1320
rect 1675 1316 1676 1320
rect 2018 1319 2019 1323
rect 2023 1322 2024 1323
rect 2023 1320 2410 1322
rect 2023 1319 2024 1320
rect 2018 1318 2024 1319
rect 1670 1315 1676 1316
rect 1766 1317 1772 1318
rect 110 1312 116 1313
rect 1766 1313 1767 1317
rect 1771 1313 1772 1317
rect 1830 1316 1836 1317
rect 1766 1312 1772 1313
rect 1806 1313 1812 1314
rect 206 1311 212 1312
rect 206 1307 207 1311
rect 211 1307 212 1311
rect 206 1306 212 1307
rect 318 1311 324 1312
rect 318 1307 319 1311
rect 323 1307 324 1311
rect 318 1306 324 1307
rect 470 1311 476 1312
rect 470 1307 471 1311
rect 475 1307 476 1311
rect 470 1306 476 1307
rect 498 1311 504 1312
rect 498 1307 499 1311
rect 503 1310 504 1311
rect 798 1311 804 1312
rect 503 1308 601 1310
rect 503 1307 504 1308
rect 498 1306 504 1307
rect 798 1307 799 1311
rect 803 1307 804 1311
rect 798 1306 804 1307
rect 966 1311 972 1312
rect 966 1307 967 1311
rect 971 1307 972 1311
rect 966 1306 972 1307
rect 974 1311 980 1312
rect 974 1307 975 1311
rect 979 1310 980 1311
rect 1294 1311 1300 1312
rect 979 1308 1105 1310
rect 979 1307 980 1308
rect 974 1306 980 1307
rect 1294 1307 1295 1311
rect 1299 1307 1300 1311
rect 1294 1306 1300 1307
rect 1446 1311 1452 1312
rect 1446 1307 1447 1311
rect 1451 1307 1452 1311
rect 1446 1306 1452 1307
rect 1606 1311 1612 1312
rect 1606 1307 1607 1311
rect 1611 1307 1612 1311
rect 1606 1306 1612 1307
rect 1622 1311 1628 1312
rect 1622 1307 1623 1311
rect 1627 1310 1628 1311
rect 1627 1308 1713 1310
rect 1806 1309 1807 1313
rect 1811 1309 1812 1313
rect 1830 1312 1831 1316
rect 1835 1312 1836 1316
rect 1830 1311 1836 1312
rect 1966 1316 1972 1317
rect 1966 1312 1967 1316
rect 1971 1312 1972 1316
rect 1966 1311 1972 1312
rect 2142 1316 2148 1317
rect 2142 1312 2143 1316
rect 2147 1312 2148 1316
rect 2142 1311 2148 1312
rect 2326 1316 2332 1317
rect 2326 1312 2327 1316
rect 2331 1312 2332 1316
rect 2326 1311 2332 1312
rect 1806 1308 1812 1309
rect 1627 1307 1628 1308
rect 1622 1306 1628 1307
rect 1894 1307 1900 1308
rect 1894 1303 1895 1307
rect 1899 1303 1900 1307
rect 1894 1302 1900 1303
rect 1910 1307 1916 1308
rect 1910 1303 1911 1307
rect 1915 1306 1916 1307
rect 2214 1307 2220 1308
rect 1915 1304 2009 1306
rect 1915 1303 1916 1304
rect 1910 1302 1916 1303
rect 2214 1303 2215 1307
rect 2219 1303 2220 1307
rect 2214 1302 2220 1303
rect 2398 1307 2404 1308
rect 2398 1303 2399 1307
rect 2403 1303 2404 1307
rect 2408 1306 2410 1320
rect 2510 1316 2516 1317
rect 2510 1312 2511 1316
rect 2515 1312 2516 1316
rect 2510 1311 2516 1312
rect 2686 1316 2692 1317
rect 2686 1312 2687 1316
rect 2691 1312 2692 1316
rect 2686 1311 2692 1312
rect 2862 1316 2868 1317
rect 2862 1312 2863 1316
rect 2867 1312 2868 1316
rect 2862 1311 2868 1312
rect 3038 1316 3044 1317
rect 3038 1312 3039 1316
rect 3043 1312 3044 1316
rect 3038 1311 3044 1312
rect 3214 1316 3220 1317
rect 3214 1312 3215 1316
rect 3219 1312 3220 1316
rect 3214 1311 3220 1312
rect 3366 1316 3372 1317
rect 3366 1312 3367 1316
rect 3371 1312 3372 1316
rect 3366 1311 3372 1312
rect 3462 1313 3468 1314
rect 3462 1309 3463 1313
rect 3467 1309 3468 1313
rect 3462 1308 3468 1309
rect 2758 1307 2764 1308
rect 2408 1304 2553 1306
rect 2398 1302 2404 1303
rect 2758 1303 2759 1307
rect 2763 1303 2764 1307
rect 2758 1302 2764 1303
rect 2766 1307 2772 1308
rect 2766 1303 2767 1307
rect 2771 1306 2772 1307
rect 2942 1307 2948 1308
rect 2771 1304 2905 1306
rect 2771 1303 2772 1304
rect 2766 1302 2772 1303
rect 2942 1303 2943 1307
rect 2947 1306 2948 1307
rect 3118 1307 3124 1308
rect 2947 1304 3081 1306
rect 2947 1303 2948 1304
rect 2942 1302 2948 1303
rect 3118 1303 3119 1307
rect 3123 1306 3124 1307
rect 3430 1307 3436 1308
rect 3123 1304 3257 1306
rect 3123 1303 3124 1304
rect 3118 1302 3124 1303
rect 3430 1303 3431 1307
rect 3435 1303 3436 1307
rect 3430 1302 3436 1303
rect 134 1301 140 1302
rect 110 1300 116 1301
rect 110 1296 111 1300
rect 115 1296 116 1300
rect 134 1297 135 1301
rect 139 1297 140 1301
rect 134 1296 140 1297
rect 246 1301 252 1302
rect 246 1297 247 1301
rect 251 1297 252 1301
rect 246 1296 252 1297
rect 398 1301 404 1302
rect 398 1297 399 1301
rect 403 1297 404 1301
rect 398 1296 404 1297
rect 558 1301 564 1302
rect 558 1297 559 1301
rect 563 1297 564 1301
rect 558 1296 564 1297
rect 726 1301 732 1302
rect 726 1297 727 1301
rect 731 1297 732 1301
rect 726 1296 732 1297
rect 894 1301 900 1302
rect 894 1297 895 1301
rect 899 1297 900 1301
rect 894 1296 900 1297
rect 1062 1301 1068 1302
rect 1062 1297 1063 1301
rect 1067 1297 1068 1301
rect 1062 1296 1068 1297
rect 1222 1301 1228 1302
rect 1222 1297 1223 1301
rect 1227 1297 1228 1301
rect 1222 1296 1228 1297
rect 1374 1301 1380 1302
rect 1374 1297 1375 1301
rect 1379 1297 1380 1301
rect 1374 1296 1380 1297
rect 1534 1301 1540 1302
rect 1534 1297 1535 1301
rect 1539 1297 1540 1301
rect 1534 1296 1540 1297
rect 1670 1301 1676 1302
rect 1670 1297 1671 1301
rect 1675 1297 1676 1301
rect 1670 1296 1676 1297
rect 1766 1300 1772 1301
rect 1766 1296 1767 1300
rect 1771 1296 1772 1300
rect 1830 1297 1836 1298
rect 110 1295 116 1296
rect 1766 1295 1772 1296
rect 1806 1296 1812 1297
rect 1806 1292 1807 1296
rect 1811 1292 1812 1296
rect 1830 1293 1831 1297
rect 1835 1293 1836 1297
rect 1830 1292 1836 1293
rect 1966 1297 1972 1298
rect 1966 1293 1967 1297
rect 1971 1293 1972 1297
rect 1966 1292 1972 1293
rect 2142 1297 2148 1298
rect 2142 1293 2143 1297
rect 2147 1293 2148 1297
rect 2142 1292 2148 1293
rect 2326 1297 2332 1298
rect 2326 1293 2327 1297
rect 2331 1293 2332 1297
rect 2326 1292 2332 1293
rect 2510 1297 2516 1298
rect 2510 1293 2511 1297
rect 2515 1293 2516 1297
rect 2510 1292 2516 1293
rect 2686 1297 2692 1298
rect 2686 1293 2687 1297
rect 2691 1293 2692 1297
rect 2686 1292 2692 1293
rect 2862 1297 2868 1298
rect 2862 1293 2863 1297
rect 2867 1293 2868 1297
rect 2862 1292 2868 1293
rect 3038 1297 3044 1298
rect 3038 1293 3039 1297
rect 3043 1293 3044 1297
rect 3038 1292 3044 1293
rect 3214 1297 3220 1298
rect 3214 1293 3215 1297
rect 3219 1293 3220 1297
rect 3214 1292 3220 1293
rect 3366 1297 3372 1298
rect 3366 1293 3367 1297
rect 3371 1293 3372 1297
rect 3366 1292 3372 1293
rect 3462 1296 3468 1297
rect 3462 1292 3463 1296
rect 3467 1292 3468 1296
rect 1806 1291 1812 1292
rect 3462 1291 3468 1292
rect 183 1283 189 1284
rect 183 1279 184 1283
rect 188 1282 189 1283
rect 198 1283 204 1284
rect 198 1282 199 1283
rect 188 1280 199 1282
rect 188 1279 189 1280
rect 183 1278 189 1279
rect 198 1279 199 1280
rect 203 1279 204 1283
rect 198 1278 204 1279
rect 206 1283 212 1284
rect 206 1279 207 1283
rect 211 1282 212 1283
rect 295 1283 301 1284
rect 295 1282 296 1283
rect 211 1280 296 1282
rect 211 1279 212 1280
rect 206 1278 212 1279
rect 295 1279 296 1280
rect 300 1279 301 1283
rect 295 1278 301 1279
rect 318 1283 324 1284
rect 318 1279 319 1283
rect 323 1282 324 1283
rect 447 1283 453 1284
rect 447 1282 448 1283
rect 323 1280 448 1282
rect 323 1279 324 1280
rect 318 1278 324 1279
rect 447 1279 448 1280
rect 452 1279 453 1283
rect 447 1278 453 1279
rect 470 1283 476 1284
rect 470 1279 471 1283
rect 475 1282 476 1283
rect 607 1283 613 1284
rect 607 1282 608 1283
rect 475 1280 608 1282
rect 475 1279 476 1280
rect 470 1278 476 1279
rect 607 1279 608 1280
rect 612 1279 613 1283
rect 607 1278 613 1279
rect 750 1283 756 1284
rect 750 1279 751 1283
rect 755 1282 756 1283
rect 775 1283 781 1284
rect 775 1282 776 1283
rect 755 1280 776 1282
rect 755 1279 756 1280
rect 750 1278 756 1279
rect 775 1279 776 1280
rect 780 1279 781 1283
rect 775 1278 781 1279
rect 798 1283 804 1284
rect 798 1279 799 1283
rect 803 1282 804 1283
rect 943 1283 949 1284
rect 943 1282 944 1283
rect 803 1280 944 1282
rect 803 1279 804 1280
rect 798 1278 804 1279
rect 943 1279 944 1280
rect 948 1279 949 1283
rect 943 1278 949 1279
rect 966 1283 972 1284
rect 966 1279 967 1283
rect 971 1282 972 1283
rect 1111 1283 1117 1284
rect 1111 1282 1112 1283
rect 971 1280 1112 1282
rect 971 1279 972 1280
rect 966 1278 972 1279
rect 1111 1279 1112 1280
rect 1116 1279 1117 1283
rect 1111 1278 1117 1279
rect 1271 1283 1277 1284
rect 1271 1279 1272 1283
rect 1276 1282 1277 1283
rect 1294 1283 1300 1284
rect 1276 1280 1290 1282
rect 1276 1279 1277 1280
rect 1271 1278 1277 1279
rect 1288 1274 1290 1280
rect 1294 1279 1295 1283
rect 1299 1282 1300 1283
rect 1423 1283 1429 1284
rect 1423 1282 1424 1283
rect 1299 1280 1424 1282
rect 1299 1279 1300 1280
rect 1294 1278 1300 1279
rect 1423 1279 1424 1280
rect 1428 1279 1429 1283
rect 1423 1278 1429 1279
rect 1446 1283 1452 1284
rect 1446 1279 1447 1283
rect 1451 1282 1452 1283
rect 1583 1283 1589 1284
rect 1583 1282 1584 1283
rect 1451 1280 1584 1282
rect 1451 1279 1452 1280
rect 1446 1278 1452 1279
rect 1583 1279 1584 1280
rect 1588 1279 1589 1283
rect 1583 1278 1589 1279
rect 1606 1283 1612 1284
rect 1606 1279 1607 1283
rect 1611 1282 1612 1283
rect 1719 1283 1725 1284
rect 1719 1282 1720 1283
rect 1611 1280 1720 1282
rect 1611 1279 1612 1280
rect 1606 1278 1612 1279
rect 1719 1279 1720 1280
rect 1724 1279 1725 1283
rect 1719 1278 1725 1279
rect 1879 1279 1885 1280
rect 1510 1275 1516 1276
rect 1510 1274 1511 1275
rect 1288 1272 1511 1274
rect 1510 1271 1511 1272
rect 1515 1271 1516 1275
rect 1622 1275 1628 1276
rect 1622 1274 1623 1275
rect 1510 1270 1516 1271
rect 1568 1272 1623 1274
rect 183 1267 192 1268
rect 183 1263 184 1267
rect 191 1263 192 1267
rect 183 1262 192 1263
rect 206 1267 212 1268
rect 206 1263 207 1267
rect 211 1266 212 1267
rect 271 1267 277 1268
rect 271 1266 272 1267
rect 211 1264 272 1266
rect 211 1263 212 1264
rect 206 1262 212 1263
rect 271 1263 272 1264
rect 276 1263 277 1267
rect 271 1262 277 1263
rect 294 1267 300 1268
rect 294 1263 295 1267
rect 299 1266 300 1267
rect 367 1267 373 1268
rect 367 1266 368 1267
rect 299 1264 368 1266
rect 299 1263 300 1264
rect 294 1262 300 1263
rect 367 1263 368 1264
rect 372 1263 373 1267
rect 367 1262 373 1263
rect 390 1267 396 1268
rect 390 1263 391 1267
rect 395 1266 396 1267
rect 479 1267 485 1268
rect 479 1266 480 1267
rect 395 1264 480 1266
rect 395 1263 396 1264
rect 390 1262 396 1263
rect 479 1263 480 1264
rect 484 1263 485 1267
rect 479 1262 485 1263
rect 502 1267 508 1268
rect 502 1263 503 1267
rect 507 1266 508 1267
rect 599 1267 605 1268
rect 599 1266 600 1267
rect 507 1264 600 1266
rect 507 1263 508 1264
rect 502 1262 508 1263
rect 599 1263 600 1264
rect 604 1263 605 1267
rect 599 1262 605 1263
rect 727 1267 733 1268
rect 727 1263 728 1267
rect 732 1266 733 1267
rect 758 1267 764 1268
rect 758 1266 759 1267
rect 732 1264 759 1266
rect 732 1263 733 1264
rect 727 1262 733 1263
rect 758 1263 759 1264
rect 763 1263 764 1267
rect 758 1262 764 1263
rect 871 1267 877 1268
rect 871 1263 872 1267
rect 876 1266 877 1267
rect 902 1267 908 1268
rect 902 1266 903 1267
rect 876 1264 903 1266
rect 876 1263 877 1264
rect 871 1262 877 1263
rect 902 1263 903 1264
rect 907 1263 908 1267
rect 902 1262 908 1263
rect 1023 1267 1029 1268
rect 1023 1263 1024 1267
rect 1028 1266 1029 1267
rect 1090 1267 1096 1268
rect 1090 1266 1091 1267
rect 1028 1264 1091 1266
rect 1028 1263 1029 1264
rect 1023 1262 1029 1263
rect 1090 1263 1091 1264
rect 1095 1263 1096 1267
rect 1090 1262 1096 1263
rect 1191 1267 1197 1268
rect 1191 1263 1192 1267
rect 1196 1266 1197 1267
rect 1223 1267 1229 1268
rect 1223 1266 1224 1267
rect 1196 1264 1224 1266
rect 1196 1263 1197 1264
rect 1191 1262 1197 1263
rect 1223 1263 1224 1264
rect 1228 1263 1229 1267
rect 1223 1262 1229 1263
rect 1326 1267 1332 1268
rect 1326 1263 1327 1267
rect 1331 1266 1332 1267
rect 1367 1267 1373 1268
rect 1367 1266 1368 1267
rect 1331 1264 1368 1266
rect 1331 1263 1332 1264
rect 1326 1262 1332 1263
rect 1367 1263 1368 1264
rect 1372 1263 1373 1267
rect 1367 1262 1373 1263
rect 1551 1267 1557 1268
rect 1551 1263 1552 1267
rect 1556 1266 1557 1267
rect 1568 1266 1570 1272
rect 1622 1271 1623 1272
rect 1627 1271 1628 1275
rect 1879 1275 1880 1279
rect 1884 1278 1885 1279
rect 1910 1279 1916 1280
rect 1910 1278 1911 1279
rect 1884 1276 1911 1278
rect 1884 1275 1885 1276
rect 1879 1274 1885 1275
rect 1910 1275 1911 1276
rect 1915 1275 1916 1279
rect 1910 1274 1916 1275
rect 2015 1279 2024 1280
rect 2015 1275 2016 1279
rect 2023 1275 2024 1279
rect 2015 1274 2024 1275
rect 2166 1279 2172 1280
rect 2166 1275 2167 1279
rect 2171 1278 2172 1279
rect 2191 1279 2197 1280
rect 2191 1278 2192 1279
rect 2171 1276 2192 1278
rect 2171 1275 2172 1276
rect 2166 1274 2172 1275
rect 2191 1275 2192 1276
rect 2196 1275 2197 1279
rect 2191 1274 2197 1275
rect 2214 1279 2220 1280
rect 2214 1275 2215 1279
rect 2219 1278 2220 1279
rect 2375 1279 2381 1280
rect 2375 1278 2376 1279
rect 2219 1276 2376 1278
rect 2219 1275 2220 1276
rect 2214 1274 2220 1275
rect 2375 1275 2376 1276
rect 2380 1275 2381 1279
rect 2375 1274 2381 1275
rect 2398 1279 2404 1280
rect 2398 1275 2399 1279
rect 2403 1278 2404 1279
rect 2559 1279 2565 1280
rect 2559 1278 2560 1279
rect 2403 1276 2560 1278
rect 2403 1275 2404 1276
rect 2398 1274 2404 1275
rect 2559 1275 2560 1276
rect 2564 1275 2565 1279
rect 2735 1279 2741 1280
rect 2559 1274 2565 1275
rect 2678 1275 2684 1276
rect 2678 1274 2679 1275
rect 1622 1270 1628 1271
rect 2424 1272 2554 1274
rect 1556 1264 1570 1266
rect 1574 1267 1580 1268
rect 1556 1263 1557 1264
rect 1551 1262 1557 1263
rect 1574 1263 1575 1267
rect 1579 1266 1580 1267
rect 1719 1267 1725 1268
rect 1719 1266 1720 1267
rect 1579 1264 1720 1266
rect 1579 1263 1580 1264
rect 1574 1262 1580 1263
rect 1719 1263 1720 1264
rect 1724 1263 1725 1267
rect 1719 1262 1725 1263
rect 1742 1267 1748 1268
rect 1742 1263 1743 1267
rect 1747 1266 1748 1267
rect 1879 1267 1885 1268
rect 1879 1266 1880 1267
rect 1747 1264 1880 1266
rect 1747 1263 1748 1264
rect 1742 1262 1748 1263
rect 1879 1263 1880 1264
rect 1884 1263 1885 1267
rect 1879 1262 1885 1263
rect 1902 1267 1908 1268
rect 1902 1263 1903 1267
rect 1907 1266 1908 1267
rect 2143 1267 2149 1268
rect 2143 1266 2144 1267
rect 1907 1264 2144 1266
rect 1907 1263 1908 1264
rect 1902 1262 1908 1263
rect 2143 1263 2144 1264
rect 2148 1263 2149 1267
rect 2143 1262 2149 1263
rect 2407 1267 2413 1268
rect 2407 1263 2408 1267
rect 2412 1266 2413 1267
rect 2424 1266 2426 1272
rect 2552 1270 2554 1272
rect 2624 1272 2679 1274
rect 2624 1270 2626 1272
rect 2678 1271 2679 1272
rect 2683 1271 2684 1275
rect 2735 1275 2736 1279
rect 2740 1278 2741 1279
rect 2766 1279 2772 1280
rect 2766 1278 2767 1279
rect 2740 1276 2767 1278
rect 2740 1275 2741 1276
rect 2735 1274 2741 1275
rect 2766 1275 2767 1276
rect 2771 1275 2772 1279
rect 2766 1274 2772 1275
rect 2911 1279 2917 1280
rect 2911 1275 2912 1279
rect 2916 1278 2917 1279
rect 2942 1279 2948 1280
rect 2942 1278 2943 1279
rect 2916 1276 2943 1278
rect 2916 1275 2917 1276
rect 2911 1274 2917 1275
rect 2942 1275 2943 1276
rect 2947 1275 2948 1279
rect 2942 1274 2948 1275
rect 3087 1279 3093 1280
rect 3087 1275 3088 1279
rect 3092 1278 3093 1279
rect 3118 1279 3124 1280
rect 3118 1278 3119 1279
rect 3092 1276 3119 1278
rect 3092 1275 3093 1276
rect 3087 1274 3093 1275
rect 3118 1275 3119 1276
rect 3123 1275 3124 1279
rect 3118 1274 3124 1275
rect 3262 1279 3269 1280
rect 3262 1275 3263 1279
rect 3268 1275 3269 1279
rect 3262 1274 3269 1275
rect 3415 1279 3421 1280
rect 3415 1275 3416 1279
rect 3420 1278 3421 1279
rect 3438 1279 3444 1280
rect 3438 1278 3439 1279
rect 3420 1276 3439 1278
rect 3420 1275 3421 1276
rect 3415 1274 3421 1275
rect 3438 1275 3439 1276
rect 3443 1275 3444 1279
rect 3438 1274 3444 1275
rect 2678 1270 2684 1271
rect 2552 1268 2626 1270
rect 2412 1264 2426 1266
rect 2430 1267 2436 1268
rect 2412 1263 2413 1264
rect 2407 1262 2413 1263
rect 2430 1263 2431 1267
rect 2435 1266 2436 1267
rect 2647 1267 2653 1268
rect 2647 1266 2648 1267
rect 2435 1264 2648 1266
rect 2435 1263 2436 1264
rect 2430 1262 2436 1263
rect 2647 1263 2648 1264
rect 2652 1263 2653 1267
rect 2647 1262 2653 1263
rect 2758 1267 2764 1268
rect 2758 1263 2759 1267
rect 2763 1266 2764 1267
rect 2855 1267 2861 1268
rect 2855 1266 2856 1267
rect 2763 1264 2856 1266
rect 2763 1263 2764 1264
rect 2758 1262 2764 1263
rect 2855 1263 2856 1264
rect 2860 1263 2861 1267
rect 2855 1262 2861 1263
rect 3055 1267 3061 1268
rect 3055 1263 3056 1267
rect 3060 1266 3061 1267
rect 3086 1267 3092 1268
rect 3086 1266 3087 1267
rect 3060 1264 3087 1266
rect 3060 1263 3061 1264
rect 3055 1262 3061 1263
rect 3086 1263 3087 1264
rect 3091 1263 3092 1267
rect 3086 1262 3092 1263
rect 3146 1267 3152 1268
rect 3146 1263 3147 1267
rect 3151 1266 3152 1267
rect 3247 1267 3253 1268
rect 3247 1266 3248 1267
rect 3151 1264 3248 1266
rect 3151 1263 3152 1264
rect 3146 1262 3152 1263
rect 3247 1263 3248 1264
rect 3252 1263 3253 1267
rect 3247 1262 3253 1263
rect 3415 1267 3421 1268
rect 3415 1263 3416 1267
rect 3420 1266 3421 1267
rect 3430 1267 3436 1268
rect 3430 1266 3431 1267
rect 3420 1264 3431 1266
rect 3420 1263 3421 1264
rect 3415 1262 3421 1263
rect 3430 1263 3431 1264
rect 3435 1263 3436 1267
rect 3430 1262 3436 1263
rect 110 1252 116 1253
rect 1766 1252 1772 1253
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 110 1247 116 1248
rect 134 1251 140 1252
rect 134 1247 135 1251
rect 139 1247 140 1251
rect 134 1246 140 1247
rect 222 1251 228 1252
rect 222 1247 223 1251
rect 227 1247 228 1251
rect 222 1246 228 1247
rect 318 1251 324 1252
rect 318 1247 319 1251
rect 323 1247 324 1251
rect 318 1246 324 1247
rect 430 1251 436 1252
rect 430 1247 431 1251
rect 435 1247 436 1251
rect 430 1246 436 1247
rect 550 1251 556 1252
rect 550 1247 551 1251
rect 555 1247 556 1251
rect 550 1246 556 1247
rect 678 1251 684 1252
rect 678 1247 679 1251
rect 683 1247 684 1251
rect 678 1246 684 1247
rect 822 1251 828 1252
rect 822 1247 823 1251
rect 827 1247 828 1251
rect 822 1246 828 1247
rect 974 1251 980 1252
rect 974 1247 975 1251
rect 979 1247 980 1251
rect 974 1246 980 1247
rect 1142 1251 1148 1252
rect 1142 1247 1143 1251
rect 1147 1247 1148 1251
rect 1142 1246 1148 1247
rect 1318 1251 1324 1252
rect 1318 1247 1319 1251
rect 1323 1247 1324 1251
rect 1318 1246 1324 1247
rect 1502 1251 1508 1252
rect 1502 1247 1503 1251
rect 1507 1247 1508 1251
rect 1502 1246 1508 1247
rect 1670 1251 1676 1252
rect 1670 1247 1671 1251
rect 1675 1247 1676 1251
rect 1766 1248 1767 1252
rect 1771 1248 1772 1252
rect 1766 1247 1772 1248
rect 1806 1252 1812 1253
rect 3462 1252 3468 1253
rect 1806 1248 1807 1252
rect 1811 1248 1812 1252
rect 1806 1247 1812 1248
rect 1830 1251 1836 1252
rect 1830 1247 1831 1251
rect 1835 1247 1836 1251
rect 1670 1246 1676 1247
rect 1830 1246 1836 1247
rect 2094 1251 2100 1252
rect 2094 1247 2095 1251
rect 2099 1247 2100 1251
rect 2094 1246 2100 1247
rect 2358 1251 2364 1252
rect 2358 1247 2359 1251
rect 2363 1247 2364 1251
rect 2358 1246 2364 1247
rect 2598 1251 2604 1252
rect 2598 1247 2599 1251
rect 2603 1247 2604 1251
rect 2598 1246 2604 1247
rect 2806 1251 2812 1252
rect 2806 1247 2807 1251
rect 2811 1247 2812 1251
rect 2806 1246 2812 1247
rect 3006 1251 3012 1252
rect 3006 1247 3007 1251
rect 3011 1247 3012 1251
rect 3006 1246 3012 1247
rect 3198 1251 3204 1252
rect 3198 1247 3199 1251
rect 3203 1247 3204 1251
rect 3366 1251 3372 1252
rect 3198 1246 3204 1247
rect 3262 1247 3268 1248
rect 206 1243 212 1244
rect 206 1239 207 1243
rect 211 1239 212 1243
rect 206 1238 212 1239
rect 294 1243 300 1244
rect 294 1239 295 1243
rect 299 1239 300 1243
rect 294 1238 300 1239
rect 390 1243 396 1244
rect 390 1239 391 1243
rect 395 1239 396 1243
rect 390 1238 396 1239
rect 502 1243 508 1244
rect 502 1239 503 1243
rect 507 1239 508 1243
rect 502 1238 508 1239
rect 510 1243 516 1244
rect 510 1239 511 1243
rect 515 1242 516 1243
rect 750 1243 756 1244
rect 515 1240 593 1242
rect 515 1239 516 1240
rect 510 1238 516 1239
rect 750 1239 751 1243
rect 755 1239 756 1243
rect 750 1238 756 1239
rect 758 1243 764 1244
rect 758 1239 759 1243
rect 763 1242 764 1243
rect 902 1243 908 1244
rect 763 1240 865 1242
rect 763 1239 764 1240
rect 758 1238 764 1239
rect 902 1239 903 1243
rect 907 1242 908 1243
rect 1090 1243 1096 1244
rect 907 1240 1017 1242
rect 907 1239 908 1240
rect 902 1238 908 1239
rect 1090 1239 1091 1243
rect 1095 1242 1096 1243
rect 1223 1243 1229 1244
rect 1095 1240 1185 1242
rect 1095 1239 1096 1240
rect 1090 1238 1096 1239
rect 1223 1239 1224 1243
rect 1228 1242 1229 1243
rect 1574 1243 1580 1244
rect 1228 1240 1361 1242
rect 1228 1239 1229 1240
rect 1223 1238 1229 1239
rect 1574 1239 1575 1243
rect 1579 1239 1580 1243
rect 1574 1238 1580 1239
rect 1742 1243 1748 1244
rect 1742 1239 1743 1243
rect 1747 1239 1748 1243
rect 1742 1238 1748 1239
rect 1902 1243 1908 1244
rect 1902 1239 1903 1243
rect 1907 1239 1908 1243
rect 1902 1238 1908 1239
rect 2166 1243 2172 1244
rect 2166 1239 2167 1243
rect 2171 1239 2172 1243
rect 2166 1238 2172 1239
rect 2430 1243 2436 1244
rect 2430 1239 2431 1243
rect 2435 1239 2436 1243
rect 2678 1243 2684 1244
rect 2430 1238 2436 1239
rect 2670 1239 2676 1240
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 1766 1235 1772 1236
rect 110 1230 116 1231
rect 134 1232 140 1233
rect 134 1228 135 1232
rect 139 1228 140 1232
rect 134 1227 140 1228
rect 222 1232 228 1233
rect 222 1228 223 1232
rect 227 1228 228 1232
rect 222 1227 228 1228
rect 318 1232 324 1233
rect 318 1228 319 1232
rect 323 1228 324 1232
rect 318 1227 324 1228
rect 430 1232 436 1233
rect 430 1228 431 1232
rect 435 1228 436 1232
rect 430 1227 436 1228
rect 550 1232 556 1233
rect 550 1228 551 1232
rect 555 1228 556 1232
rect 550 1227 556 1228
rect 678 1232 684 1233
rect 678 1228 679 1232
rect 683 1228 684 1232
rect 678 1227 684 1228
rect 822 1232 828 1233
rect 822 1228 823 1232
rect 827 1228 828 1232
rect 822 1227 828 1228
rect 974 1232 980 1233
rect 974 1228 975 1232
rect 979 1228 980 1232
rect 974 1227 980 1228
rect 1142 1232 1148 1233
rect 1142 1228 1143 1232
rect 1147 1228 1148 1232
rect 1142 1227 1148 1228
rect 1318 1232 1324 1233
rect 1318 1228 1319 1232
rect 1323 1228 1324 1232
rect 1318 1227 1324 1228
rect 1502 1232 1508 1233
rect 1502 1228 1503 1232
rect 1507 1228 1508 1232
rect 1502 1227 1508 1228
rect 1670 1232 1676 1233
rect 1670 1228 1671 1232
rect 1675 1228 1676 1232
rect 1766 1231 1767 1235
rect 1771 1231 1772 1235
rect 1766 1230 1772 1231
rect 1806 1235 1812 1236
rect 1806 1231 1807 1235
rect 1811 1231 1812 1235
rect 2670 1235 2671 1239
rect 2675 1235 2676 1239
rect 2678 1239 2679 1243
rect 2683 1242 2684 1243
rect 3146 1243 3152 1244
rect 3146 1242 3147 1243
rect 2683 1240 2849 1242
rect 3081 1240 3147 1242
rect 2683 1239 2684 1240
rect 2678 1238 2684 1239
rect 3146 1239 3147 1240
rect 3151 1239 3152 1243
rect 3262 1243 3263 1247
rect 3267 1243 3268 1247
rect 3366 1247 3367 1251
rect 3371 1247 3372 1251
rect 3462 1248 3463 1252
rect 3467 1248 3468 1252
rect 3462 1247 3468 1248
rect 3366 1246 3372 1247
rect 3262 1242 3268 1243
rect 3264 1240 3273 1242
rect 3146 1238 3152 1239
rect 3438 1239 3444 1240
rect 2670 1234 2676 1235
rect 3438 1235 3439 1239
rect 3443 1235 3444 1239
rect 3438 1234 3444 1235
rect 3462 1235 3468 1236
rect 1806 1230 1812 1231
rect 1830 1232 1836 1233
rect 1670 1227 1676 1228
rect 1830 1228 1831 1232
rect 1835 1228 1836 1232
rect 1830 1227 1836 1228
rect 2094 1232 2100 1233
rect 2094 1228 2095 1232
rect 2099 1228 2100 1232
rect 2094 1227 2100 1228
rect 2358 1232 2364 1233
rect 2358 1228 2359 1232
rect 2363 1228 2364 1232
rect 2358 1227 2364 1228
rect 2598 1232 2604 1233
rect 2598 1228 2599 1232
rect 2603 1228 2604 1232
rect 2598 1227 2604 1228
rect 2806 1232 2812 1233
rect 2806 1228 2807 1232
rect 2811 1228 2812 1232
rect 2806 1227 2812 1228
rect 3006 1232 3012 1233
rect 3006 1228 3007 1232
rect 3011 1228 3012 1232
rect 3006 1227 3012 1228
rect 3198 1232 3204 1233
rect 3198 1228 3199 1232
rect 3203 1228 3204 1232
rect 3198 1227 3204 1228
rect 3366 1232 3372 1233
rect 3366 1228 3367 1232
rect 3371 1228 3372 1232
rect 3462 1231 3463 1235
rect 3467 1231 3468 1235
rect 3462 1230 3468 1231
rect 3366 1227 3372 1228
rect 186 1195 192 1196
rect 186 1191 187 1195
rect 191 1194 192 1195
rect 510 1195 516 1196
rect 510 1194 511 1195
rect 191 1192 511 1194
rect 191 1191 192 1192
rect 186 1190 192 1191
rect 510 1191 511 1192
rect 515 1191 516 1195
rect 510 1190 516 1191
rect 134 1180 140 1181
rect 110 1177 116 1178
rect 110 1173 111 1177
rect 115 1173 116 1177
rect 134 1176 135 1180
rect 139 1176 140 1180
rect 134 1175 140 1176
rect 230 1180 236 1181
rect 230 1176 231 1180
rect 235 1176 236 1180
rect 230 1175 236 1176
rect 358 1180 364 1181
rect 358 1176 359 1180
rect 363 1176 364 1180
rect 358 1175 364 1176
rect 486 1180 492 1181
rect 486 1176 487 1180
rect 491 1176 492 1180
rect 486 1175 492 1176
rect 614 1180 620 1181
rect 614 1176 615 1180
rect 619 1176 620 1180
rect 614 1175 620 1176
rect 742 1180 748 1181
rect 742 1176 743 1180
rect 747 1176 748 1180
rect 742 1175 748 1176
rect 870 1180 876 1181
rect 870 1176 871 1180
rect 875 1176 876 1180
rect 870 1175 876 1176
rect 990 1180 996 1181
rect 990 1176 991 1180
rect 995 1176 996 1180
rect 990 1175 996 1176
rect 1118 1180 1124 1181
rect 1118 1176 1119 1180
rect 1123 1176 1124 1180
rect 1118 1175 1124 1176
rect 1246 1180 1252 1181
rect 1246 1176 1247 1180
rect 1251 1176 1252 1180
rect 1934 1180 1940 1181
rect 1246 1175 1252 1176
rect 1766 1177 1772 1178
rect 110 1172 116 1173
rect 1766 1173 1767 1177
rect 1771 1173 1772 1177
rect 1766 1172 1772 1173
rect 1806 1177 1812 1178
rect 1806 1173 1807 1177
rect 1811 1173 1812 1177
rect 1934 1176 1935 1180
rect 1939 1176 1940 1180
rect 1934 1175 1940 1176
rect 2038 1180 2044 1181
rect 2038 1176 2039 1180
rect 2043 1176 2044 1180
rect 2038 1175 2044 1176
rect 2158 1180 2164 1181
rect 2158 1176 2159 1180
rect 2163 1176 2164 1180
rect 2158 1175 2164 1176
rect 2286 1180 2292 1181
rect 2286 1176 2287 1180
rect 2291 1176 2292 1180
rect 2286 1175 2292 1176
rect 2422 1180 2428 1181
rect 2422 1176 2423 1180
rect 2427 1176 2428 1180
rect 2422 1175 2428 1176
rect 2566 1180 2572 1181
rect 2566 1176 2567 1180
rect 2571 1176 2572 1180
rect 2566 1175 2572 1176
rect 2702 1180 2708 1181
rect 2702 1176 2703 1180
rect 2707 1176 2708 1180
rect 2702 1175 2708 1176
rect 2838 1180 2844 1181
rect 2838 1176 2839 1180
rect 2843 1176 2844 1180
rect 2838 1175 2844 1176
rect 2974 1180 2980 1181
rect 2974 1176 2975 1180
rect 2979 1176 2980 1180
rect 2974 1175 2980 1176
rect 3110 1180 3116 1181
rect 3110 1176 3111 1180
rect 3115 1176 3116 1180
rect 3110 1175 3116 1176
rect 3246 1180 3252 1181
rect 3246 1176 3247 1180
rect 3251 1176 3252 1180
rect 3246 1175 3252 1176
rect 3366 1180 3372 1181
rect 3366 1176 3367 1180
rect 3371 1176 3372 1180
rect 3366 1175 3372 1176
rect 3462 1177 3468 1178
rect 1806 1172 1812 1173
rect 3462 1173 3463 1177
rect 3467 1173 3468 1177
rect 3462 1172 3468 1173
rect 206 1171 212 1172
rect 206 1167 207 1171
rect 211 1167 212 1171
rect 206 1166 212 1167
rect 302 1171 308 1172
rect 302 1167 303 1171
rect 307 1167 308 1171
rect 302 1166 308 1167
rect 430 1171 436 1172
rect 430 1167 431 1171
rect 435 1167 436 1171
rect 430 1166 436 1167
rect 558 1171 564 1172
rect 558 1167 559 1171
rect 563 1167 564 1171
rect 558 1166 564 1167
rect 566 1171 572 1172
rect 566 1167 567 1171
rect 571 1170 572 1171
rect 814 1171 820 1172
rect 571 1168 657 1170
rect 571 1167 572 1168
rect 566 1166 572 1167
rect 814 1167 815 1171
rect 819 1167 820 1171
rect 814 1166 820 1167
rect 942 1171 948 1172
rect 942 1167 943 1171
rect 947 1167 948 1171
rect 942 1166 948 1167
rect 1062 1171 1068 1172
rect 1062 1167 1063 1171
rect 1067 1167 1068 1171
rect 1062 1166 1068 1167
rect 1190 1171 1196 1172
rect 1190 1167 1191 1171
rect 1195 1167 1196 1171
rect 1326 1171 1332 1172
rect 1326 1170 1327 1171
rect 1321 1168 1327 1170
rect 1190 1166 1196 1167
rect 1326 1167 1327 1168
rect 1331 1167 1332 1171
rect 1326 1166 1332 1167
rect 2002 1171 2008 1172
rect 2002 1167 2003 1171
rect 2007 1167 2008 1171
rect 2002 1166 2008 1167
rect 2014 1171 2020 1172
rect 2014 1167 2015 1171
rect 2019 1170 2020 1171
rect 2118 1171 2124 1172
rect 2019 1168 2081 1170
rect 2019 1167 2020 1168
rect 2014 1166 2020 1167
rect 2118 1167 2119 1171
rect 2123 1170 2124 1171
rect 2238 1171 2244 1172
rect 2123 1168 2201 1170
rect 2123 1167 2124 1168
rect 2118 1166 2124 1167
rect 2238 1167 2239 1171
rect 2243 1170 2244 1171
rect 2366 1171 2372 1172
rect 2243 1168 2329 1170
rect 2243 1167 2244 1168
rect 2238 1166 2244 1167
rect 2366 1167 2367 1171
rect 2371 1170 2372 1171
rect 2502 1171 2508 1172
rect 2371 1168 2465 1170
rect 2371 1167 2372 1168
rect 2366 1166 2372 1167
rect 2502 1167 2503 1171
rect 2507 1170 2508 1171
rect 2774 1171 2780 1172
rect 2507 1168 2609 1170
rect 2507 1167 2508 1168
rect 2502 1166 2508 1167
rect 2774 1167 2775 1171
rect 2779 1167 2780 1171
rect 2774 1166 2780 1167
rect 2910 1171 2916 1172
rect 2910 1167 2911 1171
rect 2915 1167 2916 1171
rect 2910 1166 2916 1167
rect 3046 1171 3052 1172
rect 3046 1167 3047 1171
rect 3051 1167 3052 1171
rect 3046 1166 3052 1167
rect 3086 1171 3092 1172
rect 3086 1167 3087 1171
rect 3091 1170 3092 1171
rect 3190 1171 3196 1172
rect 3091 1168 3153 1170
rect 3091 1167 3092 1168
rect 3086 1166 3092 1167
rect 3190 1167 3191 1171
rect 3195 1170 3196 1171
rect 3430 1171 3436 1172
rect 3195 1168 3289 1170
rect 3195 1167 3196 1168
rect 3190 1166 3196 1167
rect 3430 1167 3431 1171
rect 3435 1167 3436 1171
rect 3430 1166 3436 1167
rect 134 1161 140 1162
rect 110 1160 116 1161
rect 110 1156 111 1160
rect 115 1156 116 1160
rect 134 1157 135 1161
rect 139 1157 140 1161
rect 134 1156 140 1157
rect 230 1161 236 1162
rect 230 1157 231 1161
rect 235 1157 236 1161
rect 230 1156 236 1157
rect 358 1161 364 1162
rect 358 1157 359 1161
rect 363 1157 364 1161
rect 358 1156 364 1157
rect 486 1161 492 1162
rect 486 1157 487 1161
rect 491 1157 492 1161
rect 486 1156 492 1157
rect 614 1161 620 1162
rect 614 1157 615 1161
rect 619 1157 620 1161
rect 614 1156 620 1157
rect 742 1161 748 1162
rect 742 1157 743 1161
rect 747 1157 748 1161
rect 742 1156 748 1157
rect 870 1161 876 1162
rect 870 1157 871 1161
rect 875 1157 876 1161
rect 870 1156 876 1157
rect 990 1161 996 1162
rect 990 1157 991 1161
rect 995 1157 996 1161
rect 990 1156 996 1157
rect 1118 1161 1124 1162
rect 1118 1157 1119 1161
rect 1123 1157 1124 1161
rect 1118 1156 1124 1157
rect 1246 1161 1252 1162
rect 1934 1161 1940 1162
rect 1246 1157 1247 1161
rect 1251 1157 1252 1161
rect 1246 1156 1252 1157
rect 1766 1160 1772 1161
rect 1766 1156 1767 1160
rect 1771 1156 1772 1160
rect 110 1155 116 1156
rect 1766 1155 1772 1156
rect 1806 1160 1812 1161
rect 1806 1156 1807 1160
rect 1811 1156 1812 1160
rect 1934 1157 1935 1161
rect 1939 1157 1940 1161
rect 1934 1156 1940 1157
rect 2038 1161 2044 1162
rect 2038 1157 2039 1161
rect 2043 1157 2044 1161
rect 2038 1156 2044 1157
rect 2158 1161 2164 1162
rect 2158 1157 2159 1161
rect 2163 1157 2164 1161
rect 2158 1156 2164 1157
rect 2286 1161 2292 1162
rect 2286 1157 2287 1161
rect 2291 1157 2292 1161
rect 2286 1156 2292 1157
rect 2422 1161 2428 1162
rect 2422 1157 2423 1161
rect 2427 1157 2428 1161
rect 2422 1156 2428 1157
rect 2566 1161 2572 1162
rect 2566 1157 2567 1161
rect 2571 1157 2572 1161
rect 2566 1156 2572 1157
rect 2702 1161 2708 1162
rect 2702 1157 2703 1161
rect 2707 1157 2708 1161
rect 2702 1156 2708 1157
rect 2838 1161 2844 1162
rect 2838 1157 2839 1161
rect 2843 1157 2844 1161
rect 2838 1156 2844 1157
rect 2974 1161 2980 1162
rect 2974 1157 2975 1161
rect 2979 1157 2980 1161
rect 2974 1156 2980 1157
rect 3110 1161 3116 1162
rect 3110 1157 3111 1161
rect 3115 1157 3116 1161
rect 3110 1156 3116 1157
rect 3246 1161 3252 1162
rect 3246 1157 3247 1161
rect 3251 1157 3252 1161
rect 3246 1156 3252 1157
rect 3366 1161 3372 1162
rect 3366 1157 3367 1161
rect 3371 1157 3372 1161
rect 3366 1156 3372 1157
rect 3462 1160 3468 1161
rect 3462 1156 3463 1160
rect 3467 1156 3468 1160
rect 1806 1155 1812 1156
rect 3462 1155 3468 1156
rect 183 1143 192 1144
rect 183 1139 184 1143
rect 191 1139 192 1143
rect 183 1138 192 1139
rect 206 1143 212 1144
rect 206 1139 207 1143
rect 211 1142 212 1143
rect 279 1143 285 1144
rect 279 1142 280 1143
rect 211 1140 280 1142
rect 211 1139 212 1140
rect 206 1138 212 1139
rect 279 1139 280 1140
rect 284 1139 285 1143
rect 279 1138 285 1139
rect 302 1143 308 1144
rect 302 1139 303 1143
rect 307 1142 308 1143
rect 407 1143 413 1144
rect 407 1142 408 1143
rect 307 1140 408 1142
rect 307 1139 308 1140
rect 302 1138 308 1139
rect 407 1139 408 1140
rect 412 1139 413 1143
rect 407 1138 413 1139
rect 430 1143 436 1144
rect 430 1139 431 1143
rect 435 1142 436 1143
rect 535 1143 541 1144
rect 535 1142 536 1143
rect 435 1140 536 1142
rect 435 1139 436 1140
rect 430 1138 436 1139
rect 535 1139 536 1140
rect 540 1139 541 1143
rect 535 1138 541 1139
rect 558 1143 564 1144
rect 558 1139 559 1143
rect 563 1142 564 1143
rect 663 1143 669 1144
rect 663 1142 664 1143
rect 563 1140 664 1142
rect 563 1139 564 1140
rect 558 1138 564 1139
rect 663 1139 664 1140
rect 668 1139 669 1143
rect 663 1138 669 1139
rect 791 1143 797 1144
rect 791 1139 792 1143
rect 796 1142 797 1143
rect 814 1143 820 1144
rect 796 1140 810 1142
rect 796 1139 797 1140
rect 791 1138 797 1139
rect 566 1135 572 1136
rect 566 1134 567 1135
rect 308 1132 567 1134
rect 295 1127 301 1128
rect 295 1123 296 1127
rect 300 1126 301 1127
rect 308 1126 310 1132
rect 566 1131 567 1132
rect 571 1131 572 1135
rect 808 1134 810 1140
rect 814 1139 815 1143
rect 819 1142 820 1143
rect 919 1143 925 1144
rect 919 1142 920 1143
rect 819 1140 920 1142
rect 819 1139 820 1140
rect 814 1138 820 1139
rect 919 1139 920 1140
rect 924 1139 925 1143
rect 919 1138 925 1139
rect 942 1143 948 1144
rect 942 1139 943 1143
rect 947 1142 948 1143
rect 1039 1143 1045 1144
rect 1039 1142 1040 1143
rect 947 1140 1040 1142
rect 947 1139 948 1140
rect 942 1138 948 1139
rect 1039 1139 1040 1140
rect 1044 1139 1045 1143
rect 1039 1138 1045 1139
rect 1062 1143 1068 1144
rect 1062 1139 1063 1143
rect 1067 1142 1068 1143
rect 1167 1143 1173 1144
rect 1167 1142 1168 1143
rect 1067 1140 1168 1142
rect 1067 1139 1068 1140
rect 1062 1138 1068 1139
rect 1167 1139 1168 1140
rect 1172 1139 1173 1143
rect 1167 1138 1173 1139
rect 1190 1143 1196 1144
rect 1190 1139 1191 1143
rect 1195 1142 1196 1143
rect 1295 1143 1301 1144
rect 1295 1142 1296 1143
rect 1195 1140 1296 1142
rect 1195 1139 1196 1140
rect 1190 1138 1196 1139
rect 1295 1139 1296 1140
rect 1300 1139 1301 1143
rect 1295 1138 1301 1139
rect 1983 1143 1989 1144
rect 1983 1139 1984 1143
rect 1988 1142 1989 1143
rect 2014 1143 2020 1144
rect 2014 1142 2015 1143
rect 1988 1140 2015 1142
rect 1988 1139 1989 1140
rect 1983 1138 1989 1139
rect 2014 1139 2015 1140
rect 2019 1139 2020 1143
rect 2014 1138 2020 1139
rect 2087 1143 2093 1144
rect 2087 1139 2088 1143
rect 2092 1142 2093 1143
rect 2118 1143 2124 1144
rect 2118 1142 2119 1143
rect 2092 1140 2119 1142
rect 2092 1139 2093 1140
rect 2087 1138 2093 1139
rect 2118 1139 2119 1140
rect 2123 1139 2124 1143
rect 2118 1138 2124 1139
rect 2207 1143 2213 1144
rect 2207 1139 2208 1143
rect 2212 1142 2213 1143
rect 2238 1143 2244 1144
rect 2238 1142 2239 1143
rect 2212 1140 2239 1142
rect 2212 1139 2213 1140
rect 2207 1138 2213 1139
rect 2238 1139 2239 1140
rect 2243 1139 2244 1143
rect 2238 1138 2244 1139
rect 2335 1143 2341 1144
rect 2335 1139 2336 1143
rect 2340 1142 2341 1143
rect 2366 1143 2372 1144
rect 2366 1142 2367 1143
rect 2340 1140 2367 1142
rect 2340 1139 2341 1140
rect 2335 1138 2341 1139
rect 2366 1139 2367 1140
rect 2371 1139 2372 1143
rect 2366 1138 2372 1139
rect 2471 1143 2477 1144
rect 2471 1139 2472 1143
rect 2476 1142 2477 1143
rect 2502 1143 2508 1144
rect 2502 1142 2503 1143
rect 2476 1140 2503 1142
rect 2476 1139 2477 1140
rect 2471 1138 2477 1139
rect 2502 1139 2503 1140
rect 2507 1139 2508 1143
rect 2502 1138 2508 1139
rect 2526 1143 2532 1144
rect 2526 1139 2527 1143
rect 2531 1142 2532 1143
rect 2615 1143 2621 1144
rect 2615 1142 2616 1143
rect 2531 1140 2616 1142
rect 2531 1139 2532 1140
rect 2526 1138 2532 1139
rect 2615 1139 2616 1140
rect 2620 1139 2621 1143
rect 2615 1138 2621 1139
rect 2670 1143 2676 1144
rect 2670 1139 2671 1143
rect 2675 1142 2676 1143
rect 2751 1143 2757 1144
rect 2751 1142 2752 1143
rect 2675 1140 2752 1142
rect 2675 1139 2676 1140
rect 2670 1138 2676 1139
rect 2751 1139 2752 1140
rect 2756 1139 2757 1143
rect 2751 1138 2757 1139
rect 2774 1143 2780 1144
rect 2774 1139 2775 1143
rect 2779 1142 2780 1143
rect 2887 1143 2893 1144
rect 2887 1142 2888 1143
rect 2779 1140 2888 1142
rect 2779 1139 2780 1140
rect 2774 1138 2780 1139
rect 2887 1139 2888 1140
rect 2892 1139 2893 1143
rect 2887 1138 2893 1139
rect 2910 1143 2916 1144
rect 2910 1139 2911 1143
rect 2915 1142 2916 1143
rect 3023 1143 3029 1144
rect 3023 1142 3024 1143
rect 2915 1140 3024 1142
rect 2915 1139 2916 1140
rect 2910 1138 2916 1139
rect 3023 1139 3024 1140
rect 3028 1139 3029 1143
rect 3023 1138 3029 1139
rect 3159 1143 3165 1144
rect 3159 1139 3160 1143
rect 3164 1142 3165 1143
rect 3190 1143 3196 1144
rect 3190 1142 3191 1143
rect 3164 1140 3191 1142
rect 3164 1139 3165 1140
rect 3159 1138 3165 1139
rect 3190 1139 3191 1140
rect 3195 1139 3196 1143
rect 3190 1138 3196 1139
rect 3294 1143 3301 1144
rect 3294 1139 3295 1143
rect 3300 1139 3301 1143
rect 3294 1138 3301 1139
rect 3415 1143 3421 1144
rect 3415 1139 3416 1143
rect 3420 1142 3421 1143
rect 3438 1143 3444 1144
rect 3438 1142 3439 1143
rect 3420 1140 3439 1142
rect 3420 1139 3421 1140
rect 3415 1138 3421 1139
rect 3438 1139 3439 1140
rect 3443 1139 3444 1143
rect 3438 1138 3444 1139
rect 838 1135 844 1136
rect 838 1134 839 1135
rect 808 1132 839 1134
rect 566 1130 572 1131
rect 838 1131 839 1132
rect 843 1131 844 1135
rect 838 1130 844 1131
rect 2830 1131 2836 1132
rect 2830 1130 2831 1131
rect 2664 1128 2831 1130
rect 300 1124 310 1126
rect 318 1127 324 1128
rect 300 1123 301 1124
rect 295 1122 301 1123
rect 318 1123 319 1127
rect 323 1126 324 1127
rect 415 1127 421 1128
rect 415 1126 416 1127
rect 323 1124 416 1126
rect 323 1123 324 1124
rect 318 1122 324 1123
rect 415 1123 416 1124
rect 420 1123 421 1127
rect 415 1122 421 1123
rect 438 1127 444 1128
rect 438 1123 439 1127
rect 443 1126 444 1127
rect 543 1127 549 1128
rect 543 1126 544 1127
rect 443 1124 544 1126
rect 443 1123 444 1124
rect 438 1122 444 1123
rect 543 1123 544 1124
rect 548 1123 549 1127
rect 543 1122 549 1123
rect 566 1127 572 1128
rect 566 1123 567 1127
rect 571 1126 572 1127
rect 671 1127 677 1128
rect 671 1126 672 1127
rect 571 1124 672 1126
rect 571 1123 572 1124
rect 566 1122 572 1123
rect 671 1123 672 1124
rect 676 1123 677 1127
rect 671 1122 677 1123
rect 694 1127 700 1128
rect 694 1123 695 1127
rect 699 1126 700 1127
rect 807 1127 813 1128
rect 807 1126 808 1127
rect 699 1124 808 1126
rect 699 1123 700 1124
rect 694 1122 700 1123
rect 807 1123 808 1124
rect 812 1123 813 1127
rect 807 1122 813 1123
rect 935 1127 941 1128
rect 935 1123 936 1127
rect 940 1126 941 1127
rect 998 1127 1004 1128
rect 998 1126 999 1127
rect 940 1124 999 1126
rect 940 1123 941 1124
rect 935 1122 941 1123
rect 998 1123 999 1124
rect 1003 1123 1004 1127
rect 998 1122 1004 1123
rect 1063 1127 1069 1128
rect 1063 1123 1064 1127
rect 1068 1126 1069 1127
rect 1110 1127 1116 1128
rect 1110 1126 1111 1127
rect 1068 1124 1111 1126
rect 1068 1123 1069 1124
rect 1063 1122 1069 1123
rect 1110 1123 1111 1124
rect 1115 1123 1116 1127
rect 1110 1122 1116 1123
rect 1191 1127 1197 1128
rect 1191 1123 1192 1127
rect 1196 1126 1197 1127
rect 1222 1127 1228 1128
rect 1222 1126 1223 1127
rect 1196 1124 1223 1126
rect 1196 1123 1197 1124
rect 1191 1122 1197 1123
rect 1222 1123 1223 1124
rect 1227 1123 1228 1127
rect 1222 1122 1228 1123
rect 1319 1127 1325 1128
rect 1319 1123 1320 1127
rect 1324 1126 1325 1127
rect 1350 1127 1356 1128
rect 1350 1126 1351 1127
rect 1324 1124 1351 1126
rect 1324 1123 1325 1124
rect 1319 1122 1325 1123
rect 1350 1123 1351 1124
rect 1355 1123 1356 1127
rect 1350 1122 1356 1123
rect 1382 1127 1388 1128
rect 1382 1123 1383 1127
rect 1387 1126 1388 1127
rect 1447 1127 1453 1128
rect 1447 1126 1448 1127
rect 1387 1124 1448 1126
rect 1387 1123 1388 1124
rect 1382 1122 1388 1123
rect 1447 1123 1448 1124
rect 1452 1123 1453 1127
rect 2002 1127 2008 1128
rect 2002 1126 2003 1127
rect 1447 1122 1453 1123
rect 1991 1125 2003 1126
rect 1991 1121 1992 1125
rect 1996 1124 2003 1125
rect 1996 1121 1997 1124
rect 2002 1123 2003 1124
rect 2007 1123 2008 1127
rect 2002 1122 2008 1123
rect 2014 1123 2020 1124
rect 1991 1120 1997 1121
rect 2014 1119 2015 1123
rect 2019 1122 2020 1123
rect 2111 1123 2117 1124
rect 2111 1122 2112 1123
rect 2019 1120 2112 1122
rect 2019 1119 2020 1120
rect 2014 1118 2020 1119
rect 2111 1119 2112 1120
rect 2116 1119 2117 1123
rect 2111 1118 2117 1119
rect 2134 1123 2140 1124
rect 2134 1119 2135 1123
rect 2139 1122 2140 1123
rect 2239 1123 2245 1124
rect 2239 1122 2240 1123
rect 2139 1120 2240 1122
rect 2139 1119 2140 1120
rect 2134 1118 2140 1119
rect 2239 1119 2240 1120
rect 2244 1119 2245 1123
rect 2239 1118 2245 1119
rect 2367 1123 2376 1124
rect 2367 1119 2368 1123
rect 2375 1119 2376 1123
rect 2367 1118 2376 1119
rect 2390 1123 2396 1124
rect 2390 1119 2391 1123
rect 2395 1122 2396 1123
rect 2503 1123 2509 1124
rect 2503 1122 2504 1123
rect 2395 1120 2504 1122
rect 2395 1119 2396 1120
rect 2390 1118 2396 1119
rect 2503 1119 2504 1120
rect 2508 1119 2509 1123
rect 2503 1118 2509 1119
rect 2647 1123 2653 1124
rect 2647 1119 2648 1123
rect 2652 1122 2653 1123
rect 2664 1122 2666 1128
rect 2830 1127 2831 1128
rect 2835 1127 2836 1131
rect 2830 1126 2836 1127
rect 2652 1120 2666 1122
rect 2670 1123 2676 1124
rect 2652 1119 2653 1120
rect 2647 1118 2653 1119
rect 2670 1119 2671 1123
rect 2675 1122 2676 1123
rect 2799 1123 2805 1124
rect 2799 1122 2800 1123
rect 2675 1120 2800 1122
rect 2675 1119 2676 1120
rect 2670 1118 2676 1119
rect 2799 1119 2800 1120
rect 2804 1119 2805 1123
rect 2799 1118 2805 1119
rect 2951 1123 2957 1124
rect 2951 1119 2952 1123
rect 2956 1122 2957 1123
rect 2982 1123 2988 1124
rect 2982 1122 2983 1123
rect 2956 1120 2983 1122
rect 2956 1119 2957 1120
rect 2951 1118 2957 1119
rect 2982 1119 2983 1120
rect 2987 1119 2988 1123
rect 2982 1118 2988 1119
rect 3046 1123 3052 1124
rect 3046 1119 3047 1123
rect 3051 1122 3052 1123
rect 3111 1123 3117 1124
rect 3111 1122 3112 1123
rect 3051 1120 3112 1122
rect 3051 1119 3052 1120
rect 3046 1118 3052 1119
rect 3111 1119 3112 1120
rect 3116 1119 3117 1123
rect 3111 1118 3117 1119
rect 3270 1123 3277 1124
rect 3270 1119 3271 1123
rect 3276 1119 3277 1123
rect 3270 1118 3277 1119
rect 3415 1123 3421 1124
rect 3415 1119 3416 1123
rect 3420 1122 3421 1123
rect 3430 1123 3436 1124
rect 3430 1122 3431 1123
rect 3420 1120 3431 1122
rect 3420 1119 3421 1120
rect 3415 1118 3421 1119
rect 3430 1119 3431 1120
rect 3435 1119 3436 1123
rect 3430 1118 3436 1119
rect 110 1112 116 1113
rect 1766 1112 1772 1113
rect 110 1108 111 1112
rect 115 1108 116 1112
rect 110 1107 116 1108
rect 246 1111 252 1112
rect 246 1107 247 1111
rect 251 1107 252 1111
rect 246 1106 252 1107
rect 366 1111 372 1112
rect 366 1107 367 1111
rect 371 1107 372 1111
rect 366 1106 372 1107
rect 494 1111 500 1112
rect 494 1107 495 1111
rect 499 1107 500 1111
rect 494 1106 500 1107
rect 622 1111 628 1112
rect 622 1107 623 1111
rect 627 1107 628 1111
rect 622 1106 628 1107
rect 758 1111 764 1112
rect 758 1107 759 1111
rect 763 1107 764 1111
rect 758 1106 764 1107
rect 886 1111 892 1112
rect 886 1107 887 1111
rect 891 1107 892 1111
rect 886 1106 892 1107
rect 1014 1111 1020 1112
rect 1014 1107 1015 1111
rect 1019 1107 1020 1111
rect 1014 1106 1020 1107
rect 1142 1111 1148 1112
rect 1142 1107 1143 1111
rect 1147 1107 1148 1111
rect 1142 1106 1148 1107
rect 1270 1111 1276 1112
rect 1270 1107 1271 1111
rect 1275 1107 1276 1111
rect 1270 1106 1276 1107
rect 1398 1111 1404 1112
rect 1398 1107 1399 1111
rect 1403 1107 1404 1111
rect 1766 1108 1767 1112
rect 1771 1108 1772 1112
rect 1766 1107 1772 1108
rect 1806 1108 1812 1109
rect 3462 1108 3468 1109
rect 1398 1106 1404 1107
rect 1806 1104 1807 1108
rect 1811 1104 1812 1108
rect 318 1103 324 1104
rect 318 1099 319 1103
rect 323 1099 324 1103
rect 318 1098 324 1099
rect 438 1103 444 1104
rect 438 1099 439 1103
rect 443 1099 444 1103
rect 438 1098 444 1099
rect 566 1103 572 1104
rect 566 1099 567 1103
rect 571 1099 572 1103
rect 566 1098 572 1099
rect 694 1103 700 1104
rect 694 1099 695 1103
rect 699 1099 700 1103
rect 694 1098 700 1099
rect 702 1103 708 1104
rect 702 1099 703 1103
rect 707 1102 708 1103
rect 838 1103 844 1104
rect 707 1100 801 1102
rect 707 1099 708 1100
rect 702 1098 708 1099
rect 838 1099 839 1103
rect 843 1102 844 1103
rect 998 1103 1004 1104
rect 843 1100 929 1102
rect 843 1099 844 1100
rect 838 1098 844 1099
rect 998 1099 999 1103
rect 1003 1102 1004 1103
rect 1110 1103 1116 1104
rect 1003 1100 1057 1102
rect 1003 1099 1004 1100
rect 998 1098 1004 1099
rect 1110 1099 1111 1103
rect 1115 1102 1116 1103
rect 1222 1103 1228 1104
rect 1115 1100 1185 1102
rect 1115 1099 1116 1100
rect 1110 1098 1116 1099
rect 1222 1099 1223 1103
rect 1227 1102 1228 1103
rect 1350 1103 1356 1104
rect 1806 1103 1812 1104
rect 1942 1107 1948 1108
rect 1942 1103 1943 1107
rect 1947 1103 1948 1107
rect 1227 1100 1313 1102
rect 1227 1099 1228 1100
rect 1222 1098 1228 1099
rect 1350 1099 1351 1103
rect 1355 1102 1356 1103
rect 1942 1102 1948 1103
rect 2062 1107 2068 1108
rect 2062 1103 2063 1107
rect 2067 1103 2068 1107
rect 2062 1102 2068 1103
rect 2190 1107 2196 1108
rect 2190 1103 2191 1107
rect 2195 1103 2196 1107
rect 2190 1102 2196 1103
rect 2318 1107 2324 1108
rect 2318 1103 2319 1107
rect 2323 1103 2324 1107
rect 2318 1102 2324 1103
rect 2454 1107 2460 1108
rect 2454 1103 2455 1107
rect 2459 1103 2460 1107
rect 2454 1102 2460 1103
rect 2598 1107 2604 1108
rect 2598 1103 2599 1107
rect 2603 1103 2604 1107
rect 2598 1102 2604 1103
rect 2750 1107 2756 1108
rect 2750 1103 2751 1107
rect 2755 1103 2756 1107
rect 2750 1102 2756 1103
rect 2902 1107 2908 1108
rect 2902 1103 2903 1107
rect 2907 1103 2908 1107
rect 2902 1102 2908 1103
rect 3062 1107 3068 1108
rect 3062 1103 3063 1107
rect 3067 1103 3068 1107
rect 3062 1102 3068 1103
rect 3222 1107 3228 1108
rect 3222 1103 3223 1107
rect 3227 1103 3228 1107
rect 3222 1102 3228 1103
rect 3366 1107 3372 1108
rect 3366 1103 3367 1107
rect 3371 1103 3372 1107
rect 3462 1104 3463 1108
rect 3467 1104 3468 1108
rect 3462 1103 3468 1104
rect 3366 1102 3372 1103
rect 1355 1100 1441 1102
rect 1355 1099 1356 1100
rect 1350 1098 1356 1099
rect 2014 1099 2020 1100
rect 110 1095 116 1096
rect 110 1091 111 1095
rect 115 1091 116 1095
rect 1766 1095 1772 1096
rect 110 1090 116 1091
rect 246 1092 252 1093
rect 246 1088 247 1092
rect 251 1088 252 1092
rect 246 1087 252 1088
rect 366 1092 372 1093
rect 366 1088 367 1092
rect 371 1088 372 1092
rect 366 1087 372 1088
rect 494 1092 500 1093
rect 494 1088 495 1092
rect 499 1088 500 1092
rect 494 1087 500 1088
rect 622 1092 628 1093
rect 622 1088 623 1092
rect 627 1088 628 1092
rect 622 1087 628 1088
rect 758 1092 764 1093
rect 758 1088 759 1092
rect 763 1088 764 1092
rect 758 1087 764 1088
rect 886 1092 892 1093
rect 886 1088 887 1092
rect 891 1088 892 1092
rect 886 1087 892 1088
rect 1014 1092 1020 1093
rect 1014 1088 1015 1092
rect 1019 1088 1020 1092
rect 1014 1087 1020 1088
rect 1142 1092 1148 1093
rect 1142 1088 1143 1092
rect 1147 1088 1148 1092
rect 1142 1087 1148 1088
rect 1270 1092 1276 1093
rect 1270 1088 1271 1092
rect 1275 1088 1276 1092
rect 1270 1087 1276 1088
rect 1398 1092 1404 1093
rect 1398 1088 1399 1092
rect 1403 1088 1404 1092
rect 1766 1091 1767 1095
rect 1771 1091 1772 1095
rect 2014 1095 2015 1099
rect 2019 1095 2020 1099
rect 2014 1094 2020 1095
rect 2134 1099 2140 1100
rect 2134 1095 2135 1099
rect 2139 1095 2140 1099
rect 2134 1094 2140 1095
rect 2170 1099 2176 1100
rect 2170 1095 2171 1099
rect 2175 1098 2176 1099
rect 2390 1099 2396 1100
rect 2175 1096 2233 1098
rect 2175 1095 2176 1096
rect 2170 1094 2176 1095
rect 2390 1095 2391 1099
rect 2395 1095 2396 1099
rect 2390 1094 2396 1095
rect 2526 1099 2532 1100
rect 2526 1095 2527 1099
rect 2531 1095 2532 1099
rect 2526 1094 2532 1095
rect 2670 1099 2676 1100
rect 2670 1095 2671 1099
rect 2675 1095 2676 1099
rect 2830 1099 2836 1100
rect 2670 1094 2676 1095
rect 2822 1095 2828 1096
rect 1766 1090 1772 1091
rect 1806 1091 1812 1092
rect 1398 1087 1404 1088
rect 1806 1087 1807 1091
rect 1811 1087 1812 1091
rect 2822 1091 2823 1095
rect 2827 1091 2828 1095
rect 2830 1095 2831 1099
rect 2835 1098 2836 1099
rect 2982 1099 2988 1100
rect 2835 1096 2945 1098
rect 2835 1095 2836 1096
rect 2830 1094 2836 1095
rect 2982 1095 2983 1099
rect 2987 1098 2988 1099
rect 3294 1099 3300 1100
rect 2987 1096 3105 1098
rect 2987 1095 2988 1096
rect 2982 1094 2988 1095
rect 3294 1095 3295 1099
rect 3299 1095 3300 1099
rect 3294 1094 3300 1095
rect 3438 1095 3444 1096
rect 2822 1090 2828 1091
rect 3438 1091 3439 1095
rect 3443 1091 3444 1095
rect 3438 1090 3444 1091
rect 3462 1091 3468 1092
rect 1806 1086 1812 1087
rect 1942 1088 1948 1089
rect 1942 1084 1943 1088
rect 1947 1084 1948 1088
rect 1942 1083 1948 1084
rect 2062 1088 2068 1089
rect 2062 1084 2063 1088
rect 2067 1084 2068 1088
rect 2062 1083 2068 1084
rect 2190 1088 2196 1089
rect 2190 1084 2191 1088
rect 2195 1084 2196 1088
rect 2190 1083 2196 1084
rect 2318 1088 2324 1089
rect 2318 1084 2319 1088
rect 2323 1084 2324 1088
rect 2318 1083 2324 1084
rect 2454 1088 2460 1089
rect 2454 1084 2455 1088
rect 2459 1084 2460 1088
rect 2454 1083 2460 1084
rect 2598 1088 2604 1089
rect 2598 1084 2599 1088
rect 2603 1084 2604 1088
rect 2598 1083 2604 1084
rect 2750 1088 2756 1089
rect 2750 1084 2751 1088
rect 2755 1084 2756 1088
rect 2750 1083 2756 1084
rect 2902 1088 2908 1089
rect 2902 1084 2903 1088
rect 2907 1084 2908 1088
rect 2902 1083 2908 1084
rect 3062 1088 3068 1089
rect 3062 1084 3063 1088
rect 3067 1084 3068 1088
rect 3062 1083 3068 1084
rect 3222 1088 3228 1089
rect 3222 1084 3223 1088
rect 3227 1084 3228 1088
rect 3222 1083 3228 1084
rect 3366 1088 3372 1089
rect 3366 1084 3367 1088
rect 3371 1084 3372 1088
rect 3462 1087 3463 1091
rect 3467 1087 3468 1091
rect 3462 1086 3468 1087
rect 3366 1083 3372 1084
rect 482 1059 488 1060
rect 482 1055 483 1059
rect 487 1058 488 1059
rect 702 1059 708 1060
rect 702 1058 703 1059
rect 487 1056 703 1058
rect 487 1055 488 1056
rect 482 1054 488 1055
rect 702 1055 703 1056
rect 707 1055 708 1059
rect 702 1054 708 1055
rect 1090 1051 1096 1052
rect 1090 1047 1091 1051
rect 1095 1050 1096 1051
rect 1095 1048 1490 1050
rect 1095 1047 1096 1048
rect 1090 1046 1096 1047
rect 430 1044 436 1045
rect 110 1041 116 1042
rect 110 1037 111 1041
rect 115 1037 116 1041
rect 430 1040 431 1044
rect 435 1040 436 1044
rect 430 1039 436 1040
rect 542 1044 548 1045
rect 542 1040 543 1044
rect 547 1040 548 1044
rect 542 1039 548 1040
rect 662 1044 668 1045
rect 662 1040 663 1044
rect 667 1040 668 1044
rect 662 1039 668 1040
rect 790 1044 796 1045
rect 790 1040 791 1044
rect 795 1040 796 1044
rect 790 1039 796 1040
rect 918 1044 924 1045
rect 918 1040 919 1044
rect 923 1040 924 1044
rect 918 1039 924 1040
rect 1038 1044 1044 1045
rect 1038 1040 1039 1044
rect 1043 1040 1044 1044
rect 1038 1039 1044 1040
rect 1158 1044 1164 1045
rect 1158 1040 1159 1044
rect 1163 1040 1164 1044
rect 1158 1039 1164 1040
rect 1278 1044 1284 1045
rect 1278 1040 1279 1044
rect 1283 1040 1284 1044
rect 1278 1039 1284 1040
rect 1406 1044 1412 1045
rect 1406 1040 1407 1044
rect 1411 1040 1412 1044
rect 1406 1039 1412 1040
rect 110 1036 116 1037
rect 502 1035 508 1036
rect 502 1031 503 1035
rect 507 1031 508 1035
rect 502 1030 508 1031
rect 614 1035 620 1036
rect 614 1031 615 1035
rect 619 1031 620 1035
rect 614 1030 620 1031
rect 734 1035 740 1036
rect 734 1031 735 1035
rect 739 1031 740 1035
rect 734 1030 740 1031
rect 862 1035 868 1036
rect 862 1031 863 1035
rect 867 1031 868 1035
rect 862 1030 868 1031
rect 870 1035 876 1036
rect 870 1031 871 1035
rect 875 1034 876 1035
rect 1110 1035 1116 1036
rect 875 1032 961 1034
rect 875 1031 876 1032
rect 870 1030 876 1031
rect 1110 1031 1111 1035
rect 1115 1031 1116 1035
rect 1110 1030 1116 1031
rect 1230 1035 1236 1036
rect 1230 1031 1231 1035
rect 1235 1031 1236 1035
rect 1382 1035 1388 1036
rect 1382 1034 1383 1035
rect 1353 1032 1383 1034
rect 1230 1030 1236 1031
rect 1382 1031 1383 1032
rect 1387 1031 1388 1035
rect 1382 1030 1388 1031
rect 1478 1035 1484 1036
rect 1478 1031 1479 1035
rect 1483 1031 1484 1035
rect 1488 1034 1490 1048
rect 2594 1047 2600 1048
rect 1534 1044 1540 1045
rect 1534 1040 1535 1044
rect 1539 1040 1540 1044
rect 2594 1043 2595 1047
rect 2599 1046 2600 1047
rect 2599 1044 2962 1046
rect 2599 1043 2600 1044
rect 2594 1042 2600 1043
rect 1534 1039 1540 1040
rect 1766 1041 1772 1042
rect 1766 1037 1767 1041
rect 1771 1037 1772 1041
rect 1846 1040 1852 1041
rect 1766 1036 1772 1037
rect 1806 1037 1812 1038
rect 1488 1032 1577 1034
rect 1806 1033 1807 1037
rect 1811 1033 1812 1037
rect 1846 1036 1847 1040
rect 1851 1036 1852 1040
rect 1846 1035 1852 1036
rect 1982 1040 1988 1041
rect 1982 1036 1983 1040
rect 1987 1036 1988 1040
rect 1982 1035 1988 1036
rect 2118 1040 2124 1041
rect 2118 1036 2119 1040
rect 2123 1036 2124 1040
rect 2118 1035 2124 1036
rect 2254 1040 2260 1041
rect 2254 1036 2255 1040
rect 2259 1036 2260 1040
rect 2254 1035 2260 1036
rect 2390 1040 2396 1041
rect 2390 1036 2391 1040
rect 2395 1036 2396 1040
rect 2390 1035 2396 1036
rect 2542 1040 2548 1041
rect 2542 1036 2543 1040
rect 2547 1036 2548 1040
rect 2542 1035 2548 1036
rect 2702 1040 2708 1041
rect 2702 1036 2703 1040
rect 2707 1036 2708 1040
rect 2702 1035 2708 1036
rect 2862 1040 2868 1041
rect 2862 1036 2863 1040
rect 2867 1036 2868 1040
rect 2862 1035 2868 1036
rect 1806 1032 1812 1033
rect 1478 1030 1484 1031
rect 1926 1031 1932 1032
rect 1926 1027 1927 1031
rect 1931 1030 1932 1031
rect 2062 1031 2068 1032
rect 1931 1028 2025 1030
rect 1931 1027 1932 1028
rect 1926 1026 1932 1027
rect 2062 1027 2063 1031
rect 2067 1030 2068 1031
rect 2370 1031 2376 1032
rect 2067 1028 2161 1030
rect 2067 1027 2068 1028
rect 2062 1026 2068 1027
rect 2370 1027 2371 1031
rect 2375 1030 2376 1031
rect 2614 1031 2620 1032
rect 2375 1028 2433 1030
rect 2375 1027 2376 1028
rect 2370 1026 2376 1027
rect 2614 1027 2615 1031
rect 2619 1027 2620 1031
rect 2614 1026 2620 1027
rect 2774 1031 2780 1032
rect 2774 1027 2775 1031
rect 2779 1027 2780 1031
rect 2774 1026 2780 1027
rect 2934 1031 2940 1032
rect 2934 1027 2935 1031
rect 2939 1027 2940 1031
rect 2960 1030 2962 1044
rect 3030 1040 3036 1041
rect 3030 1036 3031 1040
rect 3035 1036 3036 1040
rect 3030 1035 3036 1036
rect 3206 1040 3212 1041
rect 3206 1036 3207 1040
rect 3211 1036 3212 1040
rect 3206 1035 3212 1036
rect 3366 1040 3372 1041
rect 3366 1036 3367 1040
rect 3371 1036 3372 1040
rect 3366 1035 3372 1036
rect 3462 1037 3468 1038
rect 3462 1033 3463 1037
rect 3467 1033 3468 1037
rect 3462 1032 3468 1033
rect 3270 1031 3276 1032
rect 2960 1028 3073 1030
rect 2934 1026 2940 1027
rect 3270 1027 3271 1031
rect 3275 1027 3276 1031
rect 3270 1026 3276 1027
rect 3430 1031 3436 1032
rect 3430 1027 3431 1031
rect 3435 1027 3436 1031
rect 3430 1026 3436 1027
rect 430 1025 436 1026
rect 110 1024 116 1025
rect 110 1020 111 1024
rect 115 1020 116 1024
rect 430 1021 431 1025
rect 435 1021 436 1025
rect 430 1020 436 1021
rect 542 1025 548 1026
rect 542 1021 543 1025
rect 547 1021 548 1025
rect 542 1020 548 1021
rect 662 1025 668 1026
rect 662 1021 663 1025
rect 667 1021 668 1025
rect 662 1020 668 1021
rect 790 1025 796 1026
rect 790 1021 791 1025
rect 795 1021 796 1025
rect 790 1020 796 1021
rect 918 1025 924 1026
rect 918 1021 919 1025
rect 923 1021 924 1025
rect 918 1020 924 1021
rect 1038 1025 1044 1026
rect 1038 1021 1039 1025
rect 1043 1021 1044 1025
rect 1038 1020 1044 1021
rect 1158 1025 1164 1026
rect 1158 1021 1159 1025
rect 1163 1021 1164 1025
rect 1158 1020 1164 1021
rect 1278 1025 1284 1026
rect 1278 1021 1279 1025
rect 1283 1021 1284 1025
rect 1278 1020 1284 1021
rect 1406 1025 1412 1026
rect 1406 1021 1407 1025
rect 1411 1021 1412 1025
rect 1406 1020 1412 1021
rect 1534 1025 1540 1026
rect 1534 1021 1535 1025
rect 1539 1021 1540 1025
rect 1534 1020 1540 1021
rect 1766 1024 1772 1025
rect 1766 1020 1767 1024
rect 1771 1020 1772 1024
rect 1919 1023 1925 1024
rect 1846 1021 1852 1022
rect 110 1019 116 1020
rect 1766 1019 1772 1020
rect 1806 1020 1812 1021
rect 1806 1016 1807 1020
rect 1811 1016 1812 1020
rect 1846 1017 1847 1021
rect 1851 1017 1852 1021
rect 1919 1019 1920 1023
rect 1924 1022 1925 1023
rect 1951 1023 1957 1024
rect 1951 1022 1952 1023
rect 1924 1020 1952 1022
rect 1924 1019 1925 1020
rect 1919 1018 1925 1019
rect 1951 1019 1952 1020
rect 1956 1019 1957 1023
rect 2327 1023 2333 1024
rect 1951 1018 1957 1019
rect 1982 1021 1988 1022
rect 1846 1016 1852 1017
rect 1982 1017 1983 1021
rect 1987 1017 1988 1021
rect 1982 1016 1988 1017
rect 2118 1021 2124 1022
rect 2118 1017 2119 1021
rect 2123 1017 2124 1021
rect 2118 1016 2124 1017
rect 2254 1021 2260 1022
rect 2254 1017 2255 1021
rect 2259 1017 2260 1021
rect 2327 1019 2328 1023
rect 2332 1022 2333 1023
rect 2375 1023 2381 1024
rect 2375 1022 2376 1023
rect 2332 1020 2376 1022
rect 2332 1019 2333 1020
rect 2327 1018 2333 1019
rect 2375 1019 2376 1020
rect 2380 1019 2381 1023
rect 2375 1018 2381 1019
rect 2390 1021 2396 1022
rect 2254 1016 2260 1017
rect 2390 1017 2391 1021
rect 2395 1017 2396 1021
rect 2390 1016 2396 1017
rect 2542 1021 2548 1022
rect 2542 1017 2543 1021
rect 2547 1017 2548 1021
rect 2542 1016 2548 1017
rect 2702 1021 2708 1022
rect 2702 1017 2703 1021
rect 2707 1017 2708 1021
rect 2702 1016 2708 1017
rect 2862 1021 2868 1022
rect 2862 1017 2863 1021
rect 2867 1017 2868 1021
rect 2862 1016 2868 1017
rect 3030 1021 3036 1022
rect 3030 1017 3031 1021
rect 3035 1017 3036 1021
rect 3030 1016 3036 1017
rect 3206 1021 3212 1022
rect 3206 1017 3207 1021
rect 3211 1017 3212 1021
rect 3206 1016 3212 1017
rect 3366 1021 3372 1022
rect 3366 1017 3367 1021
rect 3371 1017 3372 1021
rect 3366 1016 3372 1017
rect 3462 1020 3468 1021
rect 3462 1016 3463 1020
rect 3467 1016 3468 1020
rect 1806 1015 1812 1016
rect 3462 1015 3468 1016
rect 479 1007 488 1008
rect 479 1003 480 1007
rect 487 1003 488 1007
rect 479 1002 488 1003
rect 502 1007 508 1008
rect 502 1003 503 1007
rect 507 1006 508 1007
rect 591 1007 597 1008
rect 591 1006 592 1007
rect 507 1004 592 1006
rect 507 1003 508 1004
rect 502 1002 508 1003
rect 591 1003 592 1004
rect 596 1003 597 1007
rect 591 1002 597 1003
rect 614 1007 620 1008
rect 614 1003 615 1007
rect 619 1006 620 1007
rect 711 1007 717 1008
rect 711 1006 712 1007
rect 619 1004 712 1006
rect 619 1003 620 1004
rect 614 1002 620 1003
rect 711 1003 712 1004
rect 716 1003 717 1007
rect 711 1002 717 1003
rect 734 1007 740 1008
rect 734 1003 735 1007
rect 739 1006 740 1007
rect 839 1007 845 1008
rect 839 1006 840 1007
rect 739 1004 840 1006
rect 739 1003 740 1004
rect 734 1002 740 1003
rect 839 1003 840 1004
rect 844 1003 845 1007
rect 839 1002 845 1003
rect 862 1007 868 1008
rect 862 1003 863 1007
rect 867 1006 868 1007
rect 967 1007 973 1008
rect 967 1006 968 1007
rect 867 1004 968 1006
rect 867 1003 868 1004
rect 862 1002 868 1003
rect 967 1003 968 1004
rect 972 1003 973 1007
rect 967 1002 973 1003
rect 1087 1007 1096 1008
rect 1087 1003 1088 1007
rect 1095 1003 1096 1007
rect 1087 1002 1096 1003
rect 1110 1007 1116 1008
rect 1110 1003 1111 1007
rect 1115 1006 1116 1007
rect 1207 1007 1213 1008
rect 1207 1006 1208 1007
rect 1115 1004 1208 1006
rect 1115 1003 1116 1004
rect 1110 1002 1116 1003
rect 1207 1003 1208 1004
rect 1212 1003 1213 1007
rect 1207 1002 1213 1003
rect 1230 1007 1236 1008
rect 1230 1003 1231 1007
rect 1235 1006 1236 1007
rect 1327 1007 1333 1008
rect 1327 1006 1328 1007
rect 1235 1004 1328 1006
rect 1235 1003 1236 1004
rect 1230 1002 1236 1003
rect 1327 1003 1328 1004
rect 1332 1003 1333 1007
rect 1327 1002 1333 1003
rect 1430 1007 1436 1008
rect 1430 1003 1431 1007
rect 1435 1006 1436 1007
rect 1455 1007 1461 1008
rect 1455 1006 1456 1007
rect 1435 1004 1456 1006
rect 1435 1003 1436 1004
rect 1430 1002 1436 1003
rect 1455 1003 1456 1004
rect 1460 1003 1461 1007
rect 1455 1002 1461 1003
rect 1478 1007 1484 1008
rect 1478 1003 1479 1007
rect 1483 1006 1484 1007
rect 1583 1007 1589 1008
rect 1583 1006 1584 1007
rect 1483 1004 1584 1006
rect 1483 1003 1484 1004
rect 1478 1002 1484 1003
rect 1583 1003 1584 1004
rect 1588 1003 1589 1007
rect 1583 1002 1589 1003
rect 1895 1003 1901 1004
rect 1895 999 1896 1003
rect 1900 1002 1901 1003
rect 1926 1003 1932 1004
rect 1926 1002 1927 1003
rect 1900 1000 1927 1002
rect 1900 999 1901 1000
rect 1895 998 1901 999
rect 1926 999 1927 1000
rect 1931 999 1932 1003
rect 1926 998 1932 999
rect 2031 1003 2037 1004
rect 2031 999 2032 1003
rect 2036 1002 2037 1003
rect 2062 1003 2068 1004
rect 2062 1002 2063 1003
rect 2036 1000 2063 1002
rect 2036 999 2037 1000
rect 2031 998 2037 999
rect 2062 999 2063 1000
rect 2067 999 2068 1003
rect 2062 998 2068 999
rect 2167 1003 2176 1004
rect 2167 999 2168 1003
rect 2175 999 2176 1003
rect 2167 998 2176 999
rect 2303 1003 2309 1004
rect 2303 999 2304 1003
rect 2308 1002 2309 1003
rect 2366 1003 2372 1004
rect 2366 1002 2367 1003
rect 2308 1000 2367 1002
rect 2308 999 2309 1000
rect 2303 998 2309 999
rect 2366 999 2367 1000
rect 2371 999 2372 1003
rect 2366 998 2372 999
rect 2375 1003 2381 1004
rect 2375 999 2376 1003
rect 2380 1002 2381 1003
rect 2439 1003 2445 1004
rect 2439 1002 2440 1003
rect 2380 1000 2440 1002
rect 2380 999 2381 1000
rect 2375 998 2381 999
rect 2439 999 2440 1000
rect 2444 999 2445 1003
rect 2439 998 2445 999
rect 2591 1003 2600 1004
rect 2591 999 2592 1003
rect 2599 999 2600 1003
rect 2591 998 2600 999
rect 2614 1003 2620 1004
rect 2614 999 2615 1003
rect 2619 1002 2620 1003
rect 2751 1003 2757 1004
rect 2751 1002 2752 1003
rect 2619 1000 2752 1002
rect 2619 999 2620 1000
rect 2614 998 2620 999
rect 2751 999 2752 1000
rect 2756 999 2757 1003
rect 2751 998 2757 999
rect 2822 1003 2828 1004
rect 2822 999 2823 1003
rect 2827 1002 2828 1003
rect 2911 1003 2917 1004
rect 2911 1002 2912 1003
rect 2827 1000 2912 1002
rect 2827 999 2828 1000
rect 2822 998 2828 999
rect 2911 999 2912 1000
rect 2916 999 2917 1003
rect 2911 998 2917 999
rect 2934 1003 2940 1004
rect 2934 999 2935 1003
rect 2939 1002 2940 1003
rect 3079 1003 3085 1004
rect 3079 1002 3080 1003
rect 2939 1000 3080 1002
rect 2939 999 2940 1000
rect 2934 998 2940 999
rect 3079 999 3080 1000
rect 3084 999 3085 1003
rect 3079 998 3085 999
rect 3254 1003 3261 1004
rect 3254 999 3255 1003
rect 3260 999 3261 1003
rect 3254 998 3261 999
rect 3415 1003 3421 1004
rect 3415 999 3416 1003
rect 3420 1002 3421 1003
rect 3438 1003 3444 1004
rect 3438 1002 3439 1003
rect 3420 1000 3439 1002
rect 3420 999 3421 1000
rect 3415 998 3421 999
rect 3438 999 3439 1000
rect 3443 999 3444 1003
rect 3438 998 3444 999
rect 870 995 876 996
rect 870 994 871 995
rect 632 992 871 994
rect 615 987 621 988
rect 615 983 616 987
rect 620 986 621 987
rect 632 986 634 992
rect 870 991 871 992
rect 875 991 876 995
rect 1438 995 1444 996
rect 1438 994 1439 995
rect 870 990 876 991
rect 1208 992 1439 994
rect 620 984 634 986
rect 638 987 644 988
rect 620 983 621 984
rect 615 982 621 983
rect 638 983 639 987
rect 643 986 644 987
rect 727 987 733 988
rect 727 986 728 987
rect 643 984 728 986
rect 643 983 644 984
rect 638 982 644 983
rect 727 983 728 984
rect 732 983 733 987
rect 727 982 733 983
rect 750 987 756 988
rect 750 983 751 987
rect 755 986 756 987
rect 839 987 845 988
rect 839 986 840 987
rect 755 984 840 986
rect 755 983 756 984
rect 750 982 756 983
rect 839 983 840 984
rect 844 983 845 987
rect 839 982 845 983
rect 862 987 868 988
rect 862 983 863 987
rect 867 986 868 987
rect 959 987 965 988
rect 959 986 960 987
rect 867 984 960 986
rect 867 983 868 984
rect 862 982 868 983
rect 959 983 960 984
rect 964 983 965 987
rect 959 982 965 983
rect 982 987 988 988
rect 982 983 983 987
rect 987 986 988 987
rect 1079 987 1085 988
rect 1079 986 1080 987
rect 987 984 1080 986
rect 987 983 988 984
rect 982 982 988 983
rect 1079 983 1080 984
rect 1084 983 1085 987
rect 1079 982 1085 983
rect 1191 987 1197 988
rect 1191 983 1192 987
rect 1196 986 1197 987
rect 1208 986 1210 992
rect 1438 991 1439 992
rect 1443 991 1444 995
rect 2418 995 2424 996
rect 2418 994 2419 995
rect 1438 990 1444 991
rect 2336 992 2419 994
rect 1196 984 1210 986
rect 1214 987 1220 988
rect 1196 983 1197 984
rect 1191 982 1197 983
rect 1214 983 1215 987
rect 1219 986 1220 987
rect 1303 987 1309 988
rect 1303 986 1304 987
rect 1219 984 1304 986
rect 1219 983 1220 984
rect 1214 982 1220 983
rect 1303 983 1304 984
rect 1308 983 1309 987
rect 1303 982 1309 983
rect 1326 987 1332 988
rect 1326 983 1327 987
rect 1331 986 1332 987
rect 1407 987 1413 988
rect 1407 986 1408 987
rect 1331 984 1408 986
rect 1331 983 1332 984
rect 1326 982 1332 983
rect 1407 983 1408 984
rect 1412 983 1413 987
rect 1407 982 1413 983
rect 1519 987 1528 988
rect 1519 983 1520 987
rect 1527 983 1528 987
rect 1519 982 1528 983
rect 1631 987 1637 988
rect 1631 983 1632 987
rect 1636 986 1637 987
rect 1662 987 1668 988
rect 1662 986 1663 987
rect 1636 984 1663 986
rect 1636 983 1637 984
rect 1631 982 1637 983
rect 1662 983 1663 984
rect 1667 983 1668 987
rect 1662 982 1668 983
rect 1719 987 1725 988
rect 1719 983 1720 987
rect 1724 986 1725 987
rect 1750 987 1756 988
rect 1750 986 1751 987
rect 1724 984 1751 986
rect 1724 983 1725 984
rect 1719 982 1725 983
rect 1750 983 1751 984
rect 1755 983 1756 987
rect 1750 982 1756 983
rect 1879 987 1885 988
rect 1879 983 1880 987
rect 1884 986 1885 987
rect 1938 987 1944 988
rect 1938 986 1939 987
rect 1884 984 1939 986
rect 1884 983 1885 984
rect 1879 982 1885 983
rect 1938 983 1939 984
rect 1943 983 1944 987
rect 1938 982 1944 983
rect 1951 987 1957 988
rect 1951 983 1952 987
rect 1956 986 1957 987
rect 2023 987 2029 988
rect 2023 986 2024 987
rect 1956 984 2024 986
rect 1956 983 1957 984
rect 1951 982 1957 983
rect 2023 983 2024 984
rect 2028 983 2029 987
rect 2023 982 2029 983
rect 2183 987 2189 988
rect 2183 983 2184 987
rect 2188 986 2189 987
rect 2336 986 2338 992
rect 2418 991 2419 992
rect 2423 991 2424 995
rect 2958 995 2964 996
rect 2958 994 2959 995
rect 2418 990 2424 991
rect 2839 992 2959 994
rect 2839 990 2841 992
rect 2958 991 2959 992
rect 2963 991 2964 995
rect 2958 990 2964 991
rect 2696 988 2841 990
rect 2188 984 2338 986
rect 2343 987 2349 988
rect 2188 983 2189 984
rect 2183 982 2189 983
rect 2343 983 2344 987
rect 2348 986 2349 987
rect 2470 987 2476 988
rect 2470 986 2471 987
rect 2348 984 2471 986
rect 2348 983 2349 984
rect 2343 982 2349 983
rect 2470 983 2471 984
rect 2475 983 2476 987
rect 2470 982 2476 983
rect 2511 987 2517 988
rect 2511 983 2512 987
rect 2516 986 2517 987
rect 2543 987 2549 988
rect 2543 986 2544 987
rect 2516 984 2544 986
rect 2516 983 2517 984
rect 2511 982 2517 983
rect 2543 983 2544 984
rect 2548 983 2549 987
rect 2543 982 2549 983
rect 2679 987 2685 988
rect 2679 983 2680 987
rect 2684 986 2685 987
rect 2696 986 2698 988
rect 2855 987 2861 988
rect 2855 986 2856 987
rect 2684 984 2698 986
rect 2839 984 2856 986
rect 2684 983 2685 984
rect 2679 982 2685 983
rect 2774 983 2780 984
rect 2774 979 2775 983
rect 2779 982 2780 983
rect 2839 982 2841 984
rect 2855 983 2856 984
rect 2860 983 2861 987
rect 2855 982 2861 983
rect 2878 987 2884 988
rect 2878 983 2879 987
rect 2883 986 2884 987
rect 3039 987 3045 988
rect 3039 986 3040 987
rect 2883 984 3040 986
rect 2883 983 2884 984
rect 2878 982 2884 983
rect 3039 983 3040 984
rect 3044 983 3045 987
rect 3039 982 3045 983
rect 3231 987 3237 988
rect 3231 983 3232 987
rect 3236 986 3237 987
rect 3294 987 3300 988
rect 3294 986 3295 987
rect 3236 984 3295 986
rect 3236 983 3237 984
rect 3231 982 3237 983
rect 3294 983 3295 984
rect 3299 983 3300 987
rect 3294 982 3300 983
rect 3415 987 3421 988
rect 3415 983 3416 987
rect 3420 986 3421 987
rect 3430 987 3436 988
rect 3430 986 3431 987
rect 3420 984 3431 986
rect 3420 983 3421 984
rect 3415 982 3421 983
rect 3430 983 3431 984
rect 3435 983 3436 987
rect 3430 982 3436 983
rect 2779 980 2841 982
rect 2779 979 2780 980
rect 2774 978 2780 979
rect 110 972 116 973
rect 1766 972 1772 973
rect 110 968 111 972
rect 115 968 116 972
rect 110 967 116 968
rect 566 971 572 972
rect 566 967 567 971
rect 571 967 572 971
rect 566 966 572 967
rect 678 971 684 972
rect 678 967 679 971
rect 683 967 684 971
rect 678 966 684 967
rect 790 971 796 972
rect 790 967 791 971
rect 795 967 796 971
rect 790 966 796 967
rect 910 971 916 972
rect 910 967 911 971
rect 915 967 916 971
rect 910 966 916 967
rect 1030 971 1036 972
rect 1030 967 1031 971
rect 1035 967 1036 971
rect 1030 966 1036 967
rect 1142 971 1148 972
rect 1142 967 1143 971
rect 1147 967 1148 971
rect 1142 966 1148 967
rect 1254 971 1260 972
rect 1254 967 1255 971
rect 1259 967 1260 971
rect 1254 966 1260 967
rect 1358 971 1364 972
rect 1358 967 1359 971
rect 1363 967 1364 971
rect 1358 966 1364 967
rect 1470 971 1476 972
rect 1470 967 1471 971
rect 1475 967 1476 971
rect 1470 966 1476 967
rect 1582 971 1588 972
rect 1582 967 1583 971
rect 1587 967 1588 971
rect 1582 966 1588 967
rect 1670 971 1676 972
rect 1670 967 1671 971
rect 1675 967 1676 971
rect 1766 968 1767 972
rect 1771 968 1772 972
rect 1766 967 1772 968
rect 1806 972 1812 973
rect 3462 972 3468 973
rect 1806 968 1807 972
rect 1811 968 1812 972
rect 1806 967 1812 968
rect 1830 971 1836 972
rect 1830 967 1831 971
rect 1835 967 1836 971
rect 1670 966 1676 967
rect 1830 966 1836 967
rect 1974 971 1980 972
rect 1974 967 1975 971
rect 1979 967 1980 971
rect 1974 966 1980 967
rect 2134 971 2140 972
rect 2134 967 2135 971
rect 2139 967 2140 971
rect 2134 966 2140 967
rect 2294 971 2300 972
rect 2294 967 2295 971
rect 2299 967 2300 971
rect 2294 966 2300 967
rect 2462 971 2468 972
rect 2462 967 2463 971
rect 2467 967 2468 971
rect 2462 966 2468 967
rect 2630 971 2636 972
rect 2630 967 2631 971
rect 2635 967 2636 971
rect 2630 966 2636 967
rect 2806 971 2812 972
rect 2806 967 2807 971
rect 2811 967 2812 971
rect 2806 966 2812 967
rect 2990 971 2996 972
rect 2990 967 2991 971
rect 2995 967 2996 971
rect 2990 966 2996 967
rect 3182 971 3188 972
rect 3182 967 3183 971
rect 3187 967 3188 971
rect 3182 966 3188 967
rect 3366 971 3372 972
rect 3366 967 3367 971
rect 3371 967 3372 971
rect 3462 968 3463 972
rect 3467 968 3468 972
rect 3462 967 3468 968
rect 3366 966 3372 967
rect 638 963 644 964
rect 638 959 639 963
rect 643 959 644 963
rect 638 958 644 959
rect 750 963 756 964
rect 750 959 751 963
rect 755 959 756 963
rect 750 958 756 959
rect 862 963 868 964
rect 862 959 863 963
rect 867 959 868 963
rect 862 958 868 959
rect 982 963 988 964
rect 982 959 983 963
rect 987 959 988 963
rect 982 958 988 959
rect 990 963 996 964
rect 990 959 991 963
rect 995 962 996 963
rect 1214 963 1220 964
rect 995 960 1073 962
rect 995 959 996 960
rect 990 958 996 959
rect 1214 959 1215 963
rect 1219 959 1220 963
rect 1214 958 1220 959
rect 1326 963 1332 964
rect 1326 959 1327 963
rect 1331 959 1332 963
rect 1326 958 1332 959
rect 1430 963 1436 964
rect 1430 959 1431 963
rect 1435 959 1436 963
rect 1430 958 1436 959
rect 1438 963 1444 964
rect 1438 959 1439 963
rect 1443 962 1444 963
rect 1662 963 1668 964
rect 1443 960 1513 962
rect 1443 959 1444 960
rect 1438 958 1444 959
rect 1654 959 1660 960
rect 110 955 116 956
rect 110 951 111 955
rect 115 951 116 955
rect 1654 955 1655 959
rect 1659 955 1660 959
rect 1662 959 1663 963
rect 1667 962 1668 963
rect 1750 963 1756 964
rect 1667 960 1713 962
rect 1667 959 1668 960
rect 1662 958 1668 959
rect 1750 959 1751 963
rect 1755 962 1756 963
rect 1938 963 1944 964
rect 1755 960 1873 962
rect 1755 959 1756 960
rect 1750 958 1756 959
rect 1938 959 1939 963
rect 1943 962 1944 963
rect 2366 963 2372 964
rect 1943 960 2017 962
rect 1943 959 1944 960
rect 1938 958 1944 959
rect 2206 959 2212 960
rect 1654 954 1660 955
rect 1766 955 1772 956
rect 110 950 116 951
rect 566 952 572 953
rect 566 948 567 952
rect 571 948 572 952
rect 566 947 572 948
rect 678 952 684 953
rect 678 948 679 952
rect 683 948 684 952
rect 678 947 684 948
rect 790 952 796 953
rect 790 948 791 952
rect 795 948 796 952
rect 790 947 796 948
rect 910 952 916 953
rect 910 948 911 952
rect 915 948 916 952
rect 910 947 916 948
rect 1030 952 1036 953
rect 1030 948 1031 952
rect 1035 948 1036 952
rect 1030 947 1036 948
rect 1142 952 1148 953
rect 1142 948 1143 952
rect 1147 948 1148 952
rect 1142 947 1148 948
rect 1254 952 1260 953
rect 1254 948 1255 952
rect 1259 948 1260 952
rect 1254 947 1260 948
rect 1358 952 1364 953
rect 1358 948 1359 952
rect 1363 948 1364 952
rect 1358 947 1364 948
rect 1470 952 1476 953
rect 1470 948 1471 952
rect 1475 948 1476 952
rect 1470 947 1476 948
rect 1582 952 1588 953
rect 1582 948 1583 952
rect 1587 948 1588 952
rect 1582 947 1588 948
rect 1670 952 1676 953
rect 1670 948 1671 952
rect 1675 948 1676 952
rect 1766 951 1767 955
rect 1771 951 1772 955
rect 1766 950 1772 951
rect 1806 955 1812 956
rect 1806 951 1807 955
rect 1811 951 1812 955
rect 2206 955 2207 959
rect 2211 955 2212 959
rect 2366 959 2367 963
rect 2371 959 2372 963
rect 2366 958 2372 959
rect 2418 963 2424 964
rect 2418 959 2419 963
rect 2423 962 2424 963
rect 2543 963 2549 964
rect 2423 960 2505 962
rect 2423 959 2424 960
rect 2418 958 2424 959
rect 2543 959 2544 963
rect 2548 962 2549 963
rect 2878 963 2884 964
rect 2548 960 2673 962
rect 2548 959 2549 960
rect 2543 958 2549 959
rect 2878 959 2879 963
rect 2883 959 2884 963
rect 2878 958 2884 959
rect 2958 963 2964 964
rect 2958 959 2959 963
rect 2963 962 2964 963
rect 3254 963 3260 964
rect 2963 960 3033 962
rect 2963 959 2964 960
rect 2958 958 2964 959
rect 3254 959 3255 963
rect 3259 959 3260 963
rect 3254 958 3260 959
rect 3438 959 3444 960
rect 2206 954 2212 955
rect 3438 955 3439 959
rect 3443 955 3444 959
rect 3438 954 3444 955
rect 3462 955 3468 956
rect 1806 950 1812 951
rect 1830 952 1836 953
rect 1670 947 1676 948
rect 1830 948 1831 952
rect 1835 948 1836 952
rect 1830 947 1836 948
rect 1974 952 1980 953
rect 1974 948 1975 952
rect 1979 948 1980 952
rect 1974 947 1980 948
rect 2134 952 2140 953
rect 2134 948 2135 952
rect 2139 948 2140 952
rect 2134 947 2140 948
rect 2294 952 2300 953
rect 2294 948 2295 952
rect 2299 948 2300 952
rect 2294 947 2300 948
rect 2462 952 2468 953
rect 2462 948 2463 952
rect 2467 948 2468 952
rect 2462 947 2468 948
rect 2630 952 2636 953
rect 2630 948 2631 952
rect 2635 948 2636 952
rect 2630 947 2636 948
rect 2806 952 2812 953
rect 2806 948 2807 952
rect 2811 948 2812 952
rect 2806 947 2812 948
rect 2990 952 2996 953
rect 2990 948 2991 952
rect 2995 948 2996 952
rect 2990 947 2996 948
rect 3182 952 3188 953
rect 3182 948 3183 952
rect 3187 948 3188 952
rect 3182 947 3188 948
rect 3366 952 3372 953
rect 3366 948 3367 952
rect 3371 948 3372 952
rect 3462 951 3463 955
rect 3467 951 3468 955
rect 3462 950 3468 951
rect 3366 947 3372 948
rect 2126 908 2132 909
rect 1806 905 1812 906
rect 414 904 420 905
rect 110 901 116 902
rect 110 897 111 901
rect 115 897 116 901
rect 414 900 415 904
rect 419 900 420 904
rect 414 899 420 900
rect 558 904 564 905
rect 558 900 559 904
rect 563 900 564 904
rect 558 899 564 900
rect 726 904 732 905
rect 726 900 727 904
rect 731 900 732 904
rect 726 899 732 900
rect 910 904 916 905
rect 910 900 911 904
rect 915 900 916 904
rect 910 899 916 900
rect 1118 904 1124 905
rect 1118 900 1119 904
rect 1123 900 1124 904
rect 1118 899 1124 900
rect 1334 904 1340 905
rect 1334 900 1335 904
rect 1339 900 1340 904
rect 1334 899 1340 900
rect 1558 904 1564 905
rect 1558 900 1559 904
rect 1563 900 1564 904
rect 1558 899 1564 900
rect 1766 901 1772 902
rect 110 896 116 897
rect 1766 897 1767 901
rect 1771 897 1772 901
rect 1806 901 1807 905
rect 1811 901 1812 905
rect 2126 904 2127 908
rect 2131 904 2132 908
rect 2126 903 2132 904
rect 2214 908 2220 909
rect 2214 904 2215 908
rect 2219 904 2220 908
rect 2214 903 2220 904
rect 2302 908 2308 909
rect 2302 904 2303 908
rect 2307 904 2308 908
rect 2302 903 2308 904
rect 2390 908 2396 909
rect 2390 904 2391 908
rect 2395 904 2396 908
rect 2390 903 2396 904
rect 2478 908 2484 909
rect 2478 904 2479 908
rect 2483 904 2484 908
rect 2478 903 2484 904
rect 2566 908 2572 909
rect 2566 904 2567 908
rect 2571 904 2572 908
rect 2566 903 2572 904
rect 2654 908 2660 909
rect 2654 904 2655 908
rect 2659 904 2660 908
rect 2654 903 2660 904
rect 2742 908 2748 909
rect 2742 904 2743 908
rect 2747 904 2748 908
rect 2742 903 2748 904
rect 2830 908 2836 909
rect 2830 904 2831 908
rect 2835 904 2836 908
rect 2830 903 2836 904
rect 3462 905 3468 906
rect 1806 900 1812 901
rect 3462 901 3463 905
rect 3467 901 3468 905
rect 3462 900 3468 901
rect 1766 896 1772 897
rect 2286 899 2292 900
rect 486 895 492 896
rect 486 891 487 895
rect 491 891 492 895
rect 486 890 492 891
rect 630 895 636 896
rect 630 891 631 895
rect 635 891 636 895
rect 630 890 636 891
rect 678 895 684 896
rect 678 891 679 895
rect 683 894 684 895
rect 806 895 812 896
rect 683 892 769 894
rect 683 891 684 892
rect 678 890 684 891
rect 806 891 807 895
rect 811 894 812 895
rect 1190 895 1196 896
rect 811 892 953 894
rect 811 891 812 892
rect 806 890 812 891
rect 1190 891 1191 895
rect 1195 891 1196 895
rect 1190 890 1196 891
rect 1322 895 1328 896
rect 1322 891 1323 895
rect 1327 894 1328 895
rect 1522 895 1528 896
rect 1327 892 1377 894
rect 1327 891 1328 892
rect 1322 890 1328 891
rect 1522 891 1523 895
rect 1527 894 1528 895
rect 2286 895 2287 899
rect 2291 895 2292 899
rect 2286 894 2292 895
rect 2374 899 2380 900
rect 2374 895 2375 899
rect 2379 895 2380 899
rect 2374 894 2380 895
rect 2462 899 2468 900
rect 2462 895 2463 899
rect 2467 895 2468 899
rect 2462 894 2468 895
rect 2470 899 2476 900
rect 2470 895 2471 899
rect 2475 898 2476 899
rect 2638 899 2644 900
rect 2475 896 2521 898
rect 2475 895 2476 896
rect 2470 894 2476 895
rect 2638 895 2639 899
rect 2643 895 2644 899
rect 2638 894 2644 895
rect 2726 899 2732 900
rect 2726 895 2727 899
rect 2731 895 2732 899
rect 2726 894 2732 895
rect 2814 899 2820 900
rect 2814 895 2815 899
rect 2819 895 2820 899
rect 2814 894 2820 895
rect 2822 899 2828 900
rect 2822 895 2823 899
rect 2827 898 2828 899
rect 2827 896 2873 898
rect 2827 895 2828 896
rect 2822 894 2828 895
rect 1527 892 1601 894
rect 1527 891 1528 892
rect 1522 890 1528 891
rect 2199 891 2205 892
rect 2126 889 2132 890
rect 1806 888 1812 889
rect 414 885 420 886
rect 110 884 116 885
rect 110 880 111 884
rect 115 880 116 884
rect 414 881 415 885
rect 419 881 420 885
rect 414 880 420 881
rect 558 885 564 886
rect 558 881 559 885
rect 563 881 564 885
rect 558 880 564 881
rect 726 885 732 886
rect 726 881 727 885
rect 731 881 732 885
rect 726 880 732 881
rect 910 885 916 886
rect 910 881 911 885
rect 915 881 916 885
rect 910 880 916 881
rect 1118 885 1124 886
rect 1118 881 1119 885
rect 1123 881 1124 885
rect 1118 880 1124 881
rect 1334 885 1340 886
rect 1334 881 1335 885
rect 1339 881 1340 885
rect 1334 880 1340 881
rect 1558 885 1564 886
rect 1558 881 1559 885
rect 1563 881 1564 885
rect 1558 880 1564 881
rect 1766 884 1772 885
rect 1766 880 1767 884
rect 1771 880 1772 884
rect 1806 884 1807 888
rect 1811 884 1812 888
rect 2126 885 2127 889
rect 2131 885 2132 889
rect 2199 887 2200 891
rect 2204 890 2205 891
rect 2204 888 2210 890
rect 2204 887 2205 888
rect 2199 886 2205 887
rect 2126 884 2132 885
rect 1806 883 1812 884
rect 2208 882 2210 888
rect 2214 889 2220 890
rect 2214 885 2215 889
rect 2219 885 2220 889
rect 2214 884 2220 885
rect 2302 889 2308 890
rect 2302 885 2303 889
rect 2307 885 2308 889
rect 2302 884 2308 885
rect 2390 889 2396 890
rect 2390 885 2391 889
rect 2395 885 2396 889
rect 2390 884 2396 885
rect 2478 889 2484 890
rect 2478 885 2479 889
rect 2483 885 2484 889
rect 2478 884 2484 885
rect 2566 889 2572 890
rect 2566 885 2567 889
rect 2571 885 2572 889
rect 2566 884 2572 885
rect 2654 889 2660 890
rect 2654 885 2655 889
rect 2659 885 2660 889
rect 2654 884 2660 885
rect 2742 889 2748 890
rect 2742 885 2743 889
rect 2747 885 2748 889
rect 2742 884 2748 885
rect 2830 889 2836 890
rect 2830 885 2831 889
rect 2835 885 2836 889
rect 2830 884 2836 885
rect 3462 888 3468 889
rect 3462 884 3463 888
rect 3467 884 3468 888
rect 3462 883 3468 884
rect 2208 880 2222 882
rect 110 879 116 880
rect 1766 879 1772 880
rect 2175 871 2181 872
rect 463 867 469 868
rect 463 863 464 867
rect 468 866 469 867
rect 486 867 492 868
rect 468 864 482 866
rect 468 863 469 864
rect 463 862 469 863
rect 480 858 482 864
rect 486 863 487 867
rect 491 866 492 867
rect 607 867 613 868
rect 607 866 608 867
rect 491 864 608 866
rect 491 863 492 864
rect 486 862 492 863
rect 607 863 608 864
rect 612 863 613 867
rect 607 862 613 863
rect 775 867 781 868
rect 775 863 776 867
rect 780 866 781 867
rect 806 867 812 868
rect 806 866 807 867
rect 780 864 807 866
rect 780 863 781 864
rect 775 862 781 863
rect 806 863 807 864
rect 811 863 812 867
rect 806 862 812 863
rect 959 867 965 868
rect 959 863 960 867
rect 964 866 965 867
rect 990 867 996 868
rect 990 866 991 867
rect 964 864 991 866
rect 964 863 965 864
rect 959 862 965 863
rect 990 863 991 864
rect 995 863 996 867
rect 990 862 996 863
rect 999 867 1005 868
rect 999 863 1000 867
rect 1004 866 1005 867
rect 1167 867 1173 868
rect 1167 866 1168 867
rect 1004 864 1168 866
rect 1004 863 1005 864
rect 999 862 1005 863
rect 1167 863 1168 864
rect 1172 863 1173 867
rect 1167 862 1173 863
rect 1190 867 1196 868
rect 1190 863 1191 867
rect 1195 866 1196 867
rect 1383 867 1389 868
rect 1383 866 1384 867
rect 1195 864 1384 866
rect 1195 863 1196 864
rect 1190 862 1196 863
rect 1383 863 1384 864
rect 1388 863 1389 867
rect 1383 862 1389 863
rect 1607 867 1613 868
rect 1607 863 1608 867
rect 1612 866 1613 867
rect 1654 867 1660 868
rect 1654 866 1655 867
rect 1612 864 1655 866
rect 1612 863 1613 864
rect 1607 862 1613 863
rect 1654 863 1655 864
rect 1659 863 1660 867
rect 2175 867 2176 871
rect 2180 870 2181 871
rect 2206 871 2212 872
rect 2206 870 2207 871
rect 2180 868 2207 870
rect 2180 867 2181 868
rect 2175 866 2181 867
rect 2206 867 2207 868
rect 2211 867 2212 871
rect 2220 870 2222 880
rect 2263 871 2269 872
rect 2263 870 2264 871
rect 2220 868 2264 870
rect 2206 866 2212 867
rect 2263 867 2264 868
rect 2268 867 2269 871
rect 2263 866 2269 867
rect 2286 871 2292 872
rect 2286 867 2287 871
rect 2291 870 2292 871
rect 2351 871 2357 872
rect 2351 870 2352 871
rect 2291 868 2352 870
rect 2291 867 2292 868
rect 2286 866 2292 867
rect 2351 867 2352 868
rect 2356 867 2357 871
rect 2351 866 2357 867
rect 2374 871 2380 872
rect 2374 867 2375 871
rect 2379 870 2380 871
rect 2439 871 2445 872
rect 2439 870 2440 871
rect 2379 868 2440 870
rect 2379 867 2380 868
rect 2374 866 2380 867
rect 2439 867 2440 868
rect 2444 867 2445 871
rect 2439 866 2445 867
rect 2518 871 2524 872
rect 2518 867 2519 871
rect 2523 870 2524 871
rect 2527 871 2533 872
rect 2527 870 2528 871
rect 2523 868 2528 870
rect 2523 867 2524 868
rect 2518 866 2524 867
rect 2527 867 2528 868
rect 2532 867 2533 871
rect 2615 871 2621 872
rect 2615 870 2616 871
rect 2527 866 2533 867
rect 2536 868 2616 870
rect 1654 862 1660 863
rect 2462 863 2468 864
rect 678 859 684 860
rect 678 858 679 859
rect 480 856 679 858
rect 678 855 679 856
rect 683 855 684 859
rect 1230 859 1236 860
rect 1230 858 1231 859
rect 678 854 684 855
rect 1159 856 1231 858
rect 1159 854 1161 856
rect 1230 855 1231 856
rect 1235 855 1236 859
rect 2462 859 2463 863
rect 2467 862 2468 863
rect 2536 862 2538 868
rect 2615 867 2616 868
rect 2620 867 2621 871
rect 2615 866 2621 867
rect 2638 871 2644 872
rect 2638 867 2639 871
rect 2643 870 2644 871
rect 2703 871 2709 872
rect 2703 870 2704 871
rect 2643 868 2704 870
rect 2643 867 2644 868
rect 2638 866 2644 867
rect 2703 867 2704 868
rect 2708 867 2709 871
rect 2703 866 2709 867
rect 2726 871 2732 872
rect 2726 867 2727 871
rect 2731 870 2732 871
rect 2791 871 2797 872
rect 2791 870 2792 871
rect 2731 868 2792 870
rect 2731 867 2732 868
rect 2726 866 2732 867
rect 2791 867 2792 868
rect 2796 867 2797 871
rect 2791 866 2797 867
rect 2814 871 2820 872
rect 2814 867 2815 871
rect 2819 870 2820 871
rect 2879 871 2885 872
rect 2879 870 2880 871
rect 2819 868 2880 870
rect 2819 867 2820 868
rect 2814 866 2820 867
rect 2879 867 2880 868
rect 2884 867 2885 871
rect 2879 866 2885 867
rect 2467 860 2538 862
rect 2467 859 2468 860
rect 2462 858 2468 859
rect 2822 859 2828 860
rect 2822 858 2823 859
rect 1230 854 1236 855
rect 2704 856 2823 858
rect 1108 852 1161 854
rect 183 851 189 852
rect 183 847 184 851
rect 188 850 189 851
rect 214 851 220 852
rect 214 850 215 851
rect 188 848 215 850
rect 188 847 189 848
rect 183 846 189 847
rect 214 847 215 848
rect 219 847 220 851
rect 214 846 220 847
rect 279 851 285 852
rect 279 847 280 851
rect 284 850 285 851
rect 310 851 316 852
rect 310 850 311 851
rect 284 848 311 850
rect 284 847 285 848
rect 279 846 285 847
rect 310 847 311 848
rect 315 847 316 851
rect 310 846 316 847
rect 407 851 413 852
rect 407 847 408 851
rect 412 850 413 851
rect 447 851 453 852
rect 447 850 448 851
rect 412 848 448 850
rect 412 847 413 848
rect 407 846 413 847
rect 447 847 448 848
rect 452 847 453 851
rect 447 846 453 847
rect 535 851 541 852
rect 535 847 536 851
rect 540 850 541 851
rect 567 851 573 852
rect 567 850 568 851
rect 540 848 568 850
rect 540 847 541 848
rect 535 846 541 847
rect 567 847 568 848
rect 572 847 573 851
rect 567 846 573 847
rect 630 851 636 852
rect 630 847 631 851
rect 635 850 636 851
rect 671 851 677 852
rect 671 850 672 851
rect 635 848 672 850
rect 635 847 636 848
rect 630 846 636 847
rect 671 847 672 848
rect 676 847 677 851
rect 671 846 677 847
rect 798 851 805 852
rect 798 847 799 851
rect 804 847 805 851
rect 798 846 805 847
rect 822 851 828 852
rect 822 847 823 851
rect 827 850 828 851
rect 927 851 933 852
rect 927 850 928 851
rect 827 848 928 850
rect 827 847 828 848
rect 822 846 828 847
rect 927 847 928 848
rect 932 847 933 851
rect 927 846 933 847
rect 1055 851 1061 852
rect 1055 847 1056 851
rect 1060 850 1061 851
rect 1108 850 1110 852
rect 1183 851 1189 852
rect 1183 850 1184 851
rect 1060 848 1110 850
rect 1159 848 1184 850
rect 1060 847 1061 848
rect 1055 846 1061 847
rect 1114 847 1120 848
rect 1114 843 1115 847
rect 1119 846 1120 847
rect 1159 846 1161 848
rect 1183 847 1184 848
rect 1188 847 1189 851
rect 1183 846 1189 847
rect 1319 851 1328 852
rect 1319 847 1320 851
rect 1327 847 1328 851
rect 1319 846 1328 847
rect 2207 851 2213 852
rect 2207 847 2208 851
rect 2212 850 2213 851
rect 2222 851 2228 852
rect 2222 850 2223 851
rect 2212 848 2223 850
rect 2212 847 2213 848
rect 2207 846 2213 847
rect 2222 847 2223 848
rect 2227 847 2228 851
rect 2222 846 2228 847
rect 2230 851 2236 852
rect 2230 847 2231 851
rect 2235 850 2236 851
rect 2295 851 2301 852
rect 2295 850 2296 851
rect 2235 848 2296 850
rect 2235 847 2236 848
rect 2230 846 2236 847
rect 2295 847 2296 848
rect 2300 847 2301 851
rect 2295 846 2301 847
rect 2318 851 2324 852
rect 2318 847 2319 851
rect 2323 850 2324 851
rect 2383 851 2389 852
rect 2383 850 2384 851
rect 2323 848 2384 850
rect 2323 847 2324 848
rect 2318 846 2324 847
rect 2383 847 2384 848
rect 2388 847 2389 851
rect 2383 846 2389 847
rect 2406 851 2412 852
rect 2406 847 2407 851
rect 2411 850 2412 851
rect 2471 851 2477 852
rect 2471 850 2472 851
rect 2411 848 2472 850
rect 2411 847 2412 848
rect 2406 846 2412 847
rect 2471 847 2472 848
rect 2476 847 2477 851
rect 2471 846 2477 847
rect 2494 851 2500 852
rect 2494 847 2495 851
rect 2499 850 2500 851
rect 2575 851 2581 852
rect 2575 850 2576 851
rect 2499 848 2576 850
rect 2499 847 2500 848
rect 2494 846 2500 847
rect 2575 847 2576 848
rect 2580 847 2581 851
rect 2575 846 2581 847
rect 2687 851 2693 852
rect 2687 847 2688 851
rect 2692 850 2693 851
rect 2704 850 2706 856
rect 2822 855 2823 856
rect 2827 855 2828 859
rect 2822 854 2828 855
rect 2692 848 2706 850
rect 2710 851 2716 852
rect 2692 847 2693 848
rect 2687 846 2693 847
rect 2710 847 2711 851
rect 2715 850 2716 851
rect 2815 851 2821 852
rect 2815 850 2816 851
rect 2715 848 2816 850
rect 2715 847 2716 848
rect 2710 846 2716 847
rect 2815 847 2816 848
rect 2820 847 2821 851
rect 2815 846 2821 847
rect 2838 851 2844 852
rect 2838 847 2839 851
rect 2843 850 2844 851
rect 2959 851 2965 852
rect 2959 850 2960 851
rect 2843 848 2960 850
rect 2843 847 2844 848
rect 2838 846 2844 847
rect 2959 847 2960 848
rect 2964 847 2965 851
rect 2959 846 2965 847
rect 2982 851 2988 852
rect 2982 847 2983 851
rect 2987 850 2988 851
rect 3111 851 3117 852
rect 3111 850 3112 851
rect 2987 848 3112 850
rect 2987 847 2988 848
rect 2982 846 2988 847
rect 3111 847 3112 848
rect 3116 847 3117 851
rect 3111 846 3117 847
rect 3190 851 3196 852
rect 3190 847 3191 851
rect 3195 850 3196 851
rect 3271 851 3277 852
rect 3271 850 3272 851
rect 3195 848 3272 850
rect 3195 847 3196 848
rect 3190 846 3196 847
rect 3271 847 3272 848
rect 3276 847 3277 851
rect 3271 846 3277 847
rect 3415 851 3421 852
rect 3415 847 3416 851
rect 3420 850 3421 851
rect 3438 851 3444 852
rect 3438 850 3439 851
rect 3420 848 3439 850
rect 3420 847 3421 848
rect 3415 846 3421 847
rect 3438 847 3439 848
rect 3443 847 3444 851
rect 3438 846 3444 847
rect 1119 844 1161 846
rect 1119 843 1120 844
rect 1114 842 1120 843
rect 110 836 116 837
rect 1766 836 1772 837
rect 110 832 111 836
rect 115 832 116 836
rect 110 831 116 832
rect 134 835 140 836
rect 134 831 135 835
rect 139 831 140 835
rect 134 830 140 831
rect 230 835 236 836
rect 230 831 231 835
rect 235 831 236 835
rect 230 830 236 831
rect 358 835 364 836
rect 358 831 359 835
rect 363 831 364 835
rect 358 830 364 831
rect 486 835 492 836
rect 486 831 487 835
rect 491 831 492 835
rect 486 830 492 831
rect 622 835 628 836
rect 622 831 623 835
rect 627 831 628 835
rect 622 830 628 831
rect 750 835 756 836
rect 750 831 751 835
rect 755 831 756 835
rect 750 830 756 831
rect 878 835 884 836
rect 878 831 879 835
rect 883 831 884 835
rect 878 830 884 831
rect 1006 835 1012 836
rect 1006 831 1007 835
rect 1011 831 1012 835
rect 1006 830 1012 831
rect 1134 835 1140 836
rect 1134 831 1135 835
rect 1139 831 1140 835
rect 1134 830 1140 831
rect 1270 835 1276 836
rect 1270 831 1271 835
rect 1275 831 1276 835
rect 1766 832 1767 836
rect 1771 832 1772 836
rect 1766 831 1772 832
rect 1806 836 1812 837
rect 3462 836 3468 837
rect 1806 832 1807 836
rect 1811 832 1812 836
rect 1806 831 1812 832
rect 2158 835 2164 836
rect 2158 831 2159 835
rect 2163 831 2164 835
rect 1270 830 1276 831
rect 2158 830 2164 831
rect 2246 835 2252 836
rect 2246 831 2247 835
rect 2251 831 2252 835
rect 2246 830 2252 831
rect 2334 835 2340 836
rect 2334 831 2335 835
rect 2339 831 2340 835
rect 2334 830 2340 831
rect 2422 835 2428 836
rect 2422 831 2423 835
rect 2427 831 2428 835
rect 2422 830 2428 831
rect 2526 835 2532 836
rect 2526 831 2527 835
rect 2531 831 2532 835
rect 2526 830 2532 831
rect 2638 835 2644 836
rect 2638 831 2639 835
rect 2643 831 2644 835
rect 2638 830 2644 831
rect 2766 835 2772 836
rect 2766 831 2767 835
rect 2771 831 2772 835
rect 2766 830 2772 831
rect 2910 835 2916 836
rect 2910 831 2911 835
rect 2915 831 2916 835
rect 2910 830 2916 831
rect 3062 835 3068 836
rect 3062 831 3063 835
rect 3067 831 3068 835
rect 3062 830 3068 831
rect 3222 835 3228 836
rect 3222 831 3223 835
rect 3227 831 3228 835
rect 3222 830 3228 831
rect 3366 835 3372 836
rect 3366 831 3367 835
rect 3371 831 3372 835
rect 3462 832 3463 836
rect 3467 832 3468 836
rect 3462 831 3468 832
rect 3366 830 3372 831
rect 214 827 220 828
rect 214 823 215 827
rect 219 826 220 827
rect 310 827 316 828
rect 219 824 273 826
rect 219 823 220 824
rect 214 822 220 823
rect 310 823 311 827
rect 315 826 316 827
rect 447 827 453 828
rect 315 824 401 826
rect 315 823 316 824
rect 310 822 316 823
rect 447 823 448 827
rect 452 826 453 827
rect 567 827 573 828
rect 452 824 529 826
rect 452 823 453 824
rect 447 822 453 823
rect 567 823 568 827
rect 572 826 573 827
rect 822 827 828 828
rect 572 824 665 826
rect 572 823 573 824
rect 567 822 573 823
rect 822 823 823 827
rect 827 823 828 827
rect 999 827 1005 828
rect 999 826 1000 827
rect 953 824 1000 826
rect 822 822 828 823
rect 999 823 1000 824
rect 1004 823 1005 827
rect 1114 827 1120 828
rect 1114 826 1115 827
rect 1081 824 1115 826
rect 999 822 1005 823
rect 1114 823 1115 824
rect 1119 823 1120 827
rect 1230 827 1236 828
rect 1114 822 1120 823
rect 1206 823 1212 824
rect 110 819 116 820
rect 110 815 111 819
rect 115 815 116 819
rect 198 819 204 820
rect 110 814 116 815
rect 134 816 140 817
rect 134 812 135 816
rect 139 812 140 816
rect 198 815 199 819
rect 203 818 204 819
rect 208 818 210 821
rect 1206 819 1207 823
rect 1211 819 1212 823
rect 1230 823 1231 827
rect 1235 826 1236 827
rect 2230 827 2236 828
rect 1235 824 1313 826
rect 1235 823 1236 824
rect 1230 822 1236 823
rect 2230 823 2231 827
rect 2235 823 2236 827
rect 2230 822 2236 823
rect 2318 827 2324 828
rect 2318 823 2319 827
rect 2323 823 2324 827
rect 2318 822 2324 823
rect 2406 827 2412 828
rect 2406 823 2407 827
rect 2411 823 2412 827
rect 2406 822 2412 823
rect 2494 827 2500 828
rect 2494 823 2495 827
rect 2499 823 2500 827
rect 2494 822 2500 823
rect 2518 827 2524 828
rect 2518 823 2519 827
rect 2523 826 2524 827
rect 2710 827 2716 828
rect 2523 824 2569 826
rect 2523 823 2524 824
rect 2518 822 2524 823
rect 2710 823 2711 827
rect 2715 823 2716 827
rect 2710 822 2716 823
rect 2838 827 2844 828
rect 2838 823 2839 827
rect 2843 823 2844 827
rect 2838 822 2844 823
rect 2982 827 2988 828
rect 2982 823 2983 827
rect 2987 823 2988 827
rect 2982 822 2988 823
rect 2990 827 2996 828
rect 2990 823 2991 827
rect 2995 826 2996 827
rect 3294 827 3300 828
rect 2995 824 3105 826
rect 2995 823 2996 824
rect 2990 822 2996 823
rect 3294 823 3295 827
rect 3299 823 3300 827
rect 3294 822 3300 823
rect 3438 823 3444 824
rect 1206 818 1212 819
rect 1766 819 1772 820
rect 203 816 210 818
rect 230 816 236 817
rect 203 815 204 816
rect 198 814 204 815
rect 134 811 140 812
rect 230 812 231 816
rect 235 812 236 816
rect 230 811 236 812
rect 358 816 364 817
rect 358 812 359 816
rect 363 812 364 816
rect 358 811 364 812
rect 486 816 492 817
rect 486 812 487 816
rect 491 812 492 816
rect 486 811 492 812
rect 622 816 628 817
rect 622 812 623 816
rect 627 812 628 816
rect 622 811 628 812
rect 750 816 756 817
rect 750 812 751 816
rect 755 812 756 816
rect 750 811 756 812
rect 878 816 884 817
rect 878 812 879 816
rect 883 812 884 816
rect 878 811 884 812
rect 1006 816 1012 817
rect 1006 812 1007 816
rect 1011 812 1012 816
rect 1006 811 1012 812
rect 1134 816 1140 817
rect 1134 812 1135 816
rect 1139 812 1140 816
rect 1134 811 1140 812
rect 1270 816 1276 817
rect 1270 812 1271 816
rect 1275 812 1276 816
rect 1766 815 1767 819
rect 1771 815 1772 819
rect 1766 814 1772 815
rect 1806 819 1812 820
rect 1806 815 1807 819
rect 1811 815 1812 819
rect 3438 819 3439 823
rect 3443 819 3444 823
rect 3438 818 3444 819
rect 3462 819 3468 820
rect 1806 814 1812 815
rect 2158 816 2164 817
rect 1270 811 1276 812
rect 2158 812 2159 816
rect 2163 812 2164 816
rect 2158 811 2164 812
rect 2246 816 2252 817
rect 2246 812 2247 816
rect 2251 812 2252 816
rect 2246 811 2252 812
rect 2334 816 2340 817
rect 2334 812 2335 816
rect 2339 812 2340 816
rect 2334 811 2340 812
rect 2422 816 2428 817
rect 2422 812 2423 816
rect 2427 812 2428 816
rect 2422 811 2428 812
rect 2526 816 2532 817
rect 2526 812 2527 816
rect 2531 812 2532 816
rect 2526 811 2532 812
rect 2638 816 2644 817
rect 2638 812 2639 816
rect 2643 812 2644 816
rect 2638 811 2644 812
rect 2766 816 2772 817
rect 2766 812 2767 816
rect 2771 812 2772 816
rect 2766 811 2772 812
rect 2910 816 2916 817
rect 2910 812 2911 816
rect 2915 812 2916 816
rect 2910 811 2916 812
rect 3062 816 3068 817
rect 3062 812 3063 816
rect 3067 812 3068 816
rect 3062 811 3068 812
rect 3222 816 3228 817
rect 3222 812 3223 816
rect 3227 812 3228 816
rect 3222 811 3228 812
rect 3366 816 3372 817
rect 3366 812 3367 816
rect 3371 812 3372 816
rect 3462 815 3463 819
rect 3467 815 3468 819
rect 3462 814 3468 815
rect 3366 811 3372 812
rect 2762 779 2768 780
rect 2222 775 2228 776
rect 2222 771 2223 775
rect 2227 774 2228 775
rect 2762 775 2763 779
rect 2767 778 2768 779
rect 2990 779 2996 780
rect 2990 778 2991 779
rect 2767 776 2991 778
rect 2767 775 2768 776
rect 2762 774 2768 775
rect 2990 775 2991 776
rect 2995 775 2996 779
rect 2990 774 2996 775
rect 2227 772 2506 774
rect 2227 771 2228 772
rect 2222 770 2228 771
rect 134 768 140 769
rect 110 765 116 766
rect 110 761 111 765
rect 115 761 116 765
rect 134 764 135 768
rect 139 764 140 768
rect 134 763 140 764
rect 222 768 228 769
rect 222 764 223 768
rect 227 764 228 768
rect 222 763 228 764
rect 342 768 348 769
rect 342 764 343 768
rect 347 764 348 768
rect 342 763 348 764
rect 470 768 476 769
rect 470 764 471 768
rect 475 764 476 768
rect 470 763 476 764
rect 606 768 612 769
rect 606 764 607 768
rect 611 764 612 768
rect 606 763 612 764
rect 742 768 748 769
rect 742 764 743 768
rect 747 764 748 768
rect 742 763 748 764
rect 886 768 892 769
rect 886 764 887 768
rect 891 764 892 768
rect 886 763 892 764
rect 1038 768 1044 769
rect 1038 764 1039 768
rect 1043 764 1044 768
rect 1038 763 1044 764
rect 1190 768 1196 769
rect 1190 764 1191 768
rect 1195 764 1196 768
rect 1190 763 1196 764
rect 1350 768 1356 769
rect 1350 764 1351 768
rect 1355 764 1356 768
rect 2062 768 2068 769
rect 1350 763 1356 764
rect 1766 765 1772 766
rect 110 760 116 761
rect 1766 761 1767 765
rect 1771 761 1772 765
rect 1766 760 1772 761
rect 1806 765 1812 766
rect 1806 761 1807 765
rect 1811 761 1812 765
rect 2062 764 2063 768
rect 2067 764 2068 768
rect 2062 763 2068 764
rect 2174 768 2180 769
rect 2174 764 2175 768
rect 2179 764 2180 768
rect 2174 763 2180 764
rect 2294 768 2300 769
rect 2294 764 2295 768
rect 2299 764 2300 768
rect 2294 763 2300 764
rect 2422 768 2428 769
rect 2422 764 2423 768
rect 2427 764 2428 768
rect 2422 763 2428 764
rect 1806 760 1812 761
rect 206 759 212 760
rect 206 755 207 759
rect 211 755 212 759
rect 206 754 212 755
rect 294 759 300 760
rect 294 755 295 759
rect 299 755 300 759
rect 294 754 300 755
rect 414 759 420 760
rect 414 755 415 759
rect 419 755 420 759
rect 414 754 420 755
rect 542 759 548 760
rect 542 755 543 759
rect 547 755 548 759
rect 542 754 548 755
rect 550 759 556 760
rect 550 755 551 759
rect 555 758 556 759
rect 806 759 812 760
rect 555 756 649 758
rect 555 755 556 756
rect 550 754 556 755
rect 806 755 807 759
rect 811 755 812 759
rect 806 754 812 755
rect 822 759 828 760
rect 822 755 823 759
rect 827 758 828 759
rect 966 759 972 760
rect 827 756 929 758
rect 827 755 828 756
rect 822 754 828 755
rect 966 755 967 759
rect 971 758 972 759
rect 1262 759 1268 760
rect 971 756 1081 758
rect 971 755 972 756
rect 966 754 972 755
rect 1262 755 1263 759
rect 1267 755 1268 759
rect 1470 759 1476 760
rect 1470 758 1471 759
rect 1425 756 1471 758
rect 1262 754 1268 755
rect 1470 755 1471 756
rect 1475 755 1476 759
rect 1470 754 1476 755
rect 2134 759 2140 760
rect 2134 755 2135 759
rect 2139 755 2140 759
rect 2134 754 2140 755
rect 2246 759 2252 760
rect 2246 755 2247 759
rect 2251 755 2252 759
rect 2246 754 2252 755
rect 2366 759 2372 760
rect 2366 755 2367 759
rect 2371 755 2372 759
rect 2366 754 2372 755
rect 2494 759 2500 760
rect 2494 755 2495 759
rect 2499 755 2500 759
rect 2504 758 2506 772
rect 2558 768 2564 769
rect 2558 764 2559 768
rect 2563 764 2564 768
rect 2558 763 2564 764
rect 2710 768 2716 769
rect 2710 764 2711 768
rect 2715 764 2716 768
rect 2710 763 2716 764
rect 2870 768 2876 769
rect 2870 764 2871 768
rect 2875 764 2876 768
rect 2870 763 2876 764
rect 3038 768 3044 769
rect 3038 764 3039 768
rect 3043 764 3044 768
rect 3038 763 3044 764
rect 3214 768 3220 769
rect 3214 764 3215 768
rect 3219 764 3220 768
rect 3214 763 3220 764
rect 3366 768 3372 769
rect 3366 764 3367 768
rect 3371 764 3372 768
rect 3366 763 3372 764
rect 3462 765 3468 766
rect 3462 761 3463 765
rect 3467 761 3468 765
rect 3462 760 3468 761
rect 2782 759 2788 760
rect 2504 756 2601 758
rect 2494 754 2500 755
rect 2782 755 2783 759
rect 2787 755 2788 759
rect 2782 754 2788 755
rect 2942 759 2948 760
rect 2942 755 2943 759
rect 2947 755 2948 759
rect 2942 754 2948 755
rect 3110 759 3116 760
rect 3110 755 3111 759
rect 3115 755 3116 759
rect 3110 754 3116 755
rect 3119 759 3125 760
rect 3119 755 3120 759
rect 3124 758 3125 759
rect 3430 759 3436 760
rect 3124 756 3257 758
rect 3124 755 3125 756
rect 3119 754 3125 755
rect 3430 755 3431 759
rect 3435 755 3436 759
rect 3430 754 3436 755
rect 134 749 140 750
rect 110 748 116 749
rect 110 744 111 748
rect 115 744 116 748
rect 134 745 135 749
rect 139 745 140 749
rect 134 744 140 745
rect 222 749 228 750
rect 222 745 223 749
rect 227 745 228 749
rect 222 744 228 745
rect 342 749 348 750
rect 342 745 343 749
rect 347 745 348 749
rect 342 744 348 745
rect 470 749 476 750
rect 470 745 471 749
rect 475 745 476 749
rect 470 744 476 745
rect 606 749 612 750
rect 606 745 607 749
rect 611 745 612 749
rect 606 744 612 745
rect 742 749 748 750
rect 742 745 743 749
rect 747 745 748 749
rect 742 744 748 745
rect 886 749 892 750
rect 886 745 887 749
rect 891 745 892 749
rect 886 744 892 745
rect 1038 749 1044 750
rect 1038 745 1039 749
rect 1043 745 1044 749
rect 1038 744 1044 745
rect 1190 749 1196 750
rect 1190 745 1191 749
rect 1195 745 1196 749
rect 1190 744 1196 745
rect 1350 749 1356 750
rect 2062 749 2068 750
rect 1350 745 1351 749
rect 1355 745 1356 749
rect 1350 744 1356 745
rect 1766 748 1772 749
rect 1766 744 1767 748
rect 1771 744 1772 748
rect 110 743 116 744
rect 1766 743 1772 744
rect 1806 748 1812 749
rect 1806 744 1807 748
rect 1811 744 1812 748
rect 2062 745 2063 749
rect 2067 745 2068 749
rect 2062 744 2068 745
rect 2174 749 2180 750
rect 2174 745 2175 749
rect 2179 745 2180 749
rect 2174 744 2180 745
rect 2294 749 2300 750
rect 2294 745 2295 749
rect 2299 745 2300 749
rect 2294 744 2300 745
rect 2422 749 2428 750
rect 2422 745 2423 749
rect 2427 745 2428 749
rect 2422 744 2428 745
rect 2558 749 2564 750
rect 2558 745 2559 749
rect 2563 745 2564 749
rect 2558 744 2564 745
rect 2710 749 2716 750
rect 2710 745 2711 749
rect 2715 745 2716 749
rect 2710 744 2716 745
rect 2870 749 2876 750
rect 2870 745 2871 749
rect 2875 745 2876 749
rect 2870 744 2876 745
rect 3038 749 3044 750
rect 3038 745 3039 749
rect 3043 745 3044 749
rect 3038 744 3044 745
rect 3214 749 3220 750
rect 3214 745 3215 749
rect 3219 745 3220 749
rect 3214 744 3220 745
rect 3366 749 3372 750
rect 3366 745 3367 749
rect 3371 745 3372 749
rect 3366 744 3372 745
rect 3462 748 3468 749
rect 3462 744 3463 748
rect 3467 744 3468 748
rect 1806 743 1812 744
rect 3462 743 3468 744
rect 183 731 189 732
rect 183 727 184 731
rect 188 730 189 731
rect 198 731 204 732
rect 198 730 199 731
rect 188 728 199 730
rect 188 727 189 728
rect 183 726 189 727
rect 198 727 199 728
rect 203 727 204 731
rect 198 726 204 727
rect 206 731 212 732
rect 206 727 207 731
rect 211 730 212 731
rect 271 731 277 732
rect 271 730 272 731
rect 211 728 272 730
rect 211 727 212 728
rect 206 726 212 727
rect 271 727 272 728
rect 276 727 277 731
rect 271 726 277 727
rect 294 731 300 732
rect 294 727 295 731
rect 299 730 300 731
rect 391 731 397 732
rect 391 730 392 731
rect 299 728 392 730
rect 299 727 300 728
rect 294 726 300 727
rect 391 727 392 728
rect 396 727 397 731
rect 391 726 397 727
rect 414 731 420 732
rect 414 727 415 731
rect 419 730 420 731
rect 519 731 525 732
rect 519 730 520 731
rect 419 728 520 730
rect 419 727 420 728
rect 414 726 420 727
rect 519 727 520 728
rect 524 727 525 731
rect 519 726 525 727
rect 542 731 548 732
rect 542 727 543 731
rect 547 730 548 731
rect 655 731 661 732
rect 655 730 656 731
rect 547 728 656 730
rect 547 727 548 728
rect 542 726 548 727
rect 655 727 656 728
rect 660 727 661 731
rect 655 726 661 727
rect 791 731 797 732
rect 791 727 792 731
rect 796 730 797 731
rect 822 731 828 732
rect 822 730 823 731
rect 796 728 823 730
rect 796 727 797 728
rect 791 726 797 727
rect 822 727 823 728
rect 827 727 828 731
rect 822 726 828 727
rect 935 731 941 732
rect 935 727 936 731
rect 940 730 941 731
rect 966 731 972 732
rect 966 730 967 731
rect 940 728 967 730
rect 940 727 941 728
rect 935 726 941 727
rect 966 727 967 728
rect 971 727 972 731
rect 966 726 972 727
rect 1087 731 1093 732
rect 1087 727 1088 731
rect 1092 730 1093 731
rect 1102 731 1108 732
rect 1102 730 1103 731
rect 1092 728 1103 730
rect 1092 727 1093 728
rect 1087 726 1093 727
rect 1102 727 1103 728
rect 1107 727 1108 731
rect 1102 726 1108 727
rect 1206 731 1212 732
rect 1206 727 1207 731
rect 1211 730 1212 731
rect 1239 731 1245 732
rect 1239 730 1240 731
rect 1211 728 1240 730
rect 1211 727 1212 728
rect 1206 726 1212 727
rect 1239 727 1240 728
rect 1244 727 1245 731
rect 1239 726 1245 727
rect 1262 731 1268 732
rect 1262 727 1263 731
rect 1267 730 1268 731
rect 1399 731 1405 732
rect 1399 730 1400 731
rect 1267 728 1400 730
rect 1267 727 1268 728
rect 1262 726 1268 727
rect 1399 727 1400 728
rect 1404 727 1405 731
rect 1399 726 1405 727
rect 2111 731 2120 732
rect 2111 727 2112 731
rect 2119 727 2120 731
rect 2111 726 2120 727
rect 2134 731 2140 732
rect 2134 727 2135 731
rect 2139 730 2140 731
rect 2223 731 2229 732
rect 2223 730 2224 731
rect 2139 728 2224 730
rect 2139 727 2140 728
rect 2134 726 2140 727
rect 2223 727 2224 728
rect 2228 727 2229 731
rect 2223 726 2229 727
rect 2246 731 2252 732
rect 2246 727 2247 731
rect 2251 730 2252 731
rect 2343 731 2349 732
rect 2343 730 2344 731
rect 2251 728 2344 730
rect 2251 727 2252 728
rect 2246 726 2252 727
rect 2343 727 2344 728
rect 2348 727 2349 731
rect 2343 726 2349 727
rect 2366 731 2372 732
rect 2366 727 2367 731
rect 2371 730 2372 731
rect 2471 731 2477 732
rect 2471 730 2472 731
rect 2371 728 2472 730
rect 2371 727 2372 728
rect 2366 726 2372 727
rect 2471 727 2472 728
rect 2476 727 2477 731
rect 2471 726 2477 727
rect 2494 731 2500 732
rect 2494 727 2495 731
rect 2499 730 2500 731
rect 2607 731 2613 732
rect 2607 730 2608 731
rect 2499 728 2608 730
rect 2499 727 2500 728
rect 2494 726 2500 727
rect 2607 727 2608 728
rect 2612 727 2613 731
rect 2607 726 2613 727
rect 2759 731 2768 732
rect 2759 727 2760 731
rect 2767 727 2768 731
rect 2759 726 2768 727
rect 2782 731 2788 732
rect 2782 727 2783 731
rect 2787 730 2788 731
rect 2919 731 2925 732
rect 2919 730 2920 731
rect 2787 728 2920 730
rect 2787 727 2788 728
rect 2782 726 2788 727
rect 2919 727 2920 728
rect 2924 727 2925 731
rect 2919 726 2925 727
rect 2942 731 2948 732
rect 2942 727 2943 731
rect 2947 730 2948 731
rect 3087 731 3093 732
rect 3087 730 3088 731
rect 2947 728 3088 730
rect 2947 727 2948 728
rect 2942 726 2948 727
rect 3087 727 3088 728
rect 3092 727 3093 731
rect 3087 726 3093 727
rect 3110 731 3116 732
rect 3110 727 3111 731
rect 3115 730 3116 731
rect 3263 731 3269 732
rect 3263 730 3264 731
rect 3115 728 3264 730
rect 3115 727 3116 728
rect 3110 726 3116 727
rect 3263 727 3264 728
rect 3268 727 3269 731
rect 3263 726 3269 727
rect 3415 731 3421 732
rect 3415 727 3416 731
rect 3420 730 3421 731
rect 3438 731 3444 732
rect 3438 730 3439 731
rect 3420 728 3439 730
rect 3420 727 3421 728
rect 3415 726 3421 727
rect 3438 727 3439 728
rect 3443 727 3444 731
rect 3438 726 3444 727
rect 550 723 556 724
rect 550 722 551 723
rect 319 720 551 722
rect 319 718 321 720
rect 550 719 551 720
rect 555 719 556 723
rect 550 718 556 719
rect 1975 719 1981 720
rect 268 716 321 718
rect 215 715 221 716
rect 215 711 216 715
rect 220 714 221 715
rect 268 714 270 716
rect 343 715 349 716
rect 343 714 344 715
rect 220 712 270 714
rect 319 712 344 714
rect 220 711 221 712
rect 215 710 221 711
rect 274 711 280 712
rect 274 707 275 711
rect 279 710 280 711
rect 319 710 321 712
rect 343 711 344 712
rect 348 711 349 715
rect 343 710 349 711
rect 366 715 372 716
rect 366 711 367 715
rect 371 714 372 715
rect 479 715 485 716
rect 479 714 480 715
rect 371 712 480 714
rect 371 711 372 712
rect 366 710 372 711
rect 479 711 480 712
rect 484 711 485 715
rect 479 710 485 711
rect 502 715 508 716
rect 502 711 503 715
rect 507 714 508 715
rect 623 715 629 716
rect 623 714 624 715
rect 507 712 624 714
rect 507 711 508 712
rect 502 710 508 711
rect 623 711 624 712
rect 628 711 629 715
rect 623 710 629 711
rect 646 715 652 716
rect 646 711 647 715
rect 651 714 652 715
rect 775 715 781 716
rect 775 714 776 715
rect 651 712 776 714
rect 651 711 652 712
rect 646 710 652 711
rect 775 711 776 712
rect 780 711 781 715
rect 775 710 781 711
rect 927 715 933 716
rect 927 711 928 715
rect 932 714 933 715
rect 942 715 948 716
rect 942 714 943 715
rect 932 712 943 714
rect 932 711 933 712
rect 927 710 933 711
rect 942 711 943 712
rect 947 711 948 715
rect 942 710 948 711
rect 950 715 956 716
rect 950 711 951 715
rect 955 714 956 715
rect 1079 715 1085 716
rect 1079 714 1080 715
rect 955 712 1080 714
rect 955 711 956 712
rect 950 710 956 711
rect 1079 711 1080 712
rect 1084 711 1085 715
rect 1079 710 1085 711
rect 1231 715 1237 716
rect 1231 711 1232 715
rect 1236 714 1237 715
rect 1262 715 1268 716
rect 1262 714 1263 715
rect 1236 712 1263 714
rect 1236 711 1237 712
rect 1231 710 1237 711
rect 1262 711 1263 712
rect 1267 711 1268 715
rect 1262 710 1268 711
rect 1391 715 1397 716
rect 1391 711 1392 715
rect 1396 714 1397 715
rect 1422 715 1428 716
rect 1422 714 1423 715
rect 1396 712 1423 714
rect 1396 711 1397 712
rect 1391 710 1397 711
rect 1422 711 1423 712
rect 1427 711 1428 715
rect 1422 710 1428 711
rect 1470 715 1476 716
rect 1470 711 1471 715
rect 1475 714 1476 715
rect 1551 715 1557 716
rect 1551 714 1552 715
rect 1475 712 1552 714
rect 1475 711 1476 712
rect 1470 710 1476 711
rect 1551 711 1552 712
rect 1556 711 1557 715
rect 1975 715 1976 719
rect 1980 718 1981 719
rect 1986 719 1992 720
rect 1986 718 1987 719
rect 1980 716 1987 718
rect 1980 715 1981 716
rect 1975 714 1981 715
rect 1986 715 1987 716
rect 1991 715 1992 719
rect 1986 714 1992 715
rect 1998 719 2004 720
rect 1998 715 1999 719
rect 2003 718 2004 719
rect 2119 719 2125 720
rect 2119 718 2120 719
rect 2003 716 2120 718
rect 2003 715 2004 716
rect 1998 714 2004 715
rect 2119 715 2120 716
rect 2124 715 2125 719
rect 2119 714 2125 715
rect 2142 719 2148 720
rect 2142 715 2143 719
rect 2147 718 2148 719
rect 2279 719 2285 720
rect 2279 718 2280 719
rect 2147 716 2280 718
rect 2147 715 2148 716
rect 2142 714 2148 715
rect 2279 715 2280 716
rect 2284 715 2285 719
rect 2279 714 2285 715
rect 2302 719 2308 720
rect 2302 715 2303 719
rect 2307 718 2308 719
rect 2439 719 2445 720
rect 2439 718 2440 719
rect 2307 716 2440 718
rect 2307 715 2308 716
rect 2302 714 2308 715
rect 2439 715 2440 716
rect 2444 715 2445 719
rect 2439 714 2445 715
rect 2462 719 2468 720
rect 2462 715 2463 719
rect 2467 718 2468 719
rect 2599 719 2605 720
rect 2599 718 2600 719
rect 2467 716 2600 718
rect 2467 715 2468 716
rect 2462 714 2468 715
rect 2599 715 2600 716
rect 2604 715 2605 719
rect 2599 714 2605 715
rect 2751 719 2757 720
rect 2751 715 2752 719
rect 2756 718 2757 719
rect 2794 719 2800 720
rect 2794 718 2795 719
rect 2756 716 2795 718
rect 2756 715 2757 716
rect 2751 714 2757 715
rect 2794 715 2795 716
rect 2799 715 2800 719
rect 2794 714 2800 715
rect 2895 719 2901 720
rect 2895 715 2896 719
rect 2900 718 2901 719
rect 2927 719 2933 720
rect 2927 718 2928 719
rect 2900 716 2928 718
rect 2900 715 2901 716
rect 2895 714 2901 715
rect 2927 715 2928 716
rect 2932 715 2933 719
rect 2927 714 2933 715
rect 3031 719 3037 720
rect 3031 715 3032 719
rect 3036 718 3037 719
rect 3119 719 3125 720
rect 3119 718 3120 719
rect 3036 716 3120 718
rect 3036 715 3037 716
rect 3031 714 3037 715
rect 3119 715 3120 716
rect 3124 715 3125 719
rect 3119 714 3125 715
rect 3167 719 3173 720
rect 3167 715 3168 719
rect 3172 718 3173 719
rect 3198 719 3204 720
rect 3198 718 3199 719
rect 3172 716 3199 718
rect 3172 715 3173 716
rect 3167 714 3173 715
rect 3198 715 3199 716
rect 3203 715 3204 719
rect 3198 714 3204 715
rect 3302 719 3309 720
rect 3302 715 3303 719
rect 3308 715 3309 719
rect 3302 714 3309 715
rect 3415 719 3421 720
rect 3415 715 3416 719
rect 3420 718 3421 719
rect 3430 719 3436 720
rect 3430 718 3431 719
rect 3420 716 3431 718
rect 3420 715 3421 716
rect 3415 714 3421 715
rect 3430 715 3431 716
rect 3435 715 3436 719
rect 3430 714 3436 715
rect 1551 710 1557 711
rect 279 708 321 710
rect 279 707 280 708
rect 274 706 280 707
rect 1806 704 1812 705
rect 3462 704 3468 705
rect 110 700 116 701
rect 1766 700 1772 701
rect 110 696 111 700
rect 115 696 116 700
rect 110 695 116 696
rect 166 699 172 700
rect 166 695 167 699
rect 171 695 172 699
rect 166 694 172 695
rect 294 699 300 700
rect 294 695 295 699
rect 299 695 300 699
rect 294 694 300 695
rect 430 699 436 700
rect 430 695 431 699
rect 435 695 436 699
rect 430 694 436 695
rect 574 699 580 700
rect 574 695 575 699
rect 579 695 580 699
rect 574 694 580 695
rect 726 699 732 700
rect 726 695 727 699
rect 731 695 732 699
rect 726 694 732 695
rect 878 699 884 700
rect 878 695 879 699
rect 883 695 884 699
rect 878 694 884 695
rect 1030 699 1036 700
rect 1030 695 1031 699
rect 1035 695 1036 699
rect 1030 694 1036 695
rect 1182 699 1188 700
rect 1182 695 1183 699
rect 1187 695 1188 699
rect 1182 694 1188 695
rect 1342 699 1348 700
rect 1342 695 1343 699
rect 1347 695 1348 699
rect 1342 694 1348 695
rect 1502 699 1508 700
rect 1502 695 1503 699
rect 1507 695 1508 699
rect 1766 696 1767 700
rect 1771 696 1772 700
rect 1806 700 1807 704
rect 1811 700 1812 704
rect 1806 699 1812 700
rect 1926 703 1932 704
rect 1926 699 1927 703
rect 1931 699 1932 703
rect 1926 698 1932 699
rect 2070 703 2076 704
rect 2070 699 2071 703
rect 2075 699 2076 703
rect 2070 698 2076 699
rect 2230 703 2236 704
rect 2230 699 2231 703
rect 2235 699 2236 703
rect 2230 698 2236 699
rect 2390 703 2396 704
rect 2390 699 2391 703
rect 2395 699 2396 703
rect 2390 698 2396 699
rect 2550 703 2556 704
rect 2550 699 2551 703
rect 2555 699 2556 703
rect 2550 698 2556 699
rect 2702 703 2708 704
rect 2702 699 2703 703
rect 2707 699 2708 703
rect 2702 698 2708 699
rect 2846 703 2852 704
rect 2846 699 2847 703
rect 2851 699 2852 703
rect 2846 698 2852 699
rect 2982 703 2988 704
rect 2982 699 2983 703
rect 2987 699 2988 703
rect 2982 698 2988 699
rect 3118 703 3124 704
rect 3118 699 3119 703
rect 3123 699 3124 703
rect 3118 698 3124 699
rect 3254 703 3260 704
rect 3254 699 3255 703
rect 3259 699 3260 703
rect 3254 698 3260 699
rect 3366 703 3372 704
rect 3366 699 3367 703
rect 3371 699 3372 703
rect 3462 700 3463 704
rect 3467 700 3468 704
rect 3462 699 3468 700
rect 3366 698 3372 699
rect 1766 695 1772 696
rect 1998 695 2004 696
rect 1502 694 1508 695
rect 274 691 280 692
rect 274 690 275 691
rect 241 688 275 690
rect 274 687 275 688
rect 279 687 280 691
rect 274 686 280 687
rect 366 691 372 692
rect 366 687 367 691
rect 371 687 372 691
rect 366 686 372 687
rect 502 691 508 692
rect 502 687 503 691
rect 507 687 508 691
rect 502 686 508 687
rect 646 691 652 692
rect 646 687 647 691
rect 651 687 652 691
rect 646 686 652 687
rect 654 691 660 692
rect 654 687 655 691
rect 659 690 660 691
rect 950 691 956 692
rect 659 688 769 690
rect 659 687 660 688
rect 654 686 660 687
rect 950 687 951 691
rect 955 687 956 691
rect 950 686 956 687
rect 1102 691 1108 692
rect 1102 687 1103 691
rect 1107 687 1108 691
rect 1262 691 1268 692
rect 1102 686 1108 687
rect 1254 687 1260 688
rect 110 683 116 684
rect 110 679 111 683
rect 115 679 116 683
rect 1254 683 1255 687
rect 1259 683 1260 687
rect 1262 687 1263 691
rect 1267 690 1268 691
rect 1422 691 1428 692
rect 1267 688 1385 690
rect 1267 687 1268 688
rect 1262 686 1268 687
rect 1422 687 1423 691
rect 1427 690 1428 691
rect 1998 691 1999 695
rect 2003 691 2004 695
rect 1998 690 2004 691
rect 2142 695 2148 696
rect 2142 691 2143 695
rect 2147 691 2148 695
rect 2142 690 2148 691
rect 2302 695 2308 696
rect 2302 691 2303 695
rect 2307 691 2308 695
rect 2302 690 2308 691
rect 2462 695 2468 696
rect 2462 691 2463 695
rect 2467 691 2468 695
rect 2462 690 2468 691
rect 2470 695 2476 696
rect 2470 691 2471 695
rect 2475 694 2476 695
rect 2694 695 2700 696
rect 2475 692 2593 694
rect 2475 691 2476 692
rect 2470 690 2476 691
rect 2694 691 2695 695
rect 2699 694 2700 695
rect 2794 695 2800 696
rect 2699 692 2745 694
rect 2699 691 2700 692
rect 2694 690 2700 691
rect 2794 691 2795 695
rect 2799 694 2800 695
rect 2927 695 2933 696
rect 2799 692 2889 694
rect 2799 691 2800 692
rect 2794 690 2800 691
rect 2927 691 2928 695
rect 2932 694 2933 695
rect 3190 695 3196 696
rect 2932 692 3025 694
rect 2932 691 2933 692
rect 2927 690 2933 691
rect 3190 691 3191 695
rect 3195 691 3196 695
rect 3190 690 3196 691
rect 3198 695 3204 696
rect 3198 691 3199 695
rect 3203 694 3204 695
rect 3203 692 3297 694
rect 3203 691 3204 692
rect 3198 690 3204 691
rect 3438 691 3444 692
rect 1427 688 1545 690
rect 1427 687 1428 688
rect 1422 686 1428 687
rect 1806 687 1812 688
rect 1254 682 1260 683
rect 1766 683 1772 684
rect 110 678 116 679
rect 166 680 172 681
rect 166 676 167 680
rect 171 676 172 680
rect 166 675 172 676
rect 294 680 300 681
rect 294 676 295 680
rect 299 676 300 680
rect 294 675 300 676
rect 430 680 436 681
rect 430 676 431 680
rect 435 676 436 680
rect 430 675 436 676
rect 574 680 580 681
rect 574 676 575 680
rect 579 676 580 680
rect 574 675 580 676
rect 726 680 732 681
rect 726 676 727 680
rect 731 676 732 680
rect 726 675 732 676
rect 878 680 884 681
rect 878 676 879 680
rect 883 676 884 680
rect 878 675 884 676
rect 1030 680 1036 681
rect 1030 676 1031 680
rect 1035 676 1036 680
rect 1030 675 1036 676
rect 1182 680 1188 681
rect 1182 676 1183 680
rect 1187 676 1188 680
rect 1182 675 1188 676
rect 1342 680 1348 681
rect 1342 676 1343 680
rect 1347 676 1348 680
rect 1342 675 1348 676
rect 1502 680 1508 681
rect 1502 676 1503 680
rect 1507 676 1508 680
rect 1766 679 1767 683
rect 1771 679 1772 683
rect 1806 683 1807 687
rect 1811 683 1812 687
rect 3438 687 3439 691
rect 3443 687 3444 691
rect 3438 686 3444 687
rect 3462 687 3468 688
rect 1806 682 1812 683
rect 1926 684 1932 685
rect 1926 680 1927 684
rect 1931 680 1932 684
rect 1926 679 1932 680
rect 2070 684 2076 685
rect 2070 680 2071 684
rect 2075 680 2076 684
rect 2070 679 2076 680
rect 2230 684 2236 685
rect 2230 680 2231 684
rect 2235 680 2236 684
rect 2230 679 2236 680
rect 2390 684 2396 685
rect 2390 680 2391 684
rect 2395 680 2396 684
rect 2390 679 2396 680
rect 2550 684 2556 685
rect 2550 680 2551 684
rect 2555 680 2556 684
rect 2550 679 2556 680
rect 2702 684 2708 685
rect 2702 680 2703 684
rect 2707 680 2708 684
rect 2702 679 2708 680
rect 2846 684 2852 685
rect 2846 680 2847 684
rect 2851 680 2852 684
rect 2846 679 2852 680
rect 2982 684 2988 685
rect 2982 680 2983 684
rect 2987 680 2988 684
rect 2982 679 2988 680
rect 3118 684 3124 685
rect 3118 680 3119 684
rect 3123 680 3124 684
rect 3118 679 3124 680
rect 3254 684 3260 685
rect 3254 680 3255 684
rect 3259 680 3260 684
rect 3254 679 3260 680
rect 3366 684 3372 685
rect 3366 680 3367 684
rect 3371 680 3372 684
rect 3462 683 3463 687
rect 3467 683 3468 687
rect 3462 682 3468 683
rect 3366 679 3372 680
rect 1766 678 1772 679
rect 1502 675 1508 676
rect 2114 675 2120 676
rect 2114 671 2115 675
rect 2119 674 2120 675
rect 2470 675 2476 676
rect 2470 674 2471 675
rect 2119 672 2471 674
rect 2119 671 2120 672
rect 2114 670 2120 671
rect 2470 671 2471 672
rect 2475 671 2476 675
rect 2470 670 2476 671
rect 1986 667 1992 668
rect 1986 663 1987 667
rect 1991 666 1992 667
rect 2398 667 2404 668
rect 2398 666 2399 667
rect 1991 664 2399 666
rect 1991 663 1992 664
rect 1986 662 1992 663
rect 2398 663 2399 664
rect 2403 663 2404 667
rect 2398 662 2404 663
rect 942 639 948 640
rect 942 635 943 639
rect 947 638 948 639
rect 1882 639 1888 640
rect 947 636 1014 638
rect 947 635 948 636
rect 942 634 948 635
rect 454 632 460 633
rect 110 629 116 630
rect 110 625 111 629
rect 115 625 116 629
rect 454 628 455 632
rect 459 628 460 632
rect 454 627 460 628
rect 558 632 564 633
rect 558 628 559 632
rect 563 628 564 632
rect 558 627 564 628
rect 678 632 684 633
rect 678 628 679 632
rect 683 628 684 632
rect 678 627 684 628
rect 798 632 804 633
rect 798 628 799 632
rect 803 628 804 632
rect 798 627 804 628
rect 926 632 932 633
rect 926 628 927 632
rect 931 628 932 632
rect 926 627 932 628
rect 110 624 116 625
rect 526 623 532 624
rect 526 619 527 623
rect 531 619 532 623
rect 526 618 532 619
rect 630 623 636 624
rect 630 619 631 623
rect 635 619 636 623
rect 630 618 636 619
rect 750 623 756 624
rect 750 619 751 623
rect 755 619 756 623
rect 750 618 756 619
rect 870 623 876 624
rect 870 619 871 623
rect 875 619 876 623
rect 870 618 876 619
rect 990 623 996 624
rect 990 619 991 623
rect 995 619 996 623
rect 1012 622 1014 636
rect 1882 635 1883 639
rect 1887 638 1888 639
rect 2238 639 2244 640
rect 2238 638 2239 639
rect 1887 636 2239 638
rect 1887 635 1888 636
rect 1882 634 1888 635
rect 2238 635 2239 636
rect 2243 635 2244 639
rect 2238 634 2244 635
rect 2506 639 2512 640
rect 2506 635 2507 639
rect 2511 638 2512 639
rect 2918 639 2924 640
rect 2918 638 2919 639
rect 2511 636 2919 638
rect 2511 635 2512 636
rect 2506 634 2512 635
rect 2918 635 2919 636
rect 2923 635 2924 639
rect 2918 634 2924 635
rect 1054 632 1060 633
rect 1054 628 1055 632
rect 1059 628 1060 632
rect 1054 627 1060 628
rect 1182 632 1188 633
rect 1182 628 1183 632
rect 1187 628 1188 632
rect 1182 627 1188 628
rect 1310 632 1316 633
rect 1310 628 1311 632
rect 1315 628 1316 632
rect 1310 627 1316 628
rect 1446 632 1452 633
rect 1446 628 1447 632
rect 1451 628 1452 632
rect 1446 627 1452 628
rect 1582 632 1588 633
rect 1582 628 1583 632
rect 1587 628 1588 632
rect 1830 632 1836 633
rect 1582 627 1588 628
rect 1766 629 1772 630
rect 1766 625 1767 629
rect 1771 625 1772 629
rect 1766 624 1772 625
rect 1806 629 1812 630
rect 1806 625 1807 629
rect 1811 625 1812 629
rect 1830 628 1831 632
rect 1835 628 1836 632
rect 1830 627 1836 628
rect 1966 632 1972 633
rect 1966 628 1967 632
rect 1971 628 1972 632
rect 1966 627 1972 628
rect 2134 632 2140 633
rect 2134 628 2135 632
rect 2139 628 2140 632
rect 2134 627 2140 628
rect 2310 632 2316 633
rect 2310 628 2311 632
rect 2315 628 2316 632
rect 2310 627 2316 628
rect 2486 632 2492 633
rect 2486 628 2487 632
rect 2491 628 2492 632
rect 2486 627 2492 628
rect 2654 632 2660 633
rect 2654 628 2655 632
rect 2659 628 2660 632
rect 2654 627 2660 628
rect 2814 632 2820 633
rect 2814 628 2815 632
rect 2819 628 2820 632
rect 2814 627 2820 628
rect 2958 632 2964 633
rect 2958 628 2959 632
rect 2963 628 2964 632
rect 2958 627 2964 628
rect 3102 632 3108 633
rect 3102 628 3103 632
rect 3107 628 3108 632
rect 3102 627 3108 628
rect 3246 632 3252 633
rect 3246 628 3247 632
rect 3251 628 3252 632
rect 3246 627 3252 628
rect 3366 632 3372 633
rect 3366 628 3367 632
rect 3371 628 3372 632
rect 3366 627 3372 628
rect 3462 629 3468 630
rect 1806 624 1812 625
rect 3462 625 3463 629
rect 3467 625 3468 629
rect 3462 624 3468 625
rect 1134 623 1140 624
rect 1012 620 1097 622
rect 990 618 996 619
rect 1134 619 1135 623
rect 1139 622 1140 623
rect 1382 623 1388 624
rect 1139 620 1225 622
rect 1139 619 1140 620
rect 1134 618 1140 619
rect 1382 619 1383 623
rect 1387 619 1388 623
rect 1382 618 1388 619
rect 1518 623 1524 624
rect 1518 619 1519 623
rect 1523 619 1524 623
rect 1518 618 1524 619
rect 1646 623 1652 624
rect 1646 619 1647 623
rect 1651 619 1652 623
rect 1646 618 1652 619
rect 1902 623 1908 624
rect 1902 619 1903 623
rect 1907 619 1908 623
rect 1902 618 1908 619
rect 2038 623 2044 624
rect 2038 619 2039 623
rect 2043 619 2044 623
rect 2038 618 2044 619
rect 2206 623 2212 624
rect 2206 619 2207 623
rect 2211 619 2212 623
rect 2206 618 2212 619
rect 2382 623 2388 624
rect 2382 619 2383 623
rect 2387 619 2388 623
rect 2382 618 2388 619
rect 2398 623 2404 624
rect 2398 619 2399 623
rect 2403 622 2404 623
rect 2726 623 2732 624
rect 2403 620 2529 622
rect 2403 619 2404 620
rect 2398 618 2404 619
rect 2726 619 2727 623
rect 2731 619 2732 623
rect 2726 618 2732 619
rect 2886 623 2892 624
rect 2886 619 2887 623
rect 2891 619 2892 623
rect 2886 618 2892 619
rect 3030 623 3036 624
rect 3030 619 3031 623
rect 3035 619 3036 623
rect 3030 618 3036 619
rect 3174 623 3180 624
rect 3174 619 3175 623
rect 3179 619 3180 623
rect 3174 618 3180 619
rect 3310 623 3316 624
rect 3310 619 3311 623
rect 3315 619 3316 623
rect 3310 618 3316 619
rect 3430 623 3436 624
rect 3430 619 3431 623
rect 3435 619 3436 623
rect 3430 618 3436 619
rect 454 613 460 614
rect 110 612 116 613
rect 110 608 111 612
rect 115 608 116 612
rect 454 609 455 613
rect 459 609 460 613
rect 454 608 460 609
rect 558 613 564 614
rect 558 609 559 613
rect 563 609 564 613
rect 558 608 564 609
rect 678 613 684 614
rect 678 609 679 613
rect 683 609 684 613
rect 678 608 684 609
rect 798 613 804 614
rect 798 609 799 613
rect 803 609 804 613
rect 798 608 804 609
rect 926 613 932 614
rect 926 609 927 613
rect 931 609 932 613
rect 926 608 932 609
rect 1054 613 1060 614
rect 1054 609 1055 613
rect 1059 609 1060 613
rect 1054 608 1060 609
rect 1182 613 1188 614
rect 1182 609 1183 613
rect 1187 609 1188 613
rect 1182 608 1188 609
rect 1310 613 1316 614
rect 1310 609 1311 613
rect 1315 609 1316 613
rect 1310 608 1316 609
rect 1446 613 1452 614
rect 1446 609 1447 613
rect 1451 609 1452 613
rect 1446 608 1452 609
rect 1582 613 1588 614
rect 1830 613 1836 614
rect 1582 609 1583 613
rect 1587 609 1588 613
rect 1582 608 1588 609
rect 1766 612 1772 613
rect 1766 608 1767 612
rect 1771 608 1772 612
rect 110 607 116 608
rect 1766 607 1772 608
rect 1806 612 1812 613
rect 1806 608 1807 612
rect 1811 608 1812 612
rect 1830 609 1831 613
rect 1835 609 1836 613
rect 1830 608 1836 609
rect 1966 613 1972 614
rect 1966 609 1967 613
rect 1971 609 1972 613
rect 1966 608 1972 609
rect 2134 613 2140 614
rect 2134 609 2135 613
rect 2139 609 2140 613
rect 2134 608 2140 609
rect 2310 613 2316 614
rect 2310 609 2311 613
rect 2315 609 2316 613
rect 2310 608 2316 609
rect 2486 613 2492 614
rect 2486 609 2487 613
rect 2491 609 2492 613
rect 2486 608 2492 609
rect 2654 613 2660 614
rect 2654 609 2655 613
rect 2659 609 2660 613
rect 2654 608 2660 609
rect 2814 613 2820 614
rect 2814 609 2815 613
rect 2819 609 2820 613
rect 2814 608 2820 609
rect 2958 613 2964 614
rect 2958 609 2959 613
rect 2963 609 2964 613
rect 2958 608 2964 609
rect 3102 613 3108 614
rect 3102 609 3103 613
rect 3107 609 3108 613
rect 3102 608 3108 609
rect 3246 613 3252 614
rect 3246 609 3247 613
rect 3251 609 3252 613
rect 3246 608 3252 609
rect 3366 613 3372 614
rect 3366 609 3367 613
rect 3371 609 3372 613
rect 3366 608 3372 609
rect 3462 612 3468 613
rect 3462 608 3463 612
rect 3467 608 3468 612
rect 1806 607 1812 608
rect 3462 607 3468 608
rect 503 595 509 596
rect 503 591 504 595
rect 508 594 509 595
rect 526 595 532 596
rect 508 592 522 594
rect 508 591 509 592
rect 503 590 509 591
rect 520 586 522 592
rect 526 591 527 595
rect 531 594 532 595
rect 607 595 613 596
rect 607 594 608 595
rect 531 592 608 594
rect 531 591 532 592
rect 526 590 532 591
rect 607 591 608 592
rect 612 591 613 595
rect 607 590 613 591
rect 630 595 636 596
rect 630 591 631 595
rect 635 594 636 595
rect 727 595 733 596
rect 727 594 728 595
rect 635 592 728 594
rect 635 591 636 592
rect 630 590 636 591
rect 727 591 728 592
rect 732 591 733 595
rect 727 590 733 591
rect 750 595 756 596
rect 750 591 751 595
rect 755 594 756 595
rect 847 595 853 596
rect 847 594 848 595
rect 755 592 848 594
rect 755 591 756 592
rect 750 590 756 591
rect 847 591 848 592
rect 852 591 853 595
rect 847 590 853 591
rect 870 595 876 596
rect 870 591 871 595
rect 875 594 876 595
rect 975 595 981 596
rect 975 594 976 595
rect 875 592 976 594
rect 875 591 876 592
rect 870 590 876 591
rect 975 591 976 592
rect 980 591 981 595
rect 975 590 981 591
rect 1103 595 1109 596
rect 1103 591 1104 595
rect 1108 594 1109 595
rect 1134 595 1140 596
rect 1134 594 1135 595
rect 1108 592 1135 594
rect 1108 591 1109 592
rect 1103 590 1109 591
rect 1134 591 1135 592
rect 1139 591 1140 595
rect 1134 590 1140 591
rect 1231 595 1237 596
rect 1231 591 1232 595
rect 1236 594 1237 595
rect 1239 595 1245 596
rect 1239 594 1240 595
rect 1236 592 1240 594
rect 1236 591 1237 592
rect 1231 590 1237 591
rect 1239 591 1240 592
rect 1244 591 1245 595
rect 1239 590 1245 591
rect 1254 595 1260 596
rect 1254 591 1255 595
rect 1259 594 1260 595
rect 1359 595 1365 596
rect 1359 594 1360 595
rect 1259 592 1360 594
rect 1259 591 1260 592
rect 1254 590 1260 591
rect 1359 591 1360 592
rect 1364 591 1365 595
rect 1359 590 1365 591
rect 1382 595 1388 596
rect 1382 591 1383 595
rect 1387 594 1388 595
rect 1495 595 1501 596
rect 1495 594 1496 595
rect 1387 592 1496 594
rect 1387 591 1388 592
rect 1382 590 1388 591
rect 1495 591 1496 592
rect 1500 591 1501 595
rect 1495 590 1501 591
rect 1518 595 1524 596
rect 1518 591 1519 595
rect 1523 594 1524 595
rect 1631 595 1637 596
rect 1631 594 1632 595
rect 1523 592 1632 594
rect 1523 591 1524 592
rect 1518 590 1524 591
rect 1631 591 1632 592
rect 1636 591 1637 595
rect 1631 590 1637 591
rect 1879 595 1888 596
rect 1879 591 1880 595
rect 1887 591 1888 595
rect 1879 590 1888 591
rect 1902 595 1908 596
rect 1902 591 1903 595
rect 1907 594 1908 595
rect 2015 595 2021 596
rect 2015 594 2016 595
rect 1907 592 2016 594
rect 1907 591 1908 592
rect 1902 590 1908 591
rect 2015 591 2016 592
rect 2020 591 2021 595
rect 2015 590 2021 591
rect 2038 595 2044 596
rect 2038 591 2039 595
rect 2043 594 2044 595
rect 2183 595 2189 596
rect 2183 594 2184 595
rect 2043 592 2184 594
rect 2043 591 2044 592
rect 2038 590 2044 591
rect 2183 591 2184 592
rect 2188 591 2189 595
rect 2183 590 2189 591
rect 2206 595 2212 596
rect 2206 591 2207 595
rect 2211 594 2212 595
rect 2359 595 2365 596
rect 2359 594 2360 595
rect 2211 592 2360 594
rect 2211 591 2212 592
rect 2206 590 2212 591
rect 2359 591 2360 592
rect 2364 591 2365 595
rect 2359 590 2365 591
rect 2382 595 2388 596
rect 2382 591 2383 595
rect 2387 594 2388 595
rect 2535 595 2541 596
rect 2535 594 2536 595
rect 2387 592 2536 594
rect 2387 591 2388 592
rect 2382 590 2388 591
rect 2535 591 2536 592
rect 2540 591 2541 595
rect 2535 590 2541 591
rect 2694 595 2700 596
rect 2694 591 2695 595
rect 2699 594 2700 595
rect 2703 595 2709 596
rect 2703 594 2704 595
rect 2699 592 2704 594
rect 2699 591 2700 592
rect 2694 590 2700 591
rect 2703 591 2704 592
rect 2708 591 2709 595
rect 2703 590 2709 591
rect 2726 595 2732 596
rect 2726 591 2727 595
rect 2731 594 2732 595
rect 2863 595 2869 596
rect 2863 594 2864 595
rect 2731 592 2864 594
rect 2731 591 2732 592
rect 2726 590 2732 591
rect 2863 591 2864 592
rect 2868 591 2869 595
rect 2863 590 2869 591
rect 2886 595 2892 596
rect 2886 591 2887 595
rect 2891 594 2892 595
rect 3007 595 3013 596
rect 3007 594 3008 595
rect 2891 592 3008 594
rect 2891 591 2892 592
rect 2886 590 2892 591
rect 3007 591 3008 592
rect 3012 591 3013 595
rect 3007 590 3013 591
rect 3030 595 3036 596
rect 3030 591 3031 595
rect 3035 594 3036 595
rect 3151 595 3157 596
rect 3151 594 3152 595
rect 3035 592 3152 594
rect 3035 591 3036 592
rect 3030 590 3036 591
rect 3151 591 3152 592
rect 3156 591 3157 595
rect 3151 590 3157 591
rect 3295 595 3301 596
rect 3295 591 3296 595
rect 3300 594 3301 595
rect 3318 595 3324 596
rect 3318 594 3319 595
rect 3300 592 3319 594
rect 3300 591 3301 592
rect 3295 590 3301 591
rect 3318 591 3319 592
rect 3323 591 3324 595
rect 3318 590 3324 591
rect 3415 595 3421 596
rect 3415 591 3416 595
rect 3420 594 3421 595
rect 3438 595 3444 596
rect 3438 594 3439 595
rect 3420 592 3439 594
rect 3420 591 3421 592
rect 3415 590 3421 591
rect 3438 591 3439 592
rect 3443 591 3444 595
rect 3438 590 3444 591
rect 654 587 660 588
rect 654 586 655 587
rect 520 584 655 586
rect 654 583 655 584
rect 659 583 660 587
rect 654 582 660 583
rect 1006 583 1012 584
rect 1006 582 1007 583
rect 664 580 1007 582
rect 647 575 653 576
rect 647 571 648 575
rect 652 574 653 575
rect 664 574 666 580
rect 1006 579 1007 580
rect 1011 579 1012 583
rect 1006 578 1012 579
rect 1742 583 1748 584
rect 1742 579 1743 583
rect 1747 582 1748 583
rect 1879 583 1885 584
rect 1879 582 1880 583
rect 1747 580 1880 582
rect 1747 579 1748 580
rect 1742 578 1748 579
rect 1879 579 1880 580
rect 1884 579 1885 583
rect 1879 578 1885 579
rect 1902 583 1908 584
rect 1902 579 1903 583
rect 1907 582 1908 583
rect 2015 583 2021 584
rect 2015 582 2016 583
rect 1907 580 2016 582
rect 1907 579 1908 580
rect 1902 578 1908 579
rect 2015 579 2016 580
rect 2020 579 2021 583
rect 2015 578 2021 579
rect 2038 583 2044 584
rect 2038 579 2039 583
rect 2043 582 2044 583
rect 2175 583 2181 584
rect 2175 582 2176 583
rect 2043 580 2176 582
rect 2043 579 2044 580
rect 2038 578 2044 579
rect 2175 579 2176 580
rect 2180 579 2181 583
rect 2175 578 2181 579
rect 2198 583 2204 584
rect 2198 579 2199 583
rect 2203 582 2204 583
rect 2335 583 2341 584
rect 2335 582 2336 583
rect 2203 580 2336 582
rect 2203 579 2204 580
rect 2198 578 2204 579
rect 2335 579 2336 580
rect 2340 579 2341 583
rect 2335 578 2341 579
rect 2503 583 2512 584
rect 2503 579 2504 583
rect 2511 579 2512 583
rect 2503 578 2512 579
rect 2526 583 2532 584
rect 2526 579 2527 583
rect 2531 582 2532 583
rect 2671 583 2677 584
rect 2671 582 2672 583
rect 2531 580 2672 582
rect 2531 579 2532 580
rect 2526 578 2532 579
rect 2671 579 2672 580
rect 2676 579 2677 583
rect 2671 578 2677 579
rect 2694 583 2700 584
rect 2694 579 2695 583
rect 2699 582 2700 583
rect 2847 583 2853 584
rect 2847 582 2848 583
rect 2699 580 2848 582
rect 2699 579 2700 580
rect 2694 578 2700 579
rect 2847 579 2848 580
rect 2852 579 2853 583
rect 2847 578 2853 579
rect 3031 583 3037 584
rect 3031 579 3032 583
rect 3036 582 3037 583
rect 3062 583 3068 584
rect 3062 582 3063 583
rect 3036 580 3063 582
rect 3036 579 3037 580
rect 3031 578 3037 579
rect 3062 579 3063 580
rect 3067 579 3068 583
rect 3062 578 3068 579
rect 3174 583 3180 584
rect 3174 579 3175 583
rect 3179 582 3180 583
rect 3215 583 3221 584
rect 3215 582 3216 583
rect 3179 580 3216 582
rect 3179 579 3180 580
rect 3174 578 3180 579
rect 3215 579 3216 580
rect 3220 579 3221 583
rect 3215 578 3221 579
rect 3407 583 3413 584
rect 3407 579 3408 583
rect 3412 582 3413 583
rect 3430 583 3436 584
rect 3430 582 3431 583
rect 3412 580 3431 582
rect 3412 579 3413 580
rect 3407 578 3413 579
rect 3430 579 3431 580
rect 3435 579 3436 583
rect 3430 578 3436 579
rect 652 572 666 574
rect 670 575 676 576
rect 652 571 653 572
rect 647 570 653 571
rect 670 571 671 575
rect 675 574 676 575
rect 751 575 757 576
rect 751 574 752 575
rect 675 572 752 574
rect 675 571 676 572
rect 670 570 676 571
rect 751 571 752 572
rect 756 571 757 575
rect 751 570 757 571
rect 774 575 780 576
rect 774 571 775 575
rect 779 574 780 575
rect 863 575 869 576
rect 863 574 864 575
rect 779 572 864 574
rect 779 571 780 572
rect 774 570 780 571
rect 863 571 864 572
rect 868 571 869 575
rect 863 570 869 571
rect 975 575 981 576
rect 975 571 976 575
rect 980 574 981 575
rect 990 575 996 576
rect 990 574 991 575
rect 980 572 991 574
rect 980 571 981 572
rect 975 570 981 571
rect 990 571 991 572
rect 995 571 996 575
rect 990 570 996 571
rect 998 575 1004 576
rect 998 571 999 575
rect 1003 574 1004 575
rect 1087 575 1093 576
rect 1087 574 1088 575
rect 1003 572 1088 574
rect 1003 571 1004 572
rect 998 570 1004 571
rect 1087 571 1088 572
rect 1092 571 1093 575
rect 1087 570 1093 571
rect 1198 575 1205 576
rect 1198 571 1199 575
rect 1204 571 1205 575
rect 1198 570 1205 571
rect 1222 575 1228 576
rect 1222 571 1223 575
rect 1227 574 1228 575
rect 1303 575 1309 576
rect 1303 574 1304 575
rect 1227 572 1304 574
rect 1227 571 1228 572
rect 1222 570 1228 571
rect 1303 571 1304 572
rect 1308 571 1309 575
rect 1303 570 1309 571
rect 1407 575 1413 576
rect 1407 571 1408 575
rect 1412 574 1413 575
rect 1438 575 1444 576
rect 1438 574 1439 575
rect 1412 572 1439 574
rect 1412 571 1413 572
rect 1407 570 1413 571
rect 1438 571 1439 572
rect 1443 571 1444 575
rect 1438 570 1444 571
rect 1519 575 1525 576
rect 1519 571 1520 575
rect 1524 574 1525 575
rect 1550 575 1556 576
rect 1550 574 1551 575
rect 1524 572 1551 574
rect 1524 571 1525 572
rect 1519 570 1525 571
rect 1550 571 1551 572
rect 1555 571 1556 575
rect 1550 570 1556 571
rect 1631 575 1637 576
rect 1631 571 1632 575
rect 1636 574 1637 575
rect 1646 575 1652 576
rect 1646 574 1647 575
rect 1636 572 1647 574
rect 1636 571 1637 572
rect 1631 570 1637 571
rect 1646 571 1647 572
rect 1651 571 1652 575
rect 1646 570 1652 571
rect 1719 575 1725 576
rect 1719 571 1720 575
rect 1724 574 1725 575
rect 1734 575 1740 576
rect 1734 574 1735 575
rect 1724 572 1735 574
rect 1724 571 1725 572
rect 1719 570 1725 571
rect 1734 571 1735 572
rect 1739 571 1740 575
rect 1734 570 1740 571
rect 1806 568 1812 569
rect 3462 568 3468 569
rect 1806 564 1807 568
rect 1811 564 1812 568
rect 1806 563 1812 564
rect 1830 567 1836 568
rect 1830 563 1831 567
rect 1835 563 1836 567
rect 1830 562 1836 563
rect 1966 567 1972 568
rect 1966 563 1967 567
rect 1971 563 1972 567
rect 1966 562 1972 563
rect 2126 567 2132 568
rect 2126 563 2127 567
rect 2131 563 2132 567
rect 2126 562 2132 563
rect 2286 567 2292 568
rect 2286 563 2287 567
rect 2291 563 2292 567
rect 2286 562 2292 563
rect 2454 567 2460 568
rect 2454 563 2455 567
rect 2459 563 2460 567
rect 2454 562 2460 563
rect 2622 567 2628 568
rect 2622 563 2623 567
rect 2627 563 2628 567
rect 2622 562 2628 563
rect 2798 567 2804 568
rect 2798 563 2799 567
rect 2803 563 2804 567
rect 2798 562 2804 563
rect 2982 567 2988 568
rect 2982 563 2983 567
rect 2987 563 2988 567
rect 2982 562 2988 563
rect 3166 567 3172 568
rect 3166 563 3167 567
rect 3171 563 3172 567
rect 3166 562 3172 563
rect 3358 567 3364 568
rect 3358 563 3359 567
rect 3363 563 3364 567
rect 3462 564 3463 568
rect 3467 564 3468 568
rect 3462 563 3468 564
rect 3358 562 3364 563
rect 110 560 116 561
rect 1766 560 1772 561
rect 110 556 111 560
rect 115 556 116 560
rect 110 555 116 556
rect 598 559 604 560
rect 598 555 599 559
rect 603 555 604 559
rect 598 554 604 555
rect 702 559 708 560
rect 702 555 703 559
rect 707 555 708 559
rect 702 554 708 555
rect 814 559 820 560
rect 814 555 815 559
rect 819 555 820 559
rect 814 554 820 555
rect 926 559 932 560
rect 926 555 927 559
rect 931 555 932 559
rect 926 554 932 555
rect 1038 559 1044 560
rect 1038 555 1039 559
rect 1043 555 1044 559
rect 1038 554 1044 555
rect 1150 559 1156 560
rect 1150 555 1151 559
rect 1155 555 1156 559
rect 1150 554 1156 555
rect 1254 559 1260 560
rect 1254 555 1255 559
rect 1259 555 1260 559
rect 1254 554 1260 555
rect 1358 559 1364 560
rect 1358 555 1359 559
rect 1363 555 1364 559
rect 1358 554 1364 555
rect 1470 559 1476 560
rect 1470 555 1471 559
rect 1475 555 1476 559
rect 1470 554 1476 555
rect 1582 559 1588 560
rect 1582 555 1583 559
rect 1587 555 1588 559
rect 1582 554 1588 555
rect 1670 559 1676 560
rect 1670 555 1671 559
rect 1675 555 1676 559
rect 1766 556 1767 560
rect 1771 556 1772 560
rect 1766 555 1772 556
rect 1902 559 1908 560
rect 1902 555 1903 559
rect 1907 555 1908 559
rect 1670 554 1676 555
rect 1902 554 1908 555
rect 2038 559 2044 560
rect 2038 555 2039 559
rect 2043 555 2044 559
rect 2038 554 2044 555
rect 2198 559 2204 560
rect 2198 555 2199 559
rect 2203 555 2204 559
rect 2198 554 2204 555
rect 2238 559 2244 560
rect 2238 555 2239 559
rect 2243 558 2244 559
rect 2526 559 2532 560
rect 2243 556 2329 558
rect 2243 555 2244 556
rect 2238 554 2244 555
rect 2526 555 2527 559
rect 2531 555 2532 559
rect 2526 554 2532 555
rect 2694 559 2700 560
rect 2694 555 2695 559
rect 2699 555 2700 559
rect 2918 559 2924 560
rect 2694 554 2700 555
rect 2878 555 2884 556
rect 2878 554 2879 555
rect 2873 552 2879 554
rect 670 551 676 552
rect 670 547 671 551
rect 675 547 676 551
rect 670 546 676 547
rect 774 551 780 552
rect 774 547 775 551
rect 779 547 780 551
rect 998 551 1004 552
rect 774 546 780 547
rect 886 547 892 548
rect 110 543 116 544
rect 110 539 111 543
rect 115 539 116 543
rect 886 543 887 547
rect 891 543 892 547
rect 998 547 999 551
rect 1003 547 1004 551
rect 998 546 1004 547
rect 1006 551 1012 552
rect 1006 547 1007 551
rect 1011 550 1012 551
rect 1222 551 1228 552
rect 1011 548 1081 550
rect 1011 547 1012 548
rect 1006 546 1012 547
rect 1222 547 1223 551
rect 1227 547 1228 551
rect 1222 546 1228 547
rect 1239 551 1245 552
rect 1239 547 1240 551
rect 1244 550 1245 551
rect 1438 551 1444 552
rect 1244 548 1297 550
rect 1244 547 1245 548
rect 1239 546 1245 547
rect 1438 547 1439 551
rect 1443 550 1444 551
rect 1550 551 1556 552
rect 1443 548 1513 550
rect 1443 547 1444 548
rect 1438 546 1444 547
rect 1550 547 1551 551
rect 1555 550 1556 551
rect 1742 551 1748 552
rect 1555 548 1625 550
rect 1555 547 1556 548
rect 1550 546 1556 547
rect 1742 547 1743 551
rect 1747 547 1748 551
rect 1742 546 1748 547
rect 1806 551 1812 552
rect 1806 547 1807 551
rect 1811 547 1812 551
rect 2878 551 2879 552
rect 2883 551 2884 555
rect 2918 555 2919 559
rect 2923 558 2924 559
rect 3062 559 3068 560
rect 2923 556 3025 558
rect 2923 555 2924 556
rect 2918 554 2924 555
rect 3062 555 3063 559
rect 3067 558 3068 559
rect 3067 556 3209 558
rect 3067 555 3068 556
rect 3062 554 3068 555
rect 3430 555 3436 556
rect 2878 550 2884 551
rect 3430 551 3431 555
rect 3435 551 3436 555
rect 3430 550 3436 551
rect 3462 551 3468 552
rect 1806 546 1812 547
rect 1830 548 1836 549
rect 886 542 892 543
rect 1432 542 1434 545
rect 1830 544 1831 548
rect 1835 544 1836 548
rect 1455 543 1461 544
rect 1455 542 1456 543
rect 110 538 116 539
rect 598 540 604 541
rect 598 536 599 540
rect 603 536 604 540
rect 598 535 604 536
rect 702 540 708 541
rect 702 536 703 540
rect 707 536 708 540
rect 702 535 708 536
rect 814 540 820 541
rect 814 536 815 540
rect 819 536 820 540
rect 814 535 820 536
rect 926 540 932 541
rect 926 536 927 540
rect 931 536 932 540
rect 926 535 932 536
rect 1038 540 1044 541
rect 1038 536 1039 540
rect 1043 536 1044 540
rect 1038 535 1044 536
rect 1150 540 1156 541
rect 1150 536 1151 540
rect 1155 536 1156 540
rect 1150 535 1156 536
rect 1254 540 1260 541
rect 1254 536 1255 540
rect 1259 536 1260 540
rect 1254 535 1260 536
rect 1358 540 1364 541
rect 1432 540 1456 542
rect 1358 536 1359 540
rect 1363 536 1364 540
rect 1455 539 1456 540
rect 1460 539 1461 543
rect 1766 543 1772 544
rect 1830 543 1836 544
rect 1966 548 1972 549
rect 1966 544 1967 548
rect 1971 544 1972 548
rect 1966 543 1972 544
rect 2126 548 2132 549
rect 2126 544 2127 548
rect 2131 544 2132 548
rect 2126 543 2132 544
rect 2286 548 2292 549
rect 2286 544 2287 548
rect 2291 544 2292 548
rect 2286 543 2292 544
rect 2454 548 2460 549
rect 2454 544 2455 548
rect 2459 544 2460 548
rect 2454 543 2460 544
rect 2622 548 2628 549
rect 2622 544 2623 548
rect 2627 544 2628 548
rect 2622 543 2628 544
rect 2798 548 2804 549
rect 2798 544 2799 548
rect 2803 544 2804 548
rect 2798 543 2804 544
rect 2982 548 2988 549
rect 2982 544 2983 548
rect 2987 544 2988 548
rect 2982 543 2988 544
rect 3166 548 3172 549
rect 3166 544 3167 548
rect 3171 544 3172 548
rect 3166 543 3172 544
rect 3358 548 3364 549
rect 3358 544 3359 548
rect 3363 544 3364 548
rect 3462 547 3463 551
rect 3467 547 3468 551
rect 3462 546 3468 547
rect 3358 543 3364 544
rect 1455 538 1461 539
rect 1470 540 1476 541
rect 1358 535 1364 536
rect 1470 536 1471 540
rect 1475 536 1476 540
rect 1470 535 1476 536
rect 1582 540 1588 541
rect 1582 536 1583 540
rect 1587 536 1588 540
rect 1582 535 1588 536
rect 1670 540 1676 541
rect 1670 536 1671 540
rect 1675 536 1676 540
rect 1766 539 1767 543
rect 1771 539 1772 543
rect 1766 538 1772 539
rect 1670 535 1676 536
rect 302 496 308 497
rect 110 493 116 494
rect 110 489 111 493
rect 115 489 116 493
rect 302 492 303 496
rect 307 492 308 496
rect 302 491 308 492
rect 430 496 436 497
rect 430 492 431 496
rect 435 492 436 496
rect 430 491 436 492
rect 566 496 572 497
rect 566 492 567 496
rect 571 492 572 496
rect 566 491 572 492
rect 702 496 708 497
rect 702 492 703 496
rect 707 492 708 496
rect 702 491 708 492
rect 846 496 852 497
rect 846 492 847 496
rect 851 492 852 496
rect 846 491 852 492
rect 982 496 988 497
rect 982 492 983 496
rect 987 492 988 496
rect 982 491 988 492
rect 1110 496 1116 497
rect 1110 492 1111 496
rect 1115 492 1116 496
rect 1110 491 1116 492
rect 1230 496 1236 497
rect 1230 492 1231 496
rect 1235 492 1236 496
rect 1230 491 1236 492
rect 1350 496 1356 497
rect 1350 492 1351 496
rect 1355 492 1356 496
rect 1350 491 1356 492
rect 1462 496 1468 497
rect 1462 492 1463 496
rect 1467 492 1468 496
rect 1462 491 1468 492
rect 1574 496 1580 497
rect 1574 492 1575 496
rect 1579 492 1580 496
rect 1574 491 1580 492
rect 1670 496 1676 497
rect 1670 492 1671 496
rect 1675 492 1676 496
rect 1882 495 1888 496
rect 1670 491 1676 492
rect 1766 493 1772 494
rect 110 488 116 489
rect 1766 489 1767 493
rect 1771 489 1772 493
rect 1882 491 1883 495
rect 1887 494 1888 495
rect 2730 495 2736 496
rect 1887 492 2066 494
rect 1887 491 1888 492
rect 1882 490 1888 491
rect 1766 488 1772 489
rect 1830 488 1836 489
rect 374 487 380 488
rect 374 483 375 487
rect 379 483 380 487
rect 374 482 380 483
rect 502 487 508 488
rect 502 483 503 487
rect 507 483 508 487
rect 502 482 508 483
rect 630 487 636 488
rect 630 483 631 487
rect 635 483 636 487
rect 630 482 636 483
rect 646 487 652 488
rect 646 483 647 487
rect 651 486 652 487
rect 782 487 788 488
rect 651 484 745 486
rect 651 483 652 484
rect 646 482 652 483
rect 782 483 783 487
rect 787 486 788 487
rect 1054 487 1060 488
rect 787 484 889 486
rect 787 483 788 484
rect 782 482 788 483
rect 1054 483 1055 487
rect 1059 483 1060 487
rect 1198 487 1204 488
rect 1198 486 1199 487
rect 1185 484 1199 486
rect 1054 482 1060 483
rect 1198 483 1199 484
rect 1203 483 1204 487
rect 1198 482 1204 483
rect 1302 487 1308 488
rect 1302 483 1303 487
rect 1307 483 1308 487
rect 1302 482 1308 483
rect 1310 487 1316 488
rect 1310 483 1311 487
rect 1315 486 1316 487
rect 1430 487 1436 488
rect 1315 484 1393 486
rect 1315 483 1316 484
rect 1310 482 1316 483
rect 1430 483 1431 487
rect 1435 486 1436 487
rect 1734 487 1740 488
rect 1435 484 1505 486
rect 1435 483 1436 484
rect 1430 482 1436 483
rect 1734 483 1735 487
rect 1739 483 1740 487
rect 1734 482 1740 483
rect 1806 485 1812 486
rect 1806 481 1807 485
rect 1811 481 1812 485
rect 1830 484 1831 488
rect 1835 484 1836 488
rect 1830 483 1836 484
rect 1966 488 1972 489
rect 1966 484 1967 488
rect 1971 484 1972 488
rect 1966 483 1972 484
rect 1806 480 1812 481
rect 1647 479 1653 480
rect 302 477 308 478
rect 110 476 116 477
rect 110 472 111 476
rect 115 472 116 476
rect 302 473 303 477
rect 307 473 308 477
rect 302 472 308 473
rect 430 477 436 478
rect 430 473 431 477
rect 435 473 436 477
rect 430 472 436 473
rect 566 477 572 478
rect 566 473 567 477
rect 571 473 572 477
rect 566 472 572 473
rect 702 477 708 478
rect 702 473 703 477
rect 707 473 708 477
rect 702 472 708 473
rect 846 477 852 478
rect 846 473 847 477
rect 851 473 852 477
rect 846 472 852 473
rect 982 477 988 478
rect 982 473 983 477
rect 987 473 988 477
rect 982 472 988 473
rect 1110 477 1116 478
rect 1110 473 1111 477
rect 1115 473 1116 477
rect 1110 472 1116 473
rect 1230 477 1236 478
rect 1230 473 1231 477
rect 1235 473 1236 477
rect 1230 472 1236 473
rect 1350 477 1356 478
rect 1350 473 1351 477
rect 1355 473 1356 477
rect 1350 472 1356 473
rect 1462 477 1468 478
rect 1462 473 1463 477
rect 1467 473 1468 477
rect 1462 472 1468 473
rect 1574 477 1580 478
rect 1574 473 1575 477
rect 1579 473 1580 477
rect 1647 475 1648 479
rect 1652 478 1653 479
rect 1774 479 1780 480
rect 1652 476 1662 478
rect 1652 475 1653 476
rect 1647 474 1653 475
rect 1574 472 1580 473
rect 110 471 116 472
rect 1660 462 1662 476
rect 1670 477 1676 478
rect 1670 473 1671 477
rect 1675 473 1676 477
rect 1670 472 1676 473
rect 1766 476 1772 477
rect 1766 472 1767 476
rect 1771 472 1772 476
rect 1774 475 1775 479
rect 1779 478 1780 479
rect 2038 479 2044 480
rect 1779 476 1873 478
rect 1779 475 1780 476
rect 1774 474 1780 475
rect 2038 475 2039 479
rect 2043 475 2044 479
rect 2064 478 2066 492
rect 2730 491 2731 495
rect 2735 494 2736 495
rect 2735 492 2998 494
rect 2735 491 2736 492
rect 2730 490 2736 491
rect 2126 488 2132 489
rect 2126 484 2127 488
rect 2131 484 2132 488
rect 2126 483 2132 484
rect 2294 488 2300 489
rect 2294 484 2295 488
rect 2299 484 2300 488
rect 2294 483 2300 484
rect 2478 488 2484 489
rect 2478 484 2479 488
rect 2483 484 2484 488
rect 2478 483 2484 484
rect 2678 488 2684 489
rect 2678 484 2679 488
rect 2683 484 2684 488
rect 2678 483 2684 484
rect 2886 488 2892 489
rect 2886 484 2887 488
rect 2891 484 2892 488
rect 2886 483 2892 484
rect 2358 479 2364 480
rect 2064 476 2169 478
rect 2038 474 2044 475
rect 2358 475 2359 479
rect 2363 475 2364 479
rect 2358 474 2364 475
rect 2374 479 2380 480
rect 2374 475 2375 479
rect 2379 478 2380 479
rect 2558 479 2564 480
rect 2379 476 2521 478
rect 2379 475 2380 476
rect 2374 474 2380 475
rect 2558 475 2559 479
rect 2563 478 2564 479
rect 2958 479 2964 480
rect 2563 476 2721 478
rect 2563 475 2564 476
rect 2558 474 2564 475
rect 2958 475 2959 479
rect 2963 475 2964 479
rect 2996 478 2998 492
rect 3110 488 3116 489
rect 3110 484 3111 488
rect 3115 484 3116 488
rect 3110 483 3116 484
rect 3334 488 3340 489
rect 3334 484 3335 488
rect 3339 484 3340 488
rect 3334 483 3340 484
rect 3462 485 3468 486
rect 3462 481 3463 485
rect 3467 481 3468 485
rect 3462 480 3468 481
rect 3318 479 3324 480
rect 2996 476 3153 478
rect 2958 474 2964 475
rect 3318 475 3319 479
rect 3323 478 3324 479
rect 3323 476 3377 478
rect 3323 475 3324 476
rect 3318 474 3324 475
rect 1766 471 1772 472
rect 1830 469 1836 470
rect 1806 468 1812 469
rect 1806 464 1807 468
rect 1811 464 1812 468
rect 1830 465 1831 469
rect 1835 465 1836 469
rect 1830 464 1836 465
rect 1966 469 1972 470
rect 1966 465 1967 469
rect 1971 465 1972 469
rect 1966 464 1972 465
rect 2126 469 2132 470
rect 2126 465 2127 469
rect 2131 465 2132 469
rect 2126 464 2132 465
rect 2294 469 2300 470
rect 2294 465 2295 469
rect 2299 465 2300 469
rect 2294 464 2300 465
rect 2478 469 2484 470
rect 2478 465 2479 469
rect 2483 465 2484 469
rect 2478 464 2484 465
rect 2678 469 2684 470
rect 2678 465 2679 469
rect 2683 465 2684 469
rect 2678 464 2684 465
rect 2886 469 2892 470
rect 2886 465 2887 469
rect 2891 465 2892 469
rect 2886 464 2892 465
rect 3110 469 3116 470
rect 3110 465 3111 469
rect 3115 465 3116 469
rect 3110 464 3116 465
rect 3334 469 3340 470
rect 3334 465 3335 469
rect 3339 465 3340 469
rect 3334 464 3340 465
rect 3462 468 3468 469
rect 3462 464 3463 468
rect 3467 464 3468 468
rect 1806 463 1812 464
rect 3462 463 3468 464
rect 1660 460 1722 462
rect 351 459 357 460
rect 351 455 352 459
rect 356 458 357 459
rect 374 459 380 460
rect 356 456 370 458
rect 356 455 357 456
rect 351 454 357 455
rect 368 450 370 456
rect 374 455 375 459
rect 379 458 380 459
rect 479 459 485 460
rect 479 458 480 459
rect 379 456 480 458
rect 379 455 380 456
rect 374 454 380 455
rect 479 455 480 456
rect 484 455 485 459
rect 479 454 485 455
rect 502 459 508 460
rect 502 455 503 459
rect 507 458 508 459
rect 615 459 621 460
rect 615 458 616 459
rect 507 456 616 458
rect 507 455 508 456
rect 502 454 508 455
rect 615 455 616 456
rect 620 455 621 459
rect 751 459 757 460
rect 615 454 621 455
rect 646 455 652 456
rect 646 451 647 455
rect 651 451 652 455
rect 751 455 752 459
rect 756 458 757 459
rect 782 459 788 460
rect 782 458 783 459
rect 756 456 783 458
rect 756 455 757 456
rect 751 454 757 455
rect 782 455 783 456
rect 787 455 788 459
rect 782 454 788 455
rect 886 459 892 460
rect 886 455 887 459
rect 891 458 892 459
rect 895 459 901 460
rect 895 458 896 459
rect 891 456 896 458
rect 891 455 892 456
rect 886 454 892 455
rect 895 455 896 456
rect 900 455 901 459
rect 895 454 901 455
rect 974 459 980 460
rect 974 455 975 459
rect 979 458 980 459
rect 1031 459 1037 460
rect 1031 458 1032 459
rect 979 456 1032 458
rect 979 455 980 456
rect 974 454 980 455
rect 1031 455 1032 456
rect 1036 455 1037 459
rect 1031 454 1037 455
rect 1054 459 1060 460
rect 1054 455 1055 459
rect 1059 458 1060 459
rect 1159 459 1165 460
rect 1159 458 1160 459
rect 1059 456 1160 458
rect 1059 455 1060 456
rect 1054 454 1060 455
rect 1159 455 1160 456
rect 1164 455 1165 459
rect 1159 454 1165 455
rect 1279 459 1285 460
rect 1279 455 1280 459
rect 1284 458 1285 459
rect 1310 459 1316 460
rect 1310 458 1311 459
rect 1284 456 1311 458
rect 1284 455 1285 456
rect 1279 454 1285 455
rect 1310 455 1311 456
rect 1315 455 1316 459
rect 1310 454 1316 455
rect 1399 459 1405 460
rect 1399 455 1400 459
rect 1404 458 1405 459
rect 1430 459 1436 460
rect 1430 458 1431 459
rect 1404 456 1431 458
rect 1404 455 1405 456
rect 1399 454 1405 455
rect 1430 455 1431 456
rect 1435 455 1436 459
rect 1430 454 1436 455
rect 1455 459 1461 460
rect 1455 455 1456 459
rect 1460 458 1461 459
rect 1511 459 1517 460
rect 1511 458 1512 459
rect 1460 456 1512 458
rect 1460 455 1461 456
rect 1455 454 1461 455
rect 1511 455 1512 456
rect 1516 455 1517 459
rect 1511 454 1517 455
rect 1623 459 1629 460
rect 1623 455 1624 459
rect 1628 458 1629 459
rect 1719 459 1725 460
rect 1628 456 1714 458
rect 1628 455 1629 456
rect 1623 454 1629 455
rect 646 450 652 451
rect 1712 450 1714 456
rect 1719 455 1720 459
rect 1724 455 1725 459
rect 1719 454 1725 455
rect 1774 451 1780 452
rect 1774 450 1775 451
rect 368 448 650 450
rect 1712 448 1775 450
rect 678 447 684 448
rect 678 446 679 447
rect 624 444 679 446
rect 183 439 189 440
rect 183 435 184 439
rect 188 438 189 439
rect 214 439 220 440
rect 214 438 215 439
rect 188 436 215 438
rect 188 435 189 436
rect 183 434 189 435
rect 214 435 215 436
rect 219 435 220 439
rect 214 434 220 435
rect 303 439 309 440
rect 303 435 304 439
rect 308 438 309 439
rect 386 439 392 440
rect 386 438 387 439
rect 308 436 387 438
rect 308 435 309 436
rect 303 434 309 435
rect 386 435 387 436
rect 391 435 392 439
rect 386 434 392 435
rect 463 439 469 440
rect 463 435 464 439
rect 468 438 469 439
rect 624 438 626 444
rect 678 443 679 444
rect 683 443 684 447
rect 1774 447 1775 448
rect 1779 447 1780 451
rect 1774 446 1780 447
rect 1879 451 1888 452
rect 1879 447 1880 451
rect 1887 447 1888 451
rect 1879 446 1888 447
rect 2015 451 2021 452
rect 2015 447 2016 451
rect 2020 450 2021 451
rect 2030 451 2036 452
rect 2030 450 2031 451
rect 2020 448 2031 450
rect 2020 447 2021 448
rect 2015 446 2021 447
rect 2030 447 2031 448
rect 2035 447 2036 451
rect 2030 446 2036 447
rect 2038 451 2044 452
rect 2038 447 2039 451
rect 2043 450 2044 451
rect 2175 451 2181 452
rect 2175 450 2176 451
rect 2043 448 2176 450
rect 2043 447 2044 448
rect 2038 446 2044 447
rect 2175 447 2176 448
rect 2180 447 2181 451
rect 2175 446 2181 447
rect 2343 451 2349 452
rect 2343 447 2344 451
rect 2348 450 2349 451
rect 2374 451 2380 452
rect 2374 450 2375 451
rect 2348 448 2375 450
rect 2348 447 2349 448
rect 2343 446 2349 447
rect 2374 447 2375 448
rect 2379 447 2380 451
rect 2374 446 2380 447
rect 2527 451 2533 452
rect 2527 447 2528 451
rect 2532 450 2533 451
rect 2558 451 2564 452
rect 2558 450 2559 451
rect 2532 448 2559 450
rect 2532 447 2533 448
rect 2527 446 2533 447
rect 2558 447 2559 448
rect 2563 447 2564 451
rect 2558 446 2564 447
rect 2727 451 2736 452
rect 2727 447 2728 451
rect 2735 447 2736 451
rect 2727 446 2736 447
rect 2878 451 2884 452
rect 2878 447 2879 451
rect 2883 450 2884 451
rect 2935 451 2941 452
rect 2935 450 2936 451
rect 2883 448 2936 450
rect 2883 447 2884 448
rect 2878 446 2884 447
rect 2935 447 2936 448
rect 2940 447 2941 451
rect 2935 446 2941 447
rect 2958 451 2964 452
rect 2958 447 2959 451
rect 2963 450 2964 451
rect 3159 451 3165 452
rect 3159 450 3160 451
rect 2963 448 3160 450
rect 2963 447 2964 448
rect 2958 446 2964 447
rect 3159 447 3160 448
rect 3164 447 3165 451
rect 3159 446 3165 447
rect 3383 451 3389 452
rect 3383 447 3384 451
rect 3388 450 3389 451
rect 3430 451 3436 452
rect 3430 450 3431 451
rect 3388 448 3431 450
rect 3388 447 3389 448
rect 3383 446 3389 447
rect 3430 447 3431 448
rect 3435 447 3436 451
rect 3430 446 3436 447
rect 678 442 684 443
rect 468 436 626 438
rect 630 439 637 440
rect 468 435 469 436
rect 463 434 469 435
rect 630 435 631 439
rect 636 435 637 439
rect 630 434 637 435
rect 654 439 660 440
rect 654 435 655 439
rect 659 438 660 439
rect 791 439 797 440
rect 791 438 792 439
rect 659 436 792 438
rect 659 435 660 436
rect 654 434 660 435
rect 791 435 792 436
rect 796 435 797 439
rect 791 434 797 435
rect 951 439 957 440
rect 951 435 952 439
rect 956 438 957 439
rect 983 439 989 440
rect 983 438 984 439
rect 956 436 984 438
rect 956 435 957 436
rect 951 434 957 435
rect 983 435 984 436
rect 988 435 989 439
rect 983 434 989 435
rect 1095 439 1101 440
rect 1095 435 1096 439
rect 1100 438 1101 439
rect 1126 439 1132 440
rect 1126 438 1127 439
rect 1100 436 1127 438
rect 1100 435 1101 436
rect 1095 434 1101 435
rect 1126 435 1127 436
rect 1131 435 1132 439
rect 1126 434 1132 435
rect 1231 439 1237 440
rect 1231 435 1232 439
rect 1236 438 1237 439
rect 1294 439 1300 440
rect 1294 438 1295 439
rect 1236 436 1295 438
rect 1236 435 1237 436
rect 1231 434 1237 435
rect 1294 435 1295 436
rect 1299 435 1300 439
rect 1294 434 1300 435
rect 1302 439 1308 440
rect 1302 435 1303 439
rect 1307 438 1308 439
rect 1359 439 1365 440
rect 1359 438 1360 439
rect 1307 436 1360 438
rect 1307 435 1308 436
rect 1302 434 1308 435
rect 1359 435 1360 436
rect 1364 435 1365 439
rect 1359 434 1365 435
rect 1382 439 1388 440
rect 1382 435 1383 439
rect 1387 438 1388 439
rect 1487 439 1493 440
rect 1487 438 1488 439
rect 1387 436 1488 438
rect 1387 435 1388 436
rect 1382 434 1388 435
rect 1487 435 1488 436
rect 1492 435 1493 439
rect 1487 434 1493 435
rect 1510 439 1516 440
rect 1510 435 1511 439
rect 1515 438 1516 439
rect 1615 439 1621 440
rect 1615 438 1616 439
rect 1515 436 1616 438
rect 1515 435 1516 436
rect 1510 434 1516 435
rect 1615 435 1616 436
rect 1620 435 1621 439
rect 1615 434 1621 435
rect 1638 439 1644 440
rect 1638 435 1639 439
rect 1643 438 1644 439
rect 1719 439 1725 440
rect 1719 438 1720 439
rect 1643 436 1720 438
rect 1643 435 1644 436
rect 1638 434 1644 435
rect 1719 435 1720 436
rect 1724 435 1725 439
rect 1719 434 1725 435
rect 1742 439 1748 440
rect 1742 435 1743 439
rect 1747 438 1748 439
rect 1879 439 1885 440
rect 1879 438 1880 439
rect 1747 436 1880 438
rect 1747 435 1748 436
rect 1742 434 1748 435
rect 1879 435 1880 436
rect 1884 435 1885 439
rect 1879 434 1885 435
rect 1902 439 1908 440
rect 1902 435 1903 439
rect 1907 438 1908 439
rect 2007 439 2013 440
rect 2007 438 2008 439
rect 1907 436 2008 438
rect 1907 435 1908 436
rect 1902 434 1908 435
rect 2007 435 2008 436
rect 2012 435 2013 439
rect 2007 434 2013 435
rect 2118 439 2124 440
rect 2118 435 2119 439
rect 2123 438 2124 439
rect 2159 439 2165 440
rect 2159 438 2160 439
rect 2123 436 2160 438
rect 2123 435 2124 436
rect 2118 434 2124 435
rect 2159 435 2160 436
rect 2164 435 2165 439
rect 2159 434 2165 435
rect 2319 439 2325 440
rect 2319 435 2320 439
rect 2324 438 2325 439
rect 2358 439 2364 440
rect 2358 438 2359 439
rect 2324 436 2359 438
rect 2324 435 2325 436
rect 2319 434 2325 435
rect 2358 435 2359 436
rect 2363 435 2364 439
rect 2358 434 2364 435
rect 2402 439 2408 440
rect 2402 435 2403 439
rect 2407 438 2408 439
rect 2503 439 2509 440
rect 2503 438 2504 439
rect 2407 436 2504 438
rect 2407 435 2408 436
rect 2402 434 2408 435
rect 2503 435 2504 436
rect 2508 435 2509 439
rect 2503 434 2509 435
rect 2526 439 2532 440
rect 2526 435 2527 439
rect 2531 438 2532 439
rect 2703 439 2709 440
rect 2703 438 2704 439
rect 2531 436 2704 438
rect 2531 435 2532 436
rect 2526 434 2532 435
rect 2703 435 2704 436
rect 2708 435 2709 439
rect 2703 434 2709 435
rect 2726 439 2732 440
rect 2726 435 2727 439
rect 2731 438 2732 439
rect 2919 439 2925 440
rect 2919 438 2920 439
rect 2731 436 2920 438
rect 2731 435 2732 436
rect 2726 434 2732 435
rect 2919 435 2920 436
rect 2924 435 2925 439
rect 2919 434 2925 435
rect 2942 439 2948 440
rect 2942 435 2943 439
rect 2947 438 2948 439
rect 3151 439 3157 440
rect 3151 438 3152 439
rect 2947 436 3152 438
rect 2947 435 2948 436
rect 2942 434 2948 435
rect 3151 435 3152 436
rect 3156 435 3157 439
rect 3151 434 3157 435
rect 3342 439 3348 440
rect 3342 435 3343 439
rect 3347 438 3348 439
rect 3383 439 3389 440
rect 3383 438 3384 439
rect 3347 436 3384 438
rect 3347 435 3348 436
rect 3342 434 3348 435
rect 3383 435 3384 436
rect 3388 435 3389 439
rect 3383 434 3389 435
rect 110 424 116 425
rect 1766 424 1772 425
rect 110 420 111 424
rect 115 420 116 424
rect 110 419 116 420
rect 134 423 140 424
rect 134 419 135 423
rect 139 419 140 423
rect 134 418 140 419
rect 254 423 260 424
rect 254 419 255 423
rect 259 419 260 423
rect 254 418 260 419
rect 414 423 420 424
rect 414 419 415 423
rect 419 419 420 423
rect 414 418 420 419
rect 582 423 588 424
rect 582 419 583 423
rect 587 419 588 423
rect 582 418 588 419
rect 742 423 748 424
rect 742 419 743 423
rect 747 419 748 423
rect 742 418 748 419
rect 902 423 908 424
rect 902 419 903 423
rect 907 419 908 423
rect 902 418 908 419
rect 1046 423 1052 424
rect 1046 419 1047 423
rect 1051 419 1052 423
rect 1046 418 1052 419
rect 1182 423 1188 424
rect 1182 419 1183 423
rect 1187 419 1188 423
rect 1182 418 1188 419
rect 1310 423 1316 424
rect 1310 419 1311 423
rect 1315 419 1316 423
rect 1310 418 1316 419
rect 1438 423 1444 424
rect 1438 419 1439 423
rect 1443 419 1444 423
rect 1438 418 1444 419
rect 1566 423 1572 424
rect 1566 419 1567 423
rect 1571 419 1572 423
rect 1566 418 1572 419
rect 1670 423 1676 424
rect 1670 419 1671 423
rect 1675 419 1676 423
rect 1766 420 1767 424
rect 1771 420 1772 424
rect 1766 419 1772 420
rect 1806 424 1812 425
rect 3462 424 3468 425
rect 1806 420 1807 424
rect 1811 420 1812 424
rect 1806 419 1812 420
rect 1830 423 1836 424
rect 1830 419 1831 423
rect 1835 419 1836 423
rect 1670 418 1676 419
rect 1830 418 1836 419
rect 1958 423 1964 424
rect 1958 419 1959 423
rect 1963 419 1964 423
rect 1958 418 1964 419
rect 2110 423 2116 424
rect 2110 419 2111 423
rect 2115 419 2116 423
rect 2110 418 2116 419
rect 2270 423 2276 424
rect 2270 419 2271 423
rect 2275 419 2276 423
rect 2270 418 2276 419
rect 2454 423 2460 424
rect 2454 419 2455 423
rect 2459 419 2460 423
rect 2454 418 2460 419
rect 2654 423 2660 424
rect 2654 419 2655 423
rect 2659 419 2660 423
rect 2654 418 2660 419
rect 2870 423 2876 424
rect 2870 419 2871 423
rect 2875 419 2876 423
rect 2870 418 2876 419
rect 3102 423 3108 424
rect 3102 419 3103 423
rect 3107 419 3108 423
rect 3102 418 3108 419
rect 3334 423 3340 424
rect 3334 419 3335 423
rect 3339 419 3340 423
rect 3462 420 3463 424
rect 3467 420 3468 424
rect 3462 419 3468 420
rect 3334 418 3340 419
rect 214 415 220 416
rect 214 411 215 415
rect 219 414 220 415
rect 386 415 392 416
rect 219 412 297 414
rect 219 411 220 412
rect 214 410 220 411
rect 386 411 387 415
rect 391 414 392 415
rect 654 415 660 416
rect 391 412 457 414
rect 391 411 392 412
rect 386 410 392 411
rect 654 411 655 415
rect 659 411 660 415
rect 654 410 660 411
rect 678 415 684 416
rect 678 411 679 415
rect 683 414 684 415
rect 974 415 980 416
rect 683 412 785 414
rect 683 411 684 412
rect 678 410 684 411
rect 974 411 975 415
rect 979 411 980 415
rect 974 410 980 411
rect 983 415 989 416
rect 983 411 984 415
rect 988 414 989 415
rect 1126 415 1132 416
rect 988 412 1089 414
rect 988 411 989 412
rect 983 410 989 411
rect 1126 411 1127 415
rect 1131 414 1132 415
rect 1382 415 1388 416
rect 1131 412 1225 414
rect 1131 411 1132 412
rect 1126 410 1132 411
rect 1382 411 1383 415
rect 1387 411 1388 415
rect 1382 410 1388 411
rect 1510 415 1516 416
rect 1510 411 1511 415
rect 1515 411 1516 415
rect 1510 410 1516 411
rect 1638 415 1644 416
rect 1638 411 1639 415
rect 1643 411 1644 415
rect 1638 410 1644 411
rect 1742 415 1748 416
rect 1742 411 1743 415
rect 1747 411 1748 415
rect 1742 410 1748 411
rect 1902 415 1908 416
rect 1902 411 1903 415
rect 1907 411 1908 415
rect 1902 410 1908 411
rect 2030 415 2036 416
rect 2030 411 2031 415
rect 2035 411 2036 415
rect 2030 410 2036 411
rect 2074 415 2080 416
rect 2074 411 2075 415
rect 2079 414 2080 415
rect 2402 415 2408 416
rect 2402 414 2403 415
rect 2079 412 2153 414
rect 2345 412 2403 414
rect 2079 411 2080 412
rect 2074 410 2080 411
rect 2402 411 2403 412
rect 2407 411 2408 415
rect 2402 410 2408 411
rect 2526 415 2532 416
rect 2526 411 2527 415
rect 2531 411 2532 415
rect 2526 410 2532 411
rect 2726 415 2732 416
rect 2726 411 2727 415
rect 2731 411 2732 415
rect 2726 410 2732 411
rect 2942 415 2948 416
rect 2942 411 2943 415
rect 2947 411 2948 415
rect 2942 410 2948 411
rect 3018 415 3024 416
rect 3018 411 3019 415
rect 3023 414 3024 415
rect 3023 412 3145 414
rect 3023 411 3024 412
rect 3018 410 3024 411
rect 3406 411 3412 412
rect 110 407 116 408
rect 110 403 111 407
rect 115 403 116 407
rect 198 407 204 408
rect 110 402 116 403
rect 134 404 140 405
rect 134 400 135 404
rect 139 400 140 404
rect 198 403 199 407
rect 203 406 204 407
rect 208 406 210 409
rect 203 404 210 406
rect 1766 407 1772 408
rect 254 404 260 405
rect 203 403 204 404
rect 198 402 204 403
rect 134 399 140 400
rect 254 400 255 404
rect 259 400 260 404
rect 254 399 260 400
rect 414 404 420 405
rect 414 400 415 404
rect 419 400 420 404
rect 414 399 420 400
rect 582 404 588 405
rect 582 400 583 404
rect 587 400 588 404
rect 582 399 588 400
rect 742 404 748 405
rect 742 400 743 404
rect 747 400 748 404
rect 742 399 748 400
rect 902 404 908 405
rect 902 400 903 404
rect 907 400 908 404
rect 902 399 908 400
rect 1046 404 1052 405
rect 1046 400 1047 404
rect 1051 400 1052 404
rect 1046 399 1052 400
rect 1182 404 1188 405
rect 1182 400 1183 404
rect 1187 400 1188 404
rect 1182 399 1188 400
rect 1310 404 1316 405
rect 1310 400 1311 404
rect 1315 400 1316 404
rect 1310 399 1316 400
rect 1438 404 1444 405
rect 1438 400 1439 404
rect 1443 400 1444 404
rect 1438 399 1444 400
rect 1566 404 1572 405
rect 1566 400 1567 404
rect 1571 400 1572 404
rect 1566 399 1572 400
rect 1670 404 1676 405
rect 1670 400 1671 404
rect 1675 400 1676 404
rect 1766 403 1767 407
rect 1771 403 1772 407
rect 1766 402 1772 403
rect 1806 407 1812 408
rect 1806 403 1807 407
rect 1811 403 1812 407
rect 3406 407 3407 411
rect 3411 407 3412 411
rect 3406 406 3412 407
rect 3462 407 3468 408
rect 1806 402 1812 403
rect 1830 404 1836 405
rect 1670 399 1676 400
rect 1830 400 1831 404
rect 1835 400 1836 404
rect 1830 399 1836 400
rect 1958 404 1964 405
rect 1958 400 1959 404
rect 1963 400 1964 404
rect 1958 399 1964 400
rect 2110 404 2116 405
rect 2110 400 2111 404
rect 2115 400 2116 404
rect 2110 399 2116 400
rect 2270 404 2276 405
rect 2270 400 2271 404
rect 2275 400 2276 404
rect 2270 399 2276 400
rect 2454 404 2460 405
rect 2454 400 2455 404
rect 2459 400 2460 404
rect 2454 399 2460 400
rect 2654 404 2660 405
rect 2654 400 2655 404
rect 2659 400 2660 404
rect 2654 399 2660 400
rect 2870 404 2876 405
rect 2870 400 2871 404
rect 2875 400 2876 404
rect 2870 399 2876 400
rect 3102 404 3108 405
rect 3102 400 3103 404
rect 3107 400 3108 404
rect 3102 399 3108 400
rect 3334 404 3340 405
rect 3334 400 3335 404
rect 3339 400 3340 404
rect 3462 403 3463 407
rect 3467 403 3468 407
rect 3462 402 3468 403
rect 3334 399 3340 400
rect 1294 375 1300 376
rect 1294 371 1295 375
rect 1299 374 1300 375
rect 2074 375 2080 376
rect 2074 374 2075 375
rect 1299 372 2075 374
rect 1299 371 1300 372
rect 1294 370 1300 371
rect 2074 371 2075 372
rect 2079 371 2080 375
rect 2074 370 2080 371
rect 2730 371 2736 372
rect 2730 367 2731 371
rect 2735 370 2736 371
rect 3030 371 3036 372
rect 3030 370 3031 371
rect 2735 368 3031 370
rect 2735 367 2736 368
rect 2730 366 2736 367
rect 3030 367 3031 368
rect 3035 367 3036 371
rect 3030 366 3036 367
rect 2634 363 2640 364
rect 2634 359 2635 363
rect 2639 362 2640 363
rect 3018 363 3024 364
rect 3018 362 3019 363
rect 2639 360 3019 362
rect 2639 359 2640 360
rect 2634 358 2640 359
rect 3018 359 3019 360
rect 3023 359 3024 363
rect 3018 358 3024 359
rect 134 356 140 357
rect 110 353 116 354
rect 110 349 111 353
rect 115 349 116 353
rect 134 352 135 356
rect 139 352 140 356
rect 134 351 140 352
rect 222 356 228 357
rect 222 352 223 356
rect 227 352 228 356
rect 222 351 228 352
rect 342 356 348 357
rect 342 352 343 356
rect 347 352 348 356
rect 342 351 348 352
rect 470 356 476 357
rect 470 352 471 356
rect 475 352 476 356
rect 470 351 476 352
rect 598 356 604 357
rect 598 352 599 356
rect 603 352 604 356
rect 598 351 604 352
rect 718 356 724 357
rect 718 352 719 356
rect 723 352 724 356
rect 718 351 724 352
rect 838 356 844 357
rect 838 352 839 356
rect 843 352 844 356
rect 838 351 844 352
rect 958 356 964 357
rect 958 352 959 356
rect 963 352 964 356
rect 958 351 964 352
rect 1078 356 1084 357
rect 1078 352 1079 356
rect 1083 352 1084 356
rect 1078 351 1084 352
rect 1206 356 1212 357
rect 1206 352 1207 356
rect 1211 352 1212 356
rect 1926 356 1932 357
rect 1206 351 1212 352
rect 1766 353 1772 354
rect 110 348 116 349
rect 1766 349 1767 353
rect 1771 349 1772 353
rect 1766 348 1772 349
rect 1806 353 1812 354
rect 1806 349 1807 353
rect 1811 349 1812 353
rect 1926 352 1927 356
rect 1931 352 1932 356
rect 1926 351 1932 352
rect 2038 356 2044 357
rect 2038 352 2039 356
rect 2043 352 2044 356
rect 2038 351 2044 352
rect 2158 356 2164 357
rect 2158 352 2159 356
rect 2163 352 2164 356
rect 2158 351 2164 352
rect 2286 356 2292 357
rect 2286 352 2287 356
rect 2291 352 2292 356
rect 2286 351 2292 352
rect 2422 356 2428 357
rect 2422 352 2423 356
rect 2427 352 2428 356
rect 2422 351 2428 352
rect 2582 356 2588 357
rect 2582 352 2583 356
rect 2587 352 2588 356
rect 2582 351 2588 352
rect 2758 356 2764 357
rect 2758 352 2759 356
rect 2763 352 2764 356
rect 2758 351 2764 352
rect 2950 356 2956 357
rect 2950 352 2951 356
rect 2955 352 2956 356
rect 2950 351 2956 352
rect 3150 356 3156 357
rect 3150 352 3151 356
rect 3155 352 3156 356
rect 3150 351 3156 352
rect 3358 356 3364 357
rect 3358 352 3359 356
rect 3363 352 3364 356
rect 3358 351 3364 352
rect 3462 353 3468 354
rect 1806 348 1812 349
rect 3462 349 3463 353
rect 3467 349 3468 353
rect 3462 348 3468 349
rect 206 347 212 348
rect 206 343 207 347
rect 211 343 212 347
rect 206 342 212 343
rect 294 347 300 348
rect 294 343 295 347
rect 299 343 300 347
rect 294 342 300 343
rect 414 347 420 348
rect 414 343 415 347
rect 419 343 420 347
rect 414 342 420 343
rect 542 347 548 348
rect 542 343 543 347
rect 547 343 548 347
rect 542 342 548 343
rect 550 347 556 348
rect 550 343 551 347
rect 555 346 556 347
rect 822 347 828 348
rect 822 346 823 347
rect 555 344 641 346
rect 793 344 823 346
rect 555 343 556 344
rect 550 342 556 343
rect 822 343 823 344
rect 827 343 828 347
rect 822 342 828 343
rect 910 347 916 348
rect 910 343 911 347
rect 915 343 916 347
rect 910 342 916 343
rect 1030 347 1036 348
rect 1030 343 1031 347
rect 1035 343 1036 347
rect 1030 342 1036 343
rect 1150 347 1156 348
rect 1150 343 1151 347
rect 1155 343 1156 347
rect 1150 342 1156 343
rect 1159 347 1165 348
rect 1159 343 1160 347
rect 1164 346 1165 347
rect 1998 347 2004 348
rect 1164 344 1249 346
rect 1164 343 1165 344
rect 1159 342 1165 343
rect 1998 343 1999 347
rect 2003 343 2004 347
rect 2118 347 2124 348
rect 2118 346 2119 347
rect 2113 344 2119 346
rect 1998 342 2004 343
rect 2118 343 2119 344
rect 2123 343 2124 347
rect 2118 342 2124 343
rect 2126 347 2132 348
rect 2126 343 2127 347
rect 2131 346 2132 347
rect 2238 347 2244 348
rect 2131 344 2201 346
rect 2131 343 2132 344
rect 2126 342 2132 343
rect 2238 343 2239 347
rect 2243 346 2244 347
rect 2366 347 2372 348
rect 2243 344 2329 346
rect 2243 343 2244 344
rect 2238 342 2244 343
rect 2366 343 2367 347
rect 2371 346 2372 347
rect 2654 347 2660 348
rect 2371 344 2465 346
rect 2371 343 2372 344
rect 2366 342 2372 343
rect 2654 343 2655 347
rect 2659 343 2660 347
rect 2654 342 2660 343
rect 2830 347 2836 348
rect 2830 343 2831 347
rect 2835 343 2836 347
rect 2830 342 2836 343
rect 3022 347 3028 348
rect 3022 343 3023 347
rect 3027 343 3028 347
rect 3022 342 3028 343
rect 3030 347 3036 348
rect 3030 343 3031 347
rect 3035 346 3036 347
rect 3422 347 3428 348
rect 3035 344 3193 346
rect 3035 343 3036 344
rect 3030 342 3036 343
rect 3422 343 3423 347
rect 3427 343 3428 347
rect 3422 342 3428 343
rect 134 337 140 338
rect 110 336 116 337
rect 110 332 111 336
rect 115 332 116 336
rect 134 333 135 337
rect 139 333 140 337
rect 134 332 140 333
rect 222 337 228 338
rect 222 333 223 337
rect 227 333 228 337
rect 222 332 228 333
rect 342 337 348 338
rect 342 333 343 337
rect 347 333 348 337
rect 342 332 348 333
rect 470 337 476 338
rect 470 333 471 337
rect 475 333 476 337
rect 470 332 476 333
rect 598 337 604 338
rect 598 333 599 337
rect 603 333 604 337
rect 598 332 604 333
rect 718 337 724 338
rect 718 333 719 337
rect 723 333 724 337
rect 718 332 724 333
rect 838 337 844 338
rect 838 333 839 337
rect 843 333 844 337
rect 838 332 844 333
rect 958 337 964 338
rect 958 333 959 337
rect 963 333 964 337
rect 958 332 964 333
rect 1078 337 1084 338
rect 1078 333 1079 337
rect 1083 333 1084 337
rect 1078 332 1084 333
rect 1206 337 1212 338
rect 1926 337 1932 338
rect 1206 333 1207 337
rect 1211 333 1212 337
rect 1206 332 1212 333
rect 1766 336 1772 337
rect 1766 332 1767 336
rect 1771 332 1772 336
rect 110 331 116 332
rect 1766 331 1772 332
rect 1806 336 1812 337
rect 1806 332 1807 336
rect 1811 332 1812 336
rect 1926 333 1927 337
rect 1931 333 1932 337
rect 1926 332 1932 333
rect 2038 337 2044 338
rect 2038 333 2039 337
rect 2043 333 2044 337
rect 2038 332 2044 333
rect 2158 337 2164 338
rect 2158 333 2159 337
rect 2163 333 2164 337
rect 2158 332 2164 333
rect 2286 337 2292 338
rect 2286 333 2287 337
rect 2291 333 2292 337
rect 2286 332 2292 333
rect 2422 337 2428 338
rect 2422 333 2423 337
rect 2427 333 2428 337
rect 2422 332 2428 333
rect 2582 337 2588 338
rect 2582 333 2583 337
rect 2587 333 2588 337
rect 2582 332 2588 333
rect 2758 337 2764 338
rect 2758 333 2759 337
rect 2763 333 2764 337
rect 2758 332 2764 333
rect 2950 337 2956 338
rect 2950 333 2951 337
rect 2955 333 2956 337
rect 2950 332 2956 333
rect 3150 337 3156 338
rect 3150 333 3151 337
rect 3155 333 3156 337
rect 3150 332 3156 333
rect 3358 337 3364 338
rect 3358 333 3359 337
rect 3363 333 3364 337
rect 3358 332 3364 333
rect 3462 336 3468 337
rect 3462 332 3463 336
rect 3467 332 3468 336
rect 1806 331 1812 332
rect 3462 331 3468 332
rect 183 319 189 320
rect 183 315 184 319
rect 188 318 189 319
rect 198 319 204 320
rect 198 318 199 319
rect 188 316 199 318
rect 188 315 189 316
rect 183 314 189 315
rect 198 315 199 316
rect 203 315 204 319
rect 198 314 204 315
rect 206 319 212 320
rect 206 315 207 319
rect 211 318 212 319
rect 271 319 277 320
rect 271 318 272 319
rect 211 316 272 318
rect 211 315 212 316
rect 206 314 212 315
rect 271 315 272 316
rect 276 315 277 319
rect 271 314 277 315
rect 294 319 300 320
rect 294 315 295 319
rect 299 318 300 319
rect 391 319 397 320
rect 391 318 392 319
rect 299 316 392 318
rect 299 315 300 316
rect 294 314 300 315
rect 391 315 392 316
rect 396 315 397 319
rect 391 314 397 315
rect 414 319 420 320
rect 414 315 415 319
rect 419 318 420 319
rect 519 319 525 320
rect 519 318 520 319
rect 419 316 520 318
rect 419 315 420 316
rect 414 314 420 315
rect 519 315 520 316
rect 524 315 525 319
rect 519 314 525 315
rect 542 319 548 320
rect 542 315 543 319
rect 547 318 548 319
rect 647 319 653 320
rect 647 318 648 319
rect 547 316 648 318
rect 547 315 548 316
rect 542 314 548 315
rect 647 315 648 316
rect 652 315 653 319
rect 647 314 653 315
rect 767 319 773 320
rect 767 315 768 319
rect 772 318 773 319
rect 791 319 797 320
rect 791 318 792 319
rect 772 316 792 318
rect 772 315 773 316
rect 767 314 773 315
rect 791 315 792 316
rect 796 315 797 319
rect 791 314 797 315
rect 822 319 828 320
rect 822 315 823 319
rect 827 318 828 319
rect 887 319 893 320
rect 887 318 888 319
rect 827 316 888 318
rect 827 315 828 316
rect 822 314 828 315
rect 887 315 888 316
rect 892 315 893 319
rect 887 314 893 315
rect 910 319 916 320
rect 910 315 911 319
rect 915 318 916 319
rect 1007 319 1013 320
rect 1007 318 1008 319
rect 915 316 1008 318
rect 915 315 916 316
rect 910 314 916 315
rect 1007 315 1008 316
rect 1012 315 1013 319
rect 1007 314 1013 315
rect 1030 319 1036 320
rect 1030 315 1031 319
rect 1035 318 1036 319
rect 1127 319 1133 320
rect 1127 318 1128 319
rect 1035 316 1128 318
rect 1035 315 1036 316
rect 1030 314 1036 315
rect 1127 315 1128 316
rect 1132 315 1133 319
rect 1127 314 1133 315
rect 1150 319 1156 320
rect 1150 315 1151 319
rect 1155 318 1156 319
rect 1255 319 1261 320
rect 1255 318 1256 319
rect 1155 316 1256 318
rect 1155 315 1156 316
rect 1150 314 1156 315
rect 1255 315 1256 316
rect 1260 315 1261 319
rect 1255 314 1261 315
rect 1975 319 1981 320
rect 1975 315 1976 319
rect 1980 318 1981 319
rect 1998 319 2004 320
rect 1980 316 1994 318
rect 1980 315 1981 316
rect 1975 314 1981 315
rect 550 311 556 312
rect 550 310 551 311
rect 319 308 551 310
rect 311 303 317 304
rect 311 299 312 303
rect 316 302 317 303
rect 319 302 321 308
rect 550 307 551 308
rect 555 307 556 311
rect 550 306 556 307
rect 1159 311 1165 312
rect 1159 307 1160 311
rect 1164 307 1165 311
rect 1992 310 1994 316
rect 1998 315 1999 319
rect 2003 318 2004 319
rect 2087 319 2093 320
rect 2087 318 2088 319
rect 2003 316 2088 318
rect 2003 315 2004 316
rect 1998 314 2004 315
rect 2087 315 2088 316
rect 2092 315 2093 319
rect 2087 314 2093 315
rect 2207 319 2213 320
rect 2207 315 2208 319
rect 2212 318 2213 319
rect 2238 319 2244 320
rect 2238 318 2239 319
rect 2212 316 2239 318
rect 2212 315 2213 316
rect 2207 314 2213 315
rect 2238 315 2239 316
rect 2243 315 2244 319
rect 2238 314 2244 315
rect 2335 319 2341 320
rect 2335 315 2336 319
rect 2340 318 2341 319
rect 2366 319 2372 320
rect 2366 318 2367 319
rect 2340 316 2367 318
rect 2340 315 2341 316
rect 2335 314 2341 315
rect 2366 315 2367 316
rect 2371 315 2372 319
rect 2366 314 2372 315
rect 2470 319 2477 320
rect 2470 315 2471 319
rect 2476 315 2477 319
rect 2470 314 2477 315
rect 2631 319 2640 320
rect 2631 315 2632 319
rect 2639 315 2640 319
rect 2631 314 2640 315
rect 2654 319 2660 320
rect 2654 315 2655 319
rect 2659 318 2660 319
rect 2807 319 2813 320
rect 2807 318 2808 319
rect 2659 316 2808 318
rect 2659 315 2660 316
rect 2654 314 2660 315
rect 2807 315 2808 316
rect 2812 315 2813 319
rect 2807 314 2813 315
rect 2830 319 2836 320
rect 2830 315 2831 319
rect 2835 318 2836 319
rect 2999 319 3005 320
rect 2999 318 3000 319
rect 2835 316 3000 318
rect 2835 315 2836 316
rect 2830 314 2836 315
rect 2999 315 3000 316
rect 3004 315 3005 319
rect 2999 314 3005 315
rect 3022 319 3028 320
rect 3022 315 3023 319
rect 3027 318 3028 319
rect 3199 319 3205 320
rect 3199 318 3200 319
rect 3027 316 3200 318
rect 3027 315 3028 316
rect 3022 314 3028 315
rect 3199 315 3200 316
rect 3204 315 3205 319
rect 3199 314 3205 315
rect 3406 319 3413 320
rect 3406 315 3407 319
rect 3412 315 3413 319
rect 3406 314 3413 315
rect 2126 311 2132 312
rect 2126 310 2127 311
rect 1992 308 2127 310
rect 1159 306 1165 307
rect 2126 307 2127 308
rect 2131 307 2132 311
rect 2126 306 2132 307
rect 2271 307 2280 308
rect 1116 304 1161 306
rect 316 300 321 302
rect 334 303 340 304
rect 316 299 317 300
rect 311 298 317 299
rect 334 299 335 303
rect 339 302 340 303
rect 423 303 429 304
rect 423 302 424 303
rect 339 300 424 302
rect 339 299 340 300
rect 334 298 340 299
rect 423 299 424 300
rect 428 299 429 303
rect 423 298 429 299
rect 446 303 452 304
rect 446 299 447 303
rect 451 302 452 303
rect 535 303 541 304
rect 535 302 536 303
rect 451 300 536 302
rect 451 299 452 300
rect 446 298 452 299
rect 535 299 536 300
rect 540 299 541 303
rect 535 298 541 299
rect 558 303 564 304
rect 558 299 559 303
rect 563 302 564 303
rect 647 303 653 304
rect 647 302 648 303
rect 563 300 648 302
rect 563 299 564 300
rect 558 298 564 299
rect 647 299 648 300
rect 652 299 653 303
rect 647 298 653 299
rect 759 303 765 304
rect 759 299 760 303
rect 764 302 765 303
rect 774 303 780 304
rect 774 302 775 303
rect 764 300 775 302
rect 764 299 765 300
rect 759 298 765 299
rect 774 299 775 300
rect 779 299 780 303
rect 774 298 780 299
rect 863 303 869 304
rect 863 299 864 303
rect 868 302 869 303
rect 895 303 901 304
rect 895 302 896 303
rect 868 300 896 302
rect 868 299 869 300
rect 863 298 869 299
rect 895 299 896 300
rect 900 299 901 303
rect 895 298 901 299
rect 967 303 973 304
rect 967 299 968 303
rect 972 302 973 303
rect 982 303 988 304
rect 982 302 983 303
rect 972 300 983 302
rect 972 299 973 300
rect 967 298 973 299
rect 982 299 983 300
rect 987 299 988 303
rect 982 298 988 299
rect 1071 303 1077 304
rect 1071 299 1072 303
rect 1076 302 1077 303
rect 1116 302 1118 304
rect 1175 303 1181 304
rect 1175 302 1176 303
rect 1076 300 1118 302
rect 1159 300 1176 302
rect 1076 299 1077 300
rect 1071 298 1077 299
rect 1159 298 1161 300
rect 1175 299 1176 300
rect 1180 299 1181 303
rect 1175 298 1181 299
rect 1198 303 1204 304
rect 1198 299 1199 303
rect 1203 302 1204 303
rect 1287 303 1293 304
rect 1287 302 1288 303
rect 1203 300 1288 302
rect 1203 299 1204 300
rect 1198 298 1204 299
rect 1287 299 1288 300
rect 1292 299 1293 303
rect 2271 303 2272 307
rect 2279 303 2280 307
rect 2271 302 2280 303
rect 2294 307 2300 308
rect 2294 303 2295 307
rect 2299 306 2300 307
rect 2359 307 2365 308
rect 2359 306 2360 307
rect 2299 304 2360 306
rect 2299 303 2300 304
rect 2294 302 2300 303
rect 2359 303 2360 304
rect 2364 303 2365 307
rect 2359 302 2365 303
rect 2382 307 2388 308
rect 2382 303 2383 307
rect 2387 306 2388 307
rect 2447 307 2453 308
rect 2447 306 2448 307
rect 2387 304 2448 306
rect 2387 303 2388 304
rect 2382 302 2388 303
rect 2447 303 2448 304
rect 2452 303 2453 307
rect 2447 302 2453 303
rect 2535 307 2541 308
rect 2535 303 2536 307
rect 2540 306 2541 307
rect 2566 307 2572 308
rect 2566 306 2567 307
rect 2540 304 2567 306
rect 2540 303 2541 304
rect 2535 302 2541 303
rect 2566 303 2567 304
rect 2571 303 2572 307
rect 2566 302 2572 303
rect 2623 307 2632 308
rect 2623 303 2624 307
rect 2631 303 2632 307
rect 2623 302 2632 303
rect 2727 307 2736 308
rect 2727 303 2728 307
rect 2735 303 2736 307
rect 2727 302 2736 303
rect 2750 307 2756 308
rect 2750 303 2751 307
rect 2755 306 2756 307
rect 2847 307 2853 308
rect 2847 306 2848 307
rect 2755 304 2848 306
rect 2755 303 2756 304
rect 2750 302 2756 303
rect 2847 303 2848 304
rect 2852 303 2853 307
rect 2847 302 2853 303
rect 2870 307 2876 308
rect 2870 303 2871 307
rect 2875 306 2876 307
rect 2975 307 2981 308
rect 2975 306 2976 307
rect 2875 304 2976 306
rect 2875 303 2876 304
rect 2870 302 2876 303
rect 2975 303 2976 304
rect 2980 303 2981 307
rect 2975 302 2981 303
rect 2998 307 3004 308
rect 2998 303 2999 307
rect 3003 306 3004 307
rect 3119 307 3125 308
rect 3119 306 3120 307
rect 3003 304 3120 306
rect 3003 303 3004 304
rect 2998 302 3004 303
rect 3119 303 3120 304
rect 3124 303 3125 307
rect 3119 302 3125 303
rect 3142 307 3148 308
rect 3142 303 3143 307
rect 3147 306 3148 307
rect 3271 307 3277 308
rect 3271 306 3272 307
rect 3147 304 3272 306
rect 3147 303 3148 304
rect 3142 302 3148 303
rect 3271 303 3272 304
rect 3276 303 3277 307
rect 3271 302 3277 303
rect 3415 307 3421 308
rect 3415 303 3416 307
rect 3420 303 3421 307
rect 3415 302 3421 303
rect 1287 298 1293 299
rect 1112 296 1161 298
rect 110 288 116 289
rect 110 284 111 288
rect 115 284 116 288
rect 110 283 116 284
rect 262 287 268 288
rect 262 283 263 287
rect 267 283 268 287
rect 262 282 268 283
rect 374 287 380 288
rect 374 283 375 287
rect 379 283 380 287
rect 374 282 380 283
rect 486 287 492 288
rect 486 283 487 287
rect 491 283 492 287
rect 486 282 492 283
rect 598 287 604 288
rect 598 283 599 287
rect 603 283 604 287
rect 598 282 604 283
rect 710 287 716 288
rect 710 283 711 287
rect 715 283 716 287
rect 710 282 716 283
rect 814 287 820 288
rect 814 283 815 287
rect 819 283 820 287
rect 814 282 820 283
rect 918 287 924 288
rect 918 283 919 287
rect 923 283 924 287
rect 918 282 924 283
rect 1022 287 1028 288
rect 1022 283 1023 287
rect 1027 283 1028 287
rect 1022 282 1028 283
rect 334 279 340 280
rect 334 275 335 279
rect 339 275 340 279
rect 334 274 340 275
rect 446 279 452 280
rect 446 275 447 279
rect 451 275 452 279
rect 446 274 452 275
rect 558 279 564 280
rect 558 275 559 279
rect 563 275 564 279
rect 558 274 564 275
rect 586 279 592 280
rect 586 275 587 279
rect 591 278 592 279
rect 791 279 797 280
rect 591 276 641 278
rect 591 275 592 276
rect 586 274 592 275
rect 782 275 788 276
rect 110 271 116 272
rect 110 267 111 271
rect 115 267 116 271
rect 782 271 783 275
rect 787 271 788 275
rect 791 275 792 279
rect 796 278 797 279
rect 895 279 901 280
rect 796 276 857 278
rect 796 275 797 276
rect 791 274 797 275
rect 895 275 896 279
rect 900 278 901 279
rect 1112 278 1114 296
rect 1806 292 1812 293
rect 3462 292 3468 293
rect 1766 288 1772 289
rect 1126 287 1132 288
rect 1126 283 1127 287
rect 1131 283 1132 287
rect 1126 282 1132 283
rect 1238 287 1244 288
rect 1238 283 1239 287
rect 1243 283 1244 287
rect 1766 284 1767 288
rect 1771 284 1772 288
rect 1806 288 1807 292
rect 1811 288 1812 292
rect 1806 287 1812 288
rect 2222 291 2228 292
rect 2222 287 2223 291
rect 2227 287 2228 291
rect 2222 286 2228 287
rect 2310 291 2316 292
rect 2310 287 2311 291
rect 2315 287 2316 291
rect 2310 286 2316 287
rect 2398 291 2404 292
rect 2398 287 2399 291
rect 2403 287 2404 291
rect 2398 286 2404 287
rect 2486 291 2492 292
rect 2486 287 2487 291
rect 2491 287 2492 291
rect 2486 286 2492 287
rect 2574 291 2580 292
rect 2574 287 2575 291
rect 2579 287 2580 291
rect 2574 286 2580 287
rect 2678 291 2684 292
rect 2678 287 2679 291
rect 2683 287 2684 291
rect 2678 286 2684 287
rect 2798 291 2804 292
rect 2798 287 2799 291
rect 2803 287 2804 291
rect 2798 286 2804 287
rect 2926 291 2932 292
rect 2926 287 2927 291
rect 2931 287 2932 291
rect 2926 286 2932 287
rect 3070 291 3076 292
rect 3070 287 3071 291
rect 3075 287 3076 291
rect 3070 286 3076 287
rect 3222 291 3228 292
rect 3222 287 3223 291
rect 3227 287 3228 291
rect 3222 286 3228 287
rect 3366 291 3372 292
rect 3366 287 3367 291
rect 3371 287 3372 291
rect 3462 288 3463 292
rect 3467 288 3468 292
rect 3462 287 3468 288
rect 3366 286 3372 287
rect 1766 283 1772 284
rect 2294 283 2300 284
rect 1238 282 1244 283
rect 900 276 961 278
rect 1097 276 1114 278
rect 1198 279 1204 280
rect 900 275 901 276
rect 895 274 901 275
rect 1198 275 1199 279
rect 1203 275 1204 279
rect 2294 279 2295 283
rect 2299 279 2300 283
rect 2294 278 2300 279
rect 2382 283 2388 284
rect 2382 279 2383 283
rect 2387 279 2388 283
rect 2382 278 2388 279
rect 2470 283 2476 284
rect 2470 279 2471 283
rect 2475 279 2476 283
rect 2470 278 2476 279
rect 2478 283 2484 284
rect 2478 279 2479 283
rect 2483 282 2484 283
rect 2566 283 2572 284
rect 2483 280 2529 282
rect 2483 279 2484 280
rect 2478 278 2484 279
rect 2566 279 2567 283
rect 2571 282 2572 283
rect 2750 283 2756 284
rect 2571 280 2617 282
rect 2571 279 2572 280
rect 2566 278 2572 279
rect 2750 279 2751 283
rect 2755 279 2756 283
rect 2750 278 2756 279
rect 2870 283 2876 284
rect 2870 279 2871 283
rect 2875 279 2876 283
rect 2870 278 2876 279
rect 2998 283 3004 284
rect 2998 279 2999 283
rect 3003 279 3004 283
rect 2998 278 3004 279
rect 3142 283 3148 284
rect 3142 279 3143 283
rect 3147 279 3148 283
rect 3142 278 3148 279
rect 3150 283 3156 284
rect 3150 279 3151 283
rect 3155 282 3156 283
rect 3155 280 3265 282
rect 3155 279 3156 280
rect 3150 278 3156 279
rect 3438 279 3444 280
rect 1198 274 1204 275
rect 1318 275 1324 276
rect 1318 274 1319 275
rect 1313 272 1319 274
rect 782 270 788 271
rect 1318 271 1319 272
rect 1323 271 1324 275
rect 1806 275 1812 276
rect 1318 270 1324 271
rect 1766 271 1772 272
rect 110 266 116 267
rect 262 268 268 269
rect 262 264 263 268
rect 267 264 268 268
rect 262 263 268 264
rect 374 268 380 269
rect 374 264 375 268
rect 379 264 380 268
rect 374 263 380 264
rect 486 268 492 269
rect 486 264 487 268
rect 491 264 492 268
rect 486 263 492 264
rect 598 268 604 269
rect 598 264 599 268
rect 603 264 604 268
rect 598 263 604 264
rect 710 268 716 269
rect 710 264 711 268
rect 715 264 716 268
rect 710 263 716 264
rect 814 268 820 269
rect 814 264 815 268
rect 819 264 820 268
rect 814 263 820 264
rect 918 268 924 269
rect 918 264 919 268
rect 923 264 924 268
rect 918 263 924 264
rect 1022 268 1028 269
rect 1022 264 1023 268
rect 1027 264 1028 268
rect 1022 263 1028 264
rect 1126 268 1132 269
rect 1126 264 1127 268
rect 1131 264 1132 268
rect 1126 263 1132 264
rect 1238 268 1244 269
rect 1238 264 1239 268
rect 1243 264 1244 268
rect 1766 267 1767 271
rect 1771 267 1772 271
rect 1806 271 1807 275
rect 1811 271 1812 275
rect 3438 275 3439 279
rect 3443 275 3444 279
rect 3438 274 3444 275
rect 3462 275 3468 276
rect 1806 270 1812 271
rect 2222 272 2228 273
rect 2222 268 2223 272
rect 2227 268 2228 272
rect 2222 267 2228 268
rect 2310 272 2316 273
rect 2310 268 2311 272
rect 2315 268 2316 272
rect 2310 267 2316 268
rect 2398 272 2404 273
rect 2398 268 2399 272
rect 2403 268 2404 272
rect 2398 267 2404 268
rect 2486 272 2492 273
rect 2486 268 2487 272
rect 2491 268 2492 272
rect 2486 267 2492 268
rect 2574 272 2580 273
rect 2574 268 2575 272
rect 2579 268 2580 272
rect 2574 267 2580 268
rect 2678 272 2684 273
rect 2678 268 2679 272
rect 2683 268 2684 272
rect 2678 267 2684 268
rect 2798 272 2804 273
rect 2798 268 2799 272
rect 2803 268 2804 272
rect 2798 267 2804 268
rect 2926 272 2932 273
rect 2926 268 2927 272
rect 2931 268 2932 272
rect 2926 267 2932 268
rect 3070 272 3076 273
rect 3070 268 3071 272
rect 3075 268 3076 272
rect 3070 267 3076 268
rect 3222 272 3228 273
rect 3222 268 3223 272
rect 3227 268 3228 272
rect 3222 267 3228 268
rect 3366 272 3372 273
rect 3366 268 3367 272
rect 3371 268 3372 272
rect 3462 271 3463 275
rect 3467 271 3468 275
rect 3462 270 3468 271
rect 3366 267 3372 268
rect 1766 266 1772 267
rect 1238 263 1244 264
rect 2274 263 2280 264
rect 2274 259 2275 263
rect 2279 262 2280 263
rect 2478 263 2484 264
rect 2478 262 2479 263
rect 2279 260 2479 262
rect 2279 259 2280 260
rect 2274 258 2280 259
rect 2478 259 2479 260
rect 2483 259 2484 263
rect 2478 258 2484 259
rect 446 220 452 221
rect 110 217 116 218
rect 110 213 111 217
rect 115 213 116 217
rect 446 216 447 220
rect 451 216 452 220
rect 446 215 452 216
rect 534 220 540 221
rect 534 216 535 220
rect 539 216 540 220
rect 534 215 540 216
rect 622 220 628 221
rect 622 216 623 220
rect 627 216 628 220
rect 622 215 628 216
rect 710 220 716 221
rect 710 216 711 220
rect 715 216 716 220
rect 710 215 716 216
rect 806 220 812 221
rect 806 216 807 220
rect 811 216 812 220
rect 806 215 812 216
rect 902 220 908 221
rect 902 216 903 220
rect 907 216 908 220
rect 902 215 908 216
rect 998 220 1004 221
rect 998 216 999 220
rect 1003 216 1004 220
rect 998 215 1004 216
rect 1102 220 1108 221
rect 1102 216 1103 220
rect 1107 216 1108 220
rect 1102 215 1108 216
rect 1206 220 1212 221
rect 1206 216 1207 220
rect 1211 216 1212 220
rect 1206 215 1212 216
rect 1310 220 1316 221
rect 1310 216 1311 220
rect 1315 216 1316 220
rect 2142 220 2148 221
rect 1310 215 1316 216
rect 1766 217 1772 218
rect 110 212 116 213
rect 1766 213 1767 217
rect 1771 213 1772 217
rect 1766 212 1772 213
rect 1806 217 1812 218
rect 1806 213 1807 217
rect 1811 213 1812 217
rect 2142 216 2143 220
rect 2147 216 2148 220
rect 2142 215 2148 216
rect 2262 220 2268 221
rect 2262 216 2263 220
rect 2267 216 2268 220
rect 2262 215 2268 216
rect 2382 220 2388 221
rect 2382 216 2383 220
rect 2387 216 2388 220
rect 2382 215 2388 216
rect 2510 220 2516 221
rect 2510 216 2511 220
rect 2515 216 2516 220
rect 2510 215 2516 216
rect 2638 220 2644 221
rect 2638 216 2639 220
rect 2643 216 2644 220
rect 2638 215 2644 216
rect 2766 220 2772 221
rect 2766 216 2767 220
rect 2771 216 2772 220
rect 2766 215 2772 216
rect 2894 220 2900 221
rect 2894 216 2895 220
rect 2899 216 2900 220
rect 2894 215 2900 216
rect 3014 220 3020 221
rect 3014 216 3015 220
rect 3019 216 3020 220
rect 3014 215 3020 216
rect 3134 220 3140 221
rect 3134 216 3135 220
rect 3139 216 3140 220
rect 3134 215 3140 216
rect 3262 220 3268 221
rect 3262 216 3263 220
rect 3267 216 3268 220
rect 3262 215 3268 216
rect 3366 220 3372 221
rect 3366 216 3367 220
rect 3371 216 3372 220
rect 3366 215 3372 216
rect 3462 217 3468 218
rect 1806 212 1812 213
rect 3462 213 3463 217
rect 3467 213 3468 217
rect 3462 212 3468 213
rect 314 211 320 212
rect 314 207 315 211
rect 319 210 320 211
rect 526 211 532 212
rect 319 208 489 210
rect 319 207 320 208
rect 314 206 320 207
rect 526 207 527 211
rect 531 210 532 211
rect 694 211 700 212
rect 531 208 577 210
rect 531 207 532 208
rect 526 206 532 207
rect 694 207 695 211
rect 699 207 700 211
rect 694 206 700 207
rect 774 211 780 212
rect 774 207 775 211
rect 779 207 780 211
rect 774 206 780 207
rect 878 211 884 212
rect 878 207 879 211
rect 883 207 884 211
rect 878 206 884 207
rect 886 211 892 212
rect 886 207 887 211
rect 891 210 892 211
rect 982 211 988 212
rect 891 208 945 210
rect 891 207 892 208
rect 886 206 892 207
rect 982 207 983 211
rect 987 210 988 211
rect 1079 211 1085 212
rect 987 208 1041 210
rect 987 207 988 208
rect 982 206 988 207
rect 1079 207 1080 211
rect 1084 210 1085 211
rect 1199 211 1205 212
rect 1084 208 1145 210
rect 1084 207 1085 208
rect 1079 206 1085 207
rect 1199 207 1200 211
rect 1204 210 1205 211
rect 1286 211 1292 212
rect 1204 208 1249 210
rect 1204 207 1205 208
rect 1199 206 1205 207
rect 1286 207 1287 211
rect 1291 210 1292 211
rect 2214 211 2220 212
rect 1291 208 1353 210
rect 1291 207 1292 208
rect 1286 206 1292 207
rect 2214 207 2215 211
rect 2219 207 2220 211
rect 2214 206 2220 207
rect 2334 211 2340 212
rect 2334 207 2335 211
rect 2339 207 2340 211
rect 2334 206 2340 207
rect 2454 211 2460 212
rect 2454 207 2455 211
rect 2459 207 2460 211
rect 2454 206 2460 207
rect 2582 211 2588 212
rect 2582 207 2583 211
rect 2587 207 2588 211
rect 2582 206 2588 207
rect 2626 211 2632 212
rect 2626 207 2627 211
rect 2631 210 2632 211
rect 2719 211 2725 212
rect 2631 208 2681 210
rect 2631 207 2632 208
rect 2626 206 2632 207
rect 2719 207 2720 211
rect 2724 210 2725 211
rect 2871 211 2877 212
rect 2724 208 2809 210
rect 2724 207 2725 208
rect 2719 206 2725 207
rect 2871 207 2872 211
rect 2876 210 2877 211
rect 2974 211 2980 212
rect 2876 208 2937 210
rect 2876 207 2877 208
rect 2871 206 2877 207
rect 2974 207 2975 211
rect 2979 210 2980 211
rect 3206 211 3212 212
rect 2979 208 3057 210
rect 2979 207 2980 208
rect 2974 206 2980 207
rect 3206 207 3207 211
rect 3211 207 3212 211
rect 3342 211 3348 212
rect 3342 210 3343 211
rect 3337 208 3343 210
rect 3206 206 3212 207
rect 3342 207 3343 208
rect 3347 207 3348 211
rect 3342 206 3348 207
rect 3430 211 3436 212
rect 3430 207 3431 211
rect 3435 207 3436 211
rect 3430 206 3436 207
rect 446 201 452 202
rect 110 200 116 201
rect 110 196 111 200
rect 115 196 116 200
rect 446 197 447 201
rect 451 197 452 201
rect 446 196 452 197
rect 534 201 540 202
rect 534 197 535 201
rect 539 197 540 201
rect 534 196 540 197
rect 622 201 628 202
rect 622 197 623 201
rect 627 197 628 201
rect 622 196 628 197
rect 710 201 716 202
rect 710 197 711 201
rect 715 197 716 201
rect 710 196 716 197
rect 806 201 812 202
rect 806 197 807 201
rect 811 197 812 201
rect 806 196 812 197
rect 902 201 908 202
rect 902 197 903 201
rect 907 197 908 201
rect 902 196 908 197
rect 998 201 1004 202
rect 998 197 999 201
rect 1003 197 1004 201
rect 998 196 1004 197
rect 1102 201 1108 202
rect 1102 197 1103 201
rect 1107 197 1108 201
rect 1102 196 1108 197
rect 1206 201 1212 202
rect 1206 197 1207 201
rect 1211 197 1212 201
rect 1206 196 1212 197
rect 1310 201 1316 202
rect 2142 201 2148 202
rect 1310 197 1311 201
rect 1315 197 1316 201
rect 1310 196 1316 197
rect 1766 200 1772 201
rect 1766 196 1767 200
rect 1771 196 1772 200
rect 110 195 116 196
rect 1766 195 1772 196
rect 1806 200 1812 201
rect 1806 196 1807 200
rect 1811 196 1812 200
rect 2142 197 2143 201
rect 2147 197 2148 201
rect 2142 196 2148 197
rect 2262 201 2268 202
rect 2262 197 2263 201
rect 2267 197 2268 201
rect 2262 196 2268 197
rect 2382 201 2388 202
rect 2382 197 2383 201
rect 2387 197 2388 201
rect 2382 196 2388 197
rect 2510 201 2516 202
rect 2510 197 2511 201
rect 2515 197 2516 201
rect 2510 196 2516 197
rect 2638 201 2644 202
rect 2638 197 2639 201
rect 2643 197 2644 201
rect 2638 196 2644 197
rect 2766 201 2772 202
rect 2766 197 2767 201
rect 2771 197 2772 201
rect 2766 196 2772 197
rect 2894 201 2900 202
rect 2894 197 2895 201
rect 2899 197 2900 201
rect 2894 196 2900 197
rect 3014 201 3020 202
rect 3014 197 3015 201
rect 3019 197 3020 201
rect 3014 196 3020 197
rect 3134 201 3140 202
rect 3134 197 3135 201
rect 3139 197 3140 201
rect 3134 196 3140 197
rect 3262 201 3268 202
rect 3262 197 3263 201
rect 3267 197 3268 201
rect 3262 196 3268 197
rect 3366 201 3372 202
rect 3366 197 3367 201
rect 3371 197 3372 201
rect 3366 196 3372 197
rect 3462 200 3468 201
rect 3462 196 3463 200
rect 3467 196 3468 200
rect 1806 195 1812 196
rect 3462 195 3468 196
rect 495 183 501 184
rect 495 179 496 183
rect 500 182 501 183
rect 526 183 532 184
rect 526 182 527 183
rect 500 180 527 182
rect 500 179 501 180
rect 495 178 501 179
rect 526 179 527 180
rect 531 179 532 183
rect 526 178 532 179
rect 583 183 592 184
rect 583 179 584 183
rect 591 179 592 183
rect 583 178 592 179
rect 671 183 677 184
rect 671 179 672 183
rect 676 182 677 183
rect 694 183 700 184
rect 676 180 690 182
rect 676 179 677 180
rect 671 178 677 179
rect 688 174 690 180
rect 694 179 695 183
rect 699 182 700 183
rect 759 183 765 184
rect 759 182 760 183
rect 699 180 760 182
rect 699 179 700 180
rect 694 178 700 179
rect 759 179 760 180
rect 764 179 765 183
rect 759 178 765 179
rect 782 183 788 184
rect 782 179 783 183
rect 787 182 788 183
rect 855 183 861 184
rect 855 182 856 183
rect 787 180 856 182
rect 787 179 788 180
rect 782 178 788 179
rect 855 179 856 180
rect 860 179 861 183
rect 886 183 892 184
rect 886 182 887 183
rect 855 178 861 179
rect 864 180 887 182
rect 864 174 866 180
rect 886 179 887 180
rect 891 179 892 183
rect 886 178 892 179
rect 950 183 957 184
rect 950 179 951 183
rect 956 179 957 183
rect 1047 183 1053 184
rect 1047 182 1048 183
rect 950 178 957 179
rect 960 180 1048 182
rect 688 172 866 174
rect 878 175 884 176
rect 878 171 879 175
rect 883 174 884 175
rect 960 174 962 180
rect 1047 179 1048 180
rect 1052 179 1053 183
rect 1047 178 1053 179
rect 1151 183 1157 184
rect 1151 179 1152 183
rect 1156 182 1157 183
rect 1199 183 1205 184
rect 1199 182 1200 183
rect 1156 180 1200 182
rect 1156 179 1157 180
rect 1151 178 1157 179
rect 1199 179 1200 180
rect 1204 179 1205 183
rect 1199 178 1205 179
rect 1255 183 1261 184
rect 1255 179 1256 183
rect 1260 182 1261 183
rect 1286 183 1292 184
rect 1286 182 1287 183
rect 1260 180 1287 182
rect 1260 179 1261 180
rect 1255 178 1261 179
rect 1286 179 1287 180
rect 1291 179 1292 183
rect 1286 178 1292 179
rect 1318 183 1324 184
rect 1318 179 1319 183
rect 1323 182 1324 183
rect 1359 183 1365 184
rect 1359 182 1360 183
rect 1323 180 1360 182
rect 1323 179 1324 180
rect 1318 178 1324 179
rect 1359 179 1360 180
rect 1364 179 1365 183
rect 1359 178 1365 179
rect 2191 183 2197 184
rect 2191 179 2192 183
rect 2196 182 2197 183
rect 2214 183 2220 184
rect 2196 180 2211 182
rect 2196 179 2197 180
rect 2191 178 2197 179
rect 883 172 962 174
rect 2209 174 2211 180
rect 2214 179 2215 183
rect 2219 182 2220 183
rect 2311 183 2317 184
rect 2311 182 2312 183
rect 2219 180 2312 182
rect 2219 179 2220 180
rect 2214 178 2220 179
rect 2311 179 2312 180
rect 2316 179 2317 183
rect 2311 178 2317 179
rect 2334 183 2340 184
rect 2334 179 2335 183
rect 2339 182 2340 183
rect 2431 183 2437 184
rect 2431 182 2432 183
rect 2339 180 2432 182
rect 2339 179 2340 180
rect 2334 178 2340 179
rect 2431 179 2432 180
rect 2436 179 2437 183
rect 2431 178 2437 179
rect 2454 183 2460 184
rect 2454 179 2455 183
rect 2459 182 2460 183
rect 2559 183 2565 184
rect 2559 182 2560 183
rect 2459 180 2560 182
rect 2459 179 2460 180
rect 2454 178 2460 179
rect 2559 179 2560 180
rect 2564 179 2565 183
rect 2559 178 2565 179
rect 2582 183 2588 184
rect 2582 179 2583 183
rect 2587 182 2588 183
rect 2687 183 2693 184
rect 2687 182 2688 183
rect 2587 180 2688 182
rect 2587 179 2588 180
rect 2582 178 2588 179
rect 2687 179 2688 180
rect 2692 179 2693 183
rect 2687 178 2693 179
rect 2815 183 2821 184
rect 2815 179 2816 183
rect 2820 182 2821 183
rect 2871 183 2877 184
rect 2871 182 2872 183
rect 2820 180 2872 182
rect 2820 179 2821 180
rect 2815 178 2821 179
rect 2871 179 2872 180
rect 2876 179 2877 183
rect 2871 178 2877 179
rect 2943 183 2949 184
rect 2943 179 2944 183
rect 2948 182 2949 183
rect 2974 183 2980 184
rect 2974 182 2975 183
rect 2948 180 2975 182
rect 2948 179 2949 180
rect 2943 178 2949 179
rect 2974 179 2975 180
rect 2979 179 2980 183
rect 2974 178 2980 179
rect 3063 183 3069 184
rect 3063 179 3064 183
rect 3068 182 3069 183
rect 3150 183 3156 184
rect 3150 182 3151 183
rect 3068 180 3151 182
rect 3068 179 3069 180
rect 3063 178 3069 179
rect 3150 179 3151 180
rect 3155 179 3156 183
rect 3150 178 3156 179
rect 3182 183 3189 184
rect 3182 179 3183 183
rect 3188 179 3189 183
rect 3182 178 3189 179
rect 3206 183 3212 184
rect 3206 179 3207 183
rect 3211 182 3212 183
rect 3311 183 3317 184
rect 3311 182 3312 183
rect 3211 180 3312 182
rect 3211 179 3212 180
rect 3206 178 3212 179
rect 3311 179 3312 180
rect 3316 179 3317 183
rect 3311 178 3317 179
rect 3415 183 3421 184
rect 3415 179 3416 183
rect 3420 182 3421 183
rect 3438 183 3444 184
rect 3438 182 3439 183
rect 3420 180 3439 182
rect 3420 179 3421 180
rect 3415 178 3421 179
rect 3438 179 3439 180
rect 3443 179 3444 183
rect 3438 178 3444 179
rect 2374 175 2380 176
rect 2374 174 2375 175
rect 2209 172 2375 174
rect 883 171 884 172
rect 878 170 884 171
rect 2374 171 2375 172
rect 2379 171 2380 175
rect 2374 170 2380 171
rect 2719 155 2725 156
rect 2719 154 2720 155
rect 2576 152 2720 154
rect 1079 151 1085 152
rect 1079 150 1080 151
rect 1032 148 1080 150
rect 311 143 320 144
rect 311 139 312 143
rect 319 139 320 143
rect 311 138 320 139
rect 334 143 340 144
rect 334 139 335 143
rect 339 142 340 143
rect 399 143 405 144
rect 399 142 400 143
rect 339 140 400 142
rect 339 139 340 140
rect 334 138 340 139
rect 399 139 400 140
rect 404 139 405 143
rect 399 138 405 139
rect 422 143 428 144
rect 422 139 423 143
rect 427 142 428 143
rect 487 143 493 144
rect 487 142 488 143
rect 427 140 488 142
rect 427 139 428 140
rect 422 138 428 139
rect 487 139 488 140
rect 492 139 493 143
rect 487 138 493 139
rect 510 143 516 144
rect 510 139 511 143
rect 515 142 516 143
rect 575 143 581 144
rect 575 142 576 143
rect 515 140 576 142
rect 515 139 516 140
rect 510 138 516 139
rect 575 139 576 140
rect 580 139 581 143
rect 575 138 581 139
rect 598 143 604 144
rect 598 139 599 143
rect 603 142 604 143
rect 663 143 669 144
rect 663 142 664 143
rect 603 140 664 142
rect 603 139 604 140
rect 598 138 604 139
rect 663 139 664 140
rect 668 139 669 143
rect 663 138 669 139
rect 686 143 692 144
rect 686 139 687 143
rect 691 142 692 143
rect 751 143 757 144
rect 751 142 752 143
rect 691 140 752 142
rect 691 139 692 140
rect 686 138 692 139
rect 751 139 752 140
rect 756 139 757 143
rect 751 138 757 139
rect 774 143 780 144
rect 774 139 775 143
rect 779 142 780 143
rect 839 143 845 144
rect 839 142 840 143
rect 779 140 840 142
rect 779 139 780 140
rect 774 138 780 139
rect 839 139 840 140
rect 844 139 845 143
rect 839 138 845 139
rect 862 143 868 144
rect 862 139 863 143
rect 867 142 868 143
rect 927 143 933 144
rect 927 142 928 143
rect 867 140 928 142
rect 867 139 868 140
rect 862 138 868 139
rect 927 139 928 140
rect 932 139 933 143
rect 927 138 933 139
rect 1015 143 1021 144
rect 1015 139 1016 143
rect 1020 142 1021 143
rect 1032 142 1034 148
rect 1079 147 1080 148
rect 1084 147 1085 151
rect 1079 146 1085 147
rect 1742 147 1748 148
rect 1020 140 1034 142
rect 1038 143 1044 144
rect 1020 139 1021 140
rect 1015 138 1021 139
rect 1038 139 1039 143
rect 1043 142 1044 143
rect 1103 143 1109 144
rect 1103 142 1104 143
rect 1043 140 1104 142
rect 1043 139 1044 140
rect 1038 138 1044 139
rect 1103 139 1104 140
rect 1108 139 1109 143
rect 1103 138 1109 139
rect 1126 143 1132 144
rect 1126 139 1127 143
rect 1131 142 1132 143
rect 1191 143 1197 144
rect 1191 142 1192 143
rect 1131 140 1192 142
rect 1131 139 1132 140
rect 1126 138 1132 139
rect 1191 139 1192 140
rect 1196 139 1197 143
rect 1191 138 1197 139
rect 1214 143 1220 144
rect 1214 139 1215 143
rect 1219 142 1220 143
rect 1279 143 1285 144
rect 1279 142 1280 143
rect 1219 140 1280 142
rect 1219 139 1220 140
rect 1214 138 1220 139
rect 1279 139 1280 140
rect 1284 139 1285 143
rect 1279 138 1285 139
rect 1302 143 1308 144
rect 1302 139 1303 143
rect 1307 142 1308 143
rect 1367 143 1373 144
rect 1367 142 1368 143
rect 1307 140 1368 142
rect 1307 139 1308 140
rect 1302 138 1308 139
rect 1367 139 1368 140
rect 1372 139 1373 143
rect 1367 138 1373 139
rect 1390 143 1396 144
rect 1390 139 1391 143
rect 1395 142 1396 143
rect 1455 143 1461 144
rect 1455 142 1456 143
rect 1395 140 1456 142
rect 1395 139 1396 140
rect 1390 138 1396 139
rect 1455 139 1456 140
rect 1460 139 1461 143
rect 1455 138 1461 139
rect 1478 143 1484 144
rect 1478 139 1479 143
rect 1483 142 1484 143
rect 1543 143 1549 144
rect 1543 142 1544 143
rect 1483 140 1544 142
rect 1483 139 1484 140
rect 1478 138 1484 139
rect 1543 139 1544 140
rect 1548 139 1549 143
rect 1543 138 1549 139
rect 1566 143 1572 144
rect 1566 139 1567 143
rect 1571 142 1572 143
rect 1631 143 1637 144
rect 1631 142 1632 143
rect 1571 140 1632 142
rect 1571 139 1572 140
rect 1566 138 1572 139
rect 1631 139 1632 140
rect 1636 139 1637 143
rect 1631 138 1637 139
rect 1654 143 1660 144
rect 1654 139 1655 143
rect 1659 142 1660 143
rect 1719 143 1725 144
rect 1719 142 1720 143
rect 1659 140 1720 142
rect 1659 139 1660 140
rect 1654 138 1660 139
rect 1719 139 1720 140
rect 1724 139 1725 143
rect 1742 143 1743 147
rect 1747 146 1748 147
rect 1879 147 1885 148
rect 1879 146 1880 147
rect 1747 144 1880 146
rect 1747 143 1748 144
rect 1742 142 1748 143
rect 1879 143 1880 144
rect 1884 143 1885 147
rect 1879 142 1885 143
rect 1902 147 1908 148
rect 1902 143 1903 147
rect 1907 146 1908 147
rect 1967 147 1973 148
rect 1967 146 1968 147
rect 1907 144 1968 146
rect 1907 143 1908 144
rect 1902 142 1908 143
rect 1967 143 1968 144
rect 1972 143 1973 147
rect 1967 142 1973 143
rect 1990 147 1996 148
rect 1990 143 1991 147
rect 1995 146 1996 147
rect 2055 147 2061 148
rect 2055 146 2056 147
rect 1995 144 2056 146
rect 1995 143 1996 144
rect 1990 142 1996 143
rect 2055 143 2056 144
rect 2060 143 2061 147
rect 2055 142 2061 143
rect 2078 147 2084 148
rect 2078 143 2079 147
rect 2083 146 2084 147
rect 2143 147 2149 148
rect 2143 146 2144 147
rect 2083 144 2144 146
rect 2083 143 2084 144
rect 2078 142 2084 143
rect 2143 143 2144 144
rect 2148 143 2149 147
rect 2143 142 2149 143
rect 2166 147 2172 148
rect 2166 143 2167 147
rect 2171 146 2172 147
rect 2231 147 2237 148
rect 2231 146 2232 147
rect 2171 144 2232 146
rect 2171 143 2172 144
rect 2166 142 2172 143
rect 2231 143 2232 144
rect 2236 143 2237 147
rect 2231 142 2237 143
rect 2254 147 2260 148
rect 2254 143 2255 147
rect 2259 146 2260 147
rect 2343 147 2349 148
rect 2343 146 2344 147
rect 2259 144 2344 146
rect 2259 143 2260 144
rect 2254 142 2260 143
rect 2343 143 2344 144
rect 2348 143 2349 147
rect 2343 142 2349 143
rect 2366 147 2372 148
rect 2366 143 2367 147
rect 2371 146 2372 147
rect 2455 147 2461 148
rect 2455 146 2456 147
rect 2371 144 2456 146
rect 2371 143 2372 144
rect 2366 142 2372 143
rect 2455 143 2456 144
rect 2460 143 2461 147
rect 2455 142 2461 143
rect 2559 147 2565 148
rect 2559 143 2560 147
rect 2564 146 2565 147
rect 2576 146 2578 152
rect 2719 151 2720 152
rect 2724 151 2725 155
rect 2719 150 2725 151
rect 2564 144 2578 146
rect 2582 147 2588 148
rect 2564 143 2565 144
rect 2559 142 2565 143
rect 2582 143 2583 147
rect 2587 146 2588 147
rect 2663 147 2669 148
rect 2663 146 2664 147
rect 2587 144 2664 146
rect 2587 143 2588 144
rect 2582 142 2588 143
rect 2663 143 2664 144
rect 2668 143 2669 147
rect 2663 142 2669 143
rect 2686 147 2692 148
rect 2686 143 2687 147
rect 2691 146 2692 147
rect 2767 147 2773 148
rect 2767 146 2768 147
rect 2691 144 2768 146
rect 2691 143 2692 144
rect 2686 142 2692 143
rect 2767 143 2768 144
rect 2772 143 2773 147
rect 2767 142 2773 143
rect 2790 147 2796 148
rect 2790 143 2791 147
rect 2795 146 2796 147
rect 2863 147 2869 148
rect 2863 146 2864 147
rect 2795 144 2864 146
rect 2795 143 2796 144
rect 2790 142 2796 143
rect 2863 143 2864 144
rect 2868 143 2869 147
rect 2863 142 2869 143
rect 2886 147 2892 148
rect 2886 143 2887 147
rect 2891 146 2892 147
rect 2959 147 2965 148
rect 2959 146 2960 147
rect 2891 144 2960 146
rect 2891 143 2892 144
rect 2886 142 2892 143
rect 2959 143 2960 144
rect 2964 143 2965 147
rect 2959 142 2965 143
rect 2982 147 2988 148
rect 2982 143 2983 147
rect 2987 146 2988 147
rect 3055 147 3061 148
rect 3055 146 3056 147
rect 2987 144 3056 146
rect 2987 143 2988 144
rect 2982 142 2988 143
rect 3055 143 3056 144
rect 3060 143 3061 147
rect 3055 142 3061 143
rect 3078 147 3084 148
rect 3078 143 3079 147
rect 3083 146 3084 147
rect 3151 147 3157 148
rect 3151 146 3152 147
rect 3083 144 3152 146
rect 3083 143 3084 144
rect 3078 142 3084 143
rect 3151 143 3152 144
rect 3156 143 3157 147
rect 3151 142 3157 143
rect 3174 147 3180 148
rect 3174 143 3175 147
rect 3179 146 3180 147
rect 3239 147 3245 148
rect 3239 146 3240 147
rect 3179 144 3240 146
rect 3179 143 3180 144
rect 3174 142 3180 143
rect 3239 143 3240 144
rect 3244 143 3245 147
rect 3239 142 3245 143
rect 3327 147 3333 148
rect 3327 143 3328 147
rect 3332 146 3333 147
rect 3358 147 3364 148
rect 3358 146 3359 147
rect 3332 144 3359 146
rect 3332 143 3333 144
rect 3327 142 3333 143
rect 3358 143 3359 144
rect 3363 143 3364 147
rect 3358 142 3364 143
rect 3415 147 3421 148
rect 3415 143 3416 147
rect 3420 146 3421 147
rect 3430 147 3436 148
rect 3430 146 3431 147
rect 3420 144 3431 146
rect 3420 143 3421 144
rect 3415 142 3421 143
rect 3430 143 3431 144
rect 3435 143 3436 147
rect 3430 142 3436 143
rect 1719 138 1725 139
rect 1806 132 1812 133
rect 3462 132 3468 133
rect 110 128 116 129
rect 1766 128 1772 129
rect 110 124 111 128
rect 115 124 116 128
rect 110 123 116 124
rect 262 127 268 128
rect 262 123 263 127
rect 267 123 268 127
rect 262 122 268 123
rect 350 127 356 128
rect 350 123 351 127
rect 355 123 356 127
rect 350 122 356 123
rect 438 127 444 128
rect 438 123 439 127
rect 443 123 444 127
rect 438 122 444 123
rect 526 127 532 128
rect 526 123 527 127
rect 531 123 532 127
rect 526 122 532 123
rect 614 127 620 128
rect 614 123 615 127
rect 619 123 620 127
rect 614 122 620 123
rect 702 127 708 128
rect 702 123 703 127
rect 707 123 708 127
rect 702 122 708 123
rect 790 127 796 128
rect 790 123 791 127
rect 795 123 796 127
rect 790 122 796 123
rect 878 127 884 128
rect 878 123 879 127
rect 883 123 884 127
rect 878 122 884 123
rect 966 127 972 128
rect 966 123 967 127
rect 971 123 972 127
rect 966 122 972 123
rect 1054 127 1060 128
rect 1054 123 1055 127
rect 1059 123 1060 127
rect 1054 122 1060 123
rect 1142 127 1148 128
rect 1142 123 1143 127
rect 1147 123 1148 127
rect 1142 122 1148 123
rect 1230 127 1236 128
rect 1230 123 1231 127
rect 1235 123 1236 127
rect 1230 122 1236 123
rect 1318 127 1324 128
rect 1318 123 1319 127
rect 1323 123 1324 127
rect 1318 122 1324 123
rect 1406 127 1412 128
rect 1406 123 1407 127
rect 1411 123 1412 127
rect 1406 122 1412 123
rect 1494 127 1500 128
rect 1494 123 1495 127
rect 1499 123 1500 127
rect 1494 122 1500 123
rect 1582 127 1588 128
rect 1582 123 1583 127
rect 1587 123 1588 127
rect 1582 122 1588 123
rect 1670 127 1676 128
rect 1670 123 1671 127
rect 1675 123 1676 127
rect 1766 124 1767 128
rect 1771 124 1772 128
rect 1806 128 1807 132
rect 1811 128 1812 132
rect 1806 127 1812 128
rect 1830 131 1836 132
rect 1830 127 1831 131
rect 1835 127 1836 131
rect 1830 126 1836 127
rect 1918 131 1924 132
rect 1918 127 1919 131
rect 1923 127 1924 131
rect 1918 126 1924 127
rect 2006 131 2012 132
rect 2006 127 2007 131
rect 2011 127 2012 131
rect 2006 126 2012 127
rect 2094 131 2100 132
rect 2094 127 2095 131
rect 2099 127 2100 131
rect 2094 126 2100 127
rect 2182 131 2188 132
rect 2182 127 2183 131
rect 2187 127 2188 131
rect 2182 126 2188 127
rect 2294 131 2300 132
rect 2294 127 2295 131
rect 2299 127 2300 131
rect 2294 126 2300 127
rect 2406 131 2412 132
rect 2406 127 2407 131
rect 2411 127 2412 131
rect 2406 126 2412 127
rect 2510 131 2516 132
rect 2510 127 2511 131
rect 2515 127 2516 131
rect 2510 126 2516 127
rect 2614 131 2620 132
rect 2614 127 2615 131
rect 2619 127 2620 131
rect 2614 126 2620 127
rect 2718 131 2724 132
rect 2718 127 2719 131
rect 2723 127 2724 131
rect 2718 126 2724 127
rect 2814 131 2820 132
rect 2814 127 2815 131
rect 2819 127 2820 131
rect 2814 126 2820 127
rect 2910 131 2916 132
rect 2910 127 2911 131
rect 2915 127 2916 131
rect 2910 126 2916 127
rect 3006 131 3012 132
rect 3006 127 3007 131
rect 3011 127 3012 131
rect 3006 126 3012 127
rect 3102 131 3108 132
rect 3102 127 3103 131
rect 3107 127 3108 131
rect 3102 126 3108 127
rect 3190 131 3196 132
rect 3190 127 3191 131
rect 3195 127 3196 131
rect 3190 126 3196 127
rect 3278 131 3284 132
rect 3278 127 3279 131
rect 3283 127 3284 131
rect 3278 126 3284 127
rect 3366 131 3372 132
rect 3366 127 3367 131
rect 3371 127 3372 131
rect 3462 128 3463 132
rect 3467 128 3468 132
rect 3462 127 3468 128
rect 3366 126 3372 127
rect 1766 123 1772 124
rect 1902 123 1908 124
rect 1670 122 1676 123
rect 334 119 340 120
rect 334 115 335 119
rect 339 115 340 119
rect 334 114 340 115
rect 422 119 428 120
rect 422 115 423 119
rect 427 115 428 119
rect 422 114 428 115
rect 510 119 516 120
rect 510 115 511 119
rect 515 115 516 119
rect 510 114 516 115
rect 598 119 604 120
rect 598 115 599 119
rect 603 115 604 119
rect 598 114 604 115
rect 686 119 692 120
rect 686 115 687 119
rect 691 115 692 119
rect 686 114 692 115
rect 774 119 780 120
rect 774 115 775 119
rect 779 115 780 119
rect 774 114 780 115
rect 862 119 868 120
rect 862 115 863 119
rect 867 115 868 119
rect 862 114 868 115
rect 950 119 956 120
rect 950 115 951 119
rect 955 115 956 119
rect 950 114 956 115
rect 1038 119 1044 120
rect 1038 115 1039 119
rect 1043 115 1044 119
rect 1038 114 1044 115
rect 1126 119 1132 120
rect 1126 115 1127 119
rect 1131 115 1132 119
rect 1126 114 1132 115
rect 1214 119 1220 120
rect 1214 115 1215 119
rect 1219 115 1220 119
rect 1214 114 1220 115
rect 1302 119 1308 120
rect 1302 115 1303 119
rect 1307 115 1308 119
rect 1302 114 1308 115
rect 1390 119 1396 120
rect 1390 115 1391 119
rect 1395 115 1396 119
rect 1390 114 1396 115
rect 1478 119 1484 120
rect 1478 115 1479 119
rect 1483 115 1484 119
rect 1478 114 1484 115
rect 1566 119 1572 120
rect 1566 115 1567 119
rect 1571 115 1572 119
rect 1566 114 1572 115
rect 1654 119 1660 120
rect 1654 115 1655 119
rect 1659 115 1660 119
rect 1654 114 1660 115
rect 1742 119 1748 120
rect 1742 115 1743 119
rect 1747 115 1748 119
rect 1902 119 1903 123
rect 1907 119 1908 123
rect 1902 118 1908 119
rect 1990 123 1996 124
rect 1990 119 1991 123
rect 1995 119 1996 123
rect 1990 118 1996 119
rect 2078 123 2084 124
rect 2078 119 2079 123
rect 2083 119 2084 123
rect 2078 118 2084 119
rect 2166 123 2172 124
rect 2166 119 2167 123
rect 2171 119 2172 123
rect 2166 118 2172 119
rect 2254 123 2260 124
rect 2254 119 2255 123
rect 2259 119 2260 123
rect 2254 118 2260 119
rect 2366 123 2372 124
rect 2366 119 2367 123
rect 2371 119 2372 123
rect 2366 118 2372 119
rect 2374 123 2380 124
rect 2374 119 2375 123
rect 2379 122 2380 123
rect 2582 123 2588 124
rect 2379 120 2449 122
rect 2379 119 2380 120
rect 2374 118 2380 119
rect 2582 119 2583 123
rect 2587 119 2588 123
rect 2582 118 2588 119
rect 2686 123 2692 124
rect 2686 119 2687 123
rect 2691 119 2692 123
rect 2686 118 2692 119
rect 2790 123 2796 124
rect 2790 119 2791 123
rect 2795 119 2796 123
rect 2790 118 2796 119
rect 2886 123 2892 124
rect 2886 119 2887 123
rect 2891 119 2892 123
rect 2886 118 2892 119
rect 2982 123 2988 124
rect 2982 119 2983 123
rect 2987 119 2988 123
rect 2982 118 2988 119
rect 3078 123 3084 124
rect 3078 119 3079 123
rect 3083 119 3084 123
rect 3078 118 3084 119
rect 3174 123 3180 124
rect 3174 119 3175 123
rect 3179 119 3180 123
rect 3174 118 3180 119
rect 3182 123 3188 124
rect 3182 119 3183 123
rect 3187 122 3188 123
rect 3358 123 3364 124
rect 3187 120 3233 122
rect 3187 119 3188 120
rect 3182 118 3188 119
rect 3358 119 3359 123
rect 3363 122 3364 123
rect 3363 120 3409 122
rect 3363 119 3364 120
rect 3358 118 3364 119
rect 1742 114 1748 115
rect 1806 115 1812 116
rect 110 111 116 112
rect 110 107 111 111
rect 115 107 116 111
rect 1766 111 1772 112
rect 110 106 116 107
rect 262 108 268 109
rect 262 104 263 108
rect 267 104 268 108
rect 262 103 268 104
rect 350 108 356 109
rect 350 104 351 108
rect 355 104 356 108
rect 350 103 356 104
rect 438 108 444 109
rect 438 104 439 108
rect 443 104 444 108
rect 438 103 444 104
rect 526 108 532 109
rect 526 104 527 108
rect 531 104 532 108
rect 526 103 532 104
rect 614 108 620 109
rect 614 104 615 108
rect 619 104 620 108
rect 614 103 620 104
rect 702 108 708 109
rect 702 104 703 108
rect 707 104 708 108
rect 702 103 708 104
rect 790 108 796 109
rect 790 104 791 108
rect 795 104 796 108
rect 790 103 796 104
rect 878 108 884 109
rect 878 104 879 108
rect 883 104 884 108
rect 878 103 884 104
rect 966 108 972 109
rect 966 104 967 108
rect 971 104 972 108
rect 966 103 972 104
rect 1054 108 1060 109
rect 1054 104 1055 108
rect 1059 104 1060 108
rect 1054 103 1060 104
rect 1142 108 1148 109
rect 1142 104 1143 108
rect 1147 104 1148 108
rect 1142 103 1148 104
rect 1230 108 1236 109
rect 1230 104 1231 108
rect 1235 104 1236 108
rect 1230 103 1236 104
rect 1318 108 1324 109
rect 1318 104 1319 108
rect 1323 104 1324 108
rect 1318 103 1324 104
rect 1406 108 1412 109
rect 1406 104 1407 108
rect 1411 104 1412 108
rect 1406 103 1412 104
rect 1494 108 1500 109
rect 1494 104 1495 108
rect 1499 104 1500 108
rect 1494 103 1500 104
rect 1582 108 1588 109
rect 1582 104 1583 108
rect 1587 104 1588 108
rect 1582 103 1588 104
rect 1670 108 1676 109
rect 1670 104 1671 108
rect 1675 104 1676 108
rect 1766 107 1767 111
rect 1771 107 1772 111
rect 1806 111 1807 115
rect 1811 111 1812 115
rect 3462 115 3468 116
rect 1806 110 1812 111
rect 1830 112 1836 113
rect 1830 108 1831 112
rect 1835 108 1836 112
rect 1830 107 1836 108
rect 1918 112 1924 113
rect 1918 108 1919 112
rect 1923 108 1924 112
rect 1918 107 1924 108
rect 2006 112 2012 113
rect 2006 108 2007 112
rect 2011 108 2012 112
rect 2006 107 2012 108
rect 2094 112 2100 113
rect 2094 108 2095 112
rect 2099 108 2100 112
rect 2094 107 2100 108
rect 2182 112 2188 113
rect 2182 108 2183 112
rect 2187 108 2188 112
rect 2182 107 2188 108
rect 2294 112 2300 113
rect 2294 108 2295 112
rect 2299 108 2300 112
rect 2294 107 2300 108
rect 2406 112 2412 113
rect 2406 108 2407 112
rect 2411 108 2412 112
rect 2406 107 2412 108
rect 2510 112 2516 113
rect 2510 108 2511 112
rect 2515 108 2516 112
rect 2510 107 2516 108
rect 2614 112 2620 113
rect 2614 108 2615 112
rect 2619 108 2620 112
rect 2614 107 2620 108
rect 2718 112 2724 113
rect 2718 108 2719 112
rect 2723 108 2724 112
rect 2718 107 2724 108
rect 2814 112 2820 113
rect 2814 108 2815 112
rect 2819 108 2820 112
rect 2814 107 2820 108
rect 2910 112 2916 113
rect 2910 108 2911 112
rect 2915 108 2916 112
rect 2910 107 2916 108
rect 3006 112 3012 113
rect 3006 108 3007 112
rect 3011 108 3012 112
rect 3006 107 3012 108
rect 3102 112 3108 113
rect 3102 108 3103 112
rect 3107 108 3108 112
rect 3102 107 3108 108
rect 3190 112 3196 113
rect 3190 108 3191 112
rect 3195 108 3196 112
rect 3190 107 3196 108
rect 3278 112 3284 113
rect 3278 108 3279 112
rect 3283 108 3284 112
rect 3278 107 3284 108
rect 3366 112 3372 113
rect 3366 108 3367 112
rect 3371 108 3372 112
rect 3462 111 3463 115
rect 3467 111 3468 115
rect 3462 110 3468 111
rect 3366 107 3372 108
rect 1766 106 1772 107
rect 1670 103 1676 104
<< m3c >>
rect 1343 3503 1347 3507
rect 207 3495 211 3499
rect 343 3495 347 3499
rect 511 3495 515 3499
rect 687 3495 691 3499
rect 1091 3491 1095 3495
rect 1191 3495 1195 3499
rect 1335 3495 1339 3499
rect 1479 3495 1483 3499
rect 1623 3495 1627 3499
rect 111 3480 115 3484
rect 135 3479 139 3483
rect 271 3479 275 3483
rect 439 3479 443 3483
rect 615 3479 619 3483
rect 791 3479 795 3483
rect 959 3479 963 3483
rect 1119 3479 1123 3483
rect 1263 3479 1267 3483
rect 1407 3479 1411 3483
rect 1551 3479 1555 3483
rect 1671 3479 1675 3483
rect 1767 3480 1771 3484
rect 207 3471 211 3475
rect 343 3471 347 3475
rect 511 3471 515 3475
rect 687 3471 691 3475
rect 783 3471 787 3475
rect 1091 3471 1095 3475
rect 1191 3471 1195 3475
rect 1335 3471 1339 3475
rect 1479 3471 1483 3475
rect 1623 3471 1627 3475
rect 1903 3483 1907 3487
rect 2047 3483 2051 3487
rect 2215 3483 2219 3487
rect 2575 3483 2579 3487
rect 2587 3483 2591 3487
rect 2711 3483 2715 3487
rect 2871 3483 2875 3487
rect 1807 3468 1811 3472
rect 111 3463 115 3467
rect 1831 3467 1835 3471
rect 135 3460 139 3464
rect 271 3460 275 3464
rect 439 3460 443 3464
rect 615 3460 619 3464
rect 791 3460 795 3464
rect 959 3460 963 3464
rect 1119 3460 1123 3464
rect 1263 3460 1267 3464
rect 1407 3460 1411 3464
rect 1551 3460 1555 3464
rect 1671 3460 1675 3464
rect 1767 3463 1771 3467
rect 1975 3467 1979 3471
rect 2143 3467 2147 3471
rect 2311 3467 2315 3471
rect 2479 3467 2483 3471
rect 2639 3467 2643 3471
rect 2799 3467 2803 3471
rect 2967 3467 2971 3471
rect 3463 3468 3467 3472
rect 1903 3459 1907 3463
rect 2047 3459 2051 3463
rect 2215 3459 2219 3463
rect 2223 3459 2227 3463
rect 2587 3459 2591 3463
rect 2711 3459 2715 3463
rect 2871 3459 2875 3463
rect 2883 3459 2887 3463
rect 1807 3451 1811 3455
rect 1831 3448 1835 3452
rect 1975 3448 1979 3452
rect 2143 3448 2147 3452
rect 2311 3448 2315 3452
rect 2479 3448 2483 3452
rect 2639 3448 2643 3452
rect 2799 3448 2803 3452
rect 2967 3448 2971 3452
rect 3463 3451 3467 3455
rect 187 3419 191 3423
rect 111 3409 115 3413
rect 135 3412 139 3416
rect 255 3412 259 3416
rect 415 3412 419 3416
rect 207 3403 211 3407
rect 327 3403 331 3407
rect 487 3403 491 3407
rect 575 3412 579 3416
rect 735 3412 739 3416
rect 895 3412 899 3416
rect 1063 3412 1067 3416
rect 1231 3412 1235 3416
rect 1399 3412 1403 3416
rect 2083 3415 2087 3419
rect 2223 3415 2227 3419
rect 1767 3409 1771 3413
rect 655 3403 659 3407
rect 1023 3403 1027 3407
rect 1135 3403 1139 3407
rect 1303 3403 1307 3407
rect 1343 3403 1347 3407
rect 1807 3401 1811 3405
rect 2031 3404 2035 3408
rect 2151 3404 2155 3408
rect 2271 3404 2275 3408
rect 2391 3404 2395 3408
rect 2511 3404 2515 3408
rect 2623 3404 2627 3408
rect 2727 3404 2731 3408
rect 2831 3404 2835 3408
rect 2935 3404 2939 3408
rect 3039 3404 3043 3408
rect 3151 3404 3155 3408
rect 3463 3401 3467 3405
rect 111 3392 115 3396
rect 135 3393 139 3397
rect 255 3393 259 3397
rect 415 3393 419 3397
rect 575 3393 579 3397
rect 735 3393 739 3397
rect 895 3393 899 3397
rect 1063 3393 1067 3397
rect 1231 3393 1235 3397
rect 1399 3393 1403 3397
rect 1767 3392 1771 3396
rect 2103 3395 2107 3399
rect 2223 3395 2227 3399
rect 2343 3395 2347 3399
rect 2351 3395 2355 3399
rect 2575 3395 2579 3399
rect 2591 3395 2595 3399
rect 2703 3395 2707 3399
rect 2903 3395 2907 3399
rect 3007 3395 3011 3399
rect 3111 3395 3115 3399
rect 3215 3395 3219 3399
rect 1807 3384 1811 3388
rect 2031 3385 2035 3389
rect 2151 3385 2155 3389
rect 2271 3385 2275 3389
rect 2391 3385 2395 3389
rect 2511 3385 2515 3389
rect 2623 3385 2627 3389
rect 2727 3385 2731 3389
rect 2831 3385 2835 3389
rect 2935 3385 2939 3389
rect 3039 3385 3043 3389
rect 3151 3385 3155 3389
rect 3463 3384 3467 3388
rect 187 3375 188 3379
rect 188 3375 191 3379
rect 207 3375 211 3379
rect 327 3375 331 3379
rect 655 3375 659 3379
rect 783 3375 784 3379
rect 784 3375 787 3379
rect 1007 3375 1011 3379
rect 1023 3375 1027 3379
rect 1135 3375 1139 3379
rect 1303 3375 1307 3379
rect 615 3363 619 3367
rect 2083 3367 2084 3371
rect 2084 3367 2087 3371
rect 2103 3367 2107 3371
rect 2223 3367 2227 3371
rect 2343 3367 2347 3371
rect 2591 3367 2595 3371
rect 2703 3367 2707 3371
rect 2775 3367 2776 3371
rect 2776 3367 2779 3371
rect 2883 3367 2884 3371
rect 2884 3367 2887 3371
rect 2903 3367 2907 3371
rect 3007 3367 3011 3371
rect 3111 3367 3115 3371
rect 487 3355 491 3359
rect 607 3355 611 3359
rect 1071 3355 1075 3359
rect 1199 3355 1203 3359
rect 1375 3355 1379 3359
rect 1599 3355 1603 3359
rect 1735 3355 1739 3359
rect 2351 3359 2355 3363
rect 2231 3351 2235 3355
rect 2367 3351 2371 3355
rect 2503 3351 2507 3355
rect 2783 3351 2787 3355
rect 2919 3351 2923 3355
rect 3055 3351 3059 3355
rect 3215 3351 3219 3355
rect 111 3340 115 3344
rect 135 3339 139 3343
rect 327 3339 331 3343
rect 535 3339 539 3343
rect 743 3339 747 3343
rect 935 3339 939 3343
rect 1119 3339 1123 3343
rect 1295 3339 1299 3343
rect 1463 3339 1467 3343
rect 1639 3339 1643 3343
rect 1767 3340 1771 3344
rect 1807 3336 1811 3340
rect 607 3331 611 3335
rect 615 3331 619 3335
rect 1007 3331 1011 3335
rect 1071 3331 1075 3335
rect 1199 3331 1203 3335
rect 1375 3331 1379 3335
rect 2159 3335 2163 3339
rect 1599 3331 1603 3335
rect 2295 3335 2299 3339
rect 2431 3335 2435 3339
rect 2567 3335 2571 3339
rect 2703 3335 2707 3339
rect 2839 3335 2843 3339
rect 2975 3335 2979 3339
rect 3119 3335 3123 3339
rect 3463 3336 3467 3340
rect 111 3323 115 3327
rect 135 3320 139 3324
rect 199 3323 203 3327
rect 327 3320 331 3324
rect 535 3320 539 3324
rect 743 3320 747 3324
rect 935 3320 939 3324
rect 1119 3320 1123 3324
rect 1295 3320 1299 3324
rect 1463 3320 1467 3324
rect 1639 3320 1643 3324
rect 1767 3323 1771 3327
rect 2231 3327 2235 3331
rect 2367 3327 2371 3331
rect 2503 3327 2507 3331
rect 1807 3319 1811 3323
rect 2639 3323 2643 3327
rect 2775 3327 2779 3331
rect 2911 3323 2915 3327
rect 2919 3327 2923 3331
rect 3055 3327 3059 3331
rect 2159 3316 2163 3320
rect 2295 3316 2299 3320
rect 2431 3316 2435 3320
rect 2567 3316 2571 3320
rect 2703 3316 2707 3320
rect 2839 3316 2843 3320
rect 2975 3316 2979 3320
rect 3119 3316 3123 3320
rect 3463 3319 3467 3323
rect 235 3275 239 3279
rect 111 3265 115 3269
rect 135 3268 139 3272
rect 279 3268 283 3272
rect 463 3268 467 3272
rect 647 3268 651 3272
rect 207 3259 211 3263
rect 351 3259 355 3263
rect 535 3259 539 3263
rect 719 3259 723 3263
rect 831 3268 835 3272
rect 1007 3268 1011 3272
rect 1175 3268 1179 3272
rect 1343 3268 1347 3272
rect 1503 3268 1507 3272
rect 1671 3268 1675 3272
rect 1767 3265 1771 3269
rect 1807 3269 1811 3273
rect 2087 3272 2091 3276
rect 2239 3272 2243 3276
rect 2399 3272 2403 3276
rect 2559 3272 2563 3276
rect 2719 3272 2723 3276
rect 2879 3272 2883 3276
rect 3039 3272 3043 3276
rect 3199 3272 3203 3276
rect 3463 3269 3467 3273
rect 1115 3259 1119 3263
rect 1247 3259 1251 3263
rect 1415 3259 1419 3263
rect 1575 3259 1579 3263
rect 1735 3259 1739 3263
rect 2159 3263 2163 3267
rect 2311 3263 2315 3267
rect 2479 3263 2483 3267
rect 2783 3263 2787 3267
rect 2951 3263 2955 3267
rect 3111 3263 3115 3267
rect 3263 3263 3267 3267
rect 111 3248 115 3252
rect 135 3249 139 3253
rect 279 3249 283 3253
rect 463 3249 467 3253
rect 647 3249 651 3253
rect 831 3249 835 3253
rect 1007 3249 1011 3253
rect 1175 3249 1179 3253
rect 1343 3249 1347 3253
rect 1503 3249 1507 3253
rect 1671 3249 1675 3253
rect 1767 3248 1771 3252
rect 1807 3252 1811 3256
rect 2087 3253 2091 3257
rect 2239 3253 2243 3257
rect 2399 3253 2403 3257
rect 2559 3253 2563 3257
rect 2719 3253 2723 3257
rect 2879 3253 2883 3257
rect 3039 3253 3043 3257
rect 3199 3253 3203 3257
rect 3463 3252 3467 3256
rect 199 3231 203 3235
rect 207 3231 211 3235
rect 351 3231 355 3235
rect 535 3231 539 3235
rect 719 3231 723 3235
rect 1115 3231 1119 3235
rect 1247 3231 1251 3235
rect 1415 3231 1419 3235
rect 1575 3231 1579 3235
rect 2159 3235 2163 3239
rect 2479 3235 2483 3239
rect 2639 3235 2643 3239
rect 2759 3235 2763 3239
rect 2911 3235 2915 3239
rect 2951 3235 2955 3239
rect 3111 3235 3115 3239
rect 1279 3219 1283 3223
rect 1399 3223 1403 3227
rect 1963 3219 1964 3223
rect 1964 3219 1967 3223
rect 1983 3219 1987 3223
rect 2119 3219 2123 3223
rect 2311 3219 2315 3223
rect 2431 3219 2435 3223
rect 2807 3219 2811 3223
rect 2831 3219 2835 3223
rect 3263 3219 3267 3223
rect 3303 3219 3307 3223
rect 235 3211 236 3215
rect 236 3211 239 3215
rect 255 3211 259 3215
rect 399 3211 403 3215
rect 559 3211 563 3215
rect 719 3211 723 3215
rect 1095 3207 1099 3211
rect 1251 3211 1255 3215
rect 1375 3211 1379 3215
rect 1807 3204 1811 3208
rect 1911 3203 1915 3207
rect 2047 3203 2051 3207
rect 2199 3203 2203 3207
rect 2359 3203 2363 3207
rect 2527 3203 2531 3207
rect 2687 3203 2691 3207
rect 2847 3203 2851 3207
rect 3007 3203 3011 3207
rect 3167 3203 3171 3207
rect 3335 3203 3339 3207
rect 3463 3204 3467 3208
rect 111 3196 115 3200
rect 183 3195 187 3199
rect 327 3195 331 3199
rect 487 3195 491 3199
rect 647 3195 651 3199
rect 807 3195 811 3199
rect 967 3195 971 3199
rect 1135 3195 1139 3199
rect 1303 3195 1307 3199
rect 1471 3195 1475 3199
rect 1767 3196 1771 3200
rect 1983 3195 1987 3199
rect 2119 3195 2123 3199
rect 255 3187 259 3191
rect 399 3187 403 3191
rect 559 3187 563 3191
rect 719 3187 723 3191
rect 735 3187 739 3191
rect 1095 3187 1099 3191
rect 1251 3187 1255 3191
rect 1375 3187 1379 3191
rect 1399 3187 1403 3191
rect 1807 3187 1811 3191
rect 2271 3191 2275 3195
rect 2431 3195 2435 3199
rect 2479 3195 2483 3199
rect 2759 3195 2763 3199
rect 2807 3195 2811 3199
rect 2967 3195 2971 3199
rect 3407 3191 3411 3195
rect 1911 3184 1915 3188
rect 111 3179 115 3183
rect 2047 3184 2051 3188
rect 2199 3184 2203 3188
rect 2359 3184 2363 3188
rect 2527 3184 2531 3188
rect 2687 3184 2691 3188
rect 2847 3184 2851 3188
rect 3007 3184 3011 3188
rect 3167 3184 3171 3188
rect 3335 3184 3339 3188
rect 3463 3187 3467 3191
rect 183 3176 187 3180
rect 327 3176 331 3180
rect 487 3176 491 3180
rect 647 3176 651 3180
rect 807 3176 811 3180
rect 967 3176 971 3180
rect 1135 3176 1139 3180
rect 1303 3176 1307 3180
rect 1471 3176 1475 3180
rect 1767 3179 1771 3183
rect 1963 3175 1967 3179
rect 2479 3175 2483 3179
rect 419 3143 423 3147
rect 735 3143 739 3147
rect 1807 3137 1811 3141
rect 1831 3140 1835 3144
rect 2007 3140 2011 3144
rect 2207 3140 2211 3144
rect 2399 3140 2403 3144
rect 2583 3140 2587 3144
rect 2759 3140 2763 3144
rect 2919 3140 2923 3144
rect 3079 3140 3083 3144
rect 3231 3140 3235 3144
rect 3367 3140 3371 3144
rect 111 3129 115 3133
rect 367 3132 371 3136
rect 487 3132 491 3136
rect 607 3132 611 3136
rect 727 3132 731 3136
rect 847 3132 851 3136
rect 967 3132 971 3136
rect 1079 3132 1083 3136
rect 1199 3132 1203 3136
rect 3463 3137 3467 3141
rect 1319 3132 1323 3136
rect 1767 3129 1771 3133
rect 1895 3131 1899 3135
rect 1911 3131 1915 3135
rect 2279 3131 2283 3135
rect 2287 3131 2291 3135
rect 2743 3131 2747 3135
rect 2831 3131 2835 3135
rect 2991 3131 2995 3135
rect 3151 3131 3155 3135
rect 3303 3131 3307 3135
rect 3431 3131 3435 3135
rect 439 3123 443 3127
rect 559 3123 563 3127
rect 679 3123 683 3127
rect 687 3123 691 3127
rect 919 3123 923 3127
rect 1039 3123 1043 3127
rect 1151 3123 1155 3127
rect 1271 3123 1275 3127
rect 1279 3123 1283 3127
rect 1807 3120 1811 3124
rect 1831 3121 1835 3125
rect 2007 3121 2011 3125
rect 2207 3121 2211 3125
rect 2399 3121 2403 3125
rect 2583 3121 2587 3125
rect 2759 3121 2763 3125
rect 2919 3121 2923 3125
rect 3079 3121 3083 3125
rect 3231 3121 3235 3125
rect 3367 3121 3371 3125
rect 3463 3120 3467 3124
rect 111 3112 115 3116
rect 367 3113 371 3117
rect 487 3113 491 3117
rect 607 3113 611 3117
rect 727 3113 731 3117
rect 847 3113 851 3117
rect 967 3113 971 3117
rect 1079 3113 1083 3117
rect 1199 3113 1203 3117
rect 1319 3113 1323 3117
rect 1767 3112 1771 3116
rect 1911 3103 1915 3107
rect 419 3095 420 3099
rect 420 3095 423 3099
rect 439 3095 443 3099
rect 559 3095 563 3099
rect 679 3095 683 3099
rect 687 3087 691 3091
rect 919 3095 923 3099
rect 1039 3095 1043 3099
rect 1151 3095 1155 3099
rect 1271 3095 1275 3099
rect 2271 3103 2275 3107
rect 2279 3103 2283 3107
rect 2287 3095 2291 3099
rect 2743 3103 2747 3107
rect 2967 3103 2968 3107
rect 2968 3103 2971 3107
rect 2991 3103 2995 3107
rect 3151 3103 3155 3107
rect 3407 3103 3411 3107
rect 1135 3087 1139 3091
rect 511 3079 515 3083
rect 599 3079 603 3083
rect 687 3079 691 3083
rect 775 3079 779 3083
rect 927 3079 928 3083
rect 928 3079 931 3083
rect 951 3079 955 3083
rect 1039 3079 1043 3083
rect 1127 3079 1131 3083
rect 1895 3083 1899 3087
rect 1903 3083 1907 3087
rect 2031 3083 2035 3087
rect 2191 3083 2195 3087
rect 2551 3083 2555 3087
rect 2559 3083 2563 3087
rect 2767 3083 2771 3087
rect 2991 3083 2995 3087
rect 3431 3083 3435 3087
rect 111 3064 115 3068
rect 439 3063 443 3067
rect 527 3063 531 3067
rect 615 3063 619 3067
rect 703 3063 707 3067
rect 791 3063 795 3067
rect 879 3063 883 3067
rect 967 3063 971 3067
rect 1055 3063 1059 3067
rect 1143 3063 1147 3067
rect 1767 3064 1771 3068
rect 1807 3068 1811 3072
rect 1831 3067 1835 3071
rect 1959 3067 1963 3071
rect 2119 3067 2123 3071
rect 2295 3067 2299 3071
rect 2487 3067 2491 3071
rect 2695 3067 2699 3071
rect 2919 3067 2923 3071
rect 3151 3067 3155 3071
rect 3367 3067 3371 3071
rect 3463 3068 3467 3072
rect 511 3055 515 3059
rect 599 3055 603 3059
rect 687 3055 691 3059
rect 775 3055 779 3059
rect 111 3047 115 3051
rect 863 3051 867 3055
rect 951 3055 955 3059
rect 1039 3055 1043 3059
rect 1127 3055 1131 3059
rect 1135 3055 1139 3059
rect 1903 3059 1907 3063
rect 2031 3059 2035 3063
rect 2191 3059 2195 3063
rect 439 3044 443 3048
rect 527 3044 531 3048
rect 615 3044 619 3048
rect 703 3044 707 3048
rect 791 3044 795 3048
rect 879 3044 883 3048
rect 967 3044 971 3048
rect 1055 3044 1059 3048
rect 1143 3044 1147 3048
rect 1767 3047 1771 3051
rect 1807 3051 1811 3055
rect 1831 3048 1835 3052
rect 1959 3048 1963 3052
rect 2119 3048 2123 3052
rect 2183 3051 2187 3055
rect 2559 3059 2563 3063
rect 2767 3059 2771 3063
rect 2991 3059 2995 3063
rect 2295 3048 2299 3052
rect 2487 3048 2491 3052
rect 2695 3048 2699 3052
rect 2919 3048 2923 3052
rect 3151 3048 3155 3052
rect 3367 3048 3371 3052
rect 3431 3051 3435 3055
rect 3463 3051 3467 3055
rect 111 2989 115 2993
rect 503 2992 507 2996
rect 591 2992 595 2996
rect 679 2992 683 2996
rect 767 2992 771 2996
rect 855 2992 859 2996
rect 943 2992 947 2996
rect 1031 2992 1035 2996
rect 1119 2992 1123 2996
rect 1207 2992 1211 2996
rect 1295 2992 1299 2996
rect 2551 2995 2555 2999
rect 1767 2989 1771 2993
rect 575 2983 579 2987
rect 663 2983 667 2987
rect 751 2983 755 2987
rect 759 2983 763 2987
rect 847 2983 851 2987
rect 935 2983 939 2987
rect 1023 2983 1027 2987
rect 1191 2983 1195 2987
rect 1279 2983 1283 2987
rect 1287 2983 1291 2987
rect 1807 2985 1811 2989
rect 1831 2988 1835 2992
rect 1919 2988 1923 2992
rect 2031 2988 2035 2992
rect 2143 2988 2147 2992
rect 2247 2988 2251 2992
rect 2359 2988 2363 2992
rect 2479 2988 2483 2992
rect 2623 2988 2627 2992
rect 2791 2988 2795 2992
rect 2983 2988 2987 2992
rect 1895 2979 1899 2983
rect 1911 2979 1915 2983
rect 2215 2979 2219 2983
rect 2319 2979 2323 2983
rect 2431 2979 2435 2983
rect 2551 2979 2555 2983
rect 2695 2979 2699 2983
rect 2863 2979 2867 2983
rect 3055 2979 3059 2983
rect 3183 2988 3187 2992
rect 3367 2988 3371 2992
rect 3463 2985 3467 2989
rect 3439 2979 3443 2983
rect 111 2972 115 2976
rect 503 2973 507 2977
rect 591 2973 595 2977
rect 679 2973 683 2977
rect 767 2973 771 2977
rect 855 2973 859 2977
rect 943 2973 947 2977
rect 1031 2973 1035 2977
rect 1119 2973 1123 2977
rect 1207 2973 1211 2977
rect 1295 2973 1299 2977
rect 1767 2972 1771 2976
rect 1807 2968 1811 2972
rect 1831 2969 1835 2973
rect 1919 2969 1923 2973
rect 2031 2969 2035 2973
rect 2143 2969 2147 2973
rect 2247 2969 2251 2973
rect 2359 2969 2363 2973
rect 2479 2969 2483 2973
rect 2623 2969 2627 2973
rect 2791 2969 2795 2973
rect 2983 2969 2987 2973
rect 3183 2969 3187 2973
rect 3367 2969 3371 2973
rect 3463 2968 3467 2972
rect 575 2955 579 2959
rect 663 2955 667 2959
rect 847 2955 851 2959
rect 863 2955 867 2959
rect 1023 2955 1027 2959
rect 759 2947 763 2951
rect 1167 2955 1168 2959
rect 1168 2955 1171 2959
rect 1191 2955 1195 2959
rect 1279 2955 1283 2959
rect 1287 2947 1291 2951
rect 1911 2951 1915 2955
rect 2183 2951 2187 2955
rect 2195 2951 2196 2955
rect 2196 2951 2199 2955
rect 2215 2951 2219 2955
rect 2319 2951 2323 2955
rect 2431 2951 2435 2955
rect 2551 2951 2555 2955
rect 2695 2951 2699 2955
rect 2863 2951 2867 2955
rect 3055 2951 3059 2955
rect 3431 2951 3435 2955
rect 799 2939 803 2943
rect 399 2931 403 2935
rect 519 2931 523 2935
rect 751 2931 755 2935
rect 783 2931 787 2935
rect 1183 2939 1187 2943
rect 111 2916 115 2920
rect 327 2915 331 2919
rect 447 2915 451 2919
rect 575 2915 579 2919
rect 711 2915 715 2919
rect 847 2915 851 2919
rect 975 2915 979 2919
rect 399 2907 403 2911
rect 519 2907 523 2911
rect 783 2907 787 2911
rect 799 2907 803 2911
rect 1311 2931 1315 2935
rect 1559 2931 1563 2935
rect 1895 2927 1899 2931
rect 1903 2927 1907 2931
rect 2295 2927 2299 2931
rect 2487 2927 2491 2931
rect 2639 2927 2640 2931
rect 2640 2927 2643 2931
rect 2895 2927 2899 2931
rect 2991 2927 2995 2931
rect 3143 2927 3147 2931
rect 3287 2927 3291 2931
rect 3295 2927 3299 2931
rect 1103 2915 1107 2919
rect 1167 2911 1171 2915
rect 1231 2915 1235 2919
rect 1359 2915 1363 2919
rect 1495 2915 1499 2919
rect 1767 2916 1771 2920
rect 1807 2912 1811 2916
rect 1183 2907 1187 2911
rect 1311 2907 1315 2911
rect 1831 2911 1835 2915
rect 2015 2911 2019 2915
rect 2215 2911 2219 2915
rect 2407 2911 2411 2915
rect 2591 2911 2595 2915
rect 2759 2911 2763 2915
rect 2911 2911 2915 2915
rect 3063 2911 3067 2915
rect 3207 2911 3211 2915
rect 3359 2911 3363 2915
rect 3463 2912 3467 2916
rect 111 2899 115 2903
rect 327 2896 331 2900
rect 447 2896 451 2900
rect 575 2896 579 2900
rect 639 2899 643 2903
rect 711 2896 715 2900
rect 847 2896 851 2900
rect 975 2896 979 2900
rect 1103 2896 1107 2900
rect 1231 2896 1235 2900
rect 1359 2896 1363 2900
rect 1495 2896 1499 2900
rect 1767 2899 1771 2903
rect 1903 2903 1907 2907
rect 1807 2895 1811 2899
rect 2087 2899 2091 2903
rect 2195 2903 2199 2907
rect 2295 2903 2299 2907
rect 2487 2903 2491 2907
rect 2831 2899 2835 2903
rect 2895 2903 2899 2907
rect 2991 2903 2995 2907
rect 3143 2903 3147 2907
rect 3287 2903 3291 2907
rect 1831 2892 1835 2896
rect 2015 2892 2019 2896
rect 2215 2892 2219 2896
rect 2407 2892 2411 2896
rect 2591 2892 2595 2896
rect 2759 2892 2763 2896
rect 2911 2892 2915 2896
rect 3063 2892 3067 2896
rect 3207 2892 3211 2896
rect 3359 2892 3363 2896
rect 3463 2895 3467 2899
rect 111 2841 115 2845
rect 135 2844 139 2848
rect 255 2844 259 2848
rect 415 2844 419 2848
rect 575 2844 579 2848
rect 735 2844 739 2848
rect 895 2844 899 2848
rect 1047 2844 1051 2848
rect 1191 2844 1195 2848
rect 1343 2844 1347 2848
rect 1495 2844 1499 2848
rect 1767 2841 1771 2845
rect 1807 2845 1811 2849
rect 1831 2848 1835 2852
rect 1999 2848 2003 2852
rect 2191 2848 2195 2852
rect 2383 2848 2387 2852
rect 2567 2848 2571 2852
rect 2735 2848 2739 2852
rect 2903 2848 2907 2852
rect 3063 2848 3067 2852
rect 3223 2848 3227 2852
rect 3367 2848 3371 2852
rect 3463 2845 3467 2849
rect 199 2835 203 2839
rect 215 2835 219 2839
rect 335 2835 339 2839
rect 647 2835 651 2839
rect 727 2835 731 2839
rect 967 2835 971 2839
rect 1119 2835 1123 2839
rect 1263 2835 1267 2839
rect 1415 2835 1419 2839
rect 1559 2835 1563 2839
rect 1895 2839 1899 2843
rect 1911 2839 1915 2843
rect 2263 2839 2267 2843
rect 2455 2839 2459 2843
rect 2639 2839 2643 2843
rect 2863 2839 2867 2843
rect 2975 2839 2979 2843
rect 3127 2839 3131 2843
rect 3295 2839 3299 2843
rect 3431 2839 3435 2843
rect 111 2824 115 2828
rect 135 2825 139 2829
rect 255 2825 259 2829
rect 415 2825 419 2829
rect 575 2825 579 2829
rect 735 2825 739 2829
rect 895 2825 899 2829
rect 1047 2825 1051 2829
rect 1191 2825 1195 2829
rect 1343 2825 1347 2829
rect 1495 2825 1499 2829
rect 1767 2824 1771 2828
rect 1807 2828 1811 2832
rect 1831 2829 1835 2833
rect 1999 2829 2003 2833
rect 2191 2829 2195 2833
rect 2383 2829 2387 2833
rect 2567 2829 2571 2833
rect 2735 2829 2739 2833
rect 2903 2829 2907 2833
rect 3063 2829 3067 2833
rect 3223 2829 3227 2833
rect 3367 2829 3371 2833
rect 3463 2828 3467 2832
rect 215 2807 219 2811
rect 335 2807 339 2811
rect 639 2807 643 2811
rect 647 2807 651 2811
rect 727 2799 731 2803
rect 967 2807 971 2811
rect 1119 2807 1123 2811
rect 1263 2807 1267 2811
rect 1415 2807 1419 2811
rect 1911 2811 1915 2815
rect 2087 2811 2091 2815
rect 2147 2811 2151 2815
rect 2263 2811 2267 2815
rect 2455 2811 2459 2815
rect 2831 2811 2835 2815
rect 2863 2811 2867 2815
rect 2975 2811 2979 2815
rect 3303 2811 3307 2815
rect 3439 2811 3443 2815
rect 1279 2799 1283 2803
rect 1895 2795 1899 2799
rect 2095 2795 2099 2799
rect 2295 2795 2299 2799
rect 2471 2795 2475 2799
rect 2991 2803 2995 2807
rect 2743 2795 2747 2799
rect 2823 2795 2827 2799
rect 3120 2795 3124 2799
rect 3263 2795 3267 2799
rect 3431 2795 3435 2799
rect 199 2783 203 2787
rect 207 2783 211 2787
rect 319 2783 323 2787
rect 463 2783 467 2787
rect 615 2783 619 2787
rect 903 2783 904 2787
rect 904 2783 907 2787
rect 927 2783 931 2787
rect 1095 2783 1099 2787
rect 1263 2783 1267 2787
rect 1607 2783 1611 2787
rect 1807 2780 1811 2784
rect 1831 2779 1835 2783
rect 2015 2779 2019 2783
rect 2147 2779 2151 2783
rect 2215 2779 2219 2783
rect 2407 2779 2411 2783
rect 2583 2779 2587 2783
rect 2751 2779 2755 2783
rect 2911 2779 2915 2783
rect 3071 2779 3075 2783
rect 3231 2779 3235 2783
rect 3367 2779 3371 2783
rect 3463 2780 3467 2784
rect 111 2768 115 2772
rect 135 2767 139 2771
rect 247 2767 251 2771
rect 391 2767 395 2771
rect 543 2767 547 2771
rect 695 2767 699 2771
rect 855 2767 859 2771
rect 1023 2767 1027 2771
rect 1191 2767 1195 2771
rect 1359 2767 1363 2771
rect 1527 2767 1531 2771
rect 1671 2767 1675 2771
rect 1767 2768 1771 2772
rect 2095 2771 2099 2775
rect 2295 2771 2299 2775
rect 2743 2771 2747 2775
rect 2823 2771 2827 2775
rect 207 2759 211 2763
rect 319 2759 323 2763
rect 463 2759 467 2763
rect 615 2759 619 2763
rect 623 2759 627 2763
rect 927 2759 931 2763
rect 1095 2759 1099 2763
rect 1263 2759 1267 2763
rect 1279 2759 1283 2763
rect 111 2751 115 2755
rect 1599 2755 1603 2759
rect 1607 2759 1611 2763
rect 1807 2763 1811 2767
rect 2983 2767 2987 2771
rect 2991 2771 2995 2775
rect 3303 2771 3307 2775
rect 3439 2767 3443 2771
rect 1831 2760 1835 2764
rect 2015 2760 2019 2764
rect 2215 2760 2219 2764
rect 2407 2760 2411 2764
rect 2583 2760 2587 2764
rect 2751 2760 2755 2764
rect 2911 2760 2915 2764
rect 3071 2760 3075 2764
rect 3231 2760 3235 2764
rect 3367 2760 3371 2764
rect 3463 2763 3467 2767
rect 135 2748 139 2752
rect 247 2748 251 2752
rect 391 2748 395 2752
rect 543 2748 547 2752
rect 695 2748 699 2752
rect 855 2748 859 2752
rect 1023 2748 1027 2752
rect 1191 2748 1195 2752
rect 1359 2748 1363 2752
rect 1527 2748 1531 2752
rect 1671 2748 1675 2752
rect 1767 2751 1771 2755
rect 299 2711 303 2715
rect 623 2711 627 2715
rect 111 2693 115 2697
rect 247 2696 251 2700
rect 359 2696 363 2700
rect 479 2696 483 2700
rect 615 2696 619 2700
rect 759 2696 763 2700
rect 911 2696 915 2700
rect 1063 2696 1067 2700
rect 1215 2696 1219 2700
rect 1375 2696 1379 2700
rect 1535 2696 1539 2700
rect 1671 2696 1675 2700
rect 1767 2693 1771 2697
rect 1807 2697 1811 2701
rect 2039 2700 2043 2704
rect 2159 2700 2163 2704
rect 2279 2700 2283 2704
rect 2407 2700 2411 2704
rect 2543 2700 2547 2704
rect 2687 2700 2691 2704
rect 2847 2700 2851 2704
rect 3023 2700 3027 2704
rect 3207 2700 3211 2704
rect 3367 2700 3371 2704
rect 3463 2697 3467 2701
rect 319 2687 323 2691
rect 431 2687 435 2691
rect 551 2687 555 2691
rect 687 2687 691 2691
rect 695 2687 699 2691
rect 903 2687 907 2691
rect 1135 2687 1139 2691
rect 1447 2687 1451 2691
rect 1607 2687 1611 2691
rect 1639 2687 1643 2691
rect 2111 2691 2115 2695
rect 2231 2691 2235 2695
rect 2351 2691 2355 2695
rect 2471 2691 2475 2695
rect 2615 2691 2619 2695
rect 2767 2691 2771 2695
rect 2775 2691 2779 2695
rect 3095 2691 3099 2695
rect 3103 2691 3107 2695
rect 3431 2691 3435 2695
rect 111 2676 115 2680
rect 247 2677 251 2681
rect 359 2677 363 2681
rect 479 2677 483 2681
rect 615 2677 619 2681
rect 759 2677 763 2681
rect 911 2677 915 2681
rect 1063 2677 1067 2681
rect 1215 2677 1219 2681
rect 1375 2677 1379 2681
rect 1535 2677 1539 2681
rect 1671 2677 1675 2681
rect 1767 2676 1771 2680
rect 1807 2680 1811 2684
rect 2039 2681 2043 2685
rect 2159 2681 2163 2685
rect 2279 2681 2283 2685
rect 2407 2681 2411 2685
rect 2543 2681 2547 2685
rect 2687 2681 2691 2685
rect 2847 2681 2851 2685
rect 3023 2681 3027 2685
rect 3207 2681 3211 2685
rect 3367 2681 3371 2685
rect 3463 2680 3467 2684
rect 299 2659 300 2663
rect 300 2659 303 2663
rect 319 2659 323 2663
rect 431 2659 435 2663
rect 551 2659 555 2663
rect 687 2659 691 2663
rect 1055 2659 1059 2663
rect 1135 2659 1139 2663
rect 695 2647 699 2651
rect 1599 2659 1603 2663
rect 1607 2659 1611 2663
rect 2111 2663 2115 2667
rect 2231 2663 2235 2667
rect 2351 2663 2355 2667
rect 1639 2651 1643 2655
rect 2263 2655 2267 2659
rect 2615 2663 2619 2667
rect 2775 2655 2779 2659
rect 2983 2663 2987 2667
rect 3095 2663 3099 2667
rect 3439 2663 3443 2667
rect 3103 2655 3107 2659
rect 535 2639 539 2643
rect 623 2639 627 2643
rect 711 2639 715 2643
rect 815 2639 819 2643
rect 1107 2639 1111 2643
rect 1207 2639 1211 2643
rect 1295 2639 1299 2643
rect 1447 2639 1451 2643
rect 1511 2639 1515 2643
rect 1903 2639 1907 2643
rect 1943 2639 1947 2643
rect 2063 2639 2067 2643
rect 2143 2639 2147 2643
rect 2255 2639 2259 2643
rect 2511 2639 2515 2643
rect 3139 2647 3143 2651
rect 2767 2639 2771 2643
rect 2831 2639 2835 2643
rect 3031 2639 3035 2643
rect 3431 2639 3435 2643
rect 111 2624 115 2628
rect 463 2623 467 2627
rect 551 2623 555 2627
rect 639 2623 643 2627
rect 743 2623 747 2627
rect 855 2623 859 2627
rect 983 2623 987 2627
rect 1127 2623 1131 2627
rect 1279 2623 1283 2627
rect 1439 2623 1443 2627
rect 1607 2623 1611 2627
rect 1767 2624 1771 2628
rect 1807 2624 1811 2628
rect 1871 2623 1875 2627
rect 1967 2623 1971 2627
rect 2071 2623 2075 2627
rect 2183 2623 2187 2627
rect 2295 2623 2299 2627
rect 2431 2623 2435 2627
rect 2583 2623 2587 2627
rect 2759 2623 2763 2627
rect 2959 2623 2963 2627
rect 3167 2623 3171 2627
rect 3367 2623 3371 2627
rect 3463 2624 3467 2628
rect 535 2615 539 2619
rect 623 2615 627 2619
rect 711 2615 715 2619
rect 815 2615 819 2619
rect 823 2615 827 2619
rect 1055 2615 1059 2619
rect 1107 2615 1111 2619
rect 1207 2615 1211 2619
rect 1511 2615 1515 2619
rect 111 2607 115 2611
rect 1679 2611 1683 2615
rect 1943 2615 1947 2619
rect 2063 2615 2067 2619
rect 2143 2615 2147 2619
rect 2255 2615 2259 2619
rect 2263 2615 2267 2619
rect 2395 2615 2399 2619
rect 2511 2615 2515 2619
rect 2831 2615 2835 2619
rect 3031 2615 3035 2619
rect 3139 2615 3143 2619
rect 463 2604 467 2608
rect 551 2604 555 2608
rect 639 2604 643 2608
rect 743 2604 747 2608
rect 855 2604 859 2608
rect 983 2604 987 2608
rect 1127 2604 1131 2608
rect 1279 2604 1283 2608
rect 1439 2604 1443 2608
rect 1607 2604 1611 2608
rect 1767 2607 1771 2611
rect 1807 2607 1811 2611
rect 3439 2611 3443 2615
rect 1871 2604 1875 2608
rect 1967 2604 1971 2608
rect 2071 2604 2075 2608
rect 2183 2604 2187 2608
rect 2295 2604 2299 2608
rect 2431 2604 2435 2608
rect 2583 2604 2587 2608
rect 2759 2604 2763 2608
rect 2959 2604 2963 2608
rect 3167 2604 3171 2608
rect 3367 2604 3371 2608
rect 3463 2607 3467 2611
rect 111 2549 115 2553
rect 503 2552 507 2556
rect 591 2552 595 2556
rect 679 2552 683 2556
rect 775 2552 779 2556
rect 879 2552 883 2556
rect 991 2552 995 2556
rect 1103 2552 1107 2556
rect 1223 2552 1227 2556
rect 1351 2552 1355 2556
rect 1479 2552 1483 2556
rect 1607 2552 1611 2556
rect 2579 2555 2583 2559
rect 1767 2549 1771 2553
rect 575 2543 579 2547
rect 663 2543 667 2547
rect 751 2543 755 2547
rect 847 2543 851 2547
rect 951 2543 955 2547
rect 1063 2543 1067 2547
rect 1175 2543 1179 2547
rect 1295 2543 1299 2547
rect 1423 2543 1427 2547
rect 1431 2543 1435 2547
rect 1559 2543 1563 2547
rect 1807 2545 1811 2549
rect 1831 2548 1835 2552
rect 1919 2548 1923 2552
rect 2007 2548 2011 2552
rect 2111 2548 2115 2552
rect 2223 2548 2227 2552
rect 2343 2548 2347 2552
rect 2487 2548 2491 2552
rect 2647 2548 2651 2552
rect 2815 2548 2819 2552
rect 1903 2539 1907 2543
rect 1911 2539 1915 2543
rect 2087 2539 2091 2543
rect 2191 2539 2195 2543
rect 2415 2539 2419 2543
rect 2559 2539 2563 2543
rect 2719 2539 2723 2543
rect 2887 2539 2891 2543
rect 2999 2548 3003 2552
rect 3191 2548 3195 2552
rect 3367 2548 3371 2552
rect 3463 2545 3467 2549
rect 3263 2539 3267 2543
rect 3431 2539 3435 2543
rect 111 2532 115 2536
rect 503 2533 507 2537
rect 591 2533 595 2537
rect 679 2533 683 2537
rect 775 2533 779 2537
rect 879 2533 883 2537
rect 991 2533 995 2537
rect 1103 2533 1107 2537
rect 1223 2533 1227 2537
rect 1351 2533 1355 2537
rect 1479 2533 1483 2537
rect 1607 2533 1611 2537
rect 1767 2532 1771 2536
rect 1807 2528 1811 2532
rect 1831 2529 1835 2533
rect 1919 2529 1923 2533
rect 2007 2529 2011 2533
rect 2111 2529 2115 2533
rect 2223 2529 2227 2533
rect 2343 2529 2347 2533
rect 2487 2529 2491 2533
rect 2647 2529 2651 2533
rect 2815 2529 2819 2533
rect 2999 2529 3003 2533
rect 3191 2529 3195 2533
rect 3367 2529 3371 2533
rect 3463 2528 3467 2532
rect 575 2515 579 2519
rect 663 2515 667 2519
rect 751 2515 755 2519
rect 847 2515 851 2519
rect 951 2515 955 2519
rect 1063 2515 1067 2519
rect 1175 2515 1179 2519
rect 1431 2515 1435 2519
rect 1559 2515 1563 2519
rect 1679 2515 1683 2519
rect 823 2507 827 2511
rect 1911 2511 1915 2515
rect 2087 2511 2091 2515
rect 2191 2511 2195 2515
rect 2207 2511 2211 2515
rect 2395 2511 2396 2515
rect 2396 2511 2399 2515
rect 2415 2511 2419 2515
rect 2559 2511 2563 2515
rect 2719 2511 2723 2515
rect 2887 2511 2891 2515
rect 3243 2511 3244 2515
rect 3244 2511 3247 2515
rect 3439 2511 3443 2515
rect 631 2495 635 2499
rect 815 2495 819 2499
rect 991 2491 995 2495
rect 1519 2503 1523 2507
rect 1423 2495 1427 2499
rect 1471 2495 1475 2499
rect 2015 2499 2019 2503
rect 2023 2499 2027 2503
rect 2319 2499 2323 2503
rect 2375 2499 2379 2503
rect 2579 2499 2580 2503
rect 2580 2499 2583 2503
rect 2599 2499 2603 2503
rect 2783 2499 2787 2503
rect 2991 2499 2995 2503
rect 3431 2499 3435 2503
rect 111 2480 115 2484
rect 551 2479 555 2483
rect 735 2479 739 2483
rect 911 2479 915 2483
rect 1079 2479 1083 2483
rect 1239 2479 1243 2483
rect 1399 2479 1403 2483
rect 1567 2479 1571 2483
rect 1767 2480 1771 2484
rect 1807 2484 1811 2488
rect 1951 2483 1955 2487
rect 2039 2483 2043 2487
rect 2135 2483 2139 2487
rect 2239 2483 2243 2487
rect 2367 2483 2371 2487
rect 2527 2483 2531 2487
rect 2711 2483 2715 2487
rect 2919 2483 2923 2487
rect 3143 2483 3147 2487
rect 3367 2483 3371 2487
rect 3463 2484 3467 2488
rect 111 2463 115 2467
rect 623 2467 627 2471
rect 631 2471 635 2475
rect 815 2471 819 2475
rect 1151 2467 1155 2471
rect 1471 2471 1475 2475
rect 1519 2471 1523 2475
rect 2023 2475 2027 2479
rect 2207 2475 2211 2479
rect 2215 2475 2219 2479
rect 2319 2475 2323 2479
rect 2599 2475 2603 2479
rect 2783 2475 2787 2479
rect 2991 2475 2995 2479
rect 3079 2475 3083 2479
rect 3243 2475 3247 2479
rect 551 2460 555 2464
rect 735 2460 739 2464
rect 911 2460 915 2464
rect 1079 2460 1083 2464
rect 1239 2460 1243 2464
rect 1399 2460 1403 2464
rect 1567 2460 1571 2464
rect 1767 2463 1771 2467
rect 1807 2467 1811 2471
rect 1951 2464 1955 2468
rect 2039 2464 2043 2468
rect 2135 2464 2139 2468
rect 2239 2464 2243 2468
rect 2367 2464 2371 2468
rect 2527 2464 2531 2468
rect 2711 2464 2715 2468
rect 2919 2464 2923 2468
rect 3143 2464 3147 2468
rect 3367 2464 3371 2468
rect 3463 2467 3467 2471
rect 2619 2427 2623 2431
rect 3079 2427 3083 2431
rect 111 2413 115 2417
rect 415 2416 419 2420
rect 503 2416 507 2420
rect 599 2416 603 2420
rect 703 2416 707 2420
rect 807 2416 811 2420
rect 919 2416 923 2420
rect 1039 2416 1043 2420
rect 1167 2416 1171 2420
rect 1295 2416 1299 2420
rect 1423 2416 1427 2420
rect 2263 2419 2267 2423
rect 1767 2413 1771 2417
rect 487 2407 491 2411
rect 575 2407 579 2411
rect 583 2407 587 2411
rect 775 2407 779 2411
rect 879 2407 883 2411
rect 991 2407 995 2411
rect 999 2407 1003 2411
rect 1239 2407 1243 2411
rect 1367 2407 1371 2411
rect 1387 2407 1391 2411
rect 1807 2409 1811 2413
rect 2215 2412 2219 2416
rect 2303 2412 2307 2416
rect 2287 2403 2291 2407
rect 2375 2403 2379 2407
rect 2751 2419 2755 2423
rect 2391 2412 2395 2416
rect 2479 2412 2483 2416
rect 2567 2412 2571 2416
rect 2655 2412 2659 2416
rect 2743 2412 2747 2416
rect 2839 2412 2843 2416
rect 2639 2403 2643 2407
rect 2727 2403 2731 2407
rect 2815 2403 2819 2407
rect 2935 2412 2939 2416
rect 3463 2409 3467 2413
rect 111 2396 115 2400
rect 415 2397 419 2401
rect 503 2397 507 2401
rect 599 2397 603 2401
rect 703 2397 707 2401
rect 807 2397 811 2401
rect 919 2397 923 2401
rect 1039 2397 1043 2401
rect 1167 2397 1171 2401
rect 1295 2397 1299 2401
rect 1423 2397 1427 2401
rect 1767 2396 1771 2400
rect 1807 2392 1811 2396
rect 2215 2393 2219 2397
rect 2303 2393 2307 2397
rect 2391 2393 2395 2397
rect 2479 2393 2483 2397
rect 2567 2393 2571 2397
rect 2655 2393 2659 2397
rect 2743 2393 2747 2397
rect 2839 2393 2843 2397
rect 2927 2395 2931 2399
rect 2935 2393 2939 2397
rect 3463 2392 3467 2396
rect 487 2379 491 2383
rect 623 2379 627 2383
rect 583 2371 587 2375
rect 775 2379 779 2383
rect 879 2379 883 2383
rect 1063 2379 1067 2383
rect 1151 2379 1155 2383
rect 1239 2379 1243 2383
rect 1367 2379 1371 2383
rect 2263 2381 2267 2383
rect 2263 2379 2264 2381
rect 2264 2379 2267 2381
rect 999 2371 1003 2375
rect 2287 2375 2291 2379
rect 2551 2375 2555 2379
rect 2619 2375 2620 2379
rect 2620 2375 2623 2379
rect 2639 2375 2643 2379
rect 2727 2375 2731 2379
rect 2815 2375 2819 2379
rect 2927 2375 2931 2379
rect 399 2363 403 2367
rect 551 2363 555 2367
rect 575 2363 579 2367
rect 615 2363 619 2367
rect 847 2363 851 2367
rect 867 2363 871 2367
rect 951 2363 955 2367
rect 1207 2363 1211 2367
rect 1387 2363 1388 2367
rect 1388 2363 1391 2367
rect 2231 2363 2235 2367
rect 2239 2363 2243 2367
rect 2335 2363 2339 2367
rect 2439 2363 2443 2367
rect 2543 2363 2547 2367
rect 2751 2363 2755 2367
rect 2759 2363 2763 2367
rect 2871 2363 2875 2367
rect 2983 2363 2987 2367
rect 111 2348 115 2352
rect 319 2347 323 2351
rect 431 2347 435 2351
rect 543 2347 547 2351
rect 655 2347 659 2351
rect 767 2347 771 2351
rect 879 2347 883 2351
rect 991 2347 995 2351
rect 1103 2347 1107 2351
rect 1215 2347 1219 2351
rect 1335 2347 1339 2351
rect 1767 2348 1771 2352
rect 1807 2348 1811 2352
rect 2167 2347 2171 2351
rect 2263 2347 2267 2351
rect 2367 2347 2371 2351
rect 2471 2347 2475 2351
rect 2575 2347 2579 2351
rect 2687 2347 2691 2351
rect 2799 2347 2803 2351
rect 2911 2347 2915 2351
rect 3023 2347 3027 2351
rect 3463 2348 3467 2352
rect 399 2339 403 2343
rect 615 2339 619 2343
rect 111 2331 115 2335
rect 319 2328 323 2332
rect 399 2331 403 2335
rect 431 2328 435 2332
rect 543 2328 547 2332
rect 551 2323 555 2327
rect 867 2339 871 2343
rect 951 2339 955 2343
rect 1063 2339 1067 2343
rect 1071 2339 1075 2343
rect 1207 2339 1211 2343
rect 2239 2339 2243 2343
rect 2335 2339 2339 2343
rect 2439 2339 2443 2343
rect 2543 2339 2547 2343
rect 2551 2339 2555 2343
rect 2759 2339 2763 2343
rect 2871 2339 2875 2343
rect 2983 2339 2987 2343
rect 2991 2339 2995 2343
rect 655 2328 659 2332
rect 767 2328 771 2332
rect 879 2328 883 2332
rect 991 2328 995 2332
rect 1103 2328 1107 2332
rect 1215 2328 1219 2332
rect 1335 2328 1339 2332
rect 1767 2331 1771 2335
rect 1807 2331 1811 2335
rect 2167 2328 2171 2332
rect 2263 2328 2267 2332
rect 2367 2328 2371 2332
rect 2471 2328 2475 2332
rect 2575 2328 2579 2332
rect 2687 2328 2691 2332
rect 2799 2328 2803 2332
rect 2911 2328 2915 2332
rect 3023 2328 3027 2332
rect 3463 2331 3467 2335
rect 203 2283 207 2287
rect 111 2273 115 2277
rect 151 2276 155 2280
rect 271 2276 275 2280
rect 391 2276 395 2280
rect 519 2276 523 2280
rect 223 2267 227 2271
rect 343 2267 347 2271
rect 463 2267 467 2271
rect 591 2267 595 2271
rect 2231 2283 2235 2287
rect 647 2276 651 2280
rect 775 2276 779 2280
rect 895 2276 899 2280
rect 1015 2276 1019 2280
rect 1143 2276 1147 2280
rect 1271 2276 1275 2280
rect 1767 2273 1771 2277
rect 1807 2273 1811 2277
rect 1887 2276 1891 2280
rect 2039 2276 2043 2280
rect 2199 2276 2203 2280
rect 2375 2276 2379 2280
rect 847 2267 851 2271
rect 855 2267 859 2271
rect 1087 2267 1091 2271
rect 1215 2267 1219 2271
rect 1223 2267 1227 2271
rect 1959 2267 1963 2271
rect 2111 2267 2115 2271
rect 2271 2267 2275 2271
rect 2447 2267 2451 2271
rect 2551 2276 2555 2280
rect 2719 2276 2723 2280
rect 2887 2276 2891 2280
rect 3055 2276 3059 2280
rect 3223 2276 3227 2280
rect 3367 2276 3371 2280
rect 3463 2273 3467 2277
rect 2707 2267 2711 2271
rect 2799 2267 2803 2271
rect 3127 2267 3131 2271
rect 3295 2267 3299 2271
rect 3431 2267 3435 2271
rect 111 2256 115 2260
rect 151 2257 155 2261
rect 271 2257 275 2261
rect 391 2257 395 2261
rect 519 2257 523 2261
rect 647 2257 651 2261
rect 775 2257 779 2261
rect 895 2257 899 2261
rect 1015 2257 1019 2261
rect 1143 2257 1147 2261
rect 1271 2257 1275 2261
rect 1767 2256 1771 2260
rect 1807 2256 1811 2260
rect 1887 2257 1891 2261
rect 2039 2257 2043 2261
rect 2199 2257 2203 2261
rect 2375 2257 2379 2261
rect 2551 2257 2555 2261
rect 2719 2257 2723 2261
rect 2887 2257 2891 2261
rect 3055 2257 3059 2261
rect 3223 2257 3227 2261
rect 3367 2257 3371 2261
rect 3463 2256 3467 2260
rect 203 2239 204 2243
rect 204 2239 207 2243
rect 223 2239 227 2243
rect 399 2239 403 2243
rect 463 2239 467 2243
rect 591 2239 595 2243
rect 855 2239 859 2243
rect 943 2239 944 2243
rect 944 2239 947 2243
rect 1064 2239 1068 2243
rect 1087 2239 1091 2243
rect 1215 2239 1219 2243
rect 1951 2239 1955 2243
rect 1959 2239 1963 2243
rect 2111 2239 2115 2243
rect 2271 2239 2275 2243
rect 2447 2239 2451 2243
rect 2799 2239 2803 2243
rect 2991 2239 2995 2243
rect 3031 2239 3035 2243
rect 3127 2239 3131 2243
rect 3295 2239 3299 2243
rect 215 2223 219 2227
rect 739 2231 743 2235
rect 343 2223 347 2227
rect 479 2223 483 2227
rect 655 2223 659 2227
rect 1079 2223 1083 2227
rect 1223 2223 1227 2227
rect 1303 2223 1307 2227
rect 1391 2223 1395 2227
rect 1575 2223 1579 2227
rect 1743 2227 1747 2231
rect 1903 2227 1907 2231
rect 2207 2227 2211 2231
rect 2383 2227 2387 2231
rect 2707 2227 2708 2231
rect 2708 2227 2711 2231
rect 2727 2227 2731 2231
rect 3039 2227 3043 2231
rect 3183 2227 3187 2231
rect 3431 2227 3435 2231
rect 111 2208 115 2212
rect 135 2207 139 2211
rect 247 2207 251 2211
rect 407 2207 411 2211
rect 583 2207 587 2211
rect 767 2207 771 2211
rect 951 2207 955 2211
rect 1135 2207 1139 2211
rect 1319 2207 1323 2211
rect 1503 2207 1507 2211
rect 1671 2207 1675 2211
rect 1767 2208 1771 2212
rect 1807 2212 1811 2216
rect 1831 2211 1835 2215
rect 1967 2211 1971 2215
rect 2135 2211 2139 2215
rect 2311 2211 2315 2215
rect 2487 2211 2491 2215
rect 2655 2211 2659 2215
rect 2815 2211 2819 2215
rect 2959 2211 2963 2215
rect 3103 2211 3107 2215
rect 3247 2211 3251 2215
rect 3367 2211 3371 2215
rect 3463 2212 3467 2216
rect 215 2199 219 2203
rect 479 2199 483 2203
rect 655 2199 659 2203
rect 739 2199 743 2203
rect 943 2199 947 2203
rect 1079 2199 1083 2203
rect 1391 2199 1395 2203
rect 1575 2199 1579 2203
rect 1743 2199 1747 2203
rect 1903 2203 1907 2207
rect 2207 2203 2211 2207
rect 2383 2203 2387 2207
rect 2419 2203 2423 2207
rect 2727 2203 2731 2207
rect 111 2191 115 2195
rect 135 2188 139 2192
rect 199 2191 203 2195
rect 247 2188 251 2192
rect 407 2188 411 2192
rect 583 2188 587 2192
rect 767 2188 771 2192
rect 951 2188 955 2192
rect 1135 2188 1139 2192
rect 1319 2188 1323 2192
rect 1503 2188 1507 2192
rect 1671 2188 1675 2192
rect 1767 2191 1771 2195
rect 1807 2195 1811 2199
rect 2887 2199 2891 2203
rect 3031 2203 3035 2207
rect 3039 2203 3043 2207
rect 3183 2203 3187 2207
rect 3439 2199 3443 2203
rect 1831 2192 1835 2196
rect 1967 2192 1971 2196
rect 2135 2192 2139 2196
rect 2311 2192 2315 2196
rect 2487 2192 2491 2196
rect 2655 2192 2659 2196
rect 2815 2192 2819 2196
rect 2959 2192 2963 2196
rect 3103 2192 3107 2196
rect 3247 2192 3251 2196
rect 3367 2192 3371 2196
rect 3463 2195 3467 2199
rect 1951 2183 1955 2187
rect 2419 2183 2423 2187
rect 1807 2145 1811 2149
rect 2927 2148 2931 2152
rect 3015 2148 3019 2152
rect 3103 2148 3107 2152
rect 3191 2148 3195 2152
rect 3279 2148 3283 2152
rect 3367 2148 3371 2152
rect 3463 2145 3467 2149
rect 111 2133 115 2137
rect 135 2136 139 2140
rect 247 2136 251 2140
rect 391 2136 395 2140
rect 543 2136 547 2140
rect 695 2136 699 2140
rect 839 2136 843 2140
rect 975 2136 979 2140
rect 1103 2136 1107 2140
rect 1231 2136 1235 2140
rect 1351 2136 1355 2140
rect 1463 2136 1467 2140
rect 1575 2136 1579 2140
rect 1671 2136 1675 2140
rect 2999 2139 3003 2143
rect 3087 2139 3091 2143
rect 3255 2139 3259 2143
rect 3351 2139 3355 2143
rect 3359 2139 3363 2143
rect 1767 2133 1771 2137
rect 207 2127 211 2131
rect 319 2127 323 2131
rect 463 2127 467 2131
rect 615 2127 619 2131
rect 623 2127 627 2131
rect 951 2127 955 2131
rect 1055 2127 1059 2131
rect 1175 2127 1179 2131
rect 1303 2127 1307 2131
rect 1311 2127 1315 2131
rect 1431 2127 1435 2131
rect 1543 2127 1547 2131
rect 1655 2127 1659 2131
rect 1807 2128 1811 2132
rect 2927 2129 2931 2133
rect 3015 2129 3019 2133
rect 3103 2129 3107 2133
rect 3191 2129 3195 2133
rect 3279 2129 3283 2133
rect 3367 2129 3371 2133
rect 3463 2128 3467 2132
rect 111 2116 115 2120
rect 135 2117 139 2121
rect 247 2117 251 2121
rect 391 2117 395 2121
rect 543 2117 547 2121
rect 695 2117 699 2121
rect 839 2117 843 2121
rect 975 2117 979 2121
rect 1103 2117 1107 2121
rect 1231 2117 1235 2121
rect 1351 2117 1355 2121
rect 1463 2117 1467 2121
rect 1575 2117 1579 2121
rect 1671 2117 1675 2121
rect 1767 2116 1771 2120
rect 2887 2111 2891 2115
rect 2999 2111 3003 2115
rect 3087 2111 3091 2115
rect 3359 2111 3363 2115
rect 3439 2111 3443 2115
rect 199 2099 203 2103
rect 207 2099 211 2103
rect 319 2099 323 2103
rect 463 2099 467 2103
rect 615 2099 619 2103
rect 951 2099 955 2103
rect 623 2091 627 2095
rect 1175 2099 1179 2103
rect 1431 2099 1435 2103
rect 1543 2099 1547 2103
rect 1655 2099 1659 2103
rect 1787 2099 1791 2103
rect 1311 2091 1315 2095
rect 1939 2091 1943 2095
rect 2395 2091 2396 2095
rect 2396 2091 2399 2095
rect 2583 2091 2587 2095
rect 2735 2091 2739 2095
rect 3255 2099 3259 2103
rect 3087 2091 3088 2095
rect 3088 2091 3091 2095
rect 3111 2091 3115 2095
rect 3231 2091 3235 2095
rect 3351 2091 3355 2095
rect 295 2083 299 2087
rect 415 2083 419 2087
rect 535 2083 539 2087
rect 755 2083 756 2087
rect 756 2083 759 2087
rect 775 2083 779 2087
rect 895 2083 899 2087
rect 1055 2083 1059 2087
rect 1119 2083 1123 2087
rect 1259 2083 1263 2087
rect 1807 2076 1811 2080
rect 111 2068 115 2072
rect 135 2067 139 2071
rect 1831 2075 1835 2079
rect 1991 2075 1995 2079
rect 2167 2075 2171 2079
rect 2343 2075 2347 2079
rect 2503 2075 2507 2079
rect 2655 2075 2659 2079
rect 2791 2075 2795 2079
rect 2919 2075 2923 2079
rect 3039 2075 3043 2079
rect 3159 2075 3163 2079
rect 3271 2075 3275 2079
rect 3367 2075 3371 2079
rect 3463 2076 3467 2080
rect 223 2067 227 2071
rect 343 2067 347 2071
rect 463 2067 467 2071
rect 583 2067 587 2071
rect 703 2067 707 2071
rect 823 2067 827 2071
rect 935 2067 939 2071
rect 1047 2067 1051 2071
rect 1159 2067 1163 2071
rect 1279 2067 1283 2071
rect 1767 2068 1771 2072
rect 1787 2067 1791 2071
rect 1939 2067 1943 2071
rect 295 2059 299 2063
rect 415 2059 419 2063
rect 535 2059 539 2063
rect 543 2059 547 2063
rect 775 2059 779 2063
rect 895 2059 899 2063
rect 1119 2059 1123 2063
rect 1259 2059 1263 2063
rect 1271 2059 1275 2063
rect 1807 2059 1811 2063
rect 2575 2063 2579 2067
rect 2583 2067 2587 2071
rect 2735 2067 2739 2071
rect 3111 2067 3115 2071
rect 3231 2067 3235 2071
rect 3439 2063 3443 2067
rect 1831 2056 1835 2060
rect 111 2051 115 2055
rect 1991 2056 1995 2060
rect 2167 2056 2171 2060
rect 2343 2056 2347 2060
rect 2503 2056 2507 2060
rect 2655 2056 2659 2060
rect 2791 2056 2795 2060
rect 2919 2056 2923 2060
rect 3039 2056 3043 2060
rect 3159 2056 3163 2060
rect 3271 2056 3275 2060
rect 3367 2056 3371 2060
rect 3463 2059 3467 2063
rect 135 2048 139 2052
rect 223 2048 227 2052
rect 343 2048 347 2052
rect 463 2048 467 2052
rect 583 2048 587 2052
rect 703 2048 707 2052
rect 823 2048 827 2052
rect 935 2048 939 2052
rect 1047 2048 1051 2052
rect 1159 2048 1163 2052
rect 1279 2048 1283 2052
rect 1767 2051 1771 2055
rect 187 2011 191 2015
rect 543 2011 547 2015
rect 1807 2005 1811 2009
rect 1831 2008 1835 2012
rect 2015 2008 2019 2012
rect 2223 2008 2227 2012
rect 2431 2008 2435 2012
rect 2631 2008 2635 2012
rect 2823 2008 2827 2012
rect 3007 2008 3011 2012
rect 3199 2008 3203 2012
rect 3367 2008 3371 2012
rect 3463 2005 3467 2009
rect 111 1993 115 1997
rect 135 1996 139 2000
rect 239 1996 243 2000
rect 367 1996 371 2000
rect 503 1996 507 2000
rect 639 1996 643 2000
rect 775 1996 779 2000
rect 911 1996 915 2000
rect 1047 1996 1051 2000
rect 1183 1996 1187 2000
rect 1327 1996 1331 2000
rect 1967 1999 1971 2003
rect 2087 1999 2091 2003
rect 2295 1999 2299 2003
rect 2395 1999 2399 2003
rect 2703 1999 2707 2003
rect 2895 1999 2899 2003
rect 2999 1999 3003 2003
rect 3087 1999 3091 2003
rect 3431 1999 3435 2003
rect 1767 1993 1771 1997
rect 207 1987 211 1991
rect 311 1987 315 1991
rect 439 1987 443 1991
rect 575 1987 579 1991
rect 583 1987 587 1991
rect 755 1987 759 1991
rect 855 1987 859 1991
rect 1135 1987 1139 1991
rect 1255 1987 1259 1991
rect 1399 1987 1403 1991
rect 1807 1988 1811 1992
rect 1831 1989 1835 1993
rect 2015 1989 2019 1993
rect 2223 1989 2227 1993
rect 2431 1989 2435 1993
rect 2631 1989 2635 1993
rect 2823 1989 2827 1993
rect 3007 1989 3011 1993
rect 3199 1989 3203 1993
rect 3367 1989 3371 1993
rect 3463 1988 3467 1992
rect 111 1976 115 1980
rect 135 1977 139 1981
rect 239 1977 243 1981
rect 367 1977 371 1981
rect 503 1977 507 1981
rect 639 1977 643 1981
rect 775 1977 779 1981
rect 911 1977 915 1981
rect 1047 1977 1051 1981
rect 1183 1977 1187 1981
rect 1327 1977 1331 1981
rect 1767 1976 1771 1980
rect 1935 1971 1939 1975
rect 1967 1971 1971 1975
rect 2087 1971 2091 1975
rect 2295 1971 2299 1975
rect 2575 1971 2579 1975
rect 2703 1971 2707 1975
rect 2895 1971 2899 1975
rect 3239 1971 3243 1975
rect 3439 1971 3443 1975
rect 187 1959 188 1963
rect 188 1959 191 1963
rect 207 1959 211 1963
rect 311 1959 315 1963
rect 439 1959 443 1963
rect 575 1959 579 1963
rect 855 1959 859 1963
rect 963 1959 964 1963
rect 964 1959 967 1963
rect 583 1951 587 1955
rect 1135 1959 1139 1963
rect 1255 1959 1259 1963
rect 1271 1951 1275 1955
rect 2079 1955 2083 1959
rect 2367 1963 2371 1967
rect 2299 1955 2303 1959
rect 2359 1955 2363 1959
rect 2655 1955 2659 1959
rect 2799 1955 2803 1959
rect 2911 1955 2915 1959
rect 2999 1955 3000 1959
rect 3000 1955 3003 1959
rect 3247 1963 3251 1967
rect 3135 1955 3139 1959
rect 3359 1955 3363 1959
rect 3431 1955 3435 1959
rect 403 1943 407 1947
rect 495 1943 499 1947
rect 631 1943 635 1947
rect 951 1943 955 1947
rect 111 1928 115 1932
rect 295 1927 299 1931
rect 423 1927 427 1931
rect 559 1927 563 1931
rect 703 1927 707 1931
rect 855 1927 859 1931
rect 1239 1943 1243 1947
rect 1391 1943 1395 1947
rect 1399 1943 1403 1947
rect 1807 1940 1811 1944
rect 1863 1939 1867 1943
rect 1999 1939 2003 1943
rect 2143 1939 2147 1943
rect 2287 1939 2291 1943
rect 2431 1939 2435 1943
rect 2575 1939 2579 1943
rect 2711 1939 2715 1943
rect 2831 1939 2835 1943
rect 2951 1939 2955 1943
rect 3063 1939 3067 1943
rect 3167 1939 3171 1943
rect 3279 1939 3283 1943
rect 3367 1939 3371 1943
rect 3463 1940 3467 1944
rect 403 1919 407 1923
rect 495 1919 499 1923
rect 631 1919 635 1923
rect 1007 1927 1011 1931
rect 1159 1927 1163 1931
rect 1311 1927 1315 1931
rect 1471 1927 1475 1931
rect 1767 1928 1771 1932
rect 1935 1931 1939 1935
rect 2079 1931 2083 1935
rect 2359 1931 2363 1935
rect 2367 1931 2371 1935
rect 2655 1931 2659 1935
rect 2799 1931 2803 1935
rect 2911 1931 2915 1935
rect 3135 1931 3139 1935
rect 3239 1931 3243 1935
rect 3247 1931 3251 1935
rect 3359 1931 3363 1935
rect 111 1911 115 1915
rect 775 1915 779 1919
rect 963 1919 967 1923
rect 1231 1915 1235 1919
rect 1239 1919 1243 1923
rect 1391 1919 1395 1923
rect 1807 1923 1811 1927
rect 1863 1920 1867 1924
rect 1999 1920 2003 1924
rect 2143 1920 2147 1924
rect 2287 1920 2291 1924
rect 2431 1920 2435 1924
rect 2575 1920 2579 1924
rect 2639 1923 2643 1927
rect 2711 1920 2715 1924
rect 2831 1920 2835 1924
rect 2951 1920 2955 1924
rect 3063 1920 3067 1924
rect 3167 1920 3171 1924
rect 3279 1920 3283 1924
rect 3367 1920 3371 1924
rect 3463 1923 3467 1927
rect 295 1908 299 1912
rect 423 1908 427 1912
rect 559 1908 563 1912
rect 703 1908 707 1912
rect 855 1908 859 1912
rect 1007 1908 1011 1912
rect 1159 1908 1163 1912
rect 1311 1908 1315 1912
rect 1471 1908 1475 1912
rect 1767 1911 1771 1915
rect 1807 1869 1811 1873
rect 2015 1872 2019 1876
rect 2111 1872 2115 1876
rect 2215 1872 2219 1876
rect 2327 1872 2331 1876
rect 2439 1872 2443 1876
rect 2543 1872 2547 1876
rect 2647 1872 2651 1876
rect 2759 1872 2763 1876
rect 2871 1872 2875 1876
rect 2983 1872 2987 1876
rect 111 1861 115 1865
rect 431 1864 435 1868
rect 575 1864 579 1868
rect 727 1864 731 1868
rect 887 1864 891 1868
rect 1047 1864 1051 1868
rect 1199 1864 1203 1868
rect 1351 1864 1355 1868
rect 1511 1864 1515 1868
rect 3463 1869 3467 1873
rect 1671 1864 1675 1868
rect 1767 1861 1771 1865
rect 2087 1863 2091 1867
rect 2183 1863 2187 1867
rect 2299 1863 2303 1867
rect 2307 1863 2311 1867
rect 2407 1863 2411 1867
rect 2719 1863 2723 1867
rect 2831 1863 2835 1867
rect 2943 1863 2947 1867
rect 503 1855 507 1859
rect 511 1855 515 1859
rect 655 1855 659 1859
rect 951 1855 955 1859
rect 967 1855 971 1859
rect 1271 1855 1275 1859
rect 1423 1855 1427 1859
rect 1583 1855 1587 1859
rect 1735 1855 1739 1859
rect 1807 1852 1811 1856
rect 2015 1853 2019 1857
rect 2111 1853 2115 1857
rect 2215 1853 2219 1857
rect 2327 1853 2331 1857
rect 2439 1853 2443 1857
rect 2543 1853 2547 1857
rect 2647 1853 2651 1857
rect 2759 1853 2763 1857
rect 2871 1853 2875 1857
rect 2983 1853 2987 1857
rect 3463 1852 3467 1856
rect 111 1844 115 1848
rect 431 1845 435 1849
rect 575 1845 579 1849
rect 727 1845 731 1849
rect 887 1845 891 1849
rect 1047 1845 1051 1849
rect 1199 1845 1203 1849
rect 1351 1845 1355 1849
rect 1511 1845 1515 1849
rect 1671 1845 1675 1849
rect 1767 1844 1771 1848
rect 511 1827 515 1831
rect 655 1827 659 1831
rect 775 1827 776 1831
rect 776 1827 779 1831
rect 967 1827 971 1831
rect 1095 1827 1096 1831
rect 1096 1827 1099 1831
rect 1231 1827 1235 1831
rect 1271 1827 1275 1831
rect 1423 1827 1427 1831
rect 1583 1827 1587 1831
rect 2087 1835 2091 1839
rect 2183 1835 2187 1839
rect 2407 1835 2411 1839
rect 2527 1835 2531 1839
rect 2639 1835 2643 1839
rect 2719 1835 2723 1839
rect 2831 1835 2835 1839
rect 2943 1835 2947 1839
rect 2307 1827 2311 1831
rect 503 1811 507 1815
rect 583 1811 587 1815
rect 823 1811 827 1815
rect 831 1811 835 1815
rect 959 1811 963 1815
rect 1359 1819 1363 1823
rect 1223 1811 1227 1815
rect 1487 1811 1491 1815
rect 1615 1811 1619 1815
rect 1735 1811 1739 1815
rect 2207 1815 2211 1819
rect 2263 1815 2267 1819
rect 2351 1815 2355 1819
rect 2711 1823 2715 1827
rect 2615 1815 2619 1819
rect 2887 1815 2891 1819
rect 111 1796 115 1800
rect 511 1795 515 1799
rect 631 1795 635 1799
rect 759 1795 763 1799
rect 887 1795 891 1799
rect 1023 1795 1027 1799
rect 1151 1795 1155 1799
rect 1279 1795 1283 1799
rect 1407 1795 1411 1799
rect 1535 1795 1539 1799
rect 1671 1795 1675 1799
rect 1767 1796 1771 1800
rect 1807 1800 1811 1804
rect 2103 1799 2107 1803
rect 2191 1799 2195 1803
rect 2279 1799 2283 1803
rect 2367 1799 2371 1803
rect 2455 1799 2459 1803
rect 2543 1799 2547 1803
rect 2631 1799 2635 1803
rect 2719 1799 2723 1803
rect 2807 1799 2811 1803
rect 2895 1799 2899 1803
rect 3463 1800 3467 1804
rect 583 1787 587 1791
rect 111 1779 115 1783
rect 703 1783 707 1787
rect 831 1787 835 1791
rect 959 1787 963 1791
rect 1095 1787 1099 1791
rect 1223 1787 1227 1791
rect 1359 1787 1363 1791
rect 1487 1787 1491 1791
rect 1615 1787 1619 1791
rect 2263 1791 2267 1795
rect 2351 1791 2355 1795
rect 2527 1791 2531 1795
rect 2615 1791 2619 1795
rect 511 1776 515 1780
rect 631 1776 635 1780
rect 759 1776 763 1780
rect 887 1776 891 1780
rect 1023 1776 1027 1780
rect 1151 1776 1155 1780
rect 1279 1776 1283 1780
rect 1363 1779 1367 1783
rect 1407 1776 1411 1780
rect 1535 1776 1539 1780
rect 1671 1776 1675 1780
rect 1767 1779 1771 1783
rect 1807 1783 1811 1787
rect 2703 1787 2707 1791
rect 2711 1791 2715 1795
rect 2887 1791 2891 1795
rect 2103 1780 2107 1784
rect 2191 1780 2195 1784
rect 2279 1780 2283 1784
rect 2367 1780 2371 1784
rect 2455 1780 2459 1784
rect 2543 1780 2547 1784
rect 2631 1780 2635 1784
rect 2719 1780 2723 1784
rect 2807 1780 2811 1784
rect 2895 1780 2899 1784
rect 3463 1783 3467 1787
rect 111 1725 115 1729
rect 439 1728 443 1732
rect 535 1728 539 1732
rect 639 1728 643 1732
rect 743 1728 747 1732
rect 847 1728 851 1732
rect 951 1728 955 1732
rect 1055 1728 1059 1732
rect 1159 1728 1163 1732
rect 1271 1728 1275 1732
rect 1383 1728 1387 1732
rect 1767 1725 1771 1729
rect 503 1719 507 1723
rect 519 1719 523 1723
rect 615 1719 619 1723
rect 815 1719 819 1723
rect 823 1719 827 1723
rect 1031 1719 1035 1723
rect 1135 1719 1139 1723
rect 1239 1719 1243 1723
rect 1351 1719 1355 1723
rect 1807 1721 1811 1725
rect 2143 1724 2147 1728
rect 2231 1724 2235 1728
rect 2319 1724 2323 1728
rect 2407 1724 2411 1728
rect 2495 1724 2499 1728
rect 2583 1724 2587 1728
rect 2671 1724 2675 1728
rect 2759 1724 2763 1728
rect 2847 1724 2851 1728
rect 3463 1721 3467 1725
rect 111 1708 115 1712
rect 439 1709 443 1713
rect 535 1709 539 1713
rect 639 1709 643 1713
rect 743 1709 747 1713
rect 847 1709 851 1713
rect 951 1709 955 1713
rect 2207 1715 2211 1719
rect 2223 1715 2227 1719
rect 2311 1715 2315 1719
rect 2399 1715 2403 1719
rect 2487 1715 2491 1719
rect 2647 1715 2651 1719
rect 2743 1715 2747 1719
rect 2831 1715 2835 1719
rect 1055 1709 1059 1713
rect 1159 1709 1163 1713
rect 1271 1709 1275 1713
rect 1383 1709 1387 1713
rect 1767 1708 1771 1712
rect 1079 1703 1083 1707
rect 1807 1704 1811 1708
rect 2143 1705 2147 1709
rect 2231 1705 2235 1709
rect 2319 1705 2323 1709
rect 2407 1705 2411 1709
rect 2495 1705 2499 1709
rect 2583 1705 2587 1709
rect 2671 1705 2675 1709
rect 2759 1705 2763 1709
rect 2847 1705 2851 1709
rect 3463 1704 3467 1708
rect 519 1691 523 1695
rect 615 1691 619 1695
rect 703 1691 707 1695
rect 735 1691 739 1695
rect 815 1691 819 1695
rect 1031 1691 1035 1695
rect 1135 1691 1139 1695
rect 1239 1691 1243 1695
rect 1351 1691 1355 1695
rect 1363 1691 1367 1695
rect 503 1675 507 1679
rect 671 1675 675 1679
rect 839 1675 843 1679
rect 1127 1683 1131 1687
rect 2223 1687 2227 1691
rect 2311 1687 2315 1691
rect 2399 1687 2403 1691
rect 2487 1687 2491 1691
rect 2527 1687 2531 1691
rect 1083 1675 1087 1679
rect 1119 1675 1123 1679
rect 2447 1679 2451 1683
rect 2703 1687 2707 1691
rect 2743 1687 2747 1691
rect 2831 1687 2835 1691
rect 2175 1671 2179 1675
rect 2263 1671 2267 1675
rect 2351 1671 2355 1675
rect 2439 1671 2443 1675
rect 2647 1671 2651 1675
rect 111 1660 115 1664
rect 399 1659 403 1663
rect 487 1659 491 1663
rect 575 1659 579 1663
rect 2703 1671 2707 1675
rect 2791 1671 2795 1675
rect 2879 1671 2883 1675
rect 663 1659 667 1663
rect 759 1659 763 1663
rect 855 1659 859 1663
rect 951 1659 955 1663
rect 1047 1659 1051 1663
rect 1143 1659 1147 1663
rect 1767 1660 1771 1664
rect 1807 1656 1811 1660
rect 111 1643 115 1647
rect 559 1647 563 1651
rect 735 1651 739 1655
rect 839 1651 843 1655
rect 1119 1651 1123 1655
rect 2103 1655 2107 1659
rect 1127 1651 1131 1655
rect 2191 1655 2195 1659
rect 2279 1655 2283 1659
rect 2367 1655 2371 1659
rect 2455 1655 2459 1659
rect 2543 1655 2547 1659
rect 399 1640 403 1644
rect 487 1640 491 1644
rect 575 1640 579 1644
rect 663 1640 667 1644
rect 759 1640 763 1644
rect 839 1643 843 1647
rect 855 1640 859 1644
rect 951 1640 955 1644
rect 1047 1640 1051 1644
rect 1143 1640 1147 1644
rect 1767 1643 1771 1647
rect 2175 1647 2179 1651
rect 2263 1647 2267 1651
rect 2351 1647 2355 1651
rect 2439 1647 2443 1651
rect 2527 1647 2531 1651
rect 2631 1655 2635 1659
rect 2719 1655 2723 1659
rect 2807 1655 2811 1659
rect 2895 1655 2899 1659
rect 3463 1656 3467 1660
rect 2703 1647 2707 1651
rect 2791 1647 2795 1651
rect 2879 1647 2883 1651
rect 1807 1639 1811 1643
rect 2103 1636 2107 1640
rect 2191 1636 2195 1640
rect 2279 1636 2283 1640
rect 2367 1636 2371 1640
rect 2455 1636 2459 1640
rect 2543 1636 2547 1640
rect 2631 1636 2635 1640
rect 2719 1636 2723 1640
rect 2807 1636 2811 1640
rect 2895 1636 2899 1640
rect 3463 1639 3467 1643
rect 2619 1603 2623 1607
rect 111 1589 115 1593
rect 279 1592 283 1596
rect 383 1592 387 1596
rect 495 1592 499 1596
rect 607 1592 611 1596
rect 719 1592 723 1596
rect 831 1592 835 1596
rect 943 1592 947 1596
rect 1055 1592 1059 1596
rect 1167 1592 1171 1596
rect 1279 1592 1283 1596
rect 2603 1595 2607 1599
rect 1767 1589 1771 1593
rect 351 1583 355 1587
rect 455 1583 459 1587
rect 463 1583 467 1587
rect 671 1583 675 1587
rect 687 1583 691 1587
rect 903 1583 907 1587
rect 1015 1583 1019 1587
rect 1127 1583 1131 1587
rect 1239 1583 1243 1587
rect 1247 1583 1251 1587
rect 1807 1585 1811 1589
rect 2063 1588 2067 1592
rect 2159 1588 2163 1592
rect 2255 1588 2259 1592
rect 2359 1588 2363 1592
rect 2463 1588 2467 1592
rect 2567 1588 2571 1592
rect 2671 1588 2675 1592
rect 2775 1588 2779 1592
rect 2135 1579 2139 1583
rect 2231 1579 2235 1583
rect 2327 1579 2331 1583
rect 2431 1579 2435 1583
rect 2447 1579 2451 1583
rect 2639 1579 2643 1583
rect 2743 1579 2747 1583
rect 2847 1579 2851 1583
rect 2887 1588 2891 1592
rect 3463 1585 3467 1589
rect 111 1572 115 1576
rect 279 1573 283 1577
rect 383 1573 387 1577
rect 495 1573 499 1577
rect 607 1573 611 1577
rect 719 1573 723 1577
rect 831 1573 835 1577
rect 943 1573 947 1577
rect 1055 1573 1059 1577
rect 1167 1573 1171 1577
rect 1279 1573 1283 1577
rect 1767 1572 1771 1576
rect 1807 1568 1811 1572
rect 2063 1569 2067 1573
rect 2159 1569 2163 1573
rect 2255 1569 2259 1573
rect 2359 1569 2363 1573
rect 2463 1569 2467 1573
rect 2567 1569 2571 1573
rect 2671 1569 2675 1573
rect 2775 1569 2779 1573
rect 2887 1569 2891 1573
rect 3463 1568 3467 1572
rect 351 1555 355 1559
rect 559 1555 563 1559
rect 687 1555 691 1559
rect 695 1555 699 1559
rect 839 1555 843 1559
rect 903 1555 907 1559
rect 1015 1555 1019 1559
rect 1127 1555 1131 1559
rect 1239 1555 1243 1559
rect 463 1547 467 1551
rect 2111 1551 2112 1555
rect 2112 1551 2115 1555
rect 2135 1551 2139 1555
rect 2231 1551 2235 1555
rect 2327 1551 2331 1555
rect 2431 1551 2435 1555
rect 2619 1551 2620 1555
rect 2620 1551 2623 1555
rect 2639 1551 2643 1555
rect 2743 1551 2747 1555
rect 2847 1551 2851 1555
rect 291 1535 295 1539
rect 407 1535 411 1539
rect 455 1535 459 1539
rect 703 1535 707 1539
rect 847 1535 851 1539
rect 1247 1543 1251 1547
rect 1119 1535 1123 1539
rect 1247 1535 1251 1539
rect 1383 1535 1387 1539
rect 1983 1539 1987 1543
rect 1991 1539 1995 1543
rect 2111 1539 2115 1543
rect 2239 1539 2243 1543
rect 2367 1539 2371 1543
rect 2603 1539 2604 1543
rect 2604 1539 2607 1543
rect 2623 1539 2627 1543
rect 2751 1539 2755 1543
rect 2871 1539 2875 1543
rect 2999 1539 3003 1543
rect 111 1520 115 1524
rect 183 1519 187 1523
rect 327 1519 331 1523
rect 471 1519 475 1523
rect 623 1519 627 1523
rect 767 1519 771 1523
rect 911 1519 915 1523
rect 111 1503 115 1507
rect 255 1507 259 1511
rect 291 1511 295 1515
rect 407 1511 411 1515
rect 695 1511 699 1515
rect 703 1511 707 1515
rect 1047 1519 1051 1523
rect 1175 1519 1179 1523
rect 1311 1519 1315 1523
rect 1447 1519 1451 1523
rect 1767 1520 1771 1524
rect 1807 1524 1811 1528
rect 1919 1523 1923 1527
rect 2039 1523 2043 1527
rect 2167 1523 2171 1527
rect 2295 1523 2299 1527
rect 2423 1523 2427 1527
rect 2551 1523 2555 1527
rect 2679 1523 2683 1527
rect 2799 1523 2803 1527
rect 2927 1523 2931 1527
rect 3055 1523 3059 1527
rect 3463 1524 3467 1528
rect 1119 1511 1123 1515
rect 1247 1511 1251 1515
rect 1383 1511 1387 1515
rect 1399 1511 1403 1515
rect 1991 1515 1995 1519
rect 2111 1515 2115 1519
rect 2239 1515 2243 1519
rect 2367 1515 2371 1519
rect 2375 1515 2379 1519
rect 2623 1515 2627 1519
rect 2751 1515 2755 1519
rect 2871 1515 2875 1519
rect 2999 1515 3003 1519
rect 3019 1515 3023 1519
rect 183 1500 187 1504
rect 327 1500 331 1504
rect 471 1500 475 1504
rect 623 1500 627 1504
rect 767 1500 771 1504
rect 911 1500 915 1504
rect 1047 1500 1051 1504
rect 1175 1500 1179 1504
rect 1311 1500 1315 1504
rect 1447 1500 1451 1504
rect 1767 1503 1771 1507
rect 1807 1507 1811 1511
rect 1919 1504 1923 1508
rect 2039 1504 2043 1508
rect 2167 1504 2171 1508
rect 2295 1504 2299 1508
rect 2423 1504 2427 1508
rect 2551 1504 2555 1508
rect 2679 1504 2683 1508
rect 2799 1504 2803 1508
rect 2927 1504 2931 1508
rect 3055 1504 3059 1508
rect 3463 1507 3467 1511
rect 2119 1495 2123 1499
rect 2375 1495 2379 1499
rect 1067 1459 1071 1463
rect 111 1449 115 1453
rect 159 1452 163 1456
rect 375 1452 379 1456
rect 583 1452 587 1456
rect 783 1452 787 1456
rect 959 1452 963 1456
rect 1127 1452 1131 1456
rect 1279 1452 1283 1456
rect 1431 1452 1435 1456
rect 263 1443 267 1447
rect 447 1443 451 1447
rect 655 1443 659 1447
rect 847 1443 851 1447
rect 1091 1443 1095 1447
rect 1199 1443 1203 1447
rect 1351 1443 1355 1447
rect 1503 1443 1507 1447
rect 1983 1459 1987 1463
rect 1591 1452 1595 1456
rect 1767 1449 1771 1453
rect 1807 1449 1811 1453
rect 1831 1452 1835 1456
rect 1951 1452 1955 1456
rect 2111 1452 2115 1456
rect 2271 1452 2275 1456
rect 2023 1443 2027 1447
rect 2183 1443 2187 1447
rect 2343 1443 2347 1447
rect 2611 1459 2615 1463
rect 2431 1452 2435 1456
rect 2591 1452 2595 1456
rect 2735 1452 2739 1456
rect 2871 1452 2875 1456
rect 3007 1452 3011 1456
rect 2807 1443 2811 1447
rect 2943 1443 2947 1447
rect 3079 1443 3083 1447
rect 3135 1452 3139 1456
rect 3263 1452 3267 1456
rect 3367 1452 3371 1456
rect 3463 1449 3467 1453
rect 3335 1443 3339 1447
rect 3431 1443 3435 1447
rect 111 1432 115 1436
rect 159 1433 163 1437
rect 375 1433 379 1437
rect 583 1433 587 1437
rect 783 1433 787 1437
rect 959 1433 963 1437
rect 1127 1433 1131 1437
rect 1279 1433 1283 1437
rect 1431 1433 1435 1437
rect 1591 1433 1595 1437
rect 1767 1432 1771 1436
rect 1807 1432 1811 1436
rect 1831 1433 1835 1437
rect 1951 1433 1955 1437
rect 2111 1433 2115 1437
rect 2271 1433 2275 1437
rect 2431 1433 2435 1437
rect 2591 1433 2595 1437
rect 2735 1433 2739 1437
rect 2871 1433 2875 1437
rect 3007 1433 3011 1437
rect 3135 1433 3139 1437
rect 3263 1433 3267 1437
rect 3367 1433 3371 1437
rect 3463 1432 3467 1436
rect 255 1415 259 1419
rect 263 1415 267 1419
rect 635 1415 636 1419
rect 636 1415 639 1419
rect 655 1415 659 1419
rect 1091 1415 1095 1419
rect 1199 1415 1203 1419
rect 1351 1415 1355 1419
rect 1503 1415 1507 1419
rect 1399 1407 1403 1411
rect 1743 1407 1747 1411
rect 2023 1415 2027 1419
rect 2183 1415 2187 1419
rect 2343 1415 2347 1419
rect 283 1399 287 1403
rect 447 1399 451 1403
rect 759 1399 763 1403
rect 975 1399 979 1403
rect 1067 1399 1068 1403
rect 1068 1399 1071 1403
rect 1087 1399 1091 1403
rect 1239 1399 1243 1403
rect 1375 1399 1379 1403
rect 1503 1399 1507 1403
rect 1751 1399 1755 1403
rect 1895 1399 1899 1403
rect 2343 1407 2347 1411
rect 2807 1415 2811 1419
rect 2943 1415 2947 1419
rect 3079 1415 3083 1419
rect 3327 1415 3331 1419
rect 3335 1415 3339 1419
rect 3019 1407 3023 1411
rect 2079 1399 2083 1403
rect 2335 1399 2339 1403
rect 2611 1399 2612 1403
rect 2612 1399 2615 1403
rect 2631 1399 2635 1403
rect 2791 1399 2795 1403
rect 2935 1399 2939 1403
rect 3071 1399 3075 1403
rect 3199 1399 3203 1403
rect 3431 1399 3435 1403
rect 111 1384 115 1388
rect 135 1383 139 1387
rect 303 1383 307 1387
rect 495 1383 499 1387
rect 679 1383 683 1387
rect 855 1383 859 1387
rect 1015 1383 1019 1387
rect 1167 1383 1171 1387
rect 1303 1383 1307 1387
rect 1431 1383 1435 1387
rect 1559 1383 1563 1387
rect 1671 1383 1675 1387
rect 1767 1384 1771 1388
rect 1807 1384 1811 1388
rect 1831 1383 1835 1387
rect 2007 1383 2011 1387
rect 2199 1383 2203 1387
rect 2383 1383 2387 1387
rect 2559 1383 2563 1387
rect 2719 1383 2723 1387
rect 2863 1383 2867 1387
rect 2999 1383 3003 1387
rect 3127 1383 3131 1387
rect 3255 1383 3259 1387
rect 3367 1383 3371 1387
rect 3463 1384 3467 1388
rect 283 1375 287 1379
rect 635 1375 639 1379
rect 759 1375 763 1379
rect 1087 1375 1091 1379
rect 1239 1375 1243 1379
rect 1375 1375 1379 1379
rect 1503 1375 1507 1379
rect 1511 1375 1515 1379
rect 1743 1375 1747 1379
rect 1751 1375 1755 1379
rect 2079 1375 2083 1379
rect 2335 1375 2339 1379
rect 2343 1375 2347 1379
rect 2631 1375 2635 1379
rect 2791 1375 2795 1379
rect 2935 1375 2939 1379
rect 3071 1375 3075 1379
rect 3199 1375 3203 1379
rect 3327 1375 3331 1379
rect 111 1367 115 1371
rect 135 1364 139 1368
rect 199 1367 203 1371
rect 303 1364 307 1368
rect 495 1364 499 1368
rect 679 1364 683 1368
rect 855 1364 859 1368
rect 1015 1364 1019 1368
rect 1167 1364 1171 1368
rect 1303 1364 1307 1368
rect 1431 1364 1435 1368
rect 1559 1364 1563 1368
rect 1671 1364 1675 1368
rect 1767 1367 1771 1371
rect 1807 1367 1811 1371
rect 3439 1371 3443 1375
rect 1831 1364 1835 1368
rect 2007 1364 2011 1368
rect 2199 1364 2203 1368
rect 2383 1364 2387 1368
rect 2559 1364 2563 1368
rect 2719 1364 2723 1368
rect 2863 1364 2867 1368
rect 2999 1364 3003 1368
rect 3127 1364 3131 1368
rect 3255 1364 3259 1368
rect 3367 1364 3371 1368
rect 3463 1367 3467 1371
rect 111 1313 115 1317
rect 135 1316 139 1320
rect 247 1316 251 1320
rect 399 1316 403 1320
rect 559 1316 563 1320
rect 727 1316 731 1320
rect 895 1316 899 1320
rect 1063 1316 1067 1320
rect 1223 1316 1227 1320
rect 1375 1316 1379 1320
rect 1535 1316 1539 1320
rect 1671 1316 1675 1320
rect 2019 1319 2023 1323
rect 1767 1313 1771 1317
rect 207 1307 211 1311
rect 319 1307 323 1311
rect 471 1307 475 1311
rect 499 1307 503 1311
rect 799 1307 803 1311
rect 967 1307 971 1311
rect 975 1307 979 1311
rect 1295 1307 1299 1311
rect 1447 1307 1451 1311
rect 1607 1307 1611 1311
rect 1623 1307 1627 1311
rect 1807 1309 1811 1313
rect 1831 1312 1835 1316
rect 1967 1312 1971 1316
rect 2143 1312 2147 1316
rect 2327 1312 2331 1316
rect 1895 1303 1899 1307
rect 1911 1303 1915 1307
rect 2215 1303 2219 1307
rect 2399 1303 2403 1307
rect 2511 1312 2515 1316
rect 2687 1312 2691 1316
rect 2863 1312 2867 1316
rect 3039 1312 3043 1316
rect 3215 1312 3219 1316
rect 3367 1312 3371 1316
rect 3463 1309 3467 1313
rect 2759 1303 2763 1307
rect 2767 1303 2771 1307
rect 2943 1303 2947 1307
rect 3119 1303 3123 1307
rect 3431 1303 3435 1307
rect 111 1296 115 1300
rect 135 1297 139 1301
rect 247 1297 251 1301
rect 399 1297 403 1301
rect 559 1297 563 1301
rect 727 1297 731 1301
rect 895 1297 899 1301
rect 1063 1297 1067 1301
rect 1223 1297 1227 1301
rect 1375 1297 1379 1301
rect 1535 1297 1539 1301
rect 1671 1297 1675 1301
rect 1767 1296 1771 1300
rect 1807 1292 1811 1296
rect 1831 1293 1835 1297
rect 1967 1293 1971 1297
rect 2143 1293 2147 1297
rect 2327 1293 2331 1297
rect 2511 1293 2515 1297
rect 2687 1293 2691 1297
rect 2863 1293 2867 1297
rect 3039 1293 3043 1297
rect 3215 1293 3219 1297
rect 3367 1293 3371 1297
rect 3463 1292 3467 1296
rect 199 1279 203 1283
rect 207 1279 211 1283
rect 319 1279 323 1283
rect 471 1279 475 1283
rect 751 1279 755 1283
rect 799 1279 803 1283
rect 967 1279 971 1283
rect 1295 1279 1299 1283
rect 1447 1279 1451 1283
rect 1607 1279 1611 1283
rect 1511 1271 1515 1275
rect 187 1263 188 1267
rect 188 1263 191 1267
rect 207 1263 211 1267
rect 295 1263 299 1267
rect 391 1263 395 1267
rect 503 1263 507 1267
rect 759 1263 763 1267
rect 903 1263 907 1267
rect 1091 1263 1095 1267
rect 1327 1263 1331 1267
rect 1623 1271 1627 1275
rect 1911 1275 1915 1279
rect 2019 1275 2020 1279
rect 2020 1275 2023 1279
rect 2167 1275 2171 1279
rect 2215 1275 2219 1279
rect 2399 1275 2403 1279
rect 1575 1263 1579 1267
rect 1743 1263 1747 1267
rect 1903 1263 1907 1267
rect 2679 1271 2683 1275
rect 2767 1275 2771 1279
rect 2943 1275 2947 1279
rect 3119 1275 3123 1279
rect 3263 1275 3264 1279
rect 3264 1275 3267 1279
rect 3439 1275 3443 1279
rect 2431 1263 2435 1267
rect 2759 1263 2763 1267
rect 3087 1263 3091 1267
rect 3147 1263 3151 1267
rect 3431 1263 3435 1267
rect 111 1248 115 1252
rect 135 1247 139 1251
rect 223 1247 227 1251
rect 319 1247 323 1251
rect 431 1247 435 1251
rect 551 1247 555 1251
rect 679 1247 683 1251
rect 823 1247 827 1251
rect 975 1247 979 1251
rect 1143 1247 1147 1251
rect 1319 1247 1323 1251
rect 1503 1247 1507 1251
rect 1671 1247 1675 1251
rect 1767 1248 1771 1252
rect 1807 1248 1811 1252
rect 1831 1247 1835 1251
rect 2095 1247 2099 1251
rect 2359 1247 2363 1251
rect 2599 1247 2603 1251
rect 2807 1247 2811 1251
rect 3007 1247 3011 1251
rect 3199 1247 3203 1251
rect 207 1239 211 1243
rect 295 1239 299 1243
rect 391 1239 395 1243
rect 503 1239 507 1243
rect 511 1239 515 1243
rect 751 1239 755 1243
rect 759 1239 763 1243
rect 903 1239 907 1243
rect 1091 1239 1095 1243
rect 1575 1239 1579 1243
rect 1743 1239 1747 1243
rect 1903 1239 1907 1243
rect 2167 1239 2171 1243
rect 2431 1239 2435 1243
rect 111 1231 115 1235
rect 135 1228 139 1232
rect 223 1228 227 1232
rect 319 1228 323 1232
rect 431 1228 435 1232
rect 551 1228 555 1232
rect 679 1228 683 1232
rect 823 1228 827 1232
rect 975 1228 979 1232
rect 1143 1228 1147 1232
rect 1319 1228 1323 1232
rect 1503 1228 1507 1232
rect 1671 1228 1675 1232
rect 1767 1231 1771 1235
rect 1807 1231 1811 1235
rect 2671 1235 2675 1239
rect 2679 1239 2683 1243
rect 3147 1239 3151 1243
rect 3263 1243 3267 1247
rect 3367 1247 3371 1251
rect 3463 1248 3467 1252
rect 3439 1235 3443 1239
rect 1831 1228 1835 1232
rect 2095 1228 2099 1232
rect 2359 1228 2363 1232
rect 2599 1228 2603 1232
rect 2807 1228 2811 1232
rect 3007 1228 3011 1232
rect 3199 1228 3203 1232
rect 3367 1228 3371 1232
rect 3463 1231 3467 1235
rect 187 1191 191 1195
rect 511 1191 515 1195
rect 111 1173 115 1177
rect 135 1176 139 1180
rect 231 1176 235 1180
rect 359 1176 363 1180
rect 487 1176 491 1180
rect 615 1176 619 1180
rect 743 1176 747 1180
rect 871 1176 875 1180
rect 991 1176 995 1180
rect 1119 1176 1123 1180
rect 1247 1176 1251 1180
rect 1767 1173 1771 1177
rect 1807 1173 1811 1177
rect 1935 1176 1939 1180
rect 2039 1176 2043 1180
rect 2159 1176 2163 1180
rect 2287 1176 2291 1180
rect 2423 1176 2427 1180
rect 2567 1176 2571 1180
rect 2703 1176 2707 1180
rect 2839 1176 2843 1180
rect 2975 1176 2979 1180
rect 3111 1176 3115 1180
rect 3247 1176 3251 1180
rect 3367 1176 3371 1180
rect 3463 1173 3467 1177
rect 207 1167 211 1171
rect 303 1167 307 1171
rect 431 1167 435 1171
rect 559 1167 563 1171
rect 567 1167 571 1171
rect 815 1167 819 1171
rect 943 1167 947 1171
rect 1063 1167 1067 1171
rect 1191 1167 1195 1171
rect 1327 1167 1331 1171
rect 2003 1167 2007 1171
rect 2015 1167 2019 1171
rect 2119 1167 2123 1171
rect 2239 1167 2243 1171
rect 2367 1167 2371 1171
rect 2503 1167 2507 1171
rect 2775 1167 2779 1171
rect 2911 1167 2915 1171
rect 3047 1167 3051 1171
rect 3087 1167 3091 1171
rect 3191 1167 3195 1171
rect 3431 1167 3435 1171
rect 111 1156 115 1160
rect 135 1157 139 1161
rect 231 1157 235 1161
rect 359 1157 363 1161
rect 487 1157 491 1161
rect 615 1157 619 1161
rect 743 1157 747 1161
rect 871 1157 875 1161
rect 991 1157 995 1161
rect 1119 1157 1123 1161
rect 1247 1157 1251 1161
rect 1767 1156 1771 1160
rect 1807 1156 1811 1160
rect 1935 1157 1939 1161
rect 2039 1157 2043 1161
rect 2159 1157 2163 1161
rect 2287 1157 2291 1161
rect 2423 1157 2427 1161
rect 2567 1157 2571 1161
rect 2703 1157 2707 1161
rect 2839 1157 2843 1161
rect 2975 1157 2979 1161
rect 3111 1157 3115 1161
rect 3247 1157 3251 1161
rect 3367 1157 3371 1161
rect 3463 1156 3467 1160
rect 187 1139 188 1143
rect 188 1139 191 1143
rect 207 1139 211 1143
rect 303 1139 307 1143
rect 431 1139 435 1143
rect 559 1139 563 1143
rect 567 1131 571 1135
rect 815 1139 819 1143
rect 943 1139 947 1143
rect 1063 1139 1067 1143
rect 1191 1139 1195 1143
rect 2015 1139 2019 1143
rect 2119 1139 2123 1143
rect 2239 1139 2243 1143
rect 2367 1139 2371 1143
rect 2503 1139 2507 1143
rect 2527 1139 2531 1143
rect 2671 1139 2675 1143
rect 2775 1139 2779 1143
rect 2911 1139 2915 1143
rect 3191 1139 3195 1143
rect 3295 1139 3296 1143
rect 3296 1139 3299 1143
rect 3439 1139 3443 1143
rect 839 1131 843 1135
rect 319 1123 323 1127
rect 439 1123 443 1127
rect 567 1123 571 1127
rect 695 1123 699 1127
rect 999 1123 1003 1127
rect 1111 1123 1115 1127
rect 1223 1123 1227 1127
rect 1351 1123 1355 1127
rect 1383 1123 1387 1127
rect 2003 1123 2007 1127
rect 2015 1119 2019 1123
rect 2135 1119 2139 1123
rect 2371 1119 2372 1123
rect 2372 1119 2375 1123
rect 2391 1119 2395 1123
rect 2831 1127 2835 1131
rect 2671 1119 2675 1123
rect 2983 1119 2987 1123
rect 3047 1119 3051 1123
rect 3271 1119 3272 1123
rect 3272 1119 3275 1123
rect 3431 1119 3435 1123
rect 111 1108 115 1112
rect 247 1107 251 1111
rect 367 1107 371 1111
rect 495 1107 499 1111
rect 623 1107 627 1111
rect 759 1107 763 1111
rect 887 1107 891 1111
rect 1015 1107 1019 1111
rect 1143 1107 1147 1111
rect 1271 1107 1275 1111
rect 1399 1107 1403 1111
rect 1767 1108 1771 1112
rect 1807 1104 1811 1108
rect 319 1099 323 1103
rect 439 1099 443 1103
rect 567 1099 571 1103
rect 695 1099 699 1103
rect 703 1099 707 1103
rect 839 1099 843 1103
rect 999 1099 1003 1103
rect 1111 1099 1115 1103
rect 1223 1099 1227 1103
rect 1943 1103 1947 1107
rect 1351 1099 1355 1103
rect 2063 1103 2067 1107
rect 2191 1103 2195 1107
rect 2319 1103 2323 1107
rect 2455 1103 2459 1107
rect 2599 1103 2603 1107
rect 2751 1103 2755 1107
rect 2903 1103 2907 1107
rect 3063 1103 3067 1107
rect 3223 1103 3227 1107
rect 3367 1103 3371 1107
rect 3463 1104 3467 1108
rect 111 1091 115 1095
rect 247 1088 251 1092
rect 367 1088 371 1092
rect 495 1088 499 1092
rect 623 1088 627 1092
rect 759 1088 763 1092
rect 887 1088 891 1092
rect 1015 1088 1019 1092
rect 1143 1088 1147 1092
rect 1271 1088 1275 1092
rect 1399 1088 1403 1092
rect 1767 1091 1771 1095
rect 2015 1095 2019 1099
rect 2135 1095 2139 1099
rect 2171 1095 2175 1099
rect 2391 1095 2395 1099
rect 2527 1095 2531 1099
rect 2671 1095 2675 1099
rect 1807 1087 1811 1091
rect 2823 1091 2827 1095
rect 2831 1095 2835 1099
rect 2983 1095 2987 1099
rect 3295 1095 3299 1099
rect 3439 1091 3443 1095
rect 1943 1084 1947 1088
rect 2063 1084 2067 1088
rect 2191 1084 2195 1088
rect 2319 1084 2323 1088
rect 2455 1084 2459 1088
rect 2599 1084 2603 1088
rect 2751 1084 2755 1088
rect 2903 1084 2907 1088
rect 3063 1084 3067 1088
rect 3223 1084 3227 1088
rect 3367 1084 3371 1088
rect 3463 1087 3467 1091
rect 483 1055 487 1059
rect 703 1055 707 1059
rect 1091 1047 1095 1051
rect 111 1037 115 1041
rect 431 1040 435 1044
rect 543 1040 547 1044
rect 663 1040 667 1044
rect 791 1040 795 1044
rect 919 1040 923 1044
rect 1039 1040 1043 1044
rect 1159 1040 1163 1044
rect 1279 1040 1283 1044
rect 1407 1040 1411 1044
rect 503 1031 507 1035
rect 615 1031 619 1035
rect 735 1031 739 1035
rect 863 1031 867 1035
rect 871 1031 875 1035
rect 1111 1031 1115 1035
rect 1231 1031 1235 1035
rect 1383 1031 1387 1035
rect 1479 1031 1483 1035
rect 1535 1040 1539 1044
rect 2595 1043 2599 1047
rect 1767 1037 1771 1041
rect 1807 1033 1811 1037
rect 1847 1036 1851 1040
rect 1983 1036 1987 1040
rect 2119 1036 2123 1040
rect 2255 1036 2259 1040
rect 2391 1036 2395 1040
rect 2543 1036 2547 1040
rect 2703 1036 2707 1040
rect 2863 1036 2867 1040
rect 1927 1027 1931 1031
rect 2063 1027 2067 1031
rect 2371 1027 2375 1031
rect 2615 1027 2619 1031
rect 2775 1027 2779 1031
rect 2935 1027 2939 1031
rect 3031 1036 3035 1040
rect 3207 1036 3211 1040
rect 3367 1036 3371 1040
rect 3463 1033 3467 1037
rect 3271 1027 3275 1031
rect 3431 1027 3435 1031
rect 111 1020 115 1024
rect 431 1021 435 1025
rect 543 1021 547 1025
rect 663 1021 667 1025
rect 791 1021 795 1025
rect 919 1021 923 1025
rect 1039 1021 1043 1025
rect 1159 1021 1163 1025
rect 1279 1021 1283 1025
rect 1407 1021 1411 1025
rect 1535 1021 1539 1025
rect 1767 1020 1771 1024
rect 1807 1016 1811 1020
rect 1847 1017 1851 1021
rect 1983 1017 1987 1021
rect 2119 1017 2123 1021
rect 2255 1017 2259 1021
rect 2391 1017 2395 1021
rect 2543 1017 2547 1021
rect 2703 1017 2707 1021
rect 2863 1017 2867 1021
rect 3031 1017 3035 1021
rect 3207 1017 3211 1021
rect 3367 1017 3371 1021
rect 3463 1016 3467 1020
rect 483 1003 484 1007
rect 484 1003 487 1007
rect 503 1003 507 1007
rect 615 1003 619 1007
rect 735 1003 739 1007
rect 863 1003 867 1007
rect 1091 1003 1092 1007
rect 1092 1003 1095 1007
rect 1111 1003 1115 1007
rect 1231 1003 1235 1007
rect 1431 1003 1435 1007
rect 1479 1003 1483 1007
rect 1927 999 1931 1003
rect 2063 999 2067 1003
rect 2171 999 2172 1003
rect 2172 999 2175 1003
rect 2367 999 2371 1003
rect 2595 999 2596 1003
rect 2596 999 2599 1003
rect 2615 999 2619 1003
rect 2823 999 2827 1003
rect 2935 999 2939 1003
rect 3255 999 3256 1003
rect 3256 999 3259 1003
rect 3439 999 3443 1003
rect 871 991 875 995
rect 639 983 643 987
rect 751 983 755 987
rect 863 983 867 987
rect 983 983 987 987
rect 1439 991 1443 995
rect 1215 983 1219 987
rect 1327 983 1331 987
rect 1523 983 1524 987
rect 1524 983 1527 987
rect 1663 983 1667 987
rect 1751 983 1755 987
rect 1939 983 1943 987
rect 2419 991 2423 995
rect 2959 991 2963 995
rect 2471 983 2475 987
rect 2775 979 2779 983
rect 2879 983 2883 987
rect 3295 983 3299 987
rect 3431 983 3435 987
rect 111 968 115 972
rect 567 967 571 971
rect 679 967 683 971
rect 791 967 795 971
rect 911 967 915 971
rect 1031 967 1035 971
rect 1143 967 1147 971
rect 1255 967 1259 971
rect 1359 967 1363 971
rect 1471 967 1475 971
rect 1583 967 1587 971
rect 1671 967 1675 971
rect 1767 968 1771 972
rect 1807 968 1811 972
rect 1831 967 1835 971
rect 1975 967 1979 971
rect 2135 967 2139 971
rect 2295 967 2299 971
rect 2463 967 2467 971
rect 2631 967 2635 971
rect 2807 967 2811 971
rect 2991 967 2995 971
rect 3183 967 3187 971
rect 3367 967 3371 971
rect 3463 968 3467 972
rect 639 959 643 963
rect 751 959 755 963
rect 863 959 867 963
rect 983 959 987 963
rect 991 959 995 963
rect 1215 959 1219 963
rect 1327 959 1331 963
rect 1431 959 1435 963
rect 1439 959 1443 963
rect 111 951 115 955
rect 1655 955 1659 959
rect 1663 959 1667 963
rect 1751 959 1755 963
rect 1939 959 1943 963
rect 567 948 571 952
rect 679 948 683 952
rect 791 948 795 952
rect 911 948 915 952
rect 1031 948 1035 952
rect 1143 948 1147 952
rect 1255 948 1259 952
rect 1359 948 1363 952
rect 1471 948 1475 952
rect 1583 948 1587 952
rect 1671 948 1675 952
rect 1767 951 1771 955
rect 1807 951 1811 955
rect 2207 955 2211 959
rect 2367 959 2371 963
rect 2419 959 2423 963
rect 2879 959 2883 963
rect 2959 959 2963 963
rect 3255 959 3259 963
rect 3439 955 3443 959
rect 1831 948 1835 952
rect 1975 948 1979 952
rect 2135 948 2139 952
rect 2295 948 2299 952
rect 2463 948 2467 952
rect 2631 948 2635 952
rect 2807 948 2811 952
rect 2991 948 2995 952
rect 3183 948 3187 952
rect 3367 948 3371 952
rect 3463 951 3467 955
rect 111 897 115 901
rect 415 900 419 904
rect 559 900 563 904
rect 727 900 731 904
rect 911 900 915 904
rect 1119 900 1123 904
rect 1335 900 1339 904
rect 1559 900 1563 904
rect 1767 897 1771 901
rect 1807 901 1811 905
rect 2127 904 2131 908
rect 2215 904 2219 908
rect 2303 904 2307 908
rect 2391 904 2395 908
rect 2479 904 2483 908
rect 2567 904 2571 908
rect 2655 904 2659 908
rect 2743 904 2747 908
rect 2831 904 2835 908
rect 3463 901 3467 905
rect 487 891 491 895
rect 631 891 635 895
rect 679 891 683 895
rect 807 891 811 895
rect 1191 891 1195 895
rect 1323 891 1327 895
rect 1523 891 1527 895
rect 2287 895 2291 899
rect 2375 895 2379 899
rect 2463 895 2467 899
rect 2471 895 2475 899
rect 2639 895 2643 899
rect 2727 895 2731 899
rect 2815 895 2819 899
rect 2823 895 2827 899
rect 111 880 115 884
rect 415 881 419 885
rect 559 881 563 885
rect 727 881 731 885
rect 911 881 915 885
rect 1119 881 1123 885
rect 1335 881 1339 885
rect 1559 881 1563 885
rect 1767 880 1771 884
rect 1807 884 1811 888
rect 2127 885 2131 889
rect 2215 885 2219 889
rect 2303 885 2307 889
rect 2391 885 2395 889
rect 2479 885 2483 889
rect 2567 885 2571 889
rect 2655 885 2659 889
rect 2743 885 2747 889
rect 2831 885 2835 889
rect 3463 884 3467 888
rect 487 863 491 867
rect 807 863 811 867
rect 991 863 995 867
rect 1191 863 1195 867
rect 1655 863 1659 867
rect 2207 867 2211 871
rect 2287 867 2291 871
rect 2375 867 2379 871
rect 2519 867 2523 871
rect 679 855 683 859
rect 1231 855 1235 859
rect 2463 859 2467 863
rect 2639 867 2643 871
rect 2727 867 2731 871
rect 2815 867 2819 871
rect 215 847 219 851
rect 311 847 315 851
rect 631 847 635 851
rect 799 847 800 851
rect 800 847 803 851
rect 823 847 827 851
rect 1115 843 1119 847
rect 1323 847 1324 851
rect 1324 847 1327 851
rect 2223 847 2227 851
rect 2231 847 2235 851
rect 2319 847 2323 851
rect 2407 847 2411 851
rect 2495 847 2499 851
rect 2823 855 2827 859
rect 2711 847 2715 851
rect 2839 847 2843 851
rect 2983 847 2987 851
rect 3191 847 3195 851
rect 3439 847 3443 851
rect 111 832 115 836
rect 135 831 139 835
rect 231 831 235 835
rect 359 831 363 835
rect 487 831 491 835
rect 623 831 627 835
rect 751 831 755 835
rect 879 831 883 835
rect 1007 831 1011 835
rect 1135 831 1139 835
rect 1271 831 1275 835
rect 1767 832 1771 836
rect 1807 832 1811 836
rect 2159 831 2163 835
rect 2247 831 2251 835
rect 2335 831 2339 835
rect 2423 831 2427 835
rect 2527 831 2531 835
rect 2639 831 2643 835
rect 2767 831 2771 835
rect 2911 831 2915 835
rect 3063 831 3067 835
rect 3223 831 3227 835
rect 3367 831 3371 835
rect 3463 832 3467 836
rect 215 823 219 827
rect 311 823 315 827
rect 823 823 827 827
rect 1115 823 1119 827
rect 111 815 115 819
rect 135 812 139 816
rect 199 815 203 819
rect 1207 819 1211 823
rect 1231 823 1235 827
rect 2231 823 2235 827
rect 2319 823 2323 827
rect 2407 823 2411 827
rect 2495 823 2499 827
rect 2519 823 2523 827
rect 2711 823 2715 827
rect 2839 823 2843 827
rect 2983 823 2987 827
rect 2991 823 2995 827
rect 3295 823 3299 827
rect 231 812 235 816
rect 359 812 363 816
rect 487 812 491 816
rect 623 812 627 816
rect 751 812 755 816
rect 879 812 883 816
rect 1007 812 1011 816
rect 1135 812 1139 816
rect 1271 812 1275 816
rect 1767 815 1771 819
rect 1807 815 1811 819
rect 3439 819 3443 823
rect 2159 812 2163 816
rect 2247 812 2251 816
rect 2335 812 2339 816
rect 2423 812 2427 816
rect 2527 812 2531 816
rect 2639 812 2643 816
rect 2767 812 2771 816
rect 2911 812 2915 816
rect 3063 812 3067 816
rect 3223 812 3227 816
rect 3367 812 3371 816
rect 3463 815 3467 819
rect 2223 771 2227 775
rect 2763 775 2767 779
rect 2991 775 2995 779
rect 111 761 115 765
rect 135 764 139 768
rect 223 764 227 768
rect 343 764 347 768
rect 471 764 475 768
rect 607 764 611 768
rect 743 764 747 768
rect 887 764 891 768
rect 1039 764 1043 768
rect 1191 764 1195 768
rect 1351 764 1355 768
rect 1767 761 1771 765
rect 1807 761 1811 765
rect 2063 764 2067 768
rect 2175 764 2179 768
rect 2295 764 2299 768
rect 2423 764 2427 768
rect 207 755 211 759
rect 295 755 299 759
rect 415 755 419 759
rect 543 755 547 759
rect 551 755 555 759
rect 807 755 811 759
rect 823 755 827 759
rect 967 755 971 759
rect 1263 755 1267 759
rect 1471 755 1475 759
rect 2135 755 2139 759
rect 2247 755 2251 759
rect 2367 755 2371 759
rect 2495 755 2499 759
rect 2559 764 2563 768
rect 2711 764 2715 768
rect 2871 764 2875 768
rect 3039 764 3043 768
rect 3215 764 3219 768
rect 3367 764 3371 768
rect 3463 761 3467 765
rect 2783 755 2787 759
rect 2943 755 2947 759
rect 3111 755 3115 759
rect 3431 755 3435 759
rect 111 744 115 748
rect 135 745 139 749
rect 223 745 227 749
rect 343 745 347 749
rect 471 745 475 749
rect 607 745 611 749
rect 743 745 747 749
rect 887 745 891 749
rect 1039 745 1043 749
rect 1191 745 1195 749
rect 1351 745 1355 749
rect 1767 744 1771 748
rect 1807 744 1811 748
rect 2063 745 2067 749
rect 2175 745 2179 749
rect 2295 745 2299 749
rect 2423 745 2427 749
rect 2559 745 2563 749
rect 2711 745 2715 749
rect 2871 745 2875 749
rect 3039 745 3043 749
rect 3215 745 3219 749
rect 3367 745 3371 749
rect 3463 744 3467 748
rect 199 727 203 731
rect 207 727 211 731
rect 295 727 299 731
rect 415 727 419 731
rect 543 727 547 731
rect 823 727 827 731
rect 967 727 971 731
rect 1103 727 1107 731
rect 1207 727 1211 731
rect 1263 727 1267 731
rect 2115 727 2116 731
rect 2116 727 2119 731
rect 2135 727 2139 731
rect 2247 727 2251 731
rect 2367 727 2371 731
rect 2495 727 2499 731
rect 2763 727 2764 731
rect 2764 727 2767 731
rect 2783 727 2787 731
rect 2943 727 2947 731
rect 3111 727 3115 731
rect 3439 727 3443 731
rect 551 719 555 723
rect 275 707 279 711
rect 367 711 371 715
rect 503 711 507 715
rect 647 711 651 715
rect 943 711 947 715
rect 951 711 955 715
rect 1263 711 1267 715
rect 1423 711 1427 715
rect 1471 711 1475 715
rect 1987 715 1991 719
rect 1999 715 2003 719
rect 2143 715 2147 719
rect 2303 715 2307 719
rect 2463 715 2467 719
rect 2795 715 2799 719
rect 3199 715 3203 719
rect 3303 715 3304 719
rect 3304 715 3307 719
rect 3431 715 3435 719
rect 111 696 115 700
rect 167 695 171 699
rect 295 695 299 699
rect 431 695 435 699
rect 575 695 579 699
rect 727 695 731 699
rect 879 695 883 699
rect 1031 695 1035 699
rect 1183 695 1187 699
rect 1343 695 1347 699
rect 1503 695 1507 699
rect 1767 696 1771 700
rect 1807 700 1811 704
rect 1927 699 1931 703
rect 2071 699 2075 703
rect 2231 699 2235 703
rect 2391 699 2395 703
rect 2551 699 2555 703
rect 2703 699 2707 703
rect 2847 699 2851 703
rect 2983 699 2987 703
rect 3119 699 3123 703
rect 3255 699 3259 703
rect 3367 699 3371 703
rect 3463 700 3467 704
rect 275 687 279 691
rect 367 687 371 691
rect 503 687 507 691
rect 647 687 651 691
rect 655 687 659 691
rect 951 687 955 691
rect 1103 687 1107 691
rect 111 679 115 683
rect 1255 683 1259 687
rect 1263 687 1267 691
rect 1423 687 1427 691
rect 1999 691 2003 695
rect 2143 691 2147 695
rect 2303 691 2307 695
rect 2463 691 2467 695
rect 2471 691 2475 695
rect 2695 691 2699 695
rect 2795 691 2799 695
rect 3191 691 3195 695
rect 3199 691 3203 695
rect 167 676 171 680
rect 295 676 299 680
rect 431 676 435 680
rect 575 676 579 680
rect 727 676 731 680
rect 879 676 883 680
rect 1031 676 1035 680
rect 1183 676 1187 680
rect 1343 676 1347 680
rect 1503 676 1507 680
rect 1767 679 1771 683
rect 1807 683 1811 687
rect 3439 687 3443 691
rect 1927 680 1931 684
rect 2071 680 2075 684
rect 2231 680 2235 684
rect 2391 680 2395 684
rect 2551 680 2555 684
rect 2703 680 2707 684
rect 2847 680 2851 684
rect 2983 680 2987 684
rect 3119 680 3123 684
rect 3255 680 3259 684
rect 3367 680 3371 684
rect 3463 683 3467 687
rect 2115 671 2119 675
rect 2471 671 2475 675
rect 1987 663 1991 667
rect 2399 663 2403 667
rect 943 635 947 639
rect 111 625 115 629
rect 455 628 459 632
rect 559 628 563 632
rect 679 628 683 632
rect 799 628 803 632
rect 927 628 931 632
rect 527 619 531 623
rect 631 619 635 623
rect 751 619 755 623
rect 871 619 875 623
rect 991 619 995 623
rect 1883 635 1887 639
rect 2239 635 2243 639
rect 2507 635 2511 639
rect 2919 635 2923 639
rect 1055 628 1059 632
rect 1183 628 1187 632
rect 1311 628 1315 632
rect 1447 628 1451 632
rect 1583 628 1587 632
rect 1767 625 1771 629
rect 1807 625 1811 629
rect 1831 628 1835 632
rect 1967 628 1971 632
rect 2135 628 2139 632
rect 2311 628 2315 632
rect 2487 628 2491 632
rect 2655 628 2659 632
rect 2815 628 2819 632
rect 2959 628 2963 632
rect 3103 628 3107 632
rect 3247 628 3251 632
rect 3367 628 3371 632
rect 3463 625 3467 629
rect 1135 619 1139 623
rect 1383 619 1387 623
rect 1519 619 1523 623
rect 1647 619 1651 623
rect 1903 619 1907 623
rect 2039 619 2043 623
rect 2207 619 2211 623
rect 2383 619 2387 623
rect 2399 619 2403 623
rect 2727 619 2731 623
rect 2887 619 2891 623
rect 3031 619 3035 623
rect 3175 619 3179 623
rect 3311 619 3315 623
rect 3431 619 3435 623
rect 111 608 115 612
rect 455 609 459 613
rect 559 609 563 613
rect 679 609 683 613
rect 799 609 803 613
rect 927 609 931 613
rect 1055 609 1059 613
rect 1183 609 1187 613
rect 1311 609 1315 613
rect 1447 609 1451 613
rect 1583 609 1587 613
rect 1767 608 1771 612
rect 1807 608 1811 612
rect 1831 609 1835 613
rect 1967 609 1971 613
rect 2135 609 2139 613
rect 2311 609 2315 613
rect 2487 609 2491 613
rect 2655 609 2659 613
rect 2815 609 2819 613
rect 2959 609 2963 613
rect 3103 609 3107 613
rect 3247 609 3251 613
rect 3367 609 3371 613
rect 3463 608 3467 612
rect 527 591 531 595
rect 631 591 635 595
rect 751 591 755 595
rect 871 591 875 595
rect 1135 591 1139 595
rect 1255 591 1259 595
rect 1383 591 1387 595
rect 1519 591 1523 595
rect 1883 591 1884 595
rect 1884 591 1887 595
rect 1903 591 1907 595
rect 2039 591 2043 595
rect 2207 591 2211 595
rect 2383 591 2387 595
rect 2695 591 2699 595
rect 2727 591 2731 595
rect 2887 591 2891 595
rect 3031 591 3035 595
rect 3319 591 3323 595
rect 3439 591 3443 595
rect 655 583 659 587
rect 1007 579 1011 583
rect 1743 579 1747 583
rect 1903 579 1907 583
rect 2039 579 2043 583
rect 2199 579 2203 583
rect 2507 579 2508 583
rect 2508 579 2511 583
rect 2527 579 2531 583
rect 2695 579 2699 583
rect 3063 579 3067 583
rect 3175 579 3179 583
rect 3431 579 3435 583
rect 671 571 675 575
rect 775 571 779 575
rect 991 571 995 575
rect 999 571 1003 575
rect 1199 571 1200 575
rect 1200 571 1203 575
rect 1223 571 1227 575
rect 1439 571 1443 575
rect 1551 571 1555 575
rect 1647 571 1651 575
rect 1735 571 1739 575
rect 1807 564 1811 568
rect 1831 563 1835 567
rect 1967 563 1971 567
rect 2127 563 2131 567
rect 2287 563 2291 567
rect 2455 563 2459 567
rect 2623 563 2627 567
rect 2799 563 2803 567
rect 2983 563 2987 567
rect 3167 563 3171 567
rect 3359 563 3363 567
rect 3463 564 3467 568
rect 111 556 115 560
rect 599 555 603 559
rect 703 555 707 559
rect 815 555 819 559
rect 927 555 931 559
rect 1039 555 1043 559
rect 1151 555 1155 559
rect 1255 555 1259 559
rect 1359 555 1363 559
rect 1471 555 1475 559
rect 1583 555 1587 559
rect 1671 555 1675 559
rect 1767 556 1771 560
rect 1903 555 1907 559
rect 2039 555 2043 559
rect 2199 555 2203 559
rect 2239 555 2243 559
rect 2527 555 2531 559
rect 2695 555 2699 559
rect 671 547 675 551
rect 775 547 779 551
rect 111 539 115 543
rect 887 543 891 547
rect 999 547 1003 551
rect 1007 547 1011 551
rect 1223 547 1227 551
rect 1439 547 1443 551
rect 1551 547 1555 551
rect 1743 547 1747 551
rect 1807 547 1811 551
rect 2879 551 2883 555
rect 2919 555 2923 559
rect 3063 555 3067 559
rect 3431 551 3435 555
rect 1831 544 1835 548
rect 599 536 603 540
rect 703 536 707 540
rect 815 536 819 540
rect 927 536 931 540
rect 1039 536 1043 540
rect 1151 536 1155 540
rect 1255 536 1259 540
rect 1359 536 1363 540
rect 1967 544 1971 548
rect 2127 544 2131 548
rect 2287 544 2291 548
rect 2455 544 2459 548
rect 2623 544 2627 548
rect 2799 544 2803 548
rect 2983 544 2987 548
rect 3167 544 3171 548
rect 3359 544 3363 548
rect 3463 547 3467 551
rect 1471 536 1475 540
rect 1583 536 1587 540
rect 1671 536 1675 540
rect 1767 539 1771 543
rect 111 489 115 493
rect 303 492 307 496
rect 431 492 435 496
rect 567 492 571 496
rect 703 492 707 496
rect 847 492 851 496
rect 983 492 987 496
rect 1111 492 1115 496
rect 1231 492 1235 496
rect 1351 492 1355 496
rect 1463 492 1467 496
rect 1575 492 1579 496
rect 1671 492 1675 496
rect 1767 489 1771 493
rect 1883 491 1887 495
rect 375 483 379 487
rect 503 483 507 487
rect 631 483 635 487
rect 647 483 651 487
rect 783 483 787 487
rect 1055 483 1059 487
rect 1199 483 1203 487
rect 1303 483 1307 487
rect 1311 483 1315 487
rect 1431 483 1435 487
rect 1735 483 1739 487
rect 1807 481 1811 485
rect 1831 484 1835 488
rect 1967 484 1971 488
rect 111 472 115 476
rect 303 473 307 477
rect 431 473 435 477
rect 567 473 571 477
rect 703 473 707 477
rect 847 473 851 477
rect 983 473 987 477
rect 1111 473 1115 477
rect 1231 473 1235 477
rect 1351 473 1355 477
rect 1463 473 1467 477
rect 1575 473 1579 477
rect 1671 473 1675 477
rect 1767 472 1771 476
rect 1775 475 1779 479
rect 2039 475 2043 479
rect 2731 491 2735 495
rect 2127 484 2131 488
rect 2295 484 2299 488
rect 2479 484 2483 488
rect 2679 484 2683 488
rect 2887 484 2891 488
rect 2359 475 2363 479
rect 2375 475 2379 479
rect 2559 475 2563 479
rect 2959 475 2963 479
rect 3111 484 3115 488
rect 3335 484 3339 488
rect 3463 481 3467 485
rect 3319 475 3323 479
rect 1807 464 1811 468
rect 1831 465 1835 469
rect 1967 465 1971 469
rect 2127 465 2131 469
rect 2295 465 2299 469
rect 2479 465 2483 469
rect 2679 465 2683 469
rect 2887 465 2891 469
rect 3111 465 3115 469
rect 3335 465 3339 469
rect 3463 464 3467 468
rect 375 455 379 459
rect 503 455 507 459
rect 647 451 651 455
rect 783 455 787 459
rect 887 455 891 459
rect 975 455 979 459
rect 1055 455 1059 459
rect 1311 455 1315 459
rect 1431 455 1435 459
rect 215 435 219 439
rect 387 435 391 439
rect 679 443 683 447
rect 1775 447 1779 451
rect 1883 447 1884 451
rect 1884 447 1887 451
rect 2031 447 2035 451
rect 2039 447 2043 451
rect 2375 447 2379 451
rect 2559 447 2563 451
rect 2731 447 2732 451
rect 2732 447 2735 451
rect 2879 447 2883 451
rect 2959 447 2963 451
rect 3431 447 3435 451
rect 631 435 632 439
rect 632 435 635 439
rect 655 435 659 439
rect 1127 435 1131 439
rect 1295 435 1299 439
rect 1303 435 1307 439
rect 1383 435 1387 439
rect 1511 435 1515 439
rect 1639 435 1643 439
rect 1743 435 1747 439
rect 1903 435 1907 439
rect 2119 435 2123 439
rect 2359 435 2363 439
rect 2403 435 2407 439
rect 2527 435 2531 439
rect 2727 435 2731 439
rect 2943 435 2947 439
rect 3343 435 3347 439
rect 111 420 115 424
rect 135 419 139 423
rect 255 419 259 423
rect 415 419 419 423
rect 583 419 587 423
rect 743 419 747 423
rect 903 419 907 423
rect 1047 419 1051 423
rect 1183 419 1187 423
rect 1311 419 1315 423
rect 1439 419 1443 423
rect 1567 419 1571 423
rect 1671 419 1675 423
rect 1767 420 1771 424
rect 1807 420 1811 424
rect 1831 419 1835 423
rect 1959 419 1963 423
rect 2111 419 2115 423
rect 2271 419 2275 423
rect 2455 419 2459 423
rect 2655 419 2659 423
rect 2871 419 2875 423
rect 3103 419 3107 423
rect 3335 419 3339 423
rect 3463 420 3467 424
rect 215 411 219 415
rect 387 411 391 415
rect 655 411 659 415
rect 679 411 683 415
rect 975 411 979 415
rect 1127 411 1131 415
rect 1383 411 1387 415
rect 1511 411 1515 415
rect 1639 411 1643 415
rect 1743 411 1747 415
rect 1903 411 1907 415
rect 2031 411 2035 415
rect 2075 411 2079 415
rect 2403 411 2407 415
rect 2527 411 2531 415
rect 2727 411 2731 415
rect 2943 411 2947 415
rect 3019 411 3023 415
rect 111 403 115 407
rect 135 400 139 404
rect 199 403 203 407
rect 255 400 259 404
rect 415 400 419 404
rect 583 400 587 404
rect 743 400 747 404
rect 903 400 907 404
rect 1047 400 1051 404
rect 1183 400 1187 404
rect 1311 400 1315 404
rect 1439 400 1443 404
rect 1567 400 1571 404
rect 1671 400 1675 404
rect 1767 403 1771 407
rect 1807 403 1811 407
rect 3407 407 3411 411
rect 1831 400 1835 404
rect 1959 400 1963 404
rect 2111 400 2115 404
rect 2271 400 2275 404
rect 2455 400 2459 404
rect 2655 400 2659 404
rect 2871 400 2875 404
rect 3103 400 3107 404
rect 3335 400 3339 404
rect 3463 403 3467 407
rect 1295 371 1299 375
rect 2075 371 2079 375
rect 2731 367 2735 371
rect 3031 367 3035 371
rect 2635 359 2639 363
rect 3019 359 3023 363
rect 111 349 115 353
rect 135 352 139 356
rect 223 352 227 356
rect 343 352 347 356
rect 471 352 475 356
rect 599 352 603 356
rect 719 352 723 356
rect 839 352 843 356
rect 959 352 963 356
rect 1079 352 1083 356
rect 1207 352 1211 356
rect 1767 349 1771 353
rect 1807 349 1811 353
rect 1927 352 1931 356
rect 2039 352 2043 356
rect 2159 352 2163 356
rect 2287 352 2291 356
rect 2423 352 2427 356
rect 2583 352 2587 356
rect 2759 352 2763 356
rect 2951 352 2955 356
rect 3151 352 3155 356
rect 3359 352 3363 356
rect 3463 349 3467 353
rect 207 343 211 347
rect 295 343 299 347
rect 415 343 419 347
rect 543 343 547 347
rect 551 343 555 347
rect 823 343 827 347
rect 911 343 915 347
rect 1031 343 1035 347
rect 1151 343 1155 347
rect 1999 343 2003 347
rect 2119 343 2123 347
rect 2127 343 2131 347
rect 2239 343 2243 347
rect 2367 343 2371 347
rect 2655 343 2659 347
rect 2831 343 2835 347
rect 3023 343 3027 347
rect 3031 343 3035 347
rect 3423 343 3427 347
rect 111 332 115 336
rect 135 333 139 337
rect 223 333 227 337
rect 343 333 347 337
rect 471 333 475 337
rect 599 333 603 337
rect 719 333 723 337
rect 839 333 843 337
rect 959 333 963 337
rect 1079 333 1083 337
rect 1207 333 1211 337
rect 1767 332 1771 336
rect 1807 332 1811 336
rect 1927 333 1931 337
rect 2039 333 2043 337
rect 2159 333 2163 337
rect 2287 333 2291 337
rect 2423 333 2427 337
rect 2583 333 2587 337
rect 2759 333 2763 337
rect 2951 333 2955 337
rect 3151 333 3155 337
rect 3359 333 3363 337
rect 3463 332 3467 336
rect 199 315 203 319
rect 207 315 211 319
rect 295 315 299 319
rect 415 315 419 319
rect 543 315 547 319
rect 823 315 827 319
rect 911 315 915 319
rect 1031 315 1035 319
rect 1151 315 1155 319
rect 551 307 555 311
rect 1999 315 2003 319
rect 2239 315 2243 319
rect 2367 315 2371 319
rect 2471 315 2472 319
rect 2472 315 2475 319
rect 2635 315 2636 319
rect 2636 315 2639 319
rect 2655 315 2659 319
rect 2831 315 2835 319
rect 3023 315 3027 319
rect 3407 315 3408 319
rect 3408 315 3411 319
rect 2127 307 2131 311
rect 335 299 339 303
rect 447 299 451 303
rect 559 299 563 303
rect 775 299 779 303
rect 983 299 987 303
rect 1199 299 1203 303
rect 2275 303 2276 307
rect 2276 303 2279 307
rect 2295 303 2299 307
rect 2383 303 2387 307
rect 2567 303 2571 307
rect 2627 303 2628 307
rect 2628 303 2631 307
rect 2731 303 2732 307
rect 2732 303 2735 307
rect 2751 303 2755 307
rect 2871 303 2875 307
rect 2999 303 3003 307
rect 3143 303 3147 307
rect 3416 303 3420 307
rect 111 284 115 288
rect 263 283 267 287
rect 375 283 379 287
rect 487 283 491 287
rect 599 283 603 287
rect 711 283 715 287
rect 815 283 819 287
rect 919 283 923 287
rect 1023 283 1027 287
rect 335 275 339 279
rect 447 275 451 279
rect 559 275 563 279
rect 587 275 591 279
rect 111 267 115 271
rect 783 271 787 275
rect 1127 283 1131 287
rect 1239 283 1243 287
rect 1767 284 1771 288
rect 1807 288 1811 292
rect 2223 287 2227 291
rect 2311 287 2315 291
rect 2399 287 2403 291
rect 2487 287 2491 291
rect 2575 287 2579 291
rect 2679 287 2683 291
rect 2799 287 2803 291
rect 2927 287 2931 291
rect 3071 287 3075 291
rect 3223 287 3227 291
rect 3367 287 3371 291
rect 3463 288 3467 292
rect 1199 275 1203 279
rect 2295 279 2299 283
rect 2383 279 2387 283
rect 2471 279 2475 283
rect 2479 279 2483 283
rect 2567 279 2571 283
rect 2751 279 2755 283
rect 2871 279 2875 283
rect 2999 279 3003 283
rect 3143 279 3147 283
rect 3151 279 3155 283
rect 1319 271 1323 275
rect 263 264 267 268
rect 375 264 379 268
rect 487 264 491 268
rect 599 264 603 268
rect 711 264 715 268
rect 815 264 819 268
rect 919 264 923 268
rect 1023 264 1027 268
rect 1127 264 1131 268
rect 1239 264 1243 268
rect 1767 267 1771 271
rect 1807 271 1811 275
rect 3439 275 3443 279
rect 2223 268 2227 272
rect 2311 268 2315 272
rect 2399 268 2403 272
rect 2487 268 2491 272
rect 2575 268 2579 272
rect 2679 268 2683 272
rect 2799 268 2803 272
rect 2927 268 2931 272
rect 3071 268 3075 272
rect 3223 268 3227 272
rect 3367 268 3371 272
rect 3463 271 3467 275
rect 2275 259 2279 263
rect 2479 259 2483 263
rect 111 213 115 217
rect 447 216 451 220
rect 535 216 539 220
rect 623 216 627 220
rect 711 216 715 220
rect 807 216 811 220
rect 903 216 907 220
rect 999 216 1003 220
rect 1103 216 1107 220
rect 1207 216 1211 220
rect 1311 216 1315 220
rect 1767 213 1771 217
rect 1807 213 1811 217
rect 2143 216 2147 220
rect 2263 216 2267 220
rect 2383 216 2387 220
rect 2511 216 2515 220
rect 2639 216 2643 220
rect 2767 216 2771 220
rect 2895 216 2899 220
rect 3015 216 3019 220
rect 3135 216 3139 220
rect 3263 216 3267 220
rect 3367 216 3371 220
rect 3463 213 3467 217
rect 315 207 319 211
rect 527 207 531 211
rect 695 207 699 211
rect 775 207 779 211
rect 879 207 883 211
rect 887 207 891 211
rect 983 207 987 211
rect 1287 207 1291 211
rect 2215 207 2219 211
rect 2335 207 2339 211
rect 2455 207 2459 211
rect 2583 207 2587 211
rect 2627 207 2631 211
rect 2975 207 2979 211
rect 3207 207 3211 211
rect 3343 207 3347 211
rect 3431 207 3435 211
rect 111 196 115 200
rect 447 197 451 201
rect 535 197 539 201
rect 623 197 627 201
rect 711 197 715 201
rect 807 197 811 201
rect 903 197 907 201
rect 999 197 1003 201
rect 1103 197 1107 201
rect 1207 197 1211 201
rect 1311 197 1315 201
rect 1767 196 1771 200
rect 1807 196 1811 200
rect 2143 197 2147 201
rect 2263 197 2267 201
rect 2383 197 2387 201
rect 2511 197 2515 201
rect 2639 197 2643 201
rect 2767 197 2771 201
rect 2895 197 2899 201
rect 3015 197 3019 201
rect 3135 197 3139 201
rect 3263 197 3267 201
rect 3367 197 3371 201
rect 3463 196 3467 200
rect 527 179 531 183
rect 587 179 588 183
rect 588 179 591 183
rect 695 179 699 183
rect 783 179 787 183
rect 887 179 891 183
rect 951 179 952 183
rect 952 179 955 183
rect 879 171 883 175
rect 1287 179 1291 183
rect 1319 179 1323 183
rect 2215 179 2219 183
rect 2335 179 2339 183
rect 2455 179 2459 183
rect 2583 179 2587 183
rect 2975 179 2979 183
rect 3151 179 3155 183
rect 3183 179 3184 183
rect 3184 179 3187 183
rect 3207 179 3211 183
rect 3439 179 3443 183
rect 2375 171 2379 175
rect 315 139 316 143
rect 316 139 319 143
rect 335 139 339 143
rect 423 139 427 143
rect 511 139 515 143
rect 599 139 603 143
rect 687 139 691 143
rect 775 139 779 143
rect 863 139 867 143
rect 1039 139 1043 143
rect 1127 139 1131 143
rect 1215 139 1219 143
rect 1303 139 1307 143
rect 1391 139 1395 143
rect 1479 139 1483 143
rect 1567 139 1571 143
rect 1655 139 1659 143
rect 1743 143 1747 147
rect 1903 143 1907 147
rect 1991 143 1995 147
rect 2079 143 2083 147
rect 2167 143 2171 147
rect 2255 143 2259 147
rect 2367 143 2371 147
rect 2583 143 2587 147
rect 2687 143 2691 147
rect 2791 143 2795 147
rect 2887 143 2891 147
rect 2983 143 2987 147
rect 3079 143 3083 147
rect 3175 143 3179 147
rect 3359 143 3363 147
rect 3431 143 3435 147
rect 111 124 115 128
rect 263 123 267 127
rect 351 123 355 127
rect 439 123 443 127
rect 527 123 531 127
rect 615 123 619 127
rect 703 123 707 127
rect 791 123 795 127
rect 879 123 883 127
rect 967 123 971 127
rect 1055 123 1059 127
rect 1143 123 1147 127
rect 1231 123 1235 127
rect 1319 123 1323 127
rect 1407 123 1411 127
rect 1495 123 1499 127
rect 1583 123 1587 127
rect 1671 123 1675 127
rect 1767 124 1771 128
rect 1807 128 1811 132
rect 1831 127 1835 131
rect 1919 127 1923 131
rect 2007 127 2011 131
rect 2095 127 2099 131
rect 2183 127 2187 131
rect 2295 127 2299 131
rect 2407 127 2411 131
rect 2511 127 2515 131
rect 2615 127 2619 131
rect 2719 127 2723 131
rect 2815 127 2819 131
rect 2911 127 2915 131
rect 3007 127 3011 131
rect 3103 127 3107 131
rect 3191 127 3195 131
rect 3279 127 3283 131
rect 3367 127 3371 131
rect 3463 128 3467 132
rect 335 115 339 119
rect 423 115 427 119
rect 511 115 515 119
rect 599 115 603 119
rect 687 115 691 119
rect 775 115 779 119
rect 863 115 867 119
rect 951 115 955 119
rect 1039 115 1043 119
rect 1127 115 1131 119
rect 1215 115 1219 119
rect 1303 115 1307 119
rect 1391 115 1395 119
rect 1479 115 1483 119
rect 1567 115 1571 119
rect 1655 115 1659 119
rect 1743 115 1747 119
rect 1903 119 1907 123
rect 1991 119 1995 123
rect 2079 119 2083 123
rect 2167 119 2171 123
rect 2255 119 2259 123
rect 2367 119 2371 123
rect 2375 119 2379 123
rect 2583 119 2587 123
rect 2687 119 2691 123
rect 2791 119 2795 123
rect 2887 119 2891 123
rect 2983 119 2987 123
rect 3079 119 3083 123
rect 3175 119 3179 123
rect 3183 119 3187 123
rect 3359 119 3363 123
rect 111 107 115 111
rect 263 104 267 108
rect 351 104 355 108
rect 439 104 443 108
rect 527 104 531 108
rect 615 104 619 108
rect 703 104 707 108
rect 791 104 795 108
rect 879 104 883 108
rect 967 104 971 108
rect 1055 104 1059 108
rect 1143 104 1147 108
rect 1231 104 1235 108
rect 1319 104 1323 108
rect 1407 104 1411 108
rect 1495 104 1499 108
rect 1583 104 1587 108
rect 1671 104 1675 108
rect 1767 107 1771 111
rect 1807 111 1811 115
rect 1831 108 1835 112
rect 1919 108 1923 112
rect 2007 108 2011 112
rect 2095 108 2099 112
rect 2183 108 2187 112
rect 2295 108 2299 112
rect 2407 108 2411 112
rect 2511 108 2515 112
rect 2615 108 2619 112
rect 2719 108 2723 112
rect 2815 108 2819 112
rect 2911 108 2915 112
rect 3007 108 3011 112
rect 3103 108 3107 112
rect 3191 108 3195 112
rect 3279 108 3283 112
rect 3367 108 3371 112
rect 3463 111 3467 115
<< m3 >>
rect 1342 3507 1348 3508
rect 111 3506 115 3507
rect 111 3501 115 3502
rect 135 3506 139 3507
rect 135 3501 139 3502
rect 271 3506 275 3507
rect 271 3501 275 3502
rect 439 3506 443 3507
rect 439 3501 443 3502
rect 615 3506 619 3507
rect 615 3501 619 3502
rect 791 3506 795 3507
rect 791 3501 795 3502
rect 959 3506 963 3507
rect 959 3501 963 3502
rect 1119 3506 1123 3507
rect 1119 3501 1123 3502
rect 1263 3506 1267 3507
rect 1342 3503 1343 3507
rect 1347 3503 1348 3507
rect 1342 3502 1348 3503
rect 1407 3506 1411 3507
rect 1263 3501 1267 3502
rect 112 3485 114 3501
rect 110 3484 116 3485
rect 136 3484 138 3501
rect 206 3499 212 3500
rect 206 3495 207 3499
rect 211 3495 212 3499
rect 206 3494 212 3495
rect 110 3480 111 3484
rect 115 3480 116 3484
rect 110 3479 116 3480
rect 134 3483 140 3484
rect 134 3479 135 3483
rect 139 3479 140 3483
rect 134 3478 140 3479
rect 208 3476 210 3494
rect 272 3484 274 3501
rect 342 3499 348 3500
rect 342 3495 343 3499
rect 347 3495 348 3499
rect 342 3494 348 3495
rect 270 3483 276 3484
rect 270 3479 271 3483
rect 275 3479 276 3483
rect 270 3478 276 3479
rect 344 3476 346 3494
rect 440 3484 442 3501
rect 510 3499 516 3500
rect 510 3495 511 3499
rect 515 3495 516 3499
rect 510 3494 516 3495
rect 438 3483 444 3484
rect 438 3479 439 3483
rect 443 3479 444 3483
rect 438 3478 444 3479
rect 512 3476 514 3494
rect 616 3484 618 3501
rect 686 3499 692 3500
rect 686 3495 687 3499
rect 691 3495 692 3499
rect 686 3494 692 3495
rect 614 3483 620 3484
rect 614 3479 615 3483
rect 619 3479 620 3483
rect 614 3478 620 3479
rect 688 3476 690 3494
rect 792 3484 794 3501
rect 960 3484 962 3501
rect 1090 3495 1096 3496
rect 1090 3491 1091 3495
rect 1095 3491 1096 3495
rect 1090 3490 1096 3491
rect 790 3483 796 3484
rect 790 3479 791 3483
rect 795 3479 796 3483
rect 790 3478 796 3479
rect 958 3483 964 3484
rect 958 3479 959 3483
rect 963 3479 964 3483
rect 958 3478 964 3479
rect 1092 3476 1094 3490
rect 1120 3484 1122 3501
rect 1190 3499 1196 3500
rect 1190 3495 1191 3499
rect 1195 3495 1196 3499
rect 1190 3494 1196 3495
rect 1118 3483 1124 3484
rect 1118 3479 1119 3483
rect 1123 3479 1124 3483
rect 1118 3478 1124 3479
rect 1192 3476 1194 3494
rect 1264 3484 1266 3501
rect 1334 3499 1340 3500
rect 1334 3495 1335 3499
rect 1339 3495 1340 3499
rect 1334 3494 1340 3495
rect 1262 3483 1268 3484
rect 1262 3479 1263 3483
rect 1267 3479 1268 3483
rect 1262 3478 1268 3479
rect 1336 3476 1338 3494
rect 206 3475 212 3476
rect 206 3471 207 3475
rect 211 3471 212 3475
rect 206 3470 212 3471
rect 342 3475 348 3476
rect 342 3471 343 3475
rect 347 3471 348 3475
rect 342 3470 348 3471
rect 510 3475 516 3476
rect 510 3471 511 3475
rect 515 3471 516 3475
rect 510 3470 516 3471
rect 686 3475 692 3476
rect 686 3471 687 3475
rect 691 3471 692 3475
rect 686 3470 692 3471
rect 782 3475 788 3476
rect 782 3471 783 3475
rect 787 3471 788 3475
rect 782 3470 788 3471
rect 1090 3475 1096 3476
rect 1090 3471 1091 3475
rect 1095 3471 1096 3475
rect 1090 3470 1096 3471
rect 1190 3475 1196 3476
rect 1190 3471 1191 3475
rect 1195 3471 1196 3475
rect 1190 3470 1196 3471
rect 1334 3475 1340 3476
rect 1334 3471 1335 3475
rect 1339 3471 1340 3475
rect 1334 3470 1340 3471
rect 110 3467 116 3468
rect 110 3463 111 3467
rect 115 3463 116 3467
rect 110 3462 116 3463
rect 134 3464 140 3465
rect 112 3439 114 3462
rect 134 3460 135 3464
rect 139 3460 140 3464
rect 134 3459 140 3460
rect 270 3464 276 3465
rect 270 3460 271 3464
rect 275 3460 276 3464
rect 270 3459 276 3460
rect 438 3464 444 3465
rect 438 3460 439 3464
rect 443 3460 444 3464
rect 438 3459 444 3460
rect 614 3464 620 3465
rect 614 3460 615 3464
rect 619 3460 620 3464
rect 614 3459 620 3460
rect 136 3439 138 3459
rect 272 3439 274 3459
rect 440 3439 442 3459
rect 616 3439 618 3459
rect 111 3438 115 3439
rect 111 3433 115 3434
rect 135 3438 139 3439
rect 135 3433 139 3434
rect 255 3438 259 3439
rect 255 3433 259 3434
rect 271 3438 275 3439
rect 271 3433 275 3434
rect 415 3438 419 3439
rect 415 3433 419 3434
rect 439 3438 443 3439
rect 439 3433 443 3434
rect 575 3438 579 3439
rect 575 3433 579 3434
rect 615 3438 619 3439
rect 615 3433 619 3434
rect 735 3438 739 3439
rect 735 3433 739 3434
rect 112 3414 114 3433
rect 136 3417 138 3433
rect 186 3423 192 3424
rect 186 3419 187 3423
rect 191 3419 192 3423
rect 186 3418 192 3419
rect 134 3416 140 3417
rect 110 3413 116 3414
rect 110 3409 111 3413
rect 115 3409 116 3413
rect 134 3412 135 3416
rect 139 3412 140 3416
rect 134 3411 140 3412
rect 110 3408 116 3409
rect 134 3397 140 3398
rect 110 3396 116 3397
rect 110 3392 111 3396
rect 115 3392 116 3396
rect 134 3393 135 3397
rect 139 3393 140 3397
rect 134 3392 140 3393
rect 110 3391 116 3392
rect 112 3367 114 3391
rect 136 3367 138 3392
rect 188 3380 190 3418
rect 256 3417 258 3433
rect 416 3417 418 3433
rect 576 3417 578 3433
rect 736 3417 738 3433
rect 254 3416 260 3417
rect 254 3412 255 3416
rect 259 3412 260 3416
rect 254 3411 260 3412
rect 414 3416 420 3417
rect 414 3412 415 3416
rect 419 3412 420 3416
rect 414 3411 420 3412
rect 574 3416 580 3417
rect 574 3412 575 3416
rect 579 3412 580 3416
rect 574 3411 580 3412
rect 734 3416 740 3417
rect 734 3412 735 3416
rect 739 3412 740 3416
rect 734 3411 740 3412
rect 206 3407 212 3408
rect 206 3403 207 3407
rect 211 3403 212 3407
rect 206 3402 212 3403
rect 326 3407 332 3408
rect 326 3403 327 3407
rect 331 3403 332 3407
rect 326 3402 332 3403
rect 486 3407 492 3408
rect 486 3403 487 3407
rect 491 3403 492 3407
rect 486 3402 492 3403
rect 654 3407 660 3408
rect 654 3403 655 3407
rect 659 3403 660 3407
rect 654 3402 660 3403
rect 208 3380 210 3402
rect 254 3397 260 3398
rect 254 3393 255 3397
rect 259 3393 260 3397
rect 254 3392 260 3393
rect 186 3379 192 3380
rect 186 3375 187 3379
rect 191 3375 192 3379
rect 186 3374 192 3375
rect 206 3379 212 3380
rect 206 3375 207 3379
rect 211 3375 212 3379
rect 206 3374 212 3375
rect 256 3367 258 3392
rect 328 3380 330 3402
rect 414 3397 420 3398
rect 414 3393 415 3397
rect 419 3393 420 3397
rect 414 3392 420 3393
rect 326 3379 332 3380
rect 326 3375 327 3379
rect 331 3375 332 3379
rect 326 3374 332 3375
rect 416 3367 418 3392
rect 111 3366 115 3367
rect 111 3361 115 3362
rect 135 3366 139 3367
rect 135 3361 139 3362
rect 255 3366 259 3367
rect 255 3361 259 3362
rect 327 3366 331 3367
rect 327 3361 331 3362
rect 415 3366 419 3367
rect 415 3361 419 3362
rect 112 3345 114 3361
rect 110 3344 116 3345
rect 136 3344 138 3361
rect 328 3344 330 3361
rect 488 3360 490 3402
rect 574 3397 580 3398
rect 574 3393 575 3397
rect 579 3393 580 3397
rect 574 3392 580 3393
rect 576 3367 578 3392
rect 656 3380 658 3402
rect 734 3397 740 3398
rect 734 3393 735 3397
rect 739 3393 740 3397
rect 734 3392 740 3393
rect 654 3379 660 3380
rect 654 3375 655 3379
rect 659 3375 660 3379
rect 654 3374 660 3375
rect 614 3367 620 3368
rect 736 3367 738 3392
rect 784 3380 786 3470
rect 790 3464 796 3465
rect 790 3460 791 3464
rect 795 3460 796 3464
rect 790 3459 796 3460
rect 958 3464 964 3465
rect 958 3460 959 3464
rect 963 3460 964 3464
rect 958 3459 964 3460
rect 1118 3464 1124 3465
rect 1118 3460 1119 3464
rect 1123 3460 1124 3464
rect 1118 3459 1124 3460
rect 1262 3464 1268 3465
rect 1262 3460 1263 3464
rect 1267 3460 1268 3464
rect 1262 3459 1268 3460
rect 792 3439 794 3459
rect 960 3439 962 3459
rect 1120 3439 1122 3459
rect 1264 3439 1266 3459
rect 791 3438 795 3439
rect 791 3433 795 3434
rect 895 3438 899 3439
rect 895 3433 899 3434
rect 959 3438 963 3439
rect 959 3433 963 3434
rect 1063 3438 1067 3439
rect 1063 3433 1067 3434
rect 1119 3438 1123 3439
rect 1119 3433 1123 3434
rect 1231 3438 1235 3439
rect 1231 3433 1235 3434
rect 1263 3438 1267 3439
rect 1263 3433 1267 3434
rect 896 3417 898 3433
rect 1064 3417 1066 3433
rect 1232 3417 1234 3433
rect 894 3416 900 3417
rect 894 3412 895 3416
rect 899 3412 900 3416
rect 894 3411 900 3412
rect 1062 3416 1068 3417
rect 1062 3412 1063 3416
rect 1067 3412 1068 3416
rect 1062 3411 1068 3412
rect 1230 3416 1236 3417
rect 1230 3412 1231 3416
rect 1235 3412 1236 3416
rect 1230 3411 1236 3412
rect 1344 3408 1346 3502
rect 1407 3501 1411 3502
rect 1551 3506 1555 3507
rect 1551 3501 1555 3502
rect 1671 3506 1675 3507
rect 1671 3501 1675 3502
rect 1767 3506 1771 3507
rect 1767 3501 1771 3502
rect 1408 3484 1410 3501
rect 1478 3499 1484 3500
rect 1478 3495 1479 3499
rect 1483 3495 1484 3499
rect 1478 3494 1484 3495
rect 1406 3483 1412 3484
rect 1406 3479 1407 3483
rect 1411 3479 1412 3483
rect 1406 3478 1412 3479
rect 1480 3476 1482 3494
rect 1552 3484 1554 3501
rect 1622 3499 1628 3500
rect 1622 3495 1623 3499
rect 1627 3495 1628 3499
rect 1622 3494 1628 3495
rect 1550 3483 1556 3484
rect 1550 3479 1551 3483
rect 1555 3479 1556 3483
rect 1550 3478 1556 3479
rect 1624 3476 1626 3494
rect 1672 3484 1674 3501
rect 1768 3485 1770 3501
rect 1807 3494 1811 3495
rect 1807 3489 1811 3490
rect 1831 3494 1835 3495
rect 1831 3489 1835 3490
rect 1975 3494 1979 3495
rect 1975 3489 1979 3490
rect 2143 3494 2147 3495
rect 2143 3489 2147 3490
rect 2311 3494 2315 3495
rect 2311 3489 2315 3490
rect 2479 3494 2483 3495
rect 2479 3489 2483 3490
rect 2639 3494 2643 3495
rect 2639 3489 2643 3490
rect 2799 3494 2803 3495
rect 2799 3489 2803 3490
rect 2967 3494 2971 3495
rect 2967 3489 2971 3490
rect 3463 3494 3467 3495
rect 3463 3489 3467 3490
rect 1766 3484 1772 3485
rect 1670 3483 1676 3484
rect 1670 3479 1671 3483
rect 1675 3479 1676 3483
rect 1766 3480 1767 3484
rect 1771 3480 1772 3484
rect 1766 3479 1772 3480
rect 1670 3478 1676 3479
rect 1478 3475 1484 3476
rect 1478 3471 1479 3475
rect 1483 3471 1484 3475
rect 1478 3470 1484 3471
rect 1622 3475 1628 3476
rect 1622 3471 1623 3475
rect 1627 3471 1628 3475
rect 1808 3473 1810 3489
rect 1622 3470 1628 3471
rect 1806 3472 1812 3473
rect 1832 3472 1834 3489
rect 1902 3487 1908 3488
rect 1902 3483 1903 3487
rect 1907 3483 1908 3487
rect 1902 3482 1908 3483
rect 1806 3468 1807 3472
rect 1811 3468 1812 3472
rect 1766 3467 1772 3468
rect 1806 3467 1812 3468
rect 1830 3471 1836 3472
rect 1830 3467 1831 3471
rect 1835 3467 1836 3471
rect 1406 3464 1412 3465
rect 1406 3460 1407 3464
rect 1411 3460 1412 3464
rect 1406 3459 1412 3460
rect 1550 3464 1556 3465
rect 1550 3460 1551 3464
rect 1555 3460 1556 3464
rect 1550 3459 1556 3460
rect 1670 3464 1676 3465
rect 1670 3460 1671 3464
rect 1675 3460 1676 3464
rect 1766 3463 1767 3467
rect 1771 3463 1772 3467
rect 1830 3466 1836 3467
rect 1904 3464 1906 3482
rect 1976 3472 1978 3489
rect 2046 3487 2052 3488
rect 2046 3483 2047 3487
rect 2051 3483 2052 3487
rect 2046 3482 2052 3483
rect 1974 3471 1980 3472
rect 1974 3467 1975 3471
rect 1979 3467 1980 3471
rect 1974 3466 1980 3467
rect 2048 3464 2050 3482
rect 2144 3472 2146 3489
rect 2214 3487 2220 3488
rect 2214 3483 2215 3487
rect 2219 3483 2220 3487
rect 2214 3482 2220 3483
rect 2142 3471 2148 3472
rect 2142 3467 2143 3471
rect 2147 3467 2148 3471
rect 2142 3466 2148 3467
rect 2216 3464 2218 3482
rect 2312 3472 2314 3489
rect 2480 3472 2482 3489
rect 2574 3487 2580 3488
rect 2574 3483 2575 3487
rect 2579 3483 2580 3487
rect 2574 3482 2580 3483
rect 2586 3487 2592 3488
rect 2586 3483 2587 3487
rect 2591 3483 2592 3487
rect 2586 3482 2592 3483
rect 2310 3471 2316 3472
rect 2310 3467 2311 3471
rect 2315 3467 2316 3471
rect 2310 3466 2316 3467
rect 2478 3471 2484 3472
rect 2478 3467 2479 3471
rect 2483 3467 2484 3471
rect 2478 3466 2484 3467
rect 1766 3462 1772 3463
rect 1902 3463 1908 3464
rect 1670 3459 1676 3460
rect 1408 3439 1410 3459
rect 1552 3439 1554 3459
rect 1672 3439 1674 3459
rect 1768 3439 1770 3462
rect 1902 3459 1903 3463
rect 1907 3459 1908 3463
rect 1902 3458 1908 3459
rect 2046 3463 2052 3464
rect 2046 3459 2047 3463
rect 2051 3459 2052 3463
rect 2046 3458 2052 3459
rect 2214 3463 2220 3464
rect 2214 3459 2215 3463
rect 2219 3459 2220 3463
rect 2214 3458 2220 3459
rect 2222 3463 2228 3464
rect 2222 3459 2223 3463
rect 2227 3459 2228 3463
rect 2222 3458 2228 3459
rect 1806 3455 1812 3456
rect 1806 3451 1807 3455
rect 1811 3451 1812 3455
rect 1806 3450 1812 3451
rect 1830 3452 1836 3453
rect 1399 3438 1403 3439
rect 1399 3433 1403 3434
rect 1407 3438 1411 3439
rect 1407 3433 1411 3434
rect 1551 3438 1555 3439
rect 1551 3433 1555 3434
rect 1671 3438 1675 3439
rect 1671 3433 1675 3434
rect 1767 3438 1771 3439
rect 1767 3433 1771 3434
rect 1400 3417 1402 3433
rect 1398 3416 1404 3417
rect 1398 3412 1399 3416
rect 1403 3412 1404 3416
rect 1768 3414 1770 3433
rect 1808 3431 1810 3450
rect 1830 3448 1831 3452
rect 1835 3448 1836 3452
rect 1830 3447 1836 3448
rect 1974 3452 1980 3453
rect 1974 3448 1975 3452
rect 1979 3448 1980 3452
rect 1974 3447 1980 3448
rect 2142 3452 2148 3453
rect 2142 3448 2143 3452
rect 2147 3448 2148 3452
rect 2142 3447 2148 3448
rect 1832 3431 1834 3447
rect 1976 3431 1978 3447
rect 2144 3431 2146 3447
rect 1807 3430 1811 3431
rect 1807 3425 1811 3426
rect 1831 3430 1835 3431
rect 1831 3425 1835 3426
rect 1975 3430 1979 3431
rect 1975 3425 1979 3426
rect 2031 3430 2035 3431
rect 2031 3425 2035 3426
rect 2143 3430 2147 3431
rect 2143 3425 2147 3426
rect 2151 3430 2155 3431
rect 2151 3425 2155 3426
rect 1398 3411 1404 3412
rect 1766 3413 1772 3414
rect 1766 3409 1767 3413
rect 1771 3409 1772 3413
rect 1766 3408 1772 3409
rect 1022 3407 1028 3408
rect 1022 3403 1023 3407
rect 1027 3403 1028 3407
rect 1022 3402 1028 3403
rect 1134 3407 1140 3408
rect 1134 3403 1135 3407
rect 1139 3403 1140 3407
rect 1134 3402 1140 3403
rect 1302 3407 1308 3408
rect 1302 3403 1303 3407
rect 1307 3403 1308 3407
rect 1302 3402 1308 3403
rect 1342 3407 1348 3408
rect 1342 3403 1343 3407
rect 1347 3403 1348 3407
rect 1808 3406 1810 3425
rect 2032 3409 2034 3425
rect 2082 3419 2088 3420
rect 2082 3415 2083 3419
rect 2087 3415 2088 3419
rect 2082 3414 2088 3415
rect 2030 3408 2036 3409
rect 1342 3402 1348 3403
rect 1806 3405 1812 3406
rect 894 3397 900 3398
rect 894 3393 895 3397
rect 899 3393 900 3397
rect 894 3392 900 3393
rect 782 3379 788 3380
rect 782 3375 783 3379
rect 787 3375 788 3379
rect 782 3374 788 3375
rect 896 3367 898 3392
rect 1024 3380 1026 3402
rect 1062 3397 1068 3398
rect 1062 3393 1063 3397
rect 1067 3393 1068 3397
rect 1062 3392 1068 3393
rect 1006 3379 1012 3380
rect 1006 3375 1007 3379
rect 1011 3375 1012 3379
rect 1006 3374 1012 3375
rect 1022 3379 1028 3380
rect 1022 3375 1023 3379
rect 1027 3375 1028 3379
rect 1022 3374 1028 3375
rect 535 3366 539 3367
rect 535 3361 539 3362
rect 575 3366 579 3367
rect 614 3363 615 3367
rect 619 3363 620 3367
rect 614 3362 620 3363
rect 735 3366 739 3367
rect 575 3361 579 3362
rect 486 3359 492 3360
rect 486 3355 487 3359
rect 491 3355 492 3359
rect 486 3354 492 3355
rect 536 3344 538 3361
rect 606 3359 612 3360
rect 606 3355 607 3359
rect 611 3355 612 3359
rect 606 3354 612 3355
rect 110 3340 111 3344
rect 115 3340 116 3344
rect 110 3339 116 3340
rect 134 3343 140 3344
rect 134 3339 135 3343
rect 139 3339 140 3343
rect 134 3338 140 3339
rect 326 3343 332 3344
rect 326 3339 327 3343
rect 331 3339 332 3343
rect 326 3338 332 3339
rect 534 3343 540 3344
rect 534 3339 535 3343
rect 539 3339 540 3343
rect 534 3338 540 3339
rect 608 3336 610 3354
rect 616 3336 618 3362
rect 735 3361 739 3362
rect 743 3366 747 3367
rect 743 3361 747 3362
rect 895 3366 899 3367
rect 895 3361 899 3362
rect 935 3366 939 3367
rect 935 3361 939 3362
rect 744 3344 746 3361
rect 936 3344 938 3361
rect 742 3343 748 3344
rect 742 3339 743 3343
rect 747 3339 748 3343
rect 742 3338 748 3339
rect 934 3343 940 3344
rect 934 3339 935 3343
rect 939 3339 940 3343
rect 934 3338 940 3339
rect 1008 3336 1010 3374
rect 1064 3367 1066 3392
rect 1136 3380 1138 3402
rect 1230 3397 1236 3398
rect 1230 3393 1231 3397
rect 1235 3393 1236 3397
rect 1230 3392 1236 3393
rect 1134 3379 1140 3380
rect 1134 3375 1135 3379
rect 1139 3375 1140 3379
rect 1134 3374 1140 3375
rect 1232 3367 1234 3392
rect 1304 3380 1306 3402
rect 1806 3401 1807 3405
rect 1811 3401 1812 3405
rect 2030 3404 2031 3408
rect 2035 3404 2036 3408
rect 2030 3403 2036 3404
rect 1806 3400 1812 3401
rect 1398 3397 1404 3398
rect 1398 3393 1399 3397
rect 1403 3393 1404 3397
rect 1398 3392 1404 3393
rect 1766 3396 1772 3397
rect 1766 3392 1767 3396
rect 1771 3392 1772 3396
rect 1302 3379 1308 3380
rect 1302 3375 1303 3379
rect 1307 3375 1308 3379
rect 1302 3374 1308 3375
rect 1400 3367 1402 3392
rect 1766 3391 1772 3392
rect 1768 3367 1770 3391
rect 2030 3389 2036 3390
rect 1806 3388 1812 3389
rect 1806 3384 1807 3388
rect 1811 3384 1812 3388
rect 2030 3385 2031 3389
rect 2035 3385 2036 3389
rect 2030 3384 2036 3385
rect 1806 3383 1812 3384
rect 1063 3366 1067 3367
rect 1063 3361 1067 3362
rect 1119 3366 1123 3367
rect 1119 3361 1123 3362
rect 1231 3366 1235 3367
rect 1231 3361 1235 3362
rect 1295 3366 1299 3367
rect 1295 3361 1299 3362
rect 1399 3366 1403 3367
rect 1399 3361 1403 3362
rect 1463 3366 1467 3367
rect 1463 3361 1467 3362
rect 1639 3366 1643 3367
rect 1639 3361 1643 3362
rect 1767 3366 1771 3367
rect 1808 3363 1810 3383
rect 2032 3363 2034 3384
rect 2084 3372 2086 3414
rect 2152 3409 2154 3425
rect 2224 3420 2226 3458
rect 2310 3452 2316 3453
rect 2310 3448 2311 3452
rect 2315 3448 2316 3452
rect 2310 3447 2316 3448
rect 2478 3452 2484 3453
rect 2478 3448 2479 3452
rect 2483 3448 2484 3452
rect 2478 3447 2484 3448
rect 2312 3431 2314 3447
rect 2480 3431 2482 3447
rect 2271 3430 2275 3431
rect 2271 3425 2275 3426
rect 2311 3430 2315 3431
rect 2311 3425 2315 3426
rect 2391 3430 2395 3431
rect 2391 3425 2395 3426
rect 2479 3430 2483 3431
rect 2479 3425 2483 3426
rect 2511 3430 2515 3431
rect 2511 3425 2515 3426
rect 2222 3419 2228 3420
rect 2222 3415 2223 3419
rect 2227 3415 2228 3419
rect 2222 3414 2228 3415
rect 2272 3409 2274 3425
rect 2392 3409 2394 3425
rect 2512 3409 2514 3425
rect 2150 3408 2156 3409
rect 2150 3404 2151 3408
rect 2155 3404 2156 3408
rect 2150 3403 2156 3404
rect 2270 3408 2276 3409
rect 2270 3404 2271 3408
rect 2275 3404 2276 3408
rect 2270 3403 2276 3404
rect 2390 3408 2396 3409
rect 2390 3404 2391 3408
rect 2395 3404 2396 3408
rect 2390 3403 2396 3404
rect 2510 3408 2516 3409
rect 2510 3404 2511 3408
rect 2515 3404 2516 3408
rect 2510 3403 2516 3404
rect 2576 3400 2578 3482
rect 2588 3464 2590 3482
rect 2640 3472 2642 3489
rect 2710 3487 2716 3488
rect 2710 3483 2711 3487
rect 2715 3483 2716 3487
rect 2710 3482 2716 3483
rect 2638 3471 2644 3472
rect 2638 3467 2639 3471
rect 2643 3467 2644 3471
rect 2638 3466 2644 3467
rect 2712 3464 2714 3482
rect 2800 3472 2802 3489
rect 2870 3487 2876 3488
rect 2870 3483 2871 3487
rect 2875 3483 2876 3487
rect 2870 3482 2876 3483
rect 2798 3471 2804 3472
rect 2798 3467 2799 3471
rect 2803 3467 2804 3471
rect 2798 3466 2804 3467
rect 2872 3464 2874 3482
rect 2968 3472 2970 3489
rect 3464 3473 3466 3489
rect 3462 3472 3468 3473
rect 2966 3471 2972 3472
rect 2966 3467 2967 3471
rect 2971 3467 2972 3471
rect 3462 3468 3463 3472
rect 3467 3468 3468 3472
rect 3462 3467 3468 3468
rect 2966 3466 2972 3467
rect 2586 3463 2592 3464
rect 2586 3459 2587 3463
rect 2591 3459 2592 3463
rect 2586 3458 2592 3459
rect 2710 3463 2716 3464
rect 2710 3459 2711 3463
rect 2715 3459 2716 3463
rect 2710 3458 2716 3459
rect 2870 3463 2876 3464
rect 2870 3459 2871 3463
rect 2875 3459 2876 3463
rect 2870 3458 2876 3459
rect 2882 3463 2888 3464
rect 2882 3459 2883 3463
rect 2887 3459 2888 3463
rect 2882 3458 2888 3459
rect 2638 3452 2644 3453
rect 2638 3448 2639 3452
rect 2643 3448 2644 3452
rect 2638 3447 2644 3448
rect 2798 3452 2804 3453
rect 2798 3448 2799 3452
rect 2803 3448 2804 3452
rect 2798 3447 2804 3448
rect 2640 3431 2642 3447
rect 2800 3431 2802 3447
rect 2623 3430 2627 3431
rect 2623 3425 2627 3426
rect 2639 3430 2643 3431
rect 2639 3425 2643 3426
rect 2727 3430 2731 3431
rect 2727 3425 2731 3426
rect 2799 3430 2803 3431
rect 2799 3425 2803 3426
rect 2831 3430 2835 3431
rect 2831 3425 2835 3426
rect 2624 3409 2626 3425
rect 2728 3409 2730 3425
rect 2832 3409 2834 3425
rect 2622 3408 2628 3409
rect 2622 3404 2623 3408
rect 2627 3404 2628 3408
rect 2622 3403 2628 3404
rect 2726 3408 2732 3409
rect 2726 3404 2727 3408
rect 2731 3404 2732 3408
rect 2726 3403 2732 3404
rect 2830 3408 2836 3409
rect 2830 3404 2831 3408
rect 2835 3404 2836 3408
rect 2830 3403 2836 3404
rect 2102 3399 2108 3400
rect 2102 3395 2103 3399
rect 2107 3395 2108 3399
rect 2102 3394 2108 3395
rect 2222 3399 2228 3400
rect 2222 3395 2223 3399
rect 2227 3395 2228 3399
rect 2222 3394 2228 3395
rect 2342 3399 2348 3400
rect 2342 3395 2343 3399
rect 2347 3395 2348 3399
rect 2342 3394 2348 3395
rect 2350 3399 2356 3400
rect 2350 3395 2351 3399
rect 2355 3395 2356 3399
rect 2350 3394 2356 3395
rect 2574 3399 2580 3400
rect 2574 3395 2575 3399
rect 2579 3395 2580 3399
rect 2574 3394 2580 3395
rect 2590 3399 2596 3400
rect 2590 3395 2591 3399
rect 2595 3395 2596 3399
rect 2590 3394 2596 3395
rect 2702 3399 2708 3400
rect 2702 3395 2703 3399
rect 2707 3395 2708 3399
rect 2702 3394 2708 3395
rect 2104 3372 2106 3394
rect 2150 3389 2156 3390
rect 2150 3385 2151 3389
rect 2155 3385 2156 3389
rect 2150 3384 2156 3385
rect 2082 3371 2088 3372
rect 2082 3367 2083 3371
rect 2087 3367 2088 3371
rect 2082 3366 2088 3367
rect 2102 3371 2108 3372
rect 2102 3367 2103 3371
rect 2107 3367 2108 3371
rect 2102 3366 2108 3367
rect 2152 3363 2154 3384
rect 2224 3372 2226 3394
rect 2270 3389 2276 3390
rect 2270 3385 2271 3389
rect 2275 3385 2276 3389
rect 2270 3384 2276 3385
rect 2222 3371 2228 3372
rect 2222 3367 2223 3371
rect 2227 3367 2228 3371
rect 2222 3366 2228 3367
rect 2272 3363 2274 3384
rect 2344 3372 2346 3394
rect 2342 3371 2348 3372
rect 2342 3367 2343 3371
rect 2347 3367 2348 3371
rect 2342 3366 2348 3367
rect 2352 3364 2354 3394
rect 2390 3389 2396 3390
rect 2390 3385 2391 3389
rect 2395 3385 2396 3389
rect 2390 3384 2396 3385
rect 2510 3389 2516 3390
rect 2510 3385 2511 3389
rect 2515 3385 2516 3389
rect 2510 3384 2516 3385
rect 2350 3363 2356 3364
rect 2392 3363 2394 3384
rect 2512 3363 2514 3384
rect 2592 3372 2594 3394
rect 2622 3389 2628 3390
rect 2622 3385 2623 3389
rect 2627 3385 2628 3389
rect 2622 3384 2628 3385
rect 2590 3371 2596 3372
rect 2590 3367 2591 3371
rect 2595 3367 2596 3371
rect 2590 3366 2596 3367
rect 2624 3363 2626 3384
rect 2704 3372 2706 3394
rect 2726 3389 2732 3390
rect 2726 3385 2727 3389
rect 2731 3385 2732 3389
rect 2726 3384 2732 3385
rect 2830 3389 2836 3390
rect 2830 3385 2831 3389
rect 2835 3385 2836 3389
rect 2830 3384 2836 3385
rect 2702 3371 2708 3372
rect 2702 3367 2703 3371
rect 2707 3367 2708 3371
rect 2702 3366 2708 3367
rect 2728 3363 2730 3384
rect 2774 3371 2780 3372
rect 2774 3367 2775 3371
rect 2779 3367 2780 3371
rect 2774 3366 2780 3367
rect 1767 3361 1771 3362
rect 1807 3362 1811 3363
rect 1070 3359 1076 3360
rect 1070 3355 1071 3359
rect 1075 3355 1076 3359
rect 1070 3354 1076 3355
rect 1072 3336 1074 3354
rect 1120 3344 1122 3361
rect 1198 3359 1204 3360
rect 1198 3355 1199 3359
rect 1203 3355 1204 3359
rect 1198 3354 1204 3355
rect 1118 3343 1124 3344
rect 1118 3339 1119 3343
rect 1123 3339 1124 3343
rect 1118 3338 1124 3339
rect 1200 3336 1202 3354
rect 1296 3344 1298 3361
rect 1374 3359 1380 3360
rect 1374 3355 1375 3359
rect 1379 3355 1380 3359
rect 1374 3354 1380 3355
rect 1294 3343 1300 3344
rect 1294 3339 1295 3343
rect 1299 3339 1300 3343
rect 1294 3338 1300 3339
rect 1376 3336 1378 3354
rect 1464 3344 1466 3361
rect 1598 3359 1604 3360
rect 1598 3355 1599 3359
rect 1603 3355 1604 3359
rect 1598 3354 1604 3355
rect 1462 3343 1468 3344
rect 1462 3339 1463 3343
rect 1467 3339 1468 3343
rect 1462 3338 1468 3339
rect 1600 3336 1602 3354
rect 1640 3344 1642 3361
rect 1734 3359 1740 3360
rect 1734 3355 1735 3359
rect 1739 3355 1740 3359
rect 1734 3354 1740 3355
rect 1638 3343 1644 3344
rect 1638 3339 1639 3343
rect 1643 3339 1644 3343
rect 1638 3338 1644 3339
rect 606 3335 612 3336
rect 606 3331 607 3335
rect 611 3331 612 3335
rect 606 3330 612 3331
rect 614 3335 620 3336
rect 614 3331 615 3335
rect 619 3331 620 3335
rect 614 3330 620 3331
rect 1006 3335 1012 3336
rect 1006 3331 1007 3335
rect 1011 3331 1012 3335
rect 1006 3330 1012 3331
rect 1070 3335 1076 3336
rect 1070 3331 1071 3335
rect 1075 3331 1076 3335
rect 1070 3330 1076 3331
rect 1198 3335 1204 3336
rect 1198 3331 1199 3335
rect 1203 3331 1204 3335
rect 1198 3330 1204 3331
rect 1374 3335 1380 3336
rect 1374 3331 1375 3335
rect 1379 3331 1380 3335
rect 1374 3330 1380 3331
rect 1598 3335 1604 3336
rect 1598 3331 1599 3335
rect 1603 3331 1604 3335
rect 1598 3330 1604 3331
rect 110 3327 116 3328
rect 110 3323 111 3327
rect 115 3323 116 3327
rect 198 3327 204 3328
rect 110 3322 116 3323
rect 134 3324 140 3325
rect 112 3295 114 3322
rect 134 3320 135 3324
rect 139 3320 140 3324
rect 198 3323 199 3327
rect 203 3323 204 3327
rect 198 3322 204 3323
rect 326 3324 332 3325
rect 134 3319 140 3320
rect 136 3295 138 3319
rect 111 3294 115 3295
rect 111 3289 115 3290
rect 135 3294 139 3295
rect 135 3289 139 3290
rect 112 3270 114 3289
rect 136 3273 138 3289
rect 134 3272 140 3273
rect 110 3269 116 3270
rect 110 3265 111 3269
rect 115 3265 116 3269
rect 134 3268 135 3272
rect 139 3268 140 3272
rect 134 3267 140 3268
rect 110 3264 116 3265
rect 134 3253 140 3254
rect 110 3252 116 3253
rect 110 3248 111 3252
rect 115 3248 116 3252
rect 134 3249 135 3253
rect 139 3249 140 3253
rect 134 3248 140 3249
rect 110 3247 116 3248
rect 112 3223 114 3247
rect 136 3223 138 3248
rect 200 3236 202 3322
rect 326 3320 327 3324
rect 331 3320 332 3324
rect 326 3319 332 3320
rect 534 3324 540 3325
rect 534 3320 535 3324
rect 539 3320 540 3324
rect 534 3319 540 3320
rect 742 3324 748 3325
rect 742 3320 743 3324
rect 747 3320 748 3324
rect 742 3319 748 3320
rect 934 3324 940 3325
rect 934 3320 935 3324
rect 939 3320 940 3324
rect 934 3319 940 3320
rect 1118 3324 1124 3325
rect 1118 3320 1119 3324
rect 1123 3320 1124 3324
rect 1118 3319 1124 3320
rect 1294 3324 1300 3325
rect 1294 3320 1295 3324
rect 1299 3320 1300 3324
rect 1294 3319 1300 3320
rect 1462 3324 1468 3325
rect 1462 3320 1463 3324
rect 1467 3320 1468 3324
rect 1462 3319 1468 3320
rect 1638 3324 1644 3325
rect 1638 3320 1639 3324
rect 1643 3320 1644 3324
rect 1638 3319 1644 3320
rect 328 3295 330 3319
rect 536 3295 538 3319
rect 744 3295 746 3319
rect 936 3295 938 3319
rect 1120 3295 1122 3319
rect 1296 3295 1298 3319
rect 1464 3295 1466 3319
rect 1640 3295 1642 3319
rect 279 3294 283 3295
rect 279 3289 283 3290
rect 327 3294 331 3295
rect 327 3289 331 3290
rect 463 3294 467 3295
rect 463 3289 467 3290
rect 535 3294 539 3295
rect 535 3289 539 3290
rect 647 3294 651 3295
rect 647 3289 651 3290
rect 743 3294 747 3295
rect 743 3289 747 3290
rect 831 3294 835 3295
rect 831 3289 835 3290
rect 935 3294 939 3295
rect 935 3289 939 3290
rect 1007 3294 1011 3295
rect 1007 3289 1011 3290
rect 1119 3294 1123 3295
rect 1119 3289 1123 3290
rect 1175 3294 1179 3295
rect 1175 3289 1179 3290
rect 1295 3294 1299 3295
rect 1295 3289 1299 3290
rect 1343 3294 1347 3295
rect 1343 3289 1347 3290
rect 1463 3294 1467 3295
rect 1463 3289 1467 3290
rect 1503 3294 1507 3295
rect 1503 3289 1507 3290
rect 1639 3294 1643 3295
rect 1639 3289 1643 3290
rect 1671 3294 1675 3295
rect 1671 3289 1675 3290
rect 234 3279 240 3280
rect 234 3275 235 3279
rect 239 3275 240 3279
rect 234 3274 240 3275
rect 206 3263 212 3264
rect 206 3259 207 3263
rect 211 3259 212 3263
rect 206 3258 212 3259
rect 208 3236 210 3258
rect 198 3235 204 3236
rect 198 3231 199 3235
rect 203 3231 204 3235
rect 198 3230 204 3231
rect 206 3235 212 3236
rect 206 3231 207 3235
rect 211 3231 212 3235
rect 206 3230 212 3231
rect 111 3222 115 3223
rect 111 3217 115 3218
rect 135 3222 139 3223
rect 135 3217 139 3218
rect 183 3222 187 3223
rect 183 3217 187 3218
rect 112 3201 114 3217
rect 110 3200 116 3201
rect 184 3200 186 3217
rect 236 3216 238 3274
rect 280 3273 282 3289
rect 464 3273 466 3289
rect 648 3273 650 3289
rect 832 3273 834 3289
rect 1008 3273 1010 3289
rect 1176 3273 1178 3289
rect 1344 3273 1346 3289
rect 1504 3273 1506 3289
rect 1672 3273 1674 3289
rect 278 3272 284 3273
rect 278 3268 279 3272
rect 283 3268 284 3272
rect 278 3267 284 3268
rect 462 3272 468 3273
rect 462 3268 463 3272
rect 467 3268 468 3272
rect 462 3267 468 3268
rect 646 3272 652 3273
rect 646 3268 647 3272
rect 651 3268 652 3272
rect 646 3267 652 3268
rect 830 3272 836 3273
rect 830 3268 831 3272
rect 835 3268 836 3272
rect 830 3267 836 3268
rect 1006 3272 1012 3273
rect 1006 3268 1007 3272
rect 1011 3268 1012 3272
rect 1006 3267 1012 3268
rect 1174 3272 1180 3273
rect 1174 3268 1175 3272
rect 1179 3268 1180 3272
rect 1174 3267 1180 3268
rect 1342 3272 1348 3273
rect 1342 3268 1343 3272
rect 1347 3268 1348 3272
rect 1342 3267 1348 3268
rect 1502 3272 1508 3273
rect 1502 3268 1503 3272
rect 1507 3268 1508 3272
rect 1502 3267 1508 3268
rect 1670 3272 1676 3273
rect 1670 3268 1671 3272
rect 1675 3268 1676 3272
rect 1670 3267 1676 3268
rect 1736 3264 1738 3354
rect 1768 3345 1770 3361
rect 1807 3357 1811 3358
rect 2031 3362 2035 3363
rect 2031 3357 2035 3358
rect 2151 3362 2155 3363
rect 2151 3357 2155 3358
rect 2159 3362 2163 3363
rect 2159 3357 2163 3358
rect 2271 3362 2275 3363
rect 2271 3357 2275 3358
rect 2295 3362 2299 3363
rect 2350 3359 2351 3363
rect 2355 3359 2356 3363
rect 2350 3358 2356 3359
rect 2391 3362 2395 3363
rect 2295 3357 2299 3358
rect 2391 3357 2395 3358
rect 2431 3362 2435 3363
rect 2431 3357 2435 3358
rect 2511 3362 2515 3363
rect 2511 3357 2515 3358
rect 2567 3362 2571 3363
rect 2567 3357 2571 3358
rect 2623 3362 2627 3363
rect 2623 3357 2627 3358
rect 2703 3362 2707 3363
rect 2703 3357 2707 3358
rect 2727 3362 2731 3363
rect 2727 3357 2731 3358
rect 1766 3344 1772 3345
rect 1766 3340 1767 3344
rect 1771 3340 1772 3344
rect 1808 3341 1810 3357
rect 1766 3339 1772 3340
rect 1806 3340 1812 3341
rect 2160 3340 2162 3357
rect 2230 3355 2236 3356
rect 2230 3351 2231 3355
rect 2235 3351 2236 3355
rect 2230 3350 2236 3351
rect 1806 3336 1807 3340
rect 1811 3336 1812 3340
rect 1806 3335 1812 3336
rect 2158 3339 2164 3340
rect 2158 3335 2159 3339
rect 2163 3335 2164 3339
rect 2158 3334 2164 3335
rect 2232 3332 2234 3350
rect 2296 3340 2298 3357
rect 2366 3355 2372 3356
rect 2366 3351 2367 3355
rect 2371 3351 2372 3355
rect 2366 3350 2372 3351
rect 2294 3339 2300 3340
rect 2294 3335 2295 3339
rect 2299 3335 2300 3339
rect 2294 3334 2300 3335
rect 2368 3332 2370 3350
rect 2432 3340 2434 3357
rect 2502 3355 2508 3356
rect 2502 3351 2503 3355
rect 2507 3351 2508 3355
rect 2502 3350 2508 3351
rect 2430 3339 2436 3340
rect 2430 3335 2431 3339
rect 2435 3335 2436 3339
rect 2430 3334 2436 3335
rect 2504 3332 2506 3350
rect 2568 3340 2570 3357
rect 2704 3340 2706 3357
rect 2566 3339 2572 3340
rect 2566 3335 2567 3339
rect 2571 3335 2572 3339
rect 2566 3334 2572 3335
rect 2702 3339 2708 3340
rect 2702 3335 2703 3339
rect 2707 3335 2708 3339
rect 2702 3334 2708 3335
rect 2776 3332 2778 3366
rect 2832 3363 2834 3384
rect 2884 3372 2886 3458
rect 3462 3455 3468 3456
rect 2966 3452 2972 3453
rect 2966 3448 2967 3452
rect 2971 3448 2972 3452
rect 3462 3451 3463 3455
rect 3467 3451 3468 3455
rect 3462 3450 3468 3451
rect 2966 3447 2972 3448
rect 2968 3431 2970 3447
rect 3464 3431 3466 3450
rect 2935 3430 2939 3431
rect 2935 3425 2939 3426
rect 2967 3430 2971 3431
rect 2967 3425 2971 3426
rect 3039 3430 3043 3431
rect 3039 3425 3043 3426
rect 3151 3430 3155 3431
rect 3151 3425 3155 3426
rect 3463 3430 3467 3431
rect 3463 3425 3467 3426
rect 2936 3409 2938 3425
rect 3040 3409 3042 3425
rect 3152 3409 3154 3425
rect 2934 3408 2940 3409
rect 2934 3404 2935 3408
rect 2939 3404 2940 3408
rect 2934 3403 2940 3404
rect 3038 3408 3044 3409
rect 3038 3404 3039 3408
rect 3043 3404 3044 3408
rect 3038 3403 3044 3404
rect 3150 3408 3156 3409
rect 3150 3404 3151 3408
rect 3155 3404 3156 3408
rect 3464 3406 3466 3425
rect 3150 3403 3156 3404
rect 3462 3405 3468 3406
rect 3462 3401 3463 3405
rect 3467 3401 3468 3405
rect 3462 3400 3468 3401
rect 2902 3399 2908 3400
rect 2902 3395 2903 3399
rect 2907 3395 2908 3399
rect 2902 3394 2908 3395
rect 3006 3399 3012 3400
rect 3006 3395 3007 3399
rect 3011 3395 3012 3399
rect 3006 3394 3012 3395
rect 3110 3399 3116 3400
rect 3110 3395 3111 3399
rect 3115 3395 3116 3399
rect 3110 3394 3116 3395
rect 3214 3399 3220 3400
rect 3214 3395 3215 3399
rect 3219 3395 3220 3399
rect 3214 3394 3220 3395
rect 2904 3372 2906 3394
rect 2934 3389 2940 3390
rect 2934 3385 2935 3389
rect 2939 3385 2940 3389
rect 2934 3384 2940 3385
rect 2882 3371 2888 3372
rect 2882 3367 2883 3371
rect 2887 3367 2888 3371
rect 2882 3366 2888 3367
rect 2902 3371 2908 3372
rect 2902 3367 2903 3371
rect 2907 3367 2908 3371
rect 2902 3366 2908 3367
rect 2936 3363 2938 3384
rect 3008 3372 3010 3394
rect 3038 3389 3044 3390
rect 3038 3385 3039 3389
rect 3043 3385 3044 3389
rect 3038 3384 3044 3385
rect 3006 3371 3012 3372
rect 3006 3367 3007 3371
rect 3011 3367 3012 3371
rect 3006 3366 3012 3367
rect 3040 3363 3042 3384
rect 3112 3372 3114 3394
rect 3150 3389 3156 3390
rect 3150 3385 3151 3389
rect 3155 3385 3156 3389
rect 3150 3384 3156 3385
rect 3110 3371 3116 3372
rect 3110 3367 3111 3371
rect 3115 3367 3116 3371
rect 3110 3366 3116 3367
rect 3152 3363 3154 3384
rect 2831 3362 2835 3363
rect 2831 3357 2835 3358
rect 2839 3362 2843 3363
rect 2839 3357 2843 3358
rect 2935 3362 2939 3363
rect 2935 3357 2939 3358
rect 2975 3362 2979 3363
rect 2975 3357 2979 3358
rect 3039 3362 3043 3363
rect 3039 3357 3043 3358
rect 3119 3362 3123 3363
rect 3119 3357 3123 3358
rect 3151 3362 3155 3363
rect 3151 3357 3155 3358
rect 2782 3355 2788 3356
rect 2782 3351 2783 3355
rect 2787 3351 2788 3355
rect 2782 3350 2788 3351
rect 2230 3331 2236 3332
rect 1766 3327 1772 3328
rect 1766 3323 1767 3327
rect 1771 3323 1772 3327
rect 2230 3327 2231 3331
rect 2235 3327 2236 3331
rect 2230 3326 2236 3327
rect 2366 3331 2372 3332
rect 2366 3327 2367 3331
rect 2371 3327 2372 3331
rect 2366 3326 2372 3327
rect 2502 3331 2508 3332
rect 2502 3327 2503 3331
rect 2507 3327 2508 3331
rect 2774 3331 2780 3332
rect 2502 3326 2508 3327
rect 2638 3327 2644 3328
rect 1766 3322 1772 3323
rect 1806 3323 1812 3324
rect 1768 3295 1770 3322
rect 1806 3319 1807 3323
rect 1811 3319 1812 3323
rect 2638 3323 2639 3327
rect 2643 3323 2644 3327
rect 2774 3327 2775 3331
rect 2779 3327 2780 3331
rect 2774 3326 2780 3327
rect 2638 3322 2644 3323
rect 1806 3318 1812 3319
rect 2158 3320 2164 3321
rect 1808 3299 1810 3318
rect 2158 3316 2159 3320
rect 2163 3316 2164 3320
rect 2158 3315 2164 3316
rect 2294 3320 2300 3321
rect 2294 3316 2295 3320
rect 2299 3316 2300 3320
rect 2294 3315 2300 3316
rect 2430 3320 2436 3321
rect 2430 3316 2431 3320
rect 2435 3316 2436 3320
rect 2430 3315 2436 3316
rect 2566 3320 2572 3321
rect 2566 3316 2567 3320
rect 2571 3316 2572 3320
rect 2566 3315 2572 3316
rect 2160 3299 2162 3315
rect 2296 3299 2298 3315
rect 2432 3299 2434 3315
rect 2568 3299 2570 3315
rect 1807 3298 1811 3299
rect 1767 3294 1771 3295
rect 1807 3293 1811 3294
rect 2087 3298 2091 3299
rect 2087 3293 2091 3294
rect 2159 3298 2163 3299
rect 2159 3293 2163 3294
rect 2239 3298 2243 3299
rect 2239 3293 2243 3294
rect 2295 3298 2299 3299
rect 2295 3293 2299 3294
rect 2399 3298 2403 3299
rect 2399 3293 2403 3294
rect 2431 3298 2435 3299
rect 2431 3293 2435 3294
rect 2559 3298 2563 3299
rect 2559 3293 2563 3294
rect 2567 3298 2571 3299
rect 2567 3293 2571 3294
rect 1767 3289 1771 3290
rect 1768 3270 1770 3289
rect 1808 3274 1810 3293
rect 2088 3277 2090 3293
rect 2240 3277 2242 3293
rect 2400 3277 2402 3293
rect 2560 3277 2562 3293
rect 2086 3276 2092 3277
rect 1806 3273 1812 3274
rect 1766 3269 1772 3270
rect 1766 3265 1767 3269
rect 1771 3265 1772 3269
rect 1806 3269 1807 3273
rect 1811 3269 1812 3273
rect 2086 3272 2087 3276
rect 2091 3272 2092 3276
rect 2086 3271 2092 3272
rect 2238 3276 2244 3277
rect 2238 3272 2239 3276
rect 2243 3272 2244 3276
rect 2238 3271 2244 3272
rect 2398 3276 2404 3277
rect 2398 3272 2399 3276
rect 2403 3272 2404 3276
rect 2398 3271 2404 3272
rect 2558 3276 2564 3277
rect 2558 3272 2559 3276
rect 2563 3272 2564 3276
rect 2558 3271 2564 3272
rect 1806 3268 1812 3269
rect 1766 3264 1772 3265
rect 2158 3267 2164 3268
rect 350 3263 356 3264
rect 350 3259 351 3263
rect 355 3259 356 3263
rect 350 3258 356 3259
rect 534 3263 540 3264
rect 534 3259 535 3263
rect 539 3259 540 3263
rect 534 3258 540 3259
rect 718 3263 724 3264
rect 718 3259 719 3263
rect 723 3259 724 3263
rect 718 3258 724 3259
rect 1114 3263 1120 3264
rect 1114 3259 1115 3263
rect 1119 3259 1120 3263
rect 1114 3258 1120 3259
rect 1246 3263 1252 3264
rect 1246 3259 1247 3263
rect 1251 3259 1252 3263
rect 1246 3258 1252 3259
rect 1414 3263 1420 3264
rect 1414 3259 1415 3263
rect 1419 3259 1420 3263
rect 1414 3258 1420 3259
rect 1574 3263 1580 3264
rect 1574 3259 1575 3263
rect 1579 3259 1580 3263
rect 1574 3258 1580 3259
rect 1734 3263 1740 3264
rect 1734 3259 1735 3263
rect 1739 3259 1740 3263
rect 2158 3263 2159 3267
rect 2163 3263 2164 3267
rect 2158 3262 2164 3263
rect 2310 3267 2316 3268
rect 2310 3263 2311 3267
rect 2315 3263 2316 3267
rect 2310 3262 2316 3263
rect 2478 3267 2484 3268
rect 2478 3263 2479 3267
rect 2483 3263 2484 3267
rect 2478 3262 2484 3263
rect 1734 3258 1740 3259
rect 278 3253 284 3254
rect 278 3249 279 3253
rect 283 3249 284 3253
rect 278 3248 284 3249
rect 280 3223 282 3248
rect 352 3236 354 3258
rect 462 3253 468 3254
rect 462 3249 463 3253
rect 467 3249 468 3253
rect 462 3248 468 3249
rect 350 3235 356 3236
rect 350 3231 351 3235
rect 355 3231 356 3235
rect 350 3230 356 3231
rect 464 3223 466 3248
rect 536 3236 538 3258
rect 646 3253 652 3254
rect 646 3249 647 3253
rect 651 3249 652 3253
rect 646 3248 652 3249
rect 534 3235 540 3236
rect 534 3231 535 3235
rect 539 3231 540 3235
rect 534 3230 540 3231
rect 648 3223 650 3248
rect 720 3236 722 3258
rect 830 3253 836 3254
rect 830 3249 831 3253
rect 835 3249 836 3253
rect 830 3248 836 3249
rect 1006 3253 1012 3254
rect 1006 3249 1007 3253
rect 1011 3249 1012 3253
rect 1006 3248 1012 3249
rect 718 3235 724 3236
rect 718 3231 719 3235
rect 723 3231 724 3235
rect 718 3230 724 3231
rect 832 3223 834 3248
rect 1008 3223 1010 3248
rect 1116 3236 1118 3258
rect 1174 3253 1180 3254
rect 1174 3249 1175 3253
rect 1179 3249 1180 3253
rect 1174 3248 1180 3249
rect 1114 3235 1120 3236
rect 1114 3231 1115 3235
rect 1119 3231 1120 3235
rect 1114 3230 1120 3231
rect 1176 3223 1178 3248
rect 1248 3236 1250 3258
rect 1342 3253 1348 3254
rect 1342 3249 1343 3253
rect 1347 3249 1348 3253
rect 1342 3248 1348 3249
rect 1246 3235 1252 3236
rect 1246 3231 1247 3235
rect 1251 3231 1252 3235
rect 1246 3230 1252 3231
rect 1278 3223 1284 3224
rect 1344 3223 1346 3248
rect 1416 3236 1418 3258
rect 1502 3253 1508 3254
rect 1502 3249 1503 3253
rect 1507 3249 1508 3253
rect 1502 3248 1508 3249
rect 1414 3235 1420 3236
rect 1414 3231 1415 3235
rect 1419 3231 1420 3235
rect 1414 3230 1420 3231
rect 1398 3227 1404 3228
rect 1398 3223 1399 3227
rect 1403 3223 1404 3227
rect 1504 3223 1506 3248
rect 1576 3236 1578 3258
rect 2086 3257 2092 3258
rect 1806 3256 1812 3257
rect 1670 3253 1676 3254
rect 1670 3249 1671 3253
rect 1675 3249 1676 3253
rect 1670 3248 1676 3249
rect 1766 3252 1772 3253
rect 1766 3248 1767 3252
rect 1771 3248 1772 3252
rect 1806 3252 1807 3256
rect 1811 3252 1812 3256
rect 2086 3253 2087 3257
rect 2091 3253 2092 3257
rect 2086 3252 2092 3253
rect 1806 3251 1812 3252
rect 1574 3235 1580 3236
rect 1574 3231 1575 3235
rect 1579 3231 1580 3235
rect 1574 3230 1580 3231
rect 1672 3223 1674 3248
rect 1766 3247 1772 3248
rect 1768 3223 1770 3247
rect 1808 3231 1810 3251
rect 2088 3231 2090 3252
rect 2160 3240 2162 3262
rect 2238 3257 2244 3258
rect 2238 3253 2239 3257
rect 2243 3253 2244 3257
rect 2238 3252 2244 3253
rect 2158 3239 2164 3240
rect 2158 3235 2159 3239
rect 2163 3235 2164 3239
rect 2158 3234 2164 3235
rect 2240 3231 2242 3252
rect 1807 3230 1811 3231
rect 1807 3225 1811 3226
rect 1911 3230 1915 3231
rect 1911 3225 1915 3226
rect 2047 3230 2051 3231
rect 2047 3225 2051 3226
rect 2087 3230 2091 3231
rect 2087 3225 2091 3226
rect 2199 3230 2203 3231
rect 2199 3225 2203 3226
rect 2239 3230 2243 3231
rect 2239 3225 2243 3226
rect 279 3222 283 3223
rect 279 3217 283 3218
rect 327 3222 331 3223
rect 327 3217 331 3218
rect 463 3222 467 3223
rect 463 3217 467 3218
rect 487 3222 491 3223
rect 487 3217 491 3218
rect 647 3222 651 3223
rect 647 3217 651 3218
rect 807 3222 811 3223
rect 807 3217 811 3218
rect 831 3222 835 3223
rect 831 3217 835 3218
rect 967 3222 971 3223
rect 967 3217 971 3218
rect 1007 3222 1011 3223
rect 1007 3217 1011 3218
rect 1135 3222 1139 3223
rect 1135 3217 1139 3218
rect 1175 3222 1179 3223
rect 1278 3219 1279 3223
rect 1283 3219 1284 3223
rect 1278 3218 1284 3219
rect 1303 3222 1307 3223
rect 1175 3217 1179 3218
rect 234 3215 240 3216
rect 234 3211 235 3215
rect 239 3211 240 3215
rect 234 3210 240 3211
rect 254 3215 260 3216
rect 254 3211 255 3215
rect 259 3211 260 3215
rect 254 3210 260 3211
rect 110 3196 111 3200
rect 115 3196 116 3200
rect 110 3195 116 3196
rect 182 3199 188 3200
rect 182 3195 183 3199
rect 187 3195 188 3199
rect 182 3194 188 3195
rect 256 3192 258 3210
rect 328 3200 330 3217
rect 398 3215 404 3216
rect 398 3211 399 3215
rect 403 3211 404 3215
rect 398 3210 404 3211
rect 326 3199 332 3200
rect 326 3195 327 3199
rect 331 3195 332 3199
rect 326 3194 332 3195
rect 400 3192 402 3210
rect 488 3200 490 3217
rect 558 3215 564 3216
rect 558 3211 559 3215
rect 563 3211 564 3215
rect 558 3210 564 3211
rect 486 3199 492 3200
rect 486 3195 487 3199
rect 491 3195 492 3199
rect 486 3194 492 3195
rect 560 3192 562 3210
rect 648 3200 650 3217
rect 718 3215 724 3216
rect 718 3211 719 3215
rect 723 3211 724 3215
rect 718 3210 724 3211
rect 646 3199 652 3200
rect 646 3195 647 3199
rect 651 3195 652 3199
rect 646 3194 652 3195
rect 720 3192 722 3210
rect 808 3200 810 3217
rect 968 3200 970 3217
rect 1094 3211 1100 3212
rect 1094 3207 1095 3211
rect 1099 3207 1100 3211
rect 1094 3206 1100 3207
rect 806 3199 812 3200
rect 806 3195 807 3199
rect 811 3195 812 3199
rect 806 3194 812 3195
rect 966 3199 972 3200
rect 966 3195 967 3199
rect 971 3195 972 3199
rect 966 3194 972 3195
rect 1096 3192 1098 3206
rect 1136 3200 1138 3217
rect 1250 3215 1256 3216
rect 1250 3211 1251 3215
rect 1255 3211 1256 3215
rect 1250 3210 1256 3211
rect 1134 3199 1140 3200
rect 1134 3195 1135 3199
rect 1139 3195 1140 3199
rect 1134 3194 1140 3195
rect 1252 3192 1254 3210
rect 254 3191 260 3192
rect 254 3187 255 3191
rect 259 3187 260 3191
rect 254 3186 260 3187
rect 398 3191 404 3192
rect 398 3187 399 3191
rect 403 3187 404 3191
rect 398 3186 404 3187
rect 558 3191 564 3192
rect 558 3187 559 3191
rect 563 3187 564 3191
rect 558 3186 564 3187
rect 718 3191 724 3192
rect 718 3187 719 3191
rect 723 3187 724 3191
rect 718 3186 724 3187
rect 734 3191 740 3192
rect 734 3187 735 3191
rect 739 3187 740 3191
rect 734 3186 740 3187
rect 1094 3191 1100 3192
rect 1094 3187 1095 3191
rect 1099 3187 1100 3191
rect 1094 3186 1100 3187
rect 1250 3191 1256 3192
rect 1250 3187 1251 3191
rect 1255 3187 1256 3191
rect 1250 3186 1256 3187
rect 110 3183 116 3184
rect 110 3179 111 3183
rect 115 3179 116 3183
rect 110 3178 116 3179
rect 182 3180 188 3181
rect 112 3159 114 3178
rect 182 3176 183 3180
rect 187 3176 188 3180
rect 182 3175 188 3176
rect 326 3180 332 3181
rect 326 3176 327 3180
rect 331 3176 332 3180
rect 326 3175 332 3176
rect 486 3180 492 3181
rect 486 3176 487 3180
rect 491 3176 492 3180
rect 486 3175 492 3176
rect 646 3180 652 3181
rect 646 3176 647 3180
rect 651 3176 652 3180
rect 646 3175 652 3176
rect 184 3159 186 3175
rect 328 3159 330 3175
rect 488 3159 490 3175
rect 648 3159 650 3175
rect 111 3158 115 3159
rect 111 3153 115 3154
rect 183 3158 187 3159
rect 183 3153 187 3154
rect 327 3158 331 3159
rect 327 3153 331 3154
rect 367 3158 371 3159
rect 367 3153 371 3154
rect 487 3158 491 3159
rect 487 3153 491 3154
rect 607 3158 611 3159
rect 607 3153 611 3154
rect 647 3158 651 3159
rect 647 3153 651 3154
rect 727 3158 731 3159
rect 727 3153 731 3154
rect 112 3134 114 3153
rect 368 3137 370 3153
rect 418 3147 424 3148
rect 418 3143 419 3147
rect 423 3143 424 3147
rect 418 3142 424 3143
rect 366 3136 372 3137
rect 110 3133 116 3134
rect 110 3129 111 3133
rect 115 3129 116 3133
rect 366 3132 367 3136
rect 371 3132 372 3136
rect 366 3131 372 3132
rect 110 3128 116 3129
rect 366 3117 372 3118
rect 110 3116 116 3117
rect 110 3112 111 3116
rect 115 3112 116 3116
rect 366 3113 367 3117
rect 371 3113 372 3117
rect 366 3112 372 3113
rect 110 3111 116 3112
rect 112 3091 114 3111
rect 368 3091 370 3112
rect 420 3100 422 3142
rect 488 3137 490 3153
rect 608 3137 610 3153
rect 728 3137 730 3153
rect 736 3148 738 3186
rect 806 3180 812 3181
rect 806 3176 807 3180
rect 811 3176 812 3180
rect 806 3175 812 3176
rect 966 3180 972 3181
rect 966 3176 967 3180
rect 971 3176 972 3180
rect 966 3175 972 3176
rect 1134 3180 1140 3181
rect 1134 3176 1135 3180
rect 1139 3176 1140 3180
rect 1134 3175 1140 3176
rect 808 3159 810 3175
rect 968 3159 970 3175
rect 1136 3159 1138 3175
rect 807 3158 811 3159
rect 807 3153 811 3154
rect 847 3158 851 3159
rect 847 3153 851 3154
rect 967 3158 971 3159
rect 967 3153 971 3154
rect 1079 3158 1083 3159
rect 1079 3153 1083 3154
rect 1135 3158 1139 3159
rect 1135 3153 1139 3154
rect 1199 3158 1203 3159
rect 1199 3153 1203 3154
rect 734 3147 740 3148
rect 734 3143 735 3147
rect 739 3143 740 3147
rect 734 3142 740 3143
rect 848 3137 850 3153
rect 968 3137 970 3153
rect 1080 3137 1082 3153
rect 1200 3137 1202 3153
rect 486 3136 492 3137
rect 486 3132 487 3136
rect 491 3132 492 3136
rect 486 3131 492 3132
rect 606 3136 612 3137
rect 606 3132 607 3136
rect 611 3132 612 3136
rect 606 3131 612 3132
rect 726 3136 732 3137
rect 726 3132 727 3136
rect 731 3132 732 3136
rect 726 3131 732 3132
rect 846 3136 852 3137
rect 846 3132 847 3136
rect 851 3132 852 3136
rect 846 3131 852 3132
rect 966 3136 972 3137
rect 966 3132 967 3136
rect 971 3132 972 3136
rect 966 3131 972 3132
rect 1078 3136 1084 3137
rect 1078 3132 1079 3136
rect 1083 3132 1084 3136
rect 1078 3131 1084 3132
rect 1198 3136 1204 3137
rect 1198 3132 1199 3136
rect 1203 3132 1204 3136
rect 1198 3131 1204 3132
rect 1280 3128 1282 3218
rect 1303 3217 1307 3218
rect 1343 3222 1347 3223
rect 1398 3222 1404 3223
rect 1471 3222 1475 3223
rect 1343 3217 1347 3218
rect 1304 3200 1306 3217
rect 1374 3215 1380 3216
rect 1374 3211 1375 3215
rect 1379 3211 1380 3215
rect 1374 3210 1380 3211
rect 1302 3199 1308 3200
rect 1302 3195 1303 3199
rect 1307 3195 1308 3199
rect 1302 3194 1308 3195
rect 1376 3192 1378 3210
rect 1400 3192 1402 3222
rect 1471 3217 1475 3218
rect 1503 3222 1507 3223
rect 1503 3217 1507 3218
rect 1671 3222 1675 3223
rect 1671 3217 1675 3218
rect 1767 3222 1771 3223
rect 1767 3217 1771 3218
rect 1472 3200 1474 3217
rect 1768 3201 1770 3217
rect 1808 3209 1810 3225
rect 1806 3208 1812 3209
rect 1912 3208 1914 3225
rect 1962 3223 1968 3224
rect 1962 3219 1963 3223
rect 1967 3219 1968 3223
rect 1962 3218 1968 3219
rect 1982 3223 1988 3224
rect 1982 3219 1983 3223
rect 1987 3219 1988 3223
rect 1982 3218 1988 3219
rect 1806 3204 1807 3208
rect 1811 3204 1812 3208
rect 1806 3203 1812 3204
rect 1910 3207 1916 3208
rect 1910 3203 1911 3207
rect 1915 3203 1916 3207
rect 1910 3202 1916 3203
rect 1766 3200 1772 3201
rect 1470 3199 1476 3200
rect 1470 3195 1471 3199
rect 1475 3195 1476 3199
rect 1766 3196 1767 3200
rect 1771 3196 1772 3200
rect 1766 3195 1772 3196
rect 1470 3194 1476 3195
rect 1374 3191 1380 3192
rect 1374 3187 1375 3191
rect 1379 3187 1380 3191
rect 1374 3186 1380 3187
rect 1398 3191 1404 3192
rect 1398 3187 1399 3191
rect 1403 3187 1404 3191
rect 1398 3186 1404 3187
rect 1806 3191 1812 3192
rect 1806 3187 1807 3191
rect 1811 3187 1812 3191
rect 1806 3186 1812 3187
rect 1910 3188 1916 3189
rect 1766 3183 1772 3184
rect 1302 3180 1308 3181
rect 1302 3176 1303 3180
rect 1307 3176 1308 3180
rect 1302 3175 1308 3176
rect 1470 3180 1476 3181
rect 1470 3176 1471 3180
rect 1475 3176 1476 3180
rect 1766 3179 1767 3183
rect 1771 3179 1772 3183
rect 1766 3178 1772 3179
rect 1470 3175 1476 3176
rect 1304 3159 1306 3175
rect 1472 3159 1474 3175
rect 1768 3159 1770 3178
rect 1808 3167 1810 3186
rect 1910 3184 1911 3188
rect 1915 3184 1916 3188
rect 1910 3183 1916 3184
rect 1912 3167 1914 3183
rect 1964 3180 1966 3218
rect 1984 3200 1986 3218
rect 2048 3208 2050 3225
rect 2118 3223 2124 3224
rect 2118 3219 2119 3223
rect 2123 3219 2124 3223
rect 2118 3218 2124 3219
rect 2046 3207 2052 3208
rect 2046 3203 2047 3207
rect 2051 3203 2052 3207
rect 2046 3202 2052 3203
rect 2120 3200 2122 3218
rect 2200 3208 2202 3225
rect 2312 3224 2314 3262
rect 2398 3257 2404 3258
rect 2398 3253 2399 3257
rect 2403 3253 2404 3257
rect 2398 3252 2404 3253
rect 2400 3231 2402 3252
rect 2480 3240 2482 3262
rect 2558 3257 2564 3258
rect 2558 3253 2559 3257
rect 2563 3253 2564 3257
rect 2558 3252 2564 3253
rect 2478 3239 2484 3240
rect 2478 3235 2479 3239
rect 2483 3235 2484 3239
rect 2478 3234 2484 3235
rect 2560 3231 2562 3252
rect 2640 3240 2642 3322
rect 2702 3320 2708 3321
rect 2702 3316 2703 3320
rect 2707 3316 2708 3320
rect 2702 3315 2708 3316
rect 2704 3299 2706 3315
rect 2703 3298 2707 3299
rect 2703 3293 2707 3294
rect 2719 3298 2723 3299
rect 2719 3293 2723 3294
rect 2720 3277 2722 3293
rect 2718 3276 2724 3277
rect 2718 3272 2719 3276
rect 2723 3272 2724 3276
rect 2718 3271 2724 3272
rect 2784 3268 2786 3350
rect 2840 3340 2842 3357
rect 2918 3355 2924 3356
rect 2918 3351 2919 3355
rect 2923 3351 2924 3355
rect 2918 3350 2924 3351
rect 2838 3339 2844 3340
rect 2838 3335 2839 3339
rect 2843 3335 2844 3339
rect 2838 3334 2844 3335
rect 2920 3332 2922 3350
rect 2976 3340 2978 3357
rect 3054 3355 3060 3356
rect 3054 3351 3055 3355
rect 3059 3351 3060 3355
rect 3054 3350 3060 3351
rect 2974 3339 2980 3340
rect 2974 3335 2975 3339
rect 2979 3335 2980 3339
rect 2974 3334 2980 3335
rect 3056 3332 3058 3350
rect 3120 3340 3122 3357
rect 3216 3356 3218 3394
rect 3462 3388 3468 3389
rect 3462 3384 3463 3388
rect 3467 3384 3468 3388
rect 3462 3383 3468 3384
rect 3464 3363 3466 3383
rect 3463 3362 3467 3363
rect 3463 3357 3467 3358
rect 3214 3355 3220 3356
rect 3214 3351 3215 3355
rect 3219 3351 3220 3355
rect 3214 3350 3220 3351
rect 3464 3341 3466 3357
rect 3462 3340 3468 3341
rect 3118 3339 3124 3340
rect 3118 3335 3119 3339
rect 3123 3335 3124 3339
rect 3462 3336 3463 3340
rect 3467 3336 3468 3340
rect 3462 3335 3468 3336
rect 3118 3334 3124 3335
rect 2918 3331 2924 3332
rect 2910 3327 2916 3328
rect 2910 3323 2911 3327
rect 2915 3323 2916 3327
rect 2918 3327 2919 3331
rect 2923 3327 2924 3331
rect 2918 3326 2924 3327
rect 3054 3331 3060 3332
rect 3054 3327 3055 3331
rect 3059 3327 3060 3331
rect 3054 3326 3060 3327
rect 2910 3322 2916 3323
rect 3462 3323 3468 3324
rect 2838 3320 2844 3321
rect 2838 3316 2839 3320
rect 2843 3316 2844 3320
rect 2838 3315 2844 3316
rect 2840 3299 2842 3315
rect 2839 3298 2843 3299
rect 2839 3293 2843 3294
rect 2879 3298 2883 3299
rect 2879 3293 2883 3294
rect 2880 3277 2882 3293
rect 2878 3276 2884 3277
rect 2878 3272 2879 3276
rect 2883 3272 2884 3276
rect 2878 3271 2884 3272
rect 2782 3267 2788 3268
rect 2782 3263 2783 3267
rect 2787 3263 2788 3267
rect 2782 3262 2788 3263
rect 2718 3257 2724 3258
rect 2718 3253 2719 3257
rect 2723 3253 2724 3257
rect 2718 3252 2724 3253
rect 2878 3257 2884 3258
rect 2878 3253 2879 3257
rect 2883 3253 2884 3257
rect 2878 3252 2884 3253
rect 2638 3239 2644 3240
rect 2638 3235 2639 3239
rect 2643 3235 2644 3239
rect 2638 3234 2644 3235
rect 2720 3231 2722 3252
rect 2758 3239 2764 3240
rect 2758 3235 2759 3239
rect 2763 3235 2764 3239
rect 2758 3234 2764 3235
rect 2359 3230 2363 3231
rect 2359 3225 2363 3226
rect 2399 3230 2403 3231
rect 2399 3225 2403 3226
rect 2527 3230 2531 3231
rect 2527 3225 2531 3226
rect 2559 3230 2563 3231
rect 2559 3225 2563 3226
rect 2687 3230 2691 3231
rect 2687 3225 2691 3226
rect 2719 3230 2723 3231
rect 2719 3225 2723 3226
rect 2310 3223 2316 3224
rect 2310 3219 2311 3223
rect 2315 3219 2316 3223
rect 2310 3218 2316 3219
rect 2360 3208 2362 3225
rect 2430 3223 2436 3224
rect 2430 3219 2431 3223
rect 2435 3219 2436 3223
rect 2430 3218 2436 3219
rect 2198 3207 2204 3208
rect 2198 3203 2199 3207
rect 2203 3203 2204 3207
rect 2198 3202 2204 3203
rect 2358 3207 2364 3208
rect 2358 3203 2359 3207
rect 2363 3203 2364 3207
rect 2358 3202 2364 3203
rect 2432 3200 2434 3218
rect 2528 3208 2530 3225
rect 2688 3208 2690 3225
rect 2526 3207 2532 3208
rect 2526 3203 2527 3207
rect 2531 3203 2532 3207
rect 2526 3202 2532 3203
rect 2686 3207 2692 3208
rect 2686 3203 2687 3207
rect 2691 3203 2692 3207
rect 2686 3202 2692 3203
rect 2760 3200 2762 3234
rect 2880 3231 2882 3252
rect 2912 3240 2914 3322
rect 2974 3320 2980 3321
rect 2974 3316 2975 3320
rect 2979 3316 2980 3320
rect 2974 3315 2980 3316
rect 3118 3320 3124 3321
rect 3118 3316 3119 3320
rect 3123 3316 3124 3320
rect 3462 3319 3463 3323
rect 3467 3319 3468 3323
rect 3462 3318 3468 3319
rect 3118 3315 3124 3316
rect 2976 3299 2978 3315
rect 3120 3299 3122 3315
rect 3464 3299 3466 3318
rect 2975 3298 2979 3299
rect 2975 3293 2979 3294
rect 3039 3298 3043 3299
rect 3039 3293 3043 3294
rect 3119 3298 3123 3299
rect 3119 3293 3123 3294
rect 3199 3298 3203 3299
rect 3199 3293 3203 3294
rect 3463 3298 3467 3299
rect 3463 3293 3467 3294
rect 3040 3277 3042 3293
rect 3200 3277 3202 3293
rect 3038 3276 3044 3277
rect 3038 3272 3039 3276
rect 3043 3272 3044 3276
rect 3038 3271 3044 3272
rect 3198 3276 3204 3277
rect 3198 3272 3199 3276
rect 3203 3272 3204 3276
rect 3464 3274 3466 3293
rect 3198 3271 3204 3272
rect 3462 3273 3468 3274
rect 3462 3269 3463 3273
rect 3467 3269 3468 3273
rect 3462 3268 3468 3269
rect 2950 3267 2956 3268
rect 2950 3263 2951 3267
rect 2955 3263 2956 3267
rect 2950 3262 2956 3263
rect 3110 3267 3116 3268
rect 3110 3263 3111 3267
rect 3115 3263 3116 3267
rect 3110 3262 3116 3263
rect 3262 3267 3268 3268
rect 3262 3263 3263 3267
rect 3267 3263 3268 3267
rect 3262 3262 3268 3263
rect 2952 3240 2954 3262
rect 3038 3257 3044 3258
rect 3038 3253 3039 3257
rect 3043 3253 3044 3257
rect 3038 3252 3044 3253
rect 2910 3239 2916 3240
rect 2910 3235 2911 3239
rect 2915 3235 2916 3239
rect 2910 3234 2916 3235
rect 2950 3239 2956 3240
rect 2950 3235 2951 3239
rect 2955 3235 2956 3239
rect 2950 3234 2956 3235
rect 3040 3231 3042 3252
rect 3112 3240 3114 3262
rect 3198 3257 3204 3258
rect 3198 3253 3199 3257
rect 3203 3253 3204 3257
rect 3198 3252 3204 3253
rect 3110 3239 3116 3240
rect 3110 3235 3111 3239
rect 3115 3235 3116 3239
rect 3110 3234 3116 3235
rect 3200 3231 3202 3252
rect 2847 3230 2851 3231
rect 2847 3225 2851 3226
rect 2879 3230 2883 3231
rect 2879 3225 2883 3226
rect 3007 3230 3011 3231
rect 3007 3225 3011 3226
rect 3039 3230 3043 3231
rect 3039 3225 3043 3226
rect 3167 3230 3171 3231
rect 3167 3225 3171 3226
rect 3199 3230 3203 3231
rect 3199 3225 3203 3226
rect 2806 3223 2812 3224
rect 2806 3219 2807 3223
rect 2811 3219 2812 3223
rect 2806 3218 2812 3219
rect 2830 3223 2836 3224
rect 2830 3219 2831 3223
rect 2835 3219 2836 3223
rect 2830 3218 2836 3219
rect 2808 3200 2810 3218
rect 1982 3199 1988 3200
rect 1982 3195 1983 3199
rect 1987 3195 1988 3199
rect 1982 3194 1988 3195
rect 2118 3199 2124 3200
rect 2118 3195 2119 3199
rect 2123 3195 2124 3199
rect 2430 3199 2436 3200
rect 2118 3194 2124 3195
rect 2270 3195 2276 3196
rect 2270 3191 2271 3195
rect 2275 3191 2276 3195
rect 2430 3195 2431 3199
rect 2435 3195 2436 3199
rect 2430 3194 2436 3195
rect 2478 3199 2484 3200
rect 2478 3195 2479 3199
rect 2483 3195 2484 3199
rect 2478 3194 2484 3195
rect 2758 3199 2764 3200
rect 2758 3195 2759 3199
rect 2763 3195 2764 3199
rect 2758 3194 2764 3195
rect 2806 3199 2812 3200
rect 2806 3195 2807 3199
rect 2811 3195 2812 3199
rect 2806 3194 2812 3195
rect 2270 3190 2276 3191
rect 2046 3188 2052 3189
rect 2046 3184 2047 3188
rect 2051 3184 2052 3188
rect 2046 3183 2052 3184
rect 2198 3188 2204 3189
rect 2198 3184 2199 3188
rect 2203 3184 2204 3188
rect 2198 3183 2204 3184
rect 1962 3179 1968 3180
rect 1962 3175 1963 3179
rect 1967 3175 1968 3179
rect 1962 3174 1968 3175
rect 2048 3167 2050 3183
rect 2200 3167 2202 3183
rect 1807 3166 1811 3167
rect 1807 3161 1811 3162
rect 1831 3166 1835 3167
rect 1831 3161 1835 3162
rect 1911 3166 1915 3167
rect 1911 3161 1915 3162
rect 2007 3166 2011 3167
rect 2007 3161 2011 3162
rect 2047 3166 2051 3167
rect 2047 3161 2051 3162
rect 2199 3166 2203 3167
rect 2199 3161 2203 3162
rect 2207 3166 2211 3167
rect 2207 3161 2211 3162
rect 1303 3158 1307 3159
rect 1303 3153 1307 3154
rect 1319 3158 1323 3159
rect 1319 3153 1323 3154
rect 1471 3158 1475 3159
rect 1471 3153 1475 3154
rect 1767 3158 1771 3159
rect 1767 3153 1771 3154
rect 1320 3137 1322 3153
rect 1318 3136 1324 3137
rect 1318 3132 1319 3136
rect 1323 3132 1324 3136
rect 1768 3134 1770 3153
rect 1808 3142 1810 3161
rect 1832 3145 1834 3161
rect 2008 3145 2010 3161
rect 2208 3145 2210 3161
rect 1830 3144 1836 3145
rect 1806 3141 1812 3142
rect 1806 3137 1807 3141
rect 1811 3137 1812 3141
rect 1830 3140 1831 3144
rect 1835 3140 1836 3144
rect 1830 3139 1836 3140
rect 2006 3144 2012 3145
rect 2006 3140 2007 3144
rect 2011 3140 2012 3144
rect 2006 3139 2012 3140
rect 2206 3144 2212 3145
rect 2206 3140 2207 3144
rect 2211 3140 2212 3144
rect 2206 3139 2212 3140
rect 1806 3136 1812 3137
rect 1894 3135 1900 3136
rect 1318 3131 1324 3132
rect 1766 3133 1772 3134
rect 1766 3129 1767 3133
rect 1771 3129 1772 3133
rect 1894 3131 1895 3135
rect 1899 3131 1900 3135
rect 1894 3130 1900 3131
rect 1910 3135 1916 3136
rect 1910 3131 1911 3135
rect 1915 3131 1916 3135
rect 1910 3130 1916 3131
rect 1766 3128 1772 3129
rect 438 3127 444 3128
rect 438 3123 439 3127
rect 443 3123 444 3127
rect 438 3122 444 3123
rect 558 3127 564 3128
rect 558 3123 559 3127
rect 563 3123 564 3127
rect 558 3122 564 3123
rect 678 3127 684 3128
rect 678 3123 679 3127
rect 683 3123 684 3127
rect 678 3122 684 3123
rect 686 3127 692 3128
rect 686 3123 687 3127
rect 691 3123 692 3127
rect 686 3122 692 3123
rect 918 3127 924 3128
rect 918 3123 919 3127
rect 923 3123 924 3127
rect 918 3122 924 3123
rect 1038 3127 1044 3128
rect 1038 3123 1039 3127
rect 1043 3123 1044 3127
rect 1038 3122 1044 3123
rect 1150 3127 1156 3128
rect 1150 3123 1151 3127
rect 1155 3123 1156 3127
rect 1150 3122 1156 3123
rect 1270 3127 1276 3128
rect 1270 3123 1271 3127
rect 1275 3123 1276 3127
rect 1270 3122 1276 3123
rect 1278 3127 1284 3128
rect 1278 3123 1279 3127
rect 1283 3123 1284 3127
rect 1830 3125 1836 3126
rect 1278 3122 1284 3123
rect 1806 3124 1812 3125
rect 440 3100 442 3122
rect 486 3117 492 3118
rect 486 3113 487 3117
rect 491 3113 492 3117
rect 486 3112 492 3113
rect 418 3099 424 3100
rect 418 3095 419 3099
rect 423 3095 424 3099
rect 418 3094 424 3095
rect 438 3099 444 3100
rect 438 3095 439 3099
rect 443 3095 444 3099
rect 438 3094 444 3095
rect 488 3091 490 3112
rect 560 3100 562 3122
rect 606 3117 612 3118
rect 606 3113 607 3117
rect 611 3113 612 3117
rect 606 3112 612 3113
rect 558 3099 564 3100
rect 558 3095 559 3099
rect 563 3095 564 3099
rect 558 3094 564 3095
rect 608 3091 610 3112
rect 680 3100 682 3122
rect 678 3099 684 3100
rect 678 3095 679 3099
rect 683 3095 684 3099
rect 678 3094 684 3095
rect 688 3092 690 3122
rect 726 3117 732 3118
rect 726 3113 727 3117
rect 731 3113 732 3117
rect 726 3112 732 3113
rect 846 3117 852 3118
rect 846 3113 847 3117
rect 851 3113 852 3117
rect 846 3112 852 3113
rect 686 3091 692 3092
rect 728 3091 730 3112
rect 848 3091 850 3112
rect 920 3100 922 3122
rect 966 3117 972 3118
rect 966 3113 967 3117
rect 971 3113 972 3117
rect 966 3112 972 3113
rect 918 3099 924 3100
rect 918 3095 919 3099
rect 923 3095 924 3099
rect 918 3094 924 3095
rect 968 3091 970 3112
rect 1040 3100 1042 3122
rect 1078 3117 1084 3118
rect 1078 3113 1079 3117
rect 1083 3113 1084 3117
rect 1078 3112 1084 3113
rect 1038 3099 1044 3100
rect 1038 3095 1039 3099
rect 1043 3095 1044 3099
rect 1038 3094 1044 3095
rect 1080 3091 1082 3112
rect 1152 3100 1154 3122
rect 1198 3117 1204 3118
rect 1198 3113 1199 3117
rect 1203 3113 1204 3117
rect 1198 3112 1204 3113
rect 1150 3099 1156 3100
rect 1150 3095 1151 3099
rect 1155 3095 1156 3099
rect 1150 3094 1156 3095
rect 1134 3091 1140 3092
rect 1200 3091 1202 3112
rect 1272 3100 1274 3122
rect 1806 3120 1807 3124
rect 1811 3120 1812 3124
rect 1830 3121 1831 3125
rect 1835 3121 1836 3125
rect 1830 3120 1836 3121
rect 1806 3119 1812 3120
rect 1318 3117 1324 3118
rect 1318 3113 1319 3117
rect 1323 3113 1324 3117
rect 1318 3112 1324 3113
rect 1766 3116 1772 3117
rect 1766 3112 1767 3116
rect 1771 3112 1772 3116
rect 1270 3099 1276 3100
rect 1270 3095 1271 3099
rect 1275 3095 1276 3099
rect 1270 3094 1276 3095
rect 1320 3091 1322 3112
rect 1766 3111 1772 3112
rect 1768 3091 1770 3111
rect 1808 3095 1810 3119
rect 1832 3095 1834 3120
rect 1807 3094 1811 3095
rect 111 3090 115 3091
rect 111 3085 115 3086
rect 367 3090 371 3091
rect 367 3085 371 3086
rect 439 3090 443 3091
rect 439 3085 443 3086
rect 487 3090 491 3091
rect 487 3085 491 3086
rect 527 3090 531 3091
rect 527 3085 531 3086
rect 607 3090 611 3091
rect 607 3085 611 3086
rect 615 3090 619 3091
rect 686 3087 687 3091
rect 691 3087 692 3091
rect 686 3086 692 3087
rect 703 3090 707 3091
rect 615 3085 619 3086
rect 703 3085 707 3086
rect 727 3090 731 3091
rect 727 3085 731 3086
rect 791 3090 795 3091
rect 791 3085 795 3086
rect 847 3090 851 3091
rect 847 3085 851 3086
rect 879 3090 883 3091
rect 879 3085 883 3086
rect 967 3090 971 3091
rect 967 3085 971 3086
rect 1055 3090 1059 3091
rect 1055 3085 1059 3086
rect 1079 3090 1083 3091
rect 1134 3087 1135 3091
rect 1139 3087 1140 3091
rect 1134 3086 1140 3087
rect 1143 3090 1147 3091
rect 1079 3085 1083 3086
rect 112 3069 114 3085
rect 110 3068 116 3069
rect 440 3068 442 3085
rect 510 3083 516 3084
rect 510 3079 511 3083
rect 515 3079 516 3083
rect 510 3078 516 3079
rect 110 3064 111 3068
rect 115 3064 116 3068
rect 110 3063 116 3064
rect 438 3067 444 3068
rect 438 3063 439 3067
rect 443 3063 444 3067
rect 438 3062 444 3063
rect 512 3060 514 3078
rect 528 3068 530 3085
rect 598 3083 604 3084
rect 598 3079 599 3083
rect 603 3079 604 3083
rect 598 3078 604 3079
rect 526 3067 532 3068
rect 526 3063 527 3067
rect 531 3063 532 3067
rect 526 3062 532 3063
rect 600 3060 602 3078
rect 616 3068 618 3085
rect 686 3083 692 3084
rect 686 3079 687 3083
rect 691 3079 692 3083
rect 686 3078 692 3079
rect 614 3067 620 3068
rect 614 3063 615 3067
rect 619 3063 620 3067
rect 614 3062 620 3063
rect 688 3060 690 3078
rect 704 3068 706 3085
rect 774 3083 780 3084
rect 774 3079 775 3083
rect 779 3079 780 3083
rect 774 3078 780 3079
rect 702 3067 708 3068
rect 702 3063 703 3067
rect 707 3063 708 3067
rect 702 3062 708 3063
rect 776 3060 778 3078
rect 792 3068 794 3085
rect 880 3068 882 3085
rect 926 3083 932 3084
rect 926 3079 927 3083
rect 931 3079 932 3083
rect 926 3078 932 3079
rect 950 3083 956 3084
rect 950 3079 951 3083
rect 955 3079 956 3083
rect 950 3078 956 3079
rect 928 3075 930 3078
rect 928 3073 938 3075
rect 790 3067 796 3068
rect 790 3063 791 3067
rect 795 3063 796 3067
rect 790 3062 796 3063
rect 878 3067 884 3068
rect 878 3063 879 3067
rect 883 3063 884 3067
rect 878 3062 884 3063
rect 510 3059 516 3060
rect 510 3055 511 3059
rect 515 3055 516 3059
rect 510 3054 516 3055
rect 598 3059 604 3060
rect 598 3055 599 3059
rect 603 3055 604 3059
rect 598 3054 604 3055
rect 686 3059 692 3060
rect 686 3055 687 3059
rect 691 3055 692 3059
rect 686 3054 692 3055
rect 774 3059 780 3060
rect 774 3055 775 3059
rect 779 3055 780 3059
rect 774 3054 780 3055
rect 862 3055 868 3056
rect 110 3051 116 3052
rect 110 3047 111 3051
rect 115 3047 116 3051
rect 862 3051 863 3055
rect 867 3051 868 3055
rect 862 3050 868 3051
rect 110 3046 116 3047
rect 438 3048 444 3049
rect 112 3019 114 3046
rect 438 3044 439 3048
rect 443 3044 444 3048
rect 438 3043 444 3044
rect 526 3048 532 3049
rect 526 3044 527 3048
rect 531 3044 532 3048
rect 526 3043 532 3044
rect 614 3048 620 3049
rect 614 3044 615 3048
rect 619 3044 620 3048
rect 614 3043 620 3044
rect 702 3048 708 3049
rect 702 3044 703 3048
rect 707 3044 708 3048
rect 702 3043 708 3044
rect 790 3048 796 3049
rect 790 3044 791 3048
rect 795 3044 796 3048
rect 790 3043 796 3044
rect 440 3019 442 3043
rect 528 3019 530 3043
rect 616 3019 618 3043
rect 704 3019 706 3043
rect 792 3019 794 3043
rect 111 3018 115 3019
rect 111 3013 115 3014
rect 439 3018 443 3019
rect 439 3013 443 3014
rect 503 3018 507 3019
rect 503 3013 507 3014
rect 527 3018 531 3019
rect 527 3013 531 3014
rect 591 3018 595 3019
rect 591 3013 595 3014
rect 615 3018 619 3019
rect 615 3013 619 3014
rect 679 3018 683 3019
rect 679 3013 683 3014
rect 703 3018 707 3019
rect 703 3013 707 3014
rect 767 3018 771 3019
rect 767 3013 771 3014
rect 791 3018 795 3019
rect 791 3013 795 3014
rect 855 3018 859 3019
rect 855 3013 859 3014
rect 112 2994 114 3013
rect 504 2997 506 3013
rect 592 2997 594 3013
rect 680 2997 682 3013
rect 768 2997 770 3013
rect 856 2997 858 3013
rect 502 2996 508 2997
rect 110 2993 116 2994
rect 110 2989 111 2993
rect 115 2989 116 2993
rect 502 2992 503 2996
rect 507 2992 508 2996
rect 502 2991 508 2992
rect 590 2996 596 2997
rect 590 2992 591 2996
rect 595 2992 596 2996
rect 590 2991 596 2992
rect 678 2996 684 2997
rect 678 2992 679 2996
rect 683 2992 684 2996
rect 678 2991 684 2992
rect 766 2996 772 2997
rect 766 2992 767 2996
rect 771 2992 772 2996
rect 766 2991 772 2992
rect 854 2996 860 2997
rect 854 2992 855 2996
rect 859 2992 860 2996
rect 854 2991 860 2992
rect 110 2988 116 2989
rect 574 2987 580 2988
rect 574 2983 575 2987
rect 579 2983 580 2987
rect 574 2982 580 2983
rect 662 2987 668 2988
rect 662 2983 663 2987
rect 667 2983 668 2987
rect 662 2982 668 2983
rect 750 2987 756 2988
rect 750 2983 751 2987
rect 755 2983 756 2987
rect 750 2982 756 2983
rect 758 2987 764 2988
rect 758 2983 759 2987
rect 763 2983 764 2987
rect 758 2982 764 2983
rect 846 2987 852 2988
rect 846 2983 847 2987
rect 851 2983 852 2987
rect 846 2982 852 2983
rect 502 2977 508 2978
rect 110 2976 116 2977
rect 110 2972 111 2976
rect 115 2972 116 2976
rect 502 2973 503 2977
rect 507 2973 508 2977
rect 502 2972 508 2973
rect 110 2971 116 2972
rect 112 2943 114 2971
rect 504 2943 506 2972
rect 576 2960 578 2982
rect 590 2977 596 2978
rect 590 2973 591 2977
rect 595 2973 596 2977
rect 590 2972 596 2973
rect 574 2959 580 2960
rect 574 2955 575 2959
rect 579 2955 580 2959
rect 574 2954 580 2955
rect 592 2943 594 2972
rect 664 2960 666 2982
rect 678 2977 684 2978
rect 678 2973 679 2977
rect 683 2973 684 2977
rect 678 2972 684 2973
rect 662 2959 668 2960
rect 662 2955 663 2959
rect 667 2955 668 2959
rect 662 2954 668 2955
rect 680 2943 682 2972
rect 111 2942 115 2943
rect 111 2937 115 2938
rect 327 2942 331 2943
rect 327 2937 331 2938
rect 447 2942 451 2943
rect 447 2937 451 2938
rect 503 2942 507 2943
rect 503 2937 507 2938
rect 575 2942 579 2943
rect 575 2937 579 2938
rect 591 2942 595 2943
rect 591 2937 595 2938
rect 679 2942 683 2943
rect 679 2937 683 2938
rect 711 2942 715 2943
rect 711 2937 715 2938
rect 112 2921 114 2937
rect 110 2920 116 2921
rect 328 2920 330 2937
rect 398 2935 404 2936
rect 398 2931 399 2935
rect 403 2931 404 2935
rect 398 2930 404 2931
rect 110 2916 111 2920
rect 115 2916 116 2920
rect 110 2915 116 2916
rect 326 2919 332 2920
rect 326 2915 327 2919
rect 331 2915 332 2919
rect 326 2914 332 2915
rect 400 2912 402 2930
rect 448 2920 450 2937
rect 518 2935 524 2936
rect 518 2931 519 2935
rect 523 2931 524 2935
rect 518 2930 524 2931
rect 446 2919 452 2920
rect 446 2915 447 2919
rect 451 2915 452 2919
rect 446 2914 452 2915
rect 520 2912 522 2930
rect 576 2920 578 2937
rect 712 2920 714 2937
rect 752 2936 754 2982
rect 760 2952 762 2982
rect 766 2977 772 2978
rect 766 2973 767 2977
rect 771 2973 772 2977
rect 766 2972 772 2973
rect 758 2951 764 2952
rect 758 2947 759 2951
rect 763 2947 764 2951
rect 758 2946 764 2947
rect 768 2943 770 2972
rect 848 2960 850 2982
rect 854 2977 860 2978
rect 854 2973 855 2977
rect 859 2973 860 2977
rect 854 2972 860 2973
rect 846 2959 852 2960
rect 846 2955 847 2959
rect 851 2955 852 2959
rect 846 2954 852 2955
rect 798 2943 804 2944
rect 856 2943 858 2972
rect 864 2960 866 3050
rect 878 3048 884 3049
rect 878 3044 879 3048
rect 883 3044 884 3048
rect 878 3043 884 3044
rect 880 3019 882 3043
rect 879 3018 883 3019
rect 879 3013 883 3014
rect 936 2988 938 3073
rect 952 3060 954 3078
rect 968 3068 970 3085
rect 1038 3083 1044 3084
rect 1038 3079 1039 3083
rect 1043 3079 1044 3083
rect 1038 3078 1044 3079
rect 966 3067 972 3068
rect 966 3063 967 3067
rect 971 3063 972 3067
rect 966 3062 972 3063
rect 1040 3060 1042 3078
rect 1056 3068 1058 3085
rect 1126 3083 1132 3084
rect 1126 3079 1127 3083
rect 1131 3079 1132 3083
rect 1126 3078 1132 3079
rect 1054 3067 1060 3068
rect 1054 3063 1055 3067
rect 1059 3063 1060 3067
rect 1054 3062 1060 3063
rect 1128 3060 1130 3078
rect 1136 3060 1138 3086
rect 1143 3085 1147 3086
rect 1199 3090 1203 3091
rect 1199 3085 1203 3086
rect 1319 3090 1323 3091
rect 1319 3085 1323 3086
rect 1767 3090 1771 3091
rect 1807 3089 1811 3090
rect 1831 3094 1835 3095
rect 1831 3089 1835 3090
rect 1767 3085 1771 3086
rect 1144 3068 1146 3085
rect 1768 3069 1770 3085
rect 1808 3073 1810 3089
rect 1806 3072 1812 3073
rect 1832 3072 1834 3089
rect 1896 3088 1898 3130
rect 1912 3108 1914 3130
rect 2006 3125 2012 3126
rect 2006 3121 2007 3125
rect 2011 3121 2012 3125
rect 2006 3120 2012 3121
rect 2206 3125 2212 3126
rect 2206 3121 2207 3125
rect 2211 3121 2212 3125
rect 2206 3120 2212 3121
rect 1910 3107 1916 3108
rect 1910 3103 1911 3107
rect 1915 3103 1916 3107
rect 1910 3102 1916 3103
rect 2008 3095 2010 3120
rect 2208 3095 2210 3120
rect 2272 3108 2274 3190
rect 2358 3188 2364 3189
rect 2358 3184 2359 3188
rect 2363 3184 2364 3188
rect 2358 3183 2364 3184
rect 2360 3167 2362 3183
rect 2480 3180 2482 3194
rect 2526 3188 2532 3189
rect 2526 3184 2527 3188
rect 2531 3184 2532 3188
rect 2526 3183 2532 3184
rect 2686 3188 2692 3189
rect 2686 3184 2687 3188
rect 2691 3184 2692 3188
rect 2686 3183 2692 3184
rect 2478 3179 2484 3180
rect 2478 3175 2479 3179
rect 2483 3175 2484 3179
rect 2478 3174 2484 3175
rect 2528 3167 2530 3183
rect 2688 3167 2690 3183
rect 2359 3166 2363 3167
rect 2359 3161 2363 3162
rect 2399 3166 2403 3167
rect 2399 3161 2403 3162
rect 2527 3166 2531 3167
rect 2527 3161 2531 3162
rect 2583 3166 2587 3167
rect 2583 3161 2587 3162
rect 2687 3166 2691 3167
rect 2687 3161 2691 3162
rect 2759 3166 2763 3167
rect 2759 3161 2763 3162
rect 2400 3145 2402 3161
rect 2584 3145 2586 3161
rect 2760 3145 2762 3161
rect 2398 3144 2404 3145
rect 2398 3140 2399 3144
rect 2403 3140 2404 3144
rect 2398 3139 2404 3140
rect 2582 3144 2588 3145
rect 2582 3140 2583 3144
rect 2587 3140 2588 3144
rect 2582 3139 2588 3140
rect 2758 3144 2764 3145
rect 2758 3140 2759 3144
rect 2763 3140 2764 3144
rect 2758 3139 2764 3140
rect 2832 3136 2834 3218
rect 2848 3208 2850 3225
rect 3008 3208 3010 3225
rect 3168 3208 3170 3225
rect 3264 3224 3266 3262
rect 3462 3256 3468 3257
rect 3462 3252 3463 3256
rect 3467 3252 3468 3256
rect 3462 3251 3468 3252
rect 3464 3231 3466 3251
rect 3335 3230 3339 3231
rect 3335 3225 3339 3226
rect 3463 3230 3467 3231
rect 3463 3225 3467 3226
rect 3262 3223 3268 3224
rect 3262 3219 3263 3223
rect 3267 3219 3268 3223
rect 3262 3218 3268 3219
rect 3302 3223 3308 3224
rect 3302 3219 3303 3223
rect 3307 3219 3308 3223
rect 3302 3218 3308 3219
rect 2846 3207 2852 3208
rect 2846 3203 2847 3207
rect 2851 3203 2852 3207
rect 2846 3202 2852 3203
rect 3006 3207 3012 3208
rect 3006 3203 3007 3207
rect 3011 3203 3012 3207
rect 3006 3202 3012 3203
rect 3166 3207 3172 3208
rect 3166 3203 3167 3207
rect 3171 3203 3172 3207
rect 3166 3202 3172 3203
rect 2966 3199 2972 3200
rect 2966 3195 2967 3199
rect 2971 3195 2972 3199
rect 2966 3194 2972 3195
rect 2846 3188 2852 3189
rect 2846 3184 2847 3188
rect 2851 3184 2852 3188
rect 2846 3183 2852 3184
rect 2848 3167 2850 3183
rect 2847 3166 2851 3167
rect 2847 3161 2851 3162
rect 2919 3166 2923 3167
rect 2919 3161 2923 3162
rect 2920 3145 2922 3161
rect 2918 3144 2924 3145
rect 2918 3140 2919 3144
rect 2923 3140 2924 3144
rect 2918 3139 2924 3140
rect 2278 3135 2284 3136
rect 2278 3131 2279 3135
rect 2283 3131 2284 3135
rect 2278 3130 2284 3131
rect 2286 3135 2292 3136
rect 2286 3131 2287 3135
rect 2291 3131 2292 3135
rect 2286 3130 2292 3131
rect 2742 3135 2748 3136
rect 2742 3131 2743 3135
rect 2747 3131 2748 3135
rect 2742 3130 2748 3131
rect 2830 3135 2836 3136
rect 2830 3131 2831 3135
rect 2835 3131 2836 3135
rect 2830 3130 2836 3131
rect 2280 3108 2282 3130
rect 2270 3107 2276 3108
rect 2270 3103 2271 3107
rect 2275 3103 2276 3107
rect 2270 3102 2276 3103
rect 2278 3107 2284 3108
rect 2278 3103 2279 3107
rect 2283 3103 2284 3107
rect 2278 3102 2284 3103
rect 2288 3100 2290 3130
rect 2398 3125 2404 3126
rect 2398 3121 2399 3125
rect 2403 3121 2404 3125
rect 2398 3120 2404 3121
rect 2582 3125 2588 3126
rect 2582 3121 2583 3125
rect 2587 3121 2588 3125
rect 2582 3120 2588 3121
rect 2286 3099 2292 3100
rect 2286 3095 2287 3099
rect 2291 3095 2292 3099
rect 2400 3095 2402 3120
rect 2584 3095 2586 3120
rect 2744 3108 2746 3130
rect 2758 3125 2764 3126
rect 2758 3121 2759 3125
rect 2763 3121 2764 3125
rect 2758 3120 2764 3121
rect 2918 3125 2924 3126
rect 2918 3121 2919 3125
rect 2923 3121 2924 3125
rect 2918 3120 2924 3121
rect 2742 3107 2748 3108
rect 2742 3103 2743 3107
rect 2747 3103 2748 3107
rect 2742 3102 2748 3103
rect 2760 3095 2762 3120
rect 2920 3095 2922 3120
rect 2968 3108 2970 3194
rect 3006 3188 3012 3189
rect 3006 3184 3007 3188
rect 3011 3184 3012 3188
rect 3006 3183 3012 3184
rect 3166 3188 3172 3189
rect 3166 3184 3167 3188
rect 3171 3184 3172 3188
rect 3166 3183 3172 3184
rect 3008 3167 3010 3183
rect 3168 3167 3170 3183
rect 3007 3166 3011 3167
rect 3007 3161 3011 3162
rect 3079 3166 3083 3167
rect 3079 3161 3083 3162
rect 3167 3166 3171 3167
rect 3167 3161 3171 3162
rect 3231 3166 3235 3167
rect 3231 3161 3235 3162
rect 3080 3145 3082 3161
rect 3232 3145 3234 3161
rect 3078 3144 3084 3145
rect 3078 3140 3079 3144
rect 3083 3140 3084 3144
rect 3078 3139 3084 3140
rect 3230 3144 3236 3145
rect 3230 3140 3231 3144
rect 3235 3140 3236 3144
rect 3230 3139 3236 3140
rect 3304 3136 3306 3218
rect 3336 3208 3338 3225
rect 3464 3209 3466 3225
rect 3462 3208 3468 3209
rect 3334 3207 3340 3208
rect 3334 3203 3335 3207
rect 3339 3203 3340 3207
rect 3462 3204 3463 3208
rect 3467 3204 3468 3208
rect 3462 3203 3468 3204
rect 3334 3202 3340 3203
rect 3406 3195 3412 3196
rect 3406 3191 3407 3195
rect 3411 3191 3412 3195
rect 3406 3190 3412 3191
rect 3462 3191 3468 3192
rect 3334 3188 3340 3189
rect 3334 3184 3335 3188
rect 3339 3184 3340 3188
rect 3334 3183 3340 3184
rect 3336 3167 3338 3183
rect 3335 3166 3339 3167
rect 3335 3161 3339 3162
rect 3367 3166 3371 3167
rect 3367 3161 3371 3162
rect 3368 3145 3370 3161
rect 3366 3144 3372 3145
rect 3366 3140 3367 3144
rect 3371 3140 3372 3144
rect 3366 3139 3372 3140
rect 2990 3135 2996 3136
rect 2990 3131 2991 3135
rect 2995 3131 2996 3135
rect 2990 3130 2996 3131
rect 3150 3135 3156 3136
rect 3150 3131 3151 3135
rect 3155 3131 3156 3135
rect 3150 3130 3156 3131
rect 3302 3135 3308 3136
rect 3302 3131 3303 3135
rect 3307 3131 3308 3135
rect 3302 3130 3308 3131
rect 2992 3108 2994 3130
rect 3078 3125 3084 3126
rect 3078 3121 3079 3125
rect 3083 3121 3084 3125
rect 3078 3120 3084 3121
rect 2966 3107 2972 3108
rect 2966 3103 2967 3107
rect 2971 3103 2972 3107
rect 2966 3102 2972 3103
rect 2990 3107 2996 3108
rect 2990 3103 2991 3107
rect 2995 3103 2996 3107
rect 2990 3102 2996 3103
rect 3080 3095 3082 3120
rect 3152 3108 3154 3130
rect 3230 3125 3236 3126
rect 3230 3121 3231 3125
rect 3235 3121 3236 3125
rect 3230 3120 3236 3121
rect 3366 3125 3372 3126
rect 3366 3121 3367 3125
rect 3371 3121 3372 3125
rect 3366 3120 3372 3121
rect 3150 3107 3156 3108
rect 3150 3103 3151 3107
rect 3155 3103 3156 3107
rect 3150 3102 3156 3103
rect 3232 3095 3234 3120
rect 3368 3095 3370 3120
rect 3408 3108 3410 3190
rect 3462 3187 3463 3191
rect 3467 3187 3468 3191
rect 3462 3186 3468 3187
rect 3464 3167 3466 3186
rect 3463 3166 3467 3167
rect 3463 3161 3467 3162
rect 3464 3142 3466 3161
rect 3462 3141 3468 3142
rect 3462 3137 3463 3141
rect 3467 3137 3468 3141
rect 3462 3136 3468 3137
rect 3430 3135 3436 3136
rect 3430 3131 3431 3135
rect 3435 3131 3436 3135
rect 3430 3130 3436 3131
rect 3406 3107 3412 3108
rect 3406 3103 3407 3107
rect 3411 3103 3412 3107
rect 3406 3102 3412 3103
rect 1959 3094 1963 3095
rect 1959 3089 1963 3090
rect 2007 3094 2011 3095
rect 2007 3089 2011 3090
rect 2119 3094 2123 3095
rect 2119 3089 2123 3090
rect 2207 3094 2211 3095
rect 2286 3094 2292 3095
rect 2295 3094 2299 3095
rect 2207 3089 2211 3090
rect 2295 3089 2299 3090
rect 2399 3094 2403 3095
rect 2399 3089 2403 3090
rect 2487 3094 2491 3095
rect 2487 3089 2491 3090
rect 2583 3094 2587 3095
rect 2583 3089 2587 3090
rect 2695 3094 2699 3095
rect 2695 3089 2699 3090
rect 2759 3094 2763 3095
rect 2759 3089 2763 3090
rect 2919 3094 2923 3095
rect 2919 3089 2923 3090
rect 3079 3094 3083 3095
rect 3079 3089 3083 3090
rect 3151 3094 3155 3095
rect 3151 3089 3155 3090
rect 3231 3094 3235 3095
rect 3231 3089 3235 3090
rect 3367 3094 3371 3095
rect 3367 3089 3371 3090
rect 1894 3087 1900 3088
rect 1894 3083 1895 3087
rect 1899 3083 1900 3087
rect 1894 3082 1900 3083
rect 1902 3087 1908 3088
rect 1902 3083 1903 3087
rect 1907 3083 1908 3087
rect 1902 3082 1908 3083
rect 1766 3068 1772 3069
rect 1142 3067 1148 3068
rect 1142 3063 1143 3067
rect 1147 3063 1148 3067
rect 1766 3064 1767 3068
rect 1771 3064 1772 3068
rect 1806 3068 1807 3072
rect 1811 3068 1812 3072
rect 1806 3067 1812 3068
rect 1830 3071 1836 3072
rect 1830 3067 1831 3071
rect 1835 3067 1836 3071
rect 1830 3066 1836 3067
rect 1904 3064 1906 3082
rect 1960 3072 1962 3089
rect 2030 3087 2036 3088
rect 2030 3083 2031 3087
rect 2035 3083 2036 3087
rect 2030 3082 2036 3083
rect 1958 3071 1964 3072
rect 1958 3067 1959 3071
rect 1963 3067 1964 3071
rect 1958 3066 1964 3067
rect 2032 3064 2034 3082
rect 2120 3072 2122 3089
rect 2190 3087 2196 3088
rect 2190 3083 2191 3087
rect 2195 3083 2196 3087
rect 2190 3082 2196 3083
rect 2118 3071 2124 3072
rect 2118 3067 2119 3071
rect 2123 3067 2124 3071
rect 2118 3066 2124 3067
rect 2192 3064 2194 3082
rect 2296 3072 2298 3089
rect 2488 3072 2490 3089
rect 2550 3087 2556 3088
rect 2550 3083 2551 3087
rect 2555 3083 2556 3087
rect 2550 3082 2556 3083
rect 2558 3087 2564 3088
rect 2558 3083 2559 3087
rect 2563 3083 2564 3087
rect 2558 3082 2564 3083
rect 2294 3071 2300 3072
rect 2294 3067 2295 3071
rect 2299 3067 2300 3071
rect 2294 3066 2300 3067
rect 2486 3071 2492 3072
rect 2486 3067 2487 3071
rect 2491 3067 2492 3071
rect 2486 3066 2492 3067
rect 1766 3063 1772 3064
rect 1902 3063 1908 3064
rect 1142 3062 1148 3063
rect 950 3059 956 3060
rect 950 3055 951 3059
rect 955 3055 956 3059
rect 950 3054 956 3055
rect 1038 3059 1044 3060
rect 1038 3055 1039 3059
rect 1043 3055 1044 3059
rect 1038 3054 1044 3055
rect 1126 3059 1132 3060
rect 1126 3055 1127 3059
rect 1131 3055 1132 3059
rect 1126 3054 1132 3055
rect 1134 3059 1140 3060
rect 1134 3055 1135 3059
rect 1139 3055 1140 3059
rect 1902 3059 1903 3063
rect 1907 3059 1908 3063
rect 1902 3058 1908 3059
rect 2030 3063 2036 3064
rect 2030 3059 2031 3063
rect 2035 3059 2036 3063
rect 2030 3058 2036 3059
rect 2190 3063 2196 3064
rect 2190 3059 2191 3063
rect 2195 3059 2196 3063
rect 2190 3058 2196 3059
rect 1134 3054 1140 3055
rect 1806 3055 1812 3056
rect 1766 3051 1772 3052
rect 966 3048 972 3049
rect 966 3044 967 3048
rect 971 3044 972 3048
rect 966 3043 972 3044
rect 1054 3048 1060 3049
rect 1054 3044 1055 3048
rect 1059 3044 1060 3048
rect 1054 3043 1060 3044
rect 1142 3048 1148 3049
rect 1142 3044 1143 3048
rect 1147 3044 1148 3048
rect 1766 3047 1767 3051
rect 1771 3047 1772 3051
rect 1806 3051 1807 3055
rect 1811 3051 1812 3055
rect 2182 3055 2188 3056
rect 1806 3050 1812 3051
rect 1830 3052 1836 3053
rect 1766 3046 1772 3047
rect 1142 3043 1148 3044
rect 968 3019 970 3043
rect 1056 3019 1058 3043
rect 1144 3019 1146 3043
rect 1768 3019 1770 3046
rect 943 3018 947 3019
rect 943 3013 947 3014
rect 967 3018 971 3019
rect 967 3013 971 3014
rect 1031 3018 1035 3019
rect 1031 3013 1035 3014
rect 1055 3018 1059 3019
rect 1055 3013 1059 3014
rect 1119 3018 1123 3019
rect 1119 3013 1123 3014
rect 1143 3018 1147 3019
rect 1143 3013 1147 3014
rect 1207 3018 1211 3019
rect 1207 3013 1211 3014
rect 1295 3018 1299 3019
rect 1295 3013 1299 3014
rect 1767 3018 1771 3019
rect 1808 3015 1810 3050
rect 1830 3048 1831 3052
rect 1835 3048 1836 3052
rect 1830 3047 1836 3048
rect 1958 3052 1964 3053
rect 1958 3048 1959 3052
rect 1963 3048 1964 3052
rect 1958 3047 1964 3048
rect 2118 3052 2124 3053
rect 2118 3048 2119 3052
rect 2123 3048 2124 3052
rect 2182 3051 2183 3055
rect 2187 3051 2188 3055
rect 2182 3050 2188 3051
rect 2294 3052 2300 3053
rect 2118 3047 2124 3048
rect 1832 3015 1834 3047
rect 1960 3015 1962 3047
rect 2120 3015 2122 3047
rect 1767 3013 1771 3014
rect 1807 3014 1811 3015
rect 944 2997 946 3013
rect 1032 2997 1034 3013
rect 1120 2997 1122 3013
rect 1208 2997 1210 3013
rect 1296 2997 1298 3013
rect 942 2996 948 2997
rect 942 2992 943 2996
rect 947 2992 948 2996
rect 942 2991 948 2992
rect 1030 2996 1036 2997
rect 1030 2992 1031 2996
rect 1035 2992 1036 2996
rect 1030 2991 1036 2992
rect 1118 2996 1124 2997
rect 1118 2992 1119 2996
rect 1123 2992 1124 2996
rect 1118 2991 1124 2992
rect 1206 2996 1212 2997
rect 1206 2992 1207 2996
rect 1211 2992 1212 2996
rect 1206 2991 1212 2992
rect 1294 2996 1300 2997
rect 1294 2992 1295 2996
rect 1299 2992 1300 2996
rect 1768 2994 1770 3013
rect 1807 3009 1811 3010
rect 1831 3014 1835 3015
rect 1831 3009 1835 3010
rect 1919 3014 1923 3015
rect 1919 3009 1923 3010
rect 1959 3014 1963 3015
rect 1959 3009 1963 3010
rect 2031 3014 2035 3015
rect 2031 3009 2035 3010
rect 2119 3014 2123 3015
rect 2119 3009 2123 3010
rect 2143 3014 2147 3015
rect 2143 3009 2147 3010
rect 1294 2991 1300 2992
rect 1766 2993 1772 2994
rect 1766 2989 1767 2993
rect 1771 2989 1772 2993
rect 1808 2990 1810 3009
rect 1832 2993 1834 3009
rect 1920 2993 1922 3009
rect 2032 2993 2034 3009
rect 2144 2993 2146 3009
rect 1830 2992 1836 2993
rect 1766 2988 1772 2989
rect 1806 2989 1812 2990
rect 934 2987 940 2988
rect 934 2983 935 2987
rect 939 2983 940 2987
rect 934 2982 940 2983
rect 1022 2987 1028 2988
rect 1022 2983 1023 2987
rect 1027 2983 1028 2987
rect 1022 2982 1028 2983
rect 1190 2987 1196 2988
rect 1190 2983 1191 2987
rect 1195 2983 1196 2987
rect 1190 2982 1196 2983
rect 1278 2987 1284 2988
rect 1278 2983 1279 2987
rect 1283 2983 1284 2987
rect 1278 2982 1284 2983
rect 1286 2987 1292 2988
rect 1286 2983 1287 2987
rect 1291 2983 1292 2987
rect 1806 2985 1807 2989
rect 1811 2985 1812 2989
rect 1830 2988 1831 2992
rect 1835 2988 1836 2992
rect 1830 2987 1836 2988
rect 1918 2992 1924 2993
rect 1918 2988 1919 2992
rect 1923 2988 1924 2992
rect 1918 2987 1924 2988
rect 2030 2992 2036 2993
rect 2030 2988 2031 2992
rect 2035 2988 2036 2992
rect 2030 2987 2036 2988
rect 2142 2992 2148 2993
rect 2142 2988 2143 2992
rect 2147 2988 2148 2992
rect 2142 2987 2148 2988
rect 1806 2984 1812 2985
rect 1286 2982 1292 2983
rect 1894 2983 1900 2984
rect 942 2977 948 2978
rect 942 2973 943 2977
rect 947 2973 948 2977
rect 942 2972 948 2973
rect 862 2959 868 2960
rect 862 2955 863 2959
rect 867 2955 868 2959
rect 862 2954 868 2955
rect 944 2943 946 2972
rect 1024 2960 1026 2982
rect 1030 2977 1036 2978
rect 1030 2973 1031 2977
rect 1035 2973 1036 2977
rect 1030 2972 1036 2973
rect 1118 2977 1124 2978
rect 1118 2973 1119 2977
rect 1123 2973 1124 2977
rect 1118 2972 1124 2973
rect 1022 2959 1028 2960
rect 1022 2955 1023 2959
rect 1027 2955 1028 2959
rect 1022 2954 1028 2955
rect 1032 2943 1034 2972
rect 1120 2943 1122 2972
rect 1192 2960 1194 2982
rect 1206 2977 1212 2978
rect 1206 2973 1207 2977
rect 1211 2973 1212 2977
rect 1206 2972 1212 2973
rect 1166 2959 1172 2960
rect 1166 2955 1167 2959
rect 1171 2955 1172 2959
rect 1166 2954 1172 2955
rect 1190 2959 1196 2960
rect 1190 2955 1191 2959
rect 1195 2955 1196 2959
rect 1190 2954 1196 2955
rect 767 2942 771 2943
rect 798 2939 799 2943
rect 803 2939 804 2943
rect 798 2938 804 2939
rect 847 2942 851 2943
rect 767 2937 771 2938
rect 750 2935 756 2936
rect 750 2931 751 2935
rect 755 2931 756 2935
rect 750 2930 756 2931
rect 782 2935 788 2936
rect 782 2931 783 2935
rect 787 2931 788 2935
rect 782 2930 788 2931
rect 574 2919 580 2920
rect 574 2915 575 2919
rect 579 2915 580 2919
rect 574 2914 580 2915
rect 710 2919 716 2920
rect 710 2915 711 2919
rect 715 2915 716 2919
rect 710 2914 716 2915
rect 784 2912 786 2930
rect 800 2912 802 2938
rect 847 2937 851 2938
rect 855 2942 859 2943
rect 855 2937 859 2938
rect 943 2942 947 2943
rect 943 2937 947 2938
rect 975 2942 979 2943
rect 975 2937 979 2938
rect 1031 2942 1035 2943
rect 1031 2937 1035 2938
rect 1103 2942 1107 2943
rect 1103 2937 1107 2938
rect 1119 2942 1123 2943
rect 1119 2937 1123 2938
rect 848 2920 850 2937
rect 976 2920 978 2937
rect 1104 2920 1106 2937
rect 846 2919 852 2920
rect 846 2915 847 2919
rect 851 2915 852 2919
rect 846 2914 852 2915
rect 974 2919 980 2920
rect 974 2915 975 2919
rect 979 2915 980 2919
rect 974 2914 980 2915
rect 1102 2919 1108 2920
rect 1102 2915 1103 2919
rect 1107 2915 1108 2919
rect 1168 2916 1170 2954
rect 1182 2943 1188 2944
rect 1208 2943 1210 2972
rect 1280 2960 1282 2982
rect 1278 2959 1284 2960
rect 1278 2955 1279 2959
rect 1283 2955 1284 2959
rect 1278 2954 1284 2955
rect 1288 2952 1290 2982
rect 1894 2979 1895 2983
rect 1899 2979 1900 2983
rect 1894 2978 1900 2979
rect 1910 2983 1916 2984
rect 1910 2979 1911 2983
rect 1915 2979 1916 2983
rect 1910 2978 1916 2979
rect 1294 2977 1300 2978
rect 1294 2973 1295 2977
rect 1299 2973 1300 2977
rect 1294 2972 1300 2973
rect 1766 2976 1772 2977
rect 1766 2972 1767 2976
rect 1771 2972 1772 2976
rect 1830 2973 1836 2974
rect 1286 2951 1292 2952
rect 1286 2947 1287 2951
rect 1291 2947 1292 2951
rect 1286 2946 1292 2947
rect 1296 2943 1298 2972
rect 1766 2971 1772 2972
rect 1806 2972 1812 2973
rect 1768 2943 1770 2971
rect 1806 2968 1807 2972
rect 1811 2968 1812 2972
rect 1830 2969 1831 2973
rect 1835 2969 1836 2973
rect 1830 2968 1836 2969
rect 1806 2967 1812 2968
rect 1182 2939 1183 2943
rect 1187 2939 1188 2943
rect 1182 2938 1188 2939
rect 1207 2942 1211 2943
rect 1102 2914 1108 2915
rect 1166 2915 1172 2916
rect 398 2911 404 2912
rect 398 2907 399 2911
rect 403 2907 404 2911
rect 398 2906 404 2907
rect 518 2911 524 2912
rect 518 2907 519 2911
rect 523 2907 524 2911
rect 518 2906 524 2907
rect 782 2911 788 2912
rect 782 2907 783 2911
rect 787 2907 788 2911
rect 782 2906 788 2907
rect 798 2911 804 2912
rect 798 2907 799 2911
rect 803 2907 804 2911
rect 1166 2911 1167 2915
rect 1171 2911 1172 2915
rect 1184 2912 1186 2938
rect 1207 2937 1211 2938
rect 1231 2942 1235 2943
rect 1231 2937 1235 2938
rect 1295 2942 1299 2943
rect 1295 2937 1299 2938
rect 1359 2942 1363 2943
rect 1359 2937 1363 2938
rect 1495 2942 1499 2943
rect 1495 2937 1499 2938
rect 1767 2942 1771 2943
rect 1808 2939 1810 2967
rect 1832 2939 1834 2968
rect 1767 2937 1771 2938
rect 1807 2938 1811 2939
rect 1232 2920 1234 2937
rect 1310 2935 1316 2936
rect 1310 2931 1311 2935
rect 1315 2931 1316 2935
rect 1310 2930 1316 2931
rect 1230 2919 1236 2920
rect 1230 2915 1231 2919
rect 1235 2915 1236 2919
rect 1230 2914 1236 2915
rect 1312 2912 1314 2930
rect 1360 2920 1362 2937
rect 1496 2920 1498 2937
rect 1558 2935 1564 2936
rect 1558 2931 1559 2935
rect 1563 2931 1564 2935
rect 1558 2930 1564 2931
rect 1358 2919 1364 2920
rect 1358 2915 1359 2919
rect 1363 2915 1364 2919
rect 1358 2914 1364 2915
rect 1494 2919 1500 2920
rect 1494 2915 1495 2919
rect 1499 2915 1500 2919
rect 1494 2914 1500 2915
rect 1166 2910 1172 2911
rect 1182 2911 1188 2912
rect 798 2906 804 2907
rect 1182 2907 1183 2911
rect 1187 2907 1188 2911
rect 1182 2906 1188 2907
rect 1310 2911 1316 2912
rect 1310 2907 1311 2911
rect 1315 2907 1316 2911
rect 1310 2906 1316 2907
rect 110 2903 116 2904
rect 110 2899 111 2903
rect 115 2899 116 2903
rect 638 2903 644 2904
rect 110 2898 116 2899
rect 326 2900 332 2901
rect 112 2871 114 2898
rect 326 2896 327 2900
rect 331 2896 332 2900
rect 326 2895 332 2896
rect 446 2900 452 2901
rect 446 2896 447 2900
rect 451 2896 452 2900
rect 446 2895 452 2896
rect 574 2900 580 2901
rect 574 2896 575 2900
rect 579 2896 580 2900
rect 638 2899 639 2903
rect 643 2899 644 2903
rect 638 2898 644 2899
rect 710 2900 716 2901
rect 574 2895 580 2896
rect 328 2871 330 2895
rect 448 2871 450 2895
rect 576 2871 578 2895
rect 111 2870 115 2871
rect 111 2865 115 2866
rect 135 2870 139 2871
rect 135 2865 139 2866
rect 255 2870 259 2871
rect 255 2865 259 2866
rect 327 2870 331 2871
rect 327 2865 331 2866
rect 415 2870 419 2871
rect 415 2865 419 2866
rect 447 2870 451 2871
rect 447 2865 451 2866
rect 575 2870 579 2871
rect 575 2865 579 2866
rect 112 2846 114 2865
rect 136 2849 138 2865
rect 256 2849 258 2865
rect 416 2849 418 2865
rect 576 2849 578 2865
rect 134 2848 140 2849
rect 110 2845 116 2846
rect 110 2841 111 2845
rect 115 2841 116 2845
rect 134 2844 135 2848
rect 139 2844 140 2848
rect 134 2843 140 2844
rect 254 2848 260 2849
rect 254 2844 255 2848
rect 259 2844 260 2848
rect 254 2843 260 2844
rect 414 2848 420 2849
rect 414 2844 415 2848
rect 419 2844 420 2848
rect 414 2843 420 2844
rect 574 2848 580 2849
rect 574 2844 575 2848
rect 579 2844 580 2848
rect 574 2843 580 2844
rect 110 2840 116 2841
rect 198 2839 204 2840
rect 198 2835 199 2839
rect 203 2835 204 2839
rect 198 2834 204 2835
rect 214 2839 220 2840
rect 214 2835 215 2839
rect 219 2835 220 2839
rect 214 2834 220 2835
rect 334 2839 340 2840
rect 334 2835 335 2839
rect 339 2835 340 2839
rect 334 2834 340 2835
rect 134 2829 140 2830
rect 110 2828 116 2829
rect 110 2824 111 2828
rect 115 2824 116 2828
rect 134 2825 135 2829
rect 139 2825 140 2829
rect 134 2824 140 2825
rect 110 2823 116 2824
rect 112 2795 114 2823
rect 136 2795 138 2824
rect 111 2794 115 2795
rect 111 2789 115 2790
rect 135 2794 139 2795
rect 135 2789 139 2790
rect 112 2773 114 2789
rect 110 2772 116 2773
rect 136 2772 138 2789
rect 200 2788 202 2834
rect 216 2812 218 2834
rect 254 2829 260 2830
rect 254 2825 255 2829
rect 259 2825 260 2829
rect 254 2824 260 2825
rect 214 2811 220 2812
rect 214 2807 215 2811
rect 219 2807 220 2811
rect 214 2806 220 2807
rect 256 2795 258 2824
rect 336 2812 338 2834
rect 414 2829 420 2830
rect 414 2825 415 2829
rect 419 2825 420 2829
rect 414 2824 420 2825
rect 574 2829 580 2830
rect 574 2825 575 2829
rect 579 2825 580 2829
rect 574 2824 580 2825
rect 334 2811 340 2812
rect 334 2807 335 2811
rect 339 2807 340 2811
rect 334 2806 340 2807
rect 416 2795 418 2824
rect 576 2795 578 2824
rect 640 2812 642 2898
rect 710 2896 711 2900
rect 715 2896 716 2900
rect 710 2895 716 2896
rect 846 2900 852 2901
rect 846 2896 847 2900
rect 851 2896 852 2900
rect 846 2895 852 2896
rect 974 2900 980 2901
rect 974 2896 975 2900
rect 979 2896 980 2900
rect 974 2895 980 2896
rect 1102 2900 1108 2901
rect 1102 2896 1103 2900
rect 1107 2896 1108 2900
rect 1102 2895 1108 2896
rect 1230 2900 1236 2901
rect 1230 2896 1231 2900
rect 1235 2896 1236 2900
rect 1230 2895 1236 2896
rect 1358 2900 1364 2901
rect 1358 2896 1359 2900
rect 1363 2896 1364 2900
rect 1358 2895 1364 2896
rect 1494 2900 1500 2901
rect 1494 2896 1495 2900
rect 1499 2896 1500 2900
rect 1494 2895 1500 2896
rect 712 2871 714 2895
rect 848 2871 850 2895
rect 976 2871 978 2895
rect 1104 2871 1106 2895
rect 1232 2871 1234 2895
rect 1360 2871 1362 2895
rect 1496 2871 1498 2895
rect 711 2870 715 2871
rect 711 2865 715 2866
rect 735 2870 739 2871
rect 735 2865 739 2866
rect 847 2870 851 2871
rect 847 2865 851 2866
rect 895 2870 899 2871
rect 895 2865 899 2866
rect 975 2870 979 2871
rect 975 2865 979 2866
rect 1047 2870 1051 2871
rect 1047 2865 1051 2866
rect 1103 2870 1107 2871
rect 1103 2865 1107 2866
rect 1191 2870 1195 2871
rect 1191 2865 1195 2866
rect 1231 2870 1235 2871
rect 1231 2865 1235 2866
rect 1343 2870 1347 2871
rect 1343 2865 1347 2866
rect 1359 2870 1363 2871
rect 1359 2865 1363 2866
rect 1495 2870 1499 2871
rect 1495 2865 1499 2866
rect 736 2849 738 2865
rect 896 2849 898 2865
rect 1048 2849 1050 2865
rect 1192 2849 1194 2865
rect 1344 2849 1346 2865
rect 1496 2849 1498 2865
rect 734 2848 740 2849
rect 734 2844 735 2848
rect 739 2844 740 2848
rect 734 2843 740 2844
rect 894 2848 900 2849
rect 894 2844 895 2848
rect 899 2844 900 2848
rect 894 2843 900 2844
rect 1046 2848 1052 2849
rect 1046 2844 1047 2848
rect 1051 2844 1052 2848
rect 1046 2843 1052 2844
rect 1190 2848 1196 2849
rect 1190 2844 1191 2848
rect 1195 2844 1196 2848
rect 1190 2843 1196 2844
rect 1342 2848 1348 2849
rect 1342 2844 1343 2848
rect 1347 2844 1348 2848
rect 1342 2843 1348 2844
rect 1494 2848 1500 2849
rect 1494 2844 1495 2848
rect 1499 2844 1500 2848
rect 1494 2843 1500 2844
rect 1560 2840 1562 2930
rect 1768 2921 1770 2937
rect 1807 2933 1811 2934
rect 1831 2938 1835 2939
rect 1831 2933 1835 2934
rect 1766 2920 1772 2921
rect 1766 2916 1767 2920
rect 1771 2916 1772 2920
rect 1808 2917 1810 2933
rect 1766 2915 1772 2916
rect 1806 2916 1812 2917
rect 1832 2916 1834 2933
rect 1896 2932 1898 2978
rect 1912 2956 1914 2978
rect 1918 2973 1924 2974
rect 1918 2969 1919 2973
rect 1923 2969 1924 2973
rect 1918 2968 1924 2969
rect 2030 2973 2036 2974
rect 2030 2969 2031 2973
rect 2035 2969 2036 2973
rect 2030 2968 2036 2969
rect 2142 2973 2148 2974
rect 2142 2969 2143 2973
rect 2147 2969 2148 2973
rect 2142 2968 2148 2969
rect 1910 2955 1916 2956
rect 1910 2951 1911 2955
rect 1915 2951 1916 2955
rect 1910 2950 1916 2951
rect 1920 2939 1922 2968
rect 2032 2939 2034 2968
rect 2144 2939 2146 2968
rect 2184 2956 2186 3050
rect 2294 3048 2295 3052
rect 2299 3048 2300 3052
rect 2294 3047 2300 3048
rect 2486 3052 2492 3053
rect 2486 3048 2487 3052
rect 2491 3048 2492 3052
rect 2486 3047 2492 3048
rect 2296 3015 2298 3047
rect 2488 3015 2490 3047
rect 2247 3014 2251 3015
rect 2247 3009 2251 3010
rect 2295 3014 2299 3015
rect 2295 3009 2299 3010
rect 2359 3014 2363 3015
rect 2359 3009 2363 3010
rect 2479 3014 2483 3015
rect 2479 3009 2483 3010
rect 2487 3014 2491 3015
rect 2487 3009 2491 3010
rect 2248 2993 2250 3009
rect 2360 2993 2362 3009
rect 2480 2993 2482 3009
rect 2552 3000 2554 3082
rect 2560 3064 2562 3082
rect 2696 3072 2698 3089
rect 2766 3087 2772 3088
rect 2766 3083 2767 3087
rect 2771 3083 2772 3087
rect 2766 3082 2772 3083
rect 2694 3071 2700 3072
rect 2694 3067 2695 3071
rect 2699 3067 2700 3071
rect 2694 3066 2700 3067
rect 2768 3064 2770 3082
rect 2920 3072 2922 3089
rect 2990 3087 2996 3088
rect 2990 3083 2991 3087
rect 2995 3083 2996 3087
rect 2990 3082 2996 3083
rect 2918 3071 2924 3072
rect 2918 3067 2919 3071
rect 2923 3067 2924 3071
rect 2918 3066 2924 3067
rect 2992 3064 2994 3082
rect 3152 3072 3154 3089
rect 3368 3072 3370 3089
rect 3432 3088 3434 3130
rect 3462 3124 3468 3125
rect 3462 3120 3463 3124
rect 3467 3120 3468 3124
rect 3462 3119 3468 3120
rect 3464 3095 3466 3119
rect 3463 3094 3467 3095
rect 3463 3089 3467 3090
rect 3430 3087 3436 3088
rect 3430 3083 3431 3087
rect 3435 3083 3436 3087
rect 3430 3082 3436 3083
rect 3464 3073 3466 3089
rect 3462 3072 3468 3073
rect 3150 3071 3156 3072
rect 3150 3067 3151 3071
rect 3155 3067 3156 3071
rect 3150 3066 3156 3067
rect 3366 3071 3372 3072
rect 3366 3067 3367 3071
rect 3371 3067 3372 3071
rect 3462 3068 3463 3072
rect 3467 3068 3468 3072
rect 3462 3067 3468 3068
rect 3366 3066 3372 3067
rect 2558 3063 2564 3064
rect 2558 3059 2559 3063
rect 2563 3059 2564 3063
rect 2558 3058 2564 3059
rect 2766 3063 2772 3064
rect 2766 3059 2767 3063
rect 2771 3059 2772 3063
rect 2766 3058 2772 3059
rect 2990 3063 2996 3064
rect 2990 3059 2991 3063
rect 2995 3059 2996 3063
rect 2990 3058 2996 3059
rect 3430 3055 3436 3056
rect 2694 3052 2700 3053
rect 2694 3048 2695 3052
rect 2699 3048 2700 3052
rect 2694 3047 2700 3048
rect 2918 3052 2924 3053
rect 2918 3048 2919 3052
rect 2923 3048 2924 3052
rect 2918 3047 2924 3048
rect 3150 3052 3156 3053
rect 3150 3048 3151 3052
rect 3155 3048 3156 3052
rect 3150 3047 3156 3048
rect 3366 3052 3372 3053
rect 3366 3048 3367 3052
rect 3371 3048 3372 3052
rect 3430 3051 3431 3055
rect 3435 3051 3436 3055
rect 3430 3050 3436 3051
rect 3462 3055 3468 3056
rect 3462 3051 3463 3055
rect 3467 3051 3468 3055
rect 3462 3050 3468 3051
rect 3366 3047 3372 3048
rect 2696 3015 2698 3047
rect 2920 3015 2922 3047
rect 3152 3015 3154 3047
rect 3368 3015 3370 3047
rect 2623 3014 2627 3015
rect 2623 3009 2627 3010
rect 2695 3014 2699 3015
rect 2695 3009 2699 3010
rect 2791 3014 2795 3015
rect 2791 3009 2795 3010
rect 2919 3014 2923 3015
rect 2919 3009 2923 3010
rect 2983 3014 2987 3015
rect 2983 3009 2987 3010
rect 3151 3014 3155 3015
rect 3151 3009 3155 3010
rect 3183 3014 3187 3015
rect 3183 3009 3187 3010
rect 3367 3014 3371 3015
rect 3367 3009 3371 3010
rect 2550 2999 2556 3000
rect 2550 2995 2551 2999
rect 2555 2995 2556 2999
rect 2550 2994 2556 2995
rect 2624 2993 2626 3009
rect 2792 2993 2794 3009
rect 2984 2993 2986 3009
rect 3184 2993 3186 3009
rect 3368 2993 3370 3009
rect 2246 2992 2252 2993
rect 2246 2988 2247 2992
rect 2251 2988 2252 2992
rect 2246 2987 2252 2988
rect 2358 2992 2364 2993
rect 2358 2988 2359 2992
rect 2363 2988 2364 2992
rect 2358 2987 2364 2988
rect 2478 2992 2484 2993
rect 2478 2988 2479 2992
rect 2483 2988 2484 2992
rect 2478 2987 2484 2988
rect 2622 2992 2628 2993
rect 2622 2988 2623 2992
rect 2627 2988 2628 2992
rect 2622 2987 2628 2988
rect 2790 2992 2796 2993
rect 2790 2988 2791 2992
rect 2795 2988 2796 2992
rect 2790 2987 2796 2988
rect 2982 2992 2988 2993
rect 2982 2988 2983 2992
rect 2987 2988 2988 2992
rect 2982 2987 2988 2988
rect 3182 2992 3188 2993
rect 3182 2988 3183 2992
rect 3187 2988 3188 2992
rect 3182 2987 3188 2988
rect 3366 2992 3372 2993
rect 3366 2988 3367 2992
rect 3371 2988 3372 2992
rect 3366 2987 3372 2988
rect 2214 2983 2220 2984
rect 2214 2979 2215 2983
rect 2219 2979 2220 2983
rect 2214 2978 2220 2979
rect 2318 2983 2324 2984
rect 2318 2979 2319 2983
rect 2323 2979 2324 2983
rect 2318 2978 2324 2979
rect 2430 2983 2436 2984
rect 2430 2979 2431 2983
rect 2435 2979 2436 2983
rect 2430 2978 2436 2979
rect 2550 2983 2556 2984
rect 2550 2979 2551 2983
rect 2555 2979 2556 2983
rect 2550 2978 2556 2979
rect 2694 2983 2700 2984
rect 2694 2979 2695 2983
rect 2699 2979 2700 2983
rect 2694 2978 2700 2979
rect 2862 2983 2868 2984
rect 2862 2979 2863 2983
rect 2867 2979 2868 2983
rect 2862 2978 2868 2979
rect 3054 2983 3060 2984
rect 3054 2979 3055 2983
rect 3059 2979 3060 2983
rect 3054 2978 3060 2979
rect 2216 2956 2218 2978
rect 2246 2973 2252 2974
rect 2246 2969 2247 2973
rect 2251 2969 2252 2973
rect 2246 2968 2252 2969
rect 2182 2955 2188 2956
rect 2182 2951 2183 2955
rect 2187 2951 2188 2955
rect 2182 2950 2188 2951
rect 2194 2955 2200 2956
rect 2194 2951 2195 2955
rect 2199 2951 2200 2955
rect 2194 2950 2200 2951
rect 2214 2955 2220 2956
rect 2214 2951 2215 2955
rect 2219 2951 2220 2955
rect 2214 2950 2220 2951
rect 1919 2938 1923 2939
rect 1919 2933 1923 2934
rect 2015 2938 2019 2939
rect 2015 2933 2019 2934
rect 2031 2938 2035 2939
rect 2031 2933 2035 2934
rect 2143 2938 2147 2939
rect 2143 2933 2147 2934
rect 1894 2931 1900 2932
rect 1894 2927 1895 2931
rect 1899 2927 1900 2931
rect 1894 2926 1900 2927
rect 1902 2931 1908 2932
rect 1902 2927 1903 2931
rect 1907 2927 1908 2931
rect 1902 2926 1908 2927
rect 1806 2912 1807 2916
rect 1811 2912 1812 2916
rect 1806 2911 1812 2912
rect 1830 2915 1836 2916
rect 1830 2911 1831 2915
rect 1835 2911 1836 2915
rect 1830 2910 1836 2911
rect 1904 2908 1906 2926
rect 2016 2916 2018 2933
rect 2014 2915 2020 2916
rect 2014 2911 2015 2915
rect 2019 2911 2020 2915
rect 2014 2910 2020 2911
rect 2196 2908 2198 2950
rect 2248 2939 2250 2968
rect 2320 2956 2322 2978
rect 2358 2973 2364 2974
rect 2358 2969 2359 2973
rect 2363 2969 2364 2973
rect 2358 2968 2364 2969
rect 2318 2955 2324 2956
rect 2318 2951 2319 2955
rect 2323 2951 2324 2955
rect 2318 2950 2324 2951
rect 2360 2939 2362 2968
rect 2432 2956 2434 2978
rect 2478 2973 2484 2974
rect 2478 2969 2479 2973
rect 2483 2969 2484 2973
rect 2478 2968 2484 2969
rect 2430 2955 2436 2956
rect 2430 2951 2431 2955
rect 2435 2951 2436 2955
rect 2430 2950 2436 2951
rect 2480 2939 2482 2968
rect 2552 2956 2554 2978
rect 2622 2973 2628 2974
rect 2622 2969 2623 2973
rect 2627 2969 2628 2973
rect 2622 2968 2628 2969
rect 2550 2955 2556 2956
rect 2550 2951 2551 2955
rect 2555 2951 2556 2955
rect 2550 2950 2556 2951
rect 2624 2939 2626 2968
rect 2696 2956 2698 2978
rect 2790 2973 2796 2974
rect 2790 2969 2791 2973
rect 2795 2969 2796 2973
rect 2790 2968 2796 2969
rect 2694 2955 2700 2956
rect 2694 2951 2695 2955
rect 2699 2951 2700 2955
rect 2694 2950 2700 2951
rect 2792 2939 2794 2968
rect 2864 2956 2866 2978
rect 2982 2973 2988 2974
rect 2982 2969 2983 2973
rect 2987 2969 2988 2973
rect 2982 2968 2988 2969
rect 2862 2955 2868 2956
rect 2862 2951 2863 2955
rect 2867 2951 2868 2955
rect 2862 2950 2868 2951
rect 2984 2939 2986 2968
rect 3056 2956 3058 2978
rect 3182 2973 3188 2974
rect 3182 2969 3183 2973
rect 3187 2969 3188 2973
rect 3182 2968 3188 2969
rect 3366 2973 3372 2974
rect 3366 2969 3367 2973
rect 3371 2969 3372 2973
rect 3366 2968 3372 2969
rect 3054 2955 3060 2956
rect 3054 2951 3055 2955
rect 3059 2951 3060 2955
rect 3054 2950 3060 2951
rect 3184 2939 3186 2968
rect 3368 2939 3370 2968
rect 3432 2956 3434 3050
rect 3464 3015 3466 3050
rect 3463 3014 3467 3015
rect 3463 3009 3467 3010
rect 3464 2990 3466 3009
rect 3462 2989 3468 2990
rect 3462 2985 3463 2989
rect 3467 2985 3468 2989
rect 3462 2984 3468 2985
rect 3438 2983 3444 2984
rect 3438 2979 3439 2983
rect 3443 2979 3444 2983
rect 3438 2978 3444 2979
rect 3430 2955 3436 2956
rect 3430 2951 3431 2955
rect 3435 2951 3436 2955
rect 3430 2950 3436 2951
rect 2215 2938 2219 2939
rect 2215 2933 2219 2934
rect 2247 2938 2251 2939
rect 2247 2933 2251 2934
rect 2359 2938 2363 2939
rect 2359 2933 2363 2934
rect 2407 2938 2411 2939
rect 2407 2933 2411 2934
rect 2479 2938 2483 2939
rect 2479 2933 2483 2934
rect 2591 2938 2595 2939
rect 2591 2933 2595 2934
rect 2623 2938 2627 2939
rect 2623 2933 2627 2934
rect 2759 2938 2763 2939
rect 2759 2933 2763 2934
rect 2791 2938 2795 2939
rect 2791 2933 2795 2934
rect 2911 2938 2915 2939
rect 2911 2933 2915 2934
rect 2983 2938 2987 2939
rect 2983 2933 2987 2934
rect 3063 2938 3067 2939
rect 3063 2933 3067 2934
rect 3183 2938 3187 2939
rect 3183 2933 3187 2934
rect 3207 2938 3211 2939
rect 3207 2933 3211 2934
rect 3359 2938 3363 2939
rect 3359 2933 3363 2934
rect 3367 2938 3371 2939
rect 3367 2933 3371 2934
rect 2216 2916 2218 2933
rect 2294 2931 2300 2932
rect 2294 2927 2295 2931
rect 2299 2927 2300 2931
rect 2294 2926 2300 2927
rect 2214 2915 2220 2916
rect 2214 2911 2215 2915
rect 2219 2911 2220 2915
rect 2214 2910 2220 2911
rect 2296 2908 2298 2926
rect 2408 2916 2410 2933
rect 2486 2931 2492 2932
rect 2486 2927 2487 2931
rect 2491 2927 2492 2931
rect 2486 2926 2492 2927
rect 2406 2915 2412 2916
rect 2406 2911 2407 2915
rect 2411 2911 2412 2915
rect 2406 2910 2412 2911
rect 2488 2908 2490 2926
rect 2592 2916 2594 2933
rect 2638 2931 2644 2932
rect 2638 2927 2639 2931
rect 2643 2927 2644 2931
rect 2638 2926 2644 2927
rect 2590 2915 2596 2916
rect 2590 2911 2591 2915
rect 2595 2911 2596 2915
rect 2590 2910 2596 2911
rect 1902 2907 1908 2908
rect 1766 2903 1772 2904
rect 1766 2899 1767 2903
rect 1771 2899 1772 2903
rect 1902 2903 1903 2907
rect 1907 2903 1908 2907
rect 2194 2907 2200 2908
rect 1902 2902 1908 2903
rect 2086 2903 2092 2904
rect 1766 2898 1772 2899
rect 1806 2899 1812 2900
rect 1768 2871 1770 2898
rect 1806 2895 1807 2899
rect 1811 2895 1812 2899
rect 2086 2899 2087 2903
rect 2091 2899 2092 2903
rect 2194 2903 2195 2907
rect 2199 2903 2200 2907
rect 2194 2902 2200 2903
rect 2294 2907 2300 2908
rect 2294 2903 2295 2907
rect 2299 2903 2300 2907
rect 2294 2902 2300 2903
rect 2486 2907 2492 2908
rect 2486 2903 2487 2907
rect 2491 2903 2492 2907
rect 2486 2902 2492 2903
rect 2086 2898 2092 2899
rect 1806 2894 1812 2895
rect 1830 2896 1836 2897
rect 1808 2875 1810 2894
rect 1830 2892 1831 2896
rect 1835 2892 1836 2896
rect 1830 2891 1836 2892
rect 2014 2896 2020 2897
rect 2014 2892 2015 2896
rect 2019 2892 2020 2896
rect 2014 2891 2020 2892
rect 1832 2875 1834 2891
rect 2016 2875 2018 2891
rect 1807 2874 1811 2875
rect 1767 2870 1771 2871
rect 1807 2869 1811 2870
rect 1831 2874 1835 2875
rect 1831 2869 1835 2870
rect 1999 2874 2003 2875
rect 1999 2869 2003 2870
rect 2015 2874 2019 2875
rect 2015 2869 2019 2870
rect 1767 2865 1771 2866
rect 1768 2846 1770 2865
rect 1808 2850 1810 2869
rect 1832 2853 1834 2869
rect 2000 2853 2002 2869
rect 1830 2852 1836 2853
rect 1806 2849 1812 2850
rect 1766 2845 1772 2846
rect 1766 2841 1767 2845
rect 1771 2841 1772 2845
rect 1806 2845 1807 2849
rect 1811 2845 1812 2849
rect 1830 2848 1831 2852
rect 1835 2848 1836 2852
rect 1830 2847 1836 2848
rect 1998 2852 2004 2853
rect 1998 2848 1999 2852
rect 2003 2848 2004 2852
rect 1998 2847 2004 2848
rect 1806 2844 1812 2845
rect 1766 2840 1772 2841
rect 1894 2843 1900 2844
rect 646 2839 652 2840
rect 646 2835 647 2839
rect 651 2835 652 2839
rect 646 2834 652 2835
rect 726 2839 732 2840
rect 726 2835 727 2839
rect 731 2835 732 2839
rect 726 2834 732 2835
rect 966 2839 972 2840
rect 966 2835 967 2839
rect 971 2835 972 2839
rect 966 2834 972 2835
rect 1118 2839 1124 2840
rect 1118 2835 1119 2839
rect 1123 2835 1124 2839
rect 1118 2834 1124 2835
rect 1262 2839 1268 2840
rect 1262 2835 1263 2839
rect 1267 2835 1268 2839
rect 1262 2834 1268 2835
rect 1414 2839 1420 2840
rect 1414 2835 1415 2839
rect 1419 2835 1420 2839
rect 1414 2834 1420 2835
rect 1558 2839 1564 2840
rect 1558 2835 1559 2839
rect 1563 2835 1564 2839
rect 1894 2839 1895 2843
rect 1899 2839 1900 2843
rect 1894 2838 1900 2839
rect 1910 2843 1916 2844
rect 1910 2839 1911 2843
rect 1915 2839 1916 2843
rect 1910 2838 1916 2839
rect 1558 2834 1564 2835
rect 648 2812 650 2834
rect 638 2811 644 2812
rect 638 2807 639 2811
rect 643 2807 644 2811
rect 638 2806 644 2807
rect 646 2811 652 2812
rect 646 2807 647 2811
rect 651 2807 652 2811
rect 646 2806 652 2807
rect 728 2804 730 2834
rect 734 2829 740 2830
rect 734 2825 735 2829
rect 739 2825 740 2829
rect 734 2824 740 2825
rect 894 2829 900 2830
rect 894 2825 895 2829
rect 899 2825 900 2829
rect 894 2824 900 2825
rect 726 2803 732 2804
rect 726 2799 727 2803
rect 731 2799 732 2803
rect 726 2798 732 2799
rect 736 2795 738 2824
rect 896 2795 898 2824
rect 968 2812 970 2834
rect 1046 2829 1052 2830
rect 1046 2825 1047 2829
rect 1051 2825 1052 2829
rect 1046 2824 1052 2825
rect 966 2811 972 2812
rect 966 2807 967 2811
rect 971 2807 972 2811
rect 966 2806 972 2807
rect 1048 2795 1050 2824
rect 1120 2812 1122 2834
rect 1190 2829 1196 2830
rect 1190 2825 1191 2829
rect 1195 2825 1196 2829
rect 1190 2824 1196 2825
rect 1118 2811 1124 2812
rect 1118 2807 1119 2811
rect 1123 2807 1124 2811
rect 1118 2806 1124 2807
rect 1192 2795 1194 2824
rect 1264 2812 1266 2834
rect 1342 2829 1348 2830
rect 1342 2825 1343 2829
rect 1347 2825 1348 2829
rect 1342 2824 1348 2825
rect 1262 2811 1268 2812
rect 1262 2807 1263 2811
rect 1267 2807 1268 2811
rect 1262 2806 1268 2807
rect 1278 2803 1284 2804
rect 1278 2799 1279 2803
rect 1283 2799 1284 2803
rect 1278 2798 1284 2799
rect 247 2794 251 2795
rect 247 2789 251 2790
rect 255 2794 259 2795
rect 255 2789 259 2790
rect 391 2794 395 2795
rect 391 2789 395 2790
rect 415 2794 419 2795
rect 415 2789 419 2790
rect 543 2794 547 2795
rect 543 2789 547 2790
rect 575 2794 579 2795
rect 575 2789 579 2790
rect 695 2794 699 2795
rect 695 2789 699 2790
rect 735 2794 739 2795
rect 735 2789 739 2790
rect 855 2794 859 2795
rect 855 2789 859 2790
rect 895 2794 899 2795
rect 895 2789 899 2790
rect 1023 2794 1027 2795
rect 1023 2789 1027 2790
rect 1047 2794 1051 2795
rect 1047 2789 1051 2790
rect 1191 2794 1195 2795
rect 1191 2789 1195 2790
rect 198 2787 204 2788
rect 198 2783 199 2787
rect 203 2783 204 2787
rect 198 2782 204 2783
rect 206 2787 212 2788
rect 206 2783 207 2787
rect 211 2783 212 2787
rect 206 2782 212 2783
rect 110 2768 111 2772
rect 115 2768 116 2772
rect 110 2767 116 2768
rect 134 2771 140 2772
rect 134 2767 135 2771
rect 139 2767 140 2771
rect 134 2766 140 2767
rect 208 2764 210 2782
rect 248 2772 250 2789
rect 318 2787 324 2788
rect 318 2783 319 2787
rect 323 2783 324 2787
rect 318 2782 324 2783
rect 246 2771 252 2772
rect 246 2767 247 2771
rect 251 2767 252 2771
rect 246 2766 252 2767
rect 320 2764 322 2782
rect 392 2772 394 2789
rect 462 2787 468 2788
rect 462 2783 463 2787
rect 467 2783 468 2787
rect 462 2782 468 2783
rect 390 2771 396 2772
rect 390 2767 391 2771
rect 395 2767 396 2771
rect 390 2766 396 2767
rect 464 2764 466 2782
rect 544 2772 546 2789
rect 614 2787 620 2788
rect 614 2783 615 2787
rect 619 2783 620 2787
rect 614 2782 620 2783
rect 542 2771 548 2772
rect 542 2767 543 2771
rect 547 2767 548 2771
rect 542 2766 548 2767
rect 616 2764 618 2782
rect 696 2772 698 2789
rect 856 2772 858 2789
rect 902 2787 908 2788
rect 902 2783 903 2787
rect 907 2783 908 2787
rect 902 2782 908 2783
rect 926 2787 932 2788
rect 926 2783 927 2787
rect 931 2783 932 2787
rect 926 2782 932 2783
rect 694 2771 700 2772
rect 694 2767 695 2771
rect 699 2767 700 2771
rect 694 2766 700 2767
rect 854 2771 860 2772
rect 854 2767 855 2771
rect 859 2767 860 2771
rect 854 2766 860 2767
rect 206 2763 212 2764
rect 206 2759 207 2763
rect 211 2759 212 2763
rect 206 2758 212 2759
rect 318 2763 324 2764
rect 318 2759 319 2763
rect 323 2759 324 2763
rect 318 2758 324 2759
rect 462 2763 468 2764
rect 462 2759 463 2763
rect 467 2759 468 2763
rect 462 2758 468 2759
rect 614 2763 620 2764
rect 614 2759 615 2763
rect 619 2759 620 2763
rect 614 2758 620 2759
rect 622 2763 628 2764
rect 622 2759 623 2763
rect 627 2759 628 2763
rect 622 2758 628 2759
rect 110 2755 116 2756
rect 110 2751 111 2755
rect 115 2751 116 2755
rect 110 2750 116 2751
rect 134 2752 140 2753
rect 112 2723 114 2750
rect 134 2748 135 2752
rect 139 2748 140 2752
rect 134 2747 140 2748
rect 246 2752 252 2753
rect 246 2748 247 2752
rect 251 2748 252 2752
rect 246 2747 252 2748
rect 390 2752 396 2753
rect 390 2748 391 2752
rect 395 2748 396 2752
rect 390 2747 396 2748
rect 542 2752 548 2753
rect 542 2748 543 2752
rect 547 2748 548 2752
rect 542 2747 548 2748
rect 136 2723 138 2747
rect 248 2723 250 2747
rect 392 2723 394 2747
rect 544 2723 546 2747
rect 111 2722 115 2723
rect 111 2717 115 2718
rect 135 2722 139 2723
rect 135 2717 139 2718
rect 247 2722 251 2723
rect 247 2717 251 2718
rect 359 2722 363 2723
rect 359 2717 363 2718
rect 391 2722 395 2723
rect 391 2717 395 2718
rect 479 2722 483 2723
rect 479 2717 483 2718
rect 543 2722 547 2723
rect 543 2717 547 2718
rect 615 2722 619 2723
rect 615 2717 619 2718
rect 112 2698 114 2717
rect 248 2701 250 2717
rect 298 2715 304 2716
rect 298 2711 299 2715
rect 303 2711 304 2715
rect 298 2710 304 2711
rect 246 2700 252 2701
rect 110 2697 116 2698
rect 110 2693 111 2697
rect 115 2693 116 2697
rect 246 2696 247 2700
rect 251 2696 252 2700
rect 246 2695 252 2696
rect 110 2692 116 2693
rect 246 2681 252 2682
rect 110 2680 116 2681
rect 110 2676 111 2680
rect 115 2676 116 2680
rect 246 2677 247 2681
rect 251 2677 252 2681
rect 246 2676 252 2677
rect 110 2675 116 2676
rect 112 2651 114 2675
rect 248 2651 250 2676
rect 300 2664 302 2710
rect 360 2701 362 2717
rect 480 2701 482 2717
rect 616 2701 618 2717
rect 624 2716 626 2758
rect 694 2752 700 2753
rect 694 2748 695 2752
rect 699 2748 700 2752
rect 694 2747 700 2748
rect 854 2752 860 2753
rect 854 2748 855 2752
rect 859 2748 860 2752
rect 854 2747 860 2748
rect 696 2723 698 2747
rect 856 2723 858 2747
rect 695 2722 699 2723
rect 695 2717 699 2718
rect 759 2722 763 2723
rect 759 2717 763 2718
rect 855 2722 859 2723
rect 855 2717 859 2718
rect 622 2715 628 2716
rect 622 2711 623 2715
rect 627 2711 628 2715
rect 622 2710 628 2711
rect 760 2701 762 2717
rect 358 2700 364 2701
rect 358 2696 359 2700
rect 363 2696 364 2700
rect 358 2695 364 2696
rect 478 2700 484 2701
rect 478 2696 479 2700
rect 483 2696 484 2700
rect 478 2695 484 2696
rect 614 2700 620 2701
rect 614 2696 615 2700
rect 619 2696 620 2700
rect 614 2695 620 2696
rect 758 2700 764 2701
rect 758 2696 759 2700
rect 763 2696 764 2700
rect 758 2695 764 2696
rect 904 2692 906 2782
rect 928 2764 930 2782
rect 1024 2772 1026 2789
rect 1094 2787 1100 2788
rect 1094 2783 1095 2787
rect 1099 2783 1100 2787
rect 1094 2782 1100 2783
rect 1022 2771 1028 2772
rect 1022 2767 1023 2771
rect 1027 2767 1028 2771
rect 1022 2766 1028 2767
rect 1096 2764 1098 2782
rect 1192 2772 1194 2789
rect 1262 2787 1268 2788
rect 1262 2783 1263 2787
rect 1267 2783 1268 2787
rect 1262 2782 1268 2783
rect 1190 2771 1196 2772
rect 1190 2767 1191 2771
rect 1195 2767 1196 2771
rect 1190 2766 1196 2767
rect 1264 2764 1266 2782
rect 1280 2764 1282 2798
rect 1344 2795 1346 2824
rect 1416 2812 1418 2834
rect 1830 2833 1836 2834
rect 1806 2832 1812 2833
rect 1494 2829 1500 2830
rect 1494 2825 1495 2829
rect 1499 2825 1500 2829
rect 1494 2824 1500 2825
rect 1766 2828 1772 2829
rect 1766 2824 1767 2828
rect 1771 2824 1772 2828
rect 1806 2828 1807 2832
rect 1811 2828 1812 2832
rect 1830 2829 1831 2833
rect 1835 2829 1836 2833
rect 1830 2828 1836 2829
rect 1806 2827 1812 2828
rect 1414 2811 1420 2812
rect 1414 2807 1415 2811
rect 1419 2807 1420 2811
rect 1414 2806 1420 2807
rect 1496 2795 1498 2824
rect 1766 2823 1772 2824
rect 1768 2795 1770 2823
rect 1808 2807 1810 2827
rect 1832 2807 1834 2828
rect 1807 2806 1811 2807
rect 1807 2801 1811 2802
rect 1831 2806 1835 2807
rect 1831 2801 1835 2802
rect 1343 2794 1347 2795
rect 1343 2789 1347 2790
rect 1359 2794 1363 2795
rect 1359 2789 1363 2790
rect 1495 2794 1499 2795
rect 1495 2789 1499 2790
rect 1527 2794 1531 2795
rect 1527 2789 1531 2790
rect 1671 2794 1675 2795
rect 1671 2789 1675 2790
rect 1767 2794 1771 2795
rect 1767 2789 1771 2790
rect 1360 2772 1362 2789
rect 1528 2772 1530 2789
rect 1606 2787 1612 2788
rect 1606 2783 1607 2787
rect 1611 2783 1612 2787
rect 1606 2782 1612 2783
rect 1358 2771 1364 2772
rect 1358 2767 1359 2771
rect 1363 2767 1364 2771
rect 1358 2766 1364 2767
rect 1526 2771 1532 2772
rect 1526 2767 1527 2771
rect 1531 2767 1532 2771
rect 1526 2766 1532 2767
rect 1608 2764 1610 2782
rect 1672 2772 1674 2789
rect 1768 2773 1770 2789
rect 1808 2785 1810 2801
rect 1806 2784 1812 2785
rect 1832 2784 1834 2801
rect 1896 2800 1898 2838
rect 1912 2816 1914 2838
rect 1998 2833 2004 2834
rect 1998 2829 1999 2833
rect 2003 2829 2004 2833
rect 1998 2828 2004 2829
rect 1910 2815 1916 2816
rect 1910 2811 1911 2815
rect 1915 2811 1916 2815
rect 1910 2810 1916 2811
rect 2000 2807 2002 2828
rect 2088 2816 2090 2898
rect 2214 2896 2220 2897
rect 2214 2892 2215 2896
rect 2219 2892 2220 2896
rect 2214 2891 2220 2892
rect 2406 2896 2412 2897
rect 2406 2892 2407 2896
rect 2411 2892 2412 2896
rect 2406 2891 2412 2892
rect 2590 2896 2596 2897
rect 2590 2892 2591 2896
rect 2595 2892 2596 2896
rect 2590 2891 2596 2892
rect 2216 2875 2218 2891
rect 2408 2875 2410 2891
rect 2592 2875 2594 2891
rect 2191 2874 2195 2875
rect 2191 2869 2195 2870
rect 2215 2874 2219 2875
rect 2215 2869 2219 2870
rect 2383 2874 2387 2875
rect 2383 2869 2387 2870
rect 2407 2874 2411 2875
rect 2407 2869 2411 2870
rect 2567 2874 2571 2875
rect 2567 2869 2571 2870
rect 2591 2874 2595 2875
rect 2591 2869 2595 2870
rect 2192 2853 2194 2869
rect 2384 2853 2386 2869
rect 2568 2853 2570 2869
rect 2190 2852 2196 2853
rect 2190 2848 2191 2852
rect 2195 2848 2196 2852
rect 2190 2847 2196 2848
rect 2382 2852 2388 2853
rect 2382 2848 2383 2852
rect 2387 2848 2388 2852
rect 2382 2847 2388 2848
rect 2566 2852 2572 2853
rect 2566 2848 2567 2852
rect 2571 2848 2572 2852
rect 2566 2847 2572 2848
rect 2640 2844 2642 2926
rect 2760 2916 2762 2933
rect 2894 2931 2900 2932
rect 2894 2927 2895 2931
rect 2899 2927 2900 2931
rect 2894 2926 2900 2927
rect 2758 2915 2764 2916
rect 2758 2911 2759 2915
rect 2763 2911 2764 2915
rect 2758 2910 2764 2911
rect 2896 2908 2898 2926
rect 2912 2916 2914 2933
rect 2990 2931 2996 2932
rect 2990 2927 2991 2931
rect 2995 2927 2996 2931
rect 2990 2926 2996 2927
rect 2910 2915 2916 2916
rect 2910 2911 2911 2915
rect 2915 2911 2916 2915
rect 2910 2910 2916 2911
rect 2992 2908 2994 2926
rect 3064 2916 3066 2933
rect 3142 2931 3148 2932
rect 3142 2927 3143 2931
rect 3147 2927 3148 2931
rect 3142 2926 3148 2927
rect 3062 2915 3068 2916
rect 3062 2911 3063 2915
rect 3067 2911 3068 2915
rect 3062 2910 3068 2911
rect 3144 2908 3146 2926
rect 3208 2916 3210 2933
rect 3286 2931 3292 2932
rect 3286 2927 3287 2931
rect 3291 2927 3292 2931
rect 3286 2926 3292 2927
rect 3294 2931 3300 2932
rect 3294 2927 3295 2931
rect 3299 2927 3300 2931
rect 3294 2926 3300 2927
rect 3206 2915 3212 2916
rect 3206 2911 3207 2915
rect 3211 2911 3212 2915
rect 3206 2910 3212 2911
rect 3288 2908 3290 2926
rect 2894 2907 2900 2908
rect 2830 2903 2836 2904
rect 2830 2899 2831 2903
rect 2835 2899 2836 2903
rect 2894 2903 2895 2907
rect 2899 2903 2900 2907
rect 2894 2902 2900 2903
rect 2990 2907 2996 2908
rect 2990 2903 2991 2907
rect 2995 2903 2996 2907
rect 2990 2902 2996 2903
rect 3142 2907 3148 2908
rect 3142 2903 3143 2907
rect 3147 2903 3148 2907
rect 3142 2902 3148 2903
rect 3286 2907 3292 2908
rect 3286 2903 3287 2907
rect 3291 2903 3292 2907
rect 3286 2902 3292 2903
rect 2830 2898 2836 2899
rect 2758 2896 2764 2897
rect 2758 2892 2759 2896
rect 2763 2892 2764 2896
rect 2758 2891 2764 2892
rect 2760 2875 2762 2891
rect 2735 2874 2739 2875
rect 2735 2869 2739 2870
rect 2759 2874 2763 2875
rect 2759 2869 2763 2870
rect 2736 2853 2738 2869
rect 2734 2852 2740 2853
rect 2734 2848 2735 2852
rect 2739 2848 2740 2852
rect 2734 2847 2740 2848
rect 2262 2843 2268 2844
rect 2262 2839 2263 2843
rect 2267 2839 2268 2843
rect 2262 2838 2268 2839
rect 2454 2843 2460 2844
rect 2454 2839 2455 2843
rect 2459 2839 2460 2843
rect 2454 2838 2460 2839
rect 2638 2843 2644 2844
rect 2638 2839 2639 2843
rect 2643 2839 2644 2843
rect 2638 2838 2644 2839
rect 2190 2833 2196 2834
rect 2190 2829 2191 2833
rect 2195 2829 2196 2833
rect 2190 2828 2196 2829
rect 2086 2815 2092 2816
rect 2086 2811 2087 2815
rect 2091 2811 2092 2815
rect 2086 2810 2092 2811
rect 2146 2815 2152 2816
rect 2146 2811 2147 2815
rect 2151 2811 2152 2815
rect 2146 2810 2152 2811
rect 1999 2806 2003 2807
rect 1999 2801 2003 2802
rect 2015 2806 2019 2807
rect 2015 2801 2019 2802
rect 1894 2799 1900 2800
rect 1894 2795 1895 2799
rect 1899 2795 1900 2799
rect 1894 2794 1900 2795
rect 2016 2784 2018 2801
rect 2094 2799 2100 2800
rect 2094 2795 2095 2799
rect 2099 2795 2100 2799
rect 2094 2794 2100 2795
rect 1806 2780 1807 2784
rect 1811 2780 1812 2784
rect 1806 2779 1812 2780
rect 1830 2783 1836 2784
rect 1830 2779 1831 2783
rect 1835 2779 1836 2783
rect 1830 2778 1836 2779
rect 2014 2783 2020 2784
rect 2014 2779 2015 2783
rect 2019 2779 2020 2783
rect 2014 2778 2020 2779
rect 2096 2776 2098 2794
rect 2148 2784 2150 2810
rect 2192 2807 2194 2828
rect 2264 2816 2266 2838
rect 2382 2833 2388 2834
rect 2382 2829 2383 2833
rect 2387 2829 2388 2833
rect 2382 2828 2388 2829
rect 2262 2815 2268 2816
rect 2262 2811 2263 2815
rect 2267 2811 2268 2815
rect 2262 2810 2268 2811
rect 2384 2807 2386 2828
rect 2456 2816 2458 2838
rect 2566 2833 2572 2834
rect 2566 2829 2567 2833
rect 2571 2829 2572 2833
rect 2566 2828 2572 2829
rect 2734 2833 2740 2834
rect 2734 2829 2735 2833
rect 2739 2829 2740 2833
rect 2734 2828 2740 2829
rect 2454 2815 2460 2816
rect 2454 2811 2455 2815
rect 2459 2811 2460 2815
rect 2454 2810 2460 2811
rect 2568 2807 2570 2828
rect 2736 2807 2738 2828
rect 2832 2816 2834 2898
rect 2910 2896 2916 2897
rect 2910 2892 2911 2896
rect 2915 2892 2916 2896
rect 2910 2891 2916 2892
rect 3062 2896 3068 2897
rect 3062 2892 3063 2896
rect 3067 2892 3068 2896
rect 3062 2891 3068 2892
rect 3206 2896 3212 2897
rect 3206 2892 3207 2896
rect 3211 2892 3212 2896
rect 3206 2891 3212 2892
rect 2912 2875 2914 2891
rect 3064 2875 3066 2891
rect 3208 2875 3210 2891
rect 2903 2874 2907 2875
rect 2903 2869 2907 2870
rect 2911 2874 2915 2875
rect 2911 2869 2915 2870
rect 3063 2874 3067 2875
rect 3063 2869 3067 2870
rect 3207 2874 3211 2875
rect 3207 2869 3211 2870
rect 3223 2874 3227 2875
rect 3223 2869 3227 2870
rect 2904 2853 2906 2869
rect 3064 2853 3066 2869
rect 3224 2853 3226 2869
rect 2902 2852 2908 2853
rect 2902 2848 2903 2852
rect 2907 2848 2908 2852
rect 2902 2847 2908 2848
rect 3062 2852 3068 2853
rect 3062 2848 3063 2852
rect 3067 2848 3068 2852
rect 3062 2847 3068 2848
rect 3222 2852 3228 2853
rect 3222 2848 3223 2852
rect 3227 2848 3228 2852
rect 3222 2847 3228 2848
rect 3296 2844 3298 2926
rect 3360 2916 3362 2933
rect 3358 2915 3364 2916
rect 3358 2911 3359 2915
rect 3363 2911 3364 2915
rect 3358 2910 3364 2911
rect 3358 2896 3364 2897
rect 3358 2892 3359 2896
rect 3363 2892 3364 2896
rect 3358 2891 3364 2892
rect 3360 2875 3362 2891
rect 3359 2874 3363 2875
rect 3359 2869 3363 2870
rect 3367 2874 3371 2875
rect 3367 2869 3371 2870
rect 3368 2853 3370 2869
rect 3366 2852 3372 2853
rect 3366 2848 3367 2852
rect 3371 2848 3372 2852
rect 3366 2847 3372 2848
rect 2862 2843 2868 2844
rect 2862 2839 2863 2843
rect 2867 2839 2868 2843
rect 2862 2838 2868 2839
rect 2974 2843 2980 2844
rect 2974 2839 2975 2843
rect 2979 2839 2980 2843
rect 2974 2838 2980 2839
rect 3126 2843 3132 2844
rect 3126 2839 3127 2843
rect 3131 2839 3132 2843
rect 3126 2838 3132 2839
rect 3294 2843 3300 2844
rect 3294 2839 3295 2843
rect 3299 2839 3300 2843
rect 3294 2838 3300 2839
rect 3430 2843 3436 2844
rect 3430 2839 3431 2843
rect 3435 2839 3436 2843
rect 3430 2838 3436 2839
rect 2864 2816 2866 2838
rect 2902 2833 2908 2834
rect 2902 2829 2903 2833
rect 2907 2829 2908 2833
rect 2902 2828 2908 2829
rect 2830 2815 2836 2816
rect 2830 2811 2831 2815
rect 2835 2811 2836 2815
rect 2830 2810 2836 2811
rect 2862 2815 2868 2816
rect 2862 2811 2863 2815
rect 2867 2811 2868 2815
rect 2862 2810 2868 2811
rect 2904 2807 2906 2828
rect 2976 2816 2978 2838
rect 3062 2833 3068 2834
rect 3062 2829 3063 2833
rect 3067 2829 3068 2833
rect 3062 2828 3068 2829
rect 2974 2815 2980 2816
rect 2974 2811 2975 2815
rect 2979 2811 2980 2815
rect 2974 2810 2980 2811
rect 2990 2807 2996 2808
rect 3064 2807 3066 2828
rect 2191 2806 2195 2807
rect 2191 2801 2195 2802
rect 2215 2806 2219 2807
rect 2215 2801 2219 2802
rect 2383 2806 2387 2807
rect 2383 2801 2387 2802
rect 2407 2806 2411 2807
rect 2407 2801 2411 2802
rect 2567 2806 2571 2807
rect 2567 2801 2571 2802
rect 2583 2806 2587 2807
rect 2583 2801 2587 2802
rect 2735 2806 2739 2807
rect 2735 2801 2739 2802
rect 2751 2806 2755 2807
rect 2751 2801 2755 2802
rect 2903 2806 2907 2807
rect 2903 2801 2907 2802
rect 2911 2806 2915 2807
rect 2990 2803 2991 2807
rect 2995 2803 2996 2807
rect 2990 2802 2996 2803
rect 3063 2806 3067 2807
rect 2911 2801 2915 2802
rect 2216 2784 2218 2801
rect 2294 2799 2300 2800
rect 2294 2795 2295 2799
rect 2299 2795 2300 2799
rect 2294 2794 2300 2795
rect 2146 2783 2152 2784
rect 2146 2779 2147 2783
rect 2151 2779 2152 2783
rect 2146 2778 2152 2779
rect 2214 2783 2220 2784
rect 2214 2779 2215 2783
rect 2219 2779 2220 2783
rect 2214 2778 2220 2779
rect 2296 2776 2298 2794
rect 2408 2784 2410 2801
rect 2470 2799 2476 2800
rect 2470 2795 2471 2799
rect 2475 2795 2476 2799
rect 2470 2794 2476 2795
rect 2406 2783 2412 2784
rect 2406 2779 2407 2783
rect 2411 2779 2412 2783
rect 2406 2778 2412 2779
rect 2094 2775 2100 2776
rect 1766 2772 1772 2773
rect 1670 2771 1676 2772
rect 1670 2767 1671 2771
rect 1675 2767 1676 2771
rect 1766 2768 1767 2772
rect 1771 2768 1772 2772
rect 2094 2771 2095 2775
rect 2099 2771 2100 2775
rect 2094 2770 2100 2771
rect 2294 2775 2300 2776
rect 2294 2771 2295 2775
rect 2299 2771 2300 2775
rect 2294 2770 2300 2771
rect 1766 2767 1772 2768
rect 1806 2767 1812 2768
rect 1670 2766 1676 2767
rect 926 2763 932 2764
rect 926 2759 927 2763
rect 931 2759 932 2763
rect 926 2758 932 2759
rect 1094 2763 1100 2764
rect 1094 2759 1095 2763
rect 1099 2759 1100 2763
rect 1094 2758 1100 2759
rect 1262 2763 1268 2764
rect 1262 2759 1263 2763
rect 1267 2759 1268 2763
rect 1262 2758 1268 2759
rect 1278 2763 1284 2764
rect 1278 2759 1279 2763
rect 1283 2759 1284 2763
rect 1606 2763 1612 2764
rect 1278 2758 1284 2759
rect 1598 2759 1604 2760
rect 1598 2755 1599 2759
rect 1603 2755 1604 2759
rect 1606 2759 1607 2763
rect 1611 2759 1612 2763
rect 1806 2763 1807 2767
rect 1811 2763 1812 2767
rect 1806 2762 1812 2763
rect 1830 2764 1836 2765
rect 1606 2758 1612 2759
rect 1598 2754 1604 2755
rect 1766 2755 1772 2756
rect 1022 2752 1028 2753
rect 1022 2748 1023 2752
rect 1027 2748 1028 2752
rect 1022 2747 1028 2748
rect 1190 2752 1196 2753
rect 1190 2748 1191 2752
rect 1195 2748 1196 2752
rect 1190 2747 1196 2748
rect 1358 2752 1364 2753
rect 1358 2748 1359 2752
rect 1363 2748 1364 2752
rect 1358 2747 1364 2748
rect 1526 2752 1532 2753
rect 1526 2748 1527 2752
rect 1531 2748 1532 2752
rect 1526 2747 1532 2748
rect 1024 2723 1026 2747
rect 1192 2723 1194 2747
rect 1360 2723 1362 2747
rect 1528 2723 1530 2747
rect 911 2722 915 2723
rect 911 2717 915 2718
rect 1023 2722 1027 2723
rect 1023 2717 1027 2718
rect 1063 2722 1067 2723
rect 1063 2717 1067 2718
rect 1191 2722 1195 2723
rect 1191 2717 1195 2718
rect 1215 2722 1219 2723
rect 1215 2717 1219 2718
rect 1359 2722 1363 2723
rect 1359 2717 1363 2718
rect 1375 2722 1379 2723
rect 1375 2717 1379 2718
rect 1527 2722 1531 2723
rect 1527 2717 1531 2718
rect 1535 2722 1539 2723
rect 1535 2717 1539 2718
rect 912 2701 914 2717
rect 1064 2701 1066 2717
rect 1216 2701 1218 2717
rect 1376 2701 1378 2717
rect 1536 2701 1538 2717
rect 910 2700 916 2701
rect 910 2696 911 2700
rect 915 2696 916 2700
rect 910 2695 916 2696
rect 1062 2700 1068 2701
rect 1062 2696 1063 2700
rect 1067 2696 1068 2700
rect 1062 2695 1068 2696
rect 1214 2700 1220 2701
rect 1214 2696 1215 2700
rect 1219 2696 1220 2700
rect 1214 2695 1220 2696
rect 1374 2700 1380 2701
rect 1374 2696 1375 2700
rect 1379 2696 1380 2700
rect 1374 2695 1380 2696
rect 1534 2700 1540 2701
rect 1534 2696 1535 2700
rect 1539 2696 1540 2700
rect 1534 2695 1540 2696
rect 318 2691 324 2692
rect 318 2687 319 2691
rect 323 2687 324 2691
rect 318 2686 324 2687
rect 430 2691 436 2692
rect 430 2687 431 2691
rect 435 2687 436 2691
rect 430 2686 436 2687
rect 550 2691 556 2692
rect 550 2687 551 2691
rect 555 2687 556 2691
rect 550 2686 556 2687
rect 686 2691 692 2692
rect 686 2687 687 2691
rect 691 2687 692 2691
rect 686 2686 692 2687
rect 694 2691 700 2692
rect 694 2687 695 2691
rect 699 2687 700 2691
rect 694 2686 700 2687
rect 902 2691 908 2692
rect 902 2687 903 2691
rect 907 2687 908 2691
rect 902 2686 908 2687
rect 1134 2691 1140 2692
rect 1134 2687 1135 2691
rect 1139 2687 1140 2691
rect 1134 2686 1140 2687
rect 1446 2691 1452 2692
rect 1446 2687 1447 2691
rect 1451 2687 1452 2691
rect 1446 2686 1452 2687
rect 320 2664 322 2686
rect 358 2681 364 2682
rect 358 2677 359 2681
rect 363 2677 364 2681
rect 358 2676 364 2677
rect 298 2663 304 2664
rect 298 2659 299 2663
rect 303 2659 304 2663
rect 298 2658 304 2659
rect 318 2663 324 2664
rect 318 2659 319 2663
rect 323 2659 324 2663
rect 318 2658 324 2659
rect 360 2651 362 2676
rect 432 2664 434 2686
rect 478 2681 484 2682
rect 478 2677 479 2681
rect 483 2677 484 2681
rect 478 2676 484 2677
rect 430 2663 436 2664
rect 430 2659 431 2663
rect 435 2659 436 2663
rect 430 2658 436 2659
rect 480 2651 482 2676
rect 552 2664 554 2686
rect 614 2681 620 2682
rect 614 2677 615 2681
rect 619 2677 620 2681
rect 614 2676 620 2677
rect 550 2663 556 2664
rect 550 2659 551 2663
rect 555 2659 556 2663
rect 550 2658 556 2659
rect 616 2651 618 2676
rect 688 2664 690 2686
rect 686 2663 692 2664
rect 686 2659 687 2663
rect 691 2659 692 2663
rect 686 2658 692 2659
rect 696 2652 698 2686
rect 758 2681 764 2682
rect 758 2677 759 2681
rect 763 2677 764 2681
rect 758 2676 764 2677
rect 910 2681 916 2682
rect 910 2677 911 2681
rect 915 2677 916 2681
rect 910 2676 916 2677
rect 1062 2681 1068 2682
rect 1062 2677 1063 2681
rect 1067 2677 1068 2681
rect 1062 2676 1068 2677
rect 694 2651 700 2652
rect 760 2651 762 2676
rect 912 2651 914 2676
rect 1054 2663 1060 2664
rect 1054 2659 1055 2663
rect 1059 2659 1060 2663
rect 1054 2658 1060 2659
rect 111 2650 115 2651
rect 111 2645 115 2646
rect 247 2650 251 2651
rect 247 2645 251 2646
rect 359 2650 363 2651
rect 359 2645 363 2646
rect 463 2650 467 2651
rect 463 2645 467 2646
rect 479 2650 483 2651
rect 479 2645 483 2646
rect 551 2650 555 2651
rect 551 2645 555 2646
rect 615 2650 619 2651
rect 615 2645 619 2646
rect 639 2650 643 2651
rect 694 2647 695 2651
rect 699 2647 700 2651
rect 694 2646 700 2647
rect 743 2650 747 2651
rect 639 2645 643 2646
rect 743 2645 747 2646
rect 759 2650 763 2651
rect 759 2645 763 2646
rect 855 2650 859 2651
rect 855 2645 859 2646
rect 911 2650 915 2651
rect 911 2645 915 2646
rect 983 2650 987 2651
rect 983 2645 987 2646
rect 112 2629 114 2645
rect 110 2628 116 2629
rect 464 2628 466 2645
rect 534 2643 540 2644
rect 534 2639 535 2643
rect 539 2639 540 2643
rect 534 2638 540 2639
rect 110 2624 111 2628
rect 115 2624 116 2628
rect 110 2623 116 2624
rect 462 2627 468 2628
rect 462 2623 463 2627
rect 467 2623 468 2627
rect 462 2622 468 2623
rect 536 2620 538 2638
rect 552 2628 554 2645
rect 622 2643 628 2644
rect 622 2639 623 2643
rect 627 2639 628 2643
rect 622 2638 628 2639
rect 550 2627 556 2628
rect 550 2623 551 2627
rect 555 2623 556 2627
rect 550 2622 556 2623
rect 624 2620 626 2638
rect 640 2628 642 2645
rect 710 2643 716 2644
rect 710 2639 711 2643
rect 715 2639 716 2643
rect 710 2638 716 2639
rect 638 2627 644 2628
rect 638 2623 639 2627
rect 643 2623 644 2627
rect 638 2622 644 2623
rect 712 2620 714 2638
rect 744 2628 746 2645
rect 814 2643 820 2644
rect 814 2639 815 2643
rect 819 2639 820 2643
rect 814 2638 820 2639
rect 742 2627 748 2628
rect 742 2623 743 2627
rect 747 2623 748 2627
rect 742 2622 748 2623
rect 816 2620 818 2638
rect 856 2628 858 2645
rect 984 2628 986 2645
rect 854 2627 860 2628
rect 854 2623 855 2627
rect 859 2623 860 2627
rect 854 2622 860 2623
rect 982 2627 988 2628
rect 982 2623 983 2627
rect 987 2623 988 2627
rect 982 2622 988 2623
rect 1056 2620 1058 2658
rect 1064 2651 1066 2676
rect 1136 2664 1138 2686
rect 1214 2681 1220 2682
rect 1214 2677 1215 2681
rect 1219 2677 1220 2681
rect 1214 2676 1220 2677
rect 1374 2681 1380 2682
rect 1374 2677 1375 2681
rect 1379 2677 1380 2681
rect 1374 2676 1380 2677
rect 1134 2663 1140 2664
rect 1134 2659 1135 2663
rect 1139 2659 1140 2663
rect 1134 2658 1140 2659
rect 1216 2651 1218 2676
rect 1376 2651 1378 2676
rect 1063 2650 1067 2651
rect 1063 2645 1067 2646
rect 1127 2650 1131 2651
rect 1127 2645 1131 2646
rect 1215 2650 1219 2651
rect 1215 2645 1219 2646
rect 1279 2650 1283 2651
rect 1279 2645 1283 2646
rect 1375 2650 1379 2651
rect 1375 2645 1379 2646
rect 1439 2650 1443 2651
rect 1439 2645 1443 2646
rect 1106 2643 1112 2644
rect 1106 2639 1107 2643
rect 1111 2639 1112 2643
rect 1106 2638 1112 2639
rect 1108 2620 1110 2638
rect 1128 2628 1130 2645
rect 1206 2643 1212 2644
rect 1206 2639 1207 2643
rect 1211 2639 1212 2643
rect 1206 2638 1212 2639
rect 1126 2627 1132 2628
rect 1126 2623 1127 2627
rect 1131 2623 1132 2627
rect 1126 2622 1132 2623
rect 1208 2620 1210 2638
rect 1280 2628 1282 2645
rect 1294 2643 1300 2644
rect 1294 2639 1295 2643
rect 1299 2639 1300 2643
rect 1294 2638 1300 2639
rect 1278 2627 1284 2628
rect 1278 2623 1279 2627
rect 1283 2623 1284 2627
rect 1278 2622 1284 2623
rect 534 2619 540 2620
rect 534 2615 535 2619
rect 539 2615 540 2619
rect 534 2614 540 2615
rect 622 2619 628 2620
rect 622 2615 623 2619
rect 627 2615 628 2619
rect 622 2614 628 2615
rect 710 2619 716 2620
rect 710 2615 711 2619
rect 715 2615 716 2619
rect 710 2614 716 2615
rect 814 2619 820 2620
rect 814 2615 815 2619
rect 819 2615 820 2619
rect 814 2614 820 2615
rect 822 2619 828 2620
rect 822 2615 823 2619
rect 827 2615 828 2619
rect 822 2614 828 2615
rect 1054 2619 1060 2620
rect 1054 2615 1055 2619
rect 1059 2615 1060 2619
rect 1054 2614 1060 2615
rect 1106 2619 1112 2620
rect 1106 2615 1107 2619
rect 1111 2615 1112 2619
rect 1106 2614 1112 2615
rect 1206 2619 1212 2620
rect 1206 2615 1207 2619
rect 1211 2615 1212 2619
rect 1206 2614 1212 2615
rect 110 2611 116 2612
rect 110 2607 111 2611
rect 115 2607 116 2611
rect 110 2606 116 2607
rect 462 2608 468 2609
rect 112 2579 114 2606
rect 462 2604 463 2608
rect 467 2604 468 2608
rect 462 2603 468 2604
rect 550 2608 556 2609
rect 550 2604 551 2608
rect 555 2604 556 2608
rect 550 2603 556 2604
rect 638 2608 644 2609
rect 638 2604 639 2608
rect 643 2604 644 2608
rect 638 2603 644 2604
rect 742 2608 748 2609
rect 742 2604 743 2608
rect 747 2604 748 2608
rect 742 2603 748 2604
rect 464 2579 466 2603
rect 552 2579 554 2603
rect 640 2579 642 2603
rect 744 2579 746 2603
rect 111 2578 115 2579
rect 111 2573 115 2574
rect 463 2578 467 2579
rect 463 2573 467 2574
rect 503 2578 507 2579
rect 503 2573 507 2574
rect 551 2578 555 2579
rect 551 2573 555 2574
rect 591 2578 595 2579
rect 591 2573 595 2574
rect 639 2578 643 2579
rect 639 2573 643 2574
rect 679 2578 683 2579
rect 679 2573 683 2574
rect 743 2578 747 2579
rect 743 2573 747 2574
rect 775 2578 779 2579
rect 775 2573 779 2574
rect 112 2554 114 2573
rect 504 2557 506 2573
rect 592 2557 594 2573
rect 680 2557 682 2573
rect 776 2557 778 2573
rect 502 2556 508 2557
rect 110 2553 116 2554
rect 110 2549 111 2553
rect 115 2549 116 2553
rect 502 2552 503 2556
rect 507 2552 508 2556
rect 502 2551 508 2552
rect 590 2556 596 2557
rect 590 2552 591 2556
rect 595 2552 596 2556
rect 590 2551 596 2552
rect 678 2556 684 2557
rect 678 2552 679 2556
rect 683 2552 684 2556
rect 678 2551 684 2552
rect 774 2556 780 2557
rect 774 2552 775 2556
rect 779 2552 780 2556
rect 774 2551 780 2552
rect 110 2548 116 2549
rect 574 2547 580 2548
rect 574 2543 575 2547
rect 579 2543 580 2547
rect 574 2542 580 2543
rect 662 2547 668 2548
rect 662 2543 663 2547
rect 667 2543 668 2547
rect 662 2542 668 2543
rect 750 2547 756 2548
rect 750 2543 751 2547
rect 755 2543 756 2547
rect 750 2542 756 2543
rect 502 2537 508 2538
rect 110 2536 116 2537
rect 110 2532 111 2536
rect 115 2532 116 2536
rect 502 2533 503 2537
rect 507 2533 508 2537
rect 502 2532 508 2533
rect 110 2531 116 2532
rect 112 2507 114 2531
rect 504 2507 506 2532
rect 576 2520 578 2542
rect 590 2537 596 2538
rect 590 2533 591 2537
rect 595 2533 596 2537
rect 590 2532 596 2533
rect 574 2519 580 2520
rect 574 2515 575 2519
rect 579 2515 580 2519
rect 574 2514 580 2515
rect 592 2507 594 2532
rect 664 2520 666 2542
rect 678 2537 684 2538
rect 678 2533 679 2537
rect 683 2533 684 2537
rect 678 2532 684 2533
rect 662 2519 668 2520
rect 662 2515 663 2519
rect 667 2515 668 2519
rect 662 2514 668 2515
rect 680 2507 682 2532
rect 752 2520 754 2542
rect 774 2537 780 2538
rect 774 2533 775 2537
rect 779 2533 780 2537
rect 774 2532 780 2533
rect 750 2519 756 2520
rect 750 2515 751 2519
rect 755 2515 756 2519
rect 750 2514 756 2515
rect 776 2507 778 2532
rect 824 2512 826 2614
rect 854 2608 860 2609
rect 854 2604 855 2608
rect 859 2604 860 2608
rect 854 2603 860 2604
rect 982 2608 988 2609
rect 982 2604 983 2608
rect 987 2604 988 2608
rect 982 2603 988 2604
rect 1126 2608 1132 2609
rect 1126 2604 1127 2608
rect 1131 2604 1132 2608
rect 1126 2603 1132 2604
rect 1278 2608 1284 2609
rect 1278 2604 1279 2608
rect 1283 2604 1284 2608
rect 1278 2603 1284 2604
rect 856 2579 858 2603
rect 984 2579 986 2603
rect 1128 2579 1130 2603
rect 1280 2579 1282 2603
rect 855 2578 859 2579
rect 855 2573 859 2574
rect 879 2578 883 2579
rect 879 2573 883 2574
rect 983 2578 987 2579
rect 983 2573 987 2574
rect 991 2578 995 2579
rect 991 2573 995 2574
rect 1103 2578 1107 2579
rect 1103 2573 1107 2574
rect 1127 2578 1131 2579
rect 1127 2573 1131 2574
rect 1223 2578 1227 2579
rect 1223 2573 1227 2574
rect 1279 2578 1283 2579
rect 1279 2573 1283 2574
rect 880 2557 882 2573
rect 992 2557 994 2573
rect 1104 2557 1106 2573
rect 1224 2557 1226 2573
rect 878 2556 884 2557
rect 878 2552 879 2556
rect 883 2552 884 2556
rect 878 2551 884 2552
rect 990 2556 996 2557
rect 990 2552 991 2556
rect 995 2552 996 2556
rect 990 2551 996 2552
rect 1102 2556 1108 2557
rect 1102 2552 1103 2556
rect 1107 2552 1108 2556
rect 1102 2551 1108 2552
rect 1222 2556 1228 2557
rect 1222 2552 1223 2556
rect 1227 2552 1228 2556
rect 1222 2551 1228 2552
rect 1296 2548 1298 2638
rect 1440 2628 1442 2645
rect 1448 2644 1450 2686
rect 1534 2681 1540 2682
rect 1534 2677 1535 2681
rect 1539 2677 1540 2681
rect 1534 2676 1540 2677
rect 1536 2651 1538 2676
rect 1600 2664 1602 2754
rect 1670 2752 1676 2753
rect 1670 2748 1671 2752
rect 1675 2748 1676 2752
rect 1766 2751 1767 2755
rect 1771 2751 1772 2755
rect 1766 2750 1772 2751
rect 1670 2747 1676 2748
rect 1672 2723 1674 2747
rect 1768 2723 1770 2750
rect 1808 2727 1810 2762
rect 1830 2760 1831 2764
rect 1835 2760 1836 2764
rect 1830 2759 1836 2760
rect 2014 2764 2020 2765
rect 2014 2760 2015 2764
rect 2019 2760 2020 2764
rect 2014 2759 2020 2760
rect 2214 2764 2220 2765
rect 2214 2760 2215 2764
rect 2219 2760 2220 2764
rect 2214 2759 2220 2760
rect 2406 2764 2412 2765
rect 2406 2760 2407 2764
rect 2411 2760 2412 2764
rect 2406 2759 2412 2760
rect 1832 2727 1834 2759
rect 2016 2727 2018 2759
rect 2216 2727 2218 2759
rect 2408 2727 2410 2759
rect 1807 2726 1811 2727
rect 1671 2722 1675 2723
rect 1671 2717 1675 2718
rect 1767 2722 1771 2723
rect 1807 2721 1811 2722
rect 1831 2726 1835 2727
rect 1831 2721 1835 2722
rect 2015 2726 2019 2727
rect 2015 2721 2019 2722
rect 2039 2726 2043 2727
rect 2039 2721 2043 2722
rect 2159 2726 2163 2727
rect 2159 2721 2163 2722
rect 2215 2726 2219 2727
rect 2215 2721 2219 2722
rect 2279 2726 2283 2727
rect 2279 2721 2283 2722
rect 2407 2726 2411 2727
rect 2407 2721 2411 2722
rect 1767 2717 1771 2718
rect 1672 2701 1674 2717
rect 1670 2700 1676 2701
rect 1670 2696 1671 2700
rect 1675 2696 1676 2700
rect 1768 2698 1770 2717
rect 1808 2702 1810 2721
rect 2040 2705 2042 2721
rect 2160 2705 2162 2721
rect 2280 2705 2282 2721
rect 2408 2705 2410 2721
rect 2038 2704 2044 2705
rect 1806 2701 1812 2702
rect 1670 2695 1676 2696
rect 1766 2697 1772 2698
rect 1766 2693 1767 2697
rect 1771 2693 1772 2697
rect 1806 2697 1807 2701
rect 1811 2697 1812 2701
rect 2038 2700 2039 2704
rect 2043 2700 2044 2704
rect 2038 2699 2044 2700
rect 2158 2704 2164 2705
rect 2158 2700 2159 2704
rect 2163 2700 2164 2704
rect 2158 2699 2164 2700
rect 2278 2704 2284 2705
rect 2278 2700 2279 2704
rect 2283 2700 2284 2704
rect 2278 2699 2284 2700
rect 2406 2704 2412 2705
rect 2406 2700 2407 2704
rect 2411 2700 2412 2704
rect 2406 2699 2412 2700
rect 1806 2696 1812 2697
rect 2472 2696 2474 2794
rect 2584 2784 2586 2801
rect 2742 2799 2748 2800
rect 2742 2795 2743 2799
rect 2747 2795 2748 2799
rect 2742 2794 2748 2795
rect 2582 2783 2588 2784
rect 2582 2779 2583 2783
rect 2587 2779 2588 2783
rect 2582 2778 2588 2779
rect 2744 2776 2746 2794
rect 2752 2784 2754 2801
rect 2822 2799 2828 2800
rect 2822 2795 2823 2799
rect 2827 2795 2828 2799
rect 2822 2794 2828 2795
rect 2750 2783 2756 2784
rect 2750 2779 2751 2783
rect 2755 2779 2756 2783
rect 2750 2778 2756 2779
rect 2824 2776 2826 2794
rect 2912 2784 2914 2801
rect 2910 2783 2916 2784
rect 2910 2779 2911 2783
rect 2915 2779 2916 2783
rect 2910 2778 2916 2779
rect 2992 2776 2994 2802
rect 3063 2801 3067 2802
rect 3071 2806 3075 2807
rect 3071 2801 3075 2802
rect 3072 2784 3074 2801
rect 3119 2799 3125 2800
rect 3119 2795 3120 2799
rect 3124 2798 3125 2799
rect 3128 2798 3130 2838
rect 3222 2833 3228 2834
rect 3222 2829 3223 2833
rect 3227 2829 3228 2833
rect 3222 2828 3228 2829
rect 3366 2833 3372 2834
rect 3366 2829 3367 2833
rect 3371 2829 3372 2833
rect 3366 2828 3372 2829
rect 3224 2807 3226 2828
rect 3302 2815 3308 2816
rect 3302 2811 3303 2815
rect 3307 2811 3308 2815
rect 3302 2810 3308 2811
rect 3223 2806 3227 2807
rect 3223 2801 3227 2802
rect 3231 2806 3235 2807
rect 3231 2801 3235 2802
rect 3124 2796 3130 2798
rect 3124 2795 3125 2796
rect 3119 2794 3125 2795
rect 3232 2784 3234 2801
rect 3262 2799 3268 2800
rect 3262 2795 3263 2799
rect 3267 2795 3268 2799
rect 3262 2794 3268 2795
rect 3070 2783 3076 2784
rect 3070 2779 3071 2783
rect 3075 2779 3076 2783
rect 3070 2778 3076 2779
rect 3230 2783 3236 2784
rect 3230 2779 3231 2783
rect 3235 2779 3236 2783
rect 3230 2778 3236 2779
rect 2742 2775 2748 2776
rect 2742 2771 2743 2775
rect 2747 2771 2748 2775
rect 2742 2770 2748 2771
rect 2822 2775 2828 2776
rect 2822 2771 2823 2775
rect 2827 2771 2828 2775
rect 2990 2775 2996 2776
rect 2822 2770 2828 2771
rect 2982 2771 2988 2772
rect 2982 2767 2983 2771
rect 2987 2767 2988 2771
rect 2990 2771 2991 2775
rect 2995 2771 2996 2775
rect 2990 2770 2996 2771
rect 2982 2766 2988 2767
rect 2582 2764 2588 2765
rect 2582 2760 2583 2764
rect 2587 2760 2588 2764
rect 2582 2759 2588 2760
rect 2750 2764 2756 2765
rect 2750 2760 2751 2764
rect 2755 2760 2756 2764
rect 2750 2759 2756 2760
rect 2910 2764 2916 2765
rect 2910 2760 2911 2764
rect 2915 2760 2916 2764
rect 2910 2759 2916 2760
rect 2584 2727 2586 2759
rect 2752 2727 2754 2759
rect 2912 2727 2914 2759
rect 2543 2726 2547 2727
rect 2543 2721 2547 2722
rect 2583 2726 2587 2727
rect 2583 2721 2587 2722
rect 2687 2726 2691 2727
rect 2687 2721 2691 2722
rect 2751 2726 2755 2727
rect 2751 2721 2755 2722
rect 2847 2726 2851 2727
rect 2847 2721 2851 2722
rect 2911 2726 2915 2727
rect 2911 2721 2915 2722
rect 2544 2705 2546 2721
rect 2688 2705 2690 2721
rect 2848 2705 2850 2721
rect 2542 2704 2548 2705
rect 2542 2700 2543 2704
rect 2547 2700 2548 2704
rect 2542 2699 2548 2700
rect 2686 2704 2692 2705
rect 2686 2700 2687 2704
rect 2691 2700 2692 2704
rect 2686 2699 2692 2700
rect 2846 2704 2852 2705
rect 2846 2700 2847 2704
rect 2851 2700 2852 2704
rect 2846 2699 2852 2700
rect 1766 2692 1772 2693
rect 2110 2695 2116 2696
rect 1606 2691 1612 2692
rect 1606 2687 1607 2691
rect 1611 2687 1612 2691
rect 1606 2686 1612 2687
rect 1638 2691 1644 2692
rect 1638 2687 1639 2691
rect 1643 2687 1644 2691
rect 2110 2691 2111 2695
rect 2115 2691 2116 2695
rect 2110 2690 2116 2691
rect 2230 2695 2236 2696
rect 2230 2691 2231 2695
rect 2235 2691 2236 2695
rect 2230 2690 2236 2691
rect 2350 2695 2356 2696
rect 2350 2691 2351 2695
rect 2355 2691 2356 2695
rect 2350 2690 2356 2691
rect 2470 2695 2476 2696
rect 2470 2691 2471 2695
rect 2475 2691 2476 2695
rect 2470 2690 2476 2691
rect 2614 2695 2620 2696
rect 2614 2691 2615 2695
rect 2619 2691 2620 2695
rect 2614 2690 2620 2691
rect 2766 2695 2772 2696
rect 2766 2691 2767 2695
rect 2771 2691 2772 2695
rect 2766 2690 2772 2691
rect 2774 2695 2780 2696
rect 2774 2691 2775 2695
rect 2779 2691 2780 2695
rect 2774 2690 2780 2691
rect 1638 2686 1644 2687
rect 1608 2664 1610 2686
rect 1598 2663 1604 2664
rect 1598 2659 1599 2663
rect 1603 2659 1604 2663
rect 1598 2658 1604 2659
rect 1606 2663 1612 2664
rect 1606 2659 1607 2663
rect 1611 2659 1612 2663
rect 1606 2658 1612 2659
rect 1640 2656 1642 2686
rect 2038 2685 2044 2686
rect 1806 2684 1812 2685
rect 1670 2681 1676 2682
rect 1670 2677 1671 2681
rect 1675 2677 1676 2681
rect 1670 2676 1676 2677
rect 1766 2680 1772 2681
rect 1766 2676 1767 2680
rect 1771 2676 1772 2680
rect 1806 2680 1807 2684
rect 1811 2680 1812 2684
rect 2038 2681 2039 2685
rect 2043 2681 2044 2685
rect 2038 2680 2044 2681
rect 1806 2679 1812 2680
rect 1638 2655 1644 2656
rect 1638 2651 1639 2655
rect 1643 2651 1644 2655
rect 1672 2651 1674 2676
rect 1766 2675 1772 2676
rect 1768 2651 1770 2675
rect 1808 2651 1810 2679
rect 2040 2651 2042 2680
rect 2112 2668 2114 2690
rect 2158 2685 2164 2686
rect 2158 2681 2159 2685
rect 2163 2681 2164 2685
rect 2158 2680 2164 2681
rect 2110 2667 2116 2668
rect 2110 2663 2111 2667
rect 2115 2663 2116 2667
rect 2110 2662 2116 2663
rect 2160 2651 2162 2680
rect 2232 2668 2234 2690
rect 2278 2685 2284 2686
rect 2278 2681 2279 2685
rect 2283 2681 2284 2685
rect 2278 2680 2284 2681
rect 2230 2667 2236 2668
rect 2230 2663 2231 2667
rect 2235 2663 2236 2667
rect 2230 2662 2236 2663
rect 2262 2659 2268 2660
rect 2262 2655 2263 2659
rect 2267 2655 2268 2659
rect 2262 2654 2268 2655
rect 1535 2650 1539 2651
rect 1535 2645 1539 2646
rect 1607 2650 1611 2651
rect 1638 2650 1644 2651
rect 1671 2650 1675 2651
rect 1607 2645 1611 2646
rect 1671 2645 1675 2646
rect 1767 2650 1771 2651
rect 1767 2645 1771 2646
rect 1807 2650 1811 2651
rect 1807 2645 1811 2646
rect 1871 2650 1875 2651
rect 1871 2645 1875 2646
rect 1967 2650 1971 2651
rect 1967 2645 1971 2646
rect 2039 2650 2043 2651
rect 2039 2645 2043 2646
rect 2071 2650 2075 2651
rect 2071 2645 2075 2646
rect 2159 2650 2163 2651
rect 2159 2645 2163 2646
rect 2183 2650 2187 2651
rect 2183 2645 2187 2646
rect 1446 2643 1452 2644
rect 1446 2639 1447 2643
rect 1451 2639 1452 2643
rect 1446 2638 1452 2639
rect 1510 2643 1516 2644
rect 1510 2639 1511 2643
rect 1515 2639 1516 2643
rect 1510 2638 1516 2639
rect 1438 2627 1444 2628
rect 1438 2623 1439 2627
rect 1443 2623 1444 2627
rect 1438 2622 1444 2623
rect 1512 2620 1514 2638
rect 1608 2628 1610 2645
rect 1768 2629 1770 2645
rect 1808 2629 1810 2645
rect 1766 2628 1772 2629
rect 1606 2627 1612 2628
rect 1606 2623 1607 2627
rect 1611 2623 1612 2627
rect 1766 2624 1767 2628
rect 1771 2624 1772 2628
rect 1766 2623 1772 2624
rect 1806 2628 1812 2629
rect 1872 2628 1874 2645
rect 1902 2643 1908 2644
rect 1902 2639 1903 2643
rect 1907 2639 1908 2643
rect 1902 2638 1908 2639
rect 1942 2643 1948 2644
rect 1942 2639 1943 2643
rect 1947 2639 1948 2643
rect 1942 2638 1948 2639
rect 1806 2624 1807 2628
rect 1811 2624 1812 2628
rect 1806 2623 1812 2624
rect 1870 2627 1876 2628
rect 1870 2623 1871 2627
rect 1875 2623 1876 2627
rect 1606 2622 1612 2623
rect 1870 2622 1876 2623
rect 1510 2619 1516 2620
rect 1510 2615 1511 2619
rect 1515 2615 1516 2619
rect 1510 2614 1516 2615
rect 1678 2615 1684 2616
rect 1678 2611 1679 2615
rect 1683 2611 1684 2615
rect 1678 2610 1684 2611
rect 1766 2611 1772 2612
rect 1438 2608 1444 2609
rect 1438 2604 1439 2608
rect 1443 2604 1444 2608
rect 1438 2603 1444 2604
rect 1606 2608 1612 2609
rect 1606 2604 1607 2608
rect 1611 2604 1612 2608
rect 1606 2603 1612 2604
rect 1440 2579 1442 2603
rect 1608 2579 1610 2603
rect 1351 2578 1355 2579
rect 1351 2573 1355 2574
rect 1439 2578 1443 2579
rect 1439 2573 1443 2574
rect 1479 2578 1483 2579
rect 1479 2573 1483 2574
rect 1607 2578 1611 2579
rect 1607 2573 1611 2574
rect 1352 2557 1354 2573
rect 1480 2557 1482 2573
rect 1608 2557 1610 2573
rect 1350 2556 1356 2557
rect 1350 2552 1351 2556
rect 1355 2552 1356 2556
rect 1350 2551 1356 2552
rect 1478 2556 1484 2557
rect 1478 2552 1479 2556
rect 1483 2552 1484 2556
rect 1478 2551 1484 2552
rect 1606 2556 1612 2557
rect 1606 2552 1607 2556
rect 1611 2552 1612 2556
rect 1606 2551 1612 2552
rect 846 2547 852 2548
rect 846 2543 847 2547
rect 851 2543 852 2547
rect 846 2542 852 2543
rect 950 2547 956 2548
rect 950 2543 951 2547
rect 955 2543 956 2547
rect 950 2542 956 2543
rect 1062 2547 1068 2548
rect 1062 2543 1063 2547
rect 1067 2543 1068 2547
rect 1062 2542 1068 2543
rect 1174 2547 1180 2548
rect 1174 2543 1175 2547
rect 1179 2543 1180 2547
rect 1174 2542 1180 2543
rect 1294 2547 1300 2548
rect 1294 2543 1295 2547
rect 1299 2543 1300 2547
rect 1294 2542 1300 2543
rect 1422 2547 1428 2548
rect 1422 2543 1423 2547
rect 1427 2543 1428 2547
rect 1422 2542 1428 2543
rect 1430 2547 1436 2548
rect 1430 2543 1431 2547
rect 1435 2543 1436 2547
rect 1430 2542 1436 2543
rect 1558 2547 1564 2548
rect 1558 2543 1559 2547
rect 1563 2543 1564 2547
rect 1558 2542 1564 2543
rect 848 2520 850 2542
rect 878 2537 884 2538
rect 878 2533 879 2537
rect 883 2533 884 2537
rect 878 2532 884 2533
rect 846 2519 852 2520
rect 846 2515 847 2519
rect 851 2515 852 2519
rect 846 2514 852 2515
rect 822 2511 828 2512
rect 822 2507 823 2511
rect 827 2507 828 2511
rect 880 2507 882 2532
rect 952 2520 954 2542
rect 990 2537 996 2538
rect 990 2533 991 2537
rect 995 2533 996 2537
rect 990 2532 996 2533
rect 950 2519 956 2520
rect 950 2515 951 2519
rect 955 2515 956 2519
rect 950 2514 956 2515
rect 992 2507 994 2532
rect 1064 2520 1066 2542
rect 1102 2537 1108 2538
rect 1102 2533 1103 2537
rect 1107 2533 1108 2537
rect 1102 2532 1108 2533
rect 1062 2519 1068 2520
rect 1062 2515 1063 2519
rect 1067 2515 1068 2519
rect 1062 2514 1068 2515
rect 1104 2507 1106 2532
rect 1176 2520 1178 2542
rect 1222 2537 1228 2538
rect 1222 2533 1223 2537
rect 1227 2533 1228 2537
rect 1222 2532 1228 2533
rect 1350 2537 1356 2538
rect 1350 2533 1351 2537
rect 1355 2533 1356 2537
rect 1350 2532 1356 2533
rect 1174 2519 1180 2520
rect 1174 2515 1175 2519
rect 1179 2515 1180 2519
rect 1174 2514 1180 2515
rect 1224 2507 1226 2532
rect 1352 2507 1354 2532
rect 111 2506 115 2507
rect 111 2501 115 2502
rect 503 2506 507 2507
rect 503 2501 507 2502
rect 551 2506 555 2507
rect 551 2501 555 2502
rect 591 2506 595 2507
rect 591 2501 595 2502
rect 679 2506 683 2507
rect 679 2501 683 2502
rect 735 2506 739 2507
rect 735 2501 739 2502
rect 775 2506 779 2507
rect 822 2506 828 2507
rect 879 2506 883 2507
rect 775 2501 779 2502
rect 879 2501 883 2502
rect 911 2506 915 2507
rect 911 2501 915 2502
rect 991 2506 995 2507
rect 991 2501 995 2502
rect 1079 2506 1083 2507
rect 1079 2501 1083 2502
rect 1103 2506 1107 2507
rect 1103 2501 1107 2502
rect 1223 2506 1227 2507
rect 1223 2501 1227 2502
rect 1239 2506 1243 2507
rect 1239 2501 1243 2502
rect 1351 2506 1355 2507
rect 1351 2501 1355 2502
rect 1399 2506 1403 2507
rect 1399 2501 1403 2502
rect 112 2485 114 2501
rect 110 2484 116 2485
rect 552 2484 554 2501
rect 630 2499 636 2500
rect 630 2495 631 2499
rect 635 2495 636 2499
rect 630 2494 636 2495
rect 110 2480 111 2484
rect 115 2480 116 2484
rect 110 2479 116 2480
rect 550 2483 556 2484
rect 550 2479 551 2483
rect 555 2479 556 2483
rect 550 2478 556 2479
rect 632 2476 634 2494
rect 736 2484 738 2501
rect 814 2499 820 2500
rect 814 2495 815 2499
rect 819 2495 820 2499
rect 814 2494 820 2495
rect 734 2483 740 2484
rect 734 2479 735 2483
rect 739 2479 740 2483
rect 734 2478 740 2479
rect 816 2476 818 2494
rect 912 2484 914 2501
rect 990 2495 996 2496
rect 990 2491 991 2495
rect 995 2491 996 2495
rect 990 2490 996 2491
rect 910 2483 916 2484
rect 910 2479 911 2483
rect 915 2479 916 2483
rect 910 2478 916 2479
rect 630 2475 636 2476
rect 622 2471 628 2472
rect 110 2467 116 2468
rect 110 2463 111 2467
rect 115 2463 116 2467
rect 622 2467 623 2471
rect 627 2467 628 2471
rect 630 2471 631 2475
rect 635 2471 636 2475
rect 630 2470 636 2471
rect 814 2475 820 2476
rect 814 2471 815 2475
rect 819 2471 820 2475
rect 814 2470 820 2471
rect 622 2466 628 2467
rect 110 2462 116 2463
rect 550 2464 556 2465
rect 112 2443 114 2462
rect 550 2460 551 2464
rect 555 2460 556 2464
rect 550 2459 556 2460
rect 552 2443 554 2459
rect 111 2442 115 2443
rect 111 2437 115 2438
rect 415 2442 419 2443
rect 415 2437 419 2438
rect 503 2442 507 2443
rect 503 2437 507 2438
rect 551 2442 555 2443
rect 551 2437 555 2438
rect 599 2442 603 2443
rect 599 2437 603 2438
rect 112 2418 114 2437
rect 416 2421 418 2437
rect 504 2421 506 2437
rect 600 2421 602 2437
rect 414 2420 420 2421
rect 110 2417 116 2418
rect 110 2413 111 2417
rect 115 2413 116 2417
rect 414 2416 415 2420
rect 419 2416 420 2420
rect 414 2415 420 2416
rect 502 2420 508 2421
rect 502 2416 503 2420
rect 507 2416 508 2420
rect 502 2415 508 2416
rect 598 2420 604 2421
rect 598 2416 599 2420
rect 603 2416 604 2420
rect 598 2415 604 2416
rect 110 2412 116 2413
rect 486 2411 492 2412
rect 486 2407 487 2411
rect 491 2407 492 2411
rect 486 2406 492 2407
rect 574 2411 580 2412
rect 574 2407 575 2411
rect 579 2407 580 2411
rect 574 2406 580 2407
rect 582 2411 588 2412
rect 582 2407 583 2411
rect 587 2407 588 2411
rect 582 2406 588 2407
rect 414 2401 420 2402
rect 110 2400 116 2401
rect 110 2396 111 2400
rect 115 2396 116 2400
rect 414 2397 415 2401
rect 419 2397 420 2401
rect 414 2396 420 2397
rect 110 2395 116 2396
rect 112 2375 114 2395
rect 416 2375 418 2396
rect 488 2384 490 2406
rect 502 2401 508 2402
rect 502 2397 503 2401
rect 507 2397 508 2401
rect 502 2396 508 2397
rect 486 2383 492 2384
rect 486 2379 487 2383
rect 491 2379 492 2383
rect 486 2378 492 2379
rect 504 2375 506 2396
rect 111 2374 115 2375
rect 111 2369 115 2370
rect 319 2374 323 2375
rect 319 2369 323 2370
rect 415 2374 419 2375
rect 415 2369 419 2370
rect 431 2374 435 2375
rect 431 2369 435 2370
rect 503 2374 507 2375
rect 503 2369 507 2370
rect 543 2374 547 2375
rect 543 2369 547 2370
rect 112 2353 114 2369
rect 110 2352 116 2353
rect 320 2352 322 2369
rect 398 2367 404 2368
rect 398 2363 399 2367
rect 403 2363 404 2367
rect 398 2362 404 2363
rect 110 2348 111 2352
rect 115 2348 116 2352
rect 110 2347 116 2348
rect 318 2351 324 2352
rect 318 2347 319 2351
rect 323 2347 324 2351
rect 318 2346 324 2347
rect 400 2344 402 2362
rect 432 2352 434 2369
rect 544 2352 546 2369
rect 576 2368 578 2406
rect 584 2376 586 2406
rect 598 2401 604 2402
rect 598 2397 599 2401
rect 603 2397 604 2401
rect 598 2396 604 2397
rect 582 2375 588 2376
rect 600 2375 602 2396
rect 624 2384 626 2466
rect 734 2464 740 2465
rect 734 2460 735 2464
rect 739 2460 740 2464
rect 734 2459 740 2460
rect 910 2464 916 2465
rect 910 2460 911 2464
rect 915 2460 916 2464
rect 910 2459 916 2460
rect 736 2443 738 2459
rect 912 2443 914 2459
rect 703 2442 707 2443
rect 703 2437 707 2438
rect 735 2442 739 2443
rect 735 2437 739 2438
rect 807 2442 811 2443
rect 807 2437 811 2438
rect 911 2442 915 2443
rect 911 2437 915 2438
rect 919 2442 923 2443
rect 919 2437 923 2438
rect 704 2421 706 2437
rect 808 2421 810 2437
rect 920 2421 922 2437
rect 702 2420 708 2421
rect 702 2416 703 2420
rect 707 2416 708 2420
rect 702 2415 708 2416
rect 806 2420 812 2421
rect 806 2416 807 2420
rect 811 2416 812 2420
rect 806 2415 812 2416
rect 918 2420 924 2421
rect 918 2416 919 2420
rect 923 2416 924 2420
rect 918 2415 924 2416
rect 992 2412 994 2490
rect 1080 2484 1082 2501
rect 1240 2484 1242 2501
rect 1400 2484 1402 2501
rect 1424 2500 1426 2542
rect 1432 2520 1434 2542
rect 1478 2537 1484 2538
rect 1478 2533 1479 2537
rect 1483 2533 1484 2537
rect 1478 2532 1484 2533
rect 1430 2519 1436 2520
rect 1430 2515 1431 2519
rect 1435 2515 1436 2519
rect 1430 2514 1436 2515
rect 1480 2507 1482 2532
rect 1560 2520 1562 2542
rect 1606 2537 1612 2538
rect 1606 2533 1607 2537
rect 1611 2533 1612 2537
rect 1606 2532 1612 2533
rect 1558 2519 1564 2520
rect 1558 2515 1559 2519
rect 1563 2515 1564 2519
rect 1558 2514 1564 2515
rect 1518 2507 1524 2508
rect 1608 2507 1610 2532
rect 1680 2520 1682 2610
rect 1766 2607 1767 2611
rect 1771 2607 1772 2611
rect 1766 2606 1772 2607
rect 1806 2611 1812 2612
rect 1806 2607 1807 2611
rect 1811 2607 1812 2611
rect 1806 2606 1812 2607
rect 1870 2608 1876 2609
rect 1768 2579 1770 2606
rect 1767 2578 1771 2579
rect 1808 2575 1810 2606
rect 1870 2604 1871 2608
rect 1875 2604 1876 2608
rect 1870 2603 1876 2604
rect 1872 2575 1874 2603
rect 1767 2573 1771 2574
rect 1807 2574 1811 2575
rect 1768 2554 1770 2573
rect 1807 2569 1811 2570
rect 1831 2574 1835 2575
rect 1831 2569 1835 2570
rect 1871 2574 1875 2575
rect 1871 2569 1875 2570
rect 1766 2553 1772 2554
rect 1766 2549 1767 2553
rect 1771 2549 1772 2553
rect 1808 2550 1810 2569
rect 1832 2553 1834 2569
rect 1830 2552 1836 2553
rect 1766 2548 1772 2549
rect 1806 2549 1812 2550
rect 1806 2545 1807 2549
rect 1811 2545 1812 2549
rect 1830 2548 1831 2552
rect 1835 2548 1836 2552
rect 1830 2547 1836 2548
rect 1806 2544 1812 2545
rect 1904 2544 1906 2638
rect 1944 2620 1946 2638
rect 1968 2628 1970 2645
rect 2062 2643 2068 2644
rect 2062 2639 2063 2643
rect 2067 2639 2068 2643
rect 2062 2638 2068 2639
rect 1966 2627 1972 2628
rect 1966 2623 1967 2627
rect 1971 2623 1972 2627
rect 1966 2622 1972 2623
rect 2064 2620 2066 2638
rect 2072 2628 2074 2645
rect 2142 2643 2148 2644
rect 2142 2639 2143 2643
rect 2147 2639 2148 2643
rect 2142 2638 2148 2639
rect 2070 2627 2076 2628
rect 2070 2623 2071 2627
rect 2075 2623 2076 2627
rect 2070 2622 2076 2623
rect 2144 2620 2146 2638
rect 2184 2628 2186 2645
rect 2254 2643 2260 2644
rect 2254 2639 2255 2643
rect 2259 2639 2260 2643
rect 2254 2638 2260 2639
rect 2182 2627 2188 2628
rect 2182 2623 2183 2627
rect 2187 2623 2188 2627
rect 2182 2622 2188 2623
rect 2256 2620 2258 2638
rect 2264 2620 2266 2654
rect 2280 2651 2282 2680
rect 2352 2668 2354 2690
rect 2406 2685 2412 2686
rect 2406 2681 2407 2685
rect 2411 2681 2412 2685
rect 2406 2680 2412 2681
rect 2542 2685 2548 2686
rect 2542 2681 2543 2685
rect 2547 2681 2548 2685
rect 2542 2680 2548 2681
rect 2350 2667 2356 2668
rect 2350 2663 2351 2667
rect 2355 2663 2356 2667
rect 2350 2662 2356 2663
rect 2408 2651 2410 2680
rect 2544 2651 2546 2680
rect 2616 2668 2618 2690
rect 2686 2685 2692 2686
rect 2686 2681 2687 2685
rect 2691 2681 2692 2685
rect 2686 2680 2692 2681
rect 2614 2667 2620 2668
rect 2614 2663 2615 2667
rect 2619 2663 2620 2667
rect 2614 2662 2620 2663
rect 2688 2651 2690 2680
rect 2279 2650 2283 2651
rect 2279 2645 2283 2646
rect 2295 2650 2299 2651
rect 2295 2645 2299 2646
rect 2407 2650 2411 2651
rect 2407 2645 2411 2646
rect 2431 2650 2435 2651
rect 2431 2645 2435 2646
rect 2543 2650 2547 2651
rect 2543 2645 2547 2646
rect 2583 2650 2587 2651
rect 2583 2645 2587 2646
rect 2687 2650 2691 2651
rect 2687 2645 2691 2646
rect 2759 2650 2763 2651
rect 2759 2645 2763 2646
rect 2296 2628 2298 2645
rect 2432 2628 2434 2645
rect 2510 2643 2516 2644
rect 2510 2639 2511 2643
rect 2515 2639 2516 2643
rect 2510 2638 2516 2639
rect 2294 2627 2300 2628
rect 2294 2623 2295 2627
rect 2299 2623 2300 2627
rect 2294 2622 2300 2623
rect 2430 2627 2436 2628
rect 2430 2623 2431 2627
rect 2435 2623 2436 2627
rect 2430 2622 2436 2623
rect 2512 2620 2514 2638
rect 2584 2628 2586 2645
rect 2760 2628 2762 2645
rect 2768 2644 2770 2690
rect 2776 2660 2778 2690
rect 2846 2685 2852 2686
rect 2846 2681 2847 2685
rect 2851 2681 2852 2685
rect 2846 2680 2852 2681
rect 2774 2659 2780 2660
rect 2774 2655 2775 2659
rect 2779 2655 2780 2659
rect 2774 2654 2780 2655
rect 2848 2651 2850 2680
rect 2984 2668 2986 2766
rect 3070 2764 3076 2765
rect 3070 2760 3071 2764
rect 3075 2760 3076 2764
rect 3070 2759 3076 2760
rect 3230 2764 3236 2765
rect 3230 2760 3231 2764
rect 3235 2760 3236 2764
rect 3230 2759 3236 2760
rect 3072 2727 3074 2759
rect 3232 2727 3234 2759
rect 3023 2726 3027 2727
rect 3023 2721 3027 2722
rect 3071 2726 3075 2727
rect 3071 2721 3075 2722
rect 3207 2726 3211 2727
rect 3207 2721 3211 2722
rect 3231 2726 3235 2727
rect 3231 2721 3235 2722
rect 3024 2705 3026 2721
rect 3208 2705 3210 2721
rect 3022 2704 3028 2705
rect 3022 2700 3023 2704
rect 3027 2700 3028 2704
rect 3022 2699 3028 2700
rect 3206 2704 3212 2705
rect 3206 2700 3207 2704
rect 3211 2700 3212 2704
rect 3206 2699 3212 2700
rect 3094 2695 3100 2696
rect 3094 2691 3095 2695
rect 3099 2691 3100 2695
rect 3094 2690 3100 2691
rect 3102 2695 3108 2696
rect 3102 2691 3103 2695
rect 3107 2691 3108 2695
rect 3102 2690 3108 2691
rect 3022 2685 3028 2686
rect 3022 2681 3023 2685
rect 3027 2681 3028 2685
rect 3022 2680 3028 2681
rect 2982 2667 2988 2668
rect 2982 2663 2983 2667
rect 2987 2663 2988 2667
rect 2982 2662 2988 2663
rect 3024 2651 3026 2680
rect 3096 2668 3098 2690
rect 3094 2667 3100 2668
rect 3094 2663 3095 2667
rect 3099 2663 3100 2667
rect 3094 2662 3100 2663
rect 3104 2660 3106 2690
rect 3206 2685 3212 2686
rect 3206 2681 3207 2685
rect 3211 2681 3212 2685
rect 3206 2680 3212 2681
rect 3102 2659 3108 2660
rect 3102 2655 3103 2659
rect 3107 2655 3108 2659
rect 3102 2654 3108 2655
rect 3138 2651 3144 2652
rect 3208 2651 3210 2680
rect 2847 2650 2851 2651
rect 2847 2645 2851 2646
rect 2959 2650 2963 2651
rect 2959 2645 2963 2646
rect 3023 2650 3027 2651
rect 3138 2647 3139 2651
rect 3143 2647 3144 2651
rect 3138 2646 3144 2647
rect 3167 2650 3171 2651
rect 3023 2645 3027 2646
rect 2766 2643 2772 2644
rect 2766 2639 2767 2643
rect 2771 2639 2772 2643
rect 2766 2638 2772 2639
rect 2830 2643 2836 2644
rect 2830 2639 2831 2643
rect 2835 2639 2836 2643
rect 2830 2638 2836 2639
rect 2582 2627 2588 2628
rect 2582 2623 2583 2627
rect 2587 2623 2588 2627
rect 2582 2622 2588 2623
rect 2758 2627 2764 2628
rect 2758 2623 2759 2627
rect 2763 2623 2764 2627
rect 2758 2622 2764 2623
rect 2832 2620 2834 2638
rect 2960 2628 2962 2645
rect 3030 2643 3036 2644
rect 3030 2639 3031 2643
rect 3035 2639 3036 2643
rect 3030 2638 3036 2639
rect 2958 2627 2964 2628
rect 2958 2623 2959 2627
rect 2963 2623 2964 2627
rect 2958 2622 2964 2623
rect 3032 2620 3034 2638
rect 3140 2620 3142 2646
rect 3167 2645 3171 2646
rect 3207 2650 3211 2651
rect 3207 2645 3211 2646
rect 3168 2628 3170 2645
rect 3166 2627 3172 2628
rect 3166 2623 3167 2627
rect 3171 2623 3172 2627
rect 3166 2622 3172 2623
rect 1942 2619 1948 2620
rect 1942 2615 1943 2619
rect 1947 2615 1948 2619
rect 1942 2614 1948 2615
rect 2062 2619 2068 2620
rect 2062 2615 2063 2619
rect 2067 2615 2068 2619
rect 2062 2614 2068 2615
rect 2142 2619 2148 2620
rect 2142 2615 2143 2619
rect 2147 2615 2148 2619
rect 2142 2614 2148 2615
rect 2254 2619 2260 2620
rect 2254 2615 2255 2619
rect 2259 2615 2260 2619
rect 2254 2614 2260 2615
rect 2262 2619 2268 2620
rect 2262 2615 2263 2619
rect 2267 2615 2268 2619
rect 2262 2614 2268 2615
rect 2394 2619 2400 2620
rect 2394 2615 2395 2619
rect 2399 2615 2400 2619
rect 2394 2614 2400 2615
rect 2510 2619 2516 2620
rect 2510 2615 2511 2619
rect 2515 2615 2516 2619
rect 2510 2614 2516 2615
rect 2830 2619 2836 2620
rect 2830 2615 2831 2619
rect 2835 2615 2836 2619
rect 2830 2614 2836 2615
rect 3030 2619 3036 2620
rect 3030 2615 3031 2619
rect 3035 2615 3036 2619
rect 3030 2614 3036 2615
rect 3138 2619 3144 2620
rect 3138 2615 3139 2619
rect 3143 2615 3144 2619
rect 3138 2614 3144 2615
rect 1966 2608 1972 2609
rect 1966 2604 1967 2608
rect 1971 2604 1972 2608
rect 1966 2603 1972 2604
rect 2070 2608 2076 2609
rect 2070 2604 2071 2608
rect 2075 2604 2076 2608
rect 2070 2603 2076 2604
rect 2182 2608 2188 2609
rect 2182 2604 2183 2608
rect 2187 2604 2188 2608
rect 2182 2603 2188 2604
rect 2294 2608 2300 2609
rect 2294 2604 2295 2608
rect 2299 2604 2300 2608
rect 2294 2603 2300 2604
rect 1968 2575 1970 2603
rect 2072 2575 2074 2603
rect 2184 2575 2186 2603
rect 2296 2575 2298 2603
rect 1919 2574 1923 2575
rect 1919 2569 1923 2570
rect 1967 2574 1971 2575
rect 1967 2569 1971 2570
rect 2007 2574 2011 2575
rect 2007 2569 2011 2570
rect 2071 2574 2075 2575
rect 2071 2569 2075 2570
rect 2111 2574 2115 2575
rect 2111 2569 2115 2570
rect 2183 2574 2187 2575
rect 2183 2569 2187 2570
rect 2223 2574 2227 2575
rect 2223 2569 2227 2570
rect 2295 2574 2299 2575
rect 2295 2569 2299 2570
rect 2343 2574 2347 2575
rect 2343 2569 2347 2570
rect 1920 2553 1922 2569
rect 2008 2553 2010 2569
rect 2112 2553 2114 2569
rect 2224 2553 2226 2569
rect 2344 2553 2346 2569
rect 1918 2552 1924 2553
rect 1918 2548 1919 2552
rect 1923 2548 1924 2552
rect 1918 2547 1924 2548
rect 2006 2552 2012 2553
rect 2006 2548 2007 2552
rect 2011 2548 2012 2552
rect 2006 2547 2012 2548
rect 2110 2552 2116 2553
rect 2110 2548 2111 2552
rect 2115 2548 2116 2552
rect 2110 2547 2116 2548
rect 2222 2552 2228 2553
rect 2222 2548 2223 2552
rect 2227 2548 2228 2552
rect 2222 2547 2228 2548
rect 2342 2552 2348 2553
rect 2342 2548 2343 2552
rect 2347 2548 2348 2552
rect 2342 2547 2348 2548
rect 1902 2543 1908 2544
rect 1902 2539 1903 2543
rect 1907 2539 1908 2543
rect 1902 2538 1908 2539
rect 1910 2543 1916 2544
rect 1910 2539 1911 2543
rect 1915 2539 1916 2543
rect 1910 2538 1916 2539
rect 2086 2543 2092 2544
rect 2086 2539 2087 2543
rect 2091 2539 2092 2543
rect 2086 2538 2092 2539
rect 2190 2543 2196 2544
rect 2190 2539 2191 2543
rect 2195 2539 2196 2543
rect 2190 2538 2196 2539
rect 1766 2536 1772 2537
rect 1766 2532 1767 2536
rect 1771 2532 1772 2536
rect 1830 2533 1836 2534
rect 1766 2531 1772 2532
rect 1806 2532 1812 2533
rect 1678 2519 1684 2520
rect 1678 2515 1679 2519
rect 1683 2515 1684 2519
rect 1678 2514 1684 2515
rect 1768 2507 1770 2531
rect 1806 2528 1807 2532
rect 1811 2528 1812 2532
rect 1830 2529 1831 2533
rect 1835 2529 1836 2533
rect 1830 2528 1836 2529
rect 1806 2527 1812 2528
rect 1808 2511 1810 2527
rect 1832 2511 1834 2528
rect 1912 2516 1914 2538
rect 1918 2533 1924 2534
rect 1918 2529 1919 2533
rect 1923 2529 1924 2533
rect 1918 2528 1924 2529
rect 2006 2533 2012 2534
rect 2006 2529 2007 2533
rect 2011 2529 2012 2533
rect 2006 2528 2012 2529
rect 1910 2515 1916 2516
rect 1910 2511 1911 2515
rect 1915 2511 1916 2515
rect 1920 2511 1922 2528
rect 2008 2511 2010 2528
rect 2088 2516 2090 2538
rect 2110 2533 2116 2534
rect 2110 2529 2111 2533
rect 2115 2529 2116 2533
rect 2110 2528 2116 2529
rect 2086 2515 2092 2516
rect 2086 2511 2087 2515
rect 2091 2511 2092 2515
rect 2112 2511 2114 2528
rect 2192 2516 2194 2538
rect 2222 2533 2228 2534
rect 2222 2529 2223 2533
rect 2227 2529 2228 2533
rect 2222 2528 2228 2529
rect 2342 2533 2348 2534
rect 2342 2529 2343 2533
rect 2347 2529 2348 2533
rect 2342 2528 2348 2529
rect 2190 2515 2196 2516
rect 2190 2511 2191 2515
rect 2195 2511 2196 2515
rect 1807 2510 1811 2511
rect 1479 2506 1483 2507
rect 1518 2503 1519 2507
rect 1523 2503 1524 2507
rect 1518 2502 1524 2503
rect 1567 2506 1571 2507
rect 1479 2501 1483 2502
rect 1422 2499 1428 2500
rect 1422 2495 1423 2499
rect 1427 2495 1428 2499
rect 1422 2494 1428 2495
rect 1470 2499 1476 2500
rect 1470 2495 1471 2499
rect 1475 2495 1476 2499
rect 1470 2494 1476 2495
rect 1078 2483 1084 2484
rect 1078 2479 1079 2483
rect 1083 2479 1084 2483
rect 1078 2478 1084 2479
rect 1238 2483 1244 2484
rect 1238 2479 1239 2483
rect 1243 2479 1244 2483
rect 1238 2478 1244 2479
rect 1398 2483 1404 2484
rect 1398 2479 1399 2483
rect 1403 2479 1404 2483
rect 1398 2478 1404 2479
rect 1472 2476 1474 2494
rect 1520 2476 1522 2502
rect 1567 2501 1571 2502
rect 1607 2506 1611 2507
rect 1607 2501 1611 2502
rect 1767 2506 1771 2507
rect 1807 2505 1811 2506
rect 1831 2510 1835 2511
rect 1910 2510 1916 2511
rect 1919 2510 1923 2511
rect 1831 2505 1835 2506
rect 1919 2505 1923 2506
rect 1951 2510 1955 2511
rect 1951 2505 1955 2506
rect 2007 2510 2011 2511
rect 2007 2505 2011 2506
rect 2039 2510 2043 2511
rect 2086 2510 2092 2511
rect 2111 2510 2115 2511
rect 2039 2505 2043 2506
rect 2111 2505 2115 2506
rect 2135 2510 2139 2511
rect 2190 2510 2196 2511
rect 2206 2515 2212 2516
rect 2206 2511 2207 2515
rect 2211 2511 2212 2515
rect 2224 2511 2226 2528
rect 2344 2511 2346 2528
rect 2396 2516 2398 2614
rect 2430 2608 2436 2609
rect 2430 2604 2431 2608
rect 2435 2604 2436 2608
rect 2430 2603 2436 2604
rect 2582 2608 2588 2609
rect 2582 2604 2583 2608
rect 2587 2604 2588 2608
rect 2582 2603 2588 2604
rect 2758 2608 2764 2609
rect 2758 2604 2759 2608
rect 2763 2604 2764 2608
rect 2758 2603 2764 2604
rect 2958 2608 2964 2609
rect 2958 2604 2959 2608
rect 2963 2604 2964 2608
rect 2958 2603 2964 2604
rect 3166 2608 3172 2609
rect 3166 2604 3167 2608
rect 3171 2604 3172 2608
rect 3166 2603 3172 2604
rect 2432 2575 2434 2603
rect 2584 2575 2586 2603
rect 2760 2575 2762 2603
rect 2960 2575 2962 2603
rect 3168 2575 3170 2603
rect 2431 2574 2435 2575
rect 2431 2569 2435 2570
rect 2487 2574 2491 2575
rect 2487 2569 2491 2570
rect 2583 2574 2587 2575
rect 2583 2569 2587 2570
rect 2647 2574 2651 2575
rect 2647 2569 2651 2570
rect 2759 2574 2763 2575
rect 2759 2569 2763 2570
rect 2815 2574 2819 2575
rect 2815 2569 2819 2570
rect 2959 2574 2963 2575
rect 2959 2569 2963 2570
rect 2999 2574 3003 2575
rect 2999 2569 3003 2570
rect 3167 2574 3171 2575
rect 3167 2569 3171 2570
rect 3191 2574 3195 2575
rect 3191 2569 3195 2570
rect 2488 2553 2490 2569
rect 2578 2559 2584 2560
rect 2578 2555 2579 2559
rect 2583 2555 2584 2559
rect 2578 2554 2584 2555
rect 2486 2552 2492 2553
rect 2486 2548 2487 2552
rect 2491 2548 2492 2552
rect 2486 2547 2492 2548
rect 2414 2543 2420 2544
rect 2414 2539 2415 2543
rect 2419 2539 2420 2543
rect 2414 2538 2420 2539
rect 2558 2543 2564 2544
rect 2558 2539 2559 2543
rect 2563 2539 2564 2543
rect 2558 2538 2564 2539
rect 2416 2516 2418 2538
rect 2486 2533 2492 2534
rect 2486 2529 2487 2533
rect 2491 2529 2492 2533
rect 2486 2528 2492 2529
rect 2394 2515 2400 2516
rect 2394 2511 2395 2515
rect 2399 2511 2400 2515
rect 2206 2510 2212 2511
rect 2223 2510 2227 2511
rect 2135 2505 2139 2506
rect 1767 2501 1771 2502
rect 1568 2484 1570 2501
rect 1768 2485 1770 2501
rect 1808 2489 1810 2505
rect 1806 2488 1812 2489
rect 1952 2488 1954 2505
rect 2014 2503 2020 2504
rect 2014 2498 2015 2503
rect 2019 2498 2020 2503
rect 2022 2503 2028 2504
rect 2022 2499 2023 2503
rect 2027 2499 2028 2503
rect 2022 2498 2028 2499
rect 2015 2495 2019 2496
rect 1766 2484 1772 2485
rect 1566 2483 1572 2484
rect 1566 2479 1567 2483
rect 1571 2479 1572 2483
rect 1766 2480 1767 2484
rect 1771 2480 1772 2484
rect 1806 2484 1807 2488
rect 1811 2484 1812 2488
rect 1806 2483 1812 2484
rect 1950 2487 1956 2488
rect 1950 2483 1951 2487
rect 1955 2483 1956 2487
rect 1950 2482 1956 2483
rect 2024 2480 2026 2498
rect 2040 2488 2042 2505
rect 2136 2488 2138 2505
rect 2038 2487 2044 2488
rect 2038 2483 2039 2487
rect 2043 2483 2044 2487
rect 2038 2482 2044 2483
rect 2134 2487 2140 2488
rect 2134 2483 2135 2487
rect 2139 2483 2140 2487
rect 2134 2482 2140 2483
rect 2208 2480 2210 2510
rect 2223 2505 2227 2506
rect 2239 2510 2243 2511
rect 2239 2505 2243 2506
rect 2343 2510 2347 2511
rect 2343 2505 2347 2506
rect 2367 2510 2371 2511
rect 2394 2510 2400 2511
rect 2414 2515 2420 2516
rect 2414 2511 2415 2515
rect 2419 2511 2420 2515
rect 2488 2511 2490 2528
rect 2560 2516 2562 2538
rect 2558 2515 2564 2516
rect 2558 2511 2559 2515
rect 2563 2511 2564 2515
rect 2414 2510 2420 2511
rect 2487 2510 2491 2511
rect 2367 2505 2371 2506
rect 2487 2505 2491 2506
rect 2527 2510 2531 2511
rect 2558 2510 2564 2511
rect 2527 2505 2531 2506
rect 2215 2500 2219 2501
rect 2215 2495 2219 2496
rect 2216 2480 2218 2495
rect 2240 2488 2242 2505
rect 2318 2503 2324 2504
rect 2318 2499 2319 2503
rect 2323 2499 2324 2503
rect 2318 2498 2324 2499
rect 2238 2487 2244 2488
rect 2238 2483 2239 2487
rect 2243 2483 2244 2487
rect 2238 2482 2244 2483
rect 2320 2480 2322 2498
rect 2368 2488 2370 2505
rect 2374 2503 2380 2504
rect 2374 2499 2375 2503
rect 2379 2499 2380 2503
rect 2374 2498 2380 2499
rect 2366 2487 2372 2488
rect 2366 2483 2367 2487
rect 2371 2483 2372 2487
rect 2366 2482 2372 2483
rect 1766 2479 1772 2480
rect 2022 2479 2028 2480
rect 1566 2478 1572 2479
rect 1470 2475 1476 2476
rect 1150 2471 1156 2472
rect 1150 2467 1151 2471
rect 1155 2467 1156 2471
rect 1470 2471 1471 2475
rect 1475 2471 1476 2475
rect 1470 2470 1476 2471
rect 1518 2475 1524 2476
rect 1518 2471 1519 2475
rect 1523 2471 1524 2475
rect 2022 2475 2023 2479
rect 2027 2475 2028 2479
rect 2022 2474 2028 2475
rect 2206 2479 2212 2480
rect 2206 2475 2207 2479
rect 2211 2475 2212 2479
rect 2206 2474 2212 2475
rect 2214 2479 2220 2480
rect 2214 2475 2215 2479
rect 2219 2475 2220 2479
rect 2214 2474 2220 2475
rect 2318 2479 2324 2480
rect 2318 2475 2319 2479
rect 2323 2475 2324 2479
rect 2318 2474 2324 2475
rect 1518 2470 1524 2471
rect 1806 2471 1812 2472
rect 1150 2466 1156 2467
rect 1766 2467 1772 2468
rect 1078 2464 1084 2465
rect 1078 2460 1079 2464
rect 1083 2460 1084 2464
rect 1078 2459 1084 2460
rect 1080 2443 1082 2459
rect 1039 2442 1043 2443
rect 1039 2437 1043 2438
rect 1079 2442 1083 2443
rect 1079 2437 1083 2438
rect 1040 2421 1042 2437
rect 1038 2420 1044 2421
rect 1038 2416 1039 2420
rect 1043 2416 1044 2420
rect 1038 2415 1044 2416
rect 774 2411 780 2412
rect 774 2407 775 2411
rect 779 2407 780 2411
rect 774 2406 780 2407
rect 878 2411 884 2412
rect 878 2407 879 2411
rect 883 2407 884 2411
rect 878 2406 884 2407
rect 990 2411 996 2412
rect 990 2407 991 2411
rect 995 2407 996 2411
rect 990 2406 996 2407
rect 998 2411 1004 2412
rect 998 2407 999 2411
rect 1003 2407 1004 2411
rect 998 2406 1004 2407
rect 702 2401 708 2402
rect 702 2397 703 2401
rect 707 2397 708 2401
rect 702 2396 708 2397
rect 622 2383 628 2384
rect 622 2379 623 2383
rect 627 2379 628 2383
rect 622 2378 628 2379
rect 704 2375 706 2396
rect 776 2384 778 2406
rect 806 2401 812 2402
rect 806 2397 807 2401
rect 811 2397 812 2401
rect 806 2396 812 2397
rect 774 2383 780 2384
rect 774 2379 775 2383
rect 779 2379 780 2383
rect 774 2378 780 2379
rect 808 2375 810 2396
rect 880 2384 882 2406
rect 918 2401 924 2402
rect 918 2397 919 2401
rect 923 2397 924 2401
rect 918 2396 924 2397
rect 878 2383 884 2384
rect 878 2379 879 2383
rect 883 2379 884 2383
rect 878 2378 884 2379
rect 920 2375 922 2396
rect 1000 2376 1002 2406
rect 1038 2401 1044 2402
rect 1038 2397 1039 2401
rect 1043 2397 1044 2401
rect 1038 2396 1044 2397
rect 998 2375 1004 2376
rect 1040 2375 1042 2396
rect 1152 2384 1154 2466
rect 1238 2464 1244 2465
rect 1238 2460 1239 2464
rect 1243 2460 1244 2464
rect 1238 2459 1244 2460
rect 1398 2464 1404 2465
rect 1398 2460 1399 2464
rect 1403 2460 1404 2464
rect 1398 2459 1404 2460
rect 1566 2464 1572 2465
rect 1566 2460 1567 2464
rect 1571 2460 1572 2464
rect 1766 2463 1767 2467
rect 1771 2463 1772 2467
rect 1806 2467 1807 2471
rect 1811 2467 1812 2471
rect 1806 2466 1812 2467
rect 1950 2468 1956 2469
rect 1766 2462 1772 2463
rect 1566 2459 1572 2460
rect 1240 2443 1242 2459
rect 1400 2443 1402 2459
rect 1568 2443 1570 2459
rect 1768 2443 1770 2462
rect 1167 2442 1171 2443
rect 1167 2437 1171 2438
rect 1239 2442 1243 2443
rect 1239 2437 1243 2438
rect 1295 2442 1299 2443
rect 1295 2437 1299 2438
rect 1399 2442 1403 2443
rect 1399 2437 1403 2438
rect 1423 2442 1427 2443
rect 1423 2437 1427 2438
rect 1567 2442 1571 2443
rect 1567 2437 1571 2438
rect 1767 2442 1771 2443
rect 1808 2439 1810 2466
rect 1950 2464 1951 2468
rect 1955 2464 1956 2468
rect 1950 2463 1956 2464
rect 2038 2468 2044 2469
rect 2038 2464 2039 2468
rect 2043 2464 2044 2468
rect 2038 2463 2044 2464
rect 2134 2468 2140 2469
rect 2134 2464 2135 2468
rect 2139 2464 2140 2468
rect 2134 2463 2140 2464
rect 2238 2468 2244 2469
rect 2238 2464 2239 2468
rect 2243 2464 2244 2468
rect 2238 2463 2244 2464
rect 2366 2468 2372 2469
rect 2366 2464 2367 2468
rect 2371 2464 2372 2468
rect 2366 2463 2372 2464
rect 1952 2439 1954 2463
rect 2040 2439 2042 2463
rect 2136 2439 2138 2463
rect 2240 2439 2242 2463
rect 2368 2439 2370 2463
rect 1767 2437 1771 2438
rect 1807 2438 1811 2439
rect 1168 2421 1170 2437
rect 1296 2421 1298 2437
rect 1424 2421 1426 2437
rect 1166 2420 1172 2421
rect 1166 2416 1167 2420
rect 1171 2416 1172 2420
rect 1166 2415 1172 2416
rect 1294 2420 1300 2421
rect 1294 2416 1295 2420
rect 1299 2416 1300 2420
rect 1294 2415 1300 2416
rect 1422 2420 1428 2421
rect 1422 2416 1423 2420
rect 1427 2416 1428 2420
rect 1768 2418 1770 2437
rect 1807 2433 1811 2434
rect 1951 2438 1955 2439
rect 1951 2433 1955 2434
rect 2039 2438 2043 2439
rect 2039 2433 2043 2434
rect 2135 2438 2139 2439
rect 2135 2433 2139 2434
rect 2215 2438 2219 2439
rect 2215 2433 2219 2434
rect 2239 2438 2243 2439
rect 2239 2433 2243 2434
rect 2303 2438 2307 2439
rect 2303 2433 2307 2434
rect 2367 2438 2371 2439
rect 2367 2433 2371 2434
rect 1422 2415 1428 2416
rect 1766 2417 1772 2418
rect 1766 2413 1767 2417
rect 1771 2413 1772 2417
rect 1808 2414 1810 2433
rect 2216 2417 2218 2433
rect 2262 2423 2268 2424
rect 2262 2419 2263 2423
rect 2267 2419 2268 2423
rect 2262 2418 2268 2419
rect 2214 2416 2220 2417
rect 1766 2412 1772 2413
rect 1806 2413 1812 2414
rect 1238 2411 1244 2412
rect 1238 2407 1239 2411
rect 1243 2407 1244 2411
rect 1238 2406 1244 2407
rect 1366 2411 1372 2412
rect 1366 2407 1367 2411
rect 1371 2407 1372 2411
rect 1366 2406 1372 2407
rect 1386 2411 1392 2412
rect 1386 2407 1387 2411
rect 1391 2407 1392 2411
rect 1806 2409 1807 2413
rect 1811 2409 1812 2413
rect 2214 2412 2215 2416
rect 2219 2412 2220 2416
rect 2214 2411 2220 2412
rect 1806 2408 1812 2409
rect 1386 2406 1392 2407
rect 1166 2401 1172 2402
rect 1166 2397 1167 2401
rect 1171 2397 1172 2401
rect 1166 2396 1172 2397
rect 1062 2383 1068 2384
rect 1062 2379 1063 2383
rect 1067 2379 1068 2383
rect 1062 2378 1068 2379
rect 1150 2383 1156 2384
rect 1150 2379 1151 2383
rect 1155 2379 1156 2383
rect 1150 2378 1156 2379
rect 582 2371 583 2375
rect 587 2371 588 2375
rect 582 2370 588 2371
rect 599 2374 603 2375
rect 599 2369 603 2370
rect 655 2374 659 2375
rect 655 2369 659 2370
rect 703 2374 707 2375
rect 703 2369 707 2370
rect 767 2374 771 2375
rect 767 2369 771 2370
rect 807 2374 811 2375
rect 807 2369 811 2370
rect 879 2374 883 2375
rect 879 2369 883 2370
rect 919 2374 923 2375
rect 919 2369 923 2370
rect 991 2374 995 2375
rect 998 2371 999 2375
rect 1003 2371 1004 2375
rect 998 2370 1004 2371
rect 1039 2374 1043 2375
rect 991 2369 995 2370
rect 1039 2369 1043 2370
rect 550 2367 556 2368
rect 550 2363 551 2367
rect 555 2363 556 2367
rect 550 2362 556 2363
rect 574 2367 580 2368
rect 574 2363 575 2367
rect 579 2363 580 2367
rect 574 2362 580 2363
rect 614 2367 620 2368
rect 614 2363 615 2367
rect 619 2363 620 2367
rect 614 2362 620 2363
rect 430 2351 436 2352
rect 430 2347 431 2351
rect 435 2347 436 2351
rect 430 2346 436 2347
rect 542 2351 548 2352
rect 542 2347 543 2351
rect 547 2347 548 2351
rect 542 2346 548 2347
rect 398 2343 404 2344
rect 398 2339 399 2343
rect 403 2339 404 2343
rect 398 2338 404 2339
rect 110 2335 116 2336
rect 110 2331 111 2335
rect 115 2331 116 2335
rect 398 2335 404 2336
rect 110 2330 116 2331
rect 318 2332 324 2333
rect 112 2303 114 2330
rect 318 2328 319 2332
rect 323 2328 324 2332
rect 398 2331 399 2335
rect 403 2331 404 2335
rect 398 2330 404 2331
rect 430 2332 436 2333
rect 318 2327 324 2328
rect 320 2303 322 2327
rect 111 2302 115 2303
rect 111 2297 115 2298
rect 151 2302 155 2303
rect 151 2297 155 2298
rect 271 2302 275 2303
rect 271 2297 275 2298
rect 319 2302 323 2303
rect 319 2297 323 2298
rect 391 2302 395 2303
rect 391 2297 395 2298
rect 112 2278 114 2297
rect 152 2281 154 2297
rect 202 2287 208 2288
rect 202 2283 203 2287
rect 207 2283 208 2287
rect 202 2282 208 2283
rect 150 2280 156 2281
rect 110 2277 116 2278
rect 110 2273 111 2277
rect 115 2273 116 2277
rect 150 2276 151 2280
rect 155 2276 156 2280
rect 150 2275 156 2276
rect 110 2272 116 2273
rect 150 2261 156 2262
rect 110 2260 116 2261
rect 110 2256 111 2260
rect 115 2256 116 2260
rect 150 2257 151 2261
rect 155 2257 156 2261
rect 150 2256 156 2257
rect 110 2255 116 2256
rect 112 2235 114 2255
rect 152 2235 154 2256
rect 204 2244 206 2282
rect 272 2281 274 2297
rect 392 2281 394 2297
rect 270 2280 276 2281
rect 270 2276 271 2280
rect 275 2276 276 2280
rect 270 2275 276 2276
rect 390 2280 396 2281
rect 390 2276 391 2280
rect 395 2276 396 2280
rect 390 2275 396 2276
rect 222 2271 228 2272
rect 222 2267 223 2271
rect 227 2267 228 2271
rect 222 2266 228 2267
rect 342 2271 348 2272
rect 342 2267 343 2271
rect 347 2267 348 2271
rect 342 2266 348 2267
rect 224 2244 226 2266
rect 270 2261 276 2262
rect 270 2257 271 2261
rect 275 2257 276 2261
rect 270 2256 276 2257
rect 202 2243 208 2244
rect 202 2239 203 2243
rect 207 2239 208 2243
rect 202 2238 208 2239
rect 222 2243 228 2244
rect 222 2239 223 2243
rect 227 2239 228 2243
rect 222 2238 228 2239
rect 272 2235 274 2256
rect 111 2234 115 2235
rect 111 2229 115 2230
rect 135 2234 139 2235
rect 135 2229 139 2230
rect 151 2234 155 2235
rect 151 2229 155 2230
rect 247 2234 251 2235
rect 247 2229 251 2230
rect 271 2234 275 2235
rect 271 2229 275 2230
rect 112 2213 114 2229
rect 110 2212 116 2213
rect 136 2212 138 2229
rect 214 2227 220 2228
rect 214 2223 215 2227
rect 219 2223 220 2227
rect 214 2222 220 2223
rect 110 2208 111 2212
rect 115 2208 116 2212
rect 110 2207 116 2208
rect 134 2211 140 2212
rect 134 2207 135 2211
rect 139 2207 140 2211
rect 134 2206 140 2207
rect 216 2204 218 2222
rect 248 2212 250 2229
rect 344 2228 346 2266
rect 390 2261 396 2262
rect 390 2257 391 2261
rect 395 2257 396 2261
rect 390 2256 396 2257
rect 392 2235 394 2256
rect 400 2244 402 2330
rect 430 2328 431 2332
rect 435 2328 436 2332
rect 430 2327 436 2328
rect 542 2332 548 2333
rect 542 2328 543 2332
rect 547 2328 548 2332
rect 552 2328 554 2362
rect 616 2344 618 2362
rect 656 2352 658 2369
rect 768 2352 770 2369
rect 846 2367 852 2368
rect 846 2363 847 2367
rect 851 2363 852 2367
rect 846 2362 852 2363
rect 866 2367 872 2368
rect 866 2363 867 2367
rect 871 2363 872 2367
rect 866 2362 872 2363
rect 654 2351 660 2352
rect 654 2347 655 2351
rect 659 2347 660 2351
rect 654 2346 660 2347
rect 766 2351 772 2352
rect 766 2347 767 2351
rect 771 2347 772 2351
rect 766 2346 772 2347
rect 614 2343 620 2344
rect 614 2339 615 2343
rect 619 2339 620 2343
rect 614 2338 620 2339
rect 654 2332 660 2333
rect 654 2328 655 2332
rect 659 2328 660 2332
rect 542 2327 548 2328
rect 550 2327 556 2328
rect 654 2327 660 2328
rect 766 2332 772 2333
rect 766 2328 767 2332
rect 771 2328 772 2332
rect 766 2327 772 2328
rect 432 2303 434 2327
rect 544 2303 546 2327
rect 550 2323 551 2327
rect 555 2323 556 2327
rect 550 2322 556 2323
rect 656 2303 658 2327
rect 768 2303 770 2327
rect 431 2302 435 2303
rect 431 2297 435 2298
rect 519 2302 523 2303
rect 519 2297 523 2298
rect 543 2302 547 2303
rect 543 2297 547 2298
rect 647 2302 651 2303
rect 647 2297 651 2298
rect 655 2302 659 2303
rect 655 2297 659 2298
rect 767 2302 771 2303
rect 767 2297 771 2298
rect 775 2302 779 2303
rect 775 2297 779 2298
rect 520 2281 522 2297
rect 648 2281 650 2297
rect 776 2281 778 2297
rect 518 2280 524 2281
rect 518 2276 519 2280
rect 523 2276 524 2280
rect 518 2275 524 2276
rect 646 2280 652 2281
rect 646 2276 647 2280
rect 651 2276 652 2280
rect 646 2275 652 2276
rect 774 2280 780 2281
rect 774 2276 775 2280
rect 779 2276 780 2280
rect 774 2275 780 2276
rect 848 2272 850 2362
rect 868 2344 870 2362
rect 880 2352 882 2369
rect 950 2367 956 2368
rect 950 2363 951 2367
rect 955 2363 956 2367
rect 950 2362 956 2363
rect 878 2351 884 2352
rect 878 2347 879 2351
rect 883 2347 884 2351
rect 878 2346 884 2347
rect 952 2344 954 2362
rect 992 2352 994 2369
rect 990 2351 996 2352
rect 990 2347 991 2351
rect 995 2347 996 2351
rect 990 2346 996 2347
rect 1064 2344 1066 2378
rect 1168 2375 1170 2396
rect 1240 2384 1242 2406
rect 1294 2401 1300 2402
rect 1294 2397 1295 2401
rect 1299 2397 1300 2401
rect 1294 2396 1300 2397
rect 1238 2383 1244 2384
rect 1238 2379 1239 2383
rect 1243 2379 1244 2383
rect 1238 2378 1244 2379
rect 1296 2375 1298 2396
rect 1368 2384 1370 2406
rect 1366 2383 1372 2384
rect 1366 2379 1367 2383
rect 1371 2379 1372 2383
rect 1366 2378 1372 2379
rect 1103 2374 1107 2375
rect 1103 2369 1107 2370
rect 1167 2374 1171 2375
rect 1167 2369 1171 2370
rect 1215 2374 1219 2375
rect 1215 2369 1219 2370
rect 1295 2374 1299 2375
rect 1295 2369 1299 2370
rect 1335 2374 1339 2375
rect 1335 2369 1339 2370
rect 1104 2352 1106 2369
rect 1206 2367 1212 2368
rect 1206 2363 1207 2367
rect 1211 2363 1212 2367
rect 1206 2362 1212 2363
rect 1102 2351 1108 2352
rect 1102 2347 1103 2351
rect 1107 2347 1108 2351
rect 1102 2346 1108 2347
rect 1208 2344 1210 2362
rect 1216 2352 1218 2369
rect 1336 2352 1338 2369
rect 1388 2368 1390 2406
rect 1422 2401 1428 2402
rect 1422 2397 1423 2401
rect 1427 2397 1428 2401
rect 1422 2396 1428 2397
rect 1766 2400 1772 2401
rect 1766 2396 1767 2400
rect 1771 2396 1772 2400
rect 2214 2397 2220 2398
rect 1424 2375 1426 2396
rect 1766 2395 1772 2396
rect 1806 2396 1812 2397
rect 1768 2375 1770 2395
rect 1806 2392 1807 2396
rect 1811 2392 1812 2396
rect 2214 2393 2215 2397
rect 2219 2393 2220 2397
rect 2214 2392 2220 2393
rect 1806 2391 1812 2392
rect 1808 2375 1810 2391
rect 2216 2375 2218 2392
rect 2264 2384 2266 2418
rect 2304 2417 2306 2433
rect 2302 2416 2308 2417
rect 2302 2412 2303 2416
rect 2307 2412 2308 2416
rect 2302 2411 2308 2412
rect 2376 2408 2378 2498
rect 2528 2488 2530 2505
rect 2580 2504 2582 2554
rect 2648 2553 2650 2569
rect 2816 2553 2818 2569
rect 3000 2553 3002 2569
rect 3192 2553 3194 2569
rect 2646 2552 2652 2553
rect 2646 2548 2647 2552
rect 2651 2548 2652 2552
rect 2646 2547 2652 2548
rect 2814 2552 2820 2553
rect 2814 2548 2815 2552
rect 2819 2548 2820 2552
rect 2814 2547 2820 2548
rect 2998 2552 3004 2553
rect 2998 2548 2999 2552
rect 3003 2548 3004 2552
rect 2998 2547 3004 2548
rect 3190 2552 3196 2553
rect 3190 2548 3191 2552
rect 3195 2548 3196 2552
rect 3190 2547 3196 2548
rect 3264 2544 3266 2794
rect 3304 2776 3306 2810
rect 3368 2807 3370 2828
rect 3367 2806 3371 2807
rect 3367 2801 3371 2802
rect 3368 2784 3370 2801
rect 3432 2800 3434 2838
rect 3440 2816 3442 2978
rect 3462 2972 3468 2973
rect 3462 2968 3463 2972
rect 3467 2968 3468 2972
rect 3462 2967 3468 2968
rect 3464 2939 3466 2967
rect 3463 2938 3467 2939
rect 3463 2933 3467 2934
rect 3464 2917 3466 2933
rect 3462 2916 3468 2917
rect 3462 2912 3463 2916
rect 3467 2912 3468 2916
rect 3462 2911 3468 2912
rect 3462 2899 3468 2900
rect 3462 2895 3463 2899
rect 3467 2895 3468 2899
rect 3462 2894 3468 2895
rect 3464 2875 3466 2894
rect 3463 2874 3467 2875
rect 3463 2869 3467 2870
rect 3464 2850 3466 2869
rect 3462 2849 3468 2850
rect 3462 2845 3463 2849
rect 3467 2845 3468 2849
rect 3462 2844 3468 2845
rect 3462 2832 3468 2833
rect 3462 2828 3463 2832
rect 3467 2828 3468 2832
rect 3462 2827 3468 2828
rect 3438 2815 3444 2816
rect 3438 2811 3439 2815
rect 3443 2811 3444 2815
rect 3438 2810 3444 2811
rect 3464 2807 3466 2827
rect 3463 2806 3467 2807
rect 3463 2801 3467 2802
rect 3430 2799 3436 2800
rect 3430 2795 3431 2799
rect 3435 2795 3436 2799
rect 3430 2794 3436 2795
rect 3464 2785 3466 2801
rect 3462 2784 3468 2785
rect 3366 2783 3372 2784
rect 3366 2779 3367 2783
rect 3371 2779 3372 2783
rect 3462 2780 3463 2784
rect 3467 2780 3468 2784
rect 3462 2779 3468 2780
rect 3366 2778 3372 2779
rect 3302 2775 3308 2776
rect 3302 2771 3303 2775
rect 3307 2771 3308 2775
rect 3302 2770 3308 2771
rect 3438 2771 3444 2772
rect 3438 2767 3439 2771
rect 3443 2767 3444 2771
rect 3438 2766 3444 2767
rect 3462 2767 3468 2768
rect 3366 2764 3372 2765
rect 3366 2760 3367 2764
rect 3371 2760 3372 2764
rect 3366 2759 3372 2760
rect 3368 2727 3370 2759
rect 3367 2726 3371 2727
rect 3367 2721 3371 2722
rect 3368 2705 3370 2721
rect 3366 2704 3372 2705
rect 3366 2700 3367 2704
rect 3371 2700 3372 2704
rect 3366 2699 3372 2700
rect 3430 2695 3436 2696
rect 3430 2691 3431 2695
rect 3435 2691 3436 2695
rect 3430 2690 3436 2691
rect 3366 2685 3372 2686
rect 3366 2681 3367 2685
rect 3371 2681 3372 2685
rect 3366 2680 3372 2681
rect 3368 2651 3370 2680
rect 3367 2650 3371 2651
rect 3367 2645 3371 2646
rect 3368 2628 3370 2645
rect 3432 2644 3434 2690
rect 3440 2668 3442 2766
rect 3462 2763 3463 2767
rect 3467 2763 3468 2767
rect 3462 2762 3468 2763
rect 3464 2727 3466 2762
rect 3463 2726 3467 2727
rect 3463 2721 3467 2722
rect 3464 2702 3466 2721
rect 3462 2701 3468 2702
rect 3462 2697 3463 2701
rect 3467 2697 3468 2701
rect 3462 2696 3468 2697
rect 3462 2684 3468 2685
rect 3462 2680 3463 2684
rect 3467 2680 3468 2684
rect 3462 2679 3468 2680
rect 3438 2667 3444 2668
rect 3438 2663 3439 2667
rect 3443 2663 3444 2667
rect 3438 2662 3444 2663
rect 3464 2651 3466 2679
rect 3463 2650 3467 2651
rect 3463 2645 3467 2646
rect 3430 2643 3436 2644
rect 3430 2639 3431 2643
rect 3435 2639 3436 2643
rect 3430 2638 3436 2639
rect 3464 2629 3466 2645
rect 3462 2628 3468 2629
rect 3366 2627 3372 2628
rect 3366 2623 3367 2627
rect 3371 2623 3372 2627
rect 3462 2624 3463 2628
rect 3467 2624 3468 2628
rect 3462 2623 3468 2624
rect 3366 2622 3372 2623
rect 3438 2615 3444 2616
rect 3438 2611 3439 2615
rect 3443 2611 3444 2615
rect 3438 2610 3444 2611
rect 3462 2611 3468 2612
rect 3366 2608 3372 2609
rect 3366 2604 3367 2608
rect 3371 2604 3372 2608
rect 3366 2603 3372 2604
rect 3368 2575 3370 2603
rect 3367 2574 3371 2575
rect 3367 2569 3371 2570
rect 3368 2553 3370 2569
rect 3366 2552 3372 2553
rect 3366 2548 3367 2552
rect 3371 2548 3372 2552
rect 3366 2547 3372 2548
rect 2718 2543 2724 2544
rect 2718 2539 2719 2543
rect 2723 2539 2724 2543
rect 2718 2538 2724 2539
rect 2886 2543 2892 2544
rect 2886 2539 2887 2543
rect 2891 2539 2892 2543
rect 2886 2538 2892 2539
rect 3262 2543 3268 2544
rect 3262 2539 3263 2543
rect 3267 2539 3268 2543
rect 3262 2538 3268 2539
rect 3430 2543 3436 2544
rect 3430 2539 3431 2543
rect 3435 2539 3436 2543
rect 3430 2538 3436 2539
rect 2646 2533 2652 2534
rect 2646 2529 2647 2533
rect 2651 2529 2652 2533
rect 2646 2528 2652 2529
rect 2648 2511 2650 2528
rect 2720 2516 2722 2538
rect 2814 2533 2820 2534
rect 2814 2529 2815 2533
rect 2819 2529 2820 2533
rect 2814 2528 2820 2529
rect 2718 2515 2724 2516
rect 2718 2511 2719 2515
rect 2723 2511 2724 2515
rect 2816 2511 2818 2528
rect 2888 2516 2890 2538
rect 2998 2533 3004 2534
rect 2998 2529 2999 2533
rect 3003 2529 3004 2533
rect 2998 2528 3004 2529
rect 3190 2533 3196 2534
rect 3190 2529 3191 2533
rect 3195 2529 3196 2533
rect 3190 2528 3196 2529
rect 3366 2533 3372 2534
rect 3366 2529 3367 2533
rect 3371 2529 3372 2533
rect 3366 2528 3372 2529
rect 2886 2515 2892 2516
rect 2886 2511 2887 2515
rect 2891 2511 2892 2515
rect 3000 2511 3002 2528
rect 3192 2511 3194 2528
rect 3242 2515 3248 2516
rect 3242 2511 3243 2515
rect 3247 2511 3248 2515
rect 3368 2511 3370 2528
rect 2647 2510 2651 2511
rect 2647 2505 2651 2506
rect 2711 2510 2715 2511
rect 2718 2510 2724 2511
rect 2815 2510 2819 2511
rect 2886 2510 2892 2511
rect 2919 2510 2923 2511
rect 2711 2505 2715 2506
rect 2815 2505 2819 2506
rect 2919 2505 2923 2506
rect 2999 2510 3003 2511
rect 2999 2505 3003 2506
rect 3143 2510 3147 2511
rect 3143 2505 3147 2506
rect 3191 2510 3195 2511
rect 3242 2510 3248 2511
rect 3367 2510 3371 2511
rect 3191 2505 3195 2506
rect 2578 2503 2584 2504
rect 2578 2499 2579 2503
rect 2583 2499 2584 2503
rect 2578 2498 2584 2499
rect 2598 2503 2604 2504
rect 2598 2499 2599 2503
rect 2603 2499 2604 2503
rect 2598 2498 2604 2499
rect 2526 2487 2532 2488
rect 2526 2483 2527 2487
rect 2531 2483 2532 2487
rect 2526 2482 2532 2483
rect 2600 2480 2602 2498
rect 2712 2488 2714 2505
rect 2782 2503 2788 2504
rect 2782 2499 2783 2503
rect 2787 2499 2788 2503
rect 2782 2498 2788 2499
rect 2710 2487 2716 2488
rect 2710 2483 2711 2487
rect 2715 2483 2716 2487
rect 2710 2482 2716 2483
rect 2784 2480 2786 2498
rect 2920 2488 2922 2505
rect 2990 2503 2996 2504
rect 2990 2499 2991 2503
rect 2995 2499 2996 2503
rect 2990 2498 2996 2499
rect 2918 2487 2924 2488
rect 2918 2483 2919 2487
rect 2923 2483 2924 2487
rect 2918 2482 2924 2483
rect 2992 2480 2994 2498
rect 3144 2488 3146 2505
rect 3142 2487 3148 2488
rect 3142 2483 3143 2487
rect 3147 2483 3148 2487
rect 3142 2482 3148 2483
rect 3244 2480 3246 2510
rect 3367 2505 3371 2506
rect 3368 2488 3370 2505
rect 3432 2504 3434 2538
rect 3440 2516 3442 2610
rect 3462 2607 3463 2611
rect 3467 2607 3468 2611
rect 3462 2606 3468 2607
rect 3464 2575 3466 2606
rect 3463 2574 3467 2575
rect 3463 2569 3467 2570
rect 3464 2550 3466 2569
rect 3462 2549 3468 2550
rect 3462 2545 3463 2549
rect 3467 2545 3468 2549
rect 3462 2544 3468 2545
rect 3462 2532 3468 2533
rect 3462 2528 3463 2532
rect 3467 2528 3468 2532
rect 3462 2527 3468 2528
rect 3438 2515 3444 2516
rect 3438 2511 3439 2515
rect 3443 2511 3444 2515
rect 3464 2511 3466 2527
rect 3438 2510 3444 2511
rect 3463 2510 3467 2511
rect 3463 2505 3467 2506
rect 3430 2503 3436 2504
rect 3430 2499 3431 2503
rect 3435 2499 3436 2503
rect 3430 2498 3436 2499
rect 3464 2489 3466 2505
rect 3462 2488 3468 2489
rect 3366 2487 3372 2488
rect 3366 2483 3367 2487
rect 3371 2483 3372 2487
rect 3462 2484 3463 2488
rect 3467 2484 3468 2488
rect 3462 2483 3468 2484
rect 3366 2482 3372 2483
rect 2598 2479 2604 2480
rect 2598 2475 2599 2479
rect 2603 2475 2604 2479
rect 2598 2474 2604 2475
rect 2782 2479 2788 2480
rect 2782 2475 2783 2479
rect 2787 2475 2788 2479
rect 2782 2474 2788 2475
rect 2990 2479 2996 2480
rect 2990 2475 2991 2479
rect 2995 2475 2996 2479
rect 2990 2474 2996 2475
rect 3078 2479 3084 2480
rect 3078 2475 3079 2479
rect 3083 2475 3084 2479
rect 3078 2474 3084 2475
rect 3242 2479 3248 2480
rect 3242 2475 3243 2479
rect 3247 2475 3248 2479
rect 3242 2474 3248 2475
rect 2526 2468 2532 2469
rect 2526 2464 2527 2468
rect 2531 2464 2532 2468
rect 2526 2463 2532 2464
rect 2710 2468 2716 2469
rect 2710 2464 2711 2468
rect 2715 2464 2716 2468
rect 2710 2463 2716 2464
rect 2918 2468 2924 2469
rect 2918 2464 2919 2468
rect 2923 2464 2924 2468
rect 2918 2463 2924 2464
rect 2528 2439 2530 2463
rect 2712 2439 2714 2463
rect 2920 2439 2922 2463
rect 2391 2438 2395 2439
rect 2391 2433 2395 2434
rect 2479 2438 2483 2439
rect 2479 2433 2483 2434
rect 2527 2438 2531 2439
rect 2527 2433 2531 2434
rect 2567 2438 2571 2439
rect 2567 2433 2571 2434
rect 2655 2438 2659 2439
rect 2655 2433 2659 2434
rect 2711 2438 2715 2439
rect 2711 2433 2715 2434
rect 2743 2438 2747 2439
rect 2743 2433 2747 2434
rect 2839 2438 2843 2439
rect 2839 2433 2843 2434
rect 2919 2438 2923 2439
rect 2919 2433 2923 2434
rect 2935 2438 2939 2439
rect 2935 2433 2939 2434
rect 2392 2417 2394 2433
rect 2480 2417 2482 2433
rect 2568 2417 2570 2433
rect 2618 2431 2624 2432
rect 2618 2427 2619 2431
rect 2623 2427 2624 2431
rect 2618 2426 2624 2427
rect 2390 2416 2396 2417
rect 2390 2412 2391 2416
rect 2395 2412 2396 2416
rect 2390 2411 2396 2412
rect 2478 2416 2484 2417
rect 2478 2412 2479 2416
rect 2483 2412 2484 2416
rect 2478 2411 2484 2412
rect 2566 2416 2572 2417
rect 2566 2412 2567 2416
rect 2571 2412 2572 2416
rect 2566 2411 2572 2412
rect 2286 2407 2292 2408
rect 2286 2403 2287 2407
rect 2291 2403 2292 2407
rect 2286 2402 2292 2403
rect 2374 2407 2380 2408
rect 2374 2403 2375 2407
rect 2379 2403 2380 2407
rect 2374 2402 2380 2403
rect 2262 2383 2268 2384
rect 2262 2379 2263 2383
rect 2267 2379 2268 2383
rect 2288 2380 2290 2402
rect 2302 2397 2308 2398
rect 2302 2393 2303 2397
rect 2307 2393 2308 2397
rect 2302 2392 2308 2393
rect 2390 2397 2396 2398
rect 2390 2393 2391 2397
rect 2395 2393 2396 2397
rect 2390 2392 2396 2393
rect 2478 2397 2484 2398
rect 2478 2393 2479 2397
rect 2483 2393 2484 2397
rect 2478 2392 2484 2393
rect 2566 2397 2572 2398
rect 2566 2393 2567 2397
rect 2571 2393 2572 2397
rect 2566 2392 2572 2393
rect 2262 2378 2268 2379
rect 2286 2379 2292 2380
rect 2286 2375 2287 2379
rect 2291 2375 2292 2379
rect 2304 2375 2306 2392
rect 2392 2375 2394 2392
rect 2480 2375 2482 2392
rect 2550 2379 2556 2380
rect 2550 2375 2551 2379
rect 2555 2375 2556 2379
rect 2568 2375 2570 2392
rect 2620 2380 2622 2426
rect 2656 2417 2658 2433
rect 2744 2417 2746 2433
rect 2750 2423 2756 2424
rect 2750 2419 2751 2423
rect 2755 2419 2756 2423
rect 2750 2418 2756 2419
rect 2654 2416 2660 2417
rect 2654 2412 2655 2416
rect 2659 2412 2660 2416
rect 2654 2411 2660 2412
rect 2742 2416 2748 2417
rect 2742 2412 2743 2416
rect 2747 2412 2748 2416
rect 2742 2411 2748 2412
rect 2638 2407 2644 2408
rect 2638 2403 2639 2407
rect 2643 2403 2644 2407
rect 2638 2402 2644 2403
rect 2726 2407 2732 2408
rect 2726 2403 2727 2407
rect 2731 2403 2732 2407
rect 2726 2402 2732 2403
rect 2640 2380 2642 2402
rect 2654 2397 2660 2398
rect 2654 2393 2655 2397
rect 2659 2393 2660 2397
rect 2654 2392 2660 2393
rect 2618 2379 2624 2380
rect 2618 2375 2619 2379
rect 2623 2375 2624 2379
rect 1423 2374 1427 2375
rect 1423 2369 1427 2370
rect 1767 2374 1771 2375
rect 1767 2369 1771 2370
rect 1807 2374 1811 2375
rect 1807 2369 1811 2370
rect 2167 2374 2171 2375
rect 2167 2369 2171 2370
rect 2215 2374 2219 2375
rect 2215 2369 2219 2370
rect 2263 2374 2267 2375
rect 2286 2374 2292 2375
rect 2303 2374 2307 2375
rect 2263 2369 2267 2370
rect 2303 2369 2307 2370
rect 2367 2374 2371 2375
rect 2367 2369 2371 2370
rect 2391 2374 2395 2375
rect 2391 2369 2395 2370
rect 2471 2374 2475 2375
rect 2471 2369 2475 2370
rect 2479 2374 2483 2375
rect 2550 2374 2556 2375
rect 2567 2374 2571 2375
rect 2479 2369 2483 2370
rect 1386 2367 1392 2368
rect 1386 2363 1387 2367
rect 1391 2363 1392 2367
rect 1386 2362 1392 2363
rect 1768 2353 1770 2369
rect 1808 2353 1810 2369
rect 1766 2352 1772 2353
rect 1214 2351 1220 2352
rect 1214 2347 1215 2351
rect 1219 2347 1220 2351
rect 1214 2346 1220 2347
rect 1334 2351 1340 2352
rect 1334 2347 1335 2351
rect 1339 2347 1340 2351
rect 1766 2348 1767 2352
rect 1771 2348 1772 2352
rect 1766 2347 1772 2348
rect 1806 2352 1812 2353
rect 2168 2352 2170 2369
rect 2230 2367 2236 2368
rect 2230 2363 2231 2367
rect 2235 2363 2236 2367
rect 2230 2362 2236 2363
rect 2238 2367 2244 2368
rect 2238 2363 2239 2367
rect 2243 2363 2244 2367
rect 2238 2362 2244 2363
rect 1806 2348 1807 2352
rect 1811 2348 1812 2352
rect 1806 2347 1812 2348
rect 2166 2351 2172 2352
rect 2166 2347 2167 2351
rect 2171 2347 2172 2351
rect 1334 2346 1340 2347
rect 2166 2346 2172 2347
rect 866 2343 872 2344
rect 866 2339 867 2343
rect 871 2339 872 2343
rect 866 2338 872 2339
rect 950 2343 956 2344
rect 950 2339 951 2343
rect 955 2339 956 2343
rect 950 2338 956 2339
rect 1062 2343 1068 2344
rect 1062 2339 1063 2343
rect 1067 2339 1068 2343
rect 1062 2338 1068 2339
rect 1070 2343 1076 2344
rect 1070 2339 1071 2343
rect 1075 2339 1076 2343
rect 1070 2338 1076 2339
rect 1206 2343 1212 2344
rect 1206 2339 1207 2343
rect 1211 2339 1212 2343
rect 1206 2338 1212 2339
rect 878 2332 884 2333
rect 878 2328 879 2332
rect 883 2328 884 2332
rect 878 2327 884 2328
rect 990 2332 996 2333
rect 990 2328 991 2332
rect 995 2328 996 2332
rect 990 2327 996 2328
rect 880 2303 882 2327
rect 992 2303 994 2327
rect 879 2302 883 2303
rect 879 2297 883 2298
rect 895 2302 899 2303
rect 895 2297 899 2298
rect 991 2302 995 2303
rect 991 2297 995 2298
rect 1015 2302 1019 2303
rect 1015 2297 1019 2298
rect 896 2281 898 2297
rect 1016 2281 1018 2297
rect 894 2280 900 2281
rect 894 2276 895 2280
rect 899 2276 900 2280
rect 894 2275 900 2276
rect 1014 2280 1020 2281
rect 1014 2276 1015 2280
rect 1019 2276 1020 2280
rect 1014 2275 1020 2276
rect 462 2271 468 2272
rect 462 2267 463 2271
rect 467 2267 468 2271
rect 462 2266 468 2267
rect 590 2271 596 2272
rect 590 2267 591 2271
rect 595 2267 596 2271
rect 590 2266 596 2267
rect 846 2271 852 2272
rect 846 2267 847 2271
rect 851 2267 852 2271
rect 846 2266 852 2267
rect 854 2271 860 2272
rect 854 2267 855 2271
rect 859 2267 860 2271
rect 854 2266 860 2267
rect 464 2244 466 2266
rect 518 2261 524 2262
rect 518 2257 519 2261
rect 523 2257 524 2261
rect 518 2256 524 2257
rect 398 2243 404 2244
rect 398 2239 399 2243
rect 403 2239 404 2243
rect 398 2238 404 2239
rect 462 2243 468 2244
rect 462 2239 463 2243
rect 467 2239 468 2243
rect 462 2238 468 2239
rect 520 2235 522 2256
rect 592 2244 594 2266
rect 646 2261 652 2262
rect 646 2257 647 2261
rect 651 2257 652 2261
rect 646 2256 652 2257
rect 774 2261 780 2262
rect 774 2257 775 2261
rect 779 2257 780 2261
rect 774 2256 780 2257
rect 590 2243 596 2244
rect 590 2239 591 2243
rect 595 2239 596 2243
rect 590 2238 596 2239
rect 648 2235 650 2256
rect 738 2235 744 2236
rect 776 2235 778 2256
rect 856 2244 858 2266
rect 894 2261 900 2262
rect 894 2257 895 2261
rect 899 2257 900 2261
rect 894 2256 900 2257
rect 1014 2261 1020 2262
rect 1014 2257 1015 2261
rect 1019 2257 1020 2261
rect 1014 2256 1020 2257
rect 854 2243 860 2244
rect 854 2239 855 2243
rect 859 2239 860 2243
rect 854 2238 860 2239
rect 896 2235 898 2256
rect 942 2243 948 2244
rect 942 2239 943 2243
rect 947 2239 948 2243
rect 942 2238 948 2239
rect 391 2234 395 2235
rect 391 2229 395 2230
rect 407 2234 411 2235
rect 407 2229 411 2230
rect 519 2234 523 2235
rect 519 2229 523 2230
rect 583 2234 587 2235
rect 583 2229 587 2230
rect 647 2234 651 2235
rect 738 2231 739 2235
rect 743 2231 744 2235
rect 738 2230 744 2231
rect 767 2234 771 2235
rect 647 2229 651 2230
rect 342 2227 348 2228
rect 342 2223 343 2227
rect 347 2223 348 2227
rect 342 2222 348 2223
rect 408 2212 410 2229
rect 478 2227 484 2228
rect 478 2223 479 2227
rect 483 2223 484 2227
rect 478 2222 484 2223
rect 246 2211 252 2212
rect 246 2207 247 2211
rect 251 2207 252 2211
rect 246 2206 252 2207
rect 406 2211 412 2212
rect 406 2207 407 2211
rect 411 2207 412 2211
rect 406 2206 412 2207
rect 480 2204 482 2222
rect 584 2212 586 2229
rect 654 2227 660 2228
rect 654 2223 655 2227
rect 659 2223 660 2227
rect 654 2222 660 2223
rect 582 2211 588 2212
rect 582 2207 583 2211
rect 587 2207 588 2211
rect 582 2206 588 2207
rect 656 2204 658 2222
rect 740 2204 742 2230
rect 767 2229 771 2230
rect 775 2234 779 2235
rect 775 2229 779 2230
rect 895 2234 899 2235
rect 895 2229 899 2230
rect 768 2212 770 2229
rect 766 2211 772 2212
rect 766 2207 767 2211
rect 771 2207 772 2211
rect 766 2206 772 2207
rect 944 2204 946 2238
rect 1016 2235 1018 2256
rect 1063 2243 1069 2244
rect 1063 2239 1064 2243
rect 1068 2242 1069 2243
rect 1072 2242 1074 2338
rect 1766 2335 1772 2336
rect 1102 2332 1108 2333
rect 1102 2328 1103 2332
rect 1107 2328 1108 2332
rect 1102 2327 1108 2328
rect 1214 2332 1220 2333
rect 1214 2328 1215 2332
rect 1219 2328 1220 2332
rect 1214 2327 1220 2328
rect 1334 2332 1340 2333
rect 1334 2328 1335 2332
rect 1339 2328 1340 2332
rect 1766 2331 1767 2335
rect 1771 2331 1772 2335
rect 1766 2330 1772 2331
rect 1806 2335 1812 2336
rect 1806 2331 1807 2335
rect 1811 2331 1812 2335
rect 1806 2330 1812 2331
rect 2166 2332 2172 2333
rect 1334 2327 1340 2328
rect 1104 2303 1106 2327
rect 1216 2303 1218 2327
rect 1336 2303 1338 2327
rect 1768 2303 1770 2330
rect 1808 2303 1810 2330
rect 2166 2328 2167 2332
rect 2171 2328 2172 2332
rect 2166 2327 2172 2328
rect 2168 2303 2170 2327
rect 1103 2302 1107 2303
rect 1103 2297 1107 2298
rect 1143 2302 1147 2303
rect 1143 2297 1147 2298
rect 1215 2302 1219 2303
rect 1215 2297 1219 2298
rect 1271 2302 1275 2303
rect 1271 2297 1275 2298
rect 1335 2302 1339 2303
rect 1335 2297 1339 2298
rect 1767 2302 1771 2303
rect 1767 2297 1771 2298
rect 1807 2302 1811 2303
rect 1807 2297 1811 2298
rect 1887 2302 1891 2303
rect 1887 2297 1891 2298
rect 2039 2302 2043 2303
rect 2039 2297 2043 2298
rect 2167 2302 2171 2303
rect 2167 2297 2171 2298
rect 2199 2302 2203 2303
rect 2199 2297 2203 2298
rect 1144 2281 1146 2297
rect 1272 2281 1274 2297
rect 1142 2280 1148 2281
rect 1142 2276 1143 2280
rect 1147 2276 1148 2280
rect 1142 2275 1148 2276
rect 1270 2280 1276 2281
rect 1270 2276 1271 2280
rect 1275 2276 1276 2280
rect 1768 2278 1770 2297
rect 1808 2278 1810 2297
rect 1888 2281 1890 2297
rect 2040 2281 2042 2297
rect 2200 2281 2202 2297
rect 2232 2288 2234 2362
rect 2240 2344 2242 2362
rect 2264 2352 2266 2369
rect 2334 2367 2340 2368
rect 2334 2363 2335 2367
rect 2339 2363 2340 2367
rect 2334 2362 2340 2363
rect 2262 2351 2268 2352
rect 2262 2347 2263 2351
rect 2267 2347 2268 2351
rect 2262 2346 2268 2347
rect 2336 2344 2338 2362
rect 2368 2352 2370 2369
rect 2438 2367 2444 2368
rect 2438 2363 2439 2367
rect 2443 2363 2444 2367
rect 2438 2362 2444 2363
rect 2366 2351 2372 2352
rect 2366 2347 2367 2351
rect 2371 2347 2372 2351
rect 2366 2346 2372 2347
rect 2440 2344 2442 2362
rect 2472 2352 2474 2369
rect 2542 2367 2548 2368
rect 2542 2363 2543 2367
rect 2547 2363 2548 2367
rect 2542 2362 2548 2363
rect 2470 2351 2476 2352
rect 2470 2347 2471 2351
rect 2475 2347 2476 2351
rect 2470 2346 2476 2347
rect 2544 2344 2546 2362
rect 2552 2344 2554 2374
rect 2567 2369 2571 2370
rect 2575 2374 2579 2375
rect 2618 2374 2624 2375
rect 2638 2379 2644 2380
rect 2638 2375 2639 2379
rect 2643 2375 2644 2379
rect 2656 2375 2658 2392
rect 2728 2380 2730 2402
rect 2742 2397 2748 2398
rect 2742 2393 2743 2397
rect 2747 2393 2748 2397
rect 2742 2392 2748 2393
rect 2726 2379 2732 2380
rect 2726 2375 2727 2379
rect 2731 2375 2732 2379
rect 2744 2375 2746 2392
rect 2638 2374 2644 2375
rect 2655 2374 2659 2375
rect 2575 2369 2579 2370
rect 2655 2369 2659 2370
rect 2687 2374 2691 2375
rect 2726 2374 2732 2375
rect 2743 2374 2747 2375
rect 2687 2369 2691 2370
rect 2743 2369 2747 2370
rect 2576 2352 2578 2369
rect 2688 2352 2690 2369
rect 2752 2368 2754 2418
rect 2840 2417 2842 2433
rect 2936 2417 2938 2433
rect 3080 2432 3082 2474
rect 3462 2471 3468 2472
rect 3142 2468 3148 2469
rect 3142 2464 3143 2468
rect 3147 2464 3148 2468
rect 3142 2463 3148 2464
rect 3366 2468 3372 2469
rect 3366 2464 3367 2468
rect 3371 2464 3372 2468
rect 3462 2467 3463 2471
rect 3467 2467 3468 2471
rect 3462 2466 3468 2467
rect 3366 2463 3372 2464
rect 3144 2439 3146 2463
rect 3368 2439 3370 2463
rect 3464 2439 3466 2466
rect 3143 2438 3147 2439
rect 3143 2433 3147 2434
rect 3367 2438 3371 2439
rect 3367 2433 3371 2434
rect 3463 2438 3467 2439
rect 3463 2433 3467 2434
rect 3078 2431 3084 2432
rect 3078 2427 3079 2431
rect 3083 2427 3084 2431
rect 3078 2426 3084 2427
rect 2838 2416 2844 2417
rect 2838 2412 2839 2416
rect 2843 2412 2844 2416
rect 2838 2411 2844 2412
rect 2934 2416 2940 2417
rect 2934 2412 2935 2416
rect 2939 2412 2940 2416
rect 3464 2414 3466 2433
rect 2934 2411 2940 2412
rect 3462 2413 3468 2414
rect 3462 2409 3463 2413
rect 3467 2409 3468 2413
rect 3462 2408 3468 2409
rect 2814 2407 2820 2408
rect 2814 2403 2815 2407
rect 2819 2403 2820 2407
rect 2814 2402 2820 2403
rect 2816 2380 2818 2402
rect 2926 2399 2932 2400
rect 2838 2397 2844 2398
rect 2838 2393 2839 2397
rect 2843 2393 2844 2397
rect 2926 2395 2927 2399
rect 2931 2395 2932 2399
rect 2926 2394 2932 2395
rect 2934 2397 2940 2398
rect 2838 2392 2844 2393
rect 2814 2379 2820 2380
rect 2814 2375 2815 2379
rect 2819 2375 2820 2379
rect 2840 2375 2842 2392
rect 2928 2380 2930 2394
rect 2934 2393 2935 2397
rect 2939 2393 2940 2397
rect 2934 2392 2940 2393
rect 3462 2396 3468 2397
rect 3462 2392 3463 2396
rect 3467 2392 3468 2396
rect 2926 2379 2932 2380
rect 2926 2375 2927 2379
rect 2931 2375 2932 2379
rect 2936 2375 2938 2392
rect 3462 2391 3468 2392
rect 3464 2375 3466 2391
rect 2799 2374 2803 2375
rect 2814 2374 2820 2375
rect 2839 2374 2843 2375
rect 2799 2369 2803 2370
rect 2839 2369 2843 2370
rect 2911 2374 2915 2375
rect 2926 2374 2932 2375
rect 2935 2374 2939 2375
rect 2911 2369 2915 2370
rect 2935 2369 2939 2370
rect 3023 2374 3027 2375
rect 3023 2369 3027 2370
rect 3463 2374 3467 2375
rect 3463 2369 3467 2370
rect 2750 2367 2756 2368
rect 2750 2363 2751 2367
rect 2755 2363 2756 2367
rect 2750 2362 2756 2363
rect 2758 2367 2764 2368
rect 2758 2363 2759 2367
rect 2763 2363 2764 2367
rect 2758 2362 2764 2363
rect 2574 2351 2580 2352
rect 2574 2347 2575 2351
rect 2579 2347 2580 2351
rect 2574 2346 2580 2347
rect 2686 2351 2692 2352
rect 2686 2347 2687 2351
rect 2691 2347 2692 2351
rect 2686 2346 2692 2347
rect 2760 2344 2762 2362
rect 2800 2352 2802 2369
rect 2870 2367 2876 2368
rect 2870 2363 2871 2367
rect 2875 2363 2876 2367
rect 2870 2362 2876 2363
rect 2798 2351 2804 2352
rect 2798 2347 2799 2351
rect 2803 2347 2804 2351
rect 2798 2346 2804 2347
rect 2872 2344 2874 2362
rect 2912 2352 2914 2369
rect 2982 2367 2988 2368
rect 2982 2363 2983 2367
rect 2987 2363 2988 2367
rect 2982 2362 2988 2363
rect 2910 2351 2916 2352
rect 2910 2347 2911 2351
rect 2915 2347 2916 2351
rect 2910 2346 2916 2347
rect 2984 2344 2986 2362
rect 3024 2352 3026 2369
rect 3464 2353 3466 2369
rect 3462 2352 3468 2353
rect 3022 2351 3028 2352
rect 3022 2347 3023 2351
rect 3027 2347 3028 2351
rect 3462 2348 3463 2352
rect 3467 2348 3468 2352
rect 3462 2347 3468 2348
rect 3022 2346 3028 2347
rect 2238 2343 2244 2344
rect 2238 2339 2239 2343
rect 2243 2339 2244 2343
rect 2238 2338 2244 2339
rect 2334 2343 2340 2344
rect 2334 2339 2335 2343
rect 2339 2339 2340 2343
rect 2334 2338 2340 2339
rect 2438 2343 2444 2344
rect 2438 2339 2439 2343
rect 2443 2339 2444 2343
rect 2438 2338 2444 2339
rect 2542 2343 2548 2344
rect 2542 2339 2543 2343
rect 2547 2339 2548 2343
rect 2542 2338 2548 2339
rect 2550 2343 2556 2344
rect 2550 2339 2551 2343
rect 2555 2339 2556 2343
rect 2550 2338 2556 2339
rect 2758 2343 2764 2344
rect 2758 2339 2759 2343
rect 2763 2339 2764 2343
rect 2758 2338 2764 2339
rect 2870 2343 2876 2344
rect 2870 2339 2871 2343
rect 2875 2339 2876 2343
rect 2870 2338 2876 2339
rect 2982 2343 2988 2344
rect 2982 2339 2983 2343
rect 2987 2339 2988 2343
rect 2982 2338 2988 2339
rect 2990 2343 2996 2344
rect 2990 2339 2991 2343
rect 2995 2339 2996 2343
rect 2990 2338 2996 2339
rect 2262 2332 2268 2333
rect 2262 2328 2263 2332
rect 2267 2328 2268 2332
rect 2262 2327 2268 2328
rect 2366 2332 2372 2333
rect 2366 2328 2367 2332
rect 2371 2328 2372 2332
rect 2366 2327 2372 2328
rect 2470 2332 2476 2333
rect 2470 2328 2471 2332
rect 2475 2328 2476 2332
rect 2470 2327 2476 2328
rect 2574 2332 2580 2333
rect 2574 2328 2575 2332
rect 2579 2328 2580 2332
rect 2574 2327 2580 2328
rect 2686 2332 2692 2333
rect 2686 2328 2687 2332
rect 2691 2328 2692 2332
rect 2686 2327 2692 2328
rect 2798 2332 2804 2333
rect 2798 2328 2799 2332
rect 2803 2328 2804 2332
rect 2798 2327 2804 2328
rect 2910 2332 2916 2333
rect 2910 2328 2911 2332
rect 2915 2328 2916 2332
rect 2910 2327 2916 2328
rect 2264 2303 2266 2327
rect 2368 2303 2370 2327
rect 2472 2303 2474 2327
rect 2576 2303 2578 2327
rect 2688 2303 2690 2327
rect 2800 2303 2802 2327
rect 2912 2303 2914 2327
rect 2263 2302 2267 2303
rect 2263 2297 2267 2298
rect 2367 2302 2371 2303
rect 2367 2297 2371 2298
rect 2375 2302 2379 2303
rect 2375 2297 2379 2298
rect 2471 2302 2475 2303
rect 2471 2297 2475 2298
rect 2551 2302 2555 2303
rect 2551 2297 2555 2298
rect 2575 2302 2579 2303
rect 2575 2297 2579 2298
rect 2687 2302 2691 2303
rect 2687 2297 2691 2298
rect 2719 2302 2723 2303
rect 2719 2297 2723 2298
rect 2799 2302 2803 2303
rect 2799 2297 2803 2298
rect 2887 2302 2891 2303
rect 2887 2297 2891 2298
rect 2911 2302 2915 2303
rect 2911 2297 2915 2298
rect 2230 2287 2236 2288
rect 2230 2283 2231 2287
rect 2235 2283 2236 2287
rect 2230 2282 2236 2283
rect 2376 2281 2378 2297
rect 2552 2281 2554 2297
rect 2720 2281 2722 2297
rect 2888 2281 2890 2297
rect 1886 2280 1892 2281
rect 1270 2275 1276 2276
rect 1766 2277 1772 2278
rect 1766 2273 1767 2277
rect 1771 2273 1772 2277
rect 1766 2272 1772 2273
rect 1806 2277 1812 2278
rect 1806 2273 1807 2277
rect 1811 2273 1812 2277
rect 1886 2276 1887 2280
rect 1891 2276 1892 2280
rect 1886 2275 1892 2276
rect 2038 2280 2044 2281
rect 2038 2276 2039 2280
rect 2043 2276 2044 2280
rect 2038 2275 2044 2276
rect 2198 2280 2204 2281
rect 2198 2276 2199 2280
rect 2203 2276 2204 2280
rect 2198 2275 2204 2276
rect 2374 2280 2380 2281
rect 2374 2276 2375 2280
rect 2379 2276 2380 2280
rect 2374 2275 2380 2276
rect 2550 2280 2556 2281
rect 2550 2276 2551 2280
rect 2555 2276 2556 2280
rect 2550 2275 2556 2276
rect 2718 2280 2724 2281
rect 2718 2276 2719 2280
rect 2723 2276 2724 2280
rect 2718 2275 2724 2276
rect 2886 2280 2892 2281
rect 2886 2276 2887 2280
rect 2891 2276 2892 2280
rect 2886 2275 2892 2276
rect 1806 2272 1812 2273
rect 1086 2271 1092 2272
rect 1086 2267 1087 2271
rect 1091 2267 1092 2271
rect 1086 2266 1092 2267
rect 1214 2271 1220 2272
rect 1214 2267 1215 2271
rect 1219 2267 1220 2271
rect 1214 2266 1220 2267
rect 1222 2271 1228 2272
rect 1222 2267 1223 2271
rect 1227 2267 1228 2271
rect 1222 2266 1228 2267
rect 1958 2271 1964 2272
rect 1958 2267 1959 2271
rect 1963 2267 1964 2271
rect 1958 2266 1964 2267
rect 2110 2271 2116 2272
rect 2110 2267 2111 2271
rect 2115 2267 2116 2271
rect 2110 2266 2116 2267
rect 2270 2271 2276 2272
rect 2270 2267 2271 2271
rect 2275 2267 2276 2271
rect 2270 2266 2276 2267
rect 2446 2271 2452 2272
rect 2446 2267 2447 2271
rect 2451 2267 2452 2271
rect 2446 2266 2452 2267
rect 2706 2271 2712 2272
rect 2706 2267 2707 2271
rect 2711 2267 2712 2271
rect 2706 2266 2712 2267
rect 2798 2271 2804 2272
rect 2798 2267 2799 2271
rect 2803 2267 2804 2271
rect 2798 2266 2804 2267
rect 1088 2244 1090 2266
rect 1142 2261 1148 2262
rect 1142 2257 1143 2261
rect 1147 2257 1148 2261
rect 1142 2256 1148 2257
rect 1068 2240 1074 2242
rect 1086 2243 1092 2244
rect 1068 2239 1069 2240
rect 1063 2238 1069 2239
rect 1086 2239 1087 2243
rect 1091 2239 1092 2243
rect 1086 2238 1092 2239
rect 1144 2235 1146 2256
rect 1216 2244 1218 2266
rect 1214 2243 1220 2244
rect 1214 2239 1215 2243
rect 1219 2239 1220 2243
rect 1214 2238 1220 2239
rect 951 2234 955 2235
rect 951 2229 955 2230
rect 1015 2234 1019 2235
rect 1015 2229 1019 2230
rect 1135 2234 1139 2235
rect 1135 2229 1139 2230
rect 1143 2234 1147 2235
rect 1143 2229 1147 2230
rect 952 2212 954 2229
rect 1078 2227 1084 2228
rect 1078 2223 1079 2227
rect 1083 2223 1084 2227
rect 1078 2222 1084 2223
rect 950 2211 956 2212
rect 950 2207 951 2211
rect 955 2207 956 2211
rect 950 2206 956 2207
rect 1080 2204 1082 2222
rect 1136 2212 1138 2229
rect 1224 2228 1226 2266
rect 1270 2261 1276 2262
rect 1886 2261 1892 2262
rect 1270 2257 1271 2261
rect 1275 2257 1276 2261
rect 1270 2256 1276 2257
rect 1766 2260 1772 2261
rect 1766 2256 1767 2260
rect 1771 2256 1772 2260
rect 1272 2235 1274 2256
rect 1766 2255 1772 2256
rect 1806 2260 1812 2261
rect 1806 2256 1807 2260
rect 1811 2256 1812 2260
rect 1886 2257 1887 2261
rect 1891 2257 1892 2261
rect 1886 2256 1892 2257
rect 1806 2255 1812 2256
rect 1768 2235 1770 2255
rect 1808 2239 1810 2255
rect 1888 2239 1890 2256
rect 1960 2244 1962 2266
rect 2038 2261 2044 2262
rect 2038 2257 2039 2261
rect 2043 2257 2044 2261
rect 2038 2256 2044 2257
rect 1950 2243 1956 2244
rect 1950 2239 1951 2243
rect 1955 2239 1956 2243
rect 1807 2238 1811 2239
rect 1271 2234 1275 2235
rect 1271 2229 1275 2230
rect 1319 2234 1323 2235
rect 1319 2229 1323 2230
rect 1503 2234 1507 2235
rect 1503 2229 1507 2230
rect 1671 2234 1675 2235
rect 1767 2234 1771 2235
rect 1671 2229 1675 2230
rect 1742 2231 1748 2232
rect 1222 2227 1228 2228
rect 1222 2223 1223 2227
rect 1227 2223 1228 2227
rect 1222 2222 1228 2223
rect 1302 2227 1308 2228
rect 1302 2223 1303 2227
rect 1307 2223 1308 2227
rect 1302 2222 1308 2223
rect 1134 2211 1140 2212
rect 1134 2207 1135 2211
rect 1139 2207 1140 2211
rect 1134 2206 1140 2207
rect 214 2203 220 2204
rect 214 2199 215 2203
rect 219 2199 220 2203
rect 214 2198 220 2199
rect 478 2203 484 2204
rect 478 2199 479 2203
rect 483 2199 484 2203
rect 478 2198 484 2199
rect 654 2203 660 2204
rect 654 2199 655 2203
rect 659 2199 660 2203
rect 654 2198 660 2199
rect 738 2203 744 2204
rect 738 2199 739 2203
rect 743 2199 744 2203
rect 738 2198 744 2199
rect 942 2203 948 2204
rect 942 2199 943 2203
rect 947 2199 948 2203
rect 942 2198 948 2199
rect 1078 2203 1084 2204
rect 1078 2199 1079 2203
rect 1083 2199 1084 2203
rect 1078 2198 1084 2199
rect 110 2195 116 2196
rect 110 2191 111 2195
rect 115 2191 116 2195
rect 198 2195 204 2196
rect 110 2190 116 2191
rect 134 2192 140 2193
rect 112 2163 114 2190
rect 134 2188 135 2192
rect 139 2188 140 2192
rect 198 2191 199 2195
rect 203 2191 204 2195
rect 198 2190 204 2191
rect 246 2192 252 2193
rect 134 2187 140 2188
rect 136 2163 138 2187
rect 111 2162 115 2163
rect 111 2157 115 2158
rect 135 2162 139 2163
rect 135 2157 139 2158
rect 112 2138 114 2157
rect 136 2141 138 2157
rect 134 2140 140 2141
rect 110 2137 116 2138
rect 110 2133 111 2137
rect 115 2133 116 2137
rect 134 2136 135 2140
rect 139 2136 140 2140
rect 134 2135 140 2136
rect 110 2132 116 2133
rect 134 2121 140 2122
rect 110 2120 116 2121
rect 110 2116 111 2120
rect 115 2116 116 2120
rect 134 2117 135 2121
rect 139 2117 140 2121
rect 134 2116 140 2117
rect 110 2115 116 2116
rect 112 2095 114 2115
rect 136 2095 138 2116
rect 200 2104 202 2190
rect 246 2188 247 2192
rect 251 2188 252 2192
rect 246 2187 252 2188
rect 406 2192 412 2193
rect 406 2188 407 2192
rect 411 2188 412 2192
rect 406 2187 412 2188
rect 582 2192 588 2193
rect 582 2188 583 2192
rect 587 2188 588 2192
rect 582 2187 588 2188
rect 766 2192 772 2193
rect 766 2188 767 2192
rect 771 2188 772 2192
rect 766 2187 772 2188
rect 950 2192 956 2193
rect 950 2188 951 2192
rect 955 2188 956 2192
rect 950 2187 956 2188
rect 1134 2192 1140 2193
rect 1134 2188 1135 2192
rect 1139 2188 1140 2192
rect 1134 2187 1140 2188
rect 248 2163 250 2187
rect 408 2163 410 2187
rect 584 2163 586 2187
rect 768 2163 770 2187
rect 952 2163 954 2187
rect 1136 2163 1138 2187
rect 247 2162 251 2163
rect 247 2157 251 2158
rect 391 2162 395 2163
rect 391 2157 395 2158
rect 407 2162 411 2163
rect 407 2157 411 2158
rect 543 2162 547 2163
rect 543 2157 547 2158
rect 583 2162 587 2163
rect 583 2157 587 2158
rect 695 2162 699 2163
rect 695 2157 699 2158
rect 767 2162 771 2163
rect 767 2157 771 2158
rect 839 2162 843 2163
rect 839 2157 843 2158
rect 951 2162 955 2163
rect 951 2157 955 2158
rect 975 2162 979 2163
rect 975 2157 979 2158
rect 1103 2162 1107 2163
rect 1103 2157 1107 2158
rect 1135 2162 1139 2163
rect 1135 2157 1139 2158
rect 1231 2162 1235 2163
rect 1231 2157 1235 2158
rect 248 2141 250 2157
rect 392 2141 394 2157
rect 544 2141 546 2157
rect 696 2141 698 2157
rect 840 2141 842 2157
rect 976 2141 978 2157
rect 1104 2141 1106 2157
rect 1232 2141 1234 2157
rect 246 2140 252 2141
rect 246 2136 247 2140
rect 251 2136 252 2140
rect 246 2135 252 2136
rect 390 2140 396 2141
rect 390 2136 391 2140
rect 395 2136 396 2140
rect 390 2135 396 2136
rect 542 2140 548 2141
rect 542 2136 543 2140
rect 547 2136 548 2140
rect 542 2135 548 2136
rect 694 2140 700 2141
rect 694 2136 695 2140
rect 699 2136 700 2140
rect 694 2135 700 2136
rect 838 2140 844 2141
rect 838 2136 839 2140
rect 843 2136 844 2140
rect 838 2135 844 2136
rect 974 2140 980 2141
rect 974 2136 975 2140
rect 979 2136 980 2140
rect 974 2135 980 2136
rect 1102 2140 1108 2141
rect 1102 2136 1103 2140
rect 1107 2136 1108 2140
rect 1102 2135 1108 2136
rect 1230 2140 1236 2141
rect 1230 2136 1231 2140
rect 1235 2136 1236 2140
rect 1230 2135 1236 2136
rect 1304 2132 1306 2222
rect 1320 2212 1322 2229
rect 1390 2227 1396 2228
rect 1390 2223 1391 2227
rect 1395 2223 1396 2227
rect 1390 2222 1396 2223
rect 1318 2211 1324 2212
rect 1318 2207 1319 2211
rect 1323 2207 1324 2211
rect 1318 2206 1324 2207
rect 1392 2204 1394 2222
rect 1504 2212 1506 2229
rect 1574 2227 1580 2228
rect 1574 2223 1575 2227
rect 1579 2223 1580 2227
rect 1574 2222 1580 2223
rect 1502 2211 1508 2212
rect 1502 2207 1503 2211
rect 1507 2207 1508 2211
rect 1502 2206 1508 2207
rect 1576 2204 1578 2222
rect 1672 2212 1674 2229
rect 1742 2227 1743 2231
rect 1747 2227 1748 2231
rect 1807 2233 1811 2234
rect 1831 2238 1835 2239
rect 1831 2233 1835 2234
rect 1887 2238 1891 2239
rect 1950 2238 1956 2239
rect 1958 2243 1964 2244
rect 1958 2239 1959 2243
rect 1963 2239 1964 2243
rect 2040 2239 2042 2256
rect 2112 2244 2114 2266
rect 2198 2261 2204 2262
rect 2198 2257 2199 2261
rect 2203 2257 2204 2261
rect 2198 2256 2204 2257
rect 2110 2243 2116 2244
rect 2110 2239 2111 2243
rect 2115 2239 2116 2243
rect 2200 2239 2202 2256
rect 2272 2244 2274 2266
rect 2374 2261 2380 2262
rect 2374 2257 2375 2261
rect 2379 2257 2380 2261
rect 2374 2256 2380 2257
rect 2270 2243 2276 2244
rect 2270 2239 2271 2243
rect 2275 2239 2276 2243
rect 2376 2239 2378 2256
rect 2448 2244 2450 2266
rect 2550 2261 2556 2262
rect 2550 2257 2551 2261
rect 2555 2257 2556 2261
rect 2550 2256 2556 2257
rect 2446 2243 2452 2244
rect 2446 2239 2447 2243
rect 2451 2239 2452 2243
rect 2552 2239 2554 2256
rect 1958 2238 1964 2239
rect 1967 2238 1971 2239
rect 1887 2233 1891 2234
rect 1767 2229 1771 2230
rect 1742 2226 1748 2227
rect 1670 2211 1676 2212
rect 1670 2207 1671 2211
rect 1675 2207 1676 2211
rect 1670 2206 1676 2207
rect 1744 2204 1746 2226
rect 1768 2213 1770 2229
rect 1808 2217 1810 2233
rect 1806 2216 1812 2217
rect 1832 2216 1834 2233
rect 1902 2231 1908 2232
rect 1902 2227 1903 2231
rect 1907 2227 1908 2231
rect 1902 2226 1908 2227
rect 1766 2212 1772 2213
rect 1766 2208 1767 2212
rect 1771 2208 1772 2212
rect 1806 2212 1807 2216
rect 1811 2212 1812 2216
rect 1806 2211 1812 2212
rect 1830 2215 1836 2216
rect 1830 2211 1831 2215
rect 1835 2211 1836 2215
rect 1830 2210 1836 2211
rect 1904 2208 1906 2226
rect 1766 2207 1772 2208
rect 1902 2207 1908 2208
rect 1390 2203 1396 2204
rect 1390 2199 1391 2203
rect 1395 2199 1396 2203
rect 1390 2198 1396 2199
rect 1574 2203 1580 2204
rect 1574 2199 1575 2203
rect 1579 2199 1580 2203
rect 1574 2198 1580 2199
rect 1742 2203 1748 2204
rect 1742 2199 1743 2203
rect 1747 2199 1748 2203
rect 1902 2203 1903 2207
rect 1907 2203 1908 2207
rect 1902 2202 1908 2203
rect 1742 2198 1748 2199
rect 1806 2199 1812 2200
rect 1766 2195 1772 2196
rect 1318 2192 1324 2193
rect 1318 2188 1319 2192
rect 1323 2188 1324 2192
rect 1318 2187 1324 2188
rect 1502 2192 1508 2193
rect 1502 2188 1503 2192
rect 1507 2188 1508 2192
rect 1502 2187 1508 2188
rect 1670 2192 1676 2193
rect 1670 2188 1671 2192
rect 1675 2188 1676 2192
rect 1766 2191 1767 2195
rect 1771 2191 1772 2195
rect 1806 2195 1807 2199
rect 1811 2195 1812 2199
rect 1806 2194 1812 2195
rect 1830 2196 1836 2197
rect 1766 2190 1772 2191
rect 1670 2187 1676 2188
rect 1320 2163 1322 2187
rect 1504 2163 1506 2187
rect 1672 2163 1674 2187
rect 1768 2163 1770 2190
rect 1808 2175 1810 2194
rect 1830 2192 1831 2196
rect 1835 2192 1836 2196
rect 1830 2191 1836 2192
rect 1832 2175 1834 2191
rect 1952 2188 1954 2238
rect 1967 2233 1971 2234
rect 2039 2238 2043 2239
rect 2110 2238 2116 2239
rect 2135 2238 2139 2239
rect 2039 2233 2043 2234
rect 2135 2233 2139 2234
rect 2199 2238 2203 2239
rect 2270 2238 2276 2239
rect 2311 2238 2315 2239
rect 2199 2233 2203 2234
rect 2311 2233 2315 2234
rect 2375 2238 2379 2239
rect 2446 2238 2452 2239
rect 2487 2238 2491 2239
rect 2375 2233 2379 2234
rect 2487 2233 2491 2234
rect 2551 2238 2555 2239
rect 2551 2233 2555 2234
rect 2655 2238 2659 2239
rect 2655 2233 2659 2234
rect 1968 2216 1970 2233
rect 2136 2216 2138 2233
rect 2206 2231 2212 2232
rect 2206 2227 2207 2231
rect 2211 2227 2212 2231
rect 2206 2226 2212 2227
rect 1966 2215 1972 2216
rect 1966 2211 1967 2215
rect 1971 2211 1972 2215
rect 1966 2210 1972 2211
rect 2134 2215 2140 2216
rect 2134 2211 2135 2215
rect 2139 2211 2140 2215
rect 2134 2210 2140 2211
rect 2208 2208 2210 2226
rect 2312 2216 2314 2233
rect 2382 2231 2388 2232
rect 2382 2227 2383 2231
rect 2387 2227 2388 2231
rect 2382 2226 2388 2227
rect 2310 2215 2316 2216
rect 2310 2211 2311 2215
rect 2315 2211 2316 2215
rect 2310 2210 2316 2211
rect 2384 2208 2386 2226
rect 2488 2216 2490 2233
rect 2656 2216 2658 2233
rect 2708 2232 2710 2266
rect 2718 2261 2724 2262
rect 2718 2257 2719 2261
rect 2723 2257 2724 2261
rect 2718 2256 2724 2257
rect 2720 2239 2722 2256
rect 2800 2244 2802 2266
rect 2886 2261 2892 2262
rect 2886 2257 2887 2261
rect 2891 2257 2892 2261
rect 2886 2256 2892 2257
rect 2798 2243 2804 2244
rect 2798 2239 2799 2243
rect 2803 2239 2804 2243
rect 2888 2239 2890 2256
rect 2992 2244 2994 2338
rect 3462 2335 3468 2336
rect 3022 2332 3028 2333
rect 3022 2328 3023 2332
rect 3027 2328 3028 2332
rect 3462 2331 3463 2335
rect 3467 2331 3468 2335
rect 3462 2330 3468 2331
rect 3022 2327 3028 2328
rect 3024 2303 3026 2327
rect 3464 2303 3466 2330
rect 3023 2302 3027 2303
rect 3023 2297 3027 2298
rect 3055 2302 3059 2303
rect 3055 2297 3059 2298
rect 3223 2302 3227 2303
rect 3223 2297 3227 2298
rect 3367 2302 3371 2303
rect 3367 2297 3371 2298
rect 3463 2302 3467 2303
rect 3463 2297 3467 2298
rect 3056 2281 3058 2297
rect 3224 2281 3226 2297
rect 3368 2281 3370 2297
rect 3054 2280 3060 2281
rect 3054 2276 3055 2280
rect 3059 2276 3060 2280
rect 3054 2275 3060 2276
rect 3222 2280 3228 2281
rect 3222 2276 3223 2280
rect 3227 2276 3228 2280
rect 3222 2275 3228 2276
rect 3366 2280 3372 2281
rect 3366 2276 3367 2280
rect 3371 2276 3372 2280
rect 3464 2278 3466 2297
rect 3366 2275 3372 2276
rect 3462 2277 3468 2278
rect 3462 2273 3463 2277
rect 3467 2273 3468 2277
rect 3462 2272 3468 2273
rect 3126 2271 3132 2272
rect 3126 2267 3127 2271
rect 3131 2267 3132 2271
rect 3126 2266 3132 2267
rect 3294 2271 3300 2272
rect 3294 2267 3295 2271
rect 3299 2267 3300 2271
rect 3294 2266 3300 2267
rect 3430 2271 3436 2272
rect 3430 2267 3431 2271
rect 3435 2267 3436 2271
rect 3430 2266 3436 2267
rect 3054 2261 3060 2262
rect 3054 2257 3055 2261
rect 3059 2257 3060 2261
rect 3054 2256 3060 2257
rect 2990 2243 2996 2244
rect 2990 2239 2991 2243
rect 2995 2239 2996 2243
rect 2719 2238 2723 2239
rect 2798 2238 2804 2239
rect 2815 2238 2819 2239
rect 2719 2233 2723 2234
rect 2815 2233 2819 2234
rect 2887 2238 2891 2239
rect 2887 2233 2891 2234
rect 2959 2238 2963 2239
rect 2990 2238 2996 2239
rect 3030 2243 3036 2244
rect 3030 2239 3031 2243
rect 3035 2239 3036 2243
rect 3056 2239 3058 2256
rect 3128 2244 3130 2266
rect 3222 2261 3228 2262
rect 3222 2257 3223 2261
rect 3227 2257 3228 2261
rect 3222 2256 3228 2257
rect 3126 2243 3132 2244
rect 3126 2239 3127 2243
rect 3131 2239 3132 2243
rect 3224 2239 3226 2256
rect 3296 2244 3298 2266
rect 3366 2261 3372 2262
rect 3366 2257 3367 2261
rect 3371 2257 3372 2261
rect 3366 2256 3372 2257
rect 3294 2243 3300 2244
rect 3294 2239 3295 2243
rect 3299 2239 3300 2243
rect 3368 2239 3370 2256
rect 3030 2238 3036 2239
rect 3055 2238 3059 2239
rect 2959 2233 2963 2234
rect 2706 2231 2712 2232
rect 2706 2227 2707 2231
rect 2711 2227 2712 2231
rect 2706 2226 2712 2227
rect 2726 2231 2732 2232
rect 2726 2227 2727 2231
rect 2731 2227 2732 2231
rect 2726 2226 2732 2227
rect 2486 2215 2492 2216
rect 2486 2211 2487 2215
rect 2491 2211 2492 2215
rect 2486 2210 2492 2211
rect 2654 2215 2660 2216
rect 2654 2211 2655 2215
rect 2659 2211 2660 2215
rect 2654 2210 2660 2211
rect 2728 2208 2730 2226
rect 2816 2216 2818 2233
rect 2960 2216 2962 2233
rect 2814 2215 2820 2216
rect 2814 2211 2815 2215
rect 2819 2211 2820 2215
rect 2814 2210 2820 2211
rect 2958 2215 2964 2216
rect 2958 2211 2959 2215
rect 2963 2211 2964 2215
rect 2958 2210 2964 2211
rect 3032 2208 3034 2238
rect 3055 2233 3059 2234
rect 3103 2238 3107 2239
rect 3126 2238 3132 2239
rect 3223 2238 3227 2239
rect 3103 2233 3107 2234
rect 3223 2233 3227 2234
rect 3247 2238 3251 2239
rect 3294 2238 3300 2239
rect 3367 2238 3371 2239
rect 3247 2233 3251 2234
rect 3367 2233 3371 2234
rect 3038 2231 3044 2232
rect 3038 2227 3039 2231
rect 3043 2227 3044 2231
rect 3038 2226 3044 2227
rect 3040 2208 3042 2226
rect 3104 2216 3106 2233
rect 3182 2231 3188 2232
rect 3182 2227 3183 2231
rect 3187 2227 3188 2231
rect 3182 2226 3188 2227
rect 3102 2215 3108 2216
rect 3102 2211 3103 2215
rect 3107 2211 3108 2215
rect 3102 2210 3108 2211
rect 3184 2208 3186 2226
rect 3248 2216 3250 2233
rect 3368 2216 3370 2233
rect 3432 2232 3434 2266
rect 3462 2260 3468 2261
rect 3462 2256 3463 2260
rect 3467 2256 3468 2260
rect 3462 2255 3468 2256
rect 3464 2239 3466 2255
rect 3463 2238 3467 2239
rect 3463 2233 3467 2234
rect 3430 2231 3436 2232
rect 3430 2227 3431 2231
rect 3435 2227 3436 2231
rect 3430 2226 3436 2227
rect 3464 2217 3466 2233
rect 3462 2216 3468 2217
rect 3246 2215 3252 2216
rect 3246 2211 3247 2215
rect 3251 2211 3252 2215
rect 3246 2210 3252 2211
rect 3366 2215 3372 2216
rect 3366 2211 3367 2215
rect 3371 2211 3372 2215
rect 3462 2212 3463 2216
rect 3467 2212 3468 2216
rect 3462 2211 3468 2212
rect 3366 2210 3372 2211
rect 2206 2207 2212 2208
rect 2206 2203 2207 2207
rect 2211 2203 2212 2207
rect 2206 2202 2212 2203
rect 2382 2207 2388 2208
rect 2382 2203 2383 2207
rect 2387 2203 2388 2207
rect 2382 2202 2388 2203
rect 2418 2207 2424 2208
rect 2418 2203 2419 2207
rect 2423 2203 2424 2207
rect 2418 2202 2424 2203
rect 2726 2207 2732 2208
rect 2726 2203 2727 2207
rect 2731 2203 2732 2207
rect 3030 2207 3036 2208
rect 2726 2202 2732 2203
rect 2886 2203 2892 2204
rect 1966 2196 1972 2197
rect 1966 2192 1967 2196
rect 1971 2192 1972 2196
rect 1966 2191 1972 2192
rect 2134 2196 2140 2197
rect 2134 2192 2135 2196
rect 2139 2192 2140 2196
rect 2134 2191 2140 2192
rect 2310 2196 2316 2197
rect 2310 2192 2311 2196
rect 2315 2192 2316 2196
rect 2310 2191 2316 2192
rect 1950 2187 1956 2188
rect 1950 2183 1951 2187
rect 1955 2183 1956 2187
rect 1950 2182 1956 2183
rect 1968 2175 1970 2191
rect 2136 2175 2138 2191
rect 2312 2175 2314 2191
rect 2420 2188 2422 2202
rect 2886 2199 2887 2203
rect 2891 2199 2892 2203
rect 3030 2203 3031 2207
rect 3035 2203 3036 2207
rect 3030 2202 3036 2203
rect 3038 2207 3044 2208
rect 3038 2203 3039 2207
rect 3043 2203 3044 2207
rect 3038 2202 3044 2203
rect 3182 2207 3188 2208
rect 3182 2203 3183 2207
rect 3187 2203 3188 2207
rect 3182 2202 3188 2203
rect 3438 2203 3444 2204
rect 2886 2198 2892 2199
rect 3438 2199 3439 2203
rect 3443 2199 3444 2203
rect 3438 2198 3444 2199
rect 3462 2199 3468 2200
rect 2486 2196 2492 2197
rect 2486 2192 2487 2196
rect 2491 2192 2492 2196
rect 2486 2191 2492 2192
rect 2654 2196 2660 2197
rect 2654 2192 2655 2196
rect 2659 2192 2660 2196
rect 2654 2191 2660 2192
rect 2814 2196 2820 2197
rect 2814 2192 2815 2196
rect 2819 2192 2820 2196
rect 2814 2191 2820 2192
rect 2418 2187 2424 2188
rect 2418 2183 2419 2187
rect 2423 2183 2424 2187
rect 2418 2182 2424 2183
rect 2488 2175 2490 2191
rect 2656 2175 2658 2191
rect 2816 2175 2818 2191
rect 1807 2174 1811 2175
rect 1807 2169 1811 2170
rect 1831 2174 1835 2175
rect 1831 2169 1835 2170
rect 1967 2174 1971 2175
rect 1967 2169 1971 2170
rect 2135 2174 2139 2175
rect 2135 2169 2139 2170
rect 2311 2174 2315 2175
rect 2311 2169 2315 2170
rect 2487 2174 2491 2175
rect 2487 2169 2491 2170
rect 2655 2174 2659 2175
rect 2655 2169 2659 2170
rect 2815 2174 2819 2175
rect 2815 2169 2819 2170
rect 1319 2162 1323 2163
rect 1319 2157 1323 2158
rect 1351 2162 1355 2163
rect 1351 2157 1355 2158
rect 1463 2162 1467 2163
rect 1463 2157 1467 2158
rect 1503 2162 1507 2163
rect 1503 2157 1507 2158
rect 1575 2162 1579 2163
rect 1575 2157 1579 2158
rect 1671 2162 1675 2163
rect 1671 2157 1675 2158
rect 1767 2162 1771 2163
rect 1767 2157 1771 2158
rect 1352 2141 1354 2157
rect 1464 2141 1466 2157
rect 1576 2141 1578 2157
rect 1672 2141 1674 2157
rect 1350 2140 1356 2141
rect 1350 2136 1351 2140
rect 1355 2136 1356 2140
rect 1350 2135 1356 2136
rect 1462 2140 1468 2141
rect 1462 2136 1463 2140
rect 1467 2136 1468 2140
rect 1462 2135 1468 2136
rect 1574 2140 1580 2141
rect 1574 2136 1575 2140
rect 1579 2136 1580 2140
rect 1574 2135 1580 2136
rect 1670 2140 1676 2141
rect 1670 2136 1671 2140
rect 1675 2136 1676 2140
rect 1768 2138 1770 2157
rect 1808 2150 1810 2169
rect 1806 2149 1812 2150
rect 1806 2145 1807 2149
rect 1811 2145 1812 2149
rect 1806 2144 1812 2145
rect 1670 2135 1676 2136
rect 1766 2137 1772 2138
rect 1766 2133 1767 2137
rect 1771 2133 1772 2137
rect 1766 2132 1772 2133
rect 1806 2132 1812 2133
rect 206 2131 212 2132
rect 206 2127 207 2131
rect 211 2127 212 2131
rect 206 2126 212 2127
rect 318 2131 324 2132
rect 318 2127 319 2131
rect 323 2127 324 2131
rect 318 2126 324 2127
rect 462 2131 468 2132
rect 462 2127 463 2131
rect 467 2127 468 2131
rect 462 2126 468 2127
rect 614 2131 620 2132
rect 614 2127 615 2131
rect 619 2127 620 2131
rect 614 2126 620 2127
rect 622 2131 628 2132
rect 622 2127 623 2131
rect 627 2127 628 2131
rect 622 2126 628 2127
rect 950 2131 956 2132
rect 950 2127 951 2131
rect 955 2127 956 2131
rect 950 2126 956 2127
rect 1054 2131 1060 2132
rect 1054 2127 1055 2131
rect 1059 2127 1060 2131
rect 1054 2126 1060 2127
rect 1174 2131 1180 2132
rect 1174 2127 1175 2131
rect 1179 2127 1180 2131
rect 1174 2126 1180 2127
rect 1302 2131 1308 2132
rect 1302 2127 1303 2131
rect 1307 2127 1308 2131
rect 1302 2126 1308 2127
rect 1310 2131 1316 2132
rect 1310 2127 1311 2131
rect 1315 2127 1316 2131
rect 1310 2126 1316 2127
rect 1430 2131 1436 2132
rect 1430 2127 1431 2131
rect 1435 2127 1436 2131
rect 1430 2126 1436 2127
rect 1542 2131 1548 2132
rect 1542 2127 1543 2131
rect 1547 2127 1548 2131
rect 1542 2126 1548 2127
rect 1654 2131 1660 2132
rect 1654 2127 1655 2131
rect 1659 2127 1660 2131
rect 1806 2128 1807 2132
rect 1811 2128 1812 2132
rect 1806 2127 1812 2128
rect 1654 2126 1660 2127
rect 208 2104 210 2126
rect 246 2121 252 2122
rect 246 2117 247 2121
rect 251 2117 252 2121
rect 246 2116 252 2117
rect 198 2103 204 2104
rect 198 2099 199 2103
rect 203 2099 204 2103
rect 198 2098 204 2099
rect 206 2103 212 2104
rect 206 2099 207 2103
rect 211 2099 212 2103
rect 206 2098 212 2099
rect 248 2095 250 2116
rect 320 2104 322 2126
rect 390 2121 396 2122
rect 390 2117 391 2121
rect 395 2117 396 2121
rect 390 2116 396 2117
rect 318 2103 324 2104
rect 318 2099 319 2103
rect 323 2099 324 2103
rect 318 2098 324 2099
rect 392 2095 394 2116
rect 464 2104 466 2126
rect 542 2121 548 2122
rect 542 2117 543 2121
rect 547 2117 548 2121
rect 542 2116 548 2117
rect 462 2103 468 2104
rect 462 2099 463 2103
rect 467 2099 468 2103
rect 462 2098 468 2099
rect 544 2095 546 2116
rect 616 2104 618 2126
rect 614 2103 620 2104
rect 614 2099 615 2103
rect 619 2099 620 2103
rect 614 2098 620 2099
rect 624 2096 626 2126
rect 694 2121 700 2122
rect 694 2117 695 2121
rect 699 2117 700 2121
rect 694 2116 700 2117
rect 838 2121 844 2122
rect 838 2117 839 2121
rect 843 2117 844 2121
rect 838 2116 844 2117
rect 622 2095 628 2096
rect 696 2095 698 2116
rect 840 2095 842 2116
rect 952 2104 954 2126
rect 974 2121 980 2122
rect 974 2117 975 2121
rect 979 2117 980 2121
rect 974 2116 980 2117
rect 950 2103 956 2104
rect 950 2099 951 2103
rect 955 2099 956 2103
rect 950 2098 956 2099
rect 976 2095 978 2116
rect 111 2094 115 2095
rect 111 2089 115 2090
rect 135 2094 139 2095
rect 135 2089 139 2090
rect 223 2094 227 2095
rect 223 2089 227 2090
rect 247 2094 251 2095
rect 247 2089 251 2090
rect 343 2094 347 2095
rect 343 2089 347 2090
rect 391 2094 395 2095
rect 391 2089 395 2090
rect 463 2094 467 2095
rect 463 2089 467 2090
rect 543 2094 547 2095
rect 543 2089 547 2090
rect 583 2094 587 2095
rect 622 2091 623 2095
rect 627 2091 628 2095
rect 622 2090 628 2091
rect 695 2094 699 2095
rect 583 2089 587 2090
rect 695 2089 699 2090
rect 703 2094 707 2095
rect 703 2089 707 2090
rect 823 2094 827 2095
rect 823 2089 827 2090
rect 839 2094 843 2095
rect 839 2089 843 2090
rect 935 2094 939 2095
rect 935 2089 939 2090
rect 975 2094 979 2095
rect 975 2089 979 2090
rect 1047 2094 1051 2095
rect 1047 2089 1051 2090
rect 112 2073 114 2089
rect 110 2072 116 2073
rect 136 2072 138 2089
rect 224 2072 226 2089
rect 294 2087 300 2088
rect 294 2083 295 2087
rect 299 2083 300 2087
rect 294 2082 300 2083
rect 110 2068 111 2072
rect 115 2068 116 2072
rect 110 2067 116 2068
rect 134 2071 140 2072
rect 134 2067 135 2071
rect 139 2067 140 2071
rect 134 2066 140 2067
rect 222 2071 228 2072
rect 222 2067 223 2071
rect 227 2067 228 2071
rect 222 2066 228 2067
rect 296 2064 298 2082
rect 344 2072 346 2089
rect 414 2087 420 2088
rect 414 2083 415 2087
rect 419 2083 420 2087
rect 414 2082 420 2083
rect 342 2071 348 2072
rect 342 2067 343 2071
rect 347 2067 348 2071
rect 342 2066 348 2067
rect 416 2064 418 2082
rect 464 2072 466 2089
rect 534 2087 540 2088
rect 534 2083 535 2087
rect 539 2083 540 2087
rect 534 2082 540 2083
rect 462 2071 468 2072
rect 462 2067 463 2071
rect 467 2067 468 2071
rect 462 2066 468 2067
rect 536 2064 538 2082
rect 584 2072 586 2089
rect 704 2072 706 2089
rect 754 2087 760 2088
rect 754 2083 755 2087
rect 759 2083 760 2087
rect 754 2082 760 2083
rect 774 2087 780 2088
rect 774 2083 775 2087
rect 779 2083 780 2087
rect 774 2082 780 2083
rect 582 2071 588 2072
rect 582 2067 583 2071
rect 587 2067 588 2071
rect 582 2066 588 2067
rect 702 2071 708 2072
rect 702 2067 703 2071
rect 707 2067 708 2071
rect 702 2066 708 2067
rect 294 2063 300 2064
rect 294 2059 295 2063
rect 299 2059 300 2063
rect 294 2058 300 2059
rect 414 2063 420 2064
rect 414 2059 415 2063
rect 419 2059 420 2063
rect 414 2058 420 2059
rect 534 2063 540 2064
rect 534 2059 535 2063
rect 539 2059 540 2063
rect 534 2058 540 2059
rect 542 2063 548 2064
rect 542 2059 543 2063
rect 547 2059 548 2063
rect 542 2058 548 2059
rect 110 2055 116 2056
rect 110 2051 111 2055
rect 115 2051 116 2055
rect 110 2050 116 2051
rect 134 2052 140 2053
rect 112 2023 114 2050
rect 134 2048 135 2052
rect 139 2048 140 2052
rect 134 2047 140 2048
rect 222 2052 228 2053
rect 222 2048 223 2052
rect 227 2048 228 2052
rect 222 2047 228 2048
rect 342 2052 348 2053
rect 342 2048 343 2052
rect 347 2048 348 2052
rect 342 2047 348 2048
rect 462 2052 468 2053
rect 462 2048 463 2052
rect 467 2048 468 2052
rect 462 2047 468 2048
rect 136 2023 138 2047
rect 224 2023 226 2047
rect 344 2023 346 2047
rect 464 2023 466 2047
rect 111 2022 115 2023
rect 111 2017 115 2018
rect 135 2022 139 2023
rect 135 2017 139 2018
rect 223 2022 227 2023
rect 223 2017 227 2018
rect 239 2022 243 2023
rect 239 2017 243 2018
rect 343 2022 347 2023
rect 343 2017 347 2018
rect 367 2022 371 2023
rect 367 2017 371 2018
rect 463 2022 467 2023
rect 463 2017 467 2018
rect 503 2022 507 2023
rect 503 2017 507 2018
rect 112 1998 114 2017
rect 136 2001 138 2017
rect 186 2015 192 2016
rect 186 2011 187 2015
rect 191 2011 192 2015
rect 186 2010 192 2011
rect 134 2000 140 2001
rect 110 1997 116 1998
rect 110 1993 111 1997
rect 115 1993 116 1997
rect 134 1996 135 2000
rect 139 1996 140 2000
rect 134 1995 140 1996
rect 110 1992 116 1993
rect 134 1981 140 1982
rect 110 1980 116 1981
rect 110 1976 111 1980
rect 115 1976 116 1980
rect 134 1977 135 1981
rect 139 1977 140 1981
rect 134 1976 140 1977
rect 110 1975 116 1976
rect 112 1955 114 1975
rect 136 1955 138 1976
rect 188 1964 190 2010
rect 240 2001 242 2017
rect 368 2001 370 2017
rect 504 2001 506 2017
rect 544 2016 546 2058
rect 582 2052 588 2053
rect 582 2048 583 2052
rect 587 2048 588 2052
rect 582 2047 588 2048
rect 702 2052 708 2053
rect 702 2048 703 2052
rect 707 2048 708 2052
rect 702 2047 708 2048
rect 584 2023 586 2047
rect 704 2023 706 2047
rect 583 2022 587 2023
rect 583 2017 587 2018
rect 639 2022 643 2023
rect 639 2017 643 2018
rect 703 2022 707 2023
rect 703 2017 707 2018
rect 542 2015 548 2016
rect 542 2011 543 2015
rect 547 2011 548 2015
rect 542 2010 548 2011
rect 640 2001 642 2017
rect 238 2000 244 2001
rect 238 1996 239 2000
rect 243 1996 244 2000
rect 238 1995 244 1996
rect 366 2000 372 2001
rect 366 1996 367 2000
rect 371 1996 372 2000
rect 366 1995 372 1996
rect 502 2000 508 2001
rect 502 1996 503 2000
rect 507 1996 508 2000
rect 502 1995 508 1996
rect 638 2000 644 2001
rect 638 1996 639 2000
rect 643 1996 644 2000
rect 638 1995 644 1996
rect 756 1992 758 2082
rect 776 2064 778 2082
rect 824 2072 826 2089
rect 894 2087 900 2088
rect 894 2083 895 2087
rect 899 2083 900 2087
rect 894 2082 900 2083
rect 822 2071 828 2072
rect 822 2067 823 2071
rect 827 2067 828 2071
rect 822 2066 828 2067
rect 896 2064 898 2082
rect 936 2072 938 2089
rect 1048 2072 1050 2089
rect 1056 2088 1058 2126
rect 1102 2121 1108 2122
rect 1102 2117 1103 2121
rect 1107 2117 1108 2121
rect 1102 2116 1108 2117
rect 1104 2095 1106 2116
rect 1176 2104 1178 2126
rect 1230 2121 1236 2122
rect 1230 2117 1231 2121
rect 1235 2117 1236 2121
rect 1230 2116 1236 2117
rect 1174 2103 1180 2104
rect 1174 2099 1175 2103
rect 1179 2099 1180 2103
rect 1174 2098 1180 2099
rect 1232 2095 1234 2116
rect 1312 2096 1314 2126
rect 1350 2121 1356 2122
rect 1350 2117 1351 2121
rect 1355 2117 1356 2121
rect 1350 2116 1356 2117
rect 1310 2095 1316 2096
rect 1352 2095 1354 2116
rect 1432 2104 1434 2126
rect 1462 2121 1468 2122
rect 1462 2117 1463 2121
rect 1467 2117 1468 2121
rect 1462 2116 1468 2117
rect 1430 2103 1436 2104
rect 1430 2099 1431 2103
rect 1435 2099 1436 2103
rect 1430 2098 1436 2099
rect 1464 2095 1466 2116
rect 1544 2104 1546 2126
rect 1574 2121 1580 2122
rect 1574 2117 1575 2121
rect 1579 2117 1580 2121
rect 1574 2116 1580 2117
rect 1542 2103 1548 2104
rect 1542 2099 1543 2103
rect 1547 2099 1548 2103
rect 1542 2098 1548 2099
rect 1576 2095 1578 2116
rect 1656 2104 1658 2126
rect 1670 2121 1676 2122
rect 1670 2117 1671 2121
rect 1675 2117 1676 2121
rect 1670 2116 1676 2117
rect 1766 2120 1772 2121
rect 1766 2116 1767 2120
rect 1771 2116 1772 2120
rect 1654 2103 1660 2104
rect 1654 2099 1655 2103
rect 1659 2099 1660 2103
rect 1654 2098 1660 2099
rect 1672 2095 1674 2116
rect 1766 2115 1772 2116
rect 1768 2095 1770 2115
rect 1786 2103 1792 2104
rect 1808 2103 1810 2127
rect 2888 2116 2890 2198
rect 2958 2196 2964 2197
rect 2958 2192 2959 2196
rect 2963 2192 2964 2196
rect 2958 2191 2964 2192
rect 3102 2196 3108 2197
rect 3102 2192 3103 2196
rect 3107 2192 3108 2196
rect 3102 2191 3108 2192
rect 3246 2196 3252 2197
rect 3246 2192 3247 2196
rect 3251 2192 3252 2196
rect 3246 2191 3252 2192
rect 3366 2196 3372 2197
rect 3366 2192 3367 2196
rect 3371 2192 3372 2196
rect 3366 2191 3372 2192
rect 2960 2175 2962 2191
rect 3104 2175 3106 2191
rect 3248 2175 3250 2191
rect 3368 2175 3370 2191
rect 2927 2174 2931 2175
rect 2927 2169 2931 2170
rect 2959 2174 2963 2175
rect 2959 2169 2963 2170
rect 3015 2174 3019 2175
rect 3015 2169 3019 2170
rect 3103 2174 3107 2175
rect 3103 2169 3107 2170
rect 3191 2174 3195 2175
rect 3191 2169 3195 2170
rect 3247 2174 3251 2175
rect 3247 2169 3251 2170
rect 3279 2174 3283 2175
rect 3279 2169 3283 2170
rect 3367 2174 3371 2175
rect 3367 2169 3371 2170
rect 2928 2153 2930 2169
rect 3016 2153 3018 2169
rect 3104 2153 3106 2169
rect 3192 2153 3194 2169
rect 3280 2153 3282 2169
rect 3368 2153 3370 2169
rect 2926 2152 2932 2153
rect 2926 2148 2927 2152
rect 2931 2148 2932 2152
rect 2926 2147 2932 2148
rect 3014 2152 3020 2153
rect 3014 2148 3015 2152
rect 3019 2148 3020 2152
rect 3014 2147 3020 2148
rect 3102 2152 3108 2153
rect 3102 2148 3103 2152
rect 3107 2148 3108 2152
rect 3102 2147 3108 2148
rect 3190 2152 3196 2153
rect 3190 2148 3191 2152
rect 3195 2148 3196 2152
rect 3190 2147 3196 2148
rect 3278 2152 3284 2153
rect 3278 2148 3279 2152
rect 3283 2148 3284 2152
rect 3278 2147 3284 2148
rect 3366 2152 3372 2153
rect 3366 2148 3367 2152
rect 3371 2148 3372 2152
rect 3366 2147 3372 2148
rect 2998 2143 3004 2144
rect 2998 2139 2999 2143
rect 3003 2139 3004 2143
rect 2998 2138 3004 2139
rect 3086 2143 3092 2144
rect 3086 2139 3087 2143
rect 3091 2139 3092 2143
rect 3086 2138 3092 2139
rect 3254 2143 3260 2144
rect 3254 2139 3255 2143
rect 3259 2139 3260 2143
rect 3254 2138 3260 2139
rect 3350 2143 3356 2144
rect 3350 2139 3351 2143
rect 3355 2139 3356 2143
rect 3350 2138 3356 2139
rect 3358 2143 3364 2144
rect 3358 2139 3359 2143
rect 3363 2139 3364 2143
rect 3358 2138 3364 2139
rect 2926 2133 2932 2134
rect 2926 2129 2927 2133
rect 2931 2129 2932 2133
rect 2926 2128 2932 2129
rect 2886 2115 2892 2116
rect 2886 2111 2887 2115
rect 2891 2111 2892 2115
rect 2886 2110 2892 2111
rect 2928 2103 2930 2128
rect 3000 2116 3002 2138
rect 3014 2133 3020 2134
rect 3014 2129 3015 2133
rect 3019 2129 3020 2133
rect 3014 2128 3020 2129
rect 2998 2115 3004 2116
rect 2998 2111 2999 2115
rect 3003 2111 3004 2115
rect 2998 2110 3004 2111
rect 3016 2103 3018 2128
rect 3088 2116 3090 2138
rect 3102 2133 3108 2134
rect 3102 2129 3103 2133
rect 3107 2129 3108 2133
rect 3102 2128 3108 2129
rect 3190 2133 3196 2134
rect 3190 2129 3191 2133
rect 3195 2129 3196 2133
rect 3190 2128 3196 2129
rect 3086 2115 3092 2116
rect 3086 2111 3087 2115
rect 3091 2111 3092 2115
rect 3086 2110 3092 2111
rect 3104 2103 3106 2128
rect 3192 2103 3194 2128
rect 3256 2104 3258 2138
rect 3278 2133 3284 2134
rect 3278 2129 3279 2133
rect 3283 2129 3284 2133
rect 3278 2128 3284 2129
rect 3254 2103 3260 2104
rect 3280 2103 3282 2128
rect 1786 2099 1787 2103
rect 1791 2099 1792 2103
rect 1786 2098 1792 2099
rect 1807 2102 1811 2103
rect 1103 2094 1107 2095
rect 1103 2089 1107 2090
rect 1159 2094 1163 2095
rect 1159 2089 1163 2090
rect 1231 2094 1235 2095
rect 1231 2089 1235 2090
rect 1279 2094 1283 2095
rect 1310 2091 1311 2095
rect 1315 2091 1316 2095
rect 1310 2090 1316 2091
rect 1351 2094 1355 2095
rect 1279 2089 1283 2090
rect 1351 2089 1355 2090
rect 1463 2094 1467 2095
rect 1463 2089 1467 2090
rect 1575 2094 1579 2095
rect 1575 2089 1579 2090
rect 1671 2094 1675 2095
rect 1671 2089 1675 2090
rect 1767 2094 1771 2095
rect 1767 2089 1771 2090
rect 1054 2087 1060 2088
rect 1054 2083 1055 2087
rect 1059 2083 1060 2087
rect 1054 2082 1060 2083
rect 1118 2087 1124 2088
rect 1118 2083 1119 2087
rect 1123 2083 1124 2087
rect 1118 2082 1124 2083
rect 934 2071 940 2072
rect 934 2067 935 2071
rect 939 2067 940 2071
rect 934 2066 940 2067
rect 1046 2071 1052 2072
rect 1046 2067 1047 2071
rect 1051 2067 1052 2071
rect 1046 2066 1052 2067
rect 1120 2064 1122 2082
rect 1160 2072 1162 2089
rect 1258 2087 1264 2088
rect 1258 2083 1259 2087
rect 1263 2083 1264 2087
rect 1258 2082 1264 2083
rect 1158 2071 1164 2072
rect 1158 2067 1159 2071
rect 1163 2067 1164 2071
rect 1158 2066 1164 2067
rect 1260 2064 1262 2082
rect 1280 2072 1282 2089
rect 1768 2073 1770 2089
rect 1766 2072 1772 2073
rect 1788 2072 1790 2098
rect 1807 2097 1811 2098
rect 1831 2102 1835 2103
rect 1831 2097 1835 2098
rect 1991 2102 1995 2103
rect 1991 2097 1995 2098
rect 2167 2102 2171 2103
rect 2167 2097 2171 2098
rect 2343 2102 2347 2103
rect 2343 2097 2347 2098
rect 2503 2102 2507 2103
rect 2503 2097 2507 2098
rect 2655 2102 2659 2103
rect 2655 2097 2659 2098
rect 2791 2102 2795 2103
rect 2791 2097 2795 2098
rect 2919 2102 2923 2103
rect 2919 2097 2923 2098
rect 2927 2102 2931 2103
rect 2927 2097 2931 2098
rect 3015 2102 3019 2103
rect 3015 2097 3019 2098
rect 3039 2102 3043 2103
rect 3039 2097 3043 2098
rect 3103 2102 3107 2103
rect 3103 2097 3107 2098
rect 3159 2102 3163 2103
rect 3159 2097 3163 2098
rect 3191 2102 3195 2103
rect 3254 2099 3255 2103
rect 3259 2099 3260 2103
rect 3254 2098 3260 2099
rect 3271 2102 3275 2103
rect 3191 2097 3195 2098
rect 3271 2097 3275 2098
rect 3279 2102 3283 2103
rect 3279 2097 3283 2098
rect 1808 2081 1810 2097
rect 1806 2080 1812 2081
rect 1832 2080 1834 2097
rect 1938 2095 1944 2096
rect 1938 2091 1939 2095
rect 1943 2091 1944 2095
rect 1938 2090 1944 2091
rect 1806 2076 1807 2080
rect 1811 2076 1812 2080
rect 1806 2075 1812 2076
rect 1830 2079 1836 2080
rect 1830 2075 1831 2079
rect 1835 2075 1836 2079
rect 1830 2074 1836 2075
rect 1940 2072 1942 2090
rect 1992 2080 1994 2097
rect 2168 2080 2170 2097
rect 2344 2080 2346 2097
rect 2394 2095 2400 2096
rect 2394 2091 2395 2095
rect 2399 2091 2400 2095
rect 2394 2090 2400 2091
rect 1990 2079 1996 2080
rect 1990 2075 1991 2079
rect 1995 2075 1996 2079
rect 1990 2074 1996 2075
rect 2166 2079 2172 2080
rect 2166 2075 2167 2079
rect 2171 2075 2172 2079
rect 2166 2074 2172 2075
rect 2342 2079 2348 2080
rect 2342 2075 2343 2079
rect 2347 2075 2348 2079
rect 2342 2074 2348 2075
rect 1278 2071 1284 2072
rect 1278 2067 1279 2071
rect 1283 2067 1284 2071
rect 1766 2068 1767 2072
rect 1771 2068 1772 2072
rect 1766 2067 1772 2068
rect 1786 2071 1792 2072
rect 1786 2067 1787 2071
rect 1791 2067 1792 2071
rect 1278 2066 1284 2067
rect 1786 2066 1792 2067
rect 1938 2071 1944 2072
rect 1938 2067 1939 2071
rect 1943 2067 1944 2071
rect 1938 2066 1944 2067
rect 774 2063 780 2064
rect 774 2059 775 2063
rect 779 2059 780 2063
rect 774 2058 780 2059
rect 894 2063 900 2064
rect 894 2059 895 2063
rect 899 2059 900 2063
rect 894 2058 900 2059
rect 1118 2063 1124 2064
rect 1118 2059 1119 2063
rect 1123 2059 1124 2063
rect 1118 2058 1124 2059
rect 1258 2063 1264 2064
rect 1258 2059 1259 2063
rect 1263 2059 1264 2063
rect 1258 2058 1264 2059
rect 1270 2063 1276 2064
rect 1270 2059 1271 2063
rect 1275 2059 1276 2063
rect 1270 2058 1276 2059
rect 1806 2063 1812 2064
rect 1806 2059 1807 2063
rect 1811 2059 1812 2063
rect 1806 2058 1812 2059
rect 1830 2060 1836 2061
rect 822 2052 828 2053
rect 822 2048 823 2052
rect 827 2048 828 2052
rect 822 2047 828 2048
rect 934 2052 940 2053
rect 934 2048 935 2052
rect 939 2048 940 2052
rect 934 2047 940 2048
rect 1046 2052 1052 2053
rect 1046 2048 1047 2052
rect 1051 2048 1052 2052
rect 1046 2047 1052 2048
rect 1158 2052 1164 2053
rect 1158 2048 1159 2052
rect 1163 2048 1164 2052
rect 1158 2047 1164 2048
rect 824 2023 826 2047
rect 936 2023 938 2047
rect 1048 2023 1050 2047
rect 1160 2023 1162 2047
rect 775 2022 779 2023
rect 775 2017 779 2018
rect 823 2022 827 2023
rect 823 2017 827 2018
rect 911 2022 915 2023
rect 911 2017 915 2018
rect 935 2022 939 2023
rect 935 2017 939 2018
rect 1047 2022 1051 2023
rect 1047 2017 1051 2018
rect 1159 2022 1163 2023
rect 1159 2017 1163 2018
rect 1183 2022 1187 2023
rect 1183 2017 1187 2018
rect 776 2001 778 2017
rect 912 2001 914 2017
rect 1048 2001 1050 2017
rect 1184 2001 1186 2017
rect 774 2000 780 2001
rect 774 1996 775 2000
rect 779 1996 780 2000
rect 774 1995 780 1996
rect 910 2000 916 2001
rect 910 1996 911 2000
rect 915 1996 916 2000
rect 910 1995 916 1996
rect 1046 2000 1052 2001
rect 1046 1996 1047 2000
rect 1051 1996 1052 2000
rect 1046 1995 1052 1996
rect 1182 2000 1188 2001
rect 1182 1996 1183 2000
rect 1187 1996 1188 2000
rect 1182 1995 1188 1996
rect 206 1991 212 1992
rect 206 1987 207 1991
rect 211 1987 212 1991
rect 206 1986 212 1987
rect 310 1991 316 1992
rect 310 1987 311 1991
rect 315 1987 316 1991
rect 310 1986 316 1987
rect 438 1991 444 1992
rect 438 1987 439 1991
rect 443 1987 444 1991
rect 438 1986 444 1987
rect 574 1991 580 1992
rect 574 1987 575 1991
rect 579 1987 580 1991
rect 574 1986 580 1987
rect 582 1991 588 1992
rect 582 1987 583 1991
rect 587 1987 588 1991
rect 582 1986 588 1987
rect 754 1991 760 1992
rect 754 1987 755 1991
rect 759 1987 760 1991
rect 754 1986 760 1987
rect 854 1991 860 1992
rect 854 1987 855 1991
rect 859 1987 860 1991
rect 854 1986 860 1987
rect 1134 1991 1140 1992
rect 1134 1987 1135 1991
rect 1139 1987 1140 1991
rect 1134 1986 1140 1987
rect 1254 1991 1260 1992
rect 1254 1987 1255 1991
rect 1259 1987 1260 1991
rect 1254 1986 1260 1987
rect 208 1964 210 1986
rect 238 1981 244 1982
rect 238 1977 239 1981
rect 243 1977 244 1981
rect 238 1976 244 1977
rect 186 1963 192 1964
rect 186 1959 187 1963
rect 191 1959 192 1963
rect 186 1958 192 1959
rect 206 1963 212 1964
rect 206 1959 207 1963
rect 211 1959 212 1963
rect 206 1958 212 1959
rect 240 1955 242 1976
rect 312 1964 314 1986
rect 366 1981 372 1982
rect 366 1977 367 1981
rect 371 1977 372 1981
rect 366 1976 372 1977
rect 310 1963 316 1964
rect 310 1959 311 1963
rect 315 1959 316 1963
rect 310 1958 316 1959
rect 368 1955 370 1976
rect 440 1964 442 1986
rect 502 1981 508 1982
rect 502 1977 503 1981
rect 507 1977 508 1981
rect 502 1976 508 1977
rect 438 1963 444 1964
rect 438 1959 439 1963
rect 443 1959 444 1963
rect 438 1958 444 1959
rect 504 1955 506 1976
rect 576 1964 578 1986
rect 574 1963 580 1964
rect 574 1959 575 1963
rect 579 1959 580 1963
rect 574 1958 580 1959
rect 584 1956 586 1986
rect 638 1981 644 1982
rect 638 1977 639 1981
rect 643 1977 644 1981
rect 638 1976 644 1977
rect 774 1981 780 1982
rect 774 1977 775 1981
rect 779 1977 780 1981
rect 774 1976 780 1977
rect 582 1955 588 1956
rect 640 1955 642 1976
rect 776 1955 778 1976
rect 856 1964 858 1986
rect 910 1981 916 1982
rect 910 1977 911 1981
rect 915 1977 916 1981
rect 910 1976 916 1977
rect 1046 1981 1052 1982
rect 1046 1977 1047 1981
rect 1051 1977 1052 1981
rect 1046 1976 1052 1977
rect 854 1963 860 1964
rect 854 1959 855 1963
rect 859 1959 860 1963
rect 854 1958 860 1959
rect 912 1955 914 1976
rect 962 1963 968 1964
rect 962 1959 963 1963
rect 967 1959 968 1963
rect 962 1958 968 1959
rect 111 1954 115 1955
rect 111 1949 115 1950
rect 135 1954 139 1955
rect 135 1949 139 1950
rect 239 1954 243 1955
rect 239 1949 243 1950
rect 295 1954 299 1955
rect 295 1949 299 1950
rect 367 1954 371 1955
rect 367 1949 371 1950
rect 423 1954 427 1955
rect 423 1949 427 1950
rect 503 1954 507 1955
rect 503 1949 507 1950
rect 559 1954 563 1955
rect 582 1951 583 1955
rect 587 1951 588 1955
rect 582 1950 588 1951
rect 639 1954 643 1955
rect 559 1949 563 1950
rect 639 1949 643 1950
rect 703 1954 707 1955
rect 703 1949 707 1950
rect 775 1954 779 1955
rect 775 1949 779 1950
rect 855 1954 859 1955
rect 855 1949 859 1950
rect 911 1954 915 1955
rect 911 1949 915 1950
rect 112 1933 114 1949
rect 110 1932 116 1933
rect 296 1932 298 1949
rect 402 1947 408 1948
rect 402 1943 403 1947
rect 407 1943 408 1947
rect 402 1942 408 1943
rect 110 1928 111 1932
rect 115 1928 116 1932
rect 110 1927 116 1928
rect 294 1931 300 1932
rect 294 1927 295 1931
rect 299 1927 300 1931
rect 294 1926 300 1927
rect 404 1924 406 1942
rect 424 1932 426 1949
rect 494 1947 500 1948
rect 494 1943 495 1947
rect 499 1943 500 1947
rect 494 1942 500 1943
rect 422 1931 428 1932
rect 422 1927 423 1931
rect 427 1927 428 1931
rect 422 1926 428 1927
rect 496 1924 498 1942
rect 560 1932 562 1949
rect 630 1947 636 1948
rect 630 1943 631 1947
rect 635 1943 636 1947
rect 630 1942 636 1943
rect 558 1931 564 1932
rect 558 1927 559 1931
rect 563 1927 564 1931
rect 558 1926 564 1927
rect 632 1924 634 1942
rect 704 1932 706 1949
rect 856 1932 858 1949
rect 950 1947 956 1948
rect 950 1943 951 1947
rect 955 1943 956 1947
rect 950 1942 956 1943
rect 702 1931 708 1932
rect 702 1927 703 1931
rect 707 1927 708 1931
rect 702 1926 708 1927
rect 854 1931 860 1932
rect 854 1927 855 1931
rect 859 1927 860 1931
rect 854 1926 860 1927
rect 402 1923 408 1924
rect 402 1919 403 1923
rect 407 1919 408 1923
rect 402 1918 408 1919
rect 494 1923 500 1924
rect 494 1919 495 1923
rect 499 1919 500 1923
rect 494 1918 500 1919
rect 630 1923 636 1924
rect 630 1919 631 1923
rect 635 1919 636 1923
rect 630 1918 636 1919
rect 774 1919 780 1920
rect 110 1915 116 1916
rect 110 1911 111 1915
rect 115 1911 116 1915
rect 774 1915 775 1919
rect 779 1915 780 1919
rect 774 1914 780 1915
rect 110 1910 116 1911
rect 294 1912 300 1913
rect 112 1891 114 1910
rect 294 1908 295 1912
rect 299 1908 300 1912
rect 294 1907 300 1908
rect 422 1912 428 1913
rect 422 1908 423 1912
rect 427 1908 428 1912
rect 422 1907 428 1908
rect 558 1912 564 1913
rect 558 1908 559 1912
rect 563 1908 564 1912
rect 558 1907 564 1908
rect 702 1912 708 1913
rect 702 1908 703 1912
rect 707 1908 708 1912
rect 702 1907 708 1908
rect 296 1891 298 1907
rect 424 1891 426 1907
rect 560 1891 562 1907
rect 704 1891 706 1907
rect 111 1890 115 1891
rect 111 1885 115 1886
rect 295 1890 299 1891
rect 295 1885 299 1886
rect 423 1890 427 1891
rect 423 1885 427 1886
rect 431 1890 435 1891
rect 431 1885 435 1886
rect 559 1890 563 1891
rect 559 1885 563 1886
rect 575 1890 579 1891
rect 575 1885 579 1886
rect 703 1890 707 1891
rect 703 1885 707 1886
rect 727 1890 731 1891
rect 727 1885 731 1886
rect 112 1866 114 1885
rect 432 1869 434 1885
rect 576 1869 578 1885
rect 728 1869 730 1885
rect 430 1868 436 1869
rect 110 1865 116 1866
rect 110 1861 111 1865
rect 115 1861 116 1865
rect 430 1864 431 1868
rect 435 1864 436 1868
rect 430 1863 436 1864
rect 574 1868 580 1869
rect 574 1864 575 1868
rect 579 1864 580 1868
rect 574 1863 580 1864
rect 726 1868 732 1869
rect 726 1864 727 1868
rect 731 1864 732 1868
rect 726 1863 732 1864
rect 110 1860 116 1861
rect 502 1859 508 1860
rect 502 1855 503 1859
rect 507 1855 508 1859
rect 502 1854 508 1855
rect 510 1859 516 1860
rect 510 1855 511 1859
rect 515 1855 516 1859
rect 510 1854 516 1855
rect 654 1859 660 1860
rect 654 1855 655 1859
rect 659 1855 660 1859
rect 654 1854 660 1855
rect 430 1849 436 1850
rect 110 1848 116 1849
rect 110 1844 111 1848
rect 115 1844 116 1848
rect 430 1845 431 1849
rect 435 1845 436 1849
rect 430 1844 436 1845
rect 110 1843 116 1844
rect 112 1823 114 1843
rect 432 1823 434 1844
rect 111 1822 115 1823
rect 111 1817 115 1818
rect 431 1822 435 1823
rect 431 1817 435 1818
rect 112 1801 114 1817
rect 504 1816 506 1854
rect 512 1832 514 1854
rect 574 1849 580 1850
rect 574 1845 575 1849
rect 579 1845 580 1849
rect 574 1844 580 1845
rect 510 1831 516 1832
rect 510 1827 511 1831
rect 515 1827 516 1831
rect 510 1826 516 1827
rect 576 1823 578 1844
rect 656 1832 658 1854
rect 726 1849 732 1850
rect 726 1845 727 1849
rect 731 1845 732 1849
rect 726 1844 732 1845
rect 654 1831 660 1832
rect 654 1827 655 1831
rect 659 1827 660 1831
rect 654 1826 660 1827
rect 728 1823 730 1844
rect 776 1832 778 1914
rect 854 1912 860 1913
rect 854 1908 855 1912
rect 859 1908 860 1912
rect 854 1907 860 1908
rect 856 1891 858 1907
rect 855 1890 859 1891
rect 855 1885 859 1886
rect 887 1890 891 1891
rect 887 1885 891 1886
rect 888 1869 890 1885
rect 886 1868 892 1869
rect 886 1864 887 1868
rect 891 1864 892 1868
rect 886 1863 892 1864
rect 952 1860 954 1942
rect 964 1924 966 1958
rect 1048 1955 1050 1976
rect 1136 1964 1138 1986
rect 1182 1981 1188 1982
rect 1182 1977 1183 1981
rect 1187 1977 1188 1981
rect 1182 1976 1188 1977
rect 1134 1963 1140 1964
rect 1134 1959 1135 1963
rect 1139 1959 1140 1963
rect 1134 1958 1140 1959
rect 1184 1955 1186 1976
rect 1256 1964 1258 1986
rect 1254 1963 1260 1964
rect 1254 1959 1255 1963
rect 1259 1959 1260 1963
rect 1254 1958 1260 1959
rect 1272 1956 1274 2058
rect 1766 2055 1772 2056
rect 1278 2052 1284 2053
rect 1278 2048 1279 2052
rect 1283 2048 1284 2052
rect 1766 2051 1767 2055
rect 1771 2051 1772 2055
rect 1766 2050 1772 2051
rect 1278 2047 1284 2048
rect 1280 2023 1282 2047
rect 1768 2023 1770 2050
rect 1808 2035 1810 2058
rect 1830 2056 1831 2060
rect 1835 2056 1836 2060
rect 1830 2055 1836 2056
rect 1990 2060 1996 2061
rect 1990 2056 1991 2060
rect 1995 2056 1996 2060
rect 1990 2055 1996 2056
rect 2166 2060 2172 2061
rect 2166 2056 2167 2060
rect 2171 2056 2172 2060
rect 2166 2055 2172 2056
rect 2342 2060 2348 2061
rect 2342 2056 2343 2060
rect 2347 2056 2348 2060
rect 2342 2055 2348 2056
rect 1832 2035 1834 2055
rect 1992 2035 1994 2055
rect 2168 2035 2170 2055
rect 2344 2035 2346 2055
rect 1807 2034 1811 2035
rect 1807 2029 1811 2030
rect 1831 2034 1835 2035
rect 1831 2029 1835 2030
rect 1991 2034 1995 2035
rect 1991 2029 1995 2030
rect 2015 2034 2019 2035
rect 2015 2029 2019 2030
rect 2167 2034 2171 2035
rect 2167 2029 2171 2030
rect 2223 2034 2227 2035
rect 2223 2029 2227 2030
rect 2343 2034 2347 2035
rect 2343 2029 2347 2030
rect 1279 2022 1283 2023
rect 1279 2017 1283 2018
rect 1327 2022 1331 2023
rect 1327 2017 1331 2018
rect 1767 2022 1771 2023
rect 1767 2017 1771 2018
rect 1328 2001 1330 2017
rect 1326 2000 1332 2001
rect 1326 1996 1327 2000
rect 1331 1996 1332 2000
rect 1768 1998 1770 2017
rect 1808 2010 1810 2029
rect 1832 2013 1834 2029
rect 2016 2013 2018 2029
rect 2224 2013 2226 2029
rect 1830 2012 1836 2013
rect 1806 2009 1812 2010
rect 1806 2005 1807 2009
rect 1811 2005 1812 2009
rect 1830 2008 1831 2012
rect 1835 2008 1836 2012
rect 1830 2007 1836 2008
rect 2014 2012 2020 2013
rect 2014 2008 2015 2012
rect 2019 2008 2020 2012
rect 2014 2007 2020 2008
rect 2222 2012 2228 2013
rect 2222 2008 2223 2012
rect 2227 2008 2228 2012
rect 2222 2007 2228 2008
rect 1806 2004 1812 2005
rect 2396 2004 2398 2090
rect 2504 2080 2506 2097
rect 2582 2095 2588 2096
rect 2582 2091 2583 2095
rect 2587 2091 2588 2095
rect 2582 2090 2588 2091
rect 2502 2079 2508 2080
rect 2502 2075 2503 2079
rect 2507 2075 2508 2079
rect 2502 2074 2508 2075
rect 2584 2072 2586 2090
rect 2656 2080 2658 2097
rect 2734 2095 2740 2096
rect 2734 2091 2735 2095
rect 2739 2091 2740 2095
rect 2734 2090 2740 2091
rect 2654 2079 2660 2080
rect 2654 2075 2655 2079
rect 2659 2075 2660 2079
rect 2654 2074 2660 2075
rect 2736 2072 2738 2090
rect 2792 2080 2794 2097
rect 2920 2080 2922 2097
rect 3040 2080 3042 2097
rect 3086 2095 3092 2096
rect 3086 2091 3087 2095
rect 3091 2091 3092 2095
rect 3086 2090 3092 2091
rect 3110 2095 3116 2096
rect 3110 2091 3111 2095
rect 3115 2091 3116 2095
rect 3110 2090 3116 2091
rect 2790 2079 2796 2080
rect 2790 2075 2791 2079
rect 2795 2075 2796 2079
rect 2790 2074 2796 2075
rect 2918 2079 2924 2080
rect 2918 2075 2919 2079
rect 2923 2075 2924 2079
rect 2918 2074 2924 2075
rect 3038 2079 3044 2080
rect 3038 2075 3039 2079
rect 3043 2075 3044 2079
rect 3038 2074 3044 2075
rect 2582 2071 2588 2072
rect 2574 2067 2580 2068
rect 2574 2063 2575 2067
rect 2579 2063 2580 2067
rect 2582 2067 2583 2071
rect 2587 2067 2588 2071
rect 2582 2066 2588 2067
rect 2734 2071 2740 2072
rect 2734 2067 2735 2071
rect 2739 2067 2740 2071
rect 2734 2066 2740 2067
rect 2574 2062 2580 2063
rect 2502 2060 2508 2061
rect 2502 2056 2503 2060
rect 2507 2056 2508 2060
rect 2502 2055 2508 2056
rect 2504 2035 2506 2055
rect 2431 2034 2435 2035
rect 2431 2029 2435 2030
rect 2503 2034 2507 2035
rect 2503 2029 2507 2030
rect 2432 2013 2434 2029
rect 2430 2012 2436 2013
rect 2430 2008 2431 2012
rect 2435 2008 2436 2012
rect 2430 2007 2436 2008
rect 1966 2003 1972 2004
rect 1966 1999 1967 2003
rect 1971 1999 1972 2003
rect 1966 1998 1972 1999
rect 2086 2003 2092 2004
rect 2086 1999 2087 2003
rect 2091 1999 2092 2003
rect 2086 1998 2092 1999
rect 2294 2003 2300 2004
rect 2294 1999 2295 2003
rect 2299 1999 2300 2003
rect 2294 1998 2300 1999
rect 2394 2003 2400 2004
rect 2394 1999 2395 2003
rect 2399 1999 2400 2003
rect 2394 1998 2400 1999
rect 1326 1995 1332 1996
rect 1766 1997 1772 1998
rect 1766 1993 1767 1997
rect 1771 1993 1772 1997
rect 1830 1993 1836 1994
rect 1766 1992 1772 1993
rect 1806 1992 1812 1993
rect 1398 1991 1404 1992
rect 1398 1987 1399 1991
rect 1403 1987 1404 1991
rect 1806 1988 1807 1992
rect 1811 1988 1812 1992
rect 1830 1989 1831 1993
rect 1835 1989 1836 1993
rect 1830 1988 1836 1989
rect 1806 1987 1812 1988
rect 1398 1986 1404 1987
rect 1326 1981 1332 1982
rect 1326 1977 1327 1981
rect 1331 1977 1332 1981
rect 1326 1976 1332 1977
rect 1270 1955 1276 1956
rect 1328 1955 1330 1976
rect 1007 1954 1011 1955
rect 1007 1949 1011 1950
rect 1047 1954 1051 1955
rect 1047 1949 1051 1950
rect 1159 1954 1163 1955
rect 1159 1949 1163 1950
rect 1183 1954 1187 1955
rect 1270 1951 1271 1955
rect 1275 1951 1276 1955
rect 1270 1950 1276 1951
rect 1311 1954 1315 1955
rect 1183 1949 1187 1950
rect 1311 1949 1315 1950
rect 1327 1954 1331 1955
rect 1327 1949 1331 1950
rect 1008 1932 1010 1949
rect 1160 1932 1162 1949
rect 1238 1947 1244 1948
rect 1238 1943 1239 1947
rect 1243 1943 1244 1947
rect 1238 1942 1244 1943
rect 1006 1931 1012 1932
rect 1006 1927 1007 1931
rect 1011 1927 1012 1931
rect 1006 1926 1012 1927
rect 1158 1931 1164 1932
rect 1158 1927 1159 1931
rect 1163 1927 1164 1931
rect 1158 1926 1164 1927
rect 1240 1924 1242 1942
rect 1312 1932 1314 1949
rect 1400 1948 1402 1986
rect 1766 1980 1772 1981
rect 1766 1976 1767 1980
rect 1771 1976 1772 1980
rect 1766 1975 1772 1976
rect 1768 1955 1770 1975
rect 1808 1967 1810 1987
rect 1832 1967 1834 1988
rect 1968 1976 1970 1998
rect 2014 1993 2020 1994
rect 2014 1989 2015 1993
rect 2019 1989 2020 1993
rect 2014 1988 2020 1989
rect 1934 1975 1940 1976
rect 1934 1971 1935 1975
rect 1939 1971 1940 1975
rect 1934 1970 1940 1971
rect 1966 1975 1972 1976
rect 1966 1971 1967 1975
rect 1971 1971 1972 1975
rect 1966 1970 1972 1971
rect 1807 1966 1811 1967
rect 1807 1961 1811 1962
rect 1831 1966 1835 1967
rect 1831 1961 1835 1962
rect 1863 1966 1867 1967
rect 1863 1961 1867 1962
rect 1471 1954 1475 1955
rect 1471 1949 1475 1950
rect 1767 1954 1771 1955
rect 1767 1949 1771 1950
rect 1390 1947 1396 1948
rect 1390 1943 1391 1947
rect 1395 1943 1396 1947
rect 1390 1942 1396 1943
rect 1398 1947 1404 1948
rect 1398 1943 1399 1947
rect 1403 1943 1404 1947
rect 1398 1942 1404 1943
rect 1310 1931 1316 1932
rect 1310 1927 1311 1931
rect 1315 1927 1316 1931
rect 1310 1926 1316 1927
rect 1392 1924 1394 1942
rect 1472 1932 1474 1949
rect 1768 1933 1770 1949
rect 1808 1945 1810 1961
rect 1806 1944 1812 1945
rect 1864 1944 1866 1961
rect 1806 1940 1807 1944
rect 1811 1940 1812 1944
rect 1806 1939 1812 1940
rect 1862 1943 1868 1944
rect 1862 1939 1863 1943
rect 1867 1939 1868 1943
rect 1862 1938 1868 1939
rect 1936 1936 1938 1970
rect 2016 1967 2018 1988
rect 2088 1976 2090 1998
rect 2222 1993 2228 1994
rect 2222 1989 2223 1993
rect 2227 1989 2228 1993
rect 2222 1988 2228 1989
rect 2086 1975 2092 1976
rect 2086 1971 2087 1975
rect 2091 1971 2092 1975
rect 2086 1970 2092 1971
rect 2224 1967 2226 1988
rect 2296 1976 2298 1998
rect 2430 1993 2436 1994
rect 2430 1989 2431 1993
rect 2435 1989 2436 1993
rect 2430 1988 2436 1989
rect 2294 1975 2300 1976
rect 2294 1971 2295 1975
rect 2299 1971 2300 1975
rect 2294 1970 2300 1971
rect 2366 1967 2372 1968
rect 2432 1967 2434 1988
rect 2576 1976 2578 2062
rect 2654 2060 2660 2061
rect 2654 2056 2655 2060
rect 2659 2056 2660 2060
rect 2654 2055 2660 2056
rect 2790 2060 2796 2061
rect 2790 2056 2791 2060
rect 2795 2056 2796 2060
rect 2790 2055 2796 2056
rect 2918 2060 2924 2061
rect 2918 2056 2919 2060
rect 2923 2056 2924 2060
rect 2918 2055 2924 2056
rect 3038 2060 3044 2061
rect 3038 2056 3039 2060
rect 3043 2056 3044 2060
rect 3038 2055 3044 2056
rect 2656 2035 2658 2055
rect 2792 2035 2794 2055
rect 2920 2035 2922 2055
rect 3040 2035 3042 2055
rect 2631 2034 2635 2035
rect 2631 2029 2635 2030
rect 2655 2034 2659 2035
rect 2655 2029 2659 2030
rect 2791 2034 2795 2035
rect 2791 2029 2795 2030
rect 2823 2034 2827 2035
rect 2823 2029 2827 2030
rect 2919 2034 2923 2035
rect 2919 2029 2923 2030
rect 3007 2034 3011 2035
rect 3007 2029 3011 2030
rect 3039 2034 3043 2035
rect 3039 2029 3043 2030
rect 2632 2013 2634 2029
rect 2824 2013 2826 2029
rect 3008 2013 3010 2029
rect 2630 2012 2636 2013
rect 2630 2008 2631 2012
rect 2635 2008 2636 2012
rect 2630 2007 2636 2008
rect 2822 2012 2828 2013
rect 2822 2008 2823 2012
rect 2827 2008 2828 2012
rect 2822 2007 2828 2008
rect 3006 2012 3012 2013
rect 3006 2008 3007 2012
rect 3011 2008 3012 2012
rect 3006 2007 3012 2008
rect 3088 2004 3090 2090
rect 3112 2072 3114 2090
rect 3160 2080 3162 2097
rect 3230 2095 3236 2096
rect 3230 2091 3231 2095
rect 3235 2091 3236 2095
rect 3230 2090 3236 2091
rect 3158 2079 3164 2080
rect 3158 2075 3159 2079
rect 3163 2075 3164 2079
rect 3158 2074 3164 2075
rect 3232 2072 3234 2090
rect 3272 2080 3274 2097
rect 3352 2096 3354 2138
rect 3360 2116 3362 2138
rect 3366 2133 3372 2134
rect 3366 2129 3367 2133
rect 3371 2129 3372 2133
rect 3366 2128 3372 2129
rect 3358 2115 3364 2116
rect 3358 2111 3359 2115
rect 3363 2111 3364 2115
rect 3358 2110 3364 2111
rect 3368 2103 3370 2128
rect 3440 2116 3442 2198
rect 3462 2195 3463 2199
rect 3467 2195 3468 2199
rect 3462 2194 3468 2195
rect 3464 2175 3466 2194
rect 3463 2174 3467 2175
rect 3463 2169 3467 2170
rect 3464 2150 3466 2169
rect 3462 2149 3468 2150
rect 3462 2145 3463 2149
rect 3467 2145 3468 2149
rect 3462 2144 3468 2145
rect 3462 2132 3468 2133
rect 3462 2128 3463 2132
rect 3467 2128 3468 2132
rect 3462 2127 3468 2128
rect 3438 2115 3444 2116
rect 3438 2111 3439 2115
rect 3443 2111 3444 2115
rect 3438 2110 3444 2111
rect 3464 2103 3466 2127
rect 3367 2102 3371 2103
rect 3367 2097 3371 2098
rect 3463 2102 3467 2103
rect 3463 2097 3467 2098
rect 3350 2095 3356 2096
rect 3350 2091 3351 2095
rect 3355 2091 3356 2095
rect 3350 2090 3356 2091
rect 3368 2080 3370 2097
rect 3464 2081 3466 2097
rect 3462 2080 3468 2081
rect 3270 2079 3276 2080
rect 3270 2075 3271 2079
rect 3275 2075 3276 2079
rect 3270 2074 3276 2075
rect 3366 2079 3372 2080
rect 3366 2075 3367 2079
rect 3371 2075 3372 2079
rect 3462 2076 3463 2080
rect 3467 2076 3468 2080
rect 3462 2075 3468 2076
rect 3366 2074 3372 2075
rect 3110 2071 3116 2072
rect 3110 2067 3111 2071
rect 3115 2067 3116 2071
rect 3110 2066 3116 2067
rect 3230 2071 3236 2072
rect 3230 2067 3231 2071
rect 3235 2067 3236 2071
rect 3230 2066 3236 2067
rect 3438 2067 3444 2068
rect 3438 2063 3439 2067
rect 3443 2063 3444 2067
rect 3438 2062 3444 2063
rect 3462 2063 3468 2064
rect 3158 2060 3164 2061
rect 3158 2056 3159 2060
rect 3163 2056 3164 2060
rect 3158 2055 3164 2056
rect 3270 2060 3276 2061
rect 3270 2056 3271 2060
rect 3275 2056 3276 2060
rect 3270 2055 3276 2056
rect 3366 2060 3372 2061
rect 3366 2056 3367 2060
rect 3371 2056 3372 2060
rect 3366 2055 3372 2056
rect 3160 2035 3162 2055
rect 3272 2035 3274 2055
rect 3368 2035 3370 2055
rect 3159 2034 3163 2035
rect 3159 2029 3163 2030
rect 3199 2034 3203 2035
rect 3199 2029 3203 2030
rect 3271 2034 3275 2035
rect 3271 2029 3275 2030
rect 3367 2034 3371 2035
rect 3367 2029 3371 2030
rect 3200 2013 3202 2029
rect 3368 2013 3370 2029
rect 3198 2012 3204 2013
rect 3198 2008 3199 2012
rect 3203 2008 3204 2012
rect 3198 2007 3204 2008
rect 3366 2012 3372 2013
rect 3366 2008 3367 2012
rect 3371 2008 3372 2012
rect 3366 2007 3372 2008
rect 2702 2003 2708 2004
rect 2702 1999 2703 2003
rect 2707 1999 2708 2003
rect 2702 1998 2708 1999
rect 2894 2003 2900 2004
rect 2894 1999 2895 2003
rect 2899 1999 2900 2003
rect 2894 1998 2900 1999
rect 2998 2003 3004 2004
rect 2998 1999 2999 2003
rect 3003 1999 3004 2003
rect 2998 1998 3004 1999
rect 3086 2003 3092 2004
rect 3086 1999 3087 2003
rect 3091 1999 3092 2003
rect 3086 1998 3092 1999
rect 3430 2003 3436 2004
rect 3430 1999 3431 2003
rect 3435 1999 3436 2003
rect 3430 1998 3436 1999
rect 2630 1993 2636 1994
rect 2630 1989 2631 1993
rect 2635 1989 2636 1993
rect 2630 1988 2636 1989
rect 2574 1975 2580 1976
rect 2574 1971 2575 1975
rect 2579 1971 2580 1975
rect 2574 1970 2580 1971
rect 2632 1967 2634 1988
rect 2704 1976 2706 1998
rect 2822 1993 2828 1994
rect 2822 1989 2823 1993
rect 2827 1989 2828 1993
rect 2822 1988 2828 1989
rect 2702 1975 2708 1976
rect 2702 1971 2703 1975
rect 2707 1971 2708 1975
rect 2702 1970 2708 1971
rect 2824 1967 2826 1988
rect 2896 1976 2898 1998
rect 2894 1975 2900 1976
rect 2894 1971 2895 1975
rect 2899 1971 2900 1975
rect 2894 1970 2900 1971
rect 1999 1966 2003 1967
rect 1999 1961 2003 1962
rect 2015 1966 2019 1967
rect 2015 1961 2019 1962
rect 2143 1966 2147 1967
rect 2143 1961 2147 1962
rect 2223 1966 2227 1967
rect 2223 1961 2227 1962
rect 2287 1966 2291 1967
rect 2366 1963 2367 1967
rect 2371 1963 2372 1967
rect 2366 1962 2372 1963
rect 2431 1966 2435 1967
rect 2287 1961 2291 1962
rect 2000 1944 2002 1961
rect 2078 1959 2084 1960
rect 2078 1955 2079 1959
rect 2083 1955 2084 1959
rect 2078 1954 2084 1955
rect 1998 1943 2004 1944
rect 1998 1939 1999 1943
rect 2003 1939 2004 1943
rect 1998 1938 2004 1939
rect 2080 1936 2082 1954
rect 2144 1944 2146 1961
rect 2288 1944 2290 1961
rect 2298 1959 2304 1960
rect 2298 1955 2299 1959
rect 2303 1955 2304 1959
rect 2298 1954 2304 1955
rect 2358 1959 2364 1960
rect 2358 1955 2359 1959
rect 2363 1955 2364 1959
rect 2358 1954 2364 1955
rect 2142 1943 2148 1944
rect 2142 1939 2143 1943
rect 2147 1939 2148 1943
rect 2142 1938 2148 1939
rect 2286 1943 2292 1944
rect 2286 1939 2287 1943
rect 2291 1939 2292 1943
rect 2286 1938 2292 1939
rect 1934 1935 1940 1936
rect 1766 1932 1772 1933
rect 1470 1931 1476 1932
rect 1470 1927 1471 1931
rect 1475 1927 1476 1931
rect 1766 1928 1767 1932
rect 1771 1928 1772 1932
rect 1934 1931 1935 1935
rect 1939 1931 1940 1935
rect 1934 1930 1940 1931
rect 2078 1935 2084 1936
rect 2078 1931 2079 1935
rect 2083 1931 2084 1935
rect 2078 1930 2084 1931
rect 1766 1927 1772 1928
rect 1806 1927 1812 1928
rect 1470 1926 1476 1927
rect 962 1923 968 1924
rect 962 1919 963 1923
rect 967 1919 968 1923
rect 1238 1923 1244 1924
rect 962 1918 968 1919
rect 1230 1919 1236 1920
rect 1230 1915 1231 1919
rect 1235 1915 1236 1919
rect 1238 1919 1239 1923
rect 1243 1919 1244 1923
rect 1238 1918 1244 1919
rect 1390 1923 1396 1924
rect 1390 1919 1391 1923
rect 1395 1919 1396 1923
rect 1806 1923 1807 1927
rect 1811 1923 1812 1927
rect 1806 1922 1812 1923
rect 1862 1924 1868 1925
rect 1390 1918 1396 1919
rect 1230 1914 1236 1915
rect 1766 1915 1772 1916
rect 1006 1912 1012 1913
rect 1006 1908 1007 1912
rect 1011 1908 1012 1912
rect 1006 1907 1012 1908
rect 1158 1912 1164 1913
rect 1158 1908 1159 1912
rect 1163 1908 1164 1912
rect 1158 1907 1164 1908
rect 1008 1891 1010 1907
rect 1160 1891 1162 1907
rect 1007 1890 1011 1891
rect 1007 1885 1011 1886
rect 1047 1890 1051 1891
rect 1047 1885 1051 1886
rect 1159 1890 1163 1891
rect 1159 1885 1163 1886
rect 1199 1890 1203 1891
rect 1199 1885 1203 1886
rect 1048 1869 1050 1885
rect 1200 1869 1202 1885
rect 1046 1868 1052 1869
rect 1046 1864 1047 1868
rect 1051 1864 1052 1868
rect 1046 1863 1052 1864
rect 1198 1868 1204 1869
rect 1198 1864 1199 1868
rect 1203 1864 1204 1868
rect 1198 1863 1204 1864
rect 950 1859 956 1860
rect 950 1855 951 1859
rect 955 1855 956 1859
rect 950 1854 956 1855
rect 966 1859 972 1860
rect 966 1855 967 1859
rect 971 1855 972 1859
rect 966 1854 972 1855
rect 886 1849 892 1850
rect 886 1845 887 1849
rect 891 1845 892 1849
rect 886 1844 892 1845
rect 774 1831 780 1832
rect 774 1827 775 1831
rect 779 1827 780 1831
rect 774 1826 780 1827
rect 888 1823 890 1844
rect 968 1832 970 1854
rect 1046 1849 1052 1850
rect 1046 1845 1047 1849
rect 1051 1845 1052 1849
rect 1046 1844 1052 1845
rect 1198 1849 1204 1850
rect 1198 1845 1199 1849
rect 1203 1845 1204 1849
rect 1198 1844 1204 1845
rect 966 1831 972 1832
rect 966 1827 967 1831
rect 971 1827 972 1831
rect 966 1826 972 1827
rect 1048 1823 1050 1844
rect 1094 1831 1100 1832
rect 1094 1827 1095 1831
rect 1099 1827 1100 1831
rect 1094 1826 1100 1827
rect 511 1822 515 1823
rect 511 1817 515 1818
rect 575 1822 579 1823
rect 575 1817 579 1818
rect 631 1822 635 1823
rect 631 1817 635 1818
rect 727 1822 731 1823
rect 727 1817 731 1818
rect 759 1822 763 1823
rect 759 1817 763 1818
rect 887 1822 891 1823
rect 887 1817 891 1818
rect 1023 1822 1027 1823
rect 1023 1817 1027 1818
rect 1047 1822 1051 1823
rect 1047 1817 1051 1818
rect 502 1815 508 1816
rect 502 1811 503 1815
rect 507 1811 508 1815
rect 502 1810 508 1811
rect 110 1800 116 1801
rect 512 1800 514 1817
rect 582 1815 588 1816
rect 582 1811 583 1815
rect 587 1811 588 1815
rect 582 1810 588 1811
rect 110 1796 111 1800
rect 115 1796 116 1800
rect 110 1795 116 1796
rect 510 1799 516 1800
rect 510 1795 511 1799
rect 515 1795 516 1799
rect 510 1794 516 1795
rect 584 1792 586 1810
rect 632 1800 634 1817
rect 760 1800 762 1817
rect 822 1815 828 1816
rect 822 1811 823 1815
rect 827 1811 828 1815
rect 822 1810 828 1811
rect 830 1815 836 1816
rect 830 1811 831 1815
rect 835 1811 836 1815
rect 830 1810 836 1811
rect 630 1799 636 1800
rect 630 1795 631 1799
rect 635 1795 636 1799
rect 630 1794 636 1795
rect 758 1799 764 1800
rect 758 1795 759 1799
rect 763 1795 764 1799
rect 758 1794 764 1795
rect 582 1791 588 1792
rect 582 1787 583 1791
rect 587 1787 588 1791
rect 582 1786 588 1787
rect 702 1787 708 1788
rect 110 1783 116 1784
rect 110 1779 111 1783
rect 115 1779 116 1783
rect 702 1783 703 1787
rect 707 1783 708 1787
rect 702 1782 708 1783
rect 110 1778 116 1779
rect 510 1780 516 1781
rect 112 1755 114 1778
rect 510 1776 511 1780
rect 515 1776 516 1780
rect 510 1775 516 1776
rect 630 1780 636 1781
rect 630 1776 631 1780
rect 635 1776 636 1780
rect 630 1775 636 1776
rect 512 1755 514 1775
rect 632 1755 634 1775
rect 111 1754 115 1755
rect 111 1749 115 1750
rect 439 1754 443 1755
rect 439 1749 443 1750
rect 511 1754 515 1755
rect 511 1749 515 1750
rect 535 1754 539 1755
rect 535 1749 539 1750
rect 631 1754 635 1755
rect 631 1749 635 1750
rect 639 1754 643 1755
rect 639 1749 643 1750
rect 112 1730 114 1749
rect 440 1733 442 1749
rect 536 1733 538 1749
rect 640 1733 642 1749
rect 438 1732 444 1733
rect 110 1729 116 1730
rect 110 1725 111 1729
rect 115 1725 116 1729
rect 438 1728 439 1732
rect 443 1728 444 1732
rect 438 1727 444 1728
rect 534 1732 540 1733
rect 534 1728 535 1732
rect 539 1728 540 1732
rect 534 1727 540 1728
rect 638 1732 644 1733
rect 638 1728 639 1732
rect 643 1728 644 1732
rect 638 1727 644 1728
rect 110 1724 116 1725
rect 502 1723 508 1724
rect 502 1719 503 1723
rect 507 1719 508 1723
rect 502 1718 508 1719
rect 518 1723 524 1724
rect 518 1719 519 1723
rect 523 1719 524 1723
rect 518 1718 524 1719
rect 614 1723 620 1724
rect 614 1719 615 1723
rect 619 1719 620 1723
rect 614 1718 620 1719
rect 438 1713 444 1714
rect 110 1712 116 1713
rect 110 1708 111 1712
rect 115 1708 116 1712
rect 438 1709 439 1713
rect 443 1709 444 1713
rect 438 1708 444 1709
rect 110 1707 116 1708
rect 112 1687 114 1707
rect 440 1687 442 1708
rect 111 1686 115 1687
rect 111 1681 115 1682
rect 399 1686 403 1687
rect 399 1681 403 1682
rect 439 1686 443 1687
rect 439 1681 443 1682
rect 487 1686 491 1687
rect 487 1681 491 1682
rect 112 1665 114 1681
rect 110 1664 116 1665
rect 400 1664 402 1681
rect 488 1664 490 1681
rect 504 1680 506 1718
rect 520 1696 522 1718
rect 534 1713 540 1714
rect 534 1709 535 1713
rect 539 1709 540 1713
rect 534 1708 540 1709
rect 518 1695 524 1696
rect 518 1691 519 1695
rect 523 1691 524 1695
rect 518 1690 524 1691
rect 536 1687 538 1708
rect 616 1696 618 1718
rect 638 1713 644 1714
rect 638 1709 639 1713
rect 643 1709 644 1713
rect 638 1708 644 1709
rect 614 1695 620 1696
rect 614 1691 615 1695
rect 619 1691 620 1695
rect 614 1690 620 1691
rect 640 1687 642 1708
rect 704 1696 706 1782
rect 758 1780 764 1781
rect 758 1776 759 1780
rect 763 1776 764 1780
rect 758 1775 764 1776
rect 760 1755 762 1775
rect 743 1754 747 1755
rect 743 1749 747 1750
rect 759 1754 763 1755
rect 759 1749 763 1750
rect 744 1733 746 1749
rect 742 1732 748 1733
rect 742 1728 743 1732
rect 747 1728 748 1732
rect 742 1727 748 1728
rect 824 1724 826 1810
rect 832 1792 834 1810
rect 888 1800 890 1817
rect 958 1815 964 1816
rect 958 1811 959 1815
rect 963 1811 964 1815
rect 958 1810 964 1811
rect 886 1799 892 1800
rect 886 1795 887 1799
rect 891 1795 892 1799
rect 886 1794 892 1795
rect 960 1792 962 1810
rect 1024 1800 1026 1817
rect 1022 1799 1028 1800
rect 1022 1795 1023 1799
rect 1027 1795 1028 1799
rect 1022 1794 1028 1795
rect 1096 1792 1098 1826
rect 1200 1823 1202 1844
rect 1232 1832 1234 1914
rect 1310 1912 1316 1913
rect 1310 1908 1311 1912
rect 1315 1908 1316 1912
rect 1310 1907 1316 1908
rect 1470 1912 1476 1913
rect 1470 1908 1471 1912
rect 1475 1908 1476 1912
rect 1766 1911 1767 1915
rect 1771 1911 1772 1915
rect 1766 1910 1772 1911
rect 1470 1907 1476 1908
rect 1312 1891 1314 1907
rect 1472 1891 1474 1907
rect 1768 1891 1770 1910
rect 1808 1899 1810 1922
rect 1862 1920 1863 1924
rect 1867 1920 1868 1924
rect 1862 1919 1868 1920
rect 1998 1924 2004 1925
rect 1998 1920 1999 1924
rect 2003 1920 2004 1924
rect 1998 1919 2004 1920
rect 2142 1924 2148 1925
rect 2142 1920 2143 1924
rect 2147 1920 2148 1924
rect 2142 1919 2148 1920
rect 2286 1924 2292 1925
rect 2286 1920 2287 1924
rect 2291 1920 2292 1924
rect 2286 1919 2292 1920
rect 1864 1899 1866 1919
rect 2000 1899 2002 1919
rect 2144 1899 2146 1919
rect 2288 1899 2290 1919
rect 1807 1898 1811 1899
rect 1807 1893 1811 1894
rect 1863 1898 1867 1899
rect 1863 1893 1867 1894
rect 1999 1898 2003 1899
rect 1999 1893 2003 1894
rect 2015 1898 2019 1899
rect 2015 1893 2019 1894
rect 2111 1898 2115 1899
rect 2111 1893 2115 1894
rect 2143 1898 2147 1899
rect 2143 1893 2147 1894
rect 2215 1898 2219 1899
rect 2215 1893 2219 1894
rect 2287 1898 2291 1899
rect 2287 1893 2291 1894
rect 1311 1890 1315 1891
rect 1311 1885 1315 1886
rect 1351 1890 1355 1891
rect 1351 1885 1355 1886
rect 1471 1890 1475 1891
rect 1471 1885 1475 1886
rect 1511 1890 1515 1891
rect 1511 1885 1515 1886
rect 1671 1890 1675 1891
rect 1671 1885 1675 1886
rect 1767 1890 1771 1891
rect 1767 1885 1771 1886
rect 1352 1869 1354 1885
rect 1512 1869 1514 1885
rect 1672 1869 1674 1885
rect 1350 1868 1356 1869
rect 1350 1864 1351 1868
rect 1355 1864 1356 1868
rect 1350 1863 1356 1864
rect 1510 1868 1516 1869
rect 1510 1864 1511 1868
rect 1515 1864 1516 1868
rect 1510 1863 1516 1864
rect 1670 1868 1676 1869
rect 1670 1864 1671 1868
rect 1675 1864 1676 1868
rect 1768 1866 1770 1885
rect 1808 1874 1810 1893
rect 2016 1877 2018 1893
rect 2112 1877 2114 1893
rect 2216 1877 2218 1893
rect 2014 1876 2020 1877
rect 1806 1873 1812 1874
rect 1806 1869 1807 1873
rect 1811 1869 1812 1873
rect 2014 1872 2015 1876
rect 2019 1872 2020 1876
rect 2014 1871 2020 1872
rect 2110 1876 2116 1877
rect 2110 1872 2111 1876
rect 2115 1872 2116 1876
rect 2110 1871 2116 1872
rect 2214 1876 2220 1877
rect 2214 1872 2215 1876
rect 2219 1872 2220 1876
rect 2214 1871 2220 1872
rect 1806 1868 1812 1869
rect 2300 1868 2302 1954
rect 2360 1936 2362 1954
rect 2368 1936 2370 1962
rect 2431 1961 2435 1962
rect 2575 1966 2579 1967
rect 2575 1961 2579 1962
rect 2631 1966 2635 1967
rect 2631 1961 2635 1962
rect 2711 1966 2715 1967
rect 2711 1961 2715 1962
rect 2823 1966 2827 1967
rect 2823 1961 2827 1962
rect 2831 1966 2835 1967
rect 2831 1961 2835 1962
rect 2951 1966 2955 1967
rect 2951 1961 2955 1962
rect 2432 1944 2434 1961
rect 2576 1944 2578 1961
rect 2654 1959 2660 1960
rect 2654 1955 2655 1959
rect 2659 1955 2660 1959
rect 2654 1954 2660 1955
rect 2430 1943 2436 1944
rect 2430 1939 2431 1943
rect 2435 1939 2436 1943
rect 2430 1938 2436 1939
rect 2574 1943 2580 1944
rect 2574 1939 2575 1943
rect 2579 1939 2580 1943
rect 2574 1938 2580 1939
rect 2656 1936 2658 1954
rect 2712 1944 2714 1961
rect 2798 1959 2804 1960
rect 2798 1955 2799 1959
rect 2803 1955 2804 1959
rect 2798 1954 2804 1955
rect 2710 1943 2716 1944
rect 2710 1939 2711 1943
rect 2715 1939 2716 1943
rect 2710 1938 2716 1939
rect 2800 1936 2802 1954
rect 2832 1944 2834 1961
rect 2910 1959 2916 1960
rect 2910 1955 2911 1959
rect 2915 1955 2916 1959
rect 2910 1954 2916 1955
rect 2830 1943 2836 1944
rect 2830 1939 2831 1943
rect 2835 1939 2836 1943
rect 2830 1938 2836 1939
rect 2912 1936 2914 1954
rect 2952 1944 2954 1961
rect 3000 1960 3002 1998
rect 3006 1993 3012 1994
rect 3006 1989 3007 1993
rect 3011 1989 3012 1993
rect 3006 1988 3012 1989
rect 3198 1993 3204 1994
rect 3198 1989 3199 1993
rect 3203 1989 3204 1993
rect 3198 1988 3204 1989
rect 3366 1993 3372 1994
rect 3366 1989 3367 1993
rect 3371 1989 3372 1993
rect 3366 1988 3372 1989
rect 3008 1967 3010 1988
rect 3200 1967 3202 1988
rect 3238 1975 3244 1976
rect 3238 1971 3239 1975
rect 3243 1971 3244 1975
rect 3238 1970 3244 1971
rect 3007 1966 3011 1967
rect 3007 1961 3011 1962
rect 3063 1966 3067 1967
rect 3063 1961 3067 1962
rect 3167 1966 3171 1967
rect 3167 1961 3171 1962
rect 3199 1966 3203 1967
rect 3199 1961 3203 1962
rect 2998 1959 3004 1960
rect 2998 1955 2999 1959
rect 3003 1955 3004 1959
rect 2998 1954 3004 1955
rect 3064 1944 3066 1961
rect 3134 1959 3140 1960
rect 3134 1955 3135 1959
rect 3139 1955 3140 1959
rect 3134 1954 3140 1955
rect 2950 1943 2956 1944
rect 2950 1939 2951 1943
rect 2955 1939 2956 1943
rect 2950 1938 2956 1939
rect 3062 1943 3068 1944
rect 3062 1939 3063 1943
rect 3067 1939 3068 1943
rect 3062 1938 3068 1939
rect 3136 1936 3138 1954
rect 3168 1944 3170 1961
rect 3166 1943 3172 1944
rect 3166 1939 3167 1943
rect 3171 1939 3172 1943
rect 3166 1938 3172 1939
rect 3240 1936 3242 1970
rect 3246 1967 3252 1968
rect 3368 1967 3370 1988
rect 3246 1963 3247 1967
rect 3251 1963 3252 1967
rect 3246 1962 3252 1963
rect 3279 1966 3283 1967
rect 3248 1936 3250 1962
rect 3279 1961 3283 1962
rect 3367 1966 3371 1967
rect 3367 1961 3371 1962
rect 3280 1944 3282 1961
rect 3358 1959 3364 1960
rect 3358 1955 3359 1959
rect 3363 1955 3364 1959
rect 3358 1954 3364 1955
rect 3278 1943 3284 1944
rect 3278 1939 3279 1943
rect 3283 1939 3284 1943
rect 3278 1938 3284 1939
rect 3360 1936 3362 1954
rect 3368 1944 3370 1961
rect 3432 1960 3434 1998
rect 3440 1976 3442 2062
rect 3462 2059 3463 2063
rect 3467 2059 3468 2063
rect 3462 2058 3468 2059
rect 3464 2035 3466 2058
rect 3463 2034 3467 2035
rect 3463 2029 3467 2030
rect 3464 2010 3466 2029
rect 3462 2009 3468 2010
rect 3462 2005 3463 2009
rect 3467 2005 3468 2009
rect 3462 2004 3468 2005
rect 3462 1992 3468 1993
rect 3462 1988 3463 1992
rect 3467 1988 3468 1992
rect 3462 1987 3468 1988
rect 3438 1975 3444 1976
rect 3438 1971 3439 1975
rect 3443 1971 3444 1975
rect 3438 1970 3444 1971
rect 3464 1967 3466 1987
rect 3463 1966 3467 1967
rect 3463 1961 3467 1962
rect 3430 1959 3436 1960
rect 3430 1955 3431 1959
rect 3435 1955 3436 1959
rect 3430 1954 3436 1955
rect 3464 1945 3466 1961
rect 3462 1944 3468 1945
rect 3366 1943 3372 1944
rect 3366 1939 3367 1943
rect 3371 1939 3372 1943
rect 3462 1940 3463 1944
rect 3467 1940 3468 1944
rect 3462 1939 3468 1940
rect 3366 1938 3372 1939
rect 2358 1935 2364 1936
rect 2358 1931 2359 1935
rect 2363 1931 2364 1935
rect 2358 1930 2364 1931
rect 2366 1935 2372 1936
rect 2366 1931 2367 1935
rect 2371 1931 2372 1935
rect 2366 1930 2372 1931
rect 2654 1935 2660 1936
rect 2654 1931 2655 1935
rect 2659 1931 2660 1935
rect 2654 1930 2660 1931
rect 2798 1935 2804 1936
rect 2798 1931 2799 1935
rect 2803 1931 2804 1935
rect 2798 1930 2804 1931
rect 2910 1935 2916 1936
rect 2910 1931 2911 1935
rect 2915 1931 2916 1935
rect 2910 1930 2916 1931
rect 3134 1935 3140 1936
rect 3134 1931 3135 1935
rect 3139 1931 3140 1935
rect 3134 1930 3140 1931
rect 3238 1935 3244 1936
rect 3238 1931 3239 1935
rect 3243 1931 3244 1935
rect 3238 1930 3244 1931
rect 3246 1935 3252 1936
rect 3246 1931 3247 1935
rect 3251 1931 3252 1935
rect 3246 1930 3252 1931
rect 3358 1935 3364 1936
rect 3358 1931 3359 1935
rect 3363 1931 3364 1935
rect 3358 1930 3364 1931
rect 2638 1927 2644 1928
rect 2430 1924 2436 1925
rect 2430 1920 2431 1924
rect 2435 1920 2436 1924
rect 2430 1919 2436 1920
rect 2574 1924 2580 1925
rect 2574 1920 2575 1924
rect 2579 1920 2580 1924
rect 2638 1923 2639 1927
rect 2643 1923 2644 1927
rect 3462 1927 3468 1928
rect 2638 1922 2644 1923
rect 2710 1924 2716 1925
rect 2574 1919 2580 1920
rect 2432 1899 2434 1919
rect 2576 1899 2578 1919
rect 2327 1898 2331 1899
rect 2327 1893 2331 1894
rect 2431 1898 2435 1899
rect 2431 1893 2435 1894
rect 2439 1898 2443 1899
rect 2439 1893 2443 1894
rect 2543 1898 2547 1899
rect 2543 1893 2547 1894
rect 2575 1898 2579 1899
rect 2575 1893 2579 1894
rect 2328 1877 2330 1893
rect 2440 1877 2442 1893
rect 2544 1877 2546 1893
rect 2326 1876 2332 1877
rect 2326 1872 2327 1876
rect 2331 1872 2332 1876
rect 2326 1871 2332 1872
rect 2438 1876 2444 1877
rect 2438 1872 2439 1876
rect 2443 1872 2444 1876
rect 2438 1871 2444 1872
rect 2542 1876 2548 1877
rect 2542 1872 2543 1876
rect 2547 1872 2548 1876
rect 2542 1871 2548 1872
rect 2086 1867 2092 1868
rect 1670 1863 1676 1864
rect 1766 1865 1772 1866
rect 1766 1861 1767 1865
rect 1771 1861 1772 1865
rect 2086 1863 2087 1867
rect 2091 1863 2092 1867
rect 2086 1862 2092 1863
rect 2182 1867 2188 1868
rect 2182 1863 2183 1867
rect 2187 1863 2188 1867
rect 2182 1862 2188 1863
rect 2298 1867 2304 1868
rect 2298 1863 2299 1867
rect 2303 1863 2304 1867
rect 2298 1862 2304 1863
rect 2306 1867 2312 1868
rect 2306 1863 2307 1867
rect 2311 1863 2312 1867
rect 2306 1862 2312 1863
rect 2406 1867 2412 1868
rect 2406 1863 2407 1867
rect 2411 1863 2412 1867
rect 2406 1862 2412 1863
rect 1766 1860 1772 1861
rect 1270 1859 1276 1860
rect 1270 1855 1271 1859
rect 1275 1855 1276 1859
rect 1270 1854 1276 1855
rect 1422 1859 1428 1860
rect 1422 1855 1423 1859
rect 1427 1855 1428 1859
rect 1422 1854 1428 1855
rect 1582 1859 1588 1860
rect 1582 1855 1583 1859
rect 1587 1855 1588 1859
rect 1582 1854 1588 1855
rect 1734 1859 1740 1860
rect 1734 1855 1735 1859
rect 1739 1855 1740 1859
rect 2014 1857 2020 1858
rect 1734 1854 1740 1855
rect 1806 1856 1812 1857
rect 1272 1832 1274 1854
rect 1350 1849 1356 1850
rect 1350 1845 1351 1849
rect 1355 1845 1356 1849
rect 1350 1844 1356 1845
rect 1230 1831 1236 1832
rect 1230 1827 1231 1831
rect 1235 1827 1236 1831
rect 1230 1826 1236 1827
rect 1270 1831 1276 1832
rect 1270 1827 1271 1831
rect 1275 1827 1276 1831
rect 1270 1826 1276 1827
rect 1352 1823 1354 1844
rect 1424 1832 1426 1854
rect 1510 1849 1516 1850
rect 1510 1845 1511 1849
rect 1515 1845 1516 1849
rect 1510 1844 1516 1845
rect 1422 1831 1428 1832
rect 1422 1827 1423 1831
rect 1427 1827 1428 1831
rect 1422 1826 1428 1827
rect 1358 1823 1364 1824
rect 1512 1823 1514 1844
rect 1584 1832 1586 1854
rect 1670 1849 1676 1850
rect 1670 1845 1671 1849
rect 1675 1845 1676 1849
rect 1670 1844 1676 1845
rect 1582 1831 1588 1832
rect 1582 1827 1583 1831
rect 1587 1827 1588 1831
rect 1582 1826 1588 1827
rect 1672 1823 1674 1844
rect 1151 1822 1155 1823
rect 1151 1817 1155 1818
rect 1199 1822 1203 1823
rect 1199 1817 1203 1818
rect 1279 1822 1283 1823
rect 1279 1817 1283 1818
rect 1351 1822 1355 1823
rect 1358 1819 1359 1823
rect 1363 1819 1364 1823
rect 1358 1818 1364 1819
rect 1407 1822 1411 1823
rect 1351 1817 1355 1818
rect 1152 1800 1154 1817
rect 1222 1815 1228 1816
rect 1222 1811 1223 1815
rect 1227 1811 1228 1815
rect 1222 1810 1228 1811
rect 1150 1799 1156 1800
rect 1150 1795 1151 1799
rect 1155 1795 1156 1799
rect 1150 1794 1156 1795
rect 1224 1792 1226 1810
rect 1280 1800 1282 1817
rect 1278 1799 1284 1800
rect 1278 1795 1279 1799
rect 1283 1795 1284 1799
rect 1278 1794 1284 1795
rect 1360 1792 1362 1818
rect 1407 1817 1411 1818
rect 1511 1822 1515 1823
rect 1511 1817 1515 1818
rect 1535 1822 1539 1823
rect 1535 1817 1539 1818
rect 1671 1822 1675 1823
rect 1671 1817 1675 1818
rect 1408 1800 1410 1817
rect 1486 1815 1492 1816
rect 1486 1811 1487 1815
rect 1491 1811 1492 1815
rect 1486 1810 1492 1811
rect 1406 1799 1412 1800
rect 1406 1795 1407 1799
rect 1411 1795 1412 1799
rect 1406 1794 1412 1795
rect 1488 1792 1490 1810
rect 1536 1800 1538 1817
rect 1614 1815 1620 1816
rect 1614 1811 1615 1815
rect 1619 1811 1620 1815
rect 1614 1810 1620 1811
rect 1534 1799 1540 1800
rect 1534 1795 1535 1799
rect 1539 1795 1540 1799
rect 1534 1794 1540 1795
rect 1616 1792 1618 1810
rect 1672 1800 1674 1817
rect 1736 1816 1738 1854
rect 1806 1852 1807 1856
rect 1811 1852 1812 1856
rect 2014 1853 2015 1857
rect 2019 1853 2020 1857
rect 2014 1852 2020 1853
rect 1806 1851 1812 1852
rect 1766 1848 1772 1849
rect 1766 1844 1767 1848
rect 1771 1844 1772 1848
rect 1766 1843 1772 1844
rect 1768 1823 1770 1843
rect 1808 1827 1810 1851
rect 2016 1827 2018 1852
rect 2088 1840 2090 1862
rect 2110 1857 2116 1858
rect 2110 1853 2111 1857
rect 2115 1853 2116 1857
rect 2110 1852 2116 1853
rect 2086 1839 2092 1840
rect 2086 1835 2087 1839
rect 2091 1835 2092 1839
rect 2086 1834 2092 1835
rect 2112 1827 2114 1852
rect 2184 1840 2186 1862
rect 2214 1857 2220 1858
rect 2214 1853 2215 1857
rect 2219 1853 2220 1857
rect 2214 1852 2220 1853
rect 2182 1839 2188 1840
rect 2182 1835 2183 1839
rect 2187 1835 2188 1839
rect 2182 1834 2188 1835
rect 2216 1827 2218 1852
rect 2308 1832 2310 1862
rect 2326 1857 2332 1858
rect 2326 1853 2327 1857
rect 2331 1853 2332 1857
rect 2326 1852 2332 1853
rect 2306 1831 2312 1832
rect 2306 1827 2307 1831
rect 2311 1827 2312 1831
rect 2328 1827 2330 1852
rect 2408 1840 2410 1862
rect 2438 1857 2444 1858
rect 2438 1853 2439 1857
rect 2443 1853 2444 1857
rect 2438 1852 2444 1853
rect 2542 1857 2548 1858
rect 2542 1853 2543 1857
rect 2547 1853 2548 1857
rect 2542 1852 2548 1853
rect 2406 1839 2412 1840
rect 2406 1835 2407 1839
rect 2411 1835 2412 1839
rect 2406 1834 2412 1835
rect 2440 1827 2442 1852
rect 2526 1839 2532 1840
rect 2526 1835 2527 1839
rect 2531 1835 2532 1839
rect 2526 1834 2532 1835
rect 1807 1826 1811 1827
rect 1767 1822 1771 1823
rect 1807 1821 1811 1822
rect 2015 1826 2019 1827
rect 2015 1821 2019 1822
rect 2103 1826 2107 1827
rect 2103 1821 2107 1822
rect 2111 1826 2115 1827
rect 2111 1821 2115 1822
rect 2191 1826 2195 1827
rect 2191 1821 2195 1822
rect 2215 1826 2219 1827
rect 2215 1821 2219 1822
rect 2279 1826 2283 1827
rect 2306 1826 2312 1827
rect 2327 1826 2331 1827
rect 2279 1821 2283 1822
rect 2327 1821 2331 1822
rect 2367 1826 2371 1827
rect 2367 1821 2371 1822
rect 2439 1826 2443 1827
rect 2439 1821 2443 1822
rect 2455 1826 2459 1827
rect 2455 1821 2459 1822
rect 1767 1817 1771 1818
rect 1734 1815 1740 1816
rect 1734 1811 1735 1815
rect 1739 1811 1740 1815
rect 1734 1810 1740 1811
rect 1768 1801 1770 1817
rect 1808 1805 1810 1821
rect 1806 1804 1812 1805
rect 2104 1804 2106 1821
rect 2192 1804 2194 1821
rect 2206 1819 2212 1820
rect 2206 1815 2207 1819
rect 2211 1815 2212 1819
rect 2206 1814 2212 1815
rect 2262 1819 2268 1820
rect 2262 1815 2263 1819
rect 2267 1815 2268 1819
rect 2262 1814 2268 1815
rect 1766 1800 1772 1801
rect 1670 1799 1676 1800
rect 1670 1795 1671 1799
rect 1675 1795 1676 1799
rect 1766 1796 1767 1800
rect 1771 1796 1772 1800
rect 1806 1800 1807 1804
rect 1811 1800 1812 1804
rect 1806 1799 1812 1800
rect 2102 1803 2108 1804
rect 2102 1799 2103 1803
rect 2107 1799 2108 1803
rect 2102 1798 2108 1799
rect 2190 1803 2196 1804
rect 2190 1799 2191 1803
rect 2195 1799 2196 1803
rect 2190 1798 2196 1799
rect 1766 1795 1772 1796
rect 1670 1794 1676 1795
rect 830 1791 836 1792
rect 830 1787 831 1791
rect 835 1787 836 1791
rect 830 1786 836 1787
rect 958 1791 964 1792
rect 958 1787 959 1791
rect 963 1787 964 1791
rect 958 1786 964 1787
rect 1094 1791 1100 1792
rect 1094 1787 1095 1791
rect 1099 1787 1100 1791
rect 1094 1786 1100 1787
rect 1222 1791 1228 1792
rect 1222 1787 1223 1791
rect 1227 1787 1228 1791
rect 1222 1786 1228 1787
rect 1358 1791 1364 1792
rect 1358 1787 1359 1791
rect 1363 1787 1364 1791
rect 1358 1786 1364 1787
rect 1486 1791 1492 1792
rect 1486 1787 1487 1791
rect 1491 1787 1492 1791
rect 1486 1786 1492 1787
rect 1614 1791 1620 1792
rect 1614 1787 1615 1791
rect 1619 1787 1620 1791
rect 1614 1786 1620 1787
rect 1806 1787 1812 1788
rect 1362 1783 1368 1784
rect 886 1780 892 1781
rect 886 1776 887 1780
rect 891 1776 892 1780
rect 886 1775 892 1776
rect 1022 1780 1028 1781
rect 1022 1776 1023 1780
rect 1027 1776 1028 1780
rect 1022 1775 1028 1776
rect 1150 1780 1156 1781
rect 1150 1776 1151 1780
rect 1155 1776 1156 1780
rect 1150 1775 1156 1776
rect 1278 1780 1284 1781
rect 1278 1776 1279 1780
rect 1283 1776 1284 1780
rect 1362 1779 1363 1783
rect 1367 1779 1368 1783
rect 1766 1783 1772 1784
rect 1362 1778 1368 1779
rect 1406 1780 1412 1781
rect 1278 1775 1284 1776
rect 888 1755 890 1775
rect 1024 1755 1026 1775
rect 1152 1755 1154 1775
rect 1280 1755 1282 1775
rect 847 1754 851 1755
rect 847 1749 851 1750
rect 887 1754 891 1755
rect 887 1749 891 1750
rect 951 1754 955 1755
rect 951 1749 955 1750
rect 1023 1754 1027 1755
rect 1023 1749 1027 1750
rect 1055 1754 1059 1755
rect 1055 1749 1059 1750
rect 1151 1754 1155 1755
rect 1151 1749 1155 1750
rect 1159 1754 1163 1755
rect 1159 1749 1163 1750
rect 1271 1754 1275 1755
rect 1271 1749 1275 1750
rect 1279 1754 1283 1755
rect 1279 1749 1283 1750
rect 848 1733 850 1749
rect 952 1733 954 1749
rect 1056 1733 1058 1749
rect 1160 1733 1162 1749
rect 1272 1733 1274 1749
rect 846 1732 852 1733
rect 846 1728 847 1732
rect 851 1728 852 1732
rect 846 1727 852 1728
rect 950 1732 956 1733
rect 950 1728 951 1732
rect 955 1728 956 1732
rect 950 1727 956 1728
rect 1054 1732 1060 1733
rect 1054 1728 1055 1732
rect 1059 1728 1060 1732
rect 1054 1727 1060 1728
rect 1158 1732 1164 1733
rect 1158 1728 1159 1732
rect 1163 1728 1164 1732
rect 1158 1727 1164 1728
rect 1270 1732 1276 1733
rect 1270 1728 1271 1732
rect 1275 1728 1276 1732
rect 1270 1727 1276 1728
rect 814 1723 820 1724
rect 814 1719 815 1723
rect 819 1719 820 1723
rect 814 1718 820 1719
rect 822 1723 828 1724
rect 822 1719 823 1723
rect 827 1719 828 1723
rect 822 1718 828 1719
rect 1030 1723 1036 1724
rect 1030 1719 1031 1723
rect 1035 1719 1036 1723
rect 1030 1718 1036 1719
rect 1134 1723 1140 1724
rect 1134 1719 1135 1723
rect 1139 1719 1140 1723
rect 1134 1718 1140 1719
rect 1238 1723 1244 1724
rect 1238 1719 1239 1723
rect 1243 1719 1244 1723
rect 1238 1718 1244 1719
rect 1350 1723 1356 1724
rect 1350 1719 1351 1723
rect 1355 1719 1356 1723
rect 1350 1718 1356 1719
rect 742 1713 748 1714
rect 742 1709 743 1713
rect 747 1709 748 1713
rect 742 1708 748 1709
rect 702 1695 708 1696
rect 702 1691 703 1695
rect 707 1691 708 1695
rect 702 1690 708 1691
rect 734 1695 740 1696
rect 734 1691 735 1695
rect 739 1691 740 1695
rect 734 1690 740 1691
rect 535 1686 539 1687
rect 535 1681 539 1682
rect 575 1686 579 1687
rect 575 1681 579 1682
rect 639 1686 643 1687
rect 639 1681 643 1682
rect 663 1686 667 1687
rect 663 1681 667 1682
rect 502 1679 508 1680
rect 502 1675 503 1679
rect 507 1675 508 1679
rect 502 1674 508 1675
rect 576 1664 578 1681
rect 664 1664 666 1681
rect 670 1679 676 1680
rect 670 1675 671 1679
rect 675 1675 676 1679
rect 670 1674 676 1675
rect 110 1660 111 1664
rect 115 1660 116 1664
rect 110 1659 116 1660
rect 398 1663 404 1664
rect 398 1659 399 1663
rect 403 1659 404 1663
rect 398 1658 404 1659
rect 486 1663 492 1664
rect 486 1659 487 1663
rect 491 1659 492 1663
rect 486 1658 492 1659
rect 574 1663 580 1664
rect 574 1659 575 1663
rect 579 1659 580 1663
rect 574 1658 580 1659
rect 662 1663 668 1664
rect 662 1659 663 1663
rect 667 1659 668 1663
rect 662 1658 668 1659
rect 558 1651 564 1652
rect 110 1647 116 1648
rect 110 1643 111 1647
rect 115 1643 116 1647
rect 558 1647 559 1651
rect 563 1647 564 1651
rect 558 1646 564 1647
rect 110 1642 116 1643
rect 398 1644 404 1645
rect 112 1619 114 1642
rect 398 1640 399 1644
rect 403 1640 404 1644
rect 398 1639 404 1640
rect 486 1644 492 1645
rect 486 1640 487 1644
rect 491 1640 492 1644
rect 486 1639 492 1640
rect 400 1619 402 1639
rect 488 1619 490 1639
rect 111 1618 115 1619
rect 111 1613 115 1614
rect 279 1618 283 1619
rect 279 1613 283 1614
rect 383 1618 387 1619
rect 383 1613 387 1614
rect 399 1618 403 1619
rect 399 1613 403 1614
rect 487 1618 491 1619
rect 487 1613 491 1614
rect 495 1618 499 1619
rect 495 1613 499 1614
rect 112 1594 114 1613
rect 280 1597 282 1613
rect 384 1597 386 1613
rect 496 1597 498 1613
rect 278 1596 284 1597
rect 110 1593 116 1594
rect 110 1589 111 1593
rect 115 1589 116 1593
rect 278 1592 279 1596
rect 283 1592 284 1596
rect 278 1591 284 1592
rect 382 1596 388 1597
rect 382 1592 383 1596
rect 387 1592 388 1596
rect 382 1591 388 1592
rect 494 1596 500 1597
rect 494 1592 495 1596
rect 499 1592 500 1596
rect 494 1591 500 1592
rect 110 1588 116 1589
rect 350 1587 356 1588
rect 350 1583 351 1587
rect 355 1583 356 1587
rect 350 1582 356 1583
rect 454 1587 460 1588
rect 454 1583 455 1587
rect 459 1583 460 1587
rect 454 1582 460 1583
rect 462 1587 468 1588
rect 462 1583 463 1587
rect 467 1583 468 1587
rect 462 1582 468 1583
rect 278 1577 284 1578
rect 110 1576 116 1577
rect 110 1572 111 1576
rect 115 1572 116 1576
rect 278 1573 279 1577
rect 283 1573 284 1577
rect 278 1572 284 1573
rect 110 1571 116 1572
rect 112 1547 114 1571
rect 280 1547 282 1572
rect 352 1560 354 1582
rect 382 1577 388 1578
rect 382 1573 383 1577
rect 387 1573 388 1577
rect 382 1572 388 1573
rect 350 1559 356 1560
rect 350 1555 351 1559
rect 355 1555 356 1559
rect 350 1554 356 1555
rect 384 1547 386 1572
rect 111 1546 115 1547
rect 111 1541 115 1542
rect 183 1546 187 1547
rect 183 1541 187 1542
rect 279 1546 283 1547
rect 279 1541 283 1542
rect 327 1546 331 1547
rect 327 1541 331 1542
rect 383 1546 387 1547
rect 383 1541 387 1542
rect 112 1525 114 1541
rect 110 1524 116 1525
rect 184 1524 186 1541
rect 290 1539 296 1540
rect 290 1535 291 1539
rect 295 1535 296 1539
rect 290 1534 296 1535
rect 110 1520 111 1524
rect 115 1520 116 1524
rect 110 1519 116 1520
rect 182 1523 188 1524
rect 182 1519 183 1523
rect 187 1519 188 1523
rect 182 1518 188 1519
rect 292 1516 294 1534
rect 328 1524 330 1541
rect 456 1540 458 1582
rect 464 1552 466 1582
rect 494 1577 500 1578
rect 494 1573 495 1577
rect 499 1573 500 1577
rect 494 1572 500 1573
rect 462 1551 468 1552
rect 462 1547 463 1551
rect 467 1547 468 1551
rect 496 1547 498 1572
rect 560 1560 562 1646
rect 574 1644 580 1645
rect 574 1640 575 1644
rect 579 1640 580 1644
rect 574 1639 580 1640
rect 662 1644 668 1645
rect 662 1640 663 1644
rect 667 1640 668 1644
rect 662 1639 668 1640
rect 576 1619 578 1639
rect 664 1619 666 1639
rect 575 1618 579 1619
rect 575 1613 579 1614
rect 607 1618 611 1619
rect 607 1613 611 1614
rect 663 1618 667 1619
rect 663 1613 667 1614
rect 608 1597 610 1613
rect 606 1596 612 1597
rect 606 1592 607 1596
rect 611 1592 612 1596
rect 606 1591 612 1592
rect 672 1588 674 1674
rect 736 1656 738 1690
rect 744 1687 746 1708
rect 816 1696 818 1718
rect 846 1713 852 1714
rect 846 1709 847 1713
rect 851 1709 852 1713
rect 846 1708 852 1709
rect 950 1713 956 1714
rect 950 1709 951 1713
rect 955 1709 956 1713
rect 950 1708 956 1709
rect 814 1695 820 1696
rect 814 1691 815 1695
rect 819 1691 820 1695
rect 814 1690 820 1691
rect 848 1687 850 1708
rect 952 1687 954 1708
rect 1032 1696 1034 1718
rect 1054 1713 1060 1714
rect 1054 1709 1055 1713
rect 1059 1709 1060 1713
rect 1054 1708 1060 1709
rect 1030 1695 1036 1696
rect 1030 1691 1031 1695
rect 1035 1691 1036 1695
rect 1030 1690 1036 1691
rect 1056 1687 1058 1708
rect 1078 1707 1084 1708
rect 1078 1703 1079 1707
rect 1083 1703 1084 1707
rect 1078 1702 1084 1703
rect 1080 1699 1082 1702
rect 1080 1697 1086 1699
rect 743 1686 747 1687
rect 743 1681 747 1682
rect 759 1686 763 1687
rect 759 1681 763 1682
rect 847 1686 851 1687
rect 847 1681 851 1682
rect 855 1686 859 1687
rect 855 1681 859 1682
rect 951 1686 955 1687
rect 951 1681 955 1682
rect 1047 1686 1051 1687
rect 1047 1681 1051 1682
rect 1055 1686 1059 1687
rect 1055 1681 1059 1682
rect 760 1664 762 1681
rect 838 1679 844 1680
rect 838 1675 839 1679
rect 843 1675 844 1679
rect 838 1674 844 1675
rect 758 1663 764 1664
rect 758 1659 759 1663
rect 763 1659 764 1663
rect 758 1658 764 1659
rect 840 1656 842 1674
rect 856 1664 858 1681
rect 952 1664 954 1681
rect 1048 1664 1050 1681
rect 1084 1680 1086 1697
rect 1136 1696 1138 1718
rect 1158 1713 1164 1714
rect 1158 1709 1159 1713
rect 1163 1709 1164 1713
rect 1158 1708 1164 1709
rect 1134 1695 1140 1696
rect 1134 1691 1135 1695
rect 1139 1691 1140 1695
rect 1134 1690 1140 1691
rect 1126 1687 1132 1688
rect 1160 1687 1162 1708
rect 1240 1696 1242 1718
rect 1270 1713 1276 1714
rect 1270 1709 1271 1713
rect 1275 1709 1276 1713
rect 1270 1708 1276 1709
rect 1238 1695 1244 1696
rect 1238 1691 1239 1695
rect 1243 1691 1244 1695
rect 1238 1690 1244 1691
rect 1272 1687 1274 1708
rect 1352 1696 1354 1718
rect 1364 1696 1366 1778
rect 1406 1776 1407 1780
rect 1411 1776 1412 1780
rect 1406 1775 1412 1776
rect 1534 1780 1540 1781
rect 1534 1776 1535 1780
rect 1539 1776 1540 1780
rect 1534 1775 1540 1776
rect 1670 1780 1676 1781
rect 1670 1776 1671 1780
rect 1675 1776 1676 1780
rect 1766 1779 1767 1783
rect 1771 1779 1772 1783
rect 1806 1783 1807 1787
rect 1811 1783 1812 1787
rect 1806 1782 1812 1783
rect 2102 1784 2108 1785
rect 1766 1778 1772 1779
rect 1670 1775 1676 1776
rect 1408 1755 1410 1775
rect 1536 1755 1538 1775
rect 1672 1755 1674 1775
rect 1768 1755 1770 1778
rect 1383 1754 1387 1755
rect 1383 1749 1387 1750
rect 1407 1754 1411 1755
rect 1407 1749 1411 1750
rect 1535 1754 1539 1755
rect 1535 1749 1539 1750
rect 1671 1754 1675 1755
rect 1671 1749 1675 1750
rect 1767 1754 1771 1755
rect 1808 1751 1810 1782
rect 2102 1780 2103 1784
rect 2107 1780 2108 1784
rect 2102 1779 2108 1780
rect 2190 1784 2196 1785
rect 2190 1780 2191 1784
rect 2195 1780 2196 1784
rect 2190 1779 2196 1780
rect 2104 1751 2106 1779
rect 2192 1751 2194 1779
rect 1767 1749 1771 1750
rect 1807 1750 1811 1751
rect 1384 1733 1386 1749
rect 1382 1732 1388 1733
rect 1382 1728 1383 1732
rect 1387 1728 1388 1732
rect 1768 1730 1770 1749
rect 1807 1745 1811 1746
rect 2103 1750 2107 1751
rect 2103 1745 2107 1746
rect 2143 1750 2147 1751
rect 2143 1745 2147 1746
rect 2191 1750 2195 1751
rect 2191 1745 2195 1746
rect 1382 1727 1388 1728
rect 1766 1729 1772 1730
rect 1766 1725 1767 1729
rect 1771 1725 1772 1729
rect 1808 1726 1810 1745
rect 2144 1729 2146 1745
rect 2142 1728 2148 1729
rect 1766 1724 1772 1725
rect 1806 1725 1812 1726
rect 1806 1721 1807 1725
rect 1811 1721 1812 1725
rect 2142 1724 2143 1728
rect 2147 1724 2148 1728
rect 2142 1723 2148 1724
rect 1806 1720 1812 1721
rect 2208 1720 2210 1814
rect 2264 1796 2266 1814
rect 2280 1804 2282 1821
rect 2350 1819 2356 1820
rect 2350 1815 2351 1819
rect 2355 1815 2356 1819
rect 2350 1814 2356 1815
rect 2278 1803 2284 1804
rect 2278 1799 2279 1803
rect 2283 1799 2284 1803
rect 2278 1798 2284 1799
rect 2352 1796 2354 1814
rect 2368 1804 2370 1821
rect 2456 1804 2458 1821
rect 2366 1803 2372 1804
rect 2366 1799 2367 1803
rect 2371 1799 2372 1803
rect 2366 1798 2372 1799
rect 2454 1803 2460 1804
rect 2454 1799 2455 1803
rect 2459 1799 2460 1803
rect 2454 1798 2460 1799
rect 2528 1796 2530 1834
rect 2544 1827 2546 1852
rect 2640 1840 2642 1922
rect 2710 1920 2711 1924
rect 2715 1920 2716 1924
rect 2710 1919 2716 1920
rect 2830 1924 2836 1925
rect 2830 1920 2831 1924
rect 2835 1920 2836 1924
rect 2830 1919 2836 1920
rect 2950 1924 2956 1925
rect 2950 1920 2951 1924
rect 2955 1920 2956 1924
rect 2950 1919 2956 1920
rect 3062 1924 3068 1925
rect 3062 1920 3063 1924
rect 3067 1920 3068 1924
rect 3062 1919 3068 1920
rect 3166 1924 3172 1925
rect 3166 1920 3167 1924
rect 3171 1920 3172 1924
rect 3166 1919 3172 1920
rect 3278 1924 3284 1925
rect 3278 1920 3279 1924
rect 3283 1920 3284 1924
rect 3278 1919 3284 1920
rect 3366 1924 3372 1925
rect 3366 1920 3367 1924
rect 3371 1920 3372 1924
rect 3462 1923 3463 1927
rect 3467 1923 3468 1927
rect 3462 1922 3468 1923
rect 3366 1919 3372 1920
rect 2712 1899 2714 1919
rect 2832 1899 2834 1919
rect 2952 1899 2954 1919
rect 3064 1899 3066 1919
rect 3168 1899 3170 1919
rect 3280 1899 3282 1919
rect 3368 1899 3370 1919
rect 3464 1899 3466 1922
rect 2647 1898 2651 1899
rect 2647 1893 2651 1894
rect 2711 1898 2715 1899
rect 2711 1893 2715 1894
rect 2759 1898 2763 1899
rect 2759 1893 2763 1894
rect 2831 1898 2835 1899
rect 2831 1893 2835 1894
rect 2871 1898 2875 1899
rect 2871 1893 2875 1894
rect 2951 1898 2955 1899
rect 2951 1893 2955 1894
rect 2983 1898 2987 1899
rect 2983 1893 2987 1894
rect 3063 1898 3067 1899
rect 3063 1893 3067 1894
rect 3167 1898 3171 1899
rect 3167 1893 3171 1894
rect 3279 1898 3283 1899
rect 3279 1893 3283 1894
rect 3367 1898 3371 1899
rect 3367 1893 3371 1894
rect 3463 1898 3467 1899
rect 3463 1893 3467 1894
rect 2648 1877 2650 1893
rect 2760 1877 2762 1893
rect 2872 1877 2874 1893
rect 2984 1877 2986 1893
rect 2646 1876 2652 1877
rect 2646 1872 2647 1876
rect 2651 1872 2652 1876
rect 2646 1871 2652 1872
rect 2758 1876 2764 1877
rect 2758 1872 2759 1876
rect 2763 1872 2764 1876
rect 2758 1871 2764 1872
rect 2870 1876 2876 1877
rect 2870 1872 2871 1876
rect 2875 1872 2876 1876
rect 2870 1871 2876 1872
rect 2982 1876 2988 1877
rect 2982 1872 2983 1876
rect 2987 1872 2988 1876
rect 3464 1874 3466 1893
rect 2982 1871 2988 1872
rect 3462 1873 3468 1874
rect 3462 1869 3463 1873
rect 3467 1869 3468 1873
rect 3462 1868 3468 1869
rect 2718 1867 2724 1868
rect 2718 1863 2719 1867
rect 2723 1863 2724 1867
rect 2718 1862 2724 1863
rect 2830 1867 2836 1868
rect 2830 1863 2831 1867
rect 2835 1863 2836 1867
rect 2830 1862 2836 1863
rect 2942 1867 2948 1868
rect 2942 1863 2943 1867
rect 2947 1863 2948 1867
rect 2942 1862 2948 1863
rect 2646 1857 2652 1858
rect 2646 1853 2647 1857
rect 2651 1853 2652 1857
rect 2646 1852 2652 1853
rect 2638 1839 2644 1840
rect 2638 1835 2639 1839
rect 2643 1835 2644 1839
rect 2638 1834 2644 1835
rect 2648 1827 2650 1852
rect 2720 1840 2722 1862
rect 2758 1857 2764 1858
rect 2758 1853 2759 1857
rect 2763 1853 2764 1857
rect 2758 1852 2764 1853
rect 2718 1839 2724 1840
rect 2718 1835 2719 1839
rect 2723 1835 2724 1839
rect 2718 1834 2724 1835
rect 2710 1827 2716 1828
rect 2760 1827 2762 1852
rect 2832 1840 2834 1862
rect 2870 1857 2876 1858
rect 2870 1853 2871 1857
rect 2875 1853 2876 1857
rect 2870 1852 2876 1853
rect 2830 1839 2836 1840
rect 2830 1835 2831 1839
rect 2835 1835 2836 1839
rect 2830 1834 2836 1835
rect 2872 1827 2874 1852
rect 2944 1840 2946 1862
rect 2982 1857 2988 1858
rect 2982 1853 2983 1857
rect 2987 1853 2988 1857
rect 2982 1852 2988 1853
rect 3462 1856 3468 1857
rect 3462 1852 3463 1856
rect 3467 1852 3468 1856
rect 2942 1839 2948 1840
rect 2942 1835 2943 1839
rect 2947 1835 2948 1839
rect 2942 1834 2948 1835
rect 2984 1827 2986 1852
rect 3462 1851 3468 1852
rect 3464 1827 3466 1851
rect 2543 1826 2547 1827
rect 2543 1821 2547 1822
rect 2631 1826 2635 1827
rect 2631 1821 2635 1822
rect 2647 1826 2651 1827
rect 2710 1823 2711 1827
rect 2715 1823 2716 1827
rect 2710 1822 2716 1823
rect 2719 1826 2723 1827
rect 2647 1821 2651 1822
rect 2544 1804 2546 1821
rect 2614 1819 2620 1820
rect 2614 1815 2615 1819
rect 2619 1815 2620 1819
rect 2614 1814 2620 1815
rect 2542 1803 2548 1804
rect 2542 1799 2543 1803
rect 2547 1799 2548 1803
rect 2542 1798 2548 1799
rect 2616 1796 2618 1814
rect 2632 1804 2634 1821
rect 2630 1803 2636 1804
rect 2630 1799 2631 1803
rect 2635 1799 2636 1803
rect 2630 1798 2636 1799
rect 2712 1796 2714 1822
rect 2719 1821 2723 1822
rect 2759 1826 2763 1827
rect 2759 1821 2763 1822
rect 2807 1826 2811 1827
rect 2807 1821 2811 1822
rect 2871 1826 2875 1827
rect 2871 1821 2875 1822
rect 2895 1826 2899 1827
rect 2895 1821 2899 1822
rect 2983 1826 2987 1827
rect 2983 1821 2987 1822
rect 3463 1826 3467 1827
rect 3463 1821 3467 1822
rect 2720 1804 2722 1821
rect 2808 1804 2810 1821
rect 2886 1819 2892 1820
rect 2886 1815 2887 1819
rect 2891 1815 2892 1819
rect 2886 1814 2892 1815
rect 2718 1803 2724 1804
rect 2718 1799 2719 1803
rect 2723 1799 2724 1803
rect 2718 1798 2724 1799
rect 2806 1803 2812 1804
rect 2806 1799 2807 1803
rect 2811 1799 2812 1803
rect 2806 1798 2812 1799
rect 2888 1796 2890 1814
rect 2896 1804 2898 1821
rect 3464 1805 3466 1821
rect 3462 1804 3468 1805
rect 2894 1803 2900 1804
rect 2894 1799 2895 1803
rect 2899 1799 2900 1803
rect 3462 1800 3463 1804
rect 3467 1800 3468 1804
rect 3462 1799 3468 1800
rect 2894 1798 2900 1799
rect 2262 1795 2268 1796
rect 2262 1791 2263 1795
rect 2267 1791 2268 1795
rect 2262 1790 2268 1791
rect 2350 1795 2356 1796
rect 2350 1791 2351 1795
rect 2355 1791 2356 1795
rect 2350 1790 2356 1791
rect 2526 1795 2532 1796
rect 2526 1791 2527 1795
rect 2531 1791 2532 1795
rect 2526 1790 2532 1791
rect 2614 1795 2620 1796
rect 2614 1791 2615 1795
rect 2619 1791 2620 1795
rect 2710 1795 2716 1796
rect 2614 1790 2620 1791
rect 2702 1791 2708 1792
rect 2702 1787 2703 1791
rect 2707 1787 2708 1791
rect 2710 1791 2711 1795
rect 2715 1791 2716 1795
rect 2710 1790 2716 1791
rect 2886 1795 2892 1796
rect 2886 1791 2887 1795
rect 2891 1791 2892 1795
rect 2886 1790 2892 1791
rect 2702 1786 2708 1787
rect 3462 1787 3468 1788
rect 2278 1784 2284 1785
rect 2278 1780 2279 1784
rect 2283 1780 2284 1784
rect 2278 1779 2284 1780
rect 2366 1784 2372 1785
rect 2366 1780 2367 1784
rect 2371 1780 2372 1784
rect 2366 1779 2372 1780
rect 2454 1784 2460 1785
rect 2454 1780 2455 1784
rect 2459 1780 2460 1784
rect 2454 1779 2460 1780
rect 2542 1784 2548 1785
rect 2542 1780 2543 1784
rect 2547 1780 2548 1784
rect 2542 1779 2548 1780
rect 2630 1784 2636 1785
rect 2630 1780 2631 1784
rect 2635 1780 2636 1784
rect 2630 1779 2636 1780
rect 2280 1751 2282 1779
rect 2368 1751 2370 1779
rect 2456 1751 2458 1779
rect 2544 1751 2546 1779
rect 2632 1751 2634 1779
rect 2231 1750 2235 1751
rect 2231 1745 2235 1746
rect 2279 1750 2283 1751
rect 2279 1745 2283 1746
rect 2319 1750 2323 1751
rect 2319 1745 2323 1746
rect 2367 1750 2371 1751
rect 2367 1745 2371 1746
rect 2407 1750 2411 1751
rect 2407 1745 2411 1746
rect 2455 1750 2459 1751
rect 2455 1745 2459 1746
rect 2495 1750 2499 1751
rect 2495 1745 2499 1746
rect 2543 1750 2547 1751
rect 2543 1745 2547 1746
rect 2583 1750 2587 1751
rect 2583 1745 2587 1746
rect 2631 1750 2635 1751
rect 2631 1745 2635 1746
rect 2671 1750 2675 1751
rect 2671 1745 2675 1746
rect 2232 1729 2234 1745
rect 2320 1729 2322 1745
rect 2408 1729 2410 1745
rect 2496 1729 2498 1745
rect 2584 1729 2586 1745
rect 2672 1729 2674 1745
rect 2230 1728 2236 1729
rect 2230 1724 2231 1728
rect 2235 1724 2236 1728
rect 2230 1723 2236 1724
rect 2318 1728 2324 1729
rect 2318 1724 2319 1728
rect 2323 1724 2324 1728
rect 2318 1723 2324 1724
rect 2406 1728 2412 1729
rect 2406 1724 2407 1728
rect 2411 1724 2412 1728
rect 2406 1723 2412 1724
rect 2494 1728 2500 1729
rect 2494 1724 2495 1728
rect 2499 1724 2500 1728
rect 2494 1723 2500 1724
rect 2582 1728 2588 1729
rect 2582 1724 2583 1728
rect 2587 1724 2588 1728
rect 2582 1723 2588 1724
rect 2670 1728 2676 1729
rect 2670 1724 2671 1728
rect 2675 1724 2676 1728
rect 2670 1723 2676 1724
rect 2206 1719 2212 1720
rect 2206 1715 2207 1719
rect 2211 1715 2212 1719
rect 2206 1714 2212 1715
rect 2222 1719 2228 1720
rect 2222 1715 2223 1719
rect 2227 1715 2228 1719
rect 2222 1714 2228 1715
rect 2310 1719 2316 1720
rect 2310 1715 2311 1719
rect 2315 1715 2316 1719
rect 2310 1714 2316 1715
rect 2398 1719 2404 1720
rect 2398 1715 2399 1719
rect 2403 1715 2404 1719
rect 2398 1714 2404 1715
rect 2486 1719 2492 1720
rect 2486 1715 2487 1719
rect 2491 1715 2492 1719
rect 2486 1714 2492 1715
rect 2646 1719 2652 1720
rect 2646 1715 2647 1719
rect 2651 1715 2652 1719
rect 2646 1714 2652 1715
rect 1382 1713 1388 1714
rect 1382 1709 1383 1713
rect 1387 1709 1388 1713
rect 1382 1708 1388 1709
rect 1766 1712 1772 1713
rect 1766 1708 1767 1712
rect 1771 1708 1772 1712
rect 2142 1709 2148 1710
rect 1350 1695 1356 1696
rect 1350 1691 1351 1695
rect 1355 1691 1356 1695
rect 1350 1690 1356 1691
rect 1362 1695 1368 1696
rect 1362 1691 1363 1695
rect 1367 1691 1368 1695
rect 1362 1690 1368 1691
rect 1384 1687 1386 1708
rect 1766 1707 1772 1708
rect 1806 1708 1812 1709
rect 1768 1687 1770 1707
rect 1806 1704 1807 1708
rect 1811 1704 1812 1708
rect 2142 1705 2143 1709
rect 2147 1705 2148 1709
rect 2142 1704 2148 1705
rect 1806 1703 1812 1704
rect 1126 1683 1127 1687
rect 1131 1683 1132 1687
rect 1126 1682 1132 1683
rect 1143 1686 1147 1687
rect 1082 1679 1088 1680
rect 1082 1675 1083 1679
rect 1087 1675 1088 1679
rect 1082 1674 1088 1675
rect 1118 1679 1124 1680
rect 1118 1675 1119 1679
rect 1123 1675 1124 1679
rect 1118 1674 1124 1675
rect 854 1663 860 1664
rect 854 1659 855 1663
rect 859 1659 860 1663
rect 854 1658 860 1659
rect 950 1663 956 1664
rect 950 1659 951 1663
rect 955 1659 956 1663
rect 950 1658 956 1659
rect 1046 1663 1052 1664
rect 1046 1659 1047 1663
rect 1051 1659 1052 1663
rect 1046 1658 1052 1659
rect 1120 1656 1122 1674
rect 1128 1656 1130 1682
rect 1143 1681 1147 1682
rect 1159 1686 1163 1687
rect 1159 1681 1163 1682
rect 1271 1686 1275 1687
rect 1271 1681 1275 1682
rect 1383 1686 1387 1687
rect 1383 1681 1387 1682
rect 1767 1686 1771 1687
rect 1808 1683 1810 1703
rect 2144 1683 2146 1704
rect 2224 1692 2226 1714
rect 2230 1709 2236 1710
rect 2230 1705 2231 1709
rect 2235 1705 2236 1709
rect 2230 1704 2236 1705
rect 2222 1691 2228 1692
rect 2222 1687 2223 1691
rect 2227 1687 2228 1691
rect 2222 1686 2228 1687
rect 2232 1683 2234 1704
rect 2312 1692 2314 1714
rect 2318 1709 2324 1710
rect 2318 1705 2319 1709
rect 2323 1705 2324 1709
rect 2318 1704 2324 1705
rect 2310 1691 2316 1692
rect 2310 1687 2311 1691
rect 2315 1687 2316 1691
rect 2310 1686 2316 1687
rect 2320 1683 2322 1704
rect 2400 1692 2402 1714
rect 2406 1709 2412 1710
rect 2406 1705 2407 1709
rect 2411 1705 2412 1709
rect 2406 1704 2412 1705
rect 2398 1691 2404 1692
rect 2398 1687 2399 1691
rect 2403 1687 2404 1691
rect 2398 1686 2404 1687
rect 2408 1683 2410 1704
rect 2488 1692 2490 1714
rect 2494 1709 2500 1710
rect 2494 1705 2495 1709
rect 2499 1705 2500 1709
rect 2494 1704 2500 1705
rect 2582 1709 2588 1710
rect 2582 1705 2583 1709
rect 2587 1705 2588 1709
rect 2582 1704 2588 1705
rect 2486 1691 2492 1692
rect 2486 1687 2487 1691
rect 2491 1687 2492 1691
rect 2486 1686 2492 1687
rect 2446 1683 2452 1684
rect 2496 1683 2498 1704
rect 2526 1691 2532 1692
rect 2526 1687 2527 1691
rect 2531 1687 2532 1691
rect 2526 1686 2532 1687
rect 1767 1681 1771 1682
rect 1807 1682 1811 1683
rect 1144 1664 1146 1681
rect 1768 1665 1770 1681
rect 1807 1677 1811 1678
rect 2103 1682 2107 1683
rect 2103 1677 2107 1678
rect 2143 1682 2147 1683
rect 2143 1677 2147 1678
rect 2191 1682 2195 1683
rect 2191 1677 2195 1678
rect 2231 1682 2235 1683
rect 2231 1677 2235 1678
rect 2279 1682 2283 1683
rect 2279 1677 2283 1678
rect 2319 1682 2323 1683
rect 2319 1677 2323 1678
rect 2367 1682 2371 1683
rect 2367 1677 2371 1678
rect 2407 1682 2411 1683
rect 2446 1679 2447 1683
rect 2451 1679 2452 1683
rect 2446 1678 2452 1679
rect 2455 1682 2459 1683
rect 2407 1677 2411 1678
rect 1766 1664 1772 1665
rect 1142 1663 1148 1664
rect 1142 1659 1143 1663
rect 1147 1659 1148 1663
rect 1766 1660 1767 1664
rect 1771 1660 1772 1664
rect 1808 1661 1810 1677
rect 1766 1659 1772 1660
rect 1806 1660 1812 1661
rect 2104 1660 2106 1677
rect 2174 1675 2180 1676
rect 2174 1671 2175 1675
rect 2179 1671 2180 1675
rect 2174 1670 2180 1671
rect 1142 1658 1148 1659
rect 1806 1656 1807 1660
rect 1811 1656 1812 1660
rect 734 1655 740 1656
rect 734 1651 735 1655
rect 739 1651 740 1655
rect 734 1650 740 1651
rect 838 1655 844 1656
rect 838 1651 839 1655
rect 843 1651 844 1655
rect 838 1650 844 1651
rect 1118 1655 1124 1656
rect 1118 1651 1119 1655
rect 1123 1651 1124 1655
rect 1118 1650 1124 1651
rect 1126 1655 1132 1656
rect 1806 1655 1812 1656
rect 2102 1659 2108 1660
rect 2102 1655 2103 1659
rect 2107 1655 2108 1659
rect 1126 1651 1127 1655
rect 1131 1651 1132 1655
rect 2102 1654 2108 1655
rect 2176 1652 2178 1670
rect 2192 1660 2194 1677
rect 2262 1675 2268 1676
rect 2262 1671 2263 1675
rect 2267 1671 2268 1675
rect 2262 1670 2268 1671
rect 2190 1659 2196 1660
rect 2190 1655 2191 1659
rect 2195 1655 2196 1659
rect 2190 1654 2196 1655
rect 2264 1652 2266 1670
rect 2280 1660 2282 1677
rect 2350 1675 2356 1676
rect 2350 1671 2351 1675
rect 2355 1671 2356 1675
rect 2350 1670 2356 1671
rect 2278 1659 2284 1660
rect 2278 1655 2279 1659
rect 2283 1655 2284 1659
rect 2278 1654 2284 1655
rect 2352 1652 2354 1670
rect 2368 1660 2370 1677
rect 2438 1675 2444 1676
rect 2438 1671 2439 1675
rect 2443 1671 2444 1675
rect 2438 1670 2444 1671
rect 2366 1659 2372 1660
rect 2366 1655 2367 1659
rect 2371 1655 2372 1659
rect 2366 1654 2372 1655
rect 2440 1652 2442 1670
rect 1126 1650 1132 1651
rect 2174 1651 2180 1652
rect 838 1647 844 1648
rect 758 1644 764 1645
rect 758 1640 759 1644
rect 763 1640 764 1644
rect 838 1643 839 1647
rect 843 1643 844 1647
rect 1766 1647 1772 1648
rect 838 1642 844 1643
rect 854 1644 860 1645
rect 758 1639 764 1640
rect 760 1619 762 1639
rect 719 1618 723 1619
rect 719 1613 723 1614
rect 759 1618 763 1619
rect 759 1613 763 1614
rect 831 1618 835 1619
rect 831 1613 835 1614
rect 720 1597 722 1613
rect 832 1597 834 1613
rect 718 1596 724 1597
rect 718 1592 719 1596
rect 723 1592 724 1596
rect 718 1591 724 1592
rect 830 1596 836 1597
rect 830 1592 831 1596
rect 835 1592 836 1596
rect 830 1591 836 1592
rect 670 1587 676 1588
rect 670 1583 671 1587
rect 675 1583 676 1587
rect 670 1582 676 1583
rect 686 1587 692 1588
rect 686 1583 687 1587
rect 691 1583 692 1587
rect 686 1582 692 1583
rect 606 1577 612 1578
rect 606 1573 607 1577
rect 611 1573 612 1577
rect 606 1572 612 1573
rect 558 1559 564 1560
rect 558 1555 559 1559
rect 563 1555 564 1559
rect 558 1554 564 1555
rect 608 1547 610 1572
rect 688 1560 690 1582
rect 718 1577 724 1578
rect 718 1573 719 1577
rect 723 1573 724 1577
rect 718 1572 724 1573
rect 830 1577 836 1578
rect 830 1573 831 1577
rect 835 1573 836 1577
rect 830 1572 836 1573
rect 686 1559 692 1560
rect 686 1555 687 1559
rect 691 1555 692 1559
rect 686 1554 692 1555
rect 694 1559 700 1560
rect 694 1555 695 1559
rect 699 1555 700 1559
rect 694 1554 700 1555
rect 462 1546 468 1547
rect 471 1546 475 1547
rect 471 1541 475 1542
rect 495 1546 499 1547
rect 495 1541 499 1542
rect 607 1546 611 1547
rect 607 1541 611 1542
rect 623 1546 627 1547
rect 623 1541 627 1542
rect 406 1539 412 1540
rect 406 1535 407 1539
rect 411 1535 412 1539
rect 406 1534 412 1535
rect 454 1539 460 1540
rect 454 1535 455 1539
rect 459 1535 460 1539
rect 454 1534 460 1535
rect 326 1523 332 1524
rect 326 1519 327 1523
rect 331 1519 332 1523
rect 326 1518 332 1519
rect 408 1516 410 1534
rect 472 1524 474 1541
rect 624 1524 626 1541
rect 470 1523 476 1524
rect 470 1519 471 1523
rect 475 1519 476 1523
rect 470 1518 476 1519
rect 622 1523 628 1524
rect 622 1519 623 1523
rect 627 1519 628 1523
rect 622 1518 628 1519
rect 696 1516 698 1554
rect 720 1547 722 1572
rect 832 1547 834 1572
rect 840 1560 842 1642
rect 854 1640 855 1644
rect 859 1640 860 1644
rect 854 1639 860 1640
rect 950 1644 956 1645
rect 950 1640 951 1644
rect 955 1640 956 1644
rect 950 1639 956 1640
rect 1046 1644 1052 1645
rect 1046 1640 1047 1644
rect 1051 1640 1052 1644
rect 1046 1639 1052 1640
rect 1142 1644 1148 1645
rect 1142 1640 1143 1644
rect 1147 1640 1148 1644
rect 1766 1643 1767 1647
rect 1771 1643 1772 1647
rect 2174 1647 2175 1651
rect 2179 1647 2180 1651
rect 2174 1646 2180 1647
rect 2262 1651 2268 1652
rect 2262 1647 2263 1651
rect 2267 1647 2268 1651
rect 2262 1646 2268 1647
rect 2350 1651 2356 1652
rect 2350 1647 2351 1651
rect 2355 1647 2356 1651
rect 2350 1646 2356 1647
rect 2438 1651 2444 1652
rect 2438 1647 2439 1651
rect 2443 1647 2444 1651
rect 2438 1646 2444 1647
rect 1766 1642 1772 1643
rect 1806 1643 1812 1644
rect 1142 1639 1148 1640
rect 856 1619 858 1639
rect 952 1619 954 1639
rect 1048 1619 1050 1639
rect 1144 1619 1146 1639
rect 1768 1619 1770 1642
rect 1806 1639 1807 1643
rect 1811 1639 1812 1643
rect 1806 1638 1812 1639
rect 2102 1640 2108 1641
rect 855 1618 859 1619
rect 855 1613 859 1614
rect 943 1618 947 1619
rect 943 1613 947 1614
rect 951 1618 955 1619
rect 951 1613 955 1614
rect 1047 1618 1051 1619
rect 1047 1613 1051 1614
rect 1055 1618 1059 1619
rect 1055 1613 1059 1614
rect 1143 1618 1147 1619
rect 1143 1613 1147 1614
rect 1167 1618 1171 1619
rect 1167 1613 1171 1614
rect 1279 1618 1283 1619
rect 1279 1613 1283 1614
rect 1767 1618 1771 1619
rect 1808 1615 1810 1638
rect 2102 1636 2103 1640
rect 2107 1636 2108 1640
rect 2102 1635 2108 1636
rect 2190 1640 2196 1641
rect 2190 1636 2191 1640
rect 2195 1636 2196 1640
rect 2190 1635 2196 1636
rect 2278 1640 2284 1641
rect 2278 1636 2279 1640
rect 2283 1636 2284 1640
rect 2278 1635 2284 1636
rect 2366 1640 2372 1641
rect 2366 1636 2367 1640
rect 2371 1636 2372 1640
rect 2366 1635 2372 1636
rect 2104 1615 2106 1635
rect 2192 1615 2194 1635
rect 2280 1615 2282 1635
rect 2368 1615 2370 1635
rect 1767 1613 1771 1614
rect 1807 1614 1811 1615
rect 944 1597 946 1613
rect 1056 1597 1058 1613
rect 1168 1597 1170 1613
rect 1280 1597 1282 1613
rect 942 1596 948 1597
rect 942 1592 943 1596
rect 947 1592 948 1596
rect 942 1591 948 1592
rect 1054 1596 1060 1597
rect 1054 1592 1055 1596
rect 1059 1592 1060 1596
rect 1054 1591 1060 1592
rect 1166 1596 1172 1597
rect 1166 1592 1167 1596
rect 1171 1592 1172 1596
rect 1166 1591 1172 1592
rect 1278 1596 1284 1597
rect 1278 1592 1279 1596
rect 1283 1592 1284 1596
rect 1768 1594 1770 1613
rect 1807 1609 1811 1610
rect 2063 1614 2067 1615
rect 2063 1609 2067 1610
rect 2103 1614 2107 1615
rect 2103 1609 2107 1610
rect 2159 1614 2163 1615
rect 2159 1609 2163 1610
rect 2191 1614 2195 1615
rect 2191 1609 2195 1610
rect 2255 1614 2259 1615
rect 2255 1609 2259 1610
rect 2279 1614 2283 1615
rect 2279 1609 2283 1610
rect 2359 1614 2363 1615
rect 2359 1609 2363 1610
rect 2367 1614 2371 1615
rect 2367 1609 2371 1610
rect 1278 1591 1284 1592
rect 1766 1593 1772 1594
rect 1766 1589 1767 1593
rect 1771 1589 1772 1593
rect 1808 1590 1810 1609
rect 2064 1593 2066 1609
rect 2160 1593 2162 1609
rect 2256 1593 2258 1609
rect 2360 1593 2362 1609
rect 2062 1592 2068 1593
rect 1766 1588 1772 1589
rect 1806 1589 1812 1590
rect 902 1587 908 1588
rect 902 1583 903 1587
rect 907 1583 908 1587
rect 902 1582 908 1583
rect 1014 1587 1020 1588
rect 1014 1583 1015 1587
rect 1019 1583 1020 1587
rect 1014 1582 1020 1583
rect 1126 1587 1132 1588
rect 1126 1583 1127 1587
rect 1131 1583 1132 1587
rect 1126 1582 1132 1583
rect 1238 1587 1244 1588
rect 1238 1583 1239 1587
rect 1243 1583 1244 1587
rect 1238 1582 1244 1583
rect 1246 1587 1252 1588
rect 1246 1583 1247 1587
rect 1251 1583 1252 1587
rect 1806 1585 1807 1589
rect 1811 1585 1812 1589
rect 2062 1588 2063 1592
rect 2067 1588 2068 1592
rect 2062 1587 2068 1588
rect 2158 1592 2164 1593
rect 2158 1588 2159 1592
rect 2163 1588 2164 1592
rect 2158 1587 2164 1588
rect 2254 1592 2260 1593
rect 2254 1588 2255 1592
rect 2259 1588 2260 1592
rect 2254 1587 2260 1588
rect 2358 1592 2364 1593
rect 2358 1588 2359 1592
rect 2363 1588 2364 1592
rect 2358 1587 2364 1588
rect 1806 1584 1812 1585
rect 2448 1584 2450 1678
rect 2455 1677 2459 1678
rect 2495 1682 2499 1683
rect 2495 1677 2499 1678
rect 2456 1660 2458 1677
rect 2454 1659 2460 1660
rect 2454 1655 2455 1659
rect 2459 1655 2460 1659
rect 2454 1654 2460 1655
rect 2528 1652 2530 1686
rect 2584 1683 2586 1704
rect 2543 1682 2547 1683
rect 2543 1677 2547 1678
rect 2583 1682 2587 1683
rect 2583 1677 2587 1678
rect 2631 1682 2635 1683
rect 2631 1677 2635 1678
rect 2544 1660 2546 1677
rect 2632 1660 2634 1677
rect 2648 1676 2650 1714
rect 2670 1709 2676 1710
rect 2670 1705 2671 1709
rect 2675 1705 2676 1709
rect 2670 1704 2676 1705
rect 2672 1683 2674 1704
rect 2704 1692 2706 1786
rect 2718 1784 2724 1785
rect 2718 1780 2719 1784
rect 2723 1780 2724 1784
rect 2718 1779 2724 1780
rect 2806 1784 2812 1785
rect 2806 1780 2807 1784
rect 2811 1780 2812 1784
rect 2806 1779 2812 1780
rect 2894 1784 2900 1785
rect 2894 1780 2895 1784
rect 2899 1780 2900 1784
rect 3462 1783 3463 1787
rect 3467 1783 3468 1787
rect 3462 1782 3468 1783
rect 2894 1779 2900 1780
rect 2720 1751 2722 1779
rect 2808 1751 2810 1779
rect 2896 1751 2898 1779
rect 3464 1751 3466 1782
rect 2719 1750 2723 1751
rect 2719 1745 2723 1746
rect 2759 1750 2763 1751
rect 2759 1745 2763 1746
rect 2807 1750 2811 1751
rect 2807 1745 2811 1746
rect 2847 1750 2851 1751
rect 2847 1745 2851 1746
rect 2895 1750 2899 1751
rect 2895 1745 2899 1746
rect 3463 1750 3467 1751
rect 3463 1745 3467 1746
rect 2760 1729 2762 1745
rect 2848 1729 2850 1745
rect 2758 1728 2764 1729
rect 2758 1724 2759 1728
rect 2763 1724 2764 1728
rect 2758 1723 2764 1724
rect 2846 1728 2852 1729
rect 2846 1724 2847 1728
rect 2851 1724 2852 1728
rect 3464 1726 3466 1745
rect 2846 1723 2852 1724
rect 3462 1725 3468 1726
rect 3462 1721 3463 1725
rect 3467 1721 3468 1725
rect 3462 1720 3468 1721
rect 2742 1719 2748 1720
rect 2742 1715 2743 1719
rect 2747 1715 2748 1719
rect 2742 1714 2748 1715
rect 2830 1719 2836 1720
rect 2830 1715 2831 1719
rect 2835 1715 2836 1719
rect 2830 1714 2836 1715
rect 2744 1692 2746 1714
rect 2758 1709 2764 1710
rect 2758 1705 2759 1709
rect 2763 1705 2764 1709
rect 2758 1704 2764 1705
rect 2702 1691 2708 1692
rect 2702 1687 2703 1691
rect 2707 1687 2708 1691
rect 2702 1686 2708 1687
rect 2742 1691 2748 1692
rect 2742 1687 2743 1691
rect 2747 1687 2748 1691
rect 2742 1686 2748 1687
rect 2760 1683 2762 1704
rect 2832 1692 2834 1714
rect 2846 1709 2852 1710
rect 2846 1705 2847 1709
rect 2851 1705 2852 1709
rect 2846 1704 2852 1705
rect 3462 1708 3468 1709
rect 3462 1704 3463 1708
rect 3467 1704 3468 1708
rect 2830 1691 2836 1692
rect 2830 1687 2831 1691
rect 2835 1687 2836 1691
rect 2830 1686 2836 1687
rect 2848 1683 2850 1704
rect 3462 1703 3468 1704
rect 3464 1683 3466 1703
rect 2671 1682 2675 1683
rect 2671 1677 2675 1678
rect 2719 1682 2723 1683
rect 2719 1677 2723 1678
rect 2759 1682 2763 1683
rect 2759 1677 2763 1678
rect 2807 1682 2811 1683
rect 2807 1677 2811 1678
rect 2847 1682 2851 1683
rect 2847 1677 2851 1678
rect 2895 1682 2899 1683
rect 2895 1677 2899 1678
rect 3463 1682 3467 1683
rect 3463 1677 3467 1678
rect 2646 1675 2652 1676
rect 2646 1671 2647 1675
rect 2651 1671 2652 1675
rect 2646 1670 2652 1671
rect 2702 1675 2708 1676
rect 2702 1671 2703 1675
rect 2707 1671 2708 1675
rect 2702 1670 2708 1671
rect 2542 1659 2548 1660
rect 2542 1655 2543 1659
rect 2547 1655 2548 1659
rect 2542 1654 2548 1655
rect 2630 1659 2636 1660
rect 2630 1655 2631 1659
rect 2635 1655 2636 1659
rect 2630 1654 2636 1655
rect 2704 1652 2706 1670
rect 2720 1660 2722 1677
rect 2790 1675 2796 1676
rect 2790 1671 2791 1675
rect 2795 1671 2796 1675
rect 2790 1670 2796 1671
rect 2718 1659 2724 1660
rect 2718 1655 2719 1659
rect 2723 1655 2724 1659
rect 2718 1654 2724 1655
rect 2792 1652 2794 1670
rect 2808 1660 2810 1677
rect 2878 1675 2884 1676
rect 2878 1671 2879 1675
rect 2883 1671 2884 1675
rect 2878 1670 2884 1671
rect 2806 1659 2812 1660
rect 2806 1655 2807 1659
rect 2811 1655 2812 1659
rect 2806 1654 2812 1655
rect 2880 1652 2882 1670
rect 2896 1660 2898 1677
rect 3464 1661 3466 1677
rect 3462 1660 3468 1661
rect 2894 1659 2900 1660
rect 2894 1655 2895 1659
rect 2899 1655 2900 1659
rect 3462 1656 3463 1660
rect 3467 1656 3468 1660
rect 3462 1655 3468 1656
rect 2894 1654 2900 1655
rect 2526 1651 2532 1652
rect 2526 1647 2527 1651
rect 2531 1647 2532 1651
rect 2526 1646 2532 1647
rect 2702 1651 2708 1652
rect 2702 1647 2703 1651
rect 2707 1647 2708 1651
rect 2702 1646 2708 1647
rect 2790 1651 2796 1652
rect 2790 1647 2791 1651
rect 2795 1647 2796 1651
rect 2790 1646 2796 1647
rect 2878 1651 2884 1652
rect 2878 1647 2879 1651
rect 2883 1647 2884 1651
rect 2878 1646 2884 1647
rect 3462 1643 3468 1644
rect 2454 1640 2460 1641
rect 2454 1636 2455 1640
rect 2459 1636 2460 1640
rect 2454 1635 2460 1636
rect 2542 1640 2548 1641
rect 2542 1636 2543 1640
rect 2547 1636 2548 1640
rect 2542 1635 2548 1636
rect 2630 1640 2636 1641
rect 2630 1636 2631 1640
rect 2635 1636 2636 1640
rect 2630 1635 2636 1636
rect 2718 1640 2724 1641
rect 2718 1636 2719 1640
rect 2723 1636 2724 1640
rect 2718 1635 2724 1636
rect 2806 1640 2812 1641
rect 2806 1636 2807 1640
rect 2811 1636 2812 1640
rect 2806 1635 2812 1636
rect 2894 1640 2900 1641
rect 2894 1636 2895 1640
rect 2899 1636 2900 1640
rect 3462 1639 3463 1643
rect 3467 1639 3468 1643
rect 3462 1638 3468 1639
rect 2894 1635 2900 1636
rect 2456 1615 2458 1635
rect 2544 1615 2546 1635
rect 2632 1615 2634 1635
rect 2720 1615 2722 1635
rect 2808 1615 2810 1635
rect 2896 1615 2898 1635
rect 3464 1615 3466 1638
rect 2455 1614 2459 1615
rect 2455 1609 2459 1610
rect 2463 1614 2467 1615
rect 2463 1609 2467 1610
rect 2543 1614 2547 1615
rect 2543 1609 2547 1610
rect 2567 1614 2571 1615
rect 2567 1609 2571 1610
rect 2631 1614 2635 1615
rect 2631 1609 2635 1610
rect 2671 1614 2675 1615
rect 2671 1609 2675 1610
rect 2719 1614 2723 1615
rect 2719 1609 2723 1610
rect 2775 1614 2779 1615
rect 2775 1609 2779 1610
rect 2807 1614 2811 1615
rect 2807 1609 2811 1610
rect 2887 1614 2891 1615
rect 2887 1609 2891 1610
rect 2895 1614 2899 1615
rect 2895 1609 2899 1610
rect 3463 1614 3467 1615
rect 3463 1609 3467 1610
rect 2464 1593 2466 1609
rect 2568 1593 2570 1609
rect 2618 1607 2624 1608
rect 2618 1603 2619 1607
rect 2623 1603 2624 1607
rect 2618 1602 2624 1603
rect 2602 1599 2608 1600
rect 2602 1595 2603 1599
rect 2607 1595 2608 1599
rect 2602 1594 2608 1595
rect 2462 1592 2468 1593
rect 2462 1588 2463 1592
rect 2467 1588 2468 1592
rect 2462 1587 2468 1588
rect 2566 1592 2572 1593
rect 2566 1588 2567 1592
rect 2571 1588 2572 1592
rect 2566 1587 2572 1588
rect 1246 1582 1252 1583
rect 2134 1583 2140 1584
rect 904 1560 906 1582
rect 942 1577 948 1578
rect 942 1573 943 1577
rect 947 1573 948 1577
rect 942 1572 948 1573
rect 838 1559 844 1560
rect 838 1555 839 1559
rect 843 1555 844 1559
rect 838 1554 844 1555
rect 902 1559 908 1560
rect 902 1555 903 1559
rect 907 1555 908 1559
rect 902 1554 908 1555
rect 944 1547 946 1572
rect 1016 1560 1018 1582
rect 1054 1577 1060 1578
rect 1054 1573 1055 1577
rect 1059 1573 1060 1577
rect 1054 1572 1060 1573
rect 1014 1559 1020 1560
rect 1014 1555 1015 1559
rect 1019 1555 1020 1559
rect 1014 1554 1020 1555
rect 1056 1547 1058 1572
rect 1128 1560 1130 1582
rect 1166 1577 1172 1578
rect 1166 1573 1167 1577
rect 1171 1573 1172 1577
rect 1166 1572 1172 1573
rect 1126 1559 1132 1560
rect 1126 1555 1127 1559
rect 1131 1555 1132 1559
rect 1126 1554 1132 1555
rect 1168 1547 1170 1572
rect 1240 1560 1242 1582
rect 1238 1559 1244 1560
rect 1238 1555 1239 1559
rect 1243 1555 1244 1559
rect 1238 1554 1244 1555
rect 1248 1548 1250 1582
rect 2134 1579 2135 1583
rect 2139 1579 2140 1583
rect 2134 1578 2140 1579
rect 2230 1583 2236 1584
rect 2230 1579 2231 1583
rect 2235 1579 2236 1583
rect 2230 1578 2236 1579
rect 2326 1583 2332 1584
rect 2326 1579 2327 1583
rect 2331 1579 2332 1583
rect 2326 1578 2332 1579
rect 2430 1583 2436 1584
rect 2430 1579 2431 1583
rect 2435 1579 2436 1583
rect 2430 1578 2436 1579
rect 2446 1583 2452 1584
rect 2446 1579 2447 1583
rect 2451 1579 2452 1583
rect 2446 1578 2452 1579
rect 1278 1577 1284 1578
rect 1278 1573 1279 1577
rect 1283 1573 1284 1577
rect 1278 1572 1284 1573
rect 1766 1576 1772 1577
rect 1766 1572 1767 1576
rect 1771 1572 1772 1576
rect 2062 1573 2068 1574
rect 1246 1547 1252 1548
rect 1280 1547 1282 1572
rect 1766 1571 1772 1572
rect 1806 1572 1812 1573
rect 1768 1547 1770 1571
rect 1806 1568 1807 1572
rect 1811 1568 1812 1572
rect 2062 1569 2063 1573
rect 2067 1569 2068 1573
rect 2062 1568 2068 1569
rect 1806 1567 1812 1568
rect 1808 1551 1810 1567
rect 2064 1551 2066 1568
rect 2136 1556 2138 1578
rect 2158 1573 2164 1574
rect 2158 1569 2159 1573
rect 2163 1569 2164 1573
rect 2158 1568 2164 1569
rect 2110 1555 2116 1556
rect 2110 1551 2111 1555
rect 2115 1554 2116 1555
rect 2134 1555 2140 1556
rect 2115 1552 2122 1554
rect 2115 1551 2116 1552
rect 1807 1550 1811 1551
rect 719 1546 723 1547
rect 719 1541 723 1542
rect 767 1546 771 1547
rect 767 1541 771 1542
rect 831 1546 835 1547
rect 831 1541 835 1542
rect 911 1546 915 1547
rect 911 1541 915 1542
rect 943 1546 947 1547
rect 943 1541 947 1542
rect 1047 1546 1051 1547
rect 1047 1541 1051 1542
rect 1055 1546 1059 1547
rect 1055 1541 1059 1542
rect 1167 1546 1171 1547
rect 1167 1541 1171 1542
rect 1175 1546 1179 1547
rect 1246 1543 1247 1547
rect 1251 1543 1252 1547
rect 1246 1542 1252 1543
rect 1279 1546 1283 1547
rect 1175 1541 1179 1542
rect 1279 1541 1283 1542
rect 1311 1546 1315 1547
rect 1311 1541 1315 1542
rect 1447 1546 1451 1547
rect 1447 1541 1451 1542
rect 1767 1546 1771 1547
rect 1807 1545 1811 1546
rect 1919 1550 1923 1551
rect 1919 1545 1923 1546
rect 2039 1550 2043 1551
rect 2039 1545 2043 1546
rect 2063 1550 2067 1551
rect 2110 1550 2116 1551
rect 2063 1545 2067 1546
rect 1767 1541 1771 1542
rect 702 1539 708 1540
rect 702 1535 703 1539
rect 707 1535 708 1539
rect 702 1534 708 1535
rect 704 1516 706 1534
rect 768 1524 770 1541
rect 846 1539 852 1540
rect 846 1535 847 1539
rect 851 1535 852 1539
rect 846 1534 852 1535
rect 766 1523 772 1524
rect 766 1519 767 1523
rect 771 1519 772 1523
rect 766 1518 772 1519
rect 290 1515 296 1516
rect 254 1511 260 1512
rect 110 1507 116 1508
rect 110 1503 111 1507
rect 115 1503 116 1507
rect 254 1507 255 1511
rect 259 1507 260 1511
rect 290 1511 291 1515
rect 295 1511 296 1515
rect 290 1510 296 1511
rect 406 1515 412 1516
rect 406 1511 407 1515
rect 411 1511 412 1515
rect 406 1510 412 1511
rect 694 1515 700 1516
rect 694 1511 695 1515
rect 699 1511 700 1515
rect 694 1510 700 1511
rect 702 1515 708 1516
rect 702 1511 703 1515
rect 707 1511 708 1515
rect 702 1510 708 1511
rect 254 1506 260 1507
rect 110 1502 116 1503
rect 182 1504 188 1505
rect 112 1479 114 1502
rect 182 1500 183 1504
rect 187 1500 188 1504
rect 182 1499 188 1500
rect 184 1479 186 1499
rect 111 1478 115 1479
rect 111 1473 115 1474
rect 159 1478 163 1479
rect 159 1473 163 1474
rect 183 1478 187 1479
rect 183 1473 187 1474
rect 112 1454 114 1473
rect 160 1457 162 1473
rect 158 1456 164 1457
rect 110 1453 116 1454
rect 110 1449 111 1453
rect 115 1449 116 1453
rect 158 1452 159 1456
rect 163 1452 164 1456
rect 158 1451 164 1452
rect 110 1448 116 1449
rect 158 1437 164 1438
rect 110 1436 116 1437
rect 110 1432 111 1436
rect 115 1432 116 1436
rect 158 1433 159 1437
rect 163 1433 164 1437
rect 158 1432 164 1433
rect 110 1431 116 1432
rect 112 1411 114 1431
rect 160 1411 162 1432
rect 256 1420 258 1506
rect 326 1504 332 1505
rect 326 1500 327 1504
rect 331 1500 332 1504
rect 326 1499 332 1500
rect 470 1504 476 1505
rect 470 1500 471 1504
rect 475 1500 476 1504
rect 470 1499 476 1500
rect 622 1504 628 1505
rect 622 1500 623 1504
rect 627 1500 628 1504
rect 622 1499 628 1500
rect 766 1504 772 1505
rect 766 1500 767 1504
rect 771 1500 772 1504
rect 766 1499 772 1500
rect 328 1479 330 1499
rect 472 1479 474 1499
rect 624 1479 626 1499
rect 768 1479 770 1499
rect 327 1478 331 1479
rect 327 1473 331 1474
rect 375 1478 379 1479
rect 375 1473 379 1474
rect 471 1478 475 1479
rect 471 1473 475 1474
rect 583 1478 587 1479
rect 583 1473 587 1474
rect 623 1478 627 1479
rect 623 1473 627 1474
rect 767 1478 771 1479
rect 767 1473 771 1474
rect 783 1478 787 1479
rect 783 1473 787 1474
rect 376 1457 378 1473
rect 584 1457 586 1473
rect 784 1457 786 1473
rect 374 1456 380 1457
rect 374 1452 375 1456
rect 379 1452 380 1456
rect 374 1451 380 1452
rect 582 1456 588 1457
rect 582 1452 583 1456
rect 587 1452 588 1456
rect 582 1451 588 1452
rect 782 1456 788 1457
rect 782 1452 783 1456
rect 787 1452 788 1456
rect 782 1451 788 1452
rect 848 1448 850 1534
rect 912 1524 914 1541
rect 1048 1524 1050 1541
rect 1118 1539 1124 1540
rect 1118 1535 1119 1539
rect 1123 1535 1124 1539
rect 1118 1534 1124 1535
rect 910 1523 916 1524
rect 910 1519 911 1523
rect 915 1519 916 1523
rect 910 1518 916 1519
rect 1046 1523 1052 1524
rect 1046 1519 1047 1523
rect 1051 1519 1052 1523
rect 1046 1518 1052 1519
rect 1120 1516 1122 1534
rect 1176 1524 1178 1541
rect 1246 1539 1252 1540
rect 1246 1535 1247 1539
rect 1251 1535 1252 1539
rect 1246 1534 1252 1535
rect 1174 1523 1180 1524
rect 1174 1519 1175 1523
rect 1179 1519 1180 1523
rect 1174 1518 1180 1519
rect 1248 1516 1250 1534
rect 1312 1524 1314 1541
rect 1382 1539 1388 1540
rect 1382 1535 1383 1539
rect 1387 1535 1388 1539
rect 1382 1534 1388 1535
rect 1310 1523 1316 1524
rect 1310 1519 1311 1523
rect 1315 1519 1316 1523
rect 1310 1518 1316 1519
rect 1384 1516 1386 1534
rect 1448 1524 1450 1541
rect 1768 1525 1770 1541
rect 1808 1529 1810 1545
rect 1806 1528 1812 1529
rect 1920 1528 1922 1545
rect 1982 1543 1988 1544
rect 1982 1539 1983 1543
rect 1987 1539 1988 1543
rect 1982 1538 1988 1539
rect 1990 1543 1996 1544
rect 1990 1539 1991 1543
rect 1995 1539 1996 1543
rect 1990 1538 1996 1539
rect 1766 1524 1772 1525
rect 1446 1523 1452 1524
rect 1446 1519 1447 1523
rect 1451 1519 1452 1523
rect 1766 1520 1767 1524
rect 1771 1520 1772 1524
rect 1806 1524 1807 1528
rect 1811 1524 1812 1528
rect 1806 1523 1812 1524
rect 1918 1527 1924 1528
rect 1918 1523 1919 1527
rect 1923 1523 1924 1527
rect 1918 1522 1924 1523
rect 1766 1519 1772 1520
rect 1446 1518 1452 1519
rect 1118 1515 1124 1516
rect 1118 1511 1119 1515
rect 1123 1511 1124 1515
rect 1118 1510 1124 1511
rect 1246 1515 1252 1516
rect 1246 1511 1247 1515
rect 1251 1511 1252 1515
rect 1246 1510 1252 1511
rect 1382 1515 1388 1516
rect 1382 1511 1383 1515
rect 1387 1511 1388 1515
rect 1382 1510 1388 1511
rect 1398 1515 1404 1516
rect 1398 1511 1399 1515
rect 1403 1511 1404 1515
rect 1398 1510 1404 1511
rect 1806 1511 1812 1512
rect 910 1504 916 1505
rect 910 1500 911 1504
rect 915 1500 916 1504
rect 910 1499 916 1500
rect 1046 1504 1052 1505
rect 1046 1500 1047 1504
rect 1051 1500 1052 1504
rect 1046 1499 1052 1500
rect 1174 1504 1180 1505
rect 1174 1500 1175 1504
rect 1179 1500 1180 1504
rect 1174 1499 1180 1500
rect 1310 1504 1316 1505
rect 1310 1500 1311 1504
rect 1315 1500 1316 1504
rect 1310 1499 1316 1500
rect 912 1479 914 1499
rect 1048 1479 1050 1499
rect 1176 1479 1178 1499
rect 1312 1479 1314 1499
rect 911 1478 915 1479
rect 911 1473 915 1474
rect 959 1478 963 1479
rect 959 1473 963 1474
rect 1047 1478 1051 1479
rect 1047 1473 1051 1474
rect 1127 1478 1131 1479
rect 1127 1473 1131 1474
rect 1175 1478 1179 1479
rect 1175 1473 1179 1474
rect 1279 1478 1283 1479
rect 1279 1473 1283 1474
rect 1311 1478 1315 1479
rect 1311 1473 1315 1474
rect 960 1457 962 1473
rect 1066 1463 1072 1464
rect 1066 1459 1067 1463
rect 1071 1459 1072 1463
rect 1066 1458 1072 1459
rect 958 1456 964 1457
rect 958 1452 959 1456
rect 963 1452 964 1456
rect 958 1451 964 1452
rect 262 1447 268 1448
rect 262 1443 263 1447
rect 267 1443 268 1447
rect 262 1442 268 1443
rect 446 1447 452 1448
rect 446 1443 447 1447
rect 451 1443 452 1447
rect 446 1442 452 1443
rect 654 1447 660 1448
rect 654 1443 655 1447
rect 659 1443 660 1447
rect 654 1442 660 1443
rect 846 1447 852 1448
rect 846 1443 847 1447
rect 851 1443 852 1447
rect 846 1442 852 1443
rect 264 1420 266 1442
rect 374 1437 380 1438
rect 374 1433 375 1437
rect 379 1433 380 1437
rect 374 1432 380 1433
rect 254 1419 260 1420
rect 254 1415 255 1419
rect 259 1415 260 1419
rect 254 1414 260 1415
rect 262 1419 268 1420
rect 262 1415 263 1419
rect 267 1415 268 1419
rect 262 1414 268 1415
rect 376 1411 378 1432
rect 111 1410 115 1411
rect 111 1405 115 1406
rect 135 1410 139 1411
rect 135 1405 139 1406
rect 159 1410 163 1411
rect 159 1405 163 1406
rect 303 1410 307 1411
rect 303 1405 307 1406
rect 375 1410 379 1411
rect 375 1405 379 1406
rect 112 1389 114 1405
rect 110 1388 116 1389
rect 136 1388 138 1405
rect 282 1403 288 1404
rect 282 1399 283 1403
rect 287 1399 288 1403
rect 282 1398 288 1399
rect 110 1384 111 1388
rect 115 1384 116 1388
rect 110 1383 116 1384
rect 134 1387 140 1388
rect 134 1383 135 1387
rect 139 1383 140 1387
rect 134 1382 140 1383
rect 284 1380 286 1398
rect 304 1388 306 1405
rect 448 1404 450 1442
rect 582 1437 588 1438
rect 582 1433 583 1437
rect 587 1433 588 1437
rect 582 1432 588 1433
rect 584 1411 586 1432
rect 656 1420 658 1442
rect 782 1437 788 1438
rect 782 1433 783 1437
rect 787 1433 788 1437
rect 782 1432 788 1433
rect 958 1437 964 1438
rect 958 1433 959 1437
rect 963 1433 964 1437
rect 958 1432 964 1433
rect 634 1419 640 1420
rect 634 1415 635 1419
rect 639 1415 640 1419
rect 634 1414 640 1415
rect 654 1419 660 1420
rect 654 1415 655 1419
rect 659 1415 660 1419
rect 654 1414 660 1415
rect 495 1410 499 1411
rect 495 1405 499 1406
rect 583 1410 587 1411
rect 583 1405 587 1406
rect 446 1403 452 1404
rect 446 1399 447 1403
rect 451 1399 452 1403
rect 446 1398 452 1399
rect 496 1388 498 1405
rect 302 1387 308 1388
rect 302 1383 303 1387
rect 307 1383 308 1387
rect 302 1382 308 1383
rect 494 1387 500 1388
rect 494 1383 495 1387
rect 499 1383 500 1387
rect 494 1382 500 1383
rect 636 1380 638 1414
rect 784 1411 786 1432
rect 960 1411 962 1432
rect 679 1410 683 1411
rect 679 1405 683 1406
rect 783 1410 787 1411
rect 783 1405 787 1406
rect 855 1410 859 1411
rect 855 1405 859 1406
rect 959 1410 963 1411
rect 959 1405 963 1406
rect 1015 1410 1019 1411
rect 1015 1405 1019 1406
rect 680 1388 682 1405
rect 758 1403 764 1404
rect 758 1399 759 1403
rect 763 1399 764 1403
rect 758 1398 764 1399
rect 678 1387 684 1388
rect 678 1383 679 1387
rect 683 1383 684 1387
rect 678 1382 684 1383
rect 760 1380 762 1398
rect 856 1388 858 1405
rect 974 1403 980 1404
rect 974 1399 975 1403
rect 979 1399 980 1403
rect 974 1398 980 1399
rect 854 1387 860 1388
rect 854 1383 855 1387
rect 859 1383 860 1387
rect 854 1382 860 1383
rect 282 1379 288 1380
rect 282 1375 283 1379
rect 287 1375 288 1379
rect 282 1374 288 1375
rect 634 1379 640 1380
rect 634 1375 635 1379
rect 639 1375 640 1379
rect 634 1374 640 1375
rect 758 1379 764 1380
rect 758 1375 759 1379
rect 763 1375 764 1379
rect 758 1374 764 1375
rect 110 1371 116 1372
rect 110 1367 111 1371
rect 115 1367 116 1371
rect 198 1371 204 1372
rect 110 1366 116 1367
rect 134 1368 140 1369
rect 112 1343 114 1366
rect 134 1364 135 1368
rect 139 1364 140 1368
rect 198 1367 199 1371
rect 203 1367 204 1371
rect 198 1366 204 1367
rect 302 1368 308 1369
rect 134 1363 140 1364
rect 136 1343 138 1363
rect 111 1342 115 1343
rect 111 1337 115 1338
rect 135 1342 139 1343
rect 135 1337 139 1338
rect 112 1318 114 1337
rect 136 1321 138 1337
rect 134 1320 140 1321
rect 110 1317 116 1318
rect 110 1313 111 1317
rect 115 1313 116 1317
rect 134 1316 135 1320
rect 139 1316 140 1320
rect 134 1315 140 1316
rect 110 1312 116 1313
rect 134 1301 140 1302
rect 110 1300 116 1301
rect 110 1296 111 1300
rect 115 1296 116 1300
rect 134 1297 135 1301
rect 139 1297 140 1301
rect 134 1296 140 1297
rect 110 1295 116 1296
rect 112 1275 114 1295
rect 136 1275 138 1296
rect 187 1284 191 1285
rect 200 1284 202 1366
rect 302 1364 303 1368
rect 307 1364 308 1368
rect 302 1363 308 1364
rect 494 1368 500 1369
rect 494 1364 495 1368
rect 499 1364 500 1368
rect 494 1363 500 1364
rect 678 1368 684 1369
rect 678 1364 679 1368
rect 683 1364 684 1368
rect 678 1363 684 1364
rect 854 1368 860 1369
rect 854 1364 855 1368
rect 859 1364 860 1368
rect 854 1363 860 1364
rect 304 1343 306 1363
rect 496 1343 498 1363
rect 680 1343 682 1363
rect 856 1343 858 1363
rect 247 1342 251 1343
rect 247 1337 251 1338
rect 303 1342 307 1343
rect 303 1337 307 1338
rect 399 1342 403 1343
rect 399 1337 403 1338
rect 495 1342 499 1343
rect 495 1337 499 1338
rect 559 1342 563 1343
rect 559 1337 563 1338
rect 679 1342 683 1343
rect 679 1337 683 1338
rect 727 1342 731 1343
rect 727 1337 731 1338
rect 855 1342 859 1343
rect 855 1337 859 1338
rect 895 1342 899 1343
rect 895 1337 899 1338
rect 248 1321 250 1337
rect 400 1321 402 1337
rect 560 1321 562 1337
rect 728 1321 730 1337
rect 896 1321 898 1337
rect 246 1320 252 1321
rect 246 1316 247 1320
rect 251 1316 252 1320
rect 246 1315 252 1316
rect 398 1320 404 1321
rect 398 1316 399 1320
rect 403 1316 404 1320
rect 398 1315 404 1316
rect 558 1320 564 1321
rect 558 1316 559 1320
rect 563 1316 564 1320
rect 558 1315 564 1316
rect 726 1320 732 1321
rect 726 1316 727 1320
rect 731 1316 732 1320
rect 726 1315 732 1316
rect 894 1320 900 1321
rect 894 1316 895 1320
rect 899 1316 900 1320
rect 894 1315 900 1316
rect 976 1312 978 1398
rect 1016 1388 1018 1405
rect 1068 1404 1070 1458
rect 1128 1457 1130 1473
rect 1280 1457 1282 1473
rect 1126 1456 1132 1457
rect 1126 1452 1127 1456
rect 1131 1452 1132 1456
rect 1126 1451 1132 1452
rect 1278 1456 1284 1457
rect 1278 1452 1279 1456
rect 1283 1452 1284 1456
rect 1278 1451 1284 1452
rect 1090 1447 1096 1448
rect 1090 1443 1091 1447
rect 1095 1443 1096 1447
rect 1090 1442 1096 1443
rect 1198 1447 1204 1448
rect 1198 1443 1199 1447
rect 1203 1443 1204 1447
rect 1198 1442 1204 1443
rect 1350 1447 1356 1448
rect 1350 1443 1351 1447
rect 1355 1443 1356 1447
rect 1350 1442 1356 1443
rect 1092 1420 1094 1442
rect 1126 1437 1132 1438
rect 1126 1433 1127 1437
rect 1131 1433 1132 1437
rect 1126 1432 1132 1433
rect 1090 1419 1096 1420
rect 1090 1415 1091 1419
rect 1095 1415 1096 1419
rect 1090 1414 1096 1415
rect 1128 1411 1130 1432
rect 1200 1420 1202 1442
rect 1278 1437 1284 1438
rect 1278 1433 1279 1437
rect 1283 1433 1284 1437
rect 1278 1432 1284 1433
rect 1198 1419 1204 1420
rect 1198 1415 1199 1419
rect 1203 1415 1204 1419
rect 1198 1414 1204 1415
rect 1280 1411 1282 1432
rect 1352 1420 1354 1442
rect 1350 1419 1356 1420
rect 1350 1415 1351 1419
rect 1355 1415 1356 1419
rect 1350 1414 1356 1415
rect 1400 1412 1402 1510
rect 1766 1507 1772 1508
rect 1446 1504 1452 1505
rect 1446 1500 1447 1504
rect 1451 1500 1452 1504
rect 1766 1503 1767 1507
rect 1771 1503 1772 1507
rect 1806 1507 1807 1511
rect 1811 1507 1812 1511
rect 1806 1506 1812 1507
rect 1918 1508 1924 1509
rect 1766 1502 1772 1503
rect 1446 1499 1452 1500
rect 1448 1479 1450 1499
rect 1768 1479 1770 1502
rect 1808 1479 1810 1506
rect 1918 1504 1919 1508
rect 1923 1504 1924 1508
rect 1918 1503 1924 1504
rect 1920 1479 1922 1503
rect 1431 1478 1435 1479
rect 1431 1473 1435 1474
rect 1447 1478 1451 1479
rect 1447 1473 1451 1474
rect 1591 1478 1595 1479
rect 1591 1473 1595 1474
rect 1767 1478 1771 1479
rect 1767 1473 1771 1474
rect 1807 1478 1811 1479
rect 1807 1473 1811 1474
rect 1831 1478 1835 1479
rect 1831 1473 1835 1474
rect 1919 1478 1923 1479
rect 1919 1473 1923 1474
rect 1951 1478 1955 1479
rect 1951 1473 1955 1474
rect 1432 1457 1434 1473
rect 1592 1457 1594 1473
rect 1430 1456 1436 1457
rect 1430 1452 1431 1456
rect 1435 1452 1436 1456
rect 1430 1451 1436 1452
rect 1590 1456 1596 1457
rect 1590 1452 1591 1456
rect 1595 1452 1596 1456
rect 1768 1454 1770 1473
rect 1808 1454 1810 1473
rect 1832 1457 1834 1473
rect 1952 1457 1954 1473
rect 1984 1464 1986 1538
rect 1992 1520 1994 1538
rect 2040 1528 2042 1545
rect 2110 1543 2116 1544
rect 2110 1539 2111 1543
rect 2115 1539 2116 1543
rect 2110 1538 2116 1539
rect 2038 1527 2044 1528
rect 2038 1523 2039 1527
rect 2043 1523 2044 1527
rect 2038 1522 2044 1523
rect 2112 1520 2114 1538
rect 1990 1519 1996 1520
rect 1990 1515 1991 1519
rect 1995 1515 1996 1519
rect 1990 1514 1996 1515
rect 2110 1519 2116 1520
rect 2110 1515 2111 1519
rect 2115 1515 2116 1519
rect 2110 1514 2116 1515
rect 2038 1508 2044 1509
rect 2038 1504 2039 1508
rect 2043 1504 2044 1508
rect 2038 1503 2044 1504
rect 2040 1479 2042 1503
rect 2120 1500 2122 1552
rect 2134 1551 2135 1555
rect 2139 1551 2140 1555
rect 2160 1551 2162 1568
rect 2232 1556 2234 1578
rect 2254 1573 2260 1574
rect 2254 1569 2255 1573
rect 2259 1569 2260 1573
rect 2254 1568 2260 1569
rect 2230 1555 2236 1556
rect 2230 1551 2231 1555
rect 2235 1551 2236 1555
rect 2256 1551 2258 1568
rect 2328 1556 2330 1578
rect 2358 1573 2364 1574
rect 2358 1569 2359 1573
rect 2363 1569 2364 1573
rect 2358 1568 2364 1569
rect 2326 1555 2332 1556
rect 2326 1551 2327 1555
rect 2331 1551 2332 1555
rect 2360 1551 2362 1568
rect 2432 1556 2434 1578
rect 2462 1573 2468 1574
rect 2462 1569 2463 1573
rect 2467 1569 2468 1573
rect 2462 1568 2468 1569
rect 2566 1573 2572 1574
rect 2566 1569 2567 1573
rect 2571 1569 2572 1573
rect 2566 1568 2572 1569
rect 2430 1555 2436 1556
rect 2430 1551 2431 1555
rect 2435 1551 2436 1555
rect 2464 1551 2466 1568
rect 2568 1551 2570 1568
rect 2134 1550 2140 1551
rect 2159 1550 2163 1551
rect 2159 1545 2163 1546
rect 2167 1550 2171 1551
rect 2230 1550 2236 1551
rect 2255 1550 2259 1551
rect 2167 1545 2171 1546
rect 2255 1545 2259 1546
rect 2295 1550 2299 1551
rect 2326 1550 2332 1551
rect 2359 1550 2363 1551
rect 2295 1545 2299 1546
rect 2359 1545 2363 1546
rect 2423 1550 2427 1551
rect 2430 1550 2436 1551
rect 2463 1550 2467 1551
rect 2423 1545 2427 1546
rect 2463 1545 2467 1546
rect 2551 1550 2555 1551
rect 2551 1545 2555 1546
rect 2567 1550 2571 1551
rect 2567 1545 2571 1546
rect 2168 1528 2170 1545
rect 2238 1543 2244 1544
rect 2238 1539 2239 1543
rect 2243 1539 2244 1543
rect 2238 1538 2244 1539
rect 2166 1527 2172 1528
rect 2166 1523 2167 1527
rect 2171 1523 2172 1527
rect 2166 1522 2172 1523
rect 2240 1520 2242 1538
rect 2296 1528 2298 1545
rect 2366 1543 2372 1544
rect 2366 1539 2367 1543
rect 2371 1539 2372 1543
rect 2366 1538 2372 1539
rect 2294 1527 2300 1528
rect 2294 1523 2295 1527
rect 2299 1523 2300 1527
rect 2294 1522 2300 1523
rect 2368 1520 2370 1538
rect 2424 1528 2426 1545
rect 2552 1528 2554 1545
rect 2604 1544 2606 1594
rect 2620 1556 2622 1602
rect 2672 1593 2674 1609
rect 2776 1593 2778 1609
rect 2888 1593 2890 1609
rect 2670 1592 2676 1593
rect 2670 1588 2671 1592
rect 2675 1588 2676 1592
rect 2670 1587 2676 1588
rect 2774 1592 2780 1593
rect 2774 1588 2775 1592
rect 2779 1588 2780 1592
rect 2774 1587 2780 1588
rect 2886 1592 2892 1593
rect 2886 1588 2887 1592
rect 2891 1588 2892 1592
rect 3464 1590 3466 1609
rect 2886 1587 2892 1588
rect 3462 1589 3468 1590
rect 3462 1585 3463 1589
rect 3467 1585 3468 1589
rect 3462 1584 3468 1585
rect 2638 1583 2644 1584
rect 2638 1579 2639 1583
rect 2643 1579 2644 1583
rect 2638 1578 2644 1579
rect 2742 1583 2748 1584
rect 2742 1579 2743 1583
rect 2747 1579 2748 1583
rect 2742 1578 2748 1579
rect 2846 1583 2852 1584
rect 2846 1579 2847 1583
rect 2851 1579 2852 1583
rect 2846 1578 2852 1579
rect 2640 1556 2642 1578
rect 2670 1573 2676 1574
rect 2670 1569 2671 1573
rect 2675 1569 2676 1573
rect 2670 1568 2676 1569
rect 2618 1555 2624 1556
rect 2618 1551 2619 1555
rect 2623 1551 2624 1555
rect 2618 1550 2624 1551
rect 2638 1555 2644 1556
rect 2638 1551 2639 1555
rect 2643 1551 2644 1555
rect 2672 1551 2674 1568
rect 2744 1556 2746 1578
rect 2774 1573 2780 1574
rect 2774 1569 2775 1573
rect 2779 1569 2780 1573
rect 2774 1568 2780 1569
rect 2742 1555 2748 1556
rect 2742 1551 2743 1555
rect 2747 1551 2748 1555
rect 2776 1551 2778 1568
rect 2848 1556 2850 1578
rect 2886 1573 2892 1574
rect 2886 1569 2887 1573
rect 2891 1569 2892 1573
rect 2886 1568 2892 1569
rect 3462 1572 3468 1573
rect 3462 1568 3463 1572
rect 3467 1568 3468 1572
rect 2846 1555 2852 1556
rect 2846 1551 2847 1555
rect 2851 1551 2852 1555
rect 2888 1551 2890 1568
rect 3462 1567 3468 1568
rect 3464 1551 3466 1567
rect 2638 1550 2644 1551
rect 2671 1550 2675 1551
rect 2671 1545 2675 1546
rect 2679 1550 2683 1551
rect 2742 1550 2748 1551
rect 2775 1550 2779 1551
rect 2679 1545 2683 1546
rect 2775 1545 2779 1546
rect 2799 1550 2803 1551
rect 2846 1550 2852 1551
rect 2887 1550 2891 1551
rect 2799 1545 2803 1546
rect 2887 1545 2891 1546
rect 2927 1550 2931 1551
rect 2927 1545 2931 1546
rect 3055 1550 3059 1551
rect 3055 1545 3059 1546
rect 3463 1550 3467 1551
rect 3463 1545 3467 1546
rect 2602 1543 2608 1544
rect 2602 1539 2603 1543
rect 2607 1539 2608 1543
rect 2602 1538 2608 1539
rect 2622 1543 2628 1544
rect 2622 1539 2623 1543
rect 2627 1539 2628 1543
rect 2622 1538 2628 1539
rect 2422 1527 2428 1528
rect 2422 1523 2423 1527
rect 2427 1523 2428 1527
rect 2422 1522 2428 1523
rect 2550 1527 2556 1528
rect 2550 1523 2551 1527
rect 2555 1523 2556 1527
rect 2550 1522 2556 1523
rect 2624 1520 2626 1538
rect 2680 1528 2682 1545
rect 2750 1543 2756 1544
rect 2750 1539 2751 1543
rect 2755 1539 2756 1543
rect 2750 1538 2756 1539
rect 2678 1527 2684 1528
rect 2678 1523 2679 1527
rect 2683 1523 2684 1527
rect 2678 1522 2684 1523
rect 2752 1520 2754 1538
rect 2800 1528 2802 1545
rect 2870 1543 2876 1544
rect 2870 1539 2871 1543
rect 2875 1539 2876 1543
rect 2870 1538 2876 1539
rect 2798 1527 2804 1528
rect 2798 1523 2799 1527
rect 2803 1523 2804 1527
rect 2798 1522 2804 1523
rect 2872 1520 2874 1538
rect 2928 1528 2930 1545
rect 2998 1543 3004 1544
rect 2998 1539 2999 1543
rect 3003 1539 3004 1543
rect 2998 1538 3004 1539
rect 2926 1527 2932 1528
rect 2926 1523 2927 1527
rect 2931 1523 2932 1527
rect 2926 1522 2932 1523
rect 3000 1520 3002 1538
rect 3056 1528 3058 1545
rect 3464 1529 3466 1545
rect 3462 1528 3468 1529
rect 3054 1527 3060 1528
rect 3054 1523 3055 1527
rect 3059 1523 3060 1527
rect 3462 1524 3463 1528
rect 3467 1524 3468 1528
rect 3462 1523 3468 1524
rect 3054 1522 3060 1523
rect 2238 1519 2244 1520
rect 2238 1515 2239 1519
rect 2243 1515 2244 1519
rect 2238 1514 2244 1515
rect 2366 1519 2372 1520
rect 2366 1515 2367 1519
rect 2371 1515 2372 1519
rect 2366 1514 2372 1515
rect 2374 1519 2380 1520
rect 2374 1515 2375 1519
rect 2379 1515 2380 1519
rect 2374 1514 2380 1515
rect 2622 1519 2628 1520
rect 2622 1515 2623 1519
rect 2627 1515 2628 1519
rect 2622 1514 2628 1515
rect 2750 1519 2756 1520
rect 2750 1515 2751 1519
rect 2755 1515 2756 1519
rect 2750 1514 2756 1515
rect 2870 1519 2876 1520
rect 2870 1515 2871 1519
rect 2875 1515 2876 1519
rect 2870 1514 2876 1515
rect 2998 1519 3004 1520
rect 2998 1515 2999 1519
rect 3003 1515 3004 1519
rect 2998 1514 3004 1515
rect 3018 1519 3024 1520
rect 3018 1515 3019 1519
rect 3023 1515 3024 1519
rect 3018 1514 3024 1515
rect 2166 1508 2172 1509
rect 2166 1504 2167 1508
rect 2171 1504 2172 1508
rect 2166 1503 2172 1504
rect 2294 1508 2300 1509
rect 2294 1504 2295 1508
rect 2299 1504 2300 1508
rect 2294 1503 2300 1504
rect 2118 1499 2124 1500
rect 2118 1495 2119 1499
rect 2123 1495 2124 1499
rect 2118 1494 2124 1495
rect 2168 1479 2170 1503
rect 2296 1479 2298 1503
rect 2376 1500 2378 1514
rect 2422 1508 2428 1509
rect 2422 1504 2423 1508
rect 2427 1504 2428 1508
rect 2422 1503 2428 1504
rect 2550 1508 2556 1509
rect 2550 1504 2551 1508
rect 2555 1504 2556 1508
rect 2550 1503 2556 1504
rect 2678 1508 2684 1509
rect 2678 1504 2679 1508
rect 2683 1504 2684 1508
rect 2678 1503 2684 1504
rect 2798 1508 2804 1509
rect 2798 1504 2799 1508
rect 2803 1504 2804 1508
rect 2798 1503 2804 1504
rect 2926 1508 2932 1509
rect 2926 1504 2927 1508
rect 2931 1504 2932 1508
rect 2926 1503 2932 1504
rect 2374 1499 2380 1500
rect 2374 1495 2375 1499
rect 2379 1495 2380 1499
rect 2374 1494 2380 1495
rect 2424 1479 2426 1503
rect 2552 1479 2554 1503
rect 2680 1479 2682 1503
rect 2800 1479 2802 1503
rect 2928 1479 2930 1503
rect 2039 1478 2043 1479
rect 2039 1473 2043 1474
rect 2111 1478 2115 1479
rect 2111 1473 2115 1474
rect 2167 1478 2171 1479
rect 2167 1473 2171 1474
rect 2271 1478 2275 1479
rect 2271 1473 2275 1474
rect 2295 1478 2299 1479
rect 2295 1473 2299 1474
rect 2423 1478 2427 1479
rect 2423 1473 2427 1474
rect 2431 1478 2435 1479
rect 2431 1473 2435 1474
rect 2551 1478 2555 1479
rect 2551 1473 2555 1474
rect 2591 1478 2595 1479
rect 2591 1473 2595 1474
rect 2679 1478 2683 1479
rect 2679 1473 2683 1474
rect 2735 1478 2739 1479
rect 2735 1473 2739 1474
rect 2799 1478 2803 1479
rect 2799 1473 2803 1474
rect 2871 1478 2875 1479
rect 2871 1473 2875 1474
rect 2927 1478 2931 1479
rect 2927 1473 2931 1474
rect 3007 1478 3011 1479
rect 3007 1473 3011 1474
rect 1982 1463 1988 1464
rect 1982 1459 1983 1463
rect 1987 1459 1988 1463
rect 1982 1458 1988 1459
rect 2112 1457 2114 1473
rect 2272 1457 2274 1473
rect 2432 1457 2434 1473
rect 2592 1457 2594 1473
rect 2610 1463 2616 1464
rect 2610 1459 2611 1463
rect 2615 1459 2616 1463
rect 2610 1458 2616 1459
rect 1830 1456 1836 1457
rect 1590 1451 1596 1452
rect 1766 1453 1772 1454
rect 1766 1449 1767 1453
rect 1771 1449 1772 1453
rect 1766 1448 1772 1449
rect 1806 1453 1812 1454
rect 1806 1449 1807 1453
rect 1811 1449 1812 1453
rect 1830 1452 1831 1456
rect 1835 1452 1836 1456
rect 1830 1451 1836 1452
rect 1950 1456 1956 1457
rect 1950 1452 1951 1456
rect 1955 1452 1956 1456
rect 1950 1451 1956 1452
rect 2110 1456 2116 1457
rect 2110 1452 2111 1456
rect 2115 1452 2116 1456
rect 2110 1451 2116 1452
rect 2270 1456 2276 1457
rect 2270 1452 2271 1456
rect 2275 1452 2276 1456
rect 2270 1451 2276 1452
rect 2430 1456 2436 1457
rect 2430 1452 2431 1456
rect 2435 1452 2436 1456
rect 2430 1451 2436 1452
rect 2590 1456 2596 1457
rect 2590 1452 2591 1456
rect 2595 1452 2596 1456
rect 2590 1451 2596 1452
rect 1806 1448 1812 1449
rect 1502 1447 1508 1448
rect 1502 1443 1503 1447
rect 1507 1443 1508 1447
rect 1502 1442 1508 1443
rect 2022 1447 2028 1448
rect 2022 1443 2023 1447
rect 2027 1443 2028 1447
rect 2022 1442 2028 1443
rect 2182 1447 2188 1448
rect 2182 1443 2183 1447
rect 2187 1443 2188 1447
rect 2182 1442 2188 1443
rect 2342 1447 2348 1448
rect 2342 1443 2343 1447
rect 2347 1443 2348 1447
rect 2342 1442 2348 1443
rect 1430 1437 1436 1438
rect 1430 1433 1431 1437
rect 1435 1433 1436 1437
rect 1430 1432 1436 1433
rect 1398 1411 1404 1412
rect 1432 1411 1434 1432
rect 1504 1420 1506 1442
rect 1590 1437 1596 1438
rect 1830 1437 1836 1438
rect 1590 1433 1591 1437
rect 1595 1433 1596 1437
rect 1590 1432 1596 1433
rect 1766 1436 1772 1437
rect 1766 1432 1767 1436
rect 1771 1432 1772 1436
rect 1502 1419 1508 1420
rect 1502 1415 1503 1419
rect 1507 1415 1508 1419
rect 1502 1414 1508 1415
rect 1592 1411 1594 1432
rect 1766 1431 1772 1432
rect 1806 1436 1812 1437
rect 1806 1432 1807 1436
rect 1811 1432 1812 1436
rect 1830 1433 1831 1437
rect 1835 1433 1836 1437
rect 1830 1432 1836 1433
rect 1950 1437 1956 1438
rect 1950 1433 1951 1437
rect 1955 1433 1956 1437
rect 1950 1432 1956 1433
rect 1806 1431 1812 1432
rect 1742 1411 1748 1412
rect 1768 1411 1770 1431
rect 1808 1411 1810 1431
rect 1832 1411 1834 1432
rect 1952 1411 1954 1432
rect 2024 1420 2026 1442
rect 2110 1437 2116 1438
rect 2110 1433 2111 1437
rect 2115 1433 2116 1437
rect 2110 1432 2116 1433
rect 2022 1419 2028 1420
rect 2022 1415 2023 1419
rect 2027 1415 2028 1419
rect 2022 1414 2028 1415
rect 2112 1411 2114 1432
rect 2184 1420 2186 1442
rect 2270 1437 2276 1438
rect 2270 1433 2271 1437
rect 2275 1433 2276 1437
rect 2270 1432 2276 1433
rect 2182 1419 2188 1420
rect 2182 1415 2183 1419
rect 2187 1415 2188 1419
rect 2182 1414 2188 1415
rect 2272 1411 2274 1432
rect 2344 1420 2346 1442
rect 2430 1437 2436 1438
rect 2430 1433 2431 1437
rect 2435 1433 2436 1437
rect 2430 1432 2436 1433
rect 2590 1437 2596 1438
rect 2590 1433 2591 1437
rect 2595 1433 2596 1437
rect 2590 1432 2596 1433
rect 2342 1419 2348 1420
rect 2342 1415 2343 1419
rect 2347 1415 2348 1419
rect 2342 1414 2348 1415
rect 2342 1411 2348 1412
rect 2432 1411 2434 1432
rect 2592 1411 2594 1432
rect 1127 1410 1131 1411
rect 1127 1405 1131 1406
rect 1167 1410 1171 1411
rect 1167 1405 1171 1406
rect 1279 1410 1283 1411
rect 1279 1405 1283 1406
rect 1303 1410 1307 1411
rect 1398 1407 1399 1411
rect 1403 1407 1404 1411
rect 1398 1406 1404 1407
rect 1431 1410 1435 1411
rect 1303 1405 1307 1406
rect 1431 1405 1435 1406
rect 1559 1410 1563 1411
rect 1559 1405 1563 1406
rect 1591 1410 1595 1411
rect 1591 1405 1595 1406
rect 1671 1410 1675 1411
rect 1742 1407 1743 1411
rect 1747 1407 1748 1411
rect 1742 1406 1748 1407
rect 1767 1410 1771 1411
rect 1671 1405 1675 1406
rect 1066 1403 1072 1404
rect 1066 1399 1067 1403
rect 1071 1399 1072 1403
rect 1066 1398 1072 1399
rect 1086 1403 1092 1404
rect 1086 1399 1087 1403
rect 1091 1399 1092 1403
rect 1086 1398 1092 1399
rect 1014 1387 1020 1388
rect 1014 1383 1015 1387
rect 1019 1383 1020 1387
rect 1014 1382 1020 1383
rect 1088 1380 1090 1398
rect 1168 1388 1170 1405
rect 1238 1403 1244 1404
rect 1238 1399 1239 1403
rect 1243 1399 1244 1403
rect 1238 1398 1244 1399
rect 1166 1387 1172 1388
rect 1166 1383 1167 1387
rect 1171 1383 1172 1387
rect 1166 1382 1172 1383
rect 1240 1380 1242 1398
rect 1304 1388 1306 1405
rect 1374 1403 1380 1404
rect 1374 1399 1375 1403
rect 1379 1399 1380 1403
rect 1374 1398 1380 1399
rect 1302 1387 1308 1388
rect 1302 1383 1303 1387
rect 1307 1383 1308 1387
rect 1302 1382 1308 1383
rect 1376 1380 1378 1398
rect 1432 1388 1434 1405
rect 1502 1403 1508 1404
rect 1502 1399 1503 1403
rect 1507 1399 1508 1403
rect 1502 1398 1508 1399
rect 1430 1387 1436 1388
rect 1430 1383 1431 1387
rect 1435 1383 1436 1387
rect 1430 1382 1436 1383
rect 1504 1380 1506 1398
rect 1560 1388 1562 1405
rect 1672 1388 1674 1405
rect 1558 1387 1564 1388
rect 1558 1383 1559 1387
rect 1563 1383 1564 1387
rect 1558 1382 1564 1383
rect 1670 1387 1676 1388
rect 1670 1383 1671 1387
rect 1675 1383 1676 1387
rect 1670 1382 1676 1383
rect 1744 1380 1746 1406
rect 1767 1405 1771 1406
rect 1807 1410 1811 1411
rect 1807 1405 1811 1406
rect 1831 1410 1835 1411
rect 1831 1405 1835 1406
rect 1951 1410 1955 1411
rect 1951 1405 1955 1406
rect 2007 1410 2011 1411
rect 2007 1405 2011 1406
rect 2111 1410 2115 1411
rect 2111 1405 2115 1406
rect 2199 1410 2203 1411
rect 2199 1405 2203 1406
rect 2271 1410 2275 1411
rect 2342 1407 2343 1411
rect 2347 1407 2348 1411
rect 2342 1406 2348 1407
rect 2383 1410 2387 1411
rect 2271 1405 2275 1406
rect 1750 1403 1756 1404
rect 1750 1399 1751 1403
rect 1755 1399 1756 1403
rect 1750 1398 1756 1399
rect 1752 1380 1754 1398
rect 1768 1389 1770 1405
rect 1808 1389 1810 1405
rect 1766 1388 1772 1389
rect 1766 1384 1767 1388
rect 1771 1384 1772 1388
rect 1766 1383 1772 1384
rect 1806 1388 1812 1389
rect 1832 1388 1834 1405
rect 1894 1403 1900 1404
rect 1894 1399 1895 1403
rect 1899 1399 1900 1403
rect 1894 1398 1900 1399
rect 1806 1384 1807 1388
rect 1811 1384 1812 1388
rect 1806 1383 1812 1384
rect 1830 1387 1836 1388
rect 1830 1383 1831 1387
rect 1835 1383 1836 1387
rect 1830 1382 1836 1383
rect 1086 1379 1092 1380
rect 1086 1375 1087 1379
rect 1091 1375 1092 1379
rect 1086 1374 1092 1375
rect 1238 1379 1244 1380
rect 1238 1375 1239 1379
rect 1243 1375 1244 1379
rect 1238 1374 1244 1375
rect 1374 1379 1380 1380
rect 1374 1375 1375 1379
rect 1379 1375 1380 1379
rect 1374 1374 1380 1375
rect 1502 1379 1508 1380
rect 1502 1375 1503 1379
rect 1507 1375 1508 1379
rect 1502 1374 1508 1375
rect 1510 1379 1516 1380
rect 1510 1375 1511 1379
rect 1515 1375 1516 1379
rect 1510 1374 1516 1375
rect 1742 1379 1748 1380
rect 1742 1375 1743 1379
rect 1747 1375 1748 1379
rect 1742 1374 1748 1375
rect 1750 1379 1756 1380
rect 1750 1375 1751 1379
rect 1755 1375 1756 1379
rect 1750 1374 1756 1375
rect 1014 1368 1020 1369
rect 1014 1364 1015 1368
rect 1019 1364 1020 1368
rect 1014 1363 1020 1364
rect 1166 1368 1172 1369
rect 1166 1364 1167 1368
rect 1171 1364 1172 1368
rect 1166 1363 1172 1364
rect 1302 1368 1308 1369
rect 1302 1364 1303 1368
rect 1307 1364 1308 1368
rect 1302 1363 1308 1364
rect 1430 1368 1436 1369
rect 1430 1364 1431 1368
rect 1435 1364 1436 1368
rect 1430 1363 1436 1364
rect 1016 1343 1018 1363
rect 1168 1343 1170 1363
rect 1304 1343 1306 1363
rect 1432 1343 1434 1363
rect 1015 1342 1019 1343
rect 1015 1337 1019 1338
rect 1063 1342 1067 1343
rect 1063 1337 1067 1338
rect 1167 1342 1171 1343
rect 1167 1337 1171 1338
rect 1223 1342 1227 1343
rect 1223 1337 1227 1338
rect 1303 1342 1307 1343
rect 1303 1337 1307 1338
rect 1375 1342 1379 1343
rect 1375 1337 1379 1338
rect 1431 1342 1435 1343
rect 1431 1337 1435 1338
rect 1064 1321 1066 1337
rect 1224 1321 1226 1337
rect 1376 1321 1378 1337
rect 1062 1320 1068 1321
rect 1062 1316 1063 1320
rect 1067 1316 1068 1320
rect 1062 1315 1068 1316
rect 1222 1320 1228 1321
rect 1222 1316 1223 1320
rect 1227 1316 1228 1320
rect 1222 1315 1228 1316
rect 1374 1320 1380 1321
rect 1374 1316 1375 1320
rect 1379 1316 1380 1320
rect 1374 1315 1380 1316
rect 206 1311 212 1312
rect 206 1307 207 1311
rect 211 1307 212 1311
rect 206 1306 212 1307
rect 318 1311 324 1312
rect 318 1307 319 1311
rect 323 1307 324 1311
rect 318 1306 324 1307
rect 470 1311 476 1312
rect 470 1307 471 1311
rect 475 1307 476 1311
rect 470 1306 476 1307
rect 498 1311 504 1312
rect 498 1307 499 1311
rect 503 1307 504 1311
rect 498 1306 504 1307
rect 798 1311 804 1312
rect 798 1307 799 1311
rect 803 1307 804 1311
rect 798 1306 804 1307
rect 966 1311 972 1312
rect 966 1307 967 1311
rect 971 1307 972 1311
rect 966 1306 972 1307
rect 974 1311 980 1312
rect 974 1307 975 1311
rect 979 1307 980 1311
rect 974 1306 980 1307
rect 1294 1311 1300 1312
rect 1294 1307 1295 1311
rect 1299 1307 1300 1311
rect 1294 1306 1300 1307
rect 1446 1311 1452 1312
rect 1446 1307 1447 1311
rect 1451 1307 1452 1311
rect 1446 1306 1452 1307
rect 208 1284 210 1306
rect 246 1301 252 1302
rect 246 1297 247 1301
rect 251 1297 252 1301
rect 246 1296 252 1297
rect 187 1279 191 1280
rect 198 1283 204 1284
rect 198 1279 199 1283
rect 203 1279 204 1283
rect 111 1274 115 1275
rect 111 1269 115 1270
rect 135 1274 139 1275
rect 135 1269 139 1270
rect 112 1253 114 1269
rect 110 1252 116 1253
rect 136 1252 138 1269
rect 188 1268 190 1279
rect 198 1278 204 1279
rect 206 1283 212 1284
rect 206 1279 207 1283
rect 211 1279 212 1283
rect 206 1278 212 1279
rect 248 1275 250 1296
rect 320 1284 322 1306
rect 398 1301 404 1302
rect 398 1297 399 1301
rect 403 1297 404 1301
rect 398 1296 404 1297
rect 318 1283 324 1284
rect 318 1279 319 1283
rect 323 1279 324 1283
rect 318 1278 324 1279
rect 400 1275 402 1296
rect 472 1284 474 1306
rect 500 1285 502 1306
rect 558 1301 564 1302
rect 558 1297 559 1301
rect 563 1297 564 1301
rect 558 1296 564 1297
rect 726 1301 732 1302
rect 726 1297 727 1301
rect 731 1297 732 1301
rect 726 1296 732 1297
rect 499 1284 503 1285
rect 470 1283 476 1284
rect 470 1279 471 1283
rect 475 1279 476 1283
rect 499 1279 503 1280
rect 470 1278 476 1279
rect 560 1275 562 1296
rect 728 1275 730 1296
rect 800 1284 802 1306
rect 894 1301 900 1302
rect 894 1297 895 1301
rect 899 1297 900 1301
rect 894 1296 900 1297
rect 750 1283 756 1284
rect 750 1279 751 1283
rect 755 1279 756 1283
rect 750 1278 756 1279
rect 798 1283 804 1284
rect 798 1279 799 1283
rect 803 1279 804 1283
rect 798 1278 804 1279
rect 223 1274 227 1275
rect 223 1269 227 1270
rect 247 1274 251 1275
rect 247 1269 251 1270
rect 319 1274 323 1275
rect 319 1269 323 1270
rect 399 1274 403 1275
rect 399 1269 403 1270
rect 431 1274 435 1275
rect 431 1269 435 1270
rect 551 1274 555 1275
rect 551 1269 555 1270
rect 559 1274 563 1275
rect 559 1269 563 1270
rect 679 1274 683 1275
rect 679 1269 683 1270
rect 727 1274 731 1275
rect 727 1269 731 1270
rect 186 1267 192 1268
rect 186 1263 187 1267
rect 191 1263 192 1267
rect 186 1262 192 1263
rect 206 1267 212 1268
rect 206 1263 207 1267
rect 211 1263 212 1267
rect 206 1262 212 1263
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 110 1247 116 1248
rect 134 1251 140 1252
rect 134 1247 135 1251
rect 139 1247 140 1251
rect 134 1246 140 1247
rect 208 1244 210 1262
rect 224 1252 226 1269
rect 294 1267 300 1268
rect 294 1263 295 1267
rect 299 1263 300 1267
rect 294 1262 300 1263
rect 222 1251 228 1252
rect 222 1247 223 1251
rect 227 1247 228 1251
rect 222 1246 228 1247
rect 296 1244 298 1262
rect 320 1252 322 1269
rect 390 1267 396 1268
rect 390 1263 391 1267
rect 395 1263 396 1267
rect 390 1262 396 1263
rect 318 1251 324 1252
rect 318 1247 319 1251
rect 323 1247 324 1251
rect 318 1246 324 1247
rect 392 1244 394 1262
rect 432 1252 434 1269
rect 502 1267 508 1268
rect 502 1263 503 1267
rect 507 1263 508 1267
rect 502 1262 508 1263
rect 430 1251 436 1252
rect 430 1247 431 1251
rect 435 1247 436 1251
rect 430 1246 436 1247
rect 504 1244 506 1262
rect 552 1252 554 1269
rect 680 1252 682 1269
rect 550 1251 556 1252
rect 550 1247 551 1251
rect 555 1247 556 1251
rect 550 1246 556 1247
rect 678 1251 684 1252
rect 678 1247 679 1251
rect 683 1247 684 1251
rect 678 1246 684 1247
rect 752 1244 754 1278
rect 896 1275 898 1296
rect 968 1284 970 1306
rect 1062 1301 1068 1302
rect 1062 1297 1063 1301
rect 1067 1297 1068 1301
rect 1062 1296 1068 1297
rect 1222 1301 1228 1302
rect 1222 1297 1223 1301
rect 1227 1297 1228 1301
rect 1222 1296 1228 1297
rect 966 1283 972 1284
rect 966 1279 967 1283
rect 971 1279 972 1283
rect 966 1278 972 1279
rect 1064 1275 1066 1296
rect 1224 1275 1226 1296
rect 1296 1284 1298 1306
rect 1374 1301 1380 1302
rect 1374 1297 1375 1301
rect 1379 1297 1380 1301
rect 1374 1296 1380 1297
rect 1294 1283 1300 1284
rect 1294 1279 1295 1283
rect 1299 1279 1300 1283
rect 1294 1278 1300 1279
rect 1376 1275 1378 1296
rect 1448 1284 1450 1306
rect 1446 1283 1452 1284
rect 1446 1279 1447 1283
rect 1451 1279 1452 1283
rect 1446 1278 1452 1279
rect 1512 1276 1514 1374
rect 1766 1371 1772 1372
rect 1558 1368 1564 1369
rect 1558 1364 1559 1368
rect 1563 1364 1564 1368
rect 1558 1363 1564 1364
rect 1670 1368 1676 1369
rect 1670 1364 1671 1368
rect 1675 1364 1676 1368
rect 1766 1367 1767 1371
rect 1771 1367 1772 1371
rect 1766 1366 1772 1367
rect 1806 1371 1812 1372
rect 1806 1367 1807 1371
rect 1811 1367 1812 1371
rect 1806 1366 1812 1367
rect 1830 1368 1836 1369
rect 1670 1363 1676 1364
rect 1560 1343 1562 1363
rect 1672 1343 1674 1363
rect 1768 1343 1770 1366
rect 1535 1342 1539 1343
rect 1535 1337 1539 1338
rect 1559 1342 1563 1343
rect 1559 1337 1563 1338
rect 1671 1342 1675 1343
rect 1671 1337 1675 1338
rect 1767 1342 1771 1343
rect 1808 1339 1810 1366
rect 1830 1364 1831 1368
rect 1835 1364 1836 1368
rect 1830 1363 1836 1364
rect 1832 1339 1834 1363
rect 1767 1337 1771 1338
rect 1807 1338 1811 1339
rect 1536 1321 1538 1337
rect 1672 1321 1674 1337
rect 1534 1320 1540 1321
rect 1534 1316 1535 1320
rect 1539 1316 1540 1320
rect 1534 1315 1540 1316
rect 1670 1320 1676 1321
rect 1670 1316 1671 1320
rect 1675 1316 1676 1320
rect 1768 1318 1770 1337
rect 1807 1333 1811 1334
rect 1831 1338 1835 1339
rect 1831 1333 1835 1334
rect 1670 1315 1676 1316
rect 1766 1317 1772 1318
rect 1766 1313 1767 1317
rect 1771 1313 1772 1317
rect 1808 1314 1810 1333
rect 1832 1317 1834 1333
rect 1830 1316 1836 1317
rect 1766 1312 1772 1313
rect 1806 1313 1812 1314
rect 1606 1311 1612 1312
rect 1606 1307 1607 1311
rect 1611 1307 1612 1311
rect 1606 1306 1612 1307
rect 1622 1311 1628 1312
rect 1622 1307 1623 1311
rect 1627 1307 1628 1311
rect 1806 1309 1807 1313
rect 1811 1309 1812 1313
rect 1830 1312 1831 1316
rect 1835 1312 1836 1316
rect 1830 1311 1836 1312
rect 1806 1308 1812 1309
rect 1896 1308 1898 1398
rect 2008 1388 2010 1405
rect 2078 1403 2084 1404
rect 2078 1399 2079 1403
rect 2083 1399 2084 1403
rect 2078 1398 2084 1399
rect 2006 1387 2012 1388
rect 2006 1383 2007 1387
rect 2011 1383 2012 1387
rect 2006 1382 2012 1383
rect 2080 1380 2082 1398
rect 2200 1388 2202 1405
rect 2334 1403 2340 1404
rect 2334 1399 2335 1403
rect 2339 1399 2340 1403
rect 2334 1398 2340 1399
rect 2198 1387 2204 1388
rect 2198 1383 2199 1387
rect 2203 1383 2204 1387
rect 2198 1382 2204 1383
rect 2336 1380 2338 1398
rect 2344 1380 2346 1406
rect 2383 1405 2387 1406
rect 2431 1410 2435 1411
rect 2431 1405 2435 1406
rect 2559 1410 2563 1411
rect 2559 1405 2563 1406
rect 2591 1410 2595 1411
rect 2591 1405 2595 1406
rect 2384 1388 2386 1405
rect 2560 1388 2562 1405
rect 2612 1404 2614 1458
rect 2736 1457 2738 1473
rect 2872 1457 2874 1473
rect 3008 1457 3010 1473
rect 2734 1456 2740 1457
rect 2734 1452 2735 1456
rect 2739 1452 2740 1456
rect 2734 1451 2740 1452
rect 2870 1456 2876 1457
rect 2870 1452 2871 1456
rect 2875 1452 2876 1456
rect 2870 1451 2876 1452
rect 3006 1456 3012 1457
rect 3006 1452 3007 1456
rect 3011 1452 3012 1456
rect 3006 1451 3012 1452
rect 2806 1447 2812 1448
rect 2806 1443 2807 1447
rect 2811 1443 2812 1447
rect 2806 1442 2812 1443
rect 2942 1447 2948 1448
rect 2942 1443 2943 1447
rect 2947 1443 2948 1447
rect 2942 1442 2948 1443
rect 2734 1437 2740 1438
rect 2734 1433 2735 1437
rect 2739 1433 2740 1437
rect 2734 1432 2740 1433
rect 2736 1411 2738 1432
rect 2808 1420 2810 1442
rect 2870 1437 2876 1438
rect 2870 1433 2871 1437
rect 2875 1433 2876 1437
rect 2870 1432 2876 1433
rect 2806 1419 2812 1420
rect 2806 1415 2807 1419
rect 2811 1415 2812 1419
rect 2806 1414 2812 1415
rect 2872 1411 2874 1432
rect 2944 1420 2946 1442
rect 3006 1437 3012 1438
rect 3006 1433 3007 1437
rect 3011 1433 3012 1437
rect 3006 1432 3012 1433
rect 2942 1419 2948 1420
rect 2942 1415 2943 1419
rect 2947 1415 2948 1419
rect 2942 1414 2948 1415
rect 3008 1411 3010 1432
rect 3020 1412 3022 1514
rect 3462 1511 3468 1512
rect 3054 1508 3060 1509
rect 3054 1504 3055 1508
rect 3059 1504 3060 1508
rect 3462 1507 3463 1511
rect 3467 1507 3468 1511
rect 3462 1506 3468 1507
rect 3054 1503 3060 1504
rect 3056 1479 3058 1503
rect 3464 1479 3466 1506
rect 3055 1478 3059 1479
rect 3055 1473 3059 1474
rect 3135 1478 3139 1479
rect 3135 1473 3139 1474
rect 3263 1478 3267 1479
rect 3263 1473 3267 1474
rect 3367 1478 3371 1479
rect 3367 1473 3371 1474
rect 3463 1478 3467 1479
rect 3463 1473 3467 1474
rect 3136 1457 3138 1473
rect 3264 1457 3266 1473
rect 3368 1457 3370 1473
rect 3134 1456 3140 1457
rect 3134 1452 3135 1456
rect 3139 1452 3140 1456
rect 3134 1451 3140 1452
rect 3262 1456 3268 1457
rect 3262 1452 3263 1456
rect 3267 1452 3268 1456
rect 3262 1451 3268 1452
rect 3366 1456 3372 1457
rect 3366 1452 3367 1456
rect 3371 1452 3372 1456
rect 3464 1454 3466 1473
rect 3366 1451 3372 1452
rect 3462 1453 3468 1454
rect 3462 1449 3463 1453
rect 3467 1449 3468 1453
rect 3462 1448 3468 1449
rect 3078 1447 3084 1448
rect 3078 1443 3079 1447
rect 3083 1443 3084 1447
rect 3078 1442 3084 1443
rect 3334 1447 3340 1448
rect 3334 1443 3335 1447
rect 3339 1443 3340 1447
rect 3334 1442 3340 1443
rect 3430 1447 3436 1448
rect 3430 1443 3431 1447
rect 3435 1443 3436 1447
rect 3430 1442 3436 1443
rect 3080 1420 3082 1442
rect 3134 1437 3140 1438
rect 3134 1433 3135 1437
rect 3139 1433 3140 1437
rect 3134 1432 3140 1433
rect 3262 1437 3268 1438
rect 3262 1433 3263 1437
rect 3267 1433 3268 1437
rect 3262 1432 3268 1433
rect 3078 1419 3084 1420
rect 3078 1415 3079 1419
rect 3083 1415 3084 1419
rect 3078 1414 3084 1415
rect 3018 1411 3024 1412
rect 3136 1411 3138 1432
rect 3264 1411 3266 1432
rect 3336 1420 3338 1442
rect 3366 1437 3372 1438
rect 3366 1433 3367 1437
rect 3371 1433 3372 1437
rect 3366 1432 3372 1433
rect 3326 1419 3332 1420
rect 3326 1415 3327 1419
rect 3331 1415 3332 1419
rect 3326 1414 3332 1415
rect 3334 1419 3340 1420
rect 3334 1415 3335 1419
rect 3339 1415 3340 1419
rect 3334 1414 3340 1415
rect 2719 1410 2723 1411
rect 2719 1405 2723 1406
rect 2735 1410 2739 1411
rect 2735 1405 2739 1406
rect 2863 1410 2867 1411
rect 2863 1405 2867 1406
rect 2871 1410 2875 1411
rect 2871 1405 2875 1406
rect 2999 1410 3003 1411
rect 2999 1405 3003 1406
rect 3007 1410 3011 1411
rect 3018 1407 3019 1411
rect 3023 1407 3024 1411
rect 3018 1406 3024 1407
rect 3127 1410 3131 1411
rect 3007 1405 3011 1406
rect 3127 1405 3131 1406
rect 3135 1410 3139 1411
rect 3135 1405 3139 1406
rect 3255 1410 3259 1411
rect 3255 1405 3259 1406
rect 3263 1410 3267 1411
rect 3263 1405 3267 1406
rect 2610 1403 2616 1404
rect 2610 1399 2611 1403
rect 2615 1399 2616 1403
rect 2610 1398 2616 1399
rect 2630 1403 2636 1404
rect 2630 1399 2631 1403
rect 2635 1399 2636 1403
rect 2630 1398 2636 1399
rect 2382 1387 2388 1388
rect 2382 1383 2383 1387
rect 2387 1383 2388 1387
rect 2382 1382 2388 1383
rect 2558 1387 2564 1388
rect 2558 1383 2559 1387
rect 2563 1383 2564 1387
rect 2558 1382 2564 1383
rect 2632 1380 2634 1398
rect 2720 1388 2722 1405
rect 2790 1403 2796 1404
rect 2790 1399 2791 1403
rect 2795 1399 2796 1403
rect 2790 1398 2796 1399
rect 2718 1387 2724 1388
rect 2718 1383 2719 1387
rect 2723 1383 2724 1387
rect 2718 1382 2724 1383
rect 2792 1380 2794 1398
rect 2864 1388 2866 1405
rect 2934 1403 2940 1404
rect 2934 1399 2935 1403
rect 2939 1399 2940 1403
rect 2934 1398 2940 1399
rect 2862 1387 2868 1388
rect 2862 1383 2863 1387
rect 2867 1383 2868 1387
rect 2862 1382 2868 1383
rect 2936 1380 2938 1398
rect 3000 1388 3002 1405
rect 3070 1403 3076 1404
rect 3070 1399 3071 1403
rect 3075 1399 3076 1403
rect 3070 1398 3076 1399
rect 2998 1387 3004 1388
rect 2998 1383 2999 1387
rect 3003 1383 3004 1387
rect 2998 1382 3004 1383
rect 3072 1380 3074 1398
rect 3128 1388 3130 1405
rect 3198 1403 3204 1404
rect 3198 1399 3199 1403
rect 3203 1399 3204 1403
rect 3198 1398 3204 1399
rect 3126 1387 3132 1388
rect 3126 1383 3127 1387
rect 3131 1383 3132 1387
rect 3126 1382 3132 1383
rect 3200 1380 3202 1398
rect 3256 1388 3258 1405
rect 3254 1387 3260 1388
rect 3254 1383 3255 1387
rect 3259 1383 3260 1387
rect 3254 1382 3260 1383
rect 3328 1380 3330 1414
rect 3368 1411 3370 1432
rect 3367 1410 3371 1411
rect 3367 1405 3371 1406
rect 3368 1388 3370 1405
rect 3432 1404 3434 1442
rect 3462 1436 3468 1437
rect 3462 1432 3463 1436
rect 3467 1432 3468 1436
rect 3462 1431 3468 1432
rect 3464 1411 3466 1431
rect 3463 1410 3467 1411
rect 3463 1405 3467 1406
rect 3430 1403 3436 1404
rect 3430 1399 3431 1403
rect 3435 1399 3436 1403
rect 3430 1398 3436 1399
rect 3464 1389 3466 1405
rect 3462 1388 3468 1389
rect 3366 1387 3372 1388
rect 3366 1383 3367 1387
rect 3371 1383 3372 1387
rect 3462 1384 3463 1388
rect 3467 1384 3468 1388
rect 3462 1383 3468 1384
rect 3366 1382 3372 1383
rect 2078 1379 2084 1380
rect 2078 1375 2079 1379
rect 2083 1375 2084 1379
rect 2078 1374 2084 1375
rect 2334 1379 2340 1380
rect 2334 1375 2335 1379
rect 2339 1375 2340 1379
rect 2334 1374 2340 1375
rect 2342 1379 2348 1380
rect 2342 1375 2343 1379
rect 2347 1375 2348 1379
rect 2342 1374 2348 1375
rect 2630 1379 2636 1380
rect 2630 1375 2631 1379
rect 2635 1375 2636 1379
rect 2630 1374 2636 1375
rect 2790 1379 2796 1380
rect 2790 1375 2791 1379
rect 2795 1375 2796 1379
rect 2790 1374 2796 1375
rect 2934 1379 2940 1380
rect 2934 1375 2935 1379
rect 2939 1375 2940 1379
rect 2934 1374 2940 1375
rect 3070 1379 3076 1380
rect 3070 1375 3071 1379
rect 3075 1375 3076 1379
rect 3070 1374 3076 1375
rect 3198 1379 3204 1380
rect 3198 1375 3199 1379
rect 3203 1375 3204 1379
rect 3198 1374 3204 1375
rect 3326 1379 3332 1380
rect 3326 1375 3327 1379
rect 3331 1375 3332 1379
rect 3326 1374 3332 1375
rect 3438 1375 3444 1376
rect 3438 1371 3439 1375
rect 3443 1371 3444 1375
rect 3438 1370 3444 1371
rect 3462 1371 3468 1372
rect 2006 1368 2012 1369
rect 2006 1364 2007 1368
rect 2011 1364 2012 1368
rect 2006 1363 2012 1364
rect 2198 1368 2204 1369
rect 2198 1364 2199 1368
rect 2203 1364 2204 1368
rect 2198 1363 2204 1364
rect 2382 1368 2388 1369
rect 2382 1364 2383 1368
rect 2387 1364 2388 1368
rect 2382 1363 2388 1364
rect 2558 1368 2564 1369
rect 2558 1364 2559 1368
rect 2563 1364 2564 1368
rect 2558 1363 2564 1364
rect 2718 1368 2724 1369
rect 2718 1364 2719 1368
rect 2723 1364 2724 1368
rect 2718 1363 2724 1364
rect 2862 1368 2868 1369
rect 2862 1364 2863 1368
rect 2867 1364 2868 1368
rect 2862 1363 2868 1364
rect 2998 1368 3004 1369
rect 2998 1364 2999 1368
rect 3003 1364 3004 1368
rect 2998 1363 3004 1364
rect 3126 1368 3132 1369
rect 3126 1364 3127 1368
rect 3131 1364 3132 1368
rect 3126 1363 3132 1364
rect 3254 1368 3260 1369
rect 3254 1364 3255 1368
rect 3259 1364 3260 1368
rect 3254 1363 3260 1364
rect 3366 1368 3372 1369
rect 3366 1364 3367 1368
rect 3371 1364 3372 1368
rect 3366 1363 3372 1364
rect 2008 1339 2010 1363
rect 2200 1339 2202 1363
rect 2384 1339 2386 1363
rect 2560 1339 2562 1363
rect 2720 1339 2722 1363
rect 2864 1339 2866 1363
rect 3000 1339 3002 1363
rect 3128 1339 3130 1363
rect 3256 1339 3258 1363
rect 3368 1339 3370 1363
rect 1967 1338 1971 1339
rect 1967 1333 1971 1334
rect 2007 1338 2011 1339
rect 2007 1333 2011 1334
rect 2143 1338 2147 1339
rect 2143 1333 2147 1334
rect 2199 1338 2203 1339
rect 2199 1333 2203 1334
rect 2327 1338 2331 1339
rect 2327 1333 2331 1334
rect 2383 1338 2387 1339
rect 2383 1333 2387 1334
rect 2511 1338 2515 1339
rect 2511 1333 2515 1334
rect 2559 1338 2563 1339
rect 2559 1333 2563 1334
rect 2687 1338 2691 1339
rect 2687 1333 2691 1334
rect 2719 1338 2723 1339
rect 2719 1333 2723 1334
rect 2863 1338 2867 1339
rect 2863 1333 2867 1334
rect 2999 1338 3003 1339
rect 2999 1333 3003 1334
rect 3039 1338 3043 1339
rect 3039 1333 3043 1334
rect 3127 1338 3131 1339
rect 3127 1333 3131 1334
rect 3215 1338 3219 1339
rect 3215 1333 3219 1334
rect 3255 1338 3259 1339
rect 3255 1333 3259 1334
rect 3367 1338 3371 1339
rect 3367 1333 3371 1334
rect 1968 1317 1970 1333
rect 2018 1323 2024 1324
rect 2018 1319 2019 1323
rect 2023 1319 2024 1323
rect 2018 1318 2024 1319
rect 1966 1316 1972 1317
rect 1966 1312 1967 1316
rect 1971 1312 1972 1316
rect 1966 1311 1972 1312
rect 1622 1306 1628 1307
rect 1894 1307 1900 1308
rect 1534 1301 1540 1302
rect 1534 1297 1535 1301
rect 1539 1297 1540 1301
rect 1534 1296 1540 1297
rect 1510 1275 1516 1276
rect 1536 1275 1538 1296
rect 1608 1284 1610 1306
rect 1606 1283 1612 1284
rect 1606 1279 1607 1283
rect 1611 1279 1612 1283
rect 1606 1278 1612 1279
rect 1624 1276 1626 1306
rect 1894 1303 1895 1307
rect 1899 1303 1900 1307
rect 1894 1302 1900 1303
rect 1910 1307 1916 1308
rect 1910 1303 1911 1307
rect 1915 1303 1916 1307
rect 1910 1302 1916 1303
rect 1670 1301 1676 1302
rect 1670 1297 1671 1301
rect 1675 1297 1676 1301
rect 1670 1296 1676 1297
rect 1766 1300 1772 1301
rect 1766 1296 1767 1300
rect 1771 1296 1772 1300
rect 1830 1297 1836 1298
rect 1622 1275 1628 1276
rect 1672 1275 1674 1296
rect 1766 1295 1772 1296
rect 1806 1296 1812 1297
rect 1768 1275 1770 1295
rect 1806 1292 1807 1296
rect 1811 1292 1812 1296
rect 1830 1293 1831 1297
rect 1835 1293 1836 1297
rect 1830 1292 1836 1293
rect 1806 1291 1812 1292
rect 1808 1275 1810 1291
rect 1832 1275 1834 1292
rect 1912 1280 1914 1302
rect 1966 1297 1972 1298
rect 1966 1293 1967 1297
rect 1971 1293 1972 1297
rect 1966 1292 1972 1293
rect 1910 1279 1916 1280
rect 1910 1275 1911 1279
rect 1915 1275 1916 1279
rect 1968 1275 1970 1292
rect 2020 1280 2022 1318
rect 2144 1317 2146 1333
rect 2328 1317 2330 1333
rect 2512 1317 2514 1333
rect 2688 1317 2690 1333
rect 2864 1317 2866 1333
rect 3040 1317 3042 1333
rect 3216 1317 3218 1333
rect 3368 1317 3370 1333
rect 2142 1316 2148 1317
rect 2142 1312 2143 1316
rect 2147 1312 2148 1316
rect 2142 1311 2148 1312
rect 2326 1316 2332 1317
rect 2326 1312 2327 1316
rect 2331 1312 2332 1316
rect 2326 1311 2332 1312
rect 2510 1316 2516 1317
rect 2510 1312 2511 1316
rect 2515 1312 2516 1316
rect 2510 1311 2516 1312
rect 2686 1316 2692 1317
rect 2686 1312 2687 1316
rect 2691 1312 2692 1316
rect 2686 1311 2692 1312
rect 2862 1316 2868 1317
rect 2862 1312 2863 1316
rect 2867 1312 2868 1316
rect 2862 1311 2868 1312
rect 3038 1316 3044 1317
rect 3038 1312 3039 1316
rect 3043 1312 3044 1316
rect 3038 1311 3044 1312
rect 3214 1316 3220 1317
rect 3214 1312 3215 1316
rect 3219 1312 3220 1316
rect 3214 1311 3220 1312
rect 3366 1316 3372 1317
rect 3366 1312 3367 1316
rect 3371 1312 3372 1316
rect 3366 1311 3372 1312
rect 2214 1307 2220 1308
rect 2214 1303 2215 1307
rect 2219 1303 2220 1307
rect 2214 1302 2220 1303
rect 2398 1307 2404 1308
rect 2398 1303 2399 1307
rect 2403 1303 2404 1307
rect 2398 1302 2404 1303
rect 2758 1307 2764 1308
rect 2758 1303 2759 1307
rect 2763 1303 2764 1307
rect 2758 1302 2764 1303
rect 2766 1307 2772 1308
rect 2766 1303 2767 1307
rect 2771 1303 2772 1307
rect 2766 1302 2772 1303
rect 2942 1307 2948 1308
rect 2942 1303 2943 1307
rect 2947 1303 2948 1307
rect 2942 1302 2948 1303
rect 3118 1307 3124 1308
rect 3118 1303 3119 1307
rect 3123 1303 3124 1307
rect 3118 1302 3124 1303
rect 3430 1307 3436 1308
rect 3430 1303 3431 1307
rect 3435 1303 3436 1307
rect 3430 1302 3436 1303
rect 2142 1297 2148 1298
rect 2142 1293 2143 1297
rect 2147 1293 2148 1297
rect 2142 1292 2148 1293
rect 2018 1279 2024 1280
rect 2018 1275 2019 1279
rect 2023 1275 2024 1279
rect 2144 1275 2146 1292
rect 2216 1280 2218 1302
rect 2326 1297 2332 1298
rect 2326 1293 2327 1297
rect 2331 1293 2332 1297
rect 2326 1292 2332 1293
rect 2166 1279 2172 1280
rect 2166 1275 2167 1279
rect 2171 1275 2172 1279
rect 823 1274 827 1275
rect 823 1269 827 1270
rect 895 1274 899 1275
rect 895 1269 899 1270
rect 975 1274 979 1275
rect 975 1269 979 1270
rect 1063 1274 1067 1275
rect 1063 1269 1067 1270
rect 1143 1274 1147 1275
rect 1143 1269 1147 1270
rect 1223 1274 1227 1275
rect 1223 1269 1227 1270
rect 1319 1274 1323 1275
rect 1319 1269 1323 1270
rect 1375 1274 1379 1275
rect 1375 1269 1379 1270
rect 1503 1274 1507 1275
rect 1510 1271 1511 1275
rect 1515 1271 1516 1275
rect 1510 1270 1516 1271
rect 1535 1274 1539 1275
rect 1622 1271 1623 1275
rect 1627 1271 1628 1275
rect 1622 1270 1628 1271
rect 1671 1274 1675 1275
rect 1503 1269 1507 1270
rect 1535 1269 1539 1270
rect 1671 1269 1675 1270
rect 1767 1274 1771 1275
rect 1767 1269 1771 1270
rect 1807 1274 1811 1275
rect 1807 1269 1811 1270
rect 1831 1274 1835 1275
rect 1910 1274 1916 1275
rect 1967 1274 1971 1275
rect 2018 1274 2024 1275
rect 2095 1274 2099 1275
rect 1831 1269 1835 1270
rect 1967 1269 1971 1270
rect 2095 1269 2099 1270
rect 2143 1274 2147 1275
rect 2166 1274 2172 1275
rect 2214 1279 2220 1280
rect 2214 1275 2215 1279
rect 2219 1275 2220 1279
rect 2328 1275 2330 1292
rect 2400 1280 2402 1302
rect 2510 1297 2516 1298
rect 2510 1293 2511 1297
rect 2515 1293 2516 1297
rect 2510 1292 2516 1293
rect 2686 1297 2692 1298
rect 2686 1293 2687 1297
rect 2691 1293 2692 1297
rect 2686 1292 2692 1293
rect 2398 1279 2404 1280
rect 2398 1275 2399 1279
rect 2403 1275 2404 1279
rect 2512 1275 2514 1292
rect 2678 1275 2684 1276
rect 2688 1275 2690 1292
rect 2214 1274 2220 1275
rect 2327 1274 2331 1275
rect 2143 1269 2147 1270
rect 758 1267 764 1268
rect 758 1263 759 1267
rect 763 1263 764 1267
rect 758 1262 764 1263
rect 760 1244 762 1262
rect 824 1252 826 1269
rect 902 1267 908 1268
rect 902 1263 903 1267
rect 907 1263 908 1267
rect 902 1262 908 1263
rect 822 1251 828 1252
rect 822 1247 823 1251
rect 827 1247 828 1251
rect 822 1246 828 1247
rect 904 1244 906 1262
rect 976 1252 978 1269
rect 1090 1267 1096 1268
rect 1090 1263 1091 1267
rect 1095 1263 1096 1267
rect 1090 1262 1096 1263
rect 974 1251 980 1252
rect 974 1247 975 1251
rect 979 1247 980 1251
rect 974 1246 980 1247
rect 1092 1244 1094 1262
rect 1144 1252 1146 1269
rect 1320 1252 1322 1269
rect 1326 1267 1332 1268
rect 1326 1263 1327 1267
rect 1331 1263 1332 1267
rect 1326 1262 1332 1263
rect 1142 1251 1148 1252
rect 1142 1247 1143 1251
rect 1147 1247 1148 1251
rect 1142 1246 1148 1247
rect 1318 1251 1324 1252
rect 1318 1247 1319 1251
rect 1323 1247 1324 1251
rect 1318 1246 1324 1247
rect 206 1243 212 1244
rect 206 1239 207 1243
rect 211 1239 212 1243
rect 206 1238 212 1239
rect 294 1243 300 1244
rect 294 1239 295 1243
rect 299 1239 300 1243
rect 294 1238 300 1239
rect 390 1243 396 1244
rect 390 1239 391 1243
rect 395 1239 396 1243
rect 390 1238 396 1239
rect 502 1243 508 1244
rect 502 1239 503 1243
rect 507 1239 508 1243
rect 502 1238 508 1239
rect 510 1243 516 1244
rect 510 1239 511 1243
rect 515 1239 516 1243
rect 510 1238 516 1239
rect 750 1243 756 1244
rect 750 1239 751 1243
rect 755 1239 756 1243
rect 750 1238 756 1239
rect 758 1243 764 1244
rect 758 1239 759 1243
rect 763 1239 764 1243
rect 758 1238 764 1239
rect 902 1243 908 1244
rect 902 1239 903 1243
rect 907 1239 908 1243
rect 902 1238 908 1239
rect 1090 1243 1096 1244
rect 1090 1239 1091 1243
rect 1095 1239 1096 1243
rect 1090 1238 1096 1239
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 110 1230 116 1231
rect 134 1232 140 1233
rect 112 1203 114 1230
rect 134 1228 135 1232
rect 139 1228 140 1232
rect 134 1227 140 1228
rect 222 1232 228 1233
rect 222 1228 223 1232
rect 227 1228 228 1232
rect 222 1227 228 1228
rect 318 1232 324 1233
rect 318 1228 319 1232
rect 323 1228 324 1232
rect 318 1227 324 1228
rect 430 1232 436 1233
rect 430 1228 431 1232
rect 435 1228 436 1232
rect 430 1227 436 1228
rect 136 1203 138 1227
rect 224 1203 226 1227
rect 320 1203 322 1227
rect 432 1203 434 1227
rect 111 1202 115 1203
rect 111 1197 115 1198
rect 135 1202 139 1203
rect 135 1197 139 1198
rect 223 1202 227 1203
rect 223 1197 227 1198
rect 231 1202 235 1203
rect 231 1197 235 1198
rect 319 1202 323 1203
rect 319 1197 323 1198
rect 359 1202 363 1203
rect 359 1197 363 1198
rect 431 1202 435 1203
rect 431 1197 435 1198
rect 487 1202 491 1203
rect 487 1197 491 1198
rect 112 1178 114 1197
rect 136 1181 138 1197
rect 186 1195 192 1196
rect 186 1191 187 1195
rect 191 1191 192 1195
rect 186 1190 192 1191
rect 134 1180 140 1181
rect 110 1177 116 1178
rect 110 1173 111 1177
rect 115 1173 116 1177
rect 134 1176 135 1180
rect 139 1176 140 1180
rect 134 1175 140 1176
rect 110 1172 116 1173
rect 134 1161 140 1162
rect 110 1160 116 1161
rect 110 1156 111 1160
rect 115 1156 116 1160
rect 134 1157 135 1161
rect 139 1157 140 1161
rect 134 1156 140 1157
rect 110 1155 116 1156
rect 112 1135 114 1155
rect 136 1135 138 1156
rect 188 1144 190 1190
rect 232 1181 234 1197
rect 360 1181 362 1197
rect 488 1181 490 1197
rect 512 1196 514 1238
rect 550 1232 556 1233
rect 550 1228 551 1232
rect 555 1228 556 1232
rect 550 1227 556 1228
rect 678 1232 684 1233
rect 678 1228 679 1232
rect 683 1228 684 1232
rect 678 1227 684 1228
rect 822 1232 828 1233
rect 822 1228 823 1232
rect 827 1228 828 1232
rect 822 1227 828 1228
rect 974 1232 980 1233
rect 974 1228 975 1232
rect 979 1228 980 1232
rect 974 1227 980 1228
rect 1142 1232 1148 1233
rect 1142 1228 1143 1232
rect 1147 1228 1148 1232
rect 1142 1227 1148 1228
rect 1318 1232 1324 1233
rect 1318 1228 1319 1232
rect 1323 1228 1324 1232
rect 1318 1227 1324 1228
rect 552 1203 554 1227
rect 680 1203 682 1227
rect 824 1203 826 1227
rect 976 1203 978 1227
rect 1144 1203 1146 1227
rect 1320 1203 1322 1227
rect 551 1202 555 1203
rect 551 1197 555 1198
rect 615 1202 619 1203
rect 615 1197 619 1198
rect 679 1202 683 1203
rect 679 1197 683 1198
rect 743 1202 747 1203
rect 743 1197 747 1198
rect 823 1202 827 1203
rect 823 1197 827 1198
rect 871 1202 875 1203
rect 871 1197 875 1198
rect 975 1202 979 1203
rect 975 1197 979 1198
rect 991 1202 995 1203
rect 991 1197 995 1198
rect 1119 1202 1123 1203
rect 1119 1197 1123 1198
rect 1143 1202 1147 1203
rect 1143 1197 1147 1198
rect 1247 1202 1251 1203
rect 1247 1197 1251 1198
rect 1319 1202 1323 1203
rect 1319 1197 1323 1198
rect 510 1195 516 1196
rect 510 1191 511 1195
rect 515 1191 516 1195
rect 510 1190 516 1191
rect 616 1181 618 1197
rect 744 1181 746 1197
rect 872 1181 874 1197
rect 992 1181 994 1197
rect 1120 1181 1122 1197
rect 1248 1181 1250 1197
rect 230 1180 236 1181
rect 230 1176 231 1180
rect 235 1176 236 1180
rect 230 1175 236 1176
rect 358 1180 364 1181
rect 358 1176 359 1180
rect 363 1176 364 1180
rect 358 1175 364 1176
rect 486 1180 492 1181
rect 486 1176 487 1180
rect 491 1176 492 1180
rect 486 1175 492 1176
rect 614 1180 620 1181
rect 614 1176 615 1180
rect 619 1176 620 1180
rect 614 1175 620 1176
rect 742 1180 748 1181
rect 742 1176 743 1180
rect 747 1176 748 1180
rect 742 1175 748 1176
rect 870 1180 876 1181
rect 870 1176 871 1180
rect 875 1176 876 1180
rect 870 1175 876 1176
rect 990 1180 996 1181
rect 990 1176 991 1180
rect 995 1176 996 1180
rect 990 1175 996 1176
rect 1118 1180 1124 1181
rect 1118 1176 1119 1180
rect 1123 1176 1124 1180
rect 1118 1175 1124 1176
rect 1246 1180 1252 1181
rect 1246 1176 1247 1180
rect 1251 1176 1252 1180
rect 1246 1175 1252 1176
rect 1328 1172 1330 1262
rect 1504 1252 1506 1269
rect 1574 1267 1580 1268
rect 1574 1263 1575 1267
rect 1579 1263 1580 1267
rect 1574 1262 1580 1263
rect 1502 1251 1508 1252
rect 1502 1247 1503 1251
rect 1507 1247 1508 1251
rect 1502 1246 1508 1247
rect 1576 1244 1578 1262
rect 1672 1252 1674 1269
rect 1742 1267 1748 1268
rect 1742 1263 1743 1267
rect 1747 1263 1748 1267
rect 1742 1262 1748 1263
rect 1670 1251 1676 1252
rect 1670 1247 1671 1251
rect 1675 1247 1676 1251
rect 1670 1246 1676 1247
rect 1744 1244 1746 1262
rect 1768 1253 1770 1269
rect 1808 1253 1810 1269
rect 1766 1252 1772 1253
rect 1766 1248 1767 1252
rect 1771 1248 1772 1252
rect 1766 1247 1772 1248
rect 1806 1252 1812 1253
rect 1832 1252 1834 1269
rect 1902 1267 1908 1268
rect 1902 1263 1903 1267
rect 1907 1263 1908 1267
rect 1902 1262 1908 1263
rect 1806 1248 1807 1252
rect 1811 1248 1812 1252
rect 1806 1247 1812 1248
rect 1830 1251 1836 1252
rect 1830 1247 1831 1251
rect 1835 1247 1836 1251
rect 1830 1246 1836 1247
rect 1904 1244 1906 1262
rect 2096 1252 2098 1269
rect 2094 1251 2100 1252
rect 2094 1247 2095 1251
rect 2099 1247 2100 1251
rect 2094 1246 2100 1247
rect 2168 1244 2170 1274
rect 2327 1269 2331 1270
rect 2359 1274 2363 1275
rect 2398 1274 2404 1275
rect 2511 1274 2515 1275
rect 2359 1269 2363 1270
rect 2511 1269 2515 1270
rect 2599 1274 2603 1275
rect 2678 1271 2679 1275
rect 2683 1271 2684 1275
rect 2678 1270 2684 1271
rect 2687 1274 2691 1275
rect 2599 1269 2603 1270
rect 2360 1252 2362 1269
rect 2430 1267 2436 1268
rect 2430 1263 2431 1267
rect 2435 1263 2436 1267
rect 2430 1262 2436 1263
rect 2358 1251 2364 1252
rect 2358 1247 2359 1251
rect 2363 1247 2364 1251
rect 2358 1246 2364 1247
rect 2432 1244 2434 1262
rect 2600 1252 2602 1269
rect 2598 1251 2604 1252
rect 2598 1247 2599 1251
rect 2603 1247 2604 1251
rect 2598 1246 2604 1247
rect 2680 1244 2682 1270
rect 2687 1269 2691 1270
rect 2760 1268 2762 1302
rect 2768 1280 2770 1302
rect 2862 1297 2868 1298
rect 2862 1293 2863 1297
rect 2867 1293 2868 1297
rect 2862 1292 2868 1293
rect 2766 1279 2772 1280
rect 2766 1275 2767 1279
rect 2771 1275 2772 1279
rect 2864 1275 2866 1292
rect 2944 1280 2946 1302
rect 3038 1297 3044 1298
rect 3038 1293 3039 1297
rect 3043 1293 3044 1297
rect 3038 1292 3044 1293
rect 2942 1279 2948 1280
rect 2942 1275 2943 1279
rect 2947 1275 2948 1279
rect 3040 1275 3042 1292
rect 3120 1280 3122 1302
rect 3214 1297 3220 1298
rect 3214 1293 3215 1297
rect 3219 1293 3220 1297
rect 3214 1292 3220 1293
rect 3366 1297 3372 1298
rect 3366 1293 3367 1297
rect 3371 1293 3372 1297
rect 3366 1292 3372 1293
rect 3118 1279 3124 1280
rect 3118 1275 3119 1279
rect 3123 1275 3124 1279
rect 3216 1275 3218 1292
rect 3262 1279 3268 1280
rect 3262 1275 3263 1279
rect 3267 1275 3268 1279
rect 3368 1275 3370 1292
rect 2766 1274 2772 1275
rect 2807 1274 2811 1275
rect 2807 1269 2811 1270
rect 2863 1274 2867 1275
rect 2942 1274 2948 1275
rect 3007 1274 3011 1275
rect 2863 1269 2867 1270
rect 3007 1269 3011 1270
rect 3039 1274 3043 1275
rect 3118 1274 3124 1275
rect 3199 1274 3203 1275
rect 3039 1269 3043 1270
rect 3199 1269 3203 1270
rect 3215 1274 3219 1275
rect 3262 1274 3268 1275
rect 3367 1274 3371 1275
rect 3215 1269 3219 1270
rect 2758 1267 2764 1268
rect 2758 1263 2759 1267
rect 2763 1263 2764 1267
rect 2758 1262 2764 1263
rect 2808 1252 2810 1269
rect 3008 1252 3010 1269
rect 3086 1267 3092 1268
rect 3086 1263 3087 1267
rect 3091 1263 3092 1267
rect 3086 1262 3092 1263
rect 3146 1267 3152 1268
rect 3146 1263 3147 1267
rect 3151 1263 3152 1267
rect 3146 1262 3152 1263
rect 2806 1251 2812 1252
rect 2806 1247 2807 1251
rect 2811 1247 2812 1251
rect 2806 1246 2812 1247
rect 3006 1251 3012 1252
rect 3006 1247 3007 1251
rect 3011 1247 3012 1251
rect 3006 1246 3012 1247
rect 1574 1243 1580 1244
rect 1574 1239 1575 1243
rect 1579 1239 1580 1243
rect 1574 1238 1580 1239
rect 1742 1243 1748 1244
rect 1742 1239 1743 1243
rect 1747 1239 1748 1243
rect 1742 1238 1748 1239
rect 1902 1243 1908 1244
rect 1902 1239 1903 1243
rect 1907 1239 1908 1243
rect 1902 1238 1908 1239
rect 2166 1243 2172 1244
rect 2166 1239 2167 1243
rect 2171 1239 2172 1243
rect 2166 1238 2172 1239
rect 2430 1243 2436 1244
rect 2430 1239 2431 1243
rect 2435 1239 2436 1243
rect 2678 1243 2684 1244
rect 2430 1238 2436 1239
rect 2670 1239 2676 1240
rect 1766 1235 1772 1236
rect 1502 1232 1508 1233
rect 1502 1228 1503 1232
rect 1507 1228 1508 1232
rect 1502 1227 1508 1228
rect 1670 1232 1676 1233
rect 1670 1228 1671 1232
rect 1675 1228 1676 1232
rect 1766 1231 1767 1235
rect 1771 1231 1772 1235
rect 1766 1230 1772 1231
rect 1806 1235 1812 1236
rect 1806 1231 1807 1235
rect 1811 1231 1812 1235
rect 2670 1235 2671 1239
rect 2675 1235 2676 1239
rect 2678 1239 2679 1243
rect 2683 1239 2684 1243
rect 2678 1238 2684 1239
rect 2670 1234 2676 1235
rect 1806 1230 1812 1231
rect 1830 1232 1836 1233
rect 1670 1227 1676 1228
rect 1504 1203 1506 1227
rect 1672 1203 1674 1227
rect 1768 1203 1770 1230
rect 1808 1203 1810 1230
rect 1830 1228 1831 1232
rect 1835 1228 1836 1232
rect 1830 1227 1836 1228
rect 2094 1232 2100 1233
rect 2094 1228 2095 1232
rect 2099 1228 2100 1232
rect 2094 1227 2100 1228
rect 2358 1232 2364 1233
rect 2358 1228 2359 1232
rect 2363 1228 2364 1232
rect 2358 1227 2364 1228
rect 2598 1232 2604 1233
rect 2598 1228 2599 1232
rect 2603 1228 2604 1232
rect 2598 1227 2604 1228
rect 1832 1203 1834 1227
rect 2096 1203 2098 1227
rect 2360 1203 2362 1227
rect 2600 1203 2602 1227
rect 1503 1202 1507 1203
rect 1503 1197 1507 1198
rect 1671 1202 1675 1203
rect 1671 1197 1675 1198
rect 1767 1202 1771 1203
rect 1767 1197 1771 1198
rect 1807 1202 1811 1203
rect 1807 1197 1811 1198
rect 1831 1202 1835 1203
rect 1831 1197 1835 1198
rect 1935 1202 1939 1203
rect 1935 1197 1939 1198
rect 2039 1202 2043 1203
rect 2039 1197 2043 1198
rect 2095 1202 2099 1203
rect 2095 1197 2099 1198
rect 2159 1202 2163 1203
rect 2159 1197 2163 1198
rect 2287 1202 2291 1203
rect 2287 1197 2291 1198
rect 2359 1202 2363 1203
rect 2359 1197 2363 1198
rect 2423 1202 2427 1203
rect 2423 1197 2427 1198
rect 2567 1202 2571 1203
rect 2567 1197 2571 1198
rect 2599 1202 2603 1203
rect 2599 1197 2603 1198
rect 1768 1178 1770 1197
rect 1808 1178 1810 1197
rect 1936 1181 1938 1197
rect 2040 1181 2042 1197
rect 2160 1181 2162 1197
rect 2288 1181 2290 1197
rect 2424 1181 2426 1197
rect 2568 1181 2570 1197
rect 1934 1180 1940 1181
rect 1766 1177 1772 1178
rect 1766 1173 1767 1177
rect 1771 1173 1772 1177
rect 1766 1172 1772 1173
rect 1806 1177 1812 1178
rect 1806 1173 1807 1177
rect 1811 1173 1812 1177
rect 1934 1176 1935 1180
rect 1939 1176 1940 1180
rect 1934 1175 1940 1176
rect 2038 1180 2044 1181
rect 2038 1176 2039 1180
rect 2043 1176 2044 1180
rect 2038 1175 2044 1176
rect 2158 1180 2164 1181
rect 2158 1176 2159 1180
rect 2163 1176 2164 1180
rect 2158 1175 2164 1176
rect 2286 1180 2292 1181
rect 2286 1176 2287 1180
rect 2291 1176 2292 1180
rect 2286 1175 2292 1176
rect 2422 1180 2428 1181
rect 2422 1176 2423 1180
rect 2427 1176 2428 1180
rect 2422 1175 2428 1176
rect 2566 1180 2572 1181
rect 2566 1176 2567 1180
rect 2571 1176 2572 1180
rect 2566 1175 2572 1176
rect 1806 1172 1812 1173
rect 206 1171 212 1172
rect 206 1167 207 1171
rect 211 1167 212 1171
rect 206 1166 212 1167
rect 302 1171 308 1172
rect 302 1167 303 1171
rect 307 1167 308 1171
rect 302 1166 308 1167
rect 430 1171 436 1172
rect 430 1167 431 1171
rect 435 1167 436 1171
rect 430 1166 436 1167
rect 558 1171 564 1172
rect 558 1167 559 1171
rect 563 1167 564 1171
rect 558 1166 564 1167
rect 566 1171 572 1172
rect 566 1167 567 1171
rect 571 1167 572 1171
rect 566 1166 572 1167
rect 814 1171 820 1172
rect 814 1167 815 1171
rect 819 1167 820 1171
rect 814 1166 820 1167
rect 942 1171 948 1172
rect 942 1167 943 1171
rect 947 1167 948 1171
rect 942 1166 948 1167
rect 1062 1171 1068 1172
rect 1062 1167 1063 1171
rect 1067 1167 1068 1171
rect 1062 1166 1068 1167
rect 1190 1171 1196 1172
rect 1190 1167 1191 1171
rect 1195 1167 1196 1171
rect 1190 1166 1196 1167
rect 1326 1171 1332 1172
rect 1326 1167 1327 1171
rect 1331 1167 1332 1171
rect 1326 1166 1332 1167
rect 2002 1171 2008 1172
rect 2002 1167 2003 1171
rect 2007 1167 2008 1171
rect 2002 1166 2008 1167
rect 2014 1171 2020 1172
rect 2014 1167 2015 1171
rect 2019 1167 2020 1171
rect 2014 1166 2020 1167
rect 2118 1171 2124 1172
rect 2118 1167 2119 1171
rect 2123 1167 2124 1171
rect 2118 1166 2124 1167
rect 2238 1171 2244 1172
rect 2238 1167 2239 1171
rect 2243 1167 2244 1171
rect 2238 1166 2244 1167
rect 2366 1171 2372 1172
rect 2366 1167 2367 1171
rect 2371 1167 2372 1171
rect 2366 1166 2372 1167
rect 2502 1171 2508 1172
rect 2502 1167 2503 1171
rect 2507 1167 2508 1171
rect 2502 1166 2508 1167
rect 208 1144 210 1166
rect 230 1161 236 1162
rect 230 1157 231 1161
rect 235 1157 236 1161
rect 230 1156 236 1157
rect 186 1143 192 1144
rect 186 1139 187 1143
rect 191 1139 192 1143
rect 186 1138 192 1139
rect 206 1143 212 1144
rect 206 1139 207 1143
rect 211 1139 212 1143
rect 206 1138 212 1139
rect 232 1135 234 1156
rect 304 1144 306 1166
rect 358 1161 364 1162
rect 358 1157 359 1161
rect 363 1157 364 1161
rect 358 1156 364 1157
rect 302 1143 308 1144
rect 302 1139 303 1143
rect 307 1139 308 1143
rect 302 1138 308 1139
rect 360 1135 362 1156
rect 432 1144 434 1166
rect 486 1161 492 1162
rect 486 1157 487 1161
rect 491 1157 492 1161
rect 486 1156 492 1157
rect 430 1143 436 1144
rect 430 1139 431 1143
rect 435 1139 436 1143
rect 430 1138 436 1139
rect 488 1135 490 1156
rect 560 1144 562 1166
rect 558 1143 564 1144
rect 558 1139 559 1143
rect 563 1139 564 1143
rect 558 1138 564 1139
rect 568 1136 570 1166
rect 614 1161 620 1162
rect 614 1157 615 1161
rect 619 1157 620 1161
rect 614 1156 620 1157
rect 742 1161 748 1162
rect 742 1157 743 1161
rect 747 1157 748 1161
rect 742 1156 748 1157
rect 566 1135 572 1136
rect 616 1135 618 1156
rect 744 1135 746 1156
rect 816 1144 818 1166
rect 870 1161 876 1162
rect 870 1157 871 1161
rect 875 1157 876 1161
rect 870 1156 876 1157
rect 814 1143 820 1144
rect 814 1139 815 1143
rect 819 1139 820 1143
rect 814 1138 820 1139
rect 838 1135 844 1136
rect 872 1135 874 1156
rect 944 1144 946 1166
rect 990 1161 996 1162
rect 990 1157 991 1161
rect 995 1157 996 1161
rect 990 1156 996 1157
rect 942 1143 948 1144
rect 942 1139 943 1143
rect 947 1139 948 1143
rect 942 1138 948 1139
rect 992 1135 994 1156
rect 1064 1144 1066 1166
rect 1118 1161 1124 1162
rect 1118 1157 1119 1161
rect 1123 1157 1124 1161
rect 1118 1156 1124 1157
rect 1062 1143 1068 1144
rect 1062 1139 1063 1143
rect 1067 1139 1068 1143
rect 1062 1138 1068 1139
rect 1120 1135 1122 1156
rect 1192 1144 1194 1166
rect 1246 1161 1252 1162
rect 1934 1161 1940 1162
rect 1246 1157 1247 1161
rect 1251 1157 1252 1161
rect 1246 1156 1252 1157
rect 1766 1160 1772 1161
rect 1766 1156 1767 1160
rect 1771 1156 1772 1160
rect 1190 1143 1196 1144
rect 1190 1139 1191 1143
rect 1195 1139 1196 1143
rect 1190 1138 1196 1139
rect 1248 1135 1250 1156
rect 1766 1155 1772 1156
rect 1806 1160 1812 1161
rect 1806 1156 1807 1160
rect 1811 1156 1812 1160
rect 1934 1157 1935 1161
rect 1939 1157 1940 1161
rect 1934 1156 1940 1157
rect 1806 1155 1812 1156
rect 1768 1135 1770 1155
rect 111 1134 115 1135
rect 111 1129 115 1130
rect 135 1134 139 1135
rect 135 1129 139 1130
rect 231 1134 235 1135
rect 231 1129 235 1130
rect 247 1134 251 1135
rect 247 1129 251 1130
rect 359 1134 363 1135
rect 359 1129 363 1130
rect 367 1134 371 1135
rect 367 1129 371 1130
rect 487 1134 491 1135
rect 487 1129 491 1130
rect 495 1134 499 1135
rect 566 1131 567 1135
rect 571 1131 572 1135
rect 566 1130 572 1131
rect 615 1134 619 1135
rect 495 1129 499 1130
rect 615 1129 619 1130
rect 623 1134 627 1135
rect 623 1129 627 1130
rect 743 1134 747 1135
rect 743 1129 747 1130
rect 759 1134 763 1135
rect 838 1131 839 1135
rect 843 1131 844 1135
rect 838 1130 844 1131
rect 871 1134 875 1135
rect 759 1129 763 1130
rect 112 1113 114 1129
rect 110 1112 116 1113
rect 248 1112 250 1129
rect 318 1127 324 1128
rect 318 1123 319 1127
rect 323 1123 324 1127
rect 318 1122 324 1123
rect 110 1108 111 1112
rect 115 1108 116 1112
rect 110 1107 116 1108
rect 246 1111 252 1112
rect 246 1107 247 1111
rect 251 1107 252 1111
rect 246 1106 252 1107
rect 320 1104 322 1122
rect 368 1112 370 1129
rect 438 1127 444 1128
rect 438 1123 439 1127
rect 443 1123 444 1127
rect 438 1122 444 1123
rect 366 1111 372 1112
rect 366 1107 367 1111
rect 371 1107 372 1111
rect 366 1106 372 1107
rect 440 1104 442 1122
rect 496 1112 498 1129
rect 566 1127 572 1128
rect 566 1123 567 1127
rect 571 1123 572 1127
rect 566 1122 572 1123
rect 494 1111 500 1112
rect 494 1107 495 1111
rect 499 1107 500 1111
rect 494 1106 500 1107
rect 568 1104 570 1122
rect 624 1112 626 1129
rect 694 1127 700 1128
rect 694 1123 695 1127
rect 699 1123 700 1127
rect 694 1122 700 1123
rect 622 1111 628 1112
rect 622 1107 623 1111
rect 627 1107 628 1111
rect 622 1106 628 1107
rect 696 1104 698 1122
rect 760 1112 762 1129
rect 758 1111 764 1112
rect 758 1107 759 1111
rect 763 1107 764 1111
rect 758 1106 764 1107
rect 840 1104 842 1130
rect 871 1129 875 1130
rect 887 1134 891 1135
rect 887 1129 891 1130
rect 991 1134 995 1135
rect 991 1129 995 1130
rect 1015 1134 1019 1135
rect 1015 1129 1019 1130
rect 1119 1134 1123 1135
rect 1119 1129 1123 1130
rect 1143 1134 1147 1135
rect 1143 1129 1147 1130
rect 1247 1134 1251 1135
rect 1247 1129 1251 1130
rect 1271 1134 1275 1135
rect 1271 1129 1275 1130
rect 1399 1134 1403 1135
rect 1399 1129 1403 1130
rect 1767 1134 1771 1135
rect 1808 1131 1810 1155
rect 1936 1131 1938 1156
rect 1767 1129 1771 1130
rect 1807 1130 1811 1131
rect 888 1112 890 1129
rect 998 1127 1004 1128
rect 998 1123 999 1127
rect 1003 1123 1004 1127
rect 998 1122 1004 1123
rect 886 1111 892 1112
rect 886 1107 887 1111
rect 891 1107 892 1111
rect 886 1106 892 1107
rect 1000 1104 1002 1122
rect 1016 1112 1018 1129
rect 1110 1127 1116 1128
rect 1110 1123 1111 1127
rect 1115 1123 1116 1127
rect 1110 1122 1116 1123
rect 1014 1111 1020 1112
rect 1014 1107 1015 1111
rect 1019 1107 1020 1111
rect 1014 1106 1020 1107
rect 1112 1104 1114 1122
rect 1144 1112 1146 1129
rect 1222 1127 1228 1128
rect 1222 1123 1223 1127
rect 1227 1123 1228 1127
rect 1222 1122 1228 1123
rect 1142 1111 1148 1112
rect 1142 1107 1143 1111
rect 1147 1107 1148 1111
rect 1142 1106 1148 1107
rect 1224 1104 1226 1122
rect 1272 1112 1274 1129
rect 1350 1127 1356 1128
rect 1350 1123 1351 1127
rect 1355 1123 1356 1127
rect 1350 1122 1356 1123
rect 1382 1127 1388 1128
rect 1382 1123 1383 1127
rect 1387 1123 1388 1127
rect 1382 1122 1388 1123
rect 1270 1111 1276 1112
rect 1270 1107 1271 1111
rect 1275 1107 1276 1111
rect 1270 1106 1276 1107
rect 1352 1104 1354 1122
rect 318 1103 324 1104
rect 318 1099 319 1103
rect 323 1099 324 1103
rect 318 1098 324 1099
rect 438 1103 444 1104
rect 438 1099 439 1103
rect 443 1099 444 1103
rect 438 1098 444 1099
rect 566 1103 572 1104
rect 566 1099 567 1103
rect 571 1099 572 1103
rect 566 1098 572 1099
rect 694 1103 700 1104
rect 694 1099 695 1103
rect 699 1099 700 1103
rect 694 1098 700 1099
rect 702 1103 708 1104
rect 702 1099 703 1103
rect 707 1099 708 1103
rect 702 1098 708 1099
rect 838 1103 844 1104
rect 838 1099 839 1103
rect 843 1099 844 1103
rect 838 1098 844 1099
rect 998 1103 1004 1104
rect 998 1099 999 1103
rect 1003 1099 1004 1103
rect 998 1098 1004 1099
rect 1110 1103 1116 1104
rect 1110 1099 1111 1103
rect 1115 1099 1116 1103
rect 1110 1098 1116 1099
rect 1222 1103 1228 1104
rect 1222 1099 1223 1103
rect 1227 1099 1228 1103
rect 1222 1098 1228 1099
rect 1350 1103 1356 1104
rect 1350 1099 1351 1103
rect 1355 1099 1356 1103
rect 1350 1098 1356 1099
rect 110 1095 116 1096
rect 110 1091 111 1095
rect 115 1091 116 1095
rect 110 1090 116 1091
rect 246 1092 252 1093
rect 112 1067 114 1090
rect 246 1088 247 1092
rect 251 1088 252 1092
rect 246 1087 252 1088
rect 366 1092 372 1093
rect 366 1088 367 1092
rect 371 1088 372 1092
rect 366 1087 372 1088
rect 494 1092 500 1093
rect 494 1088 495 1092
rect 499 1088 500 1092
rect 494 1087 500 1088
rect 622 1092 628 1093
rect 622 1088 623 1092
rect 627 1088 628 1092
rect 622 1087 628 1088
rect 248 1067 250 1087
rect 368 1067 370 1087
rect 496 1067 498 1087
rect 624 1067 626 1087
rect 111 1066 115 1067
rect 111 1061 115 1062
rect 247 1066 251 1067
rect 247 1061 251 1062
rect 367 1066 371 1067
rect 367 1061 371 1062
rect 431 1066 435 1067
rect 431 1061 435 1062
rect 495 1066 499 1067
rect 495 1061 499 1062
rect 543 1066 547 1067
rect 543 1061 547 1062
rect 623 1066 627 1067
rect 623 1061 627 1062
rect 663 1066 667 1067
rect 663 1061 667 1062
rect 112 1042 114 1061
rect 432 1045 434 1061
rect 482 1059 488 1060
rect 482 1055 483 1059
rect 487 1055 488 1059
rect 482 1054 488 1055
rect 430 1044 436 1045
rect 110 1041 116 1042
rect 110 1037 111 1041
rect 115 1037 116 1041
rect 430 1040 431 1044
rect 435 1040 436 1044
rect 430 1039 436 1040
rect 110 1036 116 1037
rect 430 1025 436 1026
rect 110 1024 116 1025
rect 110 1020 111 1024
rect 115 1020 116 1024
rect 430 1021 431 1025
rect 435 1021 436 1025
rect 430 1020 436 1021
rect 110 1019 116 1020
rect 112 995 114 1019
rect 432 995 434 1020
rect 484 1008 486 1054
rect 544 1045 546 1061
rect 664 1045 666 1061
rect 704 1060 706 1098
rect 758 1092 764 1093
rect 758 1088 759 1092
rect 763 1088 764 1092
rect 758 1087 764 1088
rect 886 1092 892 1093
rect 886 1088 887 1092
rect 891 1088 892 1092
rect 886 1087 892 1088
rect 1014 1092 1020 1093
rect 1014 1088 1015 1092
rect 1019 1088 1020 1092
rect 1014 1087 1020 1088
rect 1142 1092 1148 1093
rect 1142 1088 1143 1092
rect 1147 1088 1148 1092
rect 1142 1087 1148 1088
rect 1270 1092 1276 1093
rect 1270 1088 1271 1092
rect 1275 1088 1276 1092
rect 1270 1087 1276 1088
rect 760 1067 762 1087
rect 888 1067 890 1087
rect 1016 1067 1018 1087
rect 1144 1067 1146 1087
rect 1272 1067 1274 1087
rect 759 1066 763 1067
rect 759 1061 763 1062
rect 791 1066 795 1067
rect 791 1061 795 1062
rect 887 1066 891 1067
rect 887 1061 891 1062
rect 919 1066 923 1067
rect 919 1061 923 1062
rect 1015 1066 1019 1067
rect 1015 1061 1019 1062
rect 1039 1066 1043 1067
rect 1039 1061 1043 1062
rect 1143 1066 1147 1067
rect 1143 1061 1147 1062
rect 1159 1066 1163 1067
rect 1159 1061 1163 1062
rect 1271 1066 1275 1067
rect 1271 1061 1275 1062
rect 1279 1066 1283 1067
rect 1279 1061 1283 1062
rect 702 1059 708 1060
rect 702 1055 703 1059
rect 707 1055 708 1059
rect 702 1054 708 1055
rect 792 1045 794 1061
rect 920 1045 922 1061
rect 1040 1045 1042 1061
rect 1090 1051 1096 1052
rect 1090 1047 1091 1051
rect 1095 1047 1096 1051
rect 1090 1046 1096 1047
rect 542 1044 548 1045
rect 542 1040 543 1044
rect 547 1040 548 1044
rect 542 1039 548 1040
rect 662 1044 668 1045
rect 662 1040 663 1044
rect 667 1040 668 1044
rect 662 1039 668 1040
rect 790 1044 796 1045
rect 790 1040 791 1044
rect 795 1040 796 1044
rect 790 1039 796 1040
rect 918 1044 924 1045
rect 918 1040 919 1044
rect 923 1040 924 1044
rect 918 1039 924 1040
rect 1038 1044 1044 1045
rect 1038 1040 1039 1044
rect 1043 1040 1044 1044
rect 1038 1039 1044 1040
rect 502 1035 508 1036
rect 502 1031 503 1035
rect 507 1031 508 1035
rect 502 1030 508 1031
rect 614 1035 620 1036
rect 614 1031 615 1035
rect 619 1031 620 1035
rect 614 1030 620 1031
rect 734 1035 740 1036
rect 734 1031 735 1035
rect 739 1031 740 1035
rect 734 1030 740 1031
rect 862 1035 868 1036
rect 862 1031 863 1035
rect 867 1031 868 1035
rect 862 1030 868 1031
rect 870 1035 876 1036
rect 870 1031 871 1035
rect 875 1031 876 1035
rect 870 1030 876 1031
rect 504 1008 506 1030
rect 542 1025 548 1026
rect 542 1021 543 1025
rect 547 1021 548 1025
rect 542 1020 548 1021
rect 482 1007 488 1008
rect 482 1003 483 1007
rect 487 1003 488 1007
rect 482 1002 488 1003
rect 502 1007 508 1008
rect 502 1003 503 1007
rect 507 1003 508 1007
rect 502 1002 508 1003
rect 544 995 546 1020
rect 616 1008 618 1030
rect 662 1025 668 1026
rect 662 1021 663 1025
rect 667 1021 668 1025
rect 662 1020 668 1021
rect 614 1007 620 1008
rect 614 1003 615 1007
rect 619 1003 620 1007
rect 614 1002 620 1003
rect 664 995 666 1020
rect 736 1008 738 1030
rect 790 1025 796 1026
rect 790 1021 791 1025
rect 795 1021 796 1025
rect 790 1020 796 1021
rect 734 1007 740 1008
rect 734 1003 735 1007
rect 739 1003 740 1007
rect 734 1002 740 1003
rect 792 995 794 1020
rect 864 1008 866 1030
rect 862 1007 868 1008
rect 862 1003 863 1007
rect 867 1003 868 1007
rect 862 1002 868 1003
rect 872 996 874 1030
rect 918 1025 924 1026
rect 918 1021 919 1025
rect 923 1021 924 1025
rect 918 1020 924 1021
rect 1038 1025 1044 1026
rect 1038 1021 1039 1025
rect 1043 1021 1044 1025
rect 1038 1020 1044 1021
rect 870 995 876 996
rect 920 995 922 1020
rect 1040 995 1042 1020
rect 1092 1008 1094 1046
rect 1160 1045 1162 1061
rect 1280 1045 1282 1061
rect 1158 1044 1164 1045
rect 1158 1040 1159 1044
rect 1163 1040 1164 1044
rect 1158 1039 1164 1040
rect 1278 1044 1284 1045
rect 1278 1040 1279 1044
rect 1283 1040 1284 1044
rect 1278 1039 1284 1040
rect 1384 1036 1386 1122
rect 1400 1112 1402 1129
rect 1768 1113 1770 1129
rect 1807 1125 1811 1126
rect 1935 1130 1939 1131
rect 1935 1125 1939 1126
rect 1943 1130 1947 1131
rect 2004 1128 2006 1166
rect 2016 1144 2018 1166
rect 2038 1161 2044 1162
rect 2038 1157 2039 1161
rect 2043 1157 2044 1161
rect 2038 1156 2044 1157
rect 2014 1143 2020 1144
rect 2014 1139 2015 1143
rect 2019 1139 2020 1143
rect 2014 1138 2020 1139
rect 2040 1131 2042 1156
rect 2120 1144 2122 1166
rect 2158 1161 2164 1162
rect 2158 1157 2159 1161
rect 2163 1157 2164 1161
rect 2158 1156 2164 1157
rect 2118 1143 2124 1144
rect 2118 1139 2119 1143
rect 2123 1139 2124 1143
rect 2118 1138 2124 1139
rect 2160 1131 2162 1156
rect 2240 1144 2242 1166
rect 2286 1161 2292 1162
rect 2286 1157 2287 1161
rect 2291 1157 2292 1161
rect 2286 1156 2292 1157
rect 2238 1143 2244 1144
rect 2238 1139 2239 1143
rect 2243 1139 2244 1143
rect 2238 1138 2244 1139
rect 2288 1131 2290 1156
rect 2368 1144 2370 1166
rect 2422 1161 2428 1162
rect 2422 1157 2423 1161
rect 2427 1157 2428 1161
rect 2422 1156 2428 1157
rect 2366 1143 2372 1144
rect 2366 1139 2367 1143
rect 2371 1139 2372 1143
rect 2366 1138 2372 1139
rect 2424 1131 2426 1156
rect 2504 1144 2506 1166
rect 2566 1161 2572 1162
rect 2566 1157 2567 1161
rect 2571 1157 2572 1161
rect 2566 1156 2572 1157
rect 2502 1143 2508 1144
rect 2502 1139 2503 1143
rect 2507 1139 2508 1143
rect 2502 1138 2508 1139
rect 2526 1143 2532 1144
rect 2526 1139 2527 1143
rect 2531 1139 2532 1143
rect 2526 1138 2532 1139
rect 2039 1130 2043 1131
rect 1943 1125 1947 1126
rect 2002 1127 2008 1128
rect 1766 1112 1772 1113
rect 1398 1111 1404 1112
rect 1398 1107 1399 1111
rect 1403 1107 1404 1111
rect 1766 1108 1767 1112
rect 1771 1108 1772 1112
rect 1808 1109 1810 1125
rect 1766 1107 1772 1108
rect 1806 1108 1812 1109
rect 1944 1108 1946 1125
rect 2002 1123 2003 1127
rect 2007 1123 2008 1127
rect 2039 1125 2043 1126
rect 2063 1130 2067 1131
rect 2063 1125 2067 1126
rect 2159 1130 2163 1131
rect 2159 1125 2163 1126
rect 2191 1130 2195 1131
rect 2191 1125 2195 1126
rect 2287 1130 2291 1131
rect 2287 1125 2291 1126
rect 2319 1130 2323 1131
rect 2319 1125 2323 1126
rect 2423 1130 2427 1131
rect 2423 1125 2427 1126
rect 2455 1130 2459 1131
rect 2455 1125 2459 1126
rect 2002 1122 2008 1123
rect 2014 1123 2020 1124
rect 2014 1119 2015 1123
rect 2019 1119 2020 1123
rect 2014 1118 2020 1119
rect 1398 1106 1404 1107
rect 1806 1104 1807 1108
rect 1811 1104 1812 1108
rect 1806 1103 1812 1104
rect 1942 1107 1948 1108
rect 1942 1103 1943 1107
rect 1947 1103 1948 1107
rect 1942 1102 1948 1103
rect 2016 1100 2018 1118
rect 2064 1108 2066 1125
rect 2134 1123 2140 1124
rect 2134 1119 2135 1123
rect 2139 1119 2140 1123
rect 2134 1118 2140 1119
rect 2062 1107 2068 1108
rect 2062 1103 2063 1107
rect 2067 1103 2068 1107
rect 2062 1102 2068 1103
rect 2136 1100 2138 1118
rect 2192 1108 2194 1125
rect 2320 1108 2322 1125
rect 2370 1123 2376 1124
rect 2370 1119 2371 1123
rect 2375 1119 2376 1123
rect 2370 1118 2376 1119
rect 2390 1123 2396 1124
rect 2390 1119 2391 1123
rect 2395 1119 2396 1123
rect 2390 1118 2396 1119
rect 2190 1107 2196 1108
rect 2190 1103 2191 1107
rect 2195 1103 2196 1107
rect 2190 1102 2196 1103
rect 2318 1107 2324 1108
rect 2318 1103 2319 1107
rect 2323 1103 2324 1107
rect 2318 1102 2324 1103
rect 2014 1099 2020 1100
rect 1766 1095 1772 1096
rect 1398 1092 1404 1093
rect 1398 1088 1399 1092
rect 1403 1088 1404 1092
rect 1766 1091 1767 1095
rect 1771 1091 1772 1095
rect 2014 1095 2015 1099
rect 2019 1095 2020 1099
rect 2014 1094 2020 1095
rect 2134 1099 2140 1100
rect 2134 1095 2135 1099
rect 2139 1095 2140 1099
rect 2134 1094 2140 1095
rect 2170 1099 2176 1100
rect 2170 1095 2171 1099
rect 2175 1095 2176 1099
rect 2170 1094 2176 1095
rect 1766 1090 1772 1091
rect 1806 1091 1812 1092
rect 1398 1087 1404 1088
rect 1400 1067 1402 1087
rect 1768 1067 1770 1090
rect 1806 1087 1807 1091
rect 1811 1087 1812 1091
rect 1806 1086 1812 1087
rect 1942 1088 1948 1089
rect 1399 1066 1403 1067
rect 1399 1061 1403 1062
rect 1407 1066 1411 1067
rect 1407 1061 1411 1062
rect 1535 1066 1539 1067
rect 1535 1061 1539 1062
rect 1767 1066 1771 1067
rect 1808 1063 1810 1086
rect 1942 1084 1943 1088
rect 1947 1084 1948 1088
rect 1942 1083 1948 1084
rect 2062 1088 2068 1089
rect 2062 1084 2063 1088
rect 2067 1084 2068 1088
rect 2062 1083 2068 1084
rect 1944 1063 1946 1083
rect 2064 1063 2066 1083
rect 1767 1061 1771 1062
rect 1807 1062 1811 1063
rect 1408 1045 1410 1061
rect 1536 1045 1538 1061
rect 1406 1044 1412 1045
rect 1406 1040 1407 1044
rect 1411 1040 1412 1044
rect 1406 1039 1412 1040
rect 1534 1044 1540 1045
rect 1534 1040 1535 1044
rect 1539 1040 1540 1044
rect 1768 1042 1770 1061
rect 1807 1057 1811 1058
rect 1847 1062 1851 1063
rect 1847 1057 1851 1058
rect 1943 1062 1947 1063
rect 1943 1057 1947 1058
rect 1983 1062 1987 1063
rect 1983 1057 1987 1058
rect 2063 1062 2067 1063
rect 2063 1057 2067 1058
rect 2119 1062 2123 1063
rect 2119 1057 2123 1058
rect 1534 1039 1540 1040
rect 1766 1041 1772 1042
rect 1766 1037 1767 1041
rect 1771 1037 1772 1041
rect 1808 1038 1810 1057
rect 1848 1041 1850 1057
rect 1984 1041 1986 1057
rect 2120 1041 2122 1057
rect 1846 1040 1852 1041
rect 1766 1036 1772 1037
rect 1806 1037 1812 1038
rect 1110 1035 1116 1036
rect 1110 1031 1111 1035
rect 1115 1031 1116 1035
rect 1110 1030 1116 1031
rect 1230 1035 1236 1036
rect 1230 1031 1231 1035
rect 1235 1031 1236 1035
rect 1230 1030 1236 1031
rect 1382 1035 1388 1036
rect 1382 1031 1383 1035
rect 1387 1031 1388 1035
rect 1382 1030 1388 1031
rect 1478 1035 1484 1036
rect 1478 1031 1479 1035
rect 1483 1031 1484 1035
rect 1806 1033 1807 1037
rect 1811 1033 1812 1037
rect 1846 1036 1847 1040
rect 1851 1036 1852 1040
rect 1846 1035 1852 1036
rect 1982 1040 1988 1041
rect 1982 1036 1983 1040
rect 1987 1036 1988 1040
rect 1982 1035 1988 1036
rect 2118 1040 2124 1041
rect 2118 1036 2119 1040
rect 2123 1036 2124 1040
rect 2118 1035 2124 1036
rect 1806 1032 1812 1033
rect 1478 1030 1484 1031
rect 1926 1031 1932 1032
rect 1112 1008 1114 1030
rect 1158 1025 1164 1026
rect 1158 1021 1159 1025
rect 1163 1021 1164 1025
rect 1158 1020 1164 1021
rect 1090 1007 1096 1008
rect 1090 1003 1091 1007
rect 1095 1003 1096 1007
rect 1090 1002 1096 1003
rect 1110 1007 1116 1008
rect 1110 1003 1111 1007
rect 1115 1003 1116 1007
rect 1110 1002 1116 1003
rect 1160 995 1162 1020
rect 1232 1008 1234 1030
rect 1278 1025 1284 1026
rect 1278 1021 1279 1025
rect 1283 1021 1284 1025
rect 1278 1020 1284 1021
rect 1406 1025 1412 1026
rect 1406 1021 1407 1025
rect 1411 1021 1412 1025
rect 1406 1020 1412 1021
rect 1230 1007 1236 1008
rect 1230 1003 1231 1007
rect 1235 1003 1236 1007
rect 1230 1002 1236 1003
rect 1280 995 1282 1020
rect 1408 995 1410 1020
rect 1480 1008 1482 1030
rect 1926 1027 1927 1031
rect 1931 1027 1932 1031
rect 1926 1026 1932 1027
rect 2062 1031 2068 1032
rect 2062 1027 2063 1031
rect 2067 1027 2068 1031
rect 2062 1026 2068 1027
rect 1534 1025 1540 1026
rect 1534 1021 1535 1025
rect 1539 1021 1540 1025
rect 1534 1020 1540 1021
rect 1766 1024 1772 1025
rect 1766 1020 1767 1024
rect 1771 1020 1772 1024
rect 1846 1021 1852 1022
rect 1430 1007 1436 1008
rect 1430 1003 1431 1007
rect 1435 1003 1436 1007
rect 1430 1002 1436 1003
rect 1478 1007 1484 1008
rect 1478 1003 1479 1007
rect 1483 1003 1484 1007
rect 1478 1002 1484 1003
rect 111 994 115 995
rect 111 989 115 990
rect 431 994 435 995
rect 431 989 435 990
rect 543 994 547 995
rect 543 989 547 990
rect 567 994 571 995
rect 567 989 571 990
rect 663 994 667 995
rect 663 989 667 990
rect 679 994 683 995
rect 679 989 683 990
rect 791 994 795 995
rect 870 991 871 995
rect 875 991 876 995
rect 870 990 876 991
rect 911 994 915 995
rect 791 989 795 990
rect 911 989 915 990
rect 919 994 923 995
rect 919 989 923 990
rect 1031 994 1035 995
rect 1031 989 1035 990
rect 1039 994 1043 995
rect 1039 989 1043 990
rect 1143 994 1147 995
rect 1143 989 1147 990
rect 1159 994 1163 995
rect 1159 989 1163 990
rect 1255 994 1259 995
rect 1255 989 1259 990
rect 1279 994 1283 995
rect 1279 989 1283 990
rect 1359 994 1363 995
rect 1359 989 1363 990
rect 1407 994 1411 995
rect 1407 989 1411 990
rect 112 973 114 989
rect 110 972 116 973
rect 568 972 570 989
rect 638 987 644 988
rect 638 983 639 987
rect 643 983 644 987
rect 638 982 644 983
rect 110 968 111 972
rect 115 968 116 972
rect 110 967 116 968
rect 566 971 572 972
rect 566 967 567 971
rect 571 967 572 971
rect 566 966 572 967
rect 640 964 642 982
rect 680 972 682 989
rect 750 987 756 988
rect 750 983 751 987
rect 755 983 756 987
rect 750 982 756 983
rect 678 971 684 972
rect 678 967 679 971
rect 683 967 684 971
rect 678 966 684 967
rect 752 964 754 982
rect 792 972 794 989
rect 862 987 868 988
rect 862 983 863 987
rect 867 983 868 987
rect 862 982 868 983
rect 790 971 796 972
rect 790 967 791 971
rect 795 967 796 971
rect 790 966 796 967
rect 864 964 866 982
rect 912 972 914 989
rect 982 987 988 988
rect 982 983 983 987
rect 987 983 988 987
rect 982 982 988 983
rect 910 971 916 972
rect 910 967 911 971
rect 915 967 916 971
rect 910 966 916 967
rect 984 964 986 982
rect 1032 972 1034 989
rect 1144 972 1146 989
rect 1214 987 1220 988
rect 1214 983 1215 987
rect 1219 983 1220 987
rect 1214 982 1220 983
rect 1030 971 1036 972
rect 1030 967 1031 971
rect 1035 967 1036 971
rect 1030 966 1036 967
rect 1142 971 1148 972
rect 1142 967 1143 971
rect 1147 967 1148 971
rect 1142 966 1148 967
rect 1216 964 1218 982
rect 1256 972 1258 989
rect 1326 987 1332 988
rect 1326 983 1327 987
rect 1331 983 1332 987
rect 1326 982 1332 983
rect 1254 971 1260 972
rect 1254 967 1255 971
rect 1259 967 1260 971
rect 1254 966 1260 967
rect 1328 964 1330 982
rect 1360 972 1362 989
rect 1358 971 1364 972
rect 1358 967 1359 971
rect 1363 967 1364 971
rect 1358 966 1364 967
rect 1432 964 1434 1002
rect 1438 995 1444 996
rect 1536 995 1538 1020
rect 1766 1019 1772 1020
rect 1806 1020 1812 1021
rect 1768 995 1770 1019
rect 1806 1016 1807 1020
rect 1811 1016 1812 1020
rect 1846 1017 1847 1021
rect 1851 1017 1852 1021
rect 1846 1016 1852 1017
rect 1806 1015 1812 1016
rect 1808 995 1810 1015
rect 1848 995 1850 1016
rect 1928 1004 1930 1026
rect 1982 1021 1988 1022
rect 1982 1017 1983 1021
rect 1987 1017 1988 1021
rect 1982 1016 1988 1017
rect 1926 1003 1932 1004
rect 1926 999 1927 1003
rect 1931 999 1932 1003
rect 1926 998 1932 999
rect 1984 995 1986 1016
rect 2064 1004 2066 1026
rect 2118 1021 2124 1022
rect 2118 1017 2119 1021
rect 2123 1017 2124 1021
rect 2118 1016 2124 1017
rect 2062 1003 2068 1004
rect 2062 999 2063 1003
rect 2067 999 2068 1003
rect 2062 998 2068 999
rect 2120 995 2122 1016
rect 2172 1004 2174 1094
rect 2190 1088 2196 1089
rect 2190 1084 2191 1088
rect 2195 1084 2196 1088
rect 2190 1083 2196 1084
rect 2318 1088 2324 1089
rect 2318 1084 2319 1088
rect 2323 1084 2324 1088
rect 2318 1083 2324 1084
rect 2192 1063 2194 1083
rect 2320 1063 2322 1083
rect 2191 1062 2195 1063
rect 2191 1057 2195 1058
rect 2255 1062 2259 1063
rect 2255 1057 2259 1058
rect 2319 1062 2323 1063
rect 2319 1057 2323 1058
rect 2256 1041 2258 1057
rect 2254 1040 2260 1041
rect 2254 1036 2255 1040
rect 2259 1036 2260 1040
rect 2254 1035 2260 1036
rect 2372 1032 2374 1118
rect 2392 1100 2394 1118
rect 2456 1108 2458 1125
rect 2454 1107 2460 1108
rect 2454 1103 2455 1107
rect 2459 1103 2460 1107
rect 2454 1102 2460 1103
rect 2528 1100 2530 1138
rect 2568 1131 2570 1156
rect 2672 1144 2674 1234
rect 2806 1232 2812 1233
rect 2806 1228 2807 1232
rect 2811 1228 2812 1232
rect 2806 1227 2812 1228
rect 3006 1232 3012 1233
rect 3006 1228 3007 1232
rect 3011 1228 3012 1232
rect 3006 1227 3012 1228
rect 2808 1203 2810 1227
rect 3008 1203 3010 1227
rect 2703 1202 2707 1203
rect 2703 1197 2707 1198
rect 2807 1202 2811 1203
rect 2807 1197 2811 1198
rect 2839 1202 2843 1203
rect 2839 1197 2843 1198
rect 2975 1202 2979 1203
rect 2975 1197 2979 1198
rect 3007 1202 3011 1203
rect 3007 1197 3011 1198
rect 2704 1181 2706 1197
rect 2840 1181 2842 1197
rect 2976 1181 2978 1197
rect 2702 1180 2708 1181
rect 2702 1176 2703 1180
rect 2707 1176 2708 1180
rect 2702 1175 2708 1176
rect 2838 1180 2844 1181
rect 2838 1176 2839 1180
rect 2843 1176 2844 1180
rect 2838 1175 2844 1176
rect 2974 1180 2980 1181
rect 2974 1176 2975 1180
rect 2979 1176 2980 1180
rect 2974 1175 2980 1176
rect 3088 1172 3090 1262
rect 3148 1244 3150 1262
rect 3200 1252 3202 1269
rect 3198 1251 3204 1252
rect 3198 1247 3199 1251
rect 3203 1247 3204 1251
rect 3264 1248 3266 1274
rect 3367 1269 3371 1270
rect 3368 1252 3370 1269
rect 3432 1268 3434 1302
rect 3440 1280 3442 1370
rect 3462 1367 3463 1371
rect 3467 1367 3468 1371
rect 3462 1366 3468 1367
rect 3464 1339 3466 1366
rect 3463 1338 3467 1339
rect 3463 1333 3467 1334
rect 3464 1314 3466 1333
rect 3462 1313 3468 1314
rect 3462 1309 3463 1313
rect 3467 1309 3468 1313
rect 3462 1308 3468 1309
rect 3462 1296 3468 1297
rect 3462 1292 3463 1296
rect 3467 1292 3468 1296
rect 3462 1291 3468 1292
rect 3438 1279 3444 1280
rect 3438 1275 3439 1279
rect 3443 1275 3444 1279
rect 3464 1275 3466 1291
rect 3438 1274 3444 1275
rect 3463 1274 3467 1275
rect 3463 1269 3467 1270
rect 3430 1267 3436 1268
rect 3430 1263 3431 1267
rect 3435 1263 3436 1267
rect 3430 1262 3436 1263
rect 3464 1253 3466 1269
rect 3462 1252 3468 1253
rect 3366 1251 3372 1252
rect 3198 1246 3204 1247
rect 3262 1247 3268 1248
rect 3146 1243 3152 1244
rect 3146 1239 3147 1243
rect 3151 1239 3152 1243
rect 3262 1243 3263 1247
rect 3267 1243 3268 1247
rect 3366 1247 3367 1251
rect 3371 1247 3372 1251
rect 3462 1248 3463 1252
rect 3467 1248 3468 1252
rect 3462 1247 3468 1248
rect 3366 1246 3372 1247
rect 3262 1242 3268 1243
rect 3146 1238 3152 1239
rect 3438 1239 3444 1240
rect 3438 1235 3439 1239
rect 3443 1235 3444 1239
rect 3438 1234 3444 1235
rect 3462 1235 3468 1236
rect 3198 1232 3204 1233
rect 3198 1228 3199 1232
rect 3203 1228 3204 1232
rect 3198 1227 3204 1228
rect 3366 1232 3372 1233
rect 3366 1228 3367 1232
rect 3371 1228 3372 1232
rect 3366 1227 3372 1228
rect 3200 1203 3202 1227
rect 3368 1203 3370 1227
rect 3111 1202 3115 1203
rect 3111 1197 3115 1198
rect 3199 1202 3203 1203
rect 3199 1197 3203 1198
rect 3247 1202 3251 1203
rect 3247 1197 3251 1198
rect 3367 1202 3371 1203
rect 3367 1197 3371 1198
rect 3112 1181 3114 1197
rect 3248 1181 3250 1197
rect 3368 1181 3370 1197
rect 3110 1180 3116 1181
rect 3110 1176 3111 1180
rect 3115 1176 3116 1180
rect 3110 1175 3116 1176
rect 3246 1180 3252 1181
rect 3246 1176 3247 1180
rect 3251 1176 3252 1180
rect 3246 1175 3252 1176
rect 3366 1180 3372 1181
rect 3366 1176 3367 1180
rect 3371 1176 3372 1180
rect 3366 1175 3372 1176
rect 2774 1171 2780 1172
rect 2774 1167 2775 1171
rect 2779 1167 2780 1171
rect 2774 1166 2780 1167
rect 2910 1171 2916 1172
rect 2910 1167 2911 1171
rect 2915 1167 2916 1171
rect 2910 1166 2916 1167
rect 3046 1171 3052 1172
rect 3046 1167 3047 1171
rect 3051 1167 3052 1171
rect 3046 1166 3052 1167
rect 3086 1171 3092 1172
rect 3086 1167 3087 1171
rect 3091 1167 3092 1171
rect 3086 1166 3092 1167
rect 3190 1171 3196 1172
rect 3190 1167 3191 1171
rect 3195 1167 3196 1171
rect 3190 1166 3196 1167
rect 3430 1171 3436 1172
rect 3430 1167 3431 1171
rect 3435 1167 3436 1171
rect 3430 1166 3436 1167
rect 2702 1161 2708 1162
rect 2702 1157 2703 1161
rect 2707 1157 2708 1161
rect 2702 1156 2708 1157
rect 2670 1143 2676 1144
rect 2670 1139 2671 1143
rect 2675 1139 2676 1143
rect 2670 1138 2676 1139
rect 2704 1131 2706 1156
rect 2776 1144 2778 1166
rect 2838 1161 2844 1162
rect 2838 1157 2839 1161
rect 2843 1157 2844 1161
rect 2838 1156 2844 1157
rect 2774 1143 2780 1144
rect 2774 1139 2775 1143
rect 2779 1139 2780 1143
rect 2774 1138 2780 1139
rect 2830 1131 2836 1132
rect 2840 1131 2842 1156
rect 2912 1144 2914 1166
rect 2974 1161 2980 1162
rect 2974 1157 2975 1161
rect 2979 1157 2980 1161
rect 2974 1156 2980 1157
rect 2910 1143 2916 1144
rect 2910 1139 2911 1143
rect 2915 1139 2916 1143
rect 2910 1138 2916 1139
rect 2976 1131 2978 1156
rect 2567 1130 2571 1131
rect 2567 1125 2571 1126
rect 2599 1130 2603 1131
rect 2599 1125 2603 1126
rect 2703 1130 2707 1131
rect 2703 1125 2707 1126
rect 2751 1130 2755 1131
rect 2830 1127 2831 1131
rect 2835 1127 2836 1131
rect 2830 1126 2836 1127
rect 2839 1130 2843 1131
rect 2751 1125 2755 1126
rect 2600 1108 2602 1125
rect 2670 1123 2676 1124
rect 2670 1119 2671 1123
rect 2675 1119 2676 1123
rect 2670 1118 2676 1119
rect 2598 1107 2604 1108
rect 2598 1103 2599 1107
rect 2603 1103 2604 1107
rect 2598 1102 2604 1103
rect 2672 1100 2674 1118
rect 2752 1108 2754 1125
rect 2750 1107 2756 1108
rect 2750 1103 2751 1107
rect 2755 1103 2756 1107
rect 2750 1102 2756 1103
rect 2832 1100 2834 1126
rect 2839 1125 2843 1126
rect 2903 1130 2907 1131
rect 2903 1125 2907 1126
rect 2975 1130 2979 1131
rect 2975 1125 2979 1126
rect 2904 1108 2906 1125
rect 3048 1124 3050 1166
rect 3110 1161 3116 1162
rect 3110 1157 3111 1161
rect 3115 1157 3116 1161
rect 3110 1156 3116 1157
rect 3112 1131 3114 1156
rect 3192 1144 3194 1166
rect 3246 1161 3252 1162
rect 3246 1157 3247 1161
rect 3251 1157 3252 1161
rect 3246 1156 3252 1157
rect 3366 1161 3372 1162
rect 3366 1157 3367 1161
rect 3371 1157 3372 1161
rect 3366 1156 3372 1157
rect 3190 1143 3196 1144
rect 3190 1139 3191 1143
rect 3195 1139 3196 1143
rect 3190 1138 3196 1139
rect 3248 1131 3250 1156
rect 3294 1143 3300 1144
rect 3294 1139 3295 1143
rect 3299 1139 3300 1143
rect 3294 1138 3300 1139
rect 3063 1130 3067 1131
rect 3063 1125 3067 1126
rect 3111 1130 3115 1131
rect 3111 1125 3115 1126
rect 3223 1130 3227 1131
rect 3223 1125 3227 1126
rect 3247 1130 3251 1131
rect 3247 1125 3251 1126
rect 2982 1123 2988 1124
rect 2982 1119 2983 1123
rect 2987 1119 2988 1123
rect 2982 1118 2988 1119
rect 3046 1123 3052 1124
rect 3046 1119 3047 1123
rect 3051 1119 3052 1123
rect 3046 1118 3052 1119
rect 2902 1107 2908 1108
rect 2902 1103 2903 1107
rect 2907 1103 2908 1107
rect 2902 1102 2908 1103
rect 2984 1100 2986 1118
rect 3064 1108 3066 1125
rect 3224 1108 3226 1125
rect 3270 1123 3276 1124
rect 3270 1119 3271 1123
rect 3275 1119 3276 1123
rect 3270 1118 3276 1119
rect 3062 1107 3068 1108
rect 3062 1103 3063 1107
rect 3067 1103 3068 1107
rect 3062 1102 3068 1103
rect 3222 1107 3228 1108
rect 3222 1103 3223 1107
rect 3227 1103 3228 1107
rect 3222 1102 3228 1103
rect 2390 1099 2396 1100
rect 2390 1095 2391 1099
rect 2395 1095 2396 1099
rect 2390 1094 2396 1095
rect 2526 1099 2532 1100
rect 2526 1095 2527 1099
rect 2531 1095 2532 1099
rect 2526 1094 2532 1095
rect 2670 1099 2676 1100
rect 2670 1095 2671 1099
rect 2675 1095 2676 1099
rect 2830 1099 2836 1100
rect 2670 1094 2676 1095
rect 2822 1095 2828 1096
rect 2822 1091 2823 1095
rect 2827 1091 2828 1095
rect 2830 1095 2831 1099
rect 2835 1095 2836 1099
rect 2830 1094 2836 1095
rect 2982 1099 2988 1100
rect 2982 1095 2983 1099
rect 2987 1095 2988 1099
rect 2982 1094 2988 1095
rect 2822 1090 2828 1091
rect 2454 1088 2460 1089
rect 2454 1084 2455 1088
rect 2459 1084 2460 1088
rect 2454 1083 2460 1084
rect 2598 1088 2604 1089
rect 2598 1084 2599 1088
rect 2603 1084 2604 1088
rect 2598 1083 2604 1084
rect 2750 1088 2756 1089
rect 2750 1084 2751 1088
rect 2755 1084 2756 1088
rect 2750 1083 2756 1084
rect 2456 1063 2458 1083
rect 2600 1063 2602 1083
rect 2752 1063 2754 1083
rect 2391 1062 2395 1063
rect 2391 1057 2395 1058
rect 2455 1062 2459 1063
rect 2455 1057 2459 1058
rect 2543 1062 2547 1063
rect 2543 1057 2547 1058
rect 2599 1062 2603 1063
rect 2599 1057 2603 1058
rect 2703 1062 2707 1063
rect 2703 1057 2707 1058
rect 2751 1062 2755 1063
rect 2751 1057 2755 1058
rect 2392 1041 2394 1057
rect 2544 1041 2546 1057
rect 2594 1047 2600 1048
rect 2594 1043 2595 1047
rect 2599 1043 2600 1047
rect 2594 1042 2600 1043
rect 2390 1040 2396 1041
rect 2390 1036 2391 1040
rect 2395 1036 2396 1040
rect 2390 1035 2396 1036
rect 2542 1040 2548 1041
rect 2542 1036 2543 1040
rect 2547 1036 2548 1040
rect 2542 1035 2548 1036
rect 2370 1031 2376 1032
rect 2370 1027 2371 1031
rect 2375 1027 2376 1031
rect 2370 1026 2376 1027
rect 2254 1021 2260 1022
rect 2254 1017 2255 1021
rect 2259 1017 2260 1021
rect 2254 1016 2260 1017
rect 2390 1021 2396 1022
rect 2390 1017 2391 1021
rect 2395 1017 2396 1021
rect 2390 1016 2396 1017
rect 2542 1021 2548 1022
rect 2542 1017 2543 1021
rect 2547 1017 2548 1021
rect 2542 1016 2548 1017
rect 2170 1003 2176 1004
rect 2170 999 2171 1003
rect 2175 999 2176 1003
rect 2170 998 2176 999
rect 2256 995 2258 1016
rect 2366 1003 2372 1004
rect 2366 999 2367 1003
rect 2371 999 2372 1003
rect 2366 998 2372 999
rect 1438 991 1439 995
rect 1443 991 1444 995
rect 1438 990 1444 991
rect 1471 994 1475 995
rect 1440 964 1442 990
rect 1471 989 1475 990
rect 1535 994 1539 995
rect 1535 989 1539 990
rect 1583 994 1587 995
rect 1583 989 1587 990
rect 1671 994 1675 995
rect 1671 989 1675 990
rect 1767 994 1771 995
rect 1767 989 1771 990
rect 1807 994 1811 995
rect 1807 989 1811 990
rect 1831 994 1835 995
rect 1831 989 1835 990
rect 1847 994 1851 995
rect 1847 989 1851 990
rect 1975 994 1979 995
rect 1975 989 1979 990
rect 1983 994 1987 995
rect 1983 989 1987 990
rect 2119 994 2123 995
rect 2119 989 2123 990
rect 2135 994 2139 995
rect 2135 989 2139 990
rect 2255 994 2259 995
rect 2255 989 2259 990
rect 2295 994 2299 995
rect 2295 989 2299 990
rect 1472 972 1474 989
rect 1522 987 1528 988
rect 1522 983 1523 987
rect 1527 983 1528 987
rect 1522 982 1528 983
rect 1470 971 1476 972
rect 1470 967 1471 971
rect 1475 967 1476 971
rect 1470 966 1476 967
rect 638 963 644 964
rect 638 959 639 963
rect 643 959 644 963
rect 638 958 644 959
rect 750 963 756 964
rect 750 959 751 963
rect 755 959 756 963
rect 750 958 756 959
rect 862 963 868 964
rect 862 959 863 963
rect 867 959 868 963
rect 862 958 868 959
rect 982 963 988 964
rect 982 959 983 963
rect 987 959 988 963
rect 982 958 988 959
rect 990 963 996 964
rect 990 959 991 963
rect 995 959 996 963
rect 990 958 996 959
rect 1214 963 1220 964
rect 1214 959 1215 963
rect 1219 959 1220 963
rect 1214 958 1220 959
rect 1326 963 1332 964
rect 1326 959 1327 963
rect 1331 959 1332 963
rect 1326 958 1332 959
rect 1430 963 1436 964
rect 1430 959 1431 963
rect 1435 959 1436 963
rect 1430 958 1436 959
rect 1438 963 1444 964
rect 1438 959 1439 963
rect 1443 959 1444 963
rect 1438 958 1444 959
rect 110 955 116 956
rect 110 951 111 955
rect 115 951 116 955
rect 110 950 116 951
rect 566 952 572 953
rect 112 927 114 950
rect 566 948 567 952
rect 571 948 572 952
rect 566 947 572 948
rect 678 952 684 953
rect 678 948 679 952
rect 683 948 684 952
rect 678 947 684 948
rect 790 952 796 953
rect 790 948 791 952
rect 795 948 796 952
rect 790 947 796 948
rect 910 952 916 953
rect 910 948 911 952
rect 915 948 916 952
rect 910 947 916 948
rect 568 927 570 947
rect 680 927 682 947
rect 792 927 794 947
rect 912 927 914 947
rect 111 926 115 927
rect 111 921 115 922
rect 415 926 419 927
rect 415 921 419 922
rect 559 926 563 927
rect 559 921 563 922
rect 567 926 571 927
rect 567 921 571 922
rect 679 926 683 927
rect 679 921 683 922
rect 727 926 731 927
rect 727 921 731 922
rect 791 926 795 927
rect 791 921 795 922
rect 911 926 915 927
rect 911 921 915 922
rect 112 902 114 921
rect 416 905 418 921
rect 560 905 562 921
rect 728 905 730 921
rect 912 905 914 921
rect 414 904 420 905
rect 110 901 116 902
rect 110 897 111 901
rect 115 897 116 901
rect 414 900 415 904
rect 419 900 420 904
rect 414 899 420 900
rect 558 904 564 905
rect 558 900 559 904
rect 563 900 564 904
rect 558 899 564 900
rect 726 904 732 905
rect 726 900 727 904
rect 731 900 732 904
rect 726 899 732 900
rect 910 904 916 905
rect 910 900 911 904
rect 915 900 916 904
rect 910 899 916 900
rect 110 896 116 897
rect 486 895 492 896
rect 486 891 487 895
rect 491 891 492 895
rect 486 890 492 891
rect 630 895 636 896
rect 630 891 631 895
rect 635 891 636 895
rect 630 890 636 891
rect 678 895 684 896
rect 678 891 679 895
rect 683 891 684 895
rect 678 890 684 891
rect 806 895 812 896
rect 806 891 807 895
rect 811 891 812 895
rect 806 890 812 891
rect 414 885 420 886
rect 110 884 116 885
rect 110 880 111 884
rect 115 880 116 884
rect 414 881 415 885
rect 419 881 420 885
rect 414 880 420 881
rect 110 879 116 880
rect 112 859 114 879
rect 416 859 418 880
rect 488 868 490 890
rect 558 885 564 886
rect 558 881 559 885
rect 563 881 564 885
rect 558 880 564 881
rect 486 867 492 868
rect 486 863 487 867
rect 491 863 492 867
rect 486 862 492 863
rect 560 859 562 880
rect 111 858 115 859
rect 111 853 115 854
rect 135 858 139 859
rect 135 853 139 854
rect 231 858 235 859
rect 231 853 235 854
rect 359 858 363 859
rect 359 853 363 854
rect 415 858 419 859
rect 415 853 419 854
rect 487 858 491 859
rect 487 853 491 854
rect 559 858 563 859
rect 559 853 563 854
rect 623 858 627 859
rect 623 853 627 854
rect 112 837 114 853
rect 110 836 116 837
rect 136 836 138 853
rect 214 851 220 852
rect 214 847 215 851
rect 219 847 220 851
rect 214 846 220 847
rect 110 832 111 836
rect 115 832 116 836
rect 110 831 116 832
rect 134 835 140 836
rect 134 831 135 835
rect 139 831 140 835
rect 134 830 140 831
rect 216 828 218 846
rect 232 836 234 853
rect 310 851 316 852
rect 310 847 311 851
rect 315 847 316 851
rect 310 846 316 847
rect 230 835 236 836
rect 230 831 231 835
rect 235 831 236 835
rect 230 830 236 831
rect 312 828 314 846
rect 360 836 362 853
rect 488 836 490 853
rect 624 836 626 853
rect 632 852 634 890
rect 680 860 682 890
rect 726 885 732 886
rect 726 881 727 885
rect 731 881 732 885
rect 726 880 732 881
rect 678 859 684 860
rect 728 859 730 880
rect 808 868 810 890
rect 910 885 916 886
rect 910 881 911 885
rect 915 881 916 885
rect 910 880 916 881
rect 806 867 812 868
rect 806 863 807 867
rect 811 863 812 867
rect 806 862 812 863
rect 912 859 914 880
rect 992 868 994 958
rect 1030 952 1036 953
rect 1030 948 1031 952
rect 1035 948 1036 952
rect 1030 947 1036 948
rect 1142 952 1148 953
rect 1142 948 1143 952
rect 1147 948 1148 952
rect 1142 947 1148 948
rect 1254 952 1260 953
rect 1254 948 1255 952
rect 1259 948 1260 952
rect 1254 947 1260 948
rect 1358 952 1364 953
rect 1358 948 1359 952
rect 1363 948 1364 952
rect 1358 947 1364 948
rect 1470 952 1476 953
rect 1470 948 1471 952
rect 1475 948 1476 952
rect 1470 947 1476 948
rect 1032 927 1034 947
rect 1144 927 1146 947
rect 1256 927 1258 947
rect 1360 927 1362 947
rect 1472 927 1474 947
rect 1031 926 1035 927
rect 1031 921 1035 922
rect 1119 926 1123 927
rect 1119 921 1123 922
rect 1143 926 1147 927
rect 1143 921 1147 922
rect 1255 926 1259 927
rect 1255 921 1259 922
rect 1335 926 1339 927
rect 1335 921 1339 922
rect 1359 926 1363 927
rect 1359 921 1363 922
rect 1471 926 1475 927
rect 1471 921 1475 922
rect 1120 905 1122 921
rect 1336 905 1338 921
rect 1118 904 1124 905
rect 1118 900 1119 904
rect 1123 900 1124 904
rect 1118 899 1124 900
rect 1334 904 1340 905
rect 1334 900 1335 904
rect 1339 900 1340 904
rect 1334 899 1340 900
rect 1524 896 1526 982
rect 1584 972 1586 989
rect 1662 987 1668 988
rect 1662 983 1663 987
rect 1667 983 1668 987
rect 1662 982 1668 983
rect 1582 971 1588 972
rect 1582 967 1583 971
rect 1587 967 1588 971
rect 1582 966 1588 967
rect 1664 964 1666 982
rect 1672 972 1674 989
rect 1750 987 1756 988
rect 1750 983 1751 987
rect 1755 983 1756 987
rect 1750 982 1756 983
rect 1670 971 1676 972
rect 1670 967 1671 971
rect 1675 967 1676 971
rect 1670 966 1676 967
rect 1752 964 1754 982
rect 1768 973 1770 989
rect 1808 973 1810 989
rect 1766 972 1772 973
rect 1766 968 1767 972
rect 1771 968 1772 972
rect 1766 967 1772 968
rect 1806 972 1812 973
rect 1832 972 1834 989
rect 1938 987 1944 988
rect 1938 983 1939 987
rect 1943 983 1944 987
rect 1938 982 1944 983
rect 1806 968 1807 972
rect 1811 968 1812 972
rect 1806 967 1812 968
rect 1830 971 1836 972
rect 1830 967 1831 971
rect 1835 967 1836 971
rect 1830 966 1836 967
rect 1940 964 1942 982
rect 1976 972 1978 989
rect 2136 972 2138 989
rect 2296 972 2298 989
rect 1974 971 1980 972
rect 1974 967 1975 971
rect 1979 967 1980 971
rect 1974 966 1980 967
rect 2134 971 2140 972
rect 2134 967 2135 971
rect 2139 967 2140 971
rect 2134 966 2140 967
rect 2294 971 2300 972
rect 2294 967 2295 971
rect 2299 967 2300 971
rect 2294 966 2300 967
rect 2368 964 2370 998
rect 2392 995 2394 1016
rect 2418 995 2424 996
rect 2544 995 2546 1016
rect 2596 1004 2598 1042
rect 2704 1041 2706 1057
rect 2702 1040 2708 1041
rect 2702 1036 2703 1040
rect 2707 1036 2708 1040
rect 2702 1035 2708 1036
rect 2614 1031 2620 1032
rect 2614 1027 2615 1031
rect 2619 1027 2620 1031
rect 2614 1026 2620 1027
rect 2774 1031 2780 1032
rect 2774 1027 2775 1031
rect 2779 1027 2780 1031
rect 2774 1026 2780 1027
rect 2616 1004 2618 1026
rect 2702 1021 2708 1022
rect 2702 1017 2703 1021
rect 2707 1017 2708 1021
rect 2702 1016 2708 1017
rect 2594 1003 2600 1004
rect 2594 999 2595 1003
rect 2599 999 2600 1003
rect 2594 998 2600 999
rect 2614 1003 2620 1004
rect 2614 999 2615 1003
rect 2619 999 2620 1003
rect 2614 998 2620 999
rect 2704 995 2706 1016
rect 2391 994 2395 995
rect 2418 991 2419 995
rect 2423 991 2424 995
rect 2418 990 2424 991
rect 2463 994 2467 995
rect 2391 989 2395 990
rect 2420 964 2422 990
rect 2463 989 2467 990
rect 2543 994 2547 995
rect 2543 989 2547 990
rect 2631 994 2635 995
rect 2631 989 2635 990
rect 2703 994 2707 995
rect 2703 989 2707 990
rect 2464 972 2466 989
rect 2470 987 2476 988
rect 2470 983 2471 987
rect 2475 983 2476 987
rect 2470 982 2476 983
rect 2462 971 2468 972
rect 2462 967 2463 971
rect 2467 967 2468 971
rect 2462 966 2468 967
rect 1662 963 1668 964
rect 1654 959 1660 960
rect 1654 955 1655 959
rect 1659 955 1660 959
rect 1662 959 1663 963
rect 1667 959 1668 963
rect 1662 958 1668 959
rect 1750 963 1756 964
rect 1750 959 1751 963
rect 1755 959 1756 963
rect 1750 958 1756 959
rect 1938 963 1944 964
rect 1938 959 1939 963
rect 1943 959 1944 963
rect 2366 963 2372 964
rect 1938 958 1944 959
rect 2206 959 2212 960
rect 1654 954 1660 955
rect 1766 955 1772 956
rect 1582 952 1588 953
rect 1582 948 1583 952
rect 1587 948 1588 952
rect 1582 947 1588 948
rect 1584 927 1586 947
rect 1559 926 1563 927
rect 1559 921 1563 922
rect 1583 926 1587 927
rect 1583 921 1587 922
rect 1560 905 1562 921
rect 1558 904 1564 905
rect 1558 900 1559 904
rect 1563 900 1564 904
rect 1558 899 1564 900
rect 1190 895 1196 896
rect 1190 891 1191 895
rect 1195 891 1196 895
rect 1190 890 1196 891
rect 1322 895 1328 896
rect 1322 891 1323 895
rect 1327 891 1328 895
rect 1322 890 1328 891
rect 1522 895 1528 896
rect 1522 891 1523 895
rect 1527 891 1528 895
rect 1522 890 1528 891
rect 1118 885 1124 886
rect 1118 881 1119 885
rect 1123 881 1124 885
rect 1118 880 1124 881
rect 990 867 996 868
rect 990 863 991 867
rect 995 863 996 867
rect 990 862 996 863
rect 1120 859 1122 880
rect 1192 868 1194 890
rect 1190 867 1196 868
rect 1190 863 1191 867
rect 1195 863 1196 867
rect 1190 862 1196 863
rect 1230 859 1236 860
rect 678 855 679 859
rect 683 855 684 859
rect 678 854 684 855
rect 727 858 731 859
rect 727 853 731 854
rect 751 858 755 859
rect 751 853 755 854
rect 879 858 883 859
rect 879 853 883 854
rect 911 858 915 859
rect 911 853 915 854
rect 1007 858 1011 859
rect 1007 853 1011 854
rect 1119 858 1123 859
rect 1119 853 1123 854
rect 1135 858 1139 859
rect 1230 855 1231 859
rect 1235 855 1236 859
rect 1230 854 1236 855
rect 1271 858 1275 859
rect 1135 853 1139 854
rect 630 851 636 852
rect 630 847 631 851
rect 635 847 636 851
rect 630 846 636 847
rect 752 836 754 853
rect 798 851 804 852
rect 798 847 799 851
rect 803 850 804 851
rect 822 851 828 852
rect 803 848 810 850
rect 803 847 804 848
rect 798 846 804 847
rect 358 835 364 836
rect 358 831 359 835
rect 363 831 364 835
rect 358 830 364 831
rect 486 835 492 836
rect 486 831 487 835
rect 491 831 492 835
rect 486 830 492 831
rect 622 835 628 836
rect 622 831 623 835
rect 627 831 628 835
rect 622 830 628 831
rect 750 835 756 836
rect 750 831 751 835
rect 755 831 756 835
rect 750 830 756 831
rect 214 827 220 828
rect 214 823 215 827
rect 219 823 220 827
rect 214 822 220 823
rect 310 827 316 828
rect 310 823 311 827
rect 315 823 316 827
rect 310 822 316 823
rect 110 819 116 820
rect 110 815 111 819
rect 115 815 116 819
rect 198 819 204 820
rect 110 814 116 815
rect 134 816 140 817
rect 112 791 114 814
rect 134 812 135 816
rect 139 812 140 816
rect 198 815 199 819
rect 203 815 204 819
rect 198 814 204 815
rect 230 816 236 817
rect 134 811 140 812
rect 136 791 138 811
rect 111 790 115 791
rect 111 785 115 786
rect 135 790 139 791
rect 135 785 139 786
rect 112 766 114 785
rect 136 769 138 785
rect 134 768 140 769
rect 110 765 116 766
rect 110 761 111 765
rect 115 761 116 765
rect 134 764 135 768
rect 139 764 140 768
rect 134 763 140 764
rect 110 760 116 761
rect 134 749 140 750
rect 110 748 116 749
rect 110 744 111 748
rect 115 744 116 748
rect 134 745 135 749
rect 139 745 140 749
rect 134 744 140 745
rect 110 743 116 744
rect 112 723 114 743
rect 136 723 138 744
rect 200 732 202 814
rect 230 812 231 816
rect 235 812 236 816
rect 230 811 236 812
rect 358 816 364 817
rect 358 812 359 816
rect 363 812 364 816
rect 358 811 364 812
rect 486 816 492 817
rect 486 812 487 816
rect 491 812 492 816
rect 486 811 492 812
rect 622 816 628 817
rect 622 812 623 816
rect 627 812 628 816
rect 622 811 628 812
rect 750 816 756 817
rect 750 812 751 816
rect 755 812 756 816
rect 750 811 756 812
rect 232 791 234 811
rect 360 791 362 811
rect 488 791 490 811
rect 624 791 626 811
rect 752 791 754 811
rect 223 790 227 791
rect 223 785 227 786
rect 231 790 235 791
rect 231 785 235 786
rect 343 790 347 791
rect 343 785 347 786
rect 359 790 363 791
rect 359 785 363 786
rect 471 790 475 791
rect 471 785 475 786
rect 487 790 491 791
rect 487 785 491 786
rect 607 790 611 791
rect 607 785 611 786
rect 623 790 627 791
rect 623 785 627 786
rect 743 790 747 791
rect 743 785 747 786
rect 751 790 755 791
rect 751 785 755 786
rect 224 769 226 785
rect 344 769 346 785
rect 472 769 474 785
rect 608 769 610 785
rect 744 769 746 785
rect 222 768 228 769
rect 222 764 223 768
rect 227 764 228 768
rect 222 763 228 764
rect 342 768 348 769
rect 342 764 343 768
rect 347 764 348 768
rect 342 763 348 764
rect 470 768 476 769
rect 470 764 471 768
rect 475 764 476 768
rect 470 763 476 764
rect 606 768 612 769
rect 606 764 607 768
rect 611 764 612 768
rect 606 763 612 764
rect 742 768 748 769
rect 742 764 743 768
rect 747 764 748 768
rect 742 763 748 764
rect 808 760 810 848
rect 822 847 823 851
rect 827 847 828 851
rect 822 846 828 847
rect 824 828 826 846
rect 880 836 882 853
rect 1008 836 1010 853
rect 1114 847 1120 848
rect 1114 843 1115 847
rect 1119 843 1120 847
rect 1114 842 1120 843
rect 878 835 884 836
rect 878 831 879 835
rect 883 831 884 835
rect 878 830 884 831
rect 1006 835 1012 836
rect 1006 831 1007 835
rect 1011 831 1012 835
rect 1006 830 1012 831
rect 1116 828 1118 842
rect 1136 836 1138 853
rect 1134 835 1140 836
rect 1134 831 1135 835
rect 1139 831 1140 835
rect 1134 830 1140 831
rect 1232 828 1234 854
rect 1271 853 1275 854
rect 1272 836 1274 853
rect 1324 852 1326 890
rect 1334 885 1340 886
rect 1334 881 1335 885
rect 1339 881 1340 885
rect 1334 880 1340 881
rect 1558 885 1564 886
rect 1558 881 1559 885
rect 1563 881 1564 885
rect 1558 880 1564 881
rect 1336 859 1338 880
rect 1560 859 1562 880
rect 1656 868 1658 954
rect 1670 952 1676 953
rect 1670 948 1671 952
rect 1675 948 1676 952
rect 1766 951 1767 955
rect 1771 951 1772 955
rect 1766 950 1772 951
rect 1806 955 1812 956
rect 1806 951 1807 955
rect 1811 951 1812 955
rect 2206 955 2207 959
rect 2211 955 2212 959
rect 2366 959 2367 963
rect 2371 959 2372 963
rect 2366 958 2372 959
rect 2418 963 2424 964
rect 2418 959 2419 963
rect 2423 959 2424 963
rect 2418 958 2424 959
rect 2206 954 2212 955
rect 1806 950 1812 951
rect 1830 952 1836 953
rect 1670 947 1676 948
rect 1672 927 1674 947
rect 1768 927 1770 950
rect 1808 931 1810 950
rect 1830 948 1831 952
rect 1835 948 1836 952
rect 1830 947 1836 948
rect 1974 952 1980 953
rect 1974 948 1975 952
rect 1979 948 1980 952
rect 1974 947 1980 948
rect 2134 952 2140 953
rect 2134 948 2135 952
rect 2139 948 2140 952
rect 2134 947 2140 948
rect 1832 931 1834 947
rect 1976 931 1978 947
rect 2136 931 2138 947
rect 1807 930 1811 931
rect 1671 926 1675 927
rect 1671 921 1675 922
rect 1767 926 1771 927
rect 1807 925 1811 926
rect 1831 930 1835 931
rect 1831 925 1835 926
rect 1975 930 1979 931
rect 1975 925 1979 926
rect 2127 930 2131 931
rect 2127 925 2131 926
rect 2135 930 2139 931
rect 2135 925 2139 926
rect 1767 921 1771 922
rect 1768 902 1770 921
rect 1808 906 1810 925
rect 2128 909 2130 925
rect 2126 908 2132 909
rect 1806 905 1812 906
rect 1766 901 1772 902
rect 1766 897 1767 901
rect 1771 897 1772 901
rect 1806 901 1807 905
rect 1811 901 1812 905
rect 2126 904 2127 908
rect 2131 904 2132 908
rect 2126 903 2132 904
rect 1806 900 1812 901
rect 1766 896 1772 897
rect 2126 889 2132 890
rect 1806 888 1812 889
rect 1766 884 1772 885
rect 1766 880 1767 884
rect 1771 880 1772 884
rect 1806 884 1807 888
rect 1811 884 1812 888
rect 2126 885 2127 889
rect 2131 885 2132 889
rect 2126 884 2132 885
rect 1806 883 1812 884
rect 1766 879 1772 880
rect 1654 867 1660 868
rect 1654 863 1655 867
rect 1659 863 1660 867
rect 1654 862 1660 863
rect 1768 859 1770 879
rect 1808 859 1810 883
rect 2128 859 2130 884
rect 2208 872 2210 954
rect 2294 952 2300 953
rect 2294 948 2295 952
rect 2299 948 2300 952
rect 2294 947 2300 948
rect 2462 952 2468 953
rect 2462 948 2463 952
rect 2467 948 2468 952
rect 2462 947 2468 948
rect 2296 931 2298 947
rect 2464 931 2466 947
rect 2215 930 2219 931
rect 2215 925 2219 926
rect 2295 930 2299 931
rect 2295 925 2299 926
rect 2303 930 2307 931
rect 2303 925 2307 926
rect 2391 930 2395 931
rect 2391 925 2395 926
rect 2463 930 2467 931
rect 2463 925 2467 926
rect 2216 909 2218 925
rect 2304 909 2306 925
rect 2392 909 2394 925
rect 2214 908 2220 909
rect 2214 904 2215 908
rect 2219 904 2220 908
rect 2214 903 2220 904
rect 2302 908 2308 909
rect 2302 904 2303 908
rect 2307 904 2308 908
rect 2302 903 2308 904
rect 2390 908 2396 909
rect 2390 904 2391 908
rect 2395 904 2396 908
rect 2390 903 2396 904
rect 2472 900 2474 982
rect 2632 972 2634 989
rect 2776 984 2778 1026
rect 2824 1004 2826 1090
rect 2902 1088 2908 1089
rect 2902 1084 2903 1088
rect 2907 1084 2908 1088
rect 2902 1083 2908 1084
rect 3062 1088 3068 1089
rect 3062 1084 3063 1088
rect 3067 1084 3068 1088
rect 3062 1083 3068 1084
rect 3222 1088 3228 1089
rect 3222 1084 3223 1088
rect 3227 1084 3228 1088
rect 3222 1083 3228 1084
rect 2904 1063 2906 1083
rect 3064 1063 3066 1083
rect 3224 1063 3226 1083
rect 2863 1062 2867 1063
rect 2863 1057 2867 1058
rect 2903 1062 2907 1063
rect 2903 1057 2907 1058
rect 3031 1062 3035 1063
rect 3031 1057 3035 1058
rect 3063 1062 3067 1063
rect 3063 1057 3067 1058
rect 3207 1062 3211 1063
rect 3207 1057 3211 1058
rect 3223 1062 3227 1063
rect 3223 1057 3227 1058
rect 2864 1041 2866 1057
rect 3032 1041 3034 1057
rect 3208 1041 3210 1057
rect 2862 1040 2868 1041
rect 2862 1036 2863 1040
rect 2867 1036 2868 1040
rect 2862 1035 2868 1036
rect 3030 1040 3036 1041
rect 3030 1036 3031 1040
rect 3035 1036 3036 1040
rect 3030 1035 3036 1036
rect 3206 1040 3212 1041
rect 3206 1036 3207 1040
rect 3211 1036 3212 1040
rect 3206 1035 3212 1036
rect 3272 1032 3274 1118
rect 3296 1100 3298 1138
rect 3368 1131 3370 1156
rect 3367 1130 3371 1131
rect 3367 1125 3371 1126
rect 3368 1108 3370 1125
rect 3432 1124 3434 1166
rect 3440 1144 3442 1234
rect 3462 1231 3463 1235
rect 3467 1231 3468 1235
rect 3462 1230 3468 1231
rect 3464 1203 3466 1230
rect 3463 1202 3467 1203
rect 3463 1197 3467 1198
rect 3464 1178 3466 1197
rect 3462 1177 3468 1178
rect 3462 1173 3463 1177
rect 3467 1173 3468 1177
rect 3462 1172 3468 1173
rect 3462 1160 3468 1161
rect 3462 1156 3463 1160
rect 3467 1156 3468 1160
rect 3462 1155 3468 1156
rect 3438 1143 3444 1144
rect 3438 1139 3439 1143
rect 3443 1139 3444 1143
rect 3438 1138 3444 1139
rect 3464 1131 3466 1155
rect 3463 1130 3467 1131
rect 3463 1125 3467 1126
rect 3430 1123 3436 1124
rect 3430 1119 3431 1123
rect 3435 1119 3436 1123
rect 3430 1118 3436 1119
rect 3464 1109 3466 1125
rect 3462 1108 3468 1109
rect 3366 1107 3372 1108
rect 3366 1103 3367 1107
rect 3371 1103 3372 1107
rect 3462 1104 3463 1108
rect 3467 1104 3468 1108
rect 3462 1103 3468 1104
rect 3366 1102 3372 1103
rect 3294 1099 3300 1100
rect 3294 1095 3295 1099
rect 3299 1095 3300 1099
rect 3294 1094 3300 1095
rect 3438 1095 3444 1096
rect 3438 1091 3439 1095
rect 3443 1091 3444 1095
rect 3438 1090 3444 1091
rect 3462 1091 3468 1092
rect 3366 1088 3372 1089
rect 3366 1084 3367 1088
rect 3371 1084 3372 1088
rect 3366 1083 3372 1084
rect 3368 1063 3370 1083
rect 3367 1062 3371 1063
rect 3367 1057 3371 1058
rect 3368 1041 3370 1057
rect 3366 1040 3372 1041
rect 3366 1036 3367 1040
rect 3371 1036 3372 1040
rect 3366 1035 3372 1036
rect 2934 1031 2940 1032
rect 2934 1027 2935 1031
rect 2939 1027 2940 1031
rect 2934 1026 2940 1027
rect 3270 1031 3276 1032
rect 3270 1027 3271 1031
rect 3275 1027 3276 1031
rect 3270 1026 3276 1027
rect 3430 1031 3436 1032
rect 3430 1027 3431 1031
rect 3435 1027 3436 1031
rect 3430 1026 3436 1027
rect 2862 1021 2868 1022
rect 2862 1017 2863 1021
rect 2867 1017 2868 1021
rect 2862 1016 2868 1017
rect 2822 1003 2828 1004
rect 2822 999 2823 1003
rect 2827 999 2828 1003
rect 2822 998 2828 999
rect 2864 995 2866 1016
rect 2936 1004 2938 1026
rect 3030 1021 3036 1022
rect 3030 1017 3031 1021
rect 3035 1017 3036 1021
rect 3030 1016 3036 1017
rect 3206 1021 3212 1022
rect 3206 1017 3207 1021
rect 3211 1017 3212 1021
rect 3206 1016 3212 1017
rect 3366 1021 3372 1022
rect 3366 1017 3367 1021
rect 3371 1017 3372 1021
rect 3366 1016 3372 1017
rect 2934 1003 2940 1004
rect 2934 999 2935 1003
rect 2939 999 2940 1003
rect 2934 998 2940 999
rect 2958 995 2964 996
rect 3032 995 3034 1016
rect 3208 995 3210 1016
rect 3254 1003 3260 1004
rect 3254 999 3255 1003
rect 3259 999 3260 1003
rect 3254 998 3260 999
rect 2807 994 2811 995
rect 2807 989 2811 990
rect 2863 994 2867 995
rect 2958 991 2959 995
rect 2963 991 2964 995
rect 2958 990 2964 991
rect 2991 994 2995 995
rect 2863 989 2867 990
rect 2774 983 2780 984
rect 2774 979 2775 983
rect 2779 979 2780 983
rect 2774 978 2780 979
rect 2808 972 2810 989
rect 2878 987 2884 988
rect 2878 983 2879 987
rect 2883 983 2884 987
rect 2878 982 2884 983
rect 2630 971 2636 972
rect 2630 967 2631 971
rect 2635 967 2636 971
rect 2630 966 2636 967
rect 2806 971 2812 972
rect 2806 967 2807 971
rect 2811 967 2812 971
rect 2806 966 2812 967
rect 2880 964 2882 982
rect 2960 964 2962 990
rect 2991 989 2995 990
rect 3031 994 3035 995
rect 3031 989 3035 990
rect 3183 994 3187 995
rect 3183 989 3187 990
rect 3207 994 3211 995
rect 3207 989 3211 990
rect 2992 972 2994 989
rect 3184 972 3186 989
rect 2990 971 2996 972
rect 2990 967 2991 971
rect 2995 967 2996 971
rect 2990 966 2996 967
rect 3182 971 3188 972
rect 3182 967 3183 971
rect 3187 967 3188 971
rect 3182 966 3188 967
rect 3256 964 3258 998
rect 3368 995 3370 1016
rect 3367 994 3371 995
rect 3367 989 3371 990
rect 3294 987 3300 988
rect 3294 983 3295 987
rect 3299 983 3300 987
rect 3294 982 3300 983
rect 2878 963 2884 964
rect 2878 959 2879 963
rect 2883 959 2884 963
rect 2878 958 2884 959
rect 2958 963 2964 964
rect 2958 959 2959 963
rect 2963 959 2964 963
rect 2958 958 2964 959
rect 3254 963 3260 964
rect 3254 959 3255 963
rect 3259 959 3260 963
rect 3254 958 3260 959
rect 2630 952 2636 953
rect 2630 948 2631 952
rect 2635 948 2636 952
rect 2630 947 2636 948
rect 2806 952 2812 953
rect 2806 948 2807 952
rect 2811 948 2812 952
rect 2806 947 2812 948
rect 2990 952 2996 953
rect 2990 948 2991 952
rect 2995 948 2996 952
rect 2990 947 2996 948
rect 3182 952 3188 953
rect 3182 948 3183 952
rect 3187 948 3188 952
rect 3182 947 3188 948
rect 2632 931 2634 947
rect 2808 931 2810 947
rect 2992 931 2994 947
rect 3184 931 3186 947
rect 2479 930 2483 931
rect 2479 925 2483 926
rect 2567 930 2571 931
rect 2567 925 2571 926
rect 2631 930 2635 931
rect 2631 925 2635 926
rect 2655 930 2659 931
rect 2655 925 2659 926
rect 2743 930 2747 931
rect 2743 925 2747 926
rect 2807 930 2811 931
rect 2807 925 2811 926
rect 2831 930 2835 931
rect 2831 925 2835 926
rect 2991 930 2995 931
rect 2991 925 2995 926
rect 3183 930 3187 931
rect 3183 925 3187 926
rect 2480 909 2482 925
rect 2568 909 2570 925
rect 2656 909 2658 925
rect 2744 909 2746 925
rect 2832 909 2834 925
rect 2478 908 2484 909
rect 2478 904 2479 908
rect 2483 904 2484 908
rect 2478 903 2484 904
rect 2566 908 2572 909
rect 2566 904 2567 908
rect 2571 904 2572 908
rect 2566 903 2572 904
rect 2654 908 2660 909
rect 2654 904 2655 908
rect 2659 904 2660 908
rect 2654 903 2660 904
rect 2742 908 2748 909
rect 2742 904 2743 908
rect 2747 904 2748 908
rect 2742 903 2748 904
rect 2830 908 2836 909
rect 2830 904 2831 908
rect 2835 904 2836 908
rect 2830 903 2836 904
rect 2286 899 2292 900
rect 2286 895 2287 899
rect 2291 895 2292 899
rect 2286 894 2292 895
rect 2374 899 2380 900
rect 2374 895 2375 899
rect 2379 895 2380 899
rect 2374 894 2380 895
rect 2462 899 2468 900
rect 2462 895 2463 899
rect 2467 895 2468 899
rect 2462 894 2468 895
rect 2470 899 2476 900
rect 2470 895 2471 899
rect 2475 895 2476 899
rect 2470 894 2476 895
rect 2638 899 2644 900
rect 2638 895 2639 899
rect 2643 895 2644 899
rect 2638 894 2644 895
rect 2726 899 2732 900
rect 2726 895 2727 899
rect 2731 895 2732 899
rect 2726 894 2732 895
rect 2814 899 2820 900
rect 2814 895 2815 899
rect 2819 895 2820 899
rect 2814 894 2820 895
rect 2822 899 2828 900
rect 2822 895 2823 899
rect 2827 895 2828 899
rect 2822 894 2828 895
rect 2214 889 2220 890
rect 2214 885 2215 889
rect 2219 885 2220 889
rect 2214 884 2220 885
rect 2206 871 2212 872
rect 2206 867 2207 871
rect 2211 867 2212 871
rect 2206 866 2212 867
rect 2216 859 2218 884
rect 2288 872 2290 894
rect 2302 889 2308 890
rect 2302 885 2303 889
rect 2307 885 2308 889
rect 2302 884 2308 885
rect 2286 871 2292 872
rect 2286 867 2287 871
rect 2291 867 2292 871
rect 2286 866 2292 867
rect 2304 859 2306 884
rect 2376 872 2378 894
rect 2390 889 2396 890
rect 2390 885 2391 889
rect 2395 885 2396 889
rect 2390 884 2396 885
rect 2374 871 2380 872
rect 2374 867 2375 871
rect 2379 867 2380 871
rect 2374 866 2380 867
rect 2392 859 2394 884
rect 2464 864 2466 894
rect 2478 889 2484 890
rect 2478 885 2479 889
rect 2483 885 2484 889
rect 2478 884 2484 885
rect 2566 889 2572 890
rect 2566 885 2567 889
rect 2571 885 2572 889
rect 2566 884 2572 885
rect 2462 863 2468 864
rect 2462 859 2463 863
rect 2467 859 2468 863
rect 2480 859 2482 884
rect 2518 871 2524 872
rect 2518 867 2519 871
rect 2523 867 2524 871
rect 2518 866 2524 867
rect 1335 858 1339 859
rect 1335 853 1339 854
rect 1559 858 1563 859
rect 1559 853 1563 854
rect 1767 858 1771 859
rect 1767 853 1771 854
rect 1807 858 1811 859
rect 1807 853 1811 854
rect 2127 858 2131 859
rect 2127 853 2131 854
rect 2159 858 2163 859
rect 2159 853 2163 854
rect 2215 858 2219 859
rect 2215 853 2219 854
rect 2247 858 2251 859
rect 2247 853 2251 854
rect 2303 858 2307 859
rect 2303 853 2307 854
rect 2335 858 2339 859
rect 2335 853 2339 854
rect 2391 858 2395 859
rect 2391 853 2395 854
rect 2423 858 2427 859
rect 2462 858 2468 859
rect 2479 858 2483 859
rect 2423 853 2427 854
rect 2479 853 2483 854
rect 1322 851 1328 852
rect 1322 847 1323 851
rect 1327 847 1328 851
rect 1322 846 1328 847
rect 1768 837 1770 853
rect 1808 837 1810 853
rect 1766 836 1772 837
rect 1270 835 1276 836
rect 1270 831 1271 835
rect 1275 831 1276 835
rect 1766 832 1767 836
rect 1771 832 1772 836
rect 1766 831 1772 832
rect 1806 836 1812 837
rect 2160 836 2162 853
rect 2222 851 2228 852
rect 2222 847 2223 851
rect 2227 847 2228 851
rect 2222 846 2228 847
rect 2230 851 2236 852
rect 2230 847 2231 851
rect 2235 847 2236 851
rect 2230 846 2236 847
rect 1806 832 1807 836
rect 1811 832 1812 836
rect 1806 831 1812 832
rect 2158 835 2164 836
rect 2158 831 2159 835
rect 2163 831 2164 835
rect 1270 830 1276 831
rect 2158 830 2164 831
rect 822 827 828 828
rect 822 823 823 827
rect 827 823 828 827
rect 822 822 828 823
rect 1114 827 1120 828
rect 1114 823 1115 827
rect 1119 823 1120 827
rect 1230 827 1236 828
rect 1114 822 1120 823
rect 1206 823 1212 824
rect 1206 819 1207 823
rect 1211 819 1212 823
rect 1230 823 1231 827
rect 1235 823 1236 827
rect 1230 822 1236 823
rect 1206 818 1212 819
rect 1766 819 1772 820
rect 878 816 884 817
rect 878 812 879 816
rect 883 812 884 816
rect 878 811 884 812
rect 1006 816 1012 817
rect 1006 812 1007 816
rect 1011 812 1012 816
rect 1006 811 1012 812
rect 1134 816 1140 817
rect 1134 812 1135 816
rect 1139 812 1140 816
rect 1134 811 1140 812
rect 880 791 882 811
rect 1008 791 1010 811
rect 1136 791 1138 811
rect 879 790 883 791
rect 879 785 883 786
rect 887 790 891 791
rect 887 785 891 786
rect 1007 790 1011 791
rect 1007 785 1011 786
rect 1039 790 1043 791
rect 1039 785 1043 786
rect 1135 790 1139 791
rect 1135 785 1139 786
rect 1191 790 1195 791
rect 1191 785 1195 786
rect 888 769 890 785
rect 1040 769 1042 785
rect 1192 769 1194 785
rect 886 768 892 769
rect 886 764 887 768
rect 891 764 892 768
rect 886 763 892 764
rect 1038 768 1044 769
rect 1038 764 1039 768
rect 1043 764 1044 768
rect 1038 763 1044 764
rect 1190 768 1196 769
rect 1190 764 1191 768
rect 1195 764 1196 768
rect 1190 763 1196 764
rect 206 759 212 760
rect 206 755 207 759
rect 211 755 212 759
rect 206 754 212 755
rect 294 759 300 760
rect 294 755 295 759
rect 299 755 300 759
rect 294 754 300 755
rect 414 759 420 760
rect 414 755 415 759
rect 419 755 420 759
rect 414 754 420 755
rect 542 759 548 760
rect 542 755 543 759
rect 547 755 548 759
rect 542 754 548 755
rect 550 759 556 760
rect 550 755 551 759
rect 555 755 556 759
rect 550 754 556 755
rect 806 759 812 760
rect 806 755 807 759
rect 811 755 812 759
rect 806 754 812 755
rect 822 759 828 760
rect 822 755 823 759
rect 827 755 828 759
rect 822 754 828 755
rect 966 759 972 760
rect 966 755 967 759
rect 971 755 972 759
rect 966 754 972 755
rect 208 732 210 754
rect 222 749 228 750
rect 222 745 223 749
rect 227 745 228 749
rect 222 744 228 745
rect 198 731 204 732
rect 198 727 199 731
rect 203 727 204 731
rect 198 726 204 727
rect 206 731 212 732
rect 206 727 207 731
rect 211 727 212 731
rect 206 726 212 727
rect 224 723 226 744
rect 296 732 298 754
rect 342 749 348 750
rect 342 745 343 749
rect 347 745 348 749
rect 342 744 348 745
rect 294 731 300 732
rect 294 727 295 731
rect 299 727 300 731
rect 294 726 300 727
rect 344 723 346 744
rect 416 732 418 754
rect 470 749 476 750
rect 470 745 471 749
rect 475 745 476 749
rect 470 744 476 745
rect 414 731 420 732
rect 414 727 415 731
rect 419 727 420 731
rect 414 726 420 727
rect 472 723 474 744
rect 544 732 546 754
rect 542 731 548 732
rect 542 727 543 731
rect 547 727 548 731
rect 542 726 548 727
rect 552 724 554 754
rect 606 749 612 750
rect 606 745 607 749
rect 611 745 612 749
rect 606 744 612 745
rect 742 749 748 750
rect 742 745 743 749
rect 747 745 748 749
rect 742 744 748 745
rect 550 723 556 724
rect 608 723 610 744
rect 744 723 746 744
rect 824 732 826 754
rect 886 749 892 750
rect 886 745 887 749
rect 891 745 892 749
rect 886 744 892 745
rect 822 731 828 732
rect 822 727 823 731
rect 827 727 828 731
rect 822 726 828 727
rect 888 723 890 744
rect 968 732 970 754
rect 1038 749 1044 750
rect 1038 745 1039 749
rect 1043 745 1044 749
rect 1038 744 1044 745
rect 1190 749 1196 750
rect 1190 745 1191 749
rect 1195 745 1196 749
rect 1190 744 1196 745
rect 966 731 972 732
rect 966 727 967 731
rect 971 727 972 731
rect 966 726 972 727
rect 1040 723 1042 744
rect 1102 731 1108 732
rect 1102 727 1103 731
rect 1107 727 1108 731
rect 1102 726 1108 727
rect 111 722 115 723
rect 111 717 115 718
rect 135 722 139 723
rect 135 717 139 718
rect 167 722 171 723
rect 167 717 171 718
rect 223 722 227 723
rect 223 717 227 718
rect 295 722 299 723
rect 295 717 299 718
rect 343 722 347 723
rect 343 717 347 718
rect 431 722 435 723
rect 431 717 435 718
rect 471 722 475 723
rect 550 719 551 723
rect 555 719 556 723
rect 550 718 556 719
rect 575 722 579 723
rect 471 717 475 718
rect 575 717 579 718
rect 607 722 611 723
rect 607 717 611 718
rect 727 722 731 723
rect 727 717 731 718
rect 743 722 747 723
rect 743 717 747 718
rect 879 722 883 723
rect 879 717 883 718
rect 887 722 891 723
rect 887 717 891 718
rect 1031 722 1035 723
rect 1031 717 1035 718
rect 1039 722 1043 723
rect 1039 717 1043 718
rect 112 701 114 717
rect 110 700 116 701
rect 168 700 170 717
rect 274 711 280 712
rect 274 707 275 711
rect 279 707 280 711
rect 274 706 280 707
rect 110 696 111 700
rect 115 696 116 700
rect 110 695 116 696
rect 166 699 172 700
rect 166 695 167 699
rect 171 695 172 699
rect 166 694 172 695
rect 276 692 278 706
rect 296 700 298 717
rect 366 715 372 716
rect 366 711 367 715
rect 371 711 372 715
rect 366 710 372 711
rect 294 699 300 700
rect 294 695 295 699
rect 299 695 300 699
rect 294 694 300 695
rect 368 692 370 710
rect 432 700 434 717
rect 502 715 508 716
rect 502 711 503 715
rect 507 711 508 715
rect 502 710 508 711
rect 430 699 436 700
rect 430 695 431 699
rect 435 695 436 699
rect 430 694 436 695
rect 504 692 506 710
rect 576 700 578 717
rect 646 715 652 716
rect 646 711 647 715
rect 651 711 652 715
rect 646 710 652 711
rect 574 699 580 700
rect 574 695 575 699
rect 579 695 580 699
rect 574 694 580 695
rect 648 692 650 710
rect 728 700 730 717
rect 880 700 882 717
rect 942 715 948 716
rect 942 711 943 715
rect 947 711 948 715
rect 942 710 948 711
rect 950 715 956 716
rect 950 711 951 715
rect 955 711 956 715
rect 950 710 956 711
rect 726 699 732 700
rect 726 695 727 699
rect 731 695 732 699
rect 726 694 732 695
rect 878 699 884 700
rect 878 695 879 699
rect 883 695 884 699
rect 878 694 884 695
rect 274 691 280 692
rect 274 687 275 691
rect 279 687 280 691
rect 274 686 280 687
rect 366 691 372 692
rect 366 687 367 691
rect 371 687 372 691
rect 366 686 372 687
rect 502 691 508 692
rect 502 687 503 691
rect 507 687 508 691
rect 502 686 508 687
rect 646 691 652 692
rect 646 687 647 691
rect 651 687 652 691
rect 646 686 652 687
rect 654 691 660 692
rect 654 687 655 691
rect 659 687 660 691
rect 654 686 660 687
rect 110 683 116 684
rect 110 679 111 683
rect 115 679 116 683
rect 110 678 116 679
rect 166 680 172 681
rect 112 655 114 678
rect 166 676 167 680
rect 171 676 172 680
rect 166 675 172 676
rect 294 680 300 681
rect 294 676 295 680
rect 299 676 300 680
rect 294 675 300 676
rect 430 680 436 681
rect 430 676 431 680
rect 435 676 436 680
rect 430 675 436 676
rect 574 680 580 681
rect 574 676 575 680
rect 579 676 580 680
rect 574 675 580 676
rect 168 655 170 675
rect 296 655 298 675
rect 432 655 434 675
rect 576 655 578 675
rect 111 654 115 655
rect 111 649 115 650
rect 167 654 171 655
rect 167 649 171 650
rect 295 654 299 655
rect 295 649 299 650
rect 431 654 435 655
rect 431 649 435 650
rect 455 654 459 655
rect 455 649 459 650
rect 559 654 563 655
rect 559 649 563 650
rect 575 654 579 655
rect 575 649 579 650
rect 112 630 114 649
rect 456 633 458 649
rect 560 633 562 649
rect 454 632 460 633
rect 110 629 116 630
rect 110 625 111 629
rect 115 625 116 629
rect 454 628 455 632
rect 459 628 460 632
rect 454 627 460 628
rect 558 632 564 633
rect 558 628 559 632
rect 563 628 564 632
rect 558 627 564 628
rect 110 624 116 625
rect 526 623 532 624
rect 526 619 527 623
rect 531 619 532 623
rect 526 618 532 619
rect 630 623 636 624
rect 630 619 631 623
rect 635 619 636 623
rect 630 618 636 619
rect 454 613 460 614
rect 110 612 116 613
rect 110 608 111 612
rect 115 608 116 612
rect 454 609 455 613
rect 459 609 460 613
rect 454 608 460 609
rect 110 607 116 608
rect 112 583 114 607
rect 456 583 458 608
rect 528 596 530 618
rect 558 613 564 614
rect 558 609 559 613
rect 563 609 564 613
rect 558 608 564 609
rect 526 595 532 596
rect 526 591 527 595
rect 531 591 532 595
rect 526 590 532 591
rect 560 583 562 608
rect 632 596 634 618
rect 630 595 636 596
rect 630 591 631 595
rect 635 591 636 595
rect 630 590 636 591
rect 656 588 658 686
rect 726 680 732 681
rect 726 676 727 680
rect 731 676 732 680
rect 726 675 732 676
rect 878 680 884 681
rect 878 676 879 680
rect 883 676 884 680
rect 878 675 884 676
rect 728 655 730 675
rect 880 655 882 675
rect 679 654 683 655
rect 679 649 683 650
rect 727 654 731 655
rect 727 649 731 650
rect 799 654 803 655
rect 799 649 803 650
rect 879 654 883 655
rect 879 649 883 650
rect 927 654 931 655
rect 927 649 931 650
rect 680 633 682 649
rect 800 633 802 649
rect 928 633 930 649
rect 944 640 946 710
rect 952 692 954 710
rect 1032 700 1034 717
rect 1030 699 1036 700
rect 1030 695 1031 699
rect 1035 695 1036 699
rect 1030 694 1036 695
rect 1104 692 1106 726
rect 1192 723 1194 744
rect 1208 732 1210 818
rect 1270 816 1276 817
rect 1270 812 1271 816
rect 1275 812 1276 816
rect 1766 815 1767 819
rect 1771 815 1772 819
rect 1766 814 1772 815
rect 1806 819 1812 820
rect 1806 815 1807 819
rect 1811 815 1812 819
rect 1806 814 1812 815
rect 2158 816 2164 817
rect 1270 811 1276 812
rect 1272 791 1274 811
rect 1768 791 1770 814
rect 1808 791 1810 814
rect 2158 812 2159 816
rect 2163 812 2164 816
rect 2158 811 2164 812
rect 2160 791 2162 811
rect 1271 790 1275 791
rect 1271 785 1275 786
rect 1351 790 1355 791
rect 1351 785 1355 786
rect 1767 790 1771 791
rect 1767 785 1771 786
rect 1807 790 1811 791
rect 1807 785 1811 786
rect 2063 790 2067 791
rect 2063 785 2067 786
rect 2159 790 2163 791
rect 2159 785 2163 786
rect 2175 790 2179 791
rect 2175 785 2179 786
rect 1352 769 1354 785
rect 1350 768 1356 769
rect 1350 764 1351 768
rect 1355 764 1356 768
rect 1768 766 1770 785
rect 1808 766 1810 785
rect 2064 769 2066 785
rect 2176 769 2178 785
rect 2224 776 2226 846
rect 2232 828 2234 846
rect 2248 836 2250 853
rect 2318 851 2324 852
rect 2318 847 2319 851
rect 2323 847 2324 851
rect 2318 846 2324 847
rect 2246 835 2252 836
rect 2246 831 2247 835
rect 2251 831 2252 835
rect 2246 830 2252 831
rect 2320 828 2322 846
rect 2336 836 2338 853
rect 2406 851 2412 852
rect 2406 847 2407 851
rect 2411 847 2412 851
rect 2406 846 2412 847
rect 2334 835 2340 836
rect 2334 831 2335 835
rect 2339 831 2340 835
rect 2334 830 2340 831
rect 2408 828 2410 846
rect 2424 836 2426 853
rect 2494 851 2500 852
rect 2494 847 2495 851
rect 2499 847 2500 851
rect 2494 846 2500 847
rect 2422 835 2428 836
rect 2422 831 2423 835
rect 2427 831 2428 835
rect 2422 830 2428 831
rect 2496 828 2498 846
rect 2520 828 2522 866
rect 2568 859 2570 884
rect 2640 872 2642 894
rect 2654 889 2660 890
rect 2654 885 2655 889
rect 2659 885 2660 889
rect 2654 884 2660 885
rect 2638 871 2644 872
rect 2638 867 2639 871
rect 2643 867 2644 871
rect 2638 866 2644 867
rect 2656 859 2658 884
rect 2728 872 2730 894
rect 2742 889 2748 890
rect 2742 885 2743 889
rect 2747 885 2748 889
rect 2742 884 2748 885
rect 2726 871 2732 872
rect 2726 867 2727 871
rect 2731 867 2732 871
rect 2726 866 2732 867
rect 2744 859 2746 884
rect 2816 872 2818 894
rect 2814 871 2820 872
rect 2814 867 2815 871
rect 2819 867 2820 871
rect 2814 866 2820 867
rect 2824 860 2826 894
rect 2830 889 2836 890
rect 2830 885 2831 889
rect 2835 885 2836 889
rect 2830 884 2836 885
rect 2822 859 2828 860
rect 2832 859 2834 884
rect 2527 858 2531 859
rect 2527 853 2531 854
rect 2567 858 2571 859
rect 2567 853 2571 854
rect 2639 858 2643 859
rect 2639 853 2643 854
rect 2655 858 2659 859
rect 2655 853 2659 854
rect 2743 858 2747 859
rect 2743 853 2747 854
rect 2767 858 2771 859
rect 2822 855 2823 859
rect 2827 855 2828 859
rect 2822 854 2828 855
rect 2831 858 2835 859
rect 2767 853 2771 854
rect 2831 853 2835 854
rect 2911 858 2915 859
rect 2911 853 2915 854
rect 3063 858 3067 859
rect 3063 853 3067 854
rect 3223 858 3227 859
rect 3223 853 3227 854
rect 2528 836 2530 853
rect 2640 836 2642 853
rect 2710 851 2716 852
rect 2710 847 2711 851
rect 2715 847 2716 851
rect 2710 846 2716 847
rect 2526 835 2532 836
rect 2526 831 2527 835
rect 2531 831 2532 835
rect 2526 830 2532 831
rect 2638 835 2644 836
rect 2638 831 2639 835
rect 2643 831 2644 835
rect 2638 830 2644 831
rect 2712 828 2714 846
rect 2768 836 2770 853
rect 2838 851 2844 852
rect 2838 847 2839 851
rect 2843 847 2844 851
rect 2838 846 2844 847
rect 2766 835 2772 836
rect 2766 831 2767 835
rect 2771 831 2772 835
rect 2766 830 2772 831
rect 2840 828 2842 846
rect 2912 836 2914 853
rect 2982 851 2988 852
rect 2982 847 2983 851
rect 2987 847 2988 851
rect 2982 846 2988 847
rect 2910 835 2916 836
rect 2910 831 2911 835
rect 2915 831 2916 835
rect 2910 830 2916 831
rect 2984 828 2986 846
rect 3064 836 3066 853
rect 3190 851 3196 852
rect 3190 847 3191 851
rect 3195 847 3196 851
rect 3190 846 3196 847
rect 3062 835 3068 836
rect 3062 831 3063 835
rect 3067 831 3068 835
rect 3062 830 3068 831
rect 2230 827 2236 828
rect 2230 823 2231 827
rect 2235 823 2236 827
rect 2230 822 2236 823
rect 2318 827 2324 828
rect 2318 823 2319 827
rect 2323 823 2324 827
rect 2318 822 2324 823
rect 2406 827 2412 828
rect 2406 823 2407 827
rect 2411 823 2412 827
rect 2406 822 2412 823
rect 2494 827 2500 828
rect 2494 823 2495 827
rect 2499 823 2500 827
rect 2494 822 2500 823
rect 2518 827 2524 828
rect 2518 823 2519 827
rect 2523 823 2524 827
rect 2518 822 2524 823
rect 2710 827 2716 828
rect 2710 823 2711 827
rect 2715 823 2716 827
rect 2710 822 2716 823
rect 2838 827 2844 828
rect 2838 823 2839 827
rect 2843 823 2844 827
rect 2838 822 2844 823
rect 2982 827 2988 828
rect 2982 823 2983 827
rect 2987 823 2988 827
rect 2982 822 2988 823
rect 2990 827 2996 828
rect 2990 823 2991 827
rect 2995 823 2996 827
rect 2990 822 2996 823
rect 2246 816 2252 817
rect 2246 812 2247 816
rect 2251 812 2252 816
rect 2246 811 2252 812
rect 2334 816 2340 817
rect 2334 812 2335 816
rect 2339 812 2340 816
rect 2334 811 2340 812
rect 2422 816 2428 817
rect 2422 812 2423 816
rect 2427 812 2428 816
rect 2422 811 2428 812
rect 2526 816 2532 817
rect 2526 812 2527 816
rect 2531 812 2532 816
rect 2526 811 2532 812
rect 2638 816 2644 817
rect 2638 812 2639 816
rect 2643 812 2644 816
rect 2638 811 2644 812
rect 2766 816 2772 817
rect 2766 812 2767 816
rect 2771 812 2772 816
rect 2766 811 2772 812
rect 2910 816 2916 817
rect 2910 812 2911 816
rect 2915 812 2916 816
rect 2910 811 2916 812
rect 2248 791 2250 811
rect 2336 791 2338 811
rect 2424 791 2426 811
rect 2528 791 2530 811
rect 2640 791 2642 811
rect 2768 791 2770 811
rect 2912 791 2914 811
rect 2247 790 2251 791
rect 2247 785 2251 786
rect 2295 790 2299 791
rect 2295 785 2299 786
rect 2335 790 2339 791
rect 2335 785 2339 786
rect 2423 790 2427 791
rect 2423 785 2427 786
rect 2527 790 2531 791
rect 2527 785 2531 786
rect 2559 790 2563 791
rect 2559 785 2563 786
rect 2639 790 2643 791
rect 2639 785 2643 786
rect 2711 790 2715 791
rect 2711 785 2715 786
rect 2767 790 2771 791
rect 2767 785 2771 786
rect 2871 790 2875 791
rect 2871 785 2875 786
rect 2911 790 2915 791
rect 2911 785 2915 786
rect 2222 775 2228 776
rect 2222 771 2223 775
rect 2227 771 2228 775
rect 2222 770 2228 771
rect 2296 769 2298 785
rect 2424 769 2426 785
rect 2560 769 2562 785
rect 2712 769 2714 785
rect 2762 779 2768 780
rect 2762 775 2763 779
rect 2767 775 2768 779
rect 2762 774 2768 775
rect 2062 768 2068 769
rect 1350 763 1356 764
rect 1766 765 1772 766
rect 1766 761 1767 765
rect 1771 761 1772 765
rect 1766 760 1772 761
rect 1806 765 1812 766
rect 1806 761 1807 765
rect 1811 761 1812 765
rect 2062 764 2063 768
rect 2067 764 2068 768
rect 2062 763 2068 764
rect 2174 768 2180 769
rect 2174 764 2175 768
rect 2179 764 2180 768
rect 2174 763 2180 764
rect 2294 768 2300 769
rect 2294 764 2295 768
rect 2299 764 2300 768
rect 2294 763 2300 764
rect 2422 768 2428 769
rect 2422 764 2423 768
rect 2427 764 2428 768
rect 2422 763 2428 764
rect 2558 768 2564 769
rect 2558 764 2559 768
rect 2563 764 2564 768
rect 2558 763 2564 764
rect 2710 768 2716 769
rect 2710 764 2711 768
rect 2715 764 2716 768
rect 2710 763 2716 764
rect 1806 760 1812 761
rect 1262 759 1268 760
rect 1262 755 1263 759
rect 1267 755 1268 759
rect 1262 754 1268 755
rect 1470 759 1476 760
rect 1470 755 1471 759
rect 1475 755 1476 759
rect 1470 754 1476 755
rect 2134 759 2140 760
rect 2134 755 2135 759
rect 2139 755 2140 759
rect 2134 754 2140 755
rect 2246 759 2252 760
rect 2246 755 2247 759
rect 2251 755 2252 759
rect 2246 754 2252 755
rect 2366 759 2372 760
rect 2366 755 2367 759
rect 2371 755 2372 759
rect 2366 754 2372 755
rect 2494 759 2500 760
rect 2494 755 2495 759
rect 2499 755 2500 759
rect 2494 754 2500 755
rect 1264 732 1266 754
rect 1350 749 1356 750
rect 1350 745 1351 749
rect 1355 745 1356 749
rect 1350 744 1356 745
rect 1206 731 1212 732
rect 1206 727 1207 731
rect 1211 727 1212 731
rect 1206 726 1212 727
rect 1262 731 1268 732
rect 1262 727 1263 731
rect 1267 727 1268 731
rect 1262 726 1268 727
rect 1352 723 1354 744
rect 1183 722 1187 723
rect 1183 717 1187 718
rect 1191 722 1195 723
rect 1191 717 1195 718
rect 1343 722 1347 723
rect 1343 717 1347 718
rect 1351 722 1355 723
rect 1351 717 1355 718
rect 1184 700 1186 717
rect 1262 715 1268 716
rect 1262 711 1263 715
rect 1267 711 1268 715
rect 1262 710 1268 711
rect 1182 699 1188 700
rect 1182 695 1183 699
rect 1187 695 1188 699
rect 1182 694 1188 695
rect 1264 692 1266 710
rect 1344 700 1346 717
rect 1472 716 1474 754
rect 2062 749 2068 750
rect 1766 748 1772 749
rect 1766 744 1767 748
rect 1771 744 1772 748
rect 1766 743 1772 744
rect 1806 748 1812 749
rect 1806 744 1807 748
rect 1811 744 1812 748
rect 2062 745 2063 749
rect 2067 745 2068 749
rect 2062 744 2068 745
rect 1806 743 1812 744
rect 1768 723 1770 743
rect 1808 727 1810 743
rect 2064 727 2066 744
rect 2136 732 2138 754
rect 2174 749 2180 750
rect 2174 745 2175 749
rect 2179 745 2180 749
rect 2174 744 2180 745
rect 2114 731 2120 732
rect 2114 727 2115 731
rect 2119 727 2120 731
rect 1807 726 1811 727
rect 1503 722 1507 723
rect 1503 717 1507 718
rect 1767 722 1771 723
rect 1807 721 1811 722
rect 1927 726 1931 727
rect 1927 721 1931 722
rect 2063 726 2067 727
rect 2063 721 2067 722
rect 2071 726 2075 727
rect 2114 726 2120 727
rect 2134 731 2140 732
rect 2134 727 2135 731
rect 2139 727 2140 731
rect 2176 727 2178 744
rect 2248 732 2250 754
rect 2294 749 2300 750
rect 2294 745 2295 749
rect 2299 745 2300 749
rect 2294 744 2300 745
rect 2246 731 2252 732
rect 2246 727 2247 731
rect 2251 727 2252 731
rect 2296 727 2298 744
rect 2368 732 2370 754
rect 2422 749 2428 750
rect 2422 745 2423 749
rect 2427 745 2428 749
rect 2422 744 2428 745
rect 2366 731 2372 732
rect 2366 727 2367 731
rect 2371 727 2372 731
rect 2424 727 2426 744
rect 2496 732 2498 754
rect 2558 749 2564 750
rect 2558 745 2559 749
rect 2563 745 2564 749
rect 2558 744 2564 745
rect 2710 749 2716 750
rect 2710 745 2711 749
rect 2715 745 2716 749
rect 2710 744 2716 745
rect 2494 731 2500 732
rect 2494 727 2495 731
rect 2499 727 2500 731
rect 2560 727 2562 744
rect 2712 727 2714 744
rect 2764 732 2766 774
rect 2872 769 2874 785
rect 2992 780 2994 822
rect 3062 816 3068 817
rect 3062 812 3063 816
rect 3067 812 3068 816
rect 3062 811 3068 812
rect 3064 791 3066 811
rect 3039 790 3043 791
rect 3039 785 3043 786
rect 3063 790 3067 791
rect 3063 785 3067 786
rect 2990 779 2996 780
rect 2990 775 2991 779
rect 2995 775 2996 779
rect 2990 774 2996 775
rect 3040 769 3042 785
rect 2870 768 2876 769
rect 2870 764 2871 768
rect 2875 764 2876 768
rect 2870 763 2876 764
rect 3038 768 3044 769
rect 3038 764 3039 768
rect 3043 764 3044 768
rect 3038 763 3044 764
rect 2782 759 2788 760
rect 2782 755 2783 759
rect 2787 755 2788 759
rect 2782 754 2788 755
rect 2942 759 2948 760
rect 2942 755 2943 759
rect 2947 755 2948 759
rect 2942 754 2948 755
rect 3110 759 3116 760
rect 3110 755 3111 759
rect 3115 755 3116 759
rect 3110 754 3116 755
rect 2784 732 2786 754
rect 2870 749 2876 750
rect 2870 745 2871 749
rect 2875 745 2876 749
rect 2870 744 2876 745
rect 2762 731 2768 732
rect 2762 727 2763 731
rect 2767 727 2768 731
rect 2134 726 2140 727
rect 2175 726 2179 727
rect 2071 721 2075 722
rect 1767 717 1771 718
rect 1422 715 1428 716
rect 1422 711 1423 715
rect 1427 711 1428 715
rect 1422 710 1428 711
rect 1470 715 1476 716
rect 1470 711 1471 715
rect 1475 711 1476 715
rect 1470 710 1476 711
rect 1342 699 1348 700
rect 1342 695 1343 699
rect 1347 695 1348 699
rect 1342 694 1348 695
rect 1424 692 1426 710
rect 1504 700 1506 717
rect 1768 701 1770 717
rect 1808 705 1810 721
rect 1806 704 1812 705
rect 1928 704 1930 721
rect 1986 719 1992 720
rect 1986 715 1987 719
rect 1991 715 1992 719
rect 1986 714 1992 715
rect 1998 719 2004 720
rect 1998 715 1999 719
rect 2003 715 2004 719
rect 1998 714 2004 715
rect 1766 700 1772 701
rect 1502 699 1508 700
rect 1502 695 1503 699
rect 1507 695 1508 699
rect 1766 696 1767 700
rect 1771 696 1772 700
rect 1806 700 1807 704
rect 1811 700 1812 704
rect 1806 699 1812 700
rect 1926 703 1932 704
rect 1926 699 1927 703
rect 1931 699 1932 703
rect 1926 698 1932 699
rect 1766 695 1772 696
rect 1502 694 1508 695
rect 950 691 956 692
rect 950 687 951 691
rect 955 687 956 691
rect 950 686 956 687
rect 1102 691 1108 692
rect 1102 687 1103 691
rect 1107 687 1108 691
rect 1262 691 1268 692
rect 1102 686 1108 687
rect 1254 687 1260 688
rect 1254 683 1255 687
rect 1259 683 1260 687
rect 1262 687 1263 691
rect 1267 687 1268 691
rect 1262 686 1268 687
rect 1422 691 1428 692
rect 1422 687 1423 691
rect 1427 687 1428 691
rect 1422 686 1428 687
rect 1806 687 1812 688
rect 1254 682 1260 683
rect 1766 683 1772 684
rect 1030 680 1036 681
rect 1030 676 1031 680
rect 1035 676 1036 680
rect 1030 675 1036 676
rect 1182 680 1188 681
rect 1182 676 1183 680
rect 1187 676 1188 680
rect 1182 675 1188 676
rect 1032 655 1034 675
rect 1184 655 1186 675
rect 1031 654 1035 655
rect 1031 649 1035 650
rect 1055 654 1059 655
rect 1055 649 1059 650
rect 1183 654 1187 655
rect 1183 649 1187 650
rect 942 639 948 640
rect 942 635 943 639
rect 947 635 948 639
rect 942 634 948 635
rect 1056 633 1058 649
rect 1184 633 1186 649
rect 678 632 684 633
rect 678 628 679 632
rect 683 628 684 632
rect 678 627 684 628
rect 798 632 804 633
rect 798 628 799 632
rect 803 628 804 632
rect 798 627 804 628
rect 926 632 932 633
rect 926 628 927 632
rect 931 628 932 632
rect 926 627 932 628
rect 1054 632 1060 633
rect 1054 628 1055 632
rect 1059 628 1060 632
rect 1054 627 1060 628
rect 1182 632 1188 633
rect 1182 628 1183 632
rect 1187 628 1188 632
rect 1182 627 1188 628
rect 750 623 756 624
rect 750 619 751 623
rect 755 619 756 623
rect 750 618 756 619
rect 870 623 876 624
rect 870 619 871 623
rect 875 619 876 623
rect 870 618 876 619
rect 990 623 996 624
rect 990 619 991 623
rect 995 619 996 623
rect 990 618 996 619
rect 1134 623 1140 624
rect 1134 619 1135 623
rect 1139 619 1140 623
rect 1134 618 1140 619
rect 678 613 684 614
rect 678 609 679 613
rect 683 609 684 613
rect 678 608 684 609
rect 654 587 660 588
rect 654 583 655 587
rect 659 583 660 587
rect 680 583 682 608
rect 752 596 754 618
rect 798 613 804 614
rect 798 609 799 613
rect 803 609 804 613
rect 798 608 804 609
rect 750 595 756 596
rect 750 591 751 595
rect 755 591 756 595
rect 750 590 756 591
rect 800 583 802 608
rect 872 596 874 618
rect 926 613 932 614
rect 926 609 927 613
rect 931 609 932 613
rect 926 608 932 609
rect 870 595 876 596
rect 870 591 871 595
rect 875 591 876 595
rect 870 590 876 591
rect 928 583 930 608
rect 111 582 115 583
rect 111 577 115 578
rect 455 582 459 583
rect 455 577 459 578
rect 559 582 563 583
rect 559 577 563 578
rect 599 582 603 583
rect 654 582 660 583
rect 679 582 683 583
rect 599 577 603 578
rect 679 577 683 578
rect 703 582 707 583
rect 703 577 707 578
rect 799 582 803 583
rect 799 577 803 578
rect 815 582 819 583
rect 815 577 819 578
rect 927 582 931 583
rect 927 577 931 578
rect 112 561 114 577
rect 110 560 116 561
rect 600 560 602 577
rect 670 575 676 576
rect 670 571 671 575
rect 675 571 676 575
rect 670 570 676 571
rect 110 556 111 560
rect 115 556 116 560
rect 110 555 116 556
rect 598 559 604 560
rect 598 555 599 559
rect 603 555 604 559
rect 598 554 604 555
rect 672 552 674 570
rect 704 560 706 577
rect 774 575 780 576
rect 774 571 775 575
rect 779 571 780 575
rect 774 570 780 571
rect 702 559 708 560
rect 702 555 703 559
rect 707 555 708 559
rect 702 554 708 555
rect 776 552 778 570
rect 816 560 818 577
rect 928 560 930 577
rect 992 576 994 618
rect 1054 613 1060 614
rect 1054 609 1055 613
rect 1059 609 1060 613
rect 1054 608 1060 609
rect 1006 583 1012 584
rect 1056 583 1058 608
rect 1136 596 1138 618
rect 1182 613 1188 614
rect 1182 609 1183 613
rect 1187 609 1188 613
rect 1182 608 1188 609
rect 1134 595 1140 596
rect 1134 591 1135 595
rect 1139 591 1140 595
rect 1134 590 1140 591
rect 1184 583 1186 608
rect 1256 596 1258 682
rect 1342 680 1348 681
rect 1342 676 1343 680
rect 1347 676 1348 680
rect 1342 675 1348 676
rect 1502 680 1508 681
rect 1502 676 1503 680
rect 1507 676 1508 680
rect 1766 679 1767 683
rect 1771 679 1772 683
rect 1806 683 1807 687
rect 1811 683 1812 687
rect 1806 682 1812 683
rect 1926 684 1932 685
rect 1766 678 1772 679
rect 1502 675 1508 676
rect 1344 655 1346 675
rect 1504 655 1506 675
rect 1768 655 1770 678
rect 1808 655 1810 682
rect 1926 680 1927 684
rect 1931 680 1932 684
rect 1926 679 1932 680
rect 1928 655 1930 679
rect 1988 668 1990 714
rect 2000 696 2002 714
rect 2072 704 2074 721
rect 2070 703 2076 704
rect 2070 699 2071 703
rect 2075 699 2076 703
rect 2070 698 2076 699
rect 1998 695 2004 696
rect 1998 691 1999 695
rect 2003 691 2004 695
rect 1998 690 2004 691
rect 2070 684 2076 685
rect 2070 680 2071 684
rect 2075 680 2076 684
rect 2070 679 2076 680
rect 1986 667 1992 668
rect 1986 663 1987 667
rect 1991 663 1992 667
rect 1986 662 1992 663
rect 2072 655 2074 679
rect 2116 676 2118 726
rect 2175 721 2179 722
rect 2231 726 2235 727
rect 2246 726 2252 727
rect 2295 726 2299 727
rect 2366 726 2372 727
rect 2391 726 2395 727
rect 2231 721 2235 722
rect 2295 721 2299 722
rect 2391 721 2395 722
rect 2423 726 2427 727
rect 2494 726 2500 727
rect 2551 726 2555 727
rect 2423 721 2427 722
rect 2551 721 2555 722
rect 2559 726 2563 727
rect 2559 721 2563 722
rect 2703 726 2707 727
rect 2703 721 2707 722
rect 2711 726 2715 727
rect 2762 726 2768 727
rect 2782 731 2788 732
rect 2782 727 2783 731
rect 2787 727 2788 731
rect 2872 727 2874 744
rect 2944 732 2946 754
rect 3038 749 3044 750
rect 3038 745 3039 749
rect 3043 745 3044 749
rect 3038 744 3044 745
rect 2942 731 2948 732
rect 2942 727 2943 731
rect 2947 727 2948 731
rect 3040 727 3042 744
rect 3112 732 3114 754
rect 3110 731 3116 732
rect 3110 727 3111 731
rect 3115 727 3116 731
rect 2782 726 2788 727
rect 2847 726 2851 727
rect 2711 721 2715 722
rect 2847 721 2851 722
rect 2871 726 2875 727
rect 2942 726 2948 727
rect 2983 726 2987 727
rect 2871 721 2875 722
rect 2983 721 2987 722
rect 3039 726 3043 727
rect 3110 726 3116 727
rect 3119 726 3123 727
rect 3039 721 3043 722
rect 3119 721 3123 722
rect 2142 719 2148 720
rect 2142 715 2143 719
rect 2147 715 2148 719
rect 2142 714 2148 715
rect 2144 696 2146 714
rect 2232 704 2234 721
rect 2302 719 2308 720
rect 2302 715 2303 719
rect 2307 715 2308 719
rect 2302 714 2308 715
rect 2230 703 2236 704
rect 2230 699 2231 703
rect 2235 699 2236 703
rect 2230 698 2236 699
rect 2304 696 2306 714
rect 2392 704 2394 721
rect 2462 719 2468 720
rect 2462 715 2463 719
rect 2467 715 2468 719
rect 2462 714 2468 715
rect 2390 703 2396 704
rect 2390 699 2391 703
rect 2395 699 2396 703
rect 2390 698 2396 699
rect 2464 696 2466 714
rect 2552 704 2554 721
rect 2704 704 2706 721
rect 2794 719 2800 720
rect 2794 715 2795 719
rect 2799 715 2800 719
rect 2794 714 2800 715
rect 2550 703 2556 704
rect 2550 699 2551 703
rect 2555 699 2556 703
rect 2550 698 2556 699
rect 2702 703 2708 704
rect 2702 699 2703 703
rect 2707 699 2708 703
rect 2702 698 2708 699
rect 2796 696 2798 714
rect 2848 704 2850 721
rect 2984 704 2986 721
rect 3120 704 3122 721
rect 2846 703 2852 704
rect 2846 699 2847 703
rect 2851 699 2852 703
rect 2846 698 2852 699
rect 2982 703 2988 704
rect 2982 699 2983 703
rect 2987 699 2988 703
rect 2982 698 2988 699
rect 3118 703 3124 704
rect 3118 699 3119 703
rect 3123 699 3124 703
rect 3118 698 3124 699
rect 3192 696 3194 846
rect 3224 836 3226 853
rect 3222 835 3228 836
rect 3222 831 3223 835
rect 3227 831 3228 835
rect 3222 830 3228 831
rect 3296 828 3298 982
rect 3368 972 3370 989
rect 3432 988 3434 1026
rect 3440 1004 3442 1090
rect 3462 1087 3463 1091
rect 3467 1087 3468 1091
rect 3462 1086 3468 1087
rect 3464 1063 3466 1086
rect 3463 1062 3467 1063
rect 3463 1057 3467 1058
rect 3464 1038 3466 1057
rect 3462 1037 3468 1038
rect 3462 1033 3463 1037
rect 3467 1033 3468 1037
rect 3462 1032 3468 1033
rect 3462 1020 3468 1021
rect 3462 1016 3463 1020
rect 3467 1016 3468 1020
rect 3462 1015 3468 1016
rect 3438 1003 3444 1004
rect 3438 999 3439 1003
rect 3443 999 3444 1003
rect 3438 998 3444 999
rect 3464 995 3466 1015
rect 3463 994 3467 995
rect 3463 989 3467 990
rect 3430 987 3436 988
rect 3430 983 3431 987
rect 3435 983 3436 987
rect 3430 982 3436 983
rect 3464 973 3466 989
rect 3462 972 3468 973
rect 3366 971 3372 972
rect 3366 967 3367 971
rect 3371 967 3372 971
rect 3462 968 3463 972
rect 3467 968 3468 972
rect 3462 967 3468 968
rect 3366 966 3372 967
rect 3438 959 3444 960
rect 3438 955 3439 959
rect 3443 955 3444 959
rect 3438 954 3444 955
rect 3462 955 3468 956
rect 3366 952 3372 953
rect 3366 948 3367 952
rect 3371 948 3372 952
rect 3366 947 3372 948
rect 3368 931 3370 947
rect 3367 930 3371 931
rect 3367 925 3371 926
rect 3367 858 3371 859
rect 3367 853 3371 854
rect 3368 836 3370 853
rect 3440 852 3442 954
rect 3462 951 3463 955
rect 3467 951 3468 955
rect 3462 950 3468 951
rect 3464 931 3466 950
rect 3463 930 3467 931
rect 3463 925 3467 926
rect 3464 906 3466 925
rect 3462 905 3468 906
rect 3462 901 3463 905
rect 3467 901 3468 905
rect 3462 900 3468 901
rect 3462 888 3468 889
rect 3462 884 3463 888
rect 3467 884 3468 888
rect 3462 883 3468 884
rect 3464 859 3466 883
rect 3463 858 3467 859
rect 3463 853 3467 854
rect 3438 851 3444 852
rect 3438 847 3439 851
rect 3443 847 3444 851
rect 3438 846 3444 847
rect 3464 837 3466 853
rect 3462 836 3468 837
rect 3366 835 3372 836
rect 3366 831 3367 835
rect 3371 831 3372 835
rect 3462 832 3463 836
rect 3467 832 3468 836
rect 3462 831 3468 832
rect 3366 830 3372 831
rect 3294 827 3300 828
rect 3294 823 3295 827
rect 3299 823 3300 827
rect 3294 822 3300 823
rect 3438 823 3444 824
rect 3438 819 3439 823
rect 3443 819 3444 823
rect 3438 818 3444 819
rect 3462 819 3468 820
rect 3222 816 3228 817
rect 3222 812 3223 816
rect 3227 812 3228 816
rect 3222 811 3228 812
rect 3366 816 3372 817
rect 3366 812 3367 816
rect 3371 812 3372 816
rect 3366 811 3372 812
rect 3224 791 3226 811
rect 3368 791 3370 811
rect 3215 790 3219 791
rect 3215 785 3219 786
rect 3223 790 3227 791
rect 3223 785 3227 786
rect 3367 790 3371 791
rect 3367 785 3371 786
rect 3216 769 3218 785
rect 3368 769 3370 785
rect 3214 768 3220 769
rect 3214 764 3215 768
rect 3219 764 3220 768
rect 3214 763 3220 764
rect 3366 768 3372 769
rect 3366 764 3367 768
rect 3371 764 3372 768
rect 3366 763 3372 764
rect 3430 759 3436 760
rect 3430 755 3431 759
rect 3435 755 3436 759
rect 3430 754 3436 755
rect 3214 749 3220 750
rect 3214 745 3215 749
rect 3219 745 3220 749
rect 3214 744 3220 745
rect 3366 749 3372 750
rect 3366 745 3367 749
rect 3371 745 3372 749
rect 3366 744 3372 745
rect 3216 727 3218 744
rect 3368 727 3370 744
rect 3215 726 3219 727
rect 3215 721 3219 722
rect 3255 726 3259 727
rect 3255 721 3259 722
rect 3367 726 3371 727
rect 3367 721 3371 722
rect 3198 719 3204 720
rect 3198 715 3199 719
rect 3203 715 3204 719
rect 3198 714 3204 715
rect 3200 696 3202 714
rect 3256 704 3258 721
rect 3302 719 3308 720
rect 3302 715 3303 719
rect 3307 715 3308 719
rect 3302 714 3314 715
rect 3304 713 3314 714
rect 3254 703 3260 704
rect 3254 699 3255 703
rect 3259 699 3260 703
rect 3254 698 3260 699
rect 2142 695 2148 696
rect 2142 691 2143 695
rect 2147 691 2148 695
rect 2142 690 2148 691
rect 2302 695 2308 696
rect 2302 691 2303 695
rect 2307 691 2308 695
rect 2302 690 2308 691
rect 2462 695 2468 696
rect 2462 691 2463 695
rect 2467 691 2468 695
rect 2462 690 2468 691
rect 2470 695 2476 696
rect 2470 691 2471 695
rect 2475 691 2476 695
rect 2470 690 2476 691
rect 2694 695 2700 696
rect 2694 691 2695 695
rect 2699 691 2700 695
rect 2694 690 2700 691
rect 2794 695 2800 696
rect 2794 691 2795 695
rect 2799 691 2800 695
rect 2794 690 2800 691
rect 3190 695 3196 696
rect 3190 691 3191 695
rect 3195 691 3196 695
rect 3190 690 3196 691
rect 3198 695 3204 696
rect 3198 691 3199 695
rect 3203 691 3204 695
rect 3198 690 3204 691
rect 2230 684 2236 685
rect 2230 680 2231 684
rect 2235 680 2236 684
rect 2230 679 2236 680
rect 2390 684 2396 685
rect 2390 680 2391 684
rect 2395 680 2396 684
rect 2390 679 2396 680
rect 2114 675 2120 676
rect 2114 671 2115 675
rect 2119 671 2120 675
rect 2114 670 2120 671
rect 2232 655 2234 679
rect 2392 655 2394 679
rect 2472 676 2474 690
rect 2550 684 2556 685
rect 2550 680 2551 684
rect 2555 680 2556 684
rect 2550 679 2556 680
rect 2470 675 2476 676
rect 2470 671 2471 675
rect 2475 671 2476 675
rect 2470 670 2476 671
rect 2398 667 2404 668
rect 2398 663 2399 667
rect 2403 663 2404 667
rect 2398 662 2404 663
rect 1311 654 1315 655
rect 1311 649 1315 650
rect 1343 654 1347 655
rect 1343 649 1347 650
rect 1447 654 1451 655
rect 1447 649 1451 650
rect 1503 654 1507 655
rect 1503 649 1507 650
rect 1583 654 1587 655
rect 1583 649 1587 650
rect 1767 654 1771 655
rect 1767 649 1771 650
rect 1807 654 1811 655
rect 1807 649 1811 650
rect 1831 654 1835 655
rect 1831 649 1835 650
rect 1927 654 1931 655
rect 1927 649 1931 650
rect 1967 654 1971 655
rect 1967 649 1971 650
rect 2071 654 2075 655
rect 2071 649 2075 650
rect 2135 654 2139 655
rect 2135 649 2139 650
rect 2231 654 2235 655
rect 2231 649 2235 650
rect 2311 654 2315 655
rect 2311 649 2315 650
rect 2391 654 2395 655
rect 2391 649 2395 650
rect 1312 633 1314 649
rect 1448 633 1450 649
rect 1584 633 1586 649
rect 1310 632 1316 633
rect 1310 628 1311 632
rect 1315 628 1316 632
rect 1310 627 1316 628
rect 1446 632 1452 633
rect 1446 628 1447 632
rect 1451 628 1452 632
rect 1446 627 1452 628
rect 1582 632 1588 633
rect 1582 628 1583 632
rect 1587 628 1588 632
rect 1768 630 1770 649
rect 1808 630 1810 649
rect 1832 633 1834 649
rect 1882 639 1888 640
rect 1882 635 1883 639
rect 1887 635 1888 639
rect 1882 634 1888 635
rect 1830 632 1836 633
rect 1582 627 1588 628
rect 1766 629 1772 630
rect 1766 625 1767 629
rect 1771 625 1772 629
rect 1766 624 1772 625
rect 1806 629 1812 630
rect 1806 625 1807 629
rect 1811 625 1812 629
rect 1830 628 1831 632
rect 1835 628 1836 632
rect 1830 627 1836 628
rect 1806 624 1812 625
rect 1382 623 1388 624
rect 1382 619 1383 623
rect 1387 619 1388 623
rect 1382 618 1388 619
rect 1518 623 1524 624
rect 1518 619 1519 623
rect 1523 619 1524 623
rect 1518 618 1524 619
rect 1646 623 1652 624
rect 1646 619 1647 623
rect 1651 619 1652 623
rect 1646 618 1652 619
rect 1310 613 1316 614
rect 1310 609 1311 613
rect 1315 609 1316 613
rect 1310 608 1316 609
rect 1254 595 1260 596
rect 1254 591 1255 595
rect 1259 591 1260 595
rect 1254 590 1260 591
rect 1312 583 1314 608
rect 1384 596 1386 618
rect 1446 613 1452 614
rect 1446 609 1447 613
rect 1451 609 1452 613
rect 1446 608 1452 609
rect 1382 595 1388 596
rect 1382 591 1383 595
rect 1387 591 1388 595
rect 1382 590 1388 591
rect 1448 583 1450 608
rect 1520 596 1522 618
rect 1582 613 1588 614
rect 1582 609 1583 613
rect 1587 609 1588 613
rect 1582 608 1588 609
rect 1518 595 1524 596
rect 1518 591 1519 595
rect 1523 591 1524 595
rect 1518 590 1524 591
rect 1584 583 1586 608
rect 1006 579 1007 583
rect 1011 579 1012 583
rect 1006 578 1012 579
rect 1039 582 1043 583
rect 990 575 996 576
rect 990 571 991 575
rect 995 571 996 575
rect 990 570 996 571
rect 998 575 1004 576
rect 998 571 999 575
rect 1003 571 1004 575
rect 998 570 1004 571
rect 814 559 820 560
rect 814 555 815 559
rect 819 555 820 559
rect 814 554 820 555
rect 926 559 932 560
rect 926 555 927 559
rect 931 555 932 559
rect 926 554 932 555
rect 1000 552 1002 570
rect 1008 552 1010 578
rect 1039 577 1043 578
rect 1055 582 1059 583
rect 1055 577 1059 578
rect 1151 582 1155 583
rect 1151 577 1155 578
rect 1183 582 1187 583
rect 1183 577 1187 578
rect 1255 582 1259 583
rect 1255 577 1259 578
rect 1311 582 1315 583
rect 1311 577 1315 578
rect 1359 582 1363 583
rect 1359 577 1363 578
rect 1447 582 1451 583
rect 1447 577 1451 578
rect 1471 582 1475 583
rect 1471 577 1475 578
rect 1583 582 1587 583
rect 1583 577 1587 578
rect 1040 560 1042 577
rect 1152 560 1154 577
rect 1198 575 1204 576
rect 1198 571 1199 575
rect 1203 571 1204 575
rect 1198 570 1204 571
rect 1222 575 1228 576
rect 1222 571 1223 575
rect 1227 571 1228 575
rect 1222 570 1228 571
rect 1038 559 1044 560
rect 1038 555 1039 559
rect 1043 555 1044 559
rect 1038 554 1044 555
rect 1150 559 1156 560
rect 1150 555 1151 559
rect 1155 555 1156 559
rect 1150 554 1156 555
rect 670 551 676 552
rect 670 547 671 551
rect 675 547 676 551
rect 670 546 676 547
rect 774 551 780 552
rect 774 547 775 551
rect 779 547 780 551
rect 998 551 1004 552
rect 774 546 780 547
rect 886 547 892 548
rect 110 543 116 544
rect 110 539 111 543
rect 115 539 116 543
rect 886 543 887 547
rect 891 543 892 547
rect 998 547 999 551
rect 1003 547 1004 551
rect 998 546 1004 547
rect 1006 551 1012 552
rect 1006 547 1007 551
rect 1011 547 1012 551
rect 1006 546 1012 547
rect 886 542 892 543
rect 110 538 116 539
rect 598 540 604 541
rect 112 519 114 538
rect 598 536 599 540
rect 603 536 604 540
rect 598 535 604 536
rect 702 540 708 541
rect 702 536 703 540
rect 707 536 708 540
rect 702 535 708 536
rect 814 540 820 541
rect 814 536 815 540
rect 819 536 820 540
rect 814 535 820 536
rect 600 519 602 535
rect 704 519 706 535
rect 816 519 818 535
rect 111 518 115 519
rect 111 513 115 514
rect 303 518 307 519
rect 303 513 307 514
rect 431 518 435 519
rect 431 513 435 514
rect 567 518 571 519
rect 567 513 571 514
rect 599 518 603 519
rect 599 513 603 514
rect 703 518 707 519
rect 703 513 707 514
rect 815 518 819 519
rect 815 513 819 514
rect 847 518 851 519
rect 847 513 851 514
rect 112 494 114 513
rect 304 497 306 513
rect 432 497 434 513
rect 568 497 570 513
rect 704 497 706 513
rect 848 497 850 513
rect 302 496 308 497
rect 110 493 116 494
rect 110 489 111 493
rect 115 489 116 493
rect 302 492 303 496
rect 307 492 308 496
rect 302 491 308 492
rect 430 496 436 497
rect 430 492 431 496
rect 435 492 436 496
rect 430 491 436 492
rect 566 496 572 497
rect 566 492 567 496
rect 571 492 572 496
rect 566 491 572 492
rect 702 496 708 497
rect 702 492 703 496
rect 707 492 708 496
rect 702 491 708 492
rect 846 496 852 497
rect 846 492 847 496
rect 851 492 852 496
rect 846 491 852 492
rect 110 488 116 489
rect 374 487 380 488
rect 374 483 375 487
rect 379 483 380 487
rect 374 482 380 483
rect 502 487 508 488
rect 502 483 503 487
rect 507 483 508 487
rect 502 482 508 483
rect 630 487 636 488
rect 630 483 631 487
rect 635 483 636 487
rect 630 482 636 483
rect 646 487 652 488
rect 646 483 647 487
rect 651 483 652 487
rect 646 482 652 483
rect 782 487 788 488
rect 782 483 783 487
rect 787 483 788 487
rect 782 482 788 483
rect 302 477 308 478
rect 110 476 116 477
rect 110 472 111 476
rect 115 472 116 476
rect 302 473 303 477
rect 307 473 308 477
rect 302 472 308 473
rect 110 471 116 472
rect 112 447 114 471
rect 304 447 306 472
rect 376 460 378 482
rect 430 477 436 478
rect 430 473 431 477
rect 435 473 436 477
rect 430 472 436 473
rect 374 459 380 460
rect 374 455 375 459
rect 379 455 380 459
rect 374 454 380 455
rect 432 447 434 472
rect 504 460 506 482
rect 566 477 572 478
rect 566 473 567 477
rect 571 473 572 477
rect 566 472 572 473
rect 502 459 508 460
rect 502 455 503 459
rect 507 455 508 459
rect 502 454 508 455
rect 568 447 570 472
rect 111 446 115 447
rect 111 441 115 442
rect 135 446 139 447
rect 135 441 139 442
rect 255 446 259 447
rect 255 441 259 442
rect 303 446 307 447
rect 303 441 307 442
rect 415 446 419 447
rect 415 441 419 442
rect 431 446 435 447
rect 431 441 435 442
rect 567 446 571 447
rect 567 441 571 442
rect 583 446 587 447
rect 583 441 587 442
rect 112 425 114 441
rect 110 424 116 425
rect 136 424 138 441
rect 214 439 220 440
rect 214 435 215 439
rect 219 435 220 439
rect 214 434 220 435
rect 110 420 111 424
rect 115 420 116 424
rect 110 419 116 420
rect 134 423 140 424
rect 134 419 135 423
rect 139 419 140 423
rect 134 418 140 419
rect 216 416 218 434
rect 256 424 258 441
rect 386 439 392 440
rect 386 435 387 439
rect 391 435 392 439
rect 386 434 392 435
rect 254 423 260 424
rect 254 419 255 423
rect 259 419 260 423
rect 254 418 260 419
rect 388 416 390 434
rect 416 424 418 441
rect 584 424 586 441
rect 632 440 634 482
rect 648 456 650 482
rect 702 477 708 478
rect 702 473 703 477
rect 707 473 708 477
rect 702 472 708 473
rect 646 455 652 456
rect 646 451 647 455
rect 651 451 652 455
rect 646 450 652 451
rect 678 447 684 448
rect 704 447 706 472
rect 784 460 786 482
rect 846 477 852 478
rect 846 473 847 477
rect 851 473 852 477
rect 846 472 852 473
rect 782 459 788 460
rect 782 455 783 459
rect 787 455 788 459
rect 782 454 788 455
rect 848 447 850 472
rect 888 460 890 542
rect 926 540 932 541
rect 926 536 927 540
rect 931 536 932 540
rect 926 535 932 536
rect 1038 540 1044 541
rect 1038 536 1039 540
rect 1043 536 1044 540
rect 1038 535 1044 536
rect 1150 540 1156 541
rect 1150 536 1151 540
rect 1155 536 1156 540
rect 1150 535 1156 536
rect 928 519 930 535
rect 1040 519 1042 535
rect 1152 519 1154 535
rect 927 518 931 519
rect 927 513 931 514
rect 983 518 987 519
rect 983 513 987 514
rect 1039 518 1043 519
rect 1039 513 1043 514
rect 1111 518 1115 519
rect 1111 513 1115 514
rect 1151 518 1155 519
rect 1151 513 1155 514
rect 984 497 986 513
rect 1112 497 1114 513
rect 982 496 988 497
rect 982 492 983 496
rect 987 492 988 496
rect 982 491 988 492
rect 1110 496 1116 497
rect 1110 492 1111 496
rect 1115 492 1116 496
rect 1110 491 1116 492
rect 1200 488 1202 570
rect 1224 552 1226 570
rect 1256 560 1258 577
rect 1360 560 1362 577
rect 1438 575 1444 576
rect 1438 571 1439 575
rect 1443 571 1444 575
rect 1438 570 1444 571
rect 1254 559 1260 560
rect 1254 555 1255 559
rect 1259 555 1260 559
rect 1254 554 1260 555
rect 1358 559 1364 560
rect 1358 555 1359 559
rect 1363 555 1364 559
rect 1358 554 1364 555
rect 1440 552 1442 570
rect 1472 560 1474 577
rect 1550 575 1556 576
rect 1550 571 1551 575
rect 1555 571 1556 575
rect 1550 570 1556 571
rect 1470 559 1476 560
rect 1470 555 1471 559
rect 1475 555 1476 559
rect 1470 554 1476 555
rect 1552 552 1554 570
rect 1584 560 1586 577
rect 1648 576 1650 618
rect 1830 613 1836 614
rect 1766 612 1772 613
rect 1766 608 1767 612
rect 1771 608 1772 612
rect 1766 607 1772 608
rect 1806 612 1812 613
rect 1806 608 1807 612
rect 1811 608 1812 612
rect 1830 609 1831 613
rect 1835 609 1836 613
rect 1830 608 1836 609
rect 1806 607 1812 608
rect 1742 583 1748 584
rect 1768 583 1770 607
rect 1808 591 1810 607
rect 1832 591 1834 608
rect 1884 596 1886 634
rect 1968 633 1970 649
rect 2136 633 2138 649
rect 2238 639 2244 640
rect 2238 635 2239 639
rect 2243 635 2244 639
rect 2238 634 2244 635
rect 1966 632 1972 633
rect 1966 628 1967 632
rect 1971 628 1972 632
rect 1966 627 1972 628
rect 2134 632 2140 633
rect 2134 628 2135 632
rect 2139 628 2140 632
rect 2134 627 2140 628
rect 1902 623 1908 624
rect 1902 619 1903 623
rect 1907 619 1908 623
rect 1902 618 1908 619
rect 2038 623 2044 624
rect 2038 619 2039 623
rect 2043 619 2044 623
rect 2038 618 2044 619
rect 2206 623 2212 624
rect 2206 619 2207 623
rect 2211 619 2212 623
rect 2206 618 2212 619
rect 1904 596 1906 618
rect 1966 613 1972 614
rect 1966 609 1967 613
rect 1971 609 1972 613
rect 1966 608 1972 609
rect 1882 595 1888 596
rect 1882 591 1883 595
rect 1887 591 1888 595
rect 1807 590 1811 591
rect 1807 585 1811 586
rect 1831 590 1835 591
rect 1882 590 1888 591
rect 1902 595 1908 596
rect 1902 591 1903 595
rect 1907 591 1908 595
rect 1968 591 1970 608
rect 2040 596 2042 618
rect 2134 613 2140 614
rect 2134 609 2135 613
rect 2139 609 2140 613
rect 2134 608 2140 609
rect 2038 595 2044 596
rect 2038 591 2039 595
rect 2043 591 2044 595
rect 2136 591 2138 608
rect 2208 596 2210 618
rect 2206 595 2212 596
rect 2206 591 2207 595
rect 2211 591 2212 595
rect 1902 590 1908 591
rect 1967 590 1971 591
rect 2038 590 2044 591
rect 2127 590 2131 591
rect 1831 585 1835 586
rect 1967 585 1971 586
rect 2127 585 2131 586
rect 2135 590 2139 591
rect 2206 590 2212 591
rect 2135 585 2139 586
rect 1671 582 1675 583
rect 1742 579 1743 583
rect 1747 579 1748 583
rect 1742 578 1748 579
rect 1767 582 1771 583
rect 1671 577 1675 578
rect 1646 575 1652 576
rect 1646 571 1647 575
rect 1651 571 1652 575
rect 1646 570 1652 571
rect 1672 560 1674 577
rect 1734 575 1740 576
rect 1734 571 1735 575
rect 1739 571 1740 575
rect 1734 570 1740 571
rect 1582 559 1588 560
rect 1582 555 1583 559
rect 1587 555 1588 559
rect 1582 554 1588 555
rect 1670 559 1676 560
rect 1670 555 1671 559
rect 1675 555 1676 559
rect 1670 554 1676 555
rect 1222 551 1228 552
rect 1222 547 1223 551
rect 1227 547 1228 551
rect 1222 546 1228 547
rect 1438 551 1444 552
rect 1438 547 1439 551
rect 1443 547 1444 551
rect 1438 546 1444 547
rect 1550 551 1556 552
rect 1550 547 1551 551
rect 1555 547 1556 551
rect 1550 546 1556 547
rect 1254 540 1260 541
rect 1254 536 1255 540
rect 1259 536 1260 540
rect 1254 535 1260 536
rect 1358 540 1364 541
rect 1358 536 1359 540
rect 1363 536 1364 540
rect 1358 535 1364 536
rect 1470 540 1476 541
rect 1470 536 1471 540
rect 1475 536 1476 540
rect 1470 535 1476 536
rect 1582 540 1588 541
rect 1582 536 1583 540
rect 1587 536 1588 540
rect 1582 535 1588 536
rect 1670 540 1676 541
rect 1670 536 1671 540
rect 1675 536 1676 540
rect 1670 535 1676 536
rect 1256 519 1258 535
rect 1360 519 1362 535
rect 1472 519 1474 535
rect 1584 519 1586 535
rect 1672 519 1674 535
rect 1231 518 1235 519
rect 1231 513 1235 514
rect 1255 518 1259 519
rect 1255 513 1259 514
rect 1351 518 1355 519
rect 1351 513 1355 514
rect 1359 518 1363 519
rect 1359 513 1363 514
rect 1463 518 1467 519
rect 1463 513 1467 514
rect 1471 518 1475 519
rect 1471 513 1475 514
rect 1575 518 1579 519
rect 1575 513 1579 514
rect 1583 518 1587 519
rect 1583 513 1587 514
rect 1671 518 1675 519
rect 1671 513 1675 514
rect 1232 497 1234 513
rect 1352 497 1354 513
rect 1464 497 1466 513
rect 1576 497 1578 513
rect 1672 497 1674 513
rect 1230 496 1236 497
rect 1230 492 1231 496
rect 1235 492 1236 496
rect 1230 491 1236 492
rect 1350 496 1356 497
rect 1350 492 1351 496
rect 1355 492 1356 496
rect 1350 491 1356 492
rect 1462 496 1468 497
rect 1462 492 1463 496
rect 1467 492 1468 496
rect 1462 491 1468 492
rect 1574 496 1580 497
rect 1574 492 1575 496
rect 1579 492 1580 496
rect 1574 491 1580 492
rect 1670 496 1676 497
rect 1670 492 1671 496
rect 1675 492 1676 496
rect 1670 491 1676 492
rect 1736 488 1738 570
rect 1744 552 1746 578
rect 1767 577 1771 578
rect 1768 561 1770 577
rect 1808 569 1810 585
rect 1806 568 1812 569
rect 1832 568 1834 585
rect 1902 583 1908 584
rect 1902 579 1903 583
rect 1907 579 1908 583
rect 1902 578 1908 579
rect 1806 564 1807 568
rect 1811 564 1812 568
rect 1806 563 1812 564
rect 1830 567 1836 568
rect 1830 563 1831 567
rect 1835 563 1836 567
rect 1830 562 1836 563
rect 1766 560 1772 561
rect 1904 560 1906 578
rect 1968 568 1970 585
rect 2038 583 2044 584
rect 2038 579 2039 583
rect 2043 579 2044 583
rect 2038 578 2044 579
rect 1966 567 1972 568
rect 1966 563 1967 567
rect 1971 563 1972 567
rect 1966 562 1972 563
rect 2040 560 2042 578
rect 2128 568 2130 585
rect 2198 583 2204 584
rect 2198 579 2199 583
rect 2203 579 2204 583
rect 2198 578 2204 579
rect 2126 567 2132 568
rect 2126 563 2127 567
rect 2131 563 2132 567
rect 2126 562 2132 563
rect 2200 560 2202 578
rect 2240 560 2242 634
rect 2312 633 2314 649
rect 2310 632 2316 633
rect 2310 628 2311 632
rect 2315 628 2316 632
rect 2310 627 2316 628
rect 2400 624 2402 662
rect 2552 655 2554 679
rect 2487 654 2491 655
rect 2487 649 2491 650
rect 2551 654 2555 655
rect 2551 649 2555 650
rect 2655 654 2659 655
rect 2655 649 2659 650
rect 2488 633 2490 649
rect 2506 639 2512 640
rect 2506 635 2507 639
rect 2511 635 2512 639
rect 2506 634 2512 635
rect 2486 632 2492 633
rect 2486 628 2487 632
rect 2491 628 2492 632
rect 2486 627 2492 628
rect 2382 623 2388 624
rect 2382 619 2383 623
rect 2387 619 2388 623
rect 2382 618 2388 619
rect 2398 623 2404 624
rect 2398 619 2399 623
rect 2403 619 2404 623
rect 2398 618 2404 619
rect 2310 613 2316 614
rect 2310 609 2311 613
rect 2315 609 2316 613
rect 2310 608 2316 609
rect 2312 591 2314 608
rect 2384 596 2386 618
rect 2486 613 2492 614
rect 2486 609 2487 613
rect 2491 609 2492 613
rect 2486 608 2492 609
rect 2382 595 2388 596
rect 2382 591 2383 595
rect 2387 591 2388 595
rect 2488 591 2490 608
rect 2287 590 2291 591
rect 2287 585 2291 586
rect 2311 590 2315 591
rect 2382 590 2388 591
rect 2455 590 2459 591
rect 2311 585 2315 586
rect 2455 585 2459 586
rect 2487 590 2491 591
rect 2487 585 2491 586
rect 2288 568 2290 585
rect 2456 568 2458 585
rect 2508 584 2510 634
rect 2656 633 2658 649
rect 2654 632 2660 633
rect 2654 628 2655 632
rect 2659 628 2660 632
rect 2654 627 2660 628
rect 2654 613 2660 614
rect 2654 609 2655 613
rect 2659 609 2660 613
rect 2654 608 2660 609
rect 2656 591 2658 608
rect 2696 596 2698 690
rect 2702 684 2708 685
rect 2702 680 2703 684
rect 2707 680 2708 684
rect 2702 679 2708 680
rect 2846 684 2852 685
rect 2846 680 2847 684
rect 2851 680 2852 684
rect 2846 679 2852 680
rect 2982 684 2988 685
rect 2982 680 2983 684
rect 2987 680 2988 684
rect 2982 679 2988 680
rect 3118 684 3124 685
rect 3118 680 3119 684
rect 3123 680 3124 684
rect 3118 679 3124 680
rect 3254 684 3260 685
rect 3254 680 3255 684
rect 3259 680 3260 684
rect 3254 679 3260 680
rect 2704 655 2706 679
rect 2848 655 2850 679
rect 2984 655 2986 679
rect 3120 655 3122 679
rect 3256 655 3258 679
rect 2703 654 2707 655
rect 2703 649 2707 650
rect 2815 654 2819 655
rect 2815 649 2819 650
rect 2847 654 2851 655
rect 2847 649 2851 650
rect 2959 654 2963 655
rect 2959 649 2963 650
rect 2983 654 2987 655
rect 2983 649 2987 650
rect 3103 654 3107 655
rect 3103 649 3107 650
rect 3119 654 3123 655
rect 3119 649 3123 650
rect 3247 654 3251 655
rect 3247 649 3251 650
rect 3255 654 3259 655
rect 3255 649 3259 650
rect 2816 633 2818 649
rect 2918 639 2924 640
rect 2918 635 2919 639
rect 2923 635 2924 639
rect 2918 634 2924 635
rect 2814 632 2820 633
rect 2814 628 2815 632
rect 2819 628 2820 632
rect 2814 627 2820 628
rect 2726 623 2732 624
rect 2726 619 2727 623
rect 2731 619 2732 623
rect 2726 618 2732 619
rect 2886 623 2892 624
rect 2886 619 2887 623
rect 2891 619 2892 623
rect 2886 618 2892 619
rect 2728 596 2730 618
rect 2814 613 2820 614
rect 2814 609 2815 613
rect 2819 609 2820 613
rect 2814 608 2820 609
rect 2694 595 2700 596
rect 2694 591 2695 595
rect 2699 591 2700 595
rect 2623 590 2627 591
rect 2623 585 2627 586
rect 2655 590 2659 591
rect 2694 590 2700 591
rect 2726 595 2732 596
rect 2726 591 2727 595
rect 2731 591 2732 595
rect 2816 591 2818 608
rect 2888 596 2890 618
rect 2886 595 2892 596
rect 2886 591 2887 595
rect 2891 591 2892 595
rect 2726 590 2732 591
rect 2799 590 2803 591
rect 2655 585 2659 586
rect 2799 585 2803 586
rect 2815 590 2819 591
rect 2886 590 2892 591
rect 2815 585 2819 586
rect 2506 583 2512 584
rect 2506 579 2507 583
rect 2511 579 2512 583
rect 2506 578 2512 579
rect 2526 583 2532 584
rect 2526 579 2527 583
rect 2531 579 2532 583
rect 2526 578 2532 579
rect 2286 567 2292 568
rect 2286 563 2287 567
rect 2291 563 2292 567
rect 2286 562 2292 563
rect 2454 567 2460 568
rect 2454 563 2455 567
rect 2459 563 2460 567
rect 2454 562 2460 563
rect 2528 560 2530 578
rect 2624 568 2626 585
rect 2694 583 2700 584
rect 2694 579 2695 583
rect 2699 579 2700 583
rect 2694 578 2700 579
rect 2622 567 2628 568
rect 2622 563 2623 567
rect 2627 563 2628 567
rect 2622 562 2628 563
rect 2696 560 2698 578
rect 2800 568 2802 585
rect 2798 567 2804 568
rect 2798 563 2799 567
rect 2803 563 2804 567
rect 2798 562 2804 563
rect 2920 560 2922 634
rect 2960 633 2962 649
rect 3104 633 3106 649
rect 3248 633 3250 649
rect 2958 632 2964 633
rect 2958 628 2959 632
rect 2963 628 2964 632
rect 2958 627 2964 628
rect 3102 632 3108 633
rect 3102 628 3103 632
rect 3107 628 3108 632
rect 3102 627 3108 628
rect 3246 632 3252 633
rect 3246 628 3247 632
rect 3251 628 3252 632
rect 3246 627 3252 628
rect 3312 624 3314 713
rect 3368 704 3370 721
rect 3432 720 3434 754
rect 3440 732 3442 818
rect 3462 815 3463 819
rect 3467 815 3468 819
rect 3462 814 3468 815
rect 3464 791 3466 814
rect 3463 790 3467 791
rect 3463 785 3467 786
rect 3464 766 3466 785
rect 3462 765 3468 766
rect 3462 761 3463 765
rect 3467 761 3468 765
rect 3462 760 3468 761
rect 3462 748 3468 749
rect 3462 744 3463 748
rect 3467 744 3468 748
rect 3462 743 3468 744
rect 3438 731 3444 732
rect 3438 727 3439 731
rect 3443 727 3444 731
rect 3464 727 3466 743
rect 3438 726 3444 727
rect 3463 726 3467 727
rect 3463 721 3467 722
rect 3430 719 3436 720
rect 3430 715 3431 719
rect 3435 715 3436 719
rect 3430 714 3436 715
rect 3464 705 3466 721
rect 3462 704 3468 705
rect 3366 703 3372 704
rect 3366 699 3367 703
rect 3371 699 3372 703
rect 3462 700 3463 704
rect 3467 700 3468 704
rect 3462 699 3468 700
rect 3366 698 3372 699
rect 3438 691 3444 692
rect 3438 687 3439 691
rect 3443 687 3444 691
rect 3438 686 3444 687
rect 3462 687 3468 688
rect 3366 684 3372 685
rect 3366 680 3367 684
rect 3371 680 3372 684
rect 3366 679 3372 680
rect 3368 655 3370 679
rect 3367 654 3371 655
rect 3367 649 3371 650
rect 3368 633 3370 649
rect 3366 632 3372 633
rect 3366 628 3367 632
rect 3371 628 3372 632
rect 3366 627 3372 628
rect 3030 623 3036 624
rect 3030 619 3031 623
rect 3035 619 3036 623
rect 3030 618 3036 619
rect 3174 623 3180 624
rect 3174 619 3175 623
rect 3179 619 3180 623
rect 3174 618 3180 619
rect 3310 623 3316 624
rect 3310 619 3311 623
rect 3315 619 3316 623
rect 3310 618 3316 619
rect 3430 623 3436 624
rect 3430 619 3431 623
rect 3435 619 3436 623
rect 3430 618 3436 619
rect 2958 613 2964 614
rect 2958 609 2959 613
rect 2963 609 2964 613
rect 2958 608 2964 609
rect 2960 591 2962 608
rect 3032 596 3034 618
rect 3102 613 3108 614
rect 3102 609 3103 613
rect 3107 609 3108 613
rect 3102 608 3108 609
rect 3030 595 3036 596
rect 3030 591 3031 595
rect 3035 591 3036 595
rect 3104 591 3106 608
rect 2959 590 2963 591
rect 2959 585 2963 586
rect 2983 590 2987 591
rect 3030 590 3036 591
rect 3103 590 3107 591
rect 2983 585 2987 586
rect 3103 585 3107 586
rect 3167 590 3171 591
rect 3167 585 3171 586
rect 2984 568 2986 585
rect 3062 583 3068 584
rect 3062 579 3063 583
rect 3067 579 3068 583
rect 3062 578 3068 579
rect 2982 567 2988 568
rect 2982 563 2983 567
rect 2987 563 2988 567
rect 2982 562 2988 563
rect 3064 560 3066 578
rect 3168 568 3170 585
rect 3176 584 3178 618
rect 3246 613 3252 614
rect 3246 609 3247 613
rect 3251 609 3252 613
rect 3246 608 3252 609
rect 3366 613 3372 614
rect 3366 609 3367 613
rect 3371 609 3372 613
rect 3366 608 3372 609
rect 3248 591 3250 608
rect 3318 595 3324 596
rect 3318 591 3319 595
rect 3323 591 3324 595
rect 3368 591 3370 608
rect 3247 590 3251 591
rect 3318 590 3324 591
rect 3359 590 3363 591
rect 3247 585 3251 586
rect 3174 583 3180 584
rect 3174 579 3175 583
rect 3179 579 3180 583
rect 3174 578 3180 579
rect 3166 567 3172 568
rect 3166 563 3167 567
rect 3171 563 3172 567
rect 3166 562 3172 563
rect 1766 556 1767 560
rect 1771 556 1772 560
rect 1766 555 1772 556
rect 1902 559 1908 560
rect 1902 555 1903 559
rect 1907 555 1908 559
rect 1902 554 1908 555
rect 2038 559 2044 560
rect 2038 555 2039 559
rect 2043 555 2044 559
rect 2038 554 2044 555
rect 2198 559 2204 560
rect 2198 555 2199 559
rect 2203 555 2204 559
rect 2198 554 2204 555
rect 2238 559 2244 560
rect 2238 555 2239 559
rect 2243 555 2244 559
rect 2238 554 2244 555
rect 2526 559 2532 560
rect 2526 555 2527 559
rect 2531 555 2532 559
rect 2526 554 2532 555
rect 2694 559 2700 560
rect 2694 555 2695 559
rect 2699 555 2700 559
rect 2918 559 2924 560
rect 2694 554 2700 555
rect 2878 555 2884 556
rect 1742 551 1748 552
rect 1742 547 1743 551
rect 1747 547 1748 551
rect 1742 546 1748 547
rect 1806 551 1812 552
rect 1806 547 1807 551
rect 1811 547 1812 551
rect 2878 551 2879 555
rect 2883 551 2884 555
rect 2918 555 2919 559
rect 2923 555 2924 559
rect 2918 554 2924 555
rect 3062 559 3068 560
rect 3062 555 3063 559
rect 3067 555 3068 559
rect 3062 554 3068 555
rect 2878 550 2884 551
rect 1806 546 1812 547
rect 1830 548 1836 549
rect 1766 543 1772 544
rect 1766 539 1767 543
rect 1771 539 1772 543
rect 1766 538 1772 539
rect 1768 519 1770 538
rect 1767 518 1771 519
rect 1767 513 1771 514
rect 1768 494 1770 513
rect 1808 511 1810 546
rect 1830 544 1831 548
rect 1835 544 1836 548
rect 1830 543 1836 544
rect 1966 548 1972 549
rect 1966 544 1967 548
rect 1971 544 1972 548
rect 1966 543 1972 544
rect 2126 548 2132 549
rect 2126 544 2127 548
rect 2131 544 2132 548
rect 2126 543 2132 544
rect 2286 548 2292 549
rect 2286 544 2287 548
rect 2291 544 2292 548
rect 2286 543 2292 544
rect 2454 548 2460 549
rect 2454 544 2455 548
rect 2459 544 2460 548
rect 2454 543 2460 544
rect 2622 548 2628 549
rect 2622 544 2623 548
rect 2627 544 2628 548
rect 2622 543 2628 544
rect 2798 548 2804 549
rect 2798 544 2799 548
rect 2803 544 2804 548
rect 2798 543 2804 544
rect 1832 511 1834 543
rect 1968 511 1970 543
rect 2128 511 2130 543
rect 2288 511 2290 543
rect 2456 511 2458 543
rect 2624 511 2626 543
rect 2800 511 2802 543
rect 1807 510 1811 511
rect 1807 505 1811 506
rect 1831 510 1835 511
rect 1831 505 1835 506
rect 1967 510 1971 511
rect 1967 505 1971 506
rect 2127 510 2131 511
rect 2127 505 2131 506
rect 2287 510 2291 511
rect 2287 505 2291 506
rect 2295 510 2299 511
rect 2295 505 2299 506
rect 2455 510 2459 511
rect 2455 505 2459 506
rect 2479 510 2483 511
rect 2479 505 2483 506
rect 2623 510 2627 511
rect 2623 505 2627 506
rect 2679 510 2683 511
rect 2679 505 2683 506
rect 2799 510 2803 511
rect 2799 505 2803 506
rect 1766 493 1772 494
rect 1766 489 1767 493
rect 1771 489 1772 493
rect 1766 488 1772 489
rect 1054 487 1060 488
rect 1054 483 1055 487
rect 1059 483 1060 487
rect 1054 482 1060 483
rect 1198 487 1204 488
rect 1198 483 1199 487
rect 1203 483 1204 487
rect 1198 482 1204 483
rect 1302 487 1308 488
rect 1302 483 1303 487
rect 1307 483 1308 487
rect 1302 482 1308 483
rect 1310 487 1316 488
rect 1310 483 1311 487
rect 1315 483 1316 487
rect 1310 482 1316 483
rect 1430 487 1436 488
rect 1430 483 1431 487
rect 1435 483 1436 487
rect 1430 482 1436 483
rect 1734 487 1740 488
rect 1734 483 1735 487
rect 1739 483 1740 487
rect 1808 486 1810 505
rect 1832 489 1834 505
rect 1882 495 1888 496
rect 1882 491 1883 495
rect 1887 491 1888 495
rect 1882 490 1888 491
rect 1830 488 1836 489
rect 1734 482 1740 483
rect 1806 485 1812 486
rect 982 477 988 478
rect 982 473 983 477
rect 987 473 988 477
rect 982 472 988 473
rect 886 459 892 460
rect 886 455 887 459
rect 891 455 892 459
rect 886 454 892 455
rect 974 459 980 460
rect 974 455 975 459
rect 979 455 980 459
rect 974 454 980 455
rect 678 443 679 447
rect 683 443 684 447
rect 678 442 684 443
rect 703 446 707 447
rect 630 439 636 440
rect 630 435 631 439
rect 635 435 636 439
rect 630 434 636 435
rect 654 439 660 440
rect 654 435 655 439
rect 659 435 660 439
rect 654 434 660 435
rect 414 423 420 424
rect 414 419 415 423
rect 419 419 420 423
rect 414 418 420 419
rect 582 423 588 424
rect 582 419 583 423
rect 587 419 588 423
rect 582 418 588 419
rect 656 416 658 434
rect 680 416 682 442
rect 703 441 707 442
rect 743 446 747 447
rect 743 441 747 442
rect 847 446 851 447
rect 847 441 851 442
rect 903 446 907 447
rect 903 441 907 442
rect 744 424 746 441
rect 904 424 906 441
rect 742 423 748 424
rect 742 419 743 423
rect 747 419 748 423
rect 742 418 748 419
rect 902 423 908 424
rect 902 419 903 423
rect 907 419 908 423
rect 902 418 908 419
rect 976 416 978 454
rect 984 447 986 472
rect 1056 460 1058 482
rect 1110 477 1116 478
rect 1110 473 1111 477
rect 1115 473 1116 477
rect 1110 472 1116 473
rect 1230 477 1236 478
rect 1230 473 1231 477
rect 1235 473 1236 477
rect 1230 472 1236 473
rect 1054 459 1060 460
rect 1054 455 1055 459
rect 1059 455 1060 459
rect 1054 454 1060 455
rect 1112 447 1114 472
rect 1232 447 1234 472
rect 983 446 987 447
rect 983 441 987 442
rect 1047 446 1051 447
rect 1047 441 1051 442
rect 1111 446 1115 447
rect 1111 441 1115 442
rect 1183 446 1187 447
rect 1183 441 1187 442
rect 1231 446 1235 447
rect 1231 441 1235 442
rect 1048 424 1050 441
rect 1126 439 1132 440
rect 1126 435 1127 439
rect 1131 435 1132 439
rect 1126 434 1132 435
rect 1046 423 1052 424
rect 1046 419 1047 423
rect 1051 419 1052 423
rect 1046 418 1052 419
rect 1128 416 1130 434
rect 1184 424 1186 441
rect 1304 440 1306 482
rect 1312 460 1314 482
rect 1350 477 1356 478
rect 1350 473 1351 477
rect 1355 473 1356 477
rect 1350 472 1356 473
rect 1310 459 1316 460
rect 1310 455 1311 459
rect 1315 455 1316 459
rect 1310 454 1316 455
rect 1352 447 1354 472
rect 1432 460 1434 482
rect 1806 481 1807 485
rect 1811 481 1812 485
rect 1830 484 1831 488
rect 1835 484 1836 488
rect 1830 483 1836 484
rect 1806 480 1812 481
rect 1774 479 1780 480
rect 1462 477 1468 478
rect 1462 473 1463 477
rect 1467 473 1468 477
rect 1462 472 1468 473
rect 1574 477 1580 478
rect 1574 473 1575 477
rect 1579 473 1580 477
rect 1574 472 1580 473
rect 1670 477 1676 478
rect 1670 473 1671 477
rect 1675 473 1676 477
rect 1670 472 1676 473
rect 1766 476 1772 477
rect 1766 472 1767 476
rect 1771 472 1772 476
rect 1774 475 1775 479
rect 1779 475 1780 479
rect 1774 474 1780 475
rect 1430 459 1436 460
rect 1430 455 1431 459
rect 1435 455 1436 459
rect 1430 454 1436 455
rect 1464 447 1466 472
rect 1576 447 1578 472
rect 1672 447 1674 472
rect 1766 471 1772 472
rect 1768 447 1770 471
rect 1776 452 1778 474
rect 1830 469 1836 470
rect 1806 468 1812 469
rect 1806 464 1807 468
rect 1811 464 1812 468
rect 1830 465 1831 469
rect 1835 465 1836 469
rect 1830 464 1836 465
rect 1806 463 1812 464
rect 1774 451 1780 452
rect 1774 447 1775 451
rect 1779 447 1780 451
rect 1808 447 1810 463
rect 1832 447 1834 464
rect 1884 452 1886 490
rect 1968 489 1970 505
rect 2128 489 2130 505
rect 2296 489 2298 505
rect 2480 489 2482 505
rect 2680 489 2682 505
rect 2730 495 2736 496
rect 2730 491 2731 495
rect 2735 491 2736 495
rect 2730 490 2736 491
rect 1966 488 1972 489
rect 1966 484 1967 488
rect 1971 484 1972 488
rect 1966 483 1972 484
rect 2126 488 2132 489
rect 2126 484 2127 488
rect 2131 484 2132 488
rect 2126 483 2132 484
rect 2294 488 2300 489
rect 2294 484 2295 488
rect 2299 484 2300 488
rect 2294 483 2300 484
rect 2478 488 2484 489
rect 2478 484 2479 488
rect 2483 484 2484 488
rect 2478 483 2484 484
rect 2678 488 2684 489
rect 2678 484 2679 488
rect 2683 484 2684 488
rect 2678 483 2684 484
rect 2038 479 2044 480
rect 2038 475 2039 479
rect 2043 475 2044 479
rect 2038 474 2044 475
rect 2358 479 2364 480
rect 2358 475 2359 479
rect 2363 475 2364 479
rect 2358 474 2364 475
rect 2374 479 2380 480
rect 2374 475 2375 479
rect 2379 475 2380 479
rect 2374 474 2380 475
rect 2558 479 2564 480
rect 2558 475 2559 479
rect 2563 475 2564 479
rect 2558 474 2564 475
rect 1966 469 1972 470
rect 1966 465 1967 469
rect 1971 465 1972 469
rect 1966 464 1972 465
rect 1882 451 1888 452
rect 1882 447 1883 451
rect 1887 447 1888 451
rect 1968 447 1970 464
rect 2040 452 2042 474
rect 2126 469 2132 470
rect 2126 465 2127 469
rect 2131 465 2132 469
rect 2126 464 2132 465
rect 2294 469 2300 470
rect 2294 465 2295 469
rect 2299 465 2300 469
rect 2294 464 2300 465
rect 2030 451 2036 452
rect 2030 447 2031 451
rect 2035 447 2036 451
rect 1311 446 1315 447
rect 1311 441 1315 442
rect 1351 446 1355 447
rect 1351 441 1355 442
rect 1439 446 1443 447
rect 1439 441 1443 442
rect 1463 446 1467 447
rect 1463 441 1467 442
rect 1567 446 1571 447
rect 1567 441 1571 442
rect 1575 446 1579 447
rect 1575 441 1579 442
rect 1671 446 1675 447
rect 1671 441 1675 442
rect 1767 446 1771 447
rect 1774 446 1780 447
rect 1807 446 1811 447
rect 1767 441 1771 442
rect 1807 441 1811 442
rect 1831 446 1835 447
rect 1882 446 1888 447
rect 1959 446 1963 447
rect 1831 441 1835 442
rect 1959 441 1963 442
rect 1967 446 1971 447
rect 2030 446 2036 447
rect 2038 451 2044 452
rect 2038 447 2039 451
rect 2043 447 2044 451
rect 2128 447 2130 464
rect 2296 447 2298 464
rect 2038 446 2044 447
rect 2111 446 2115 447
rect 1967 441 1971 442
rect 1294 439 1300 440
rect 1294 435 1295 439
rect 1299 435 1300 439
rect 1294 434 1300 435
rect 1302 439 1308 440
rect 1302 435 1303 439
rect 1307 435 1308 439
rect 1302 434 1308 435
rect 1182 423 1188 424
rect 1182 419 1183 423
rect 1187 419 1188 423
rect 1182 418 1188 419
rect 214 415 220 416
rect 214 411 215 415
rect 219 411 220 415
rect 214 410 220 411
rect 386 415 392 416
rect 386 411 387 415
rect 391 411 392 415
rect 386 410 392 411
rect 654 415 660 416
rect 654 411 655 415
rect 659 411 660 415
rect 654 410 660 411
rect 678 415 684 416
rect 678 411 679 415
rect 683 411 684 415
rect 678 410 684 411
rect 974 415 980 416
rect 974 411 975 415
rect 979 411 980 415
rect 974 410 980 411
rect 1126 415 1132 416
rect 1126 411 1127 415
rect 1131 411 1132 415
rect 1126 410 1132 411
rect 110 407 116 408
rect 110 403 111 407
rect 115 403 116 407
rect 198 407 204 408
rect 110 402 116 403
rect 134 404 140 405
rect 112 379 114 402
rect 134 400 135 404
rect 139 400 140 404
rect 198 403 199 407
rect 203 403 204 407
rect 198 402 204 403
rect 254 404 260 405
rect 134 399 140 400
rect 136 379 138 399
rect 111 378 115 379
rect 111 373 115 374
rect 135 378 139 379
rect 135 373 139 374
rect 112 354 114 373
rect 136 357 138 373
rect 134 356 140 357
rect 110 353 116 354
rect 110 349 111 353
rect 115 349 116 353
rect 134 352 135 356
rect 139 352 140 356
rect 134 351 140 352
rect 110 348 116 349
rect 134 337 140 338
rect 110 336 116 337
rect 110 332 111 336
rect 115 332 116 336
rect 134 333 135 337
rect 139 333 140 337
rect 134 332 140 333
rect 110 331 116 332
rect 112 311 114 331
rect 136 311 138 332
rect 200 320 202 402
rect 254 400 255 404
rect 259 400 260 404
rect 254 399 260 400
rect 414 404 420 405
rect 414 400 415 404
rect 419 400 420 404
rect 414 399 420 400
rect 582 404 588 405
rect 582 400 583 404
rect 587 400 588 404
rect 582 399 588 400
rect 742 404 748 405
rect 742 400 743 404
rect 747 400 748 404
rect 742 399 748 400
rect 902 404 908 405
rect 902 400 903 404
rect 907 400 908 404
rect 902 399 908 400
rect 1046 404 1052 405
rect 1046 400 1047 404
rect 1051 400 1052 404
rect 1046 399 1052 400
rect 1182 404 1188 405
rect 1182 400 1183 404
rect 1187 400 1188 404
rect 1182 399 1188 400
rect 256 379 258 399
rect 416 379 418 399
rect 584 379 586 399
rect 744 379 746 399
rect 904 379 906 399
rect 1048 379 1050 399
rect 1184 379 1186 399
rect 223 378 227 379
rect 223 373 227 374
rect 255 378 259 379
rect 255 373 259 374
rect 343 378 347 379
rect 343 373 347 374
rect 415 378 419 379
rect 415 373 419 374
rect 471 378 475 379
rect 471 373 475 374
rect 583 378 587 379
rect 583 373 587 374
rect 599 378 603 379
rect 599 373 603 374
rect 719 378 723 379
rect 719 373 723 374
rect 743 378 747 379
rect 743 373 747 374
rect 839 378 843 379
rect 839 373 843 374
rect 903 378 907 379
rect 903 373 907 374
rect 959 378 963 379
rect 959 373 963 374
rect 1047 378 1051 379
rect 1047 373 1051 374
rect 1079 378 1083 379
rect 1079 373 1083 374
rect 1183 378 1187 379
rect 1183 373 1187 374
rect 1207 378 1211 379
rect 1296 376 1298 434
rect 1312 424 1314 441
rect 1382 439 1388 440
rect 1382 435 1383 439
rect 1387 435 1388 439
rect 1382 434 1388 435
rect 1310 423 1316 424
rect 1310 419 1311 423
rect 1315 419 1316 423
rect 1310 418 1316 419
rect 1384 416 1386 434
rect 1440 424 1442 441
rect 1510 439 1516 440
rect 1510 435 1511 439
rect 1515 435 1516 439
rect 1510 434 1516 435
rect 1438 423 1444 424
rect 1438 419 1439 423
rect 1443 419 1444 423
rect 1438 418 1444 419
rect 1512 416 1514 434
rect 1568 424 1570 441
rect 1638 439 1644 440
rect 1638 435 1639 439
rect 1643 435 1644 439
rect 1638 434 1644 435
rect 1566 423 1572 424
rect 1566 419 1567 423
rect 1571 419 1572 423
rect 1566 418 1572 419
rect 1640 416 1642 434
rect 1672 424 1674 441
rect 1742 439 1748 440
rect 1742 435 1743 439
rect 1747 435 1748 439
rect 1742 434 1748 435
rect 1670 423 1676 424
rect 1670 419 1671 423
rect 1675 419 1676 423
rect 1670 418 1676 419
rect 1744 416 1746 434
rect 1768 425 1770 441
rect 1808 425 1810 441
rect 1766 424 1772 425
rect 1766 420 1767 424
rect 1771 420 1772 424
rect 1766 419 1772 420
rect 1806 424 1812 425
rect 1832 424 1834 441
rect 1902 439 1908 440
rect 1902 435 1903 439
rect 1907 435 1908 439
rect 1902 434 1908 435
rect 1806 420 1807 424
rect 1811 420 1812 424
rect 1806 419 1812 420
rect 1830 423 1836 424
rect 1830 419 1831 423
rect 1835 419 1836 423
rect 1830 418 1836 419
rect 1904 416 1906 434
rect 1960 424 1962 441
rect 1958 423 1964 424
rect 1958 419 1959 423
rect 1963 419 1964 423
rect 1958 418 1964 419
rect 2032 416 2034 446
rect 2111 441 2115 442
rect 2127 446 2131 447
rect 2127 441 2131 442
rect 2271 446 2275 447
rect 2271 441 2275 442
rect 2295 446 2299 447
rect 2295 441 2299 442
rect 2112 424 2114 441
rect 2118 439 2124 440
rect 2118 435 2119 439
rect 2123 435 2124 439
rect 2118 434 2124 435
rect 2110 423 2116 424
rect 2110 419 2111 423
rect 2115 419 2116 423
rect 2110 418 2116 419
rect 1382 415 1388 416
rect 1382 411 1383 415
rect 1387 411 1388 415
rect 1382 410 1388 411
rect 1510 415 1516 416
rect 1510 411 1511 415
rect 1515 411 1516 415
rect 1510 410 1516 411
rect 1638 415 1644 416
rect 1638 411 1639 415
rect 1643 411 1644 415
rect 1638 410 1644 411
rect 1742 415 1748 416
rect 1742 411 1743 415
rect 1747 411 1748 415
rect 1742 410 1748 411
rect 1902 415 1908 416
rect 1902 411 1903 415
rect 1907 411 1908 415
rect 1902 410 1908 411
rect 2030 415 2036 416
rect 2030 411 2031 415
rect 2035 411 2036 415
rect 2030 410 2036 411
rect 2074 415 2080 416
rect 2074 411 2075 415
rect 2079 411 2080 415
rect 2074 410 2080 411
rect 1766 407 1772 408
rect 1310 404 1316 405
rect 1310 400 1311 404
rect 1315 400 1316 404
rect 1310 399 1316 400
rect 1438 404 1444 405
rect 1438 400 1439 404
rect 1443 400 1444 404
rect 1438 399 1444 400
rect 1566 404 1572 405
rect 1566 400 1567 404
rect 1571 400 1572 404
rect 1566 399 1572 400
rect 1670 404 1676 405
rect 1670 400 1671 404
rect 1675 400 1676 404
rect 1766 403 1767 407
rect 1771 403 1772 407
rect 1766 402 1772 403
rect 1806 407 1812 408
rect 1806 403 1807 407
rect 1811 403 1812 407
rect 1806 402 1812 403
rect 1830 404 1836 405
rect 1670 399 1676 400
rect 1312 379 1314 399
rect 1440 379 1442 399
rect 1568 379 1570 399
rect 1672 379 1674 399
rect 1768 379 1770 402
rect 1808 379 1810 402
rect 1830 400 1831 404
rect 1835 400 1836 404
rect 1830 399 1836 400
rect 1958 404 1964 405
rect 1958 400 1959 404
rect 1963 400 1964 404
rect 1958 399 1964 400
rect 1832 379 1834 399
rect 1960 379 1962 399
rect 1311 378 1315 379
rect 1207 373 1211 374
rect 1294 375 1300 376
rect 224 357 226 373
rect 344 357 346 373
rect 472 357 474 373
rect 600 357 602 373
rect 720 357 722 373
rect 840 357 842 373
rect 960 357 962 373
rect 1080 357 1082 373
rect 1208 357 1210 373
rect 1294 371 1295 375
rect 1299 371 1300 375
rect 1311 373 1315 374
rect 1439 378 1443 379
rect 1439 373 1443 374
rect 1567 378 1571 379
rect 1567 373 1571 374
rect 1671 378 1675 379
rect 1671 373 1675 374
rect 1767 378 1771 379
rect 1767 373 1771 374
rect 1807 378 1811 379
rect 1807 373 1811 374
rect 1831 378 1835 379
rect 1831 373 1835 374
rect 1927 378 1931 379
rect 1927 373 1931 374
rect 1959 378 1963 379
rect 1959 373 1963 374
rect 2039 378 2043 379
rect 2076 376 2078 410
rect 2110 404 2116 405
rect 2110 400 2111 404
rect 2115 400 2116 404
rect 2110 399 2116 400
rect 2112 379 2114 399
rect 2111 378 2115 379
rect 2039 373 2043 374
rect 2074 375 2080 376
rect 1294 370 1300 371
rect 222 356 228 357
rect 222 352 223 356
rect 227 352 228 356
rect 222 351 228 352
rect 342 356 348 357
rect 342 352 343 356
rect 347 352 348 356
rect 342 351 348 352
rect 470 356 476 357
rect 470 352 471 356
rect 475 352 476 356
rect 470 351 476 352
rect 598 356 604 357
rect 598 352 599 356
rect 603 352 604 356
rect 598 351 604 352
rect 718 356 724 357
rect 718 352 719 356
rect 723 352 724 356
rect 718 351 724 352
rect 838 356 844 357
rect 838 352 839 356
rect 843 352 844 356
rect 838 351 844 352
rect 958 356 964 357
rect 958 352 959 356
rect 963 352 964 356
rect 958 351 964 352
rect 1078 356 1084 357
rect 1078 352 1079 356
rect 1083 352 1084 356
rect 1078 351 1084 352
rect 1206 356 1212 357
rect 1206 352 1207 356
rect 1211 352 1212 356
rect 1768 354 1770 373
rect 1808 354 1810 373
rect 1928 357 1930 373
rect 2040 357 2042 373
rect 2074 371 2075 375
rect 2079 371 2080 375
rect 2111 373 2115 374
rect 2074 370 2080 371
rect 1926 356 1932 357
rect 1206 351 1212 352
rect 1766 353 1772 354
rect 1766 349 1767 353
rect 1771 349 1772 353
rect 1766 348 1772 349
rect 1806 353 1812 354
rect 1806 349 1807 353
rect 1811 349 1812 353
rect 1926 352 1927 356
rect 1931 352 1932 356
rect 1926 351 1932 352
rect 2038 356 2044 357
rect 2038 352 2039 356
rect 2043 352 2044 356
rect 2038 351 2044 352
rect 1806 348 1812 349
rect 2120 348 2122 434
rect 2272 424 2274 441
rect 2360 440 2362 474
rect 2376 452 2378 474
rect 2478 469 2484 470
rect 2478 465 2479 469
rect 2483 465 2484 469
rect 2478 464 2484 465
rect 2374 451 2380 452
rect 2374 447 2375 451
rect 2379 447 2380 451
rect 2480 447 2482 464
rect 2560 452 2562 474
rect 2678 469 2684 470
rect 2678 465 2679 469
rect 2683 465 2684 469
rect 2678 464 2684 465
rect 2558 451 2564 452
rect 2558 447 2559 451
rect 2563 447 2564 451
rect 2680 447 2682 464
rect 2732 452 2734 490
rect 2880 452 2882 550
rect 2982 548 2988 549
rect 2982 544 2983 548
rect 2987 544 2988 548
rect 2982 543 2988 544
rect 3166 548 3172 549
rect 3166 544 3167 548
rect 3171 544 3172 548
rect 3166 543 3172 544
rect 2984 511 2986 543
rect 3168 511 3170 543
rect 2887 510 2891 511
rect 2887 505 2891 506
rect 2983 510 2987 511
rect 2983 505 2987 506
rect 3111 510 3115 511
rect 3111 505 3115 506
rect 3167 510 3171 511
rect 3167 505 3171 506
rect 2888 489 2890 505
rect 3112 489 3114 505
rect 2886 488 2892 489
rect 2886 484 2887 488
rect 2891 484 2892 488
rect 2886 483 2892 484
rect 3110 488 3116 489
rect 3110 484 3111 488
rect 3115 484 3116 488
rect 3110 483 3116 484
rect 3320 480 3322 590
rect 3359 585 3363 586
rect 3367 590 3371 591
rect 3367 585 3371 586
rect 3360 568 3362 585
rect 3432 584 3434 618
rect 3440 596 3442 686
rect 3462 683 3463 687
rect 3467 683 3468 687
rect 3462 682 3468 683
rect 3464 655 3466 682
rect 3463 654 3467 655
rect 3463 649 3467 650
rect 3464 630 3466 649
rect 3462 629 3468 630
rect 3462 625 3463 629
rect 3467 625 3468 629
rect 3462 624 3468 625
rect 3462 612 3468 613
rect 3462 608 3463 612
rect 3467 608 3468 612
rect 3462 607 3468 608
rect 3438 595 3444 596
rect 3438 591 3439 595
rect 3443 591 3444 595
rect 3464 591 3466 607
rect 3438 590 3444 591
rect 3463 590 3467 591
rect 3463 585 3467 586
rect 3430 583 3436 584
rect 3430 579 3431 583
rect 3435 579 3436 583
rect 3430 578 3436 579
rect 3464 569 3466 585
rect 3462 568 3468 569
rect 3358 567 3364 568
rect 3358 563 3359 567
rect 3363 563 3364 567
rect 3462 564 3463 568
rect 3467 564 3468 568
rect 3462 563 3468 564
rect 3358 562 3364 563
rect 3430 555 3436 556
rect 3430 551 3431 555
rect 3435 551 3436 555
rect 3430 550 3436 551
rect 3462 551 3468 552
rect 3358 548 3364 549
rect 3358 544 3359 548
rect 3363 544 3364 548
rect 3358 543 3364 544
rect 3360 511 3362 543
rect 3335 510 3339 511
rect 3335 505 3339 506
rect 3359 510 3363 511
rect 3359 505 3363 506
rect 3336 489 3338 505
rect 3334 488 3340 489
rect 3334 484 3335 488
rect 3339 484 3340 488
rect 3334 483 3340 484
rect 2958 479 2964 480
rect 2958 475 2959 479
rect 2963 475 2964 479
rect 2958 474 2964 475
rect 3318 479 3324 480
rect 3318 475 3319 479
rect 3323 475 3324 479
rect 3318 474 3324 475
rect 2886 469 2892 470
rect 2886 465 2887 469
rect 2891 465 2892 469
rect 2886 464 2892 465
rect 2730 451 2736 452
rect 2730 447 2731 451
rect 2735 447 2736 451
rect 2878 451 2884 452
rect 2878 447 2879 451
rect 2883 447 2884 451
rect 2888 447 2890 464
rect 2960 452 2962 474
rect 3110 469 3116 470
rect 3110 465 3111 469
rect 3115 465 3116 469
rect 3110 464 3116 465
rect 3334 469 3340 470
rect 3334 465 3335 469
rect 3339 465 3340 469
rect 3334 464 3340 465
rect 2958 451 2964 452
rect 2958 447 2959 451
rect 2963 447 2964 451
rect 3112 447 3114 464
rect 3336 447 3338 464
rect 3432 452 3434 550
rect 3462 547 3463 551
rect 3467 547 3468 551
rect 3462 546 3468 547
rect 3464 511 3466 546
rect 3463 510 3467 511
rect 3463 505 3467 506
rect 3464 486 3466 505
rect 3462 485 3468 486
rect 3462 481 3463 485
rect 3467 481 3468 485
rect 3462 480 3468 481
rect 3462 468 3468 469
rect 3462 464 3463 468
rect 3467 464 3468 468
rect 3462 463 3468 464
rect 3430 451 3436 452
rect 3430 447 3431 451
rect 3435 447 3436 451
rect 3464 447 3466 463
rect 2374 446 2380 447
rect 2455 446 2459 447
rect 2455 441 2459 442
rect 2479 446 2483 447
rect 2558 446 2564 447
rect 2655 446 2659 447
rect 2479 441 2483 442
rect 2655 441 2659 442
rect 2679 446 2683 447
rect 2730 446 2736 447
rect 2871 446 2875 447
rect 2878 446 2884 447
rect 2887 446 2891 447
rect 2958 446 2964 447
rect 3103 446 3107 447
rect 2679 441 2683 442
rect 2871 441 2875 442
rect 2887 441 2891 442
rect 3103 441 3107 442
rect 3111 446 3115 447
rect 3111 441 3115 442
rect 3335 446 3339 447
rect 3430 446 3436 447
rect 3463 446 3467 447
rect 3335 441 3339 442
rect 3463 441 3467 442
rect 2358 439 2364 440
rect 2358 435 2359 439
rect 2363 435 2364 439
rect 2358 434 2364 435
rect 2402 439 2408 440
rect 2402 435 2403 439
rect 2407 435 2408 439
rect 2402 434 2408 435
rect 2270 423 2276 424
rect 2270 419 2271 423
rect 2275 419 2276 423
rect 2270 418 2276 419
rect 2404 416 2406 434
rect 2456 424 2458 441
rect 2526 439 2532 440
rect 2526 435 2527 439
rect 2531 435 2532 439
rect 2526 434 2532 435
rect 2454 423 2460 424
rect 2454 419 2455 423
rect 2459 419 2460 423
rect 2454 418 2460 419
rect 2528 416 2530 434
rect 2656 424 2658 441
rect 2726 439 2732 440
rect 2726 435 2727 439
rect 2731 435 2732 439
rect 2726 434 2732 435
rect 2654 423 2660 424
rect 2654 419 2655 423
rect 2659 419 2660 423
rect 2654 418 2660 419
rect 2728 416 2730 434
rect 2872 424 2874 441
rect 2942 439 2948 440
rect 2942 435 2943 439
rect 2947 435 2948 439
rect 2942 434 2948 435
rect 2870 423 2876 424
rect 2870 419 2871 423
rect 2875 419 2876 423
rect 2870 418 2876 419
rect 2944 416 2946 434
rect 3104 424 3106 441
rect 3336 424 3338 441
rect 3342 439 3348 440
rect 3342 435 3343 439
rect 3347 435 3348 439
rect 3342 434 3348 435
rect 3102 423 3108 424
rect 3102 419 3103 423
rect 3107 419 3108 423
rect 3102 418 3108 419
rect 3334 423 3340 424
rect 3334 419 3335 423
rect 3339 419 3340 423
rect 3334 418 3340 419
rect 2402 415 2408 416
rect 2402 411 2403 415
rect 2407 411 2408 415
rect 2402 410 2408 411
rect 2526 415 2532 416
rect 2526 411 2527 415
rect 2531 411 2532 415
rect 2526 410 2532 411
rect 2726 415 2732 416
rect 2726 411 2727 415
rect 2731 411 2732 415
rect 2726 410 2732 411
rect 2942 415 2948 416
rect 2942 411 2943 415
rect 2947 411 2948 415
rect 2942 410 2948 411
rect 3018 415 3024 416
rect 3018 411 3019 415
rect 3023 411 3024 415
rect 3018 410 3024 411
rect 2270 404 2276 405
rect 2270 400 2271 404
rect 2275 400 2276 404
rect 2270 399 2276 400
rect 2454 404 2460 405
rect 2454 400 2455 404
rect 2459 400 2460 404
rect 2454 399 2460 400
rect 2654 404 2660 405
rect 2654 400 2655 404
rect 2659 400 2660 404
rect 2654 399 2660 400
rect 2870 404 2876 405
rect 2870 400 2871 404
rect 2875 400 2876 404
rect 2870 399 2876 400
rect 2272 379 2274 399
rect 2456 379 2458 399
rect 2656 379 2658 399
rect 2872 379 2874 399
rect 2159 378 2163 379
rect 2159 373 2163 374
rect 2271 378 2275 379
rect 2271 373 2275 374
rect 2287 378 2291 379
rect 2287 373 2291 374
rect 2423 378 2427 379
rect 2423 373 2427 374
rect 2455 378 2459 379
rect 2455 373 2459 374
rect 2583 378 2587 379
rect 2583 373 2587 374
rect 2655 378 2659 379
rect 2655 373 2659 374
rect 2759 378 2763 379
rect 2759 373 2763 374
rect 2871 378 2875 379
rect 2871 373 2875 374
rect 2951 378 2955 379
rect 2951 373 2955 374
rect 2160 357 2162 373
rect 2288 357 2290 373
rect 2424 357 2426 373
rect 2584 357 2586 373
rect 2730 371 2736 372
rect 2730 367 2731 371
rect 2735 367 2736 371
rect 2730 366 2736 367
rect 2634 363 2640 364
rect 2634 359 2635 363
rect 2639 359 2640 363
rect 2634 358 2640 359
rect 2158 356 2164 357
rect 2158 352 2159 356
rect 2163 352 2164 356
rect 2158 351 2164 352
rect 2286 356 2292 357
rect 2286 352 2287 356
rect 2291 352 2292 356
rect 2286 351 2292 352
rect 2422 356 2428 357
rect 2422 352 2423 356
rect 2427 352 2428 356
rect 2422 351 2428 352
rect 2582 356 2588 357
rect 2582 352 2583 356
rect 2587 352 2588 356
rect 2582 351 2588 352
rect 206 347 212 348
rect 206 343 207 347
rect 211 343 212 347
rect 206 342 212 343
rect 294 347 300 348
rect 294 343 295 347
rect 299 343 300 347
rect 294 342 300 343
rect 414 347 420 348
rect 414 343 415 347
rect 419 343 420 347
rect 414 342 420 343
rect 542 347 548 348
rect 542 343 543 347
rect 547 343 548 347
rect 542 342 548 343
rect 550 347 556 348
rect 550 343 551 347
rect 555 343 556 347
rect 550 342 556 343
rect 822 347 828 348
rect 822 343 823 347
rect 827 343 828 347
rect 822 342 828 343
rect 910 347 916 348
rect 910 343 911 347
rect 915 343 916 347
rect 910 342 916 343
rect 1030 347 1036 348
rect 1030 343 1031 347
rect 1035 343 1036 347
rect 1030 342 1036 343
rect 1150 347 1156 348
rect 1150 343 1151 347
rect 1155 343 1156 347
rect 1150 342 1156 343
rect 1998 347 2004 348
rect 1998 343 1999 347
rect 2003 343 2004 347
rect 1998 342 2004 343
rect 2118 347 2124 348
rect 2118 343 2119 347
rect 2123 343 2124 347
rect 2118 342 2124 343
rect 2126 347 2132 348
rect 2126 343 2127 347
rect 2131 343 2132 347
rect 2126 342 2132 343
rect 2238 347 2244 348
rect 2238 343 2239 347
rect 2243 343 2244 347
rect 2238 342 2244 343
rect 2366 347 2372 348
rect 2366 343 2367 347
rect 2371 343 2372 347
rect 2366 342 2372 343
rect 208 320 210 342
rect 222 337 228 338
rect 222 333 223 337
rect 227 333 228 337
rect 222 332 228 333
rect 198 319 204 320
rect 198 315 199 319
rect 203 315 204 319
rect 198 314 204 315
rect 206 319 212 320
rect 206 315 207 319
rect 211 315 212 319
rect 206 314 212 315
rect 224 311 226 332
rect 296 320 298 342
rect 342 337 348 338
rect 342 333 343 337
rect 347 333 348 337
rect 342 332 348 333
rect 294 319 300 320
rect 294 315 295 319
rect 299 315 300 319
rect 294 314 300 315
rect 344 311 346 332
rect 416 320 418 342
rect 470 337 476 338
rect 470 333 471 337
rect 475 333 476 337
rect 470 332 476 333
rect 414 319 420 320
rect 414 315 415 319
rect 419 315 420 319
rect 414 314 420 315
rect 472 311 474 332
rect 544 320 546 342
rect 542 319 548 320
rect 542 315 543 319
rect 547 315 548 319
rect 542 314 548 315
rect 552 312 554 342
rect 598 337 604 338
rect 598 333 599 337
rect 603 333 604 337
rect 598 332 604 333
rect 718 337 724 338
rect 718 333 719 337
rect 723 333 724 337
rect 718 332 724 333
rect 550 311 556 312
rect 600 311 602 332
rect 720 311 722 332
rect 824 320 826 342
rect 838 337 844 338
rect 838 333 839 337
rect 843 333 844 337
rect 838 332 844 333
rect 822 319 828 320
rect 822 315 823 319
rect 827 315 828 319
rect 822 314 828 315
rect 840 311 842 332
rect 912 320 914 342
rect 958 337 964 338
rect 958 333 959 337
rect 963 333 964 337
rect 958 332 964 333
rect 910 319 916 320
rect 910 315 911 319
rect 915 315 916 319
rect 910 314 916 315
rect 960 311 962 332
rect 1032 320 1034 342
rect 1078 337 1084 338
rect 1078 333 1079 337
rect 1083 333 1084 337
rect 1078 332 1084 333
rect 1030 319 1036 320
rect 1030 315 1031 319
rect 1035 315 1036 319
rect 1030 314 1036 315
rect 1080 311 1082 332
rect 1152 320 1154 342
rect 1206 337 1212 338
rect 1926 337 1932 338
rect 1206 333 1207 337
rect 1211 333 1212 337
rect 1206 332 1212 333
rect 1766 336 1772 337
rect 1766 332 1767 336
rect 1771 332 1772 336
rect 1150 319 1156 320
rect 1150 315 1151 319
rect 1155 315 1156 319
rect 1150 314 1156 315
rect 1208 311 1210 332
rect 1766 331 1772 332
rect 1806 336 1812 337
rect 1806 332 1807 336
rect 1811 332 1812 336
rect 1926 333 1927 337
rect 1931 333 1932 337
rect 1926 332 1932 333
rect 1806 331 1812 332
rect 1768 311 1770 331
rect 1808 315 1810 331
rect 1928 315 1930 332
rect 2000 320 2002 342
rect 2038 337 2044 338
rect 2038 333 2039 337
rect 2043 333 2044 337
rect 2038 332 2044 333
rect 1998 319 2004 320
rect 1998 315 1999 319
rect 2003 315 2004 319
rect 2040 315 2042 332
rect 1807 314 1811 315
rect 111 310 115 311
rect 111 305 115 306
rect 135 310 139 311
rect 135 305 139 306
rect 223 310 227 311
rect 223 305 227 306
rect 263 310 267 311
rect 263 305 267 306
rect 343 310 347 311
rect 343 305 347 306
rect 375 310 379 311
rect 375 305 379 306
rect 471 310 475 311
rect 471 305 475 306
rect 487 310 491 311
rect 550 307 551 311
rect 555 307 556 311
rect 550 306 556 307
rect 599 310 603 311
rect 487 305 491 306
rect 599 305 603 306
rect 711 310 715 311
rect 711 305 715 306
rect 719 310 723 311
rect 719 305 723 306
rect 815 310 819 311
rect 815 305 819 306
rect 839 310 843 311
rect 839 305 843 306
rect 919 310 923 311
rect 919 305 923 306
rect 959 310 963 311
rect 959 305 963 306
rect 1023 310 1027 311
rect 1023 305 1027 306
rect 1079 310 1083 311
rect 1079 305 1083 306
rect 1127 310 1131 311
rect 1127 305 1131 306
rect 1207 310 1211 311
rect 1207 305 1211 306
rect 1239 310 1243 311
rect 1239 305 1243 306
rect 1767 310 1771 311
rect 1807 309 1811 310
rect 1927 314 1931 315
rect 1998 314 2004 315
rect 2039 314 2043 315
rect 1927 309 1931 310
rect 2128 312 2130 342
rect 2158 337 2164 338
rect 2158 333 2159 337
rect 2163 333 2164 337
rect 2158 332 2164 333
rect 2160 315 2162 332
rect 2240 320 2242 342
rect 2286 337 2292 338
rect 2286 333 2287 337
rect 2291 333 2292 337
rect 2286 332 2292 333
rect 2238 319 2244 320
rect 2238 315 2239 319
rect 2243 315 2244 319
rect 2288 315 2290 332
rect 2368 320 2370 342
rect 2422 337 2428 338
rect 2422 333 2423 337
rect 2427 333 2428 337
rect 2422 332 2428 333
rect 2582 337 2588 338
rect 2582 333 2583 337
rect 2587 333 2588 337
rect 2582 332 2588 333
rect 2366 319 2372 320
rect 2366 315 2367 319
rect 2371 315 2372 319
rect 2424 315 2426 332
rect 2470 319 2476 320
rect 2470 315 2471 319
rect 2475 315 2476 319
rect 2584 315 2586 332
rect 2636 320 2638 358
rect 2654 347 2660 348
rect 2654 343 2655 347
rect 2659 343 2660 347
rect 2654 342 2660 343
rect 2656 320 2658 342
rect 2634 319 2640 320
rect 2634 315 2635 319
rect 2639 315 2640 319
rect 2159 314 2163 315
rect 2039 309 2043 310
rect 2126 311 2132 312
rect 1767 305 1771 306
rect 112 289 114 305
rect 110 288 116 289
rect 264 288 266 305
rect 334 303 340 304
rect 334 299 335 303
rect 339 299 340 303
rect 334 298 340 299
rect 110 284 111 288
rect 115 284 116 288
rect 110 283 116 284
rect 262 287 268 288
rect 262 283 263 287
rect 267 283 268 287
rect 262 282 268 283
rect 336 280 338 298
rect 376 288 378 305
rect 446 303 452 304
rect 446 299 447 303
rect 451 299 452 303
rect 446 298 452 299
rect 374 287 380 288
rect 374 283 375 287
rect 379 283 380 287
rect 374 282 380 283
rect 448 280 450 298
rect 488 288 490 305
rect 558 303 564 304
rect 558 299 559 303
rect 563 299 564 303
rect 558 298 564 299
rect 486 287 492 288
rect 486 283 487 287
rect 491 283 492 287
rect 486 282 492 283
rect 560 280 562 298
rect 600 288 602 305
rect 712 288 714 305
rect 774 303 780 304
rect 774 299 775 303
rect 779 299 780 303
rect 774 298 780 299
rect 598 287 604 288
rect 598 283 599 287
rect 603 283 604 287
rect 598 282 604 283
rect 710 287 716 288
rect 710 283 711 287
rect 715 283 716 287
rect 710 282 716 283
rect 334 279 340 280
rect 334 275 335 279
rect 339 275 340 279
rect 334 274 340 275
rect 446 279 452 280
rect 446 275 447 279
rect 451 275 452 279
rect 446 274 452 275
rect 558 279 564 280
rect 558 275 559 279
rect 563 275 564 279
rect 558 274 564 275
rect 586 279 592 280
rect 586 275 587 279
rect 591 275 592 279
rect 586 274 592 275
rect 110 271 116 272
rect 110 267 111 271
rect 115 267 116 271
rect 110 266 116 267
rect 262 268 268 269
rect 112 243 114 266
rect 262 264 263 268
rect 267 264 268 268
rect 262 263 268 264
rect 374 268 380 269
rect 374 264 375 268
rect 379 264 380 268
rect 374 263 380 264
rect 486 268 492 269
rect 486 264 487 268
rect 491 264 492 268
rect 486 263 492 264
rect 264 243 266 263
rect 376 243 378 263
rect 488 243 490 263
rect 111 242 115 243
rect 111 237 115 238
rect 263 242 267 243
rect 263 237 267 238
rect 375 242 379 243
rect 375 237 379 238
rect 447 242 451 243
rect 447 237 451 238
rect 487 242 491 243
rect 487 237 491 238
rect 535 242 539 243
rect 535 237 539 238
rect 112 218 114 237
rect 448 221 450 237
rect 536 221 538 237
rect 446 220 452 221
rect 110 217 116 218
rect 110 213 111 217
rect 115 213 116 217
rect 446 216 447 220
rect 451 216 452 220
rect 446 215 452 216
rect 534 220 540 221
rect 534 216 535 220
rect 539 216 540 220
rect 534 215 540 216
rect 110 212 116 213
rect 314 211 320 212
rect 314 207 315 211
rect 319 207 320 211
rect 314 206 320 207
rect 526 211 532 212
rect 526 207 527 211
rect 531 207 532 211
rect 526 206 532 207
rect 110 200 116 201
rect 110 196 111 200
rect 115 196 116 200
rect 110 195 116 196
rect 112 151 114 195
rect 111 150 115 151
rect 111 145 115 146
rect 263 150 267 151
rect 263 145 267 146
rect 112 129 114 145
rect 110 128 116 129
rect 264 128 266 145
rect 316 144 318 206
rect 446 201 452 202
rect 446 197 447 201
rect 451 197 452 201
rect 446 196 452 197
rect 448 151 450 196
rect 528 184 530 206
rect 534 201 540 202
rect 534 197 535 201
rect 539 197 540 201
rect 534 196 540 197
rect 526 183 532 184
rect 526 179 527 183
rect 531 179 532 183
rect 526 178 532 179
rect 536 151 538 196
rect 588 184 590 274
rect 598 268 604 269
rect 598 264 599 268
rect 603 264 604 268
rect 598 263 604 264
rect 710 268 716 269
rect 710 264 711 268
rect 715 264 716 268
rect 710 263 716 264
rect 600 243 602 263
rect 712 243 714 263
rect 599 242 603 243
rect 599 237 603 238
rect 623 242 627 243
rect 623 237 627 238
rect 711 242 715 243
rect 711 237 715 238
rect 624 221 626 237
rect 712 221 714 237
rect 622 220 628 221
rect 622 216 623 220
rect 627 216 628 220
rect 622 215 628 216
rect 710 220 716 221
rect 710 216 711 220
rect 715 216 716 220
rect 710 215 716 216
rect 776 212 778 298
rect 816 288 818 305
rect 920 288 922 305
rect 982 303 988 304
rect 982 299 983 303
rect 987 299 988 303
rect 982 298 988 299
rect 814 287 820 288
rect 814 283 815 287
rect 819 283 820 287
rect 814 282 820 283
rect 918 287 924 288
rect 918 283 919 287
rect 923 283 924 287
rect 918 282 924 283
rect 782 275 788 276
rect 782 271 783 275
rect 787 271 788 275
rect 782 270 788 271
rect 694 211 700 212
rect 694 207 695 211
rect 699 207 700 211
rect 694 206 700 207
rect 774 211 780 212
rect 774 207 775 211
rect 779 207 780 211
rect 774 206 780 207
rect 622 201 628 202
rect 622 197 623 201
rect 627 197 628 201
rect 622 196 628 197
rect 586 183 592 184
rect 586 179 587 183
rect 591 179 592 183
rect 586 178 592 179
rect 624 151 626 196
rect 696 184 698 206
rect 710 201 716 202
rect 710 197 711 201
rect 715 197 716 201
rect 710 196 716 197
rect 694 183 700 184
rect 694 179 695 183
rect 699 179 700 183
rect 694 178 700 179
rect 712 151 714 196
rect 784 184 786 270
rect 814 268 820 269
rect 814 264 815 268
rect 819 264 820 268
rect 814 263 820 264
rect 918 268 924 269
rect 918 264 919 268
rect 923 264 924 268
rect 918 263 924 264
rect 816 243 818 263
rect 920 243 922 263
rect 807 242 811 243
rect 807 237 811 238
rect 815 242 819 243
rect 815 237 819 238
rect 903 242 907 243
rect 903 237 907 238
rect 919 242 923 243
rect 919 237 923 238
rect 808 221 810 237
rect 904 221 906 237
rect 806 220 812 221
rect 806 216 807 220
rect 811 216 812 220
rect 806 215 812 216
rect 902 220 908 221
rect 902 216 903 220
rect 907 216 908 220
rect 902 215 908 216
rect 984 212 986 298
rect 1024 288 1026 305
rect 1128 288 1130 305
rect 1198 303 1204 304
rect 1198 299 1199 303
rect 1203 299 1204 303
rect 1198 298 1204 299
rect 1022 287 1028 288
rect 1022 283 1023 287
rect 1027 283 1028 287
rect 1022 282 1028 283
rect 1126 287 1132 288
rect 1126 283 1127 287
rect 1131 283 1132 287
rect 1126 282 1132 283
rect 1200 280 1202 298
rect 1240 288 1242 305
rect 1768 289 1770 305
rect 1808 293 1810 309
rect 2126 307 2127 311
rect 2131 307 2132 311
rect 2159 309 2163 310
rect 2223 314 2227 315
rect 2238 314 2244 315
rect 2287 314 2291 315
rect 2223 309 2227 310
rect 2287 309 2291 310
rect 2311 314 2315 315
rect 2366 314 2372 315
rect 2399 314 2403 315
rect 2311 309 2315 310
rect 2399 309 2403 310
rect 2423 314 2427 315
rect 2470 314 2476 315
rect 2487 314 2491 315
rect 2423 309 2427 310
rect 2126 306 2132 307
rect 1806 292 1812 293
rect 2224 292 2226 309
rect 2274 307 2280 308
rect 2274 303 2275 307
rect 2279 303 2280 307
rect 2274 302 2280 303
rect 2294 307 2300 308
rect 2294 303 2295 307
rect 2299 303 2300 307
rect 2294 302 2300 303
rect 1766 288 1772 289
rect 1238 287 1244 288
rect 1238 283 1239 287
rect 1243 283 1244 287
rect 1766 284 1767 288
rect 1771 284 1772 288
rect 1806 288 1807 292
rect 1811 288 1812 292
rect 1806 287 1812 288
rect 2222 291 2228 292
rect 2222 287 2223 291
rect 2227 287 2228 291
rect 2222 286 2228 287
rect 1766 283 1772 284
rect 1238 282 1244 283
rect 1198 279 1204 280
rect 1198 275 1199 279
rect 1203 275 1204 279
rect 1198 274 1204 275
rect 1318 275 1324 276
rect 1318 271 1319 275
rect 1323 271 1324 275
rect 1806 275 1812 276
rect 1318 270 1324 271
rect 1766 271 1772 272
rect 1022 268 1028 269
rect 1022 264 1023 268
rect 1027 264 1028 268
rect 1022 263 1028 264
rect 1126 268 1132 269
rect 1126 264 1127 268
rect 1131 264 1132 268
rect 1126 263 1132 264
rect 1238 268 1244 269
rect 1238 264 1239 268
rect 1243 264 1244 268
rect 1238 263 1244 264
rect 1024 243 1026 263
rect 1128 243 1130 263
rect 1240 243 1242 263
rect 999 242 1003 243
rect 999 237 1003 238
rect 1023 242 1027 243
rect 1023 237 1027 238
rect 1103 242 1107 243
rect 1103 237 1107 238
rect 1127 242 1131 243
rect 1127 237 1131 238
rect 1207 242 1211 243
rect 1207 237 1211 238
rect 1239 242 1243 243
rect 1239 237 1243 238
rect 1311 242 1315 243
rect 1311 237 1315 238
rect 1000 221 1002 237
rect 1104 221 1106 237
rect 1208 221 1210 237
rect 1312 221 1314 237
rect 998 220 1004 221
rect 998 216 999 220
rect 1003 216 1004 220
rect 998 215 1004 216
rect 1102 220 1108 221
rect 1102 216 1103 220
rect 1107 216 1108 220
rect 1102 215 1108 216
rect 1206 220 1212 221
rect 1206 216 1207 220
rect 1211 216 1212 220
rect 1206 215 1212 216
rect 1310 220 1316 221
rect 1310 216 1311 220
rect 1315 216 1316 220
rect 1310 215 1316 216
rect 878 211 884 212
rect 878 207 879 211
rect 883 207 884 211
rect 878 206 884 207
rect 886 211 892 212
rect 886 207 887 211
rect 891 207 892 211
rect 886 206 892 207
rect 982 211 988 212
rect 982 207 983 211
rect 987 207 988 211
rect 982 206 988 207
rect 1286 211 1292 212
rect 1286 207 1287 211
rect 1291 207 1292 211
rect 1286 206 1292 207
rect 806 201 812 202
rect 806 197 807 201
rect 811 197 812 201
rect 806 196 812 197
rect 782 183 788 184
rect 782 179 783 183
rect 787 179 788 183
rect 782 178 788 179
rect 808 151 810 196
rect 880 176 882 206
rect 888 184 890 206
rect 902 201 908 202
rect 902 197 903 201
rect 907 197 908 201
rect 902 196 908 197
rect 998 201 1004 202
rect 998 197 999 201
rect 1003 197 1004 201
rect 998 196 1004 197
rect 1102 201 1108 202
rect 1102 197 1103 201
rect 1107 197 1108 201
rect 1102 196 1108 197
rect 1206 201 1212 202
rect 1206 197 1207 201
rect 1211 197 1212 201
rect 1206 196 1212 197
rect 886 183 892 184
rect 886 179 887 183
rect 891 179 892 183
rect 886 178 892 179
rect 878 175 884 176
rect 878 171 879 175
rect 883 171 884 175
rect 878 170 884 171
rect 904 151 906 196
rect 950 183 956 184
rect 950 179 951 183
rect 955 179 956 183
rect 950 178 956 179
rect 351 150 355 151
rect 351 145 355 146
rect 439 150 443 151
rect 439 145 443 146
rect 447 150 451 151
rect 447 145 451 146
rect 527 150 531 151
rect 527 145 531 146
rect 535 150 539 151
rect 535 145 539 146
rect 615 150 619 151
rect 615 145 619 146
rect 623 150 627 151
rect 623 145 627 146
rect 703 150 707 151
rect 703 145 707 146
rect 711 150 715 151
rect 711 145 715 146
rect 791 150 795 151
rect 791 145 795 146
rect 807 150 811 151
rect 807 145 811 146
rect 879 150 883 151
rect 879 145 883 146
rect 903 150 907 151
rect 903 145 907 146
rect 314 143 320 144
rect 314 139 315 143
rect 319 139 320 143
rect 314 138 320 139
rect 334 143 340 144
rect 334 139 335 143
rect 339 139 340 143
rect 334 138 340 139
rect 110 124 111 128
rect 115 124 116 128
rect 110 123 116 124
rect 262 127 268 128
rect 262 123 263 127
rect 267 123 268 127
rect 262 122 268 123
rect 336 120 338 138
rect 352 128 354 145
rect 422 143 428 144
rect 422 139 423 143
rect 427 139 428 143
rect 422 138 428 139
rect 350 127 356 128
rect 350 123 351 127
rect 355 123 356 127
rect 350 122 356 123
rect 424 120 426 138
rect 440 128 442 145
rect 510 143 516 144
rect 510 139 511 143
rect 515 139 516 143
rect 510 138 516 139
rect 438 127 444 128
rect 438 123 439 127
rect 443 123 444 127
rect 438 122 444 123
rect 512 120 514 138
rect 528 128 530 145
rect 598 143 604 144
rect 598 139 599 143
rect 603 139 604 143
rect 598 138 604 139
rect 526 127 532 128
rect 526 123 527 127
rect 531 123 532 127
rect 526 122 532 123
rect 600 120 602 138
rect 616 128 618 145
rect 686 143 692 144
rect 686 139 687 143
rect 691 139 692 143
rect 686 138 692 139
rect 614 127 620 128
rect 614 123 615 127
rect 619 123 620 127
rect 614 122 620 123
rect 688 120 690 138
rect 704 128 706 145
rect 774 143 780 144
rect 774 139 775 143
rect 779 139 780 143
rect 774 138 780 139
rect 702 127 708 128
rect 702 123 703 127
rect 707 123 708 127
rect 702 122 708 123
rect 776 120 778 138
rect 792 128 794 145
rect 862 143 868 144
rect 862 139 863 143
rect 867 139 868 143
rect 862 138 868 139
rect 790 127 796 128
rect 790 123 791 127
rect 795 123 796 127
rect 790 122 796 123
rect 864 120 866 138
rect 880 128 882 145
rect 878 127 884 128
rect 878 123 879 127
rect 883 123 884 127
rect 878 122 884 123
rect 952 120 954 178
rect 1000 151 1002 196
rect 1104 151 1106 196
rect 1208 151 1210 196
rect 1288 184 1290 206
rect 1310 201 1316 202
rect 1310 197 1311 201
rect 1315 197 1316 201
rect 1310 196 1316 197
rect 1286 183 1292 184
rect 1286 179 1287 183
rect 1291 179 1292 183
rect 1286 178 1292 179
rect 1312 151 1314 196
rect 1320 184 1322 270
rect 1766 267 1767 271
rect 1771 267 1772 271
rect 1806 271 1807 275
rect 1811 271 1812 275
rect 1806 270 1812 271
rect 2222 272 2228 273
rect 1766 266 1772 267
rect 1768 243 1770 266
rect 1808 243 1810 270
rect 2222 268 2223 272
rect 2227 268 2228 272
rect 2222 267 2228 268
rect 2224 243 2226 267
rect 2276 264 2278 302
rect 2296 284 2298 302
rect 2312 292 2314 309
rect 2382 307 2388 308
rect 2382 303 2383 307
rect 2387 303 2388 307
rect 2382 302 2388 303
rect 2310 291 2316 292
rect 2310 287 2311 291
rect 2315 287 2316 291
rect 2310 286 2316 287
rect 2384 284 2386 302
rect 2400 292 2402 309
rect 2398 291 2404 292
rect 2398 287 2399 291
rect 2403 287 2404 291
rect 2398 286 2404 287
rect 2472 284 2474 314
rect 2487 309 2491 310
rect 2575 314 2579 315
rect 2575 309 2579 310
rect 2583 314 2587 315
rect 2634 314 2640 315
rect 2654 319 2660 320
rect 2654 315 2655 319
rect 2659 315 2660 319
rect 2654 314 2660 315
rect 2679 314 2683 315
rect 2583 309 2587 310
rect 2679 309 2683 310
rect 2488 292 2490 309
rect 2566 307 2572 308
rect 2566 303 2567 307
rect 2571 303 2572 307
rect 2566 302 2572 303
rect 2486 291 2492 292
rect 2486 287 2487 291
rect 2491 287 2492 291
rect 2486 286 2492 287
rect 2568 284 2570 302
rect 2576 292 2578 309
rect 2626 307 2632 308
rect 2626 303 2627 307
rect 2631 303 2632 307
rect 2626 302 2632 303
rect 2574 291 2580 292
rect 2574 287 2575 291
rect 2579 287 2580 291
rect 2574 286 2580 287
rect 2294 283 2300 284
rect 2294 279 2295 283
rect 2299 279 2300 283
rect 2294 278 2300 279
rect 2382 283 2388 284
rect 2382 279 2383 283
rect 2387 279 2388 283
rect 2382 278 2388 279
rect 2470 283 2476 284
rect 2470 279 2471 283
rect 2475 279 2476 283
rect 2470 278 2476 279
rect 2478 283 2484 284
rect 2478 279 2479 283
rect 2483 279 2484 283
rect 2478 278 2484 279
rect 2566 283 2572 284
rect 2566 279 2567 283
rect 2571 279 2572 283
rect 2566 278 2572 279
rect 2310 272 2316 273
rect 2310 268 2311 272
rect 2315 268 2316 272
rect 2310 267 2316 268
rect 2398 272 2404 273
rect 2398 268 2399 272
rect 2403 268 2404 272
rect 2398 267 2404 268
rect 2274 263 2280 264
rect 2274 259 2275 263
rect 2279 259 2280 263
rect 2274 258 2280 259
rect 2312 243 2314 267
rect 2400 243 2402 267
rect 2480 264 2482 278
rect 2486 272 2492 273
rect 2486 268 2487 272
rect 2491 268 2492 272
rect 2486 267 2492 268
rect 2574 272 2580 273
rect 2574 268 2575 272
rect 2579 268 2580 272
rect 2574 267 2580 268
rect 2478 263 2484 264
rect 2478 259 2479 263
rect 2483 259 2484 263
rect 2478 258 2484 259
rect 2488 243 2490 267
rect 2576 243 2578 267
rect 1767 242 1771 243
rect 1767 237 1771 238
rect 1807 242 1811 243
rect 1807 237 1811 238
rect 2143 242 2147 243
rect 2143 237 2147 238
rect 2223 242 2227 243
rect 2223 237 2227 238
rect 2263 242 2267 243
rect 2263 237 2267 238
rect 2311 242 2315 243
rect 2311 237 2315 238
rect 2383 242 2387 243
rect 2383 237 2387 238
rect 2399 242 2403 243
rect 2399 237 2403 238
rect 2487 242 2491 243
rect 2487 237 2491 238
rect 2511 242 2515 243
rect 2511 237 2515 238
rect 2575 242 2579 243
rect 2575 237 2579 238
rect 1768 218 1770 237
rect 1808 218 1810 237
rect 2144 221 2146 237
rect 2264 221 2266 237
rect 2384 221 2386 237
rect 2512 221 2514 237
rect 2142 220 2148 221
rect 1766 217 1772 218
rect 1766 213 1767 217
rect 1771 213 1772 217
rect 1766 212 1772 213
rect 1806 217 1812 218
rect 1806 213 1807 217
rect 1811 213 1812 217
rect 2142 216 2143 220
rect 2147 216 2148 220
rect 2142 215 2148 216
rect 2262 220 2268 221
rect 2262 216 2263 220
rect 2267 216 2268 220
rect 2262 215 2268 216
rect 2382 220 2388 221
rect 2382 216 2383 220
rect 2387 216 2388 220
rect 2382 215 2388 216
rect 2510 220 2516 221
rect 2510 216 2511 220
rect 2515 216 2516 220
rect 2510 215 2516 216
rect 1806 212 1812 213
rect 2628 212 2630 302
rect 2680 292 2682 309
rect 2732 308 2734 366
rect 2760 357 2762 373
rect 2952 357 2954 373
rect 3020 364 3022 410
rect 3102 404 3108 405
rect 3102 400 3103 404
rect 3107 400 3108 404
rect 3102 399 3108 400
rect 3334 404 3340 405
rect 3334 400 3335 404
rect 3339 400 3340 404
rect 3334 399 3340 400
rect 3104 379 3106 399
rect 3336 379 3338 399
rect 3103 378 3107 379
rect 3103 373 3107 374
rect 3151 378 3155 379
rect 3151 373 3155 374
rect 3335 378 3339 379
rect 3335 373 3339 374
rect 3030 371 3036 372
rect 3030 367 3031 371
rect 3035 367 3036 371
rect 3030 366 3036 367
rect 3018 363 3024 364
rect 3018 359 3019 363
rect 3023 359 3024 363
rect 3018 358 3024 359
rect 2758 356 2764 357
rect 2758 352 2759 356
rect 2763 352 2764 356
rect 2758 351 2764 352
rect 2950 356 2956 357
rect 2950 352 2951 356
rect 2955 352 2956 356
rect 2950 351 2956 352
rect 3032 348 3034 366
rect 3152 357 3154 373
rect 3150 356 3156 357
rect 3150 352 3151 356
rect 3155 352 3156 356
rect 3150 351 3156 352
rect 2830 347 2836 348
rect 2830 343 2831 347
rect 2835 343 2836 347
rect 2830 342 2836 343
rect 3022 347 3028 348
rect 3022 343 3023 347
rect 3027 343 3028 347
rect 3022 342 3028 343
rect 3030 347 3036 348
rect 3030 343 3031 347
rect 3035 343 3036 347
rect 3030 342 3036 343
rect 2758 337 2764 338
rect 2758 333 2759 337
rect 2763 333 2764 337
rect 2758 332 2764 333
rect 2760 315 2762 332
rect 2832 320 2834 342
rect 2950 337 2956 338
rect 2950 333 2951 337
rect 2955 333 2956 337
rect 2950 332 2956 333
rect 2830 319 2836 320
rect 2830 315 2831 319
rect 2835 315 2836 319
rect 2952 315 2954 332
rect 3024 320 3026 342
rect 3150 337 3156 338
rect 3150 333 3151 337
rect 3155 333 3156 337
rect 3150 332 3156 333
rect 3022 319 3028 320
rect 3022 315 3023 319
rect 3027 315 3028 319
rect 3152 315 3154 332
rect 2759 314 2763 315
rect 2759 309 2763 310
rect 2799 314 2803 315
rect 2830 314 2836 315
rect 2927 314 2931 315
rect 2799 309 2803 310
rect 2927 309 2931 310
rect 2951 314 2955 315
rect 3022 314 3028 315
rect 3071 314 3075 315
rect 2951 309 2955 310
rect 3071 309 3075 310
rect 3151 314 3155 315
rect 3151 309 3155 310
rect 3223 314 3227 315
rect 3223 309 3227 310
rect 2730 307 2736 308
rect 2730 303 2731 307
rect 2735 303 2736 307
rect 2730 302 2736 303
rect 2750 307 2756 308
rect 2750 303 2751 307
rect 2755 303 2756 307
rect 2750 302 2756 303
rect 2678 291 2684 292
rect 2678 287 2679 291
rect 2683 287 2684 291
rect 2678 286 2684 287
rect 2752 284 2754 302
rect 2800 292 2802 309
rect 2870 307 2876 308
rect 2870 303 2871 307
rect 2875 303 2876 307
rect 2870 302 2876 303
rect 2798 291 2804 292
rect 2798 287 2799 291
rect 2803 287 2804 291
rect 2798 286 2804 287
rect 2872 284 2874 302
rect 2928 292 2930 309
rect 2998 307 3004 308
rect 2998 303 2999 307
rect 3003 303 3004 307
rect 2998 302 3004 303
rect 2926 291 2932 292
rect 2926 287 2927 291
rect 2931 287 2932 291
rect 2926 286 2932 287
rect 3000 284 3002 302
rect 3072 292 3074 309
rect 3142 307 3148 308
rect 3142 303 3143 307
rect 3147 303 3148 307
rect 3142 302 3148 303
rect 3070 291 3076 292
rect 3070 287 3071 291
rect 3075 287 3076 291
rect 3070 286 3076 287
rect 3144 284 3146 302
rect 3224 292 3226 309
rect 3222 291 3228 292
rect 3222 287 3223 291
rect 3227 287 3228 291
rect 3222 286 3228 287
rect 2750 283 2756 284
rect 2750 279 2751 283
rect 2755 279 2756 283
rect 2750 278 2756 279
rect 2870 283 2876 284
rect 2870 279 2871 283
rect 2875 279 2876 283
rect 2870 278 2876 279
rect 2998 283 3004 284
rect 2998 279 2999 283
rect 3003 279 3004 283
rect 2998 278 3004 279
rect 3142 283 3148 284
rect 3142 279 3143 283
rect 3147 279 3148 283
rect 3142 278 3148 279
rect 3150 283 3156 284
rect 3150 279 3151 283
rect 3155 279 3156 283
rect 3150 278 3156 279
rect 2678 272 2684 273
rect 2678 268 2679 272
rect 2683 268 2684 272
rect 2678 267 2684 268
rect 2798 272 2804 273
rect 2798 268 2799 272
rect 2803 268 2804 272
rect 2798 267 2804 268
rect 2926 272 2932 273
rect 2926 268 2927 272
rect 2931 268 2932 272
rect 2926 267 2932 268
rect 3070 272 3076 273
rect 3070 268 3071 272
rect 3075 268 3076 272
rect 3070 267 3076 268
rect 2680 243 2682 267
rect 2800 243 2802 267
rect 2928 243 2930 267
rect 3072 243 3074 267
rect 2639 242 2643 243
rect 2639 237 2643 238
rect 2679 242 2683 243
rect 2679 237 2683 238
rect 2767 242 2771 243
rect 2767 237 2771 238
rect 2799 242 2803 243
rect 2799 237 2803 238
rect 2895 242 2899 243
rect 2895 237 2899 238
rect 2927 242 2931 243
rect 2927 237 2931 238
rect 3015 242 3019 243
rect 3015 237 3019 238
rect 3071 242 3075 243
rect 3071 237 3075 238
rect 3135 242 3139 243
rect 3135 237 3139 238
rect 2640 221 2642 237
rect 2768 221 2770 237
rect 2896 221 2898 237
rect 3016 221 3018 237
rect 3136 221 3138 237
rect 2638 220 2644 221
rect 2638 216 2639 220
rect 2643 216 2644 220
rect 2638 215 2644 216
rect 2766 220 2772 221
rect 2766 216 2767 220
rect 2771 216 2772 220
rect 2766 215 2772 216
rect 2894 220 2900 221
rect 2894 216 2895 220
rect 2899 216 2900 220
rect 2894 215 2900 216
rect 3014 220 3020 221
rect 3014 216 3015 220
rect 3019 216 3020 220
rect 3014 215 3020 216
rect 3134 220 3140 221
rect 3134 216 3135 220
rect 3139 216 3140 220
rect 3134 215 3140 216
rect 2214 211 2220 212
rect 2214 207 2215 211
rect 2219 207 2220 211
rect 2214 206 2220 207
rect 2334 211 2340 212
rect 2334 207 2335 211
rect 2339 207 2340 211
rect 2334 206 2340 207
rect 2454 211 2460 212
rect 2454 207 2455 211
rect 2459 207 2460 211
rect 2454 206 2460 207
rect 2582 211 2588 212
rect 2582 207 2583 211
rect 2587 207 2588 211
rect 2582 206 2588 207
rect 2626 211 2632 212
rect 2626 207 2627 211
rect 2631 207 2632 211
rect 2626 206 2632 207
rect 2974 211 2980 212
rect 2974 207 2975 211
rect 2979 207 2980 211
rect 2974 206 2980 207
rect 2142 201 2148 202
rect 1766 200 1772 201
rect 1766 196 1767 200
rect 1771 196 1772 200
rect 1766 195 1772 196
rect 1806 200 1812 201
rect 1806 196 1807 200
rect 1811 196 1812 200
rect 2142 197 2143 201
rect 2147 197 2148 201
rect 2142 196 2148 197
rect 1806 195 1812 196
rect 1318 183 1324 184
rect 1318 179 1319 183
rect 1323 179 1324 183
rect 1318 178 1324 179
rect 1768 151 1770 195
rect 1808 155 1810 195
rect 2144 155 2146 196
rect 2216 184 2218 206
rect 2262 201 2268 202
rect 2262 197 2263 201
rect 2267 197 2268 201
rect 2262 196 2268 197
rect 2214 183 2220 184
rect 2214 179 2215 183
rect 2219 179 2220 183
rect 2214 178 2220 179
rect 2264 155 2266 196
rect 2336 184 2338 206
rect 2382 201 2388 202
rect 2382 197 2383 201
rect 2387 197 2388 201
rect 2382 196 2388 197
rect 2334 183 2340 184
rect 2334 179 2335 183
rect 2339 179 2340 183
rect 2334 178 2340 179
rect 2374 175 2380 176
rect 2374 171 2375 175
rect 2379 171 2380 175
rect 2374 170 2380 171
rect 1807 154 1811 155
rect 967 150 971 151
rect 967 145 971 146
rect 999 150 1003 151
rect 999 145 1003 146
rect 1055 150 1059 151
rect 1055 145 1059 146
rect 1103 150 1107 151
rect 1103 145 1107 146
rect 1143 150 1147 151
rect 1143 145 1147 146
rect 1207 150 1211 151
rect 1207 145 1211 146
rect 1231 150 1235 151
rect 1231 145 1235 146
rect 1311 150 1315 151
rect 1311 145 1315 146
rect 1319 150 1323 151
rect 1319 145 1323 146
rect 1407 150 1411 151
rect 1407 145 1411 146
rect 1495 150 1499 151
rect 1495 145 1499 146
rect 1583 150 1587 151
rect 1583 145 1587 146
rect 1671 150 1675 151
rect 1767 150 1771 151
rect 1671 145 1675 146
rect 1742 147 1748 148
rect 968 128 970 145
rect 1038 143 1044 144
rect 1038 139 1039 143
rect 1043 139 1044 143
rect 1038 138 1044 139
rect 966 127 972 128
rect 966 123 967 127
rect 971 123 972 127
rect 966 122 972 123
rect 1040 120 1042 138
rect 1056 128 1058 145
rect 1126 143 1132 144
rect 1126 139 1127 143
rect 1131 139 1132 143
rect 1126 138 1132 139
rect 1054 127 1060 128
rect 1054 123 1055 127
rect 1059 123 1060 127
rect 1054 122 1060 123
rect 1128 120 1130 138
rect 1144 128 1146 145
rect 1214 143 1220 144
rect 1214 139 1215 143
rect 1219 139 1220 143
rect 1214 138 1220 139
rect 1142 127 1148 128
rect 1142 123 1143 127
rect 1147 123 1148 127
rect 1142 122 1148 123
rect 1216 120 1218 138
rect 1232 128 1234 145
rect 1302 143 1308 144
rect 1302 139 1303 143
rect 1307 139 1308 143
rect 1302 138 1308 139
rect 1230 127 1236 128
rect 1230 123 1231 127
rect 1235 123 1236 127
rect 1230 122 1236 123
rect 1304 120 1306 138
rect 1320 128 1322 145
rect 1390 143 1396 144
rect 1390 139 1391 143
rect 1395 139 1396 143
rect 1390 138 1396 139
rect 1318 127 1324 128
rect 1318 123 1319 127
rect 1323 123 1324 127
rect 1318 122 1324 123
rect 1392 120 1394 138
rect 1408 128 1410 145
rect 1478 143 1484 144
rect 1478 139 1479 143
rect 1483 139 1484 143
rect 1478 138 1484 139
rect 1406 127 1412 128
rect 1406 123 1407 127
rect 1411 123 1412 127
rect 1406 122 1412 123
rect 1480 120 1482 138
rect 1496 128 1498 145
rect 1566 143 1572 144
rect 1566 139 1567 143
rect 1571 139 1572 143
rect 1566 138 1572 139
rect 1494 127 1500 128
rect 1494 123 1495 127
rect 1499 123 1500 127
rect 1494 122 1500 123
rect 1568 120 1570 138
rect 1584 128 1586 145
rect 1654 143 1660 144
rect 1654 139 1655 143
rect 1659 139 1660 143
rect 1654 138 1660 139
rect 1582 127 1588 128
rect 1582 123 1583 127
rect 1587 123 1588 127
rect 1582 122 1588 123
rect 1656 120 1658 138
rect 1672 128 1674 145
rect 1742 143 1743 147
rect 1747 143 1748 147
rect 1807 149 1811 150
rect 1831 154 1835 155
rect 1831 149 1835 150
rect 1919 154 1923 155
rect 1919 149 1923 150
rect 2007 154 2011 155
rect 2007 149 2011 150
rect 2095 154 2099 155
rect 2095 149 2099 150
rect 2143 154 2147 155
rect 2143 149 2147 150
rect 2183 154 2187 155
rect 2183 149 2187 150
rect 2263 154 2267 155
rect 2263 149 2267 150
rect 2295 154 2299 155
rect 2295 149 2299 150
rect 1767 145 1771 146
rect 1742 142 1748 143
rect 1670 127 1676 128
rect 1670 123 1671 127
rect 1675 123 1676 127
rect 1670 122 1676 123
rect 1744 120 1746 142
rect 1768 129 1770 145
rect 1808 133 1810 149
rect 1806 132 1812 133
rect 1832 132 1834 149
rect 1902 147 1908 148
rect 1902 143 1903 147
rect 1907 143 1908 147
rect 1902 142 1908 143
rect 1766 128 1772 129
rect 1766 124 1767 128
rect 1771 124 1772 128
rect 1806 128 1807 132
rect 1811 128 1812 132
rect 1806 127 1812 128
rect 1830 131 1836 132
rect 1830 127 1831 131
rect 1835 127 1836 131
rect 1830 126 1836 127
rect 1904 124 1906 142
rect 1920 132 1922 149
rect 1990 147 1996 148
rect 1990 143 1991 147
rect 1995 143 1996 147
rect 1990 142 1996 143
rect 1918 131 1924 132
rect 1918 127 1919 131
rect 1923 127 1924 131
rect 1918 126 1924 127
rect 1992 124 1994 142
rect 2008 132 2010 149
rect 2078 147 2084 148
rect 2078 143 2079 147
rect 2083 143 2084 147
rect 2078 142 2084 143
rect 2006 131 2012 132
rect 2006 127 2007 131
rect 2011 127 2012 131
rect 2006 126 2012 127
rect 2080 124 2082 142
rect 2096 132 2098 149
rect 2166 147 2172 148
rect 2166 143 2167 147
rect 2171 143 2172 147
rect 2166 142 2172 143
rect 2094 131 2100 132
rect 2094 127 2095 131
rect 2099 127 2100 131
rect 2094 126 2100 127
rect 2168 124 2170 142
rect 2184 132 2186 149
rect 2254 147 2260 148
rect 2254 143 2255 147
rect 2259 143 2260 147
rect 2254 142 2260 143
rect 2182 131 2188 132
rect 2182 127 2183 131
rect 2187 127 2188 131
rect 2182 126 2188 127
rect 2256 124 2258 142
rect 2296 132 2298 149
rect 2366 147 2372 148
rect 2366 143 2367 147
rect 2371 143 2372 147
rect 2366 142 2372 143
rect 2294 131 2300 132
rect 2294 127 2295 131
rect 2299 127 2300 131
rect 2294 126 2300 127
rect 2368 124 2370 142
rect 2376 124 2378 170
rect 2384 155 2386 196
rect 2456 184 2458 206
rect 2510 201 2516 202
rect 2510 197 2511 201
rect 2515 197 2516 201
rect 2510 196 2516 197
rect 2454 183 2460 184
rect 2454 179 2455 183
rect 2459 179 2460 183
rect 2454 178 2460 179
rect 2512 155 2514 196
rect 2584 184 2586 206
rect 2638 201 2644 202
rect 2638 197 2639 201
rect 2643 197 2644 201
rect 2638 196 2644 197
rect 2766 201 2772 202
rect 2766 197 2767 201
rect 2771 197 2772 201
rect 2766 196 2772 197
rect 2894 201 2900 202
rect 2894 197 2895 201
rect 2899 197 2900 201
rect 2894 196 2900 197
rect 2582 183 2588 184
rect 2582 179 2583 183
rect 2587 179 2588 183
rect 2582 178 2588 179
rect 2640 155 2642 196
rect 2768 155 2770 196
rect 2896 155 2898 196
rect 2976 184 2978 206
rect 3014 201 3020 202
rect 3014 197 3015 201
rect 3019 197 3020 201
rect 3014 196 3020 197
rect 3134 201 3140 202
rect 3134 197 3135 201
rect 3139 197 3140 201
rect 3134 196 3140 197
rect 2974 183 2980 184
rect 2974 179 2975 183
rect 2979 179 2980 183
rect 2974 178 2980 179
rect 3016 155 3018 196
rect 3136 155 3138 196
rect 3152 184 3154 278
rect 3222 272 3228 273
rect 3222 268 3223 272
rect 3227 268 3228 272
rect 3222 267 3228 268
rect 3224 243 3226 267
rect 3223 242 3227 243
rect 3223 237 3227 238
rect 3263 242 3267 243
rect 3263 237 3267 238
rect 3264 221 3266 237
rect 3262 220 3268 221
rect 3262 216 3263 220
rect 3267 216 3268 220
rect 3262 215 3268 216
rect 3344 212 3346 434
rect 3464 425 3466 441
rect 3462 424 3468 425
rect 3462 420 3463 424
rect 3467 420 3468 424
rect 3462 419 3468 420
rect 3406 411 3412 412
rect 3406 407 3407 411
rect 3411 407 3412 411
rect 3406 406 3412 407
rect 3462 407 3468 408
rect 3359 378 3363 379
rect 3359 373 3363 374
rect 3360 357 3362 373
rect 3358 356 3364 357
rect 3358 352 3359 356
rect 3363 352 3364 356
rect 3358 351 3364 352
rect 3358 337 3364 338
rect 3358 333 3359 337
rect 3363 333 3364 337
rect 3358 332 3364 333
rect 3360 315 3362 332
rect 3408 320 3410 406
rect 3462 403 3463 407
rect 3467 403 3468 407
rect 3462 402 3468 403
rect 3464 379 3466 402
rect 3463 378 3467 379
rect 3463 373 3467 374
rect 3464 354 3466 373
rect 3462 353 3468 354
rect 3462 349 3463 353
rect 3467 349 3468 353
rect 3462 348 3468 349
rect 3422 347 3428 348
rect 3422 343 3423 347
rect 3427 343 3428 347
rect 3422 342 3428 343
rect 3406 319 3412 320
rect 3406 315 3407 319
rect 3411 315 3412 319
rect 3359 314 3363 315
rect 3359 309 3363 310
rect 3367 314 3371 315
rect 3406 314 3412 315
rect 3367 309 3371 310
rect 3368 292 3370 309
rect 3415 307 3421 308
rect 3415 303 3416 307
rect 3420 306 3421 307
rect 3424 306 3426 342
rect 3462 336 3468 337
rect 3462 332 3463 336
rect 3467 332 3468 336
rect 3462 331 3468 332
rect 3464 315 3466 331
rect 3463 314 3467 315
rect 3463 309 3467 310
rect 3420 304 3426 306
rect 3420 303 3421 304
rect 3415 302 3421 303
rect 3464 293 3466 309
rect 3462 292 3468 293
rect 3366 291 3372 292
rect 3366 287 3367 291
rect 3371 287 3372 291
rect 3462 288 3463 292
rect 3467 288 3468 292
rect 3462 287 3468 288
rect 3366 286 3372 287
rect 3438 279 3444 280
rect 3438 275 3439 279
rect 3443 275 3444 279
rect 3438 274 3444 275
rect 3462 275 3468 276
rect 3366 272 3372 273
rect 3366 268 3367 272
rect 3371 268 3372 272
rect 3366 267 3372 268
rect 3368 243 3370 267
rect 3367 242 3371 243
rect 3367 237 3371 238
rect 3368 221 3370 237
rect 3366 220 3372 221
rect 3366 216 3367 220
rect 3371 216 3372 220
rect 3366 215 3372 216
rect 3206 211 3212 212
rect 3206 207 3207 211
rect 3211 207 3212 211
rect 3206 206 3212 207
rect 3342 211 3348 212
rect 3342 207 3343 211
rect 3347 207 3348 211
rect 3342 206 3348 207
rect 3430 211 3436 212
rect 3430 207 3431 211
rect 3435 207 3436 211
rect 3430 206 3436 207
rect 3208 184 3210 206
rect 3262 201 3268 202
rect 3262 197 3263 201
rect 3267 197 3268 201
rect 3262 196 3268 197
rect 3366 201 3372 202
rect 3366 197 3367 201
rect 3371 197 3372 201
rect 3366 196 3372 197
rect 3150 183 3156 184
rect 3150 179 3151 183
rect 3155 179 3156 183
rect 3150 178 3156 179
rect 3182 183 3188 184
rect 3182 179 3183 183
rect 3187 179 3188 183
rect 3182 178 3188 179
rect 3206 183 3212 184
rect 3206 179 3207 183
rect 3211 179 3212 183
rect 3206 178 3212 179
rect 2383 154 2387 155
rect 2383 149 2387 150
rect 2407 154 2411 155
rect 2407 149 2411 150
rect 2511 154 2515 155
rect 2511 149 2515 150
rect 2615 154 2619 155
rect 2615 149 2619 150
rect 2639 154 2643 155
rect 2639 149 2643 150
rect 2719 154 2723 155
rect 2719 149 2723 150
rect 2767 154 2771 155
rect 2767 149 2771 150
rect 2815 154 2819 155
rect 2815 149 2819 150
rect 2895 154 2899 155
rect 2895 149 2899 150
rect 2911 154 2915 155
rect 2911 149 2915 150
rect 3007 154 3011 155
rect 3007 149 3011 150
rect 3015 154 3019 155
rect 3015 149 3019 150
rect 3103 154 3107 155
rect 3103 149 3107 150
rect 3135 154 3139 155
rect 3135 149 3139 150
rect 2408 132 2410 149
rect 2512 132 2514 149
rect 2582 147 2588 148
rect 2582 143 2583 147
rect 2587 143 2588 147
rect 2582 142 2588 143
rect 2406 131 2412 132
rect 2406 127 2407 131
rect 2411 127 2412 131
rect 2406 126 2412 127
rect 2510 131 2516 132
rect 2510 127 2511 131
rect 2515 127 2516 131
rect 2510 126 2516 127
rect 2584 124 2586 142
rect 2616 132 2618 149
rect 2686 147 2692 148
rect 2686 143 2687 147
rect 2691 143 2692 147
rect 2686 142 2692 143
rect 2614 131 2620 132
rect 2614 127 2615 131
rect 2619 127 2620 131
rect 2614 126 2620 127
rect 2688 124 2690 142
rect 2720 132 2722 149
rect 2790 147 2796 148
rect 2790 143 2791 147
rect 2795 143 2796 147
rect 2790 142 2796 143
rect 2718 131 2724 132
rect 2718 127 2719 131
rect 2723 127 2724 131
rect 2718 126 2724 127
rect 2792 124 2794 142
rect 2816 132 2818 149
rect 2886 147 2892 148
rect 2886 143 2887 147
rect 2891 143 2892 147
rect 2886 142 2892 143
rect 2814 131 2820 132
rect 2814 127 2815 131
rect 2819 127 2820 131
rect 2814 126 2820 127
rect 2888 124 2890 142
rect 2912 132 2914 149
rect 2982 147 2988 148
rect 2982 143 2983 147
rect 2987 143 2988 147
rect 2982 142 2988 143
rect 2910 131 2916 132
rect 2910 127 2911 131
rect 2915 127 2916 131
rect 2910 126 2916 127
rect 2984 124 2986 142
rect 3008 132 3010 149
rect 3078 147 3084 148
rect 3078 143 3079 147
rect 3083 143 3084 147
rect 3078 142 3084 143
rect 3006 131 3012 132
rect 3006 127 3007 131
rect 3011 127 3012 131
rect 3006 126 3012 127
rect 3080 124 3082 142
rect 3104 132 3106 149
rect 3174 147 3180 148
rect 3174 143 3175 147
rect 3179 143 3180 147
rect 3174 142 3180 143
rect 3102 131 3108 132
rect 3102 127 3103 131
rect 3107 127 3108 131
rect 3102 126 3108 127
rect 3176 124 3178 142
rect 3184 124 3186 178
rect 3264 155 3266 196
rect 3368 155 3370 196
rect 3191 154 3195 155
rect 3191 149 3195 150
rect 3263 154 3267 155
rect 3263 149 3267 150
rect 3279 154 3283 155
rect 3279 149 3283 150
rect 3367 154 3371 155
rect 3367 149 3371 150
rect 3192 132 3194 149
rect 3280 132 3282 149
rect 3358 147 3364 148
rect 3358 143 3359 147
rect 3363 143 3364 147
rect 3358 142 3364 143
rect 3190 131 3196 132
rect 3190 127 3191 131
rect 3195 127 3196 131
rect 3190 126 3196 127
rect 3278 131 3284 132
rect 3278 127 3279 131
rect 3283 127 3284 131
rect 3278 126 3284 127
rect 3360 124 3362 142
rect 3368 132 3370 149
rect 3432 148 3434 206
rect 3440 184 3442 274
rect 3462 271 3463 275
rect 3467 271 3468 275
rect 3462 270 3468 271
rect 3464 243 3466 270
rect 3463 242 3467 243
rect 3463 237 3467 238
rect 3464 218 3466 237
rect 3462 217 3468 218
rect 3462 213 3463 217
rect 3467 213 3468 217
rect 3462 212 3468 213
rect 3462 200 3468 201
rect 3462 196 3463 200
rect 3467 196 3468 200
rect 3462 195 3468 196
rect 3438 183 3444 184
rect 3438 179 3439 183
rect 3443 179 3444 183
rect 3438 178 3444 179
rect 3464 155 3466 195
rect 3463 154 3467 155
rect 3463 149 3467 150
rect 3430 147 3436 148
rect 3430 143 3431 147
rect 3435 143 3436 147
rect 3430 142 3436 143
rect 3464 133 3466 149
rect 3462 132 3468 133
rect 3366 131 3372 132
rect 3366 127 3367 131
rect 3371 127 3372 131
rect 3462 128 3463 132
rect 3467 128 3468 132
rect 3462 127 3468 128
rect 3366 126 3372 127
rect 1766 123 1772 124
rect 1902 123 1908 124
rect 334 119 340 120
rect 334 115 335 119
rect 339 115 340 119
rect 334 114 340 115
rect 422 119 428 120
rect 422 115 423 119
rect 427 115 428 119
rect 422 114 428 115
rect 510 119 516 120
rect 510 115 511 119
rect 515 115 516 119
rect 510 114 516 115
rect 598 119 604 120
rect 598 115 599 119
rect 603 115 604 119
rect 598 114 604 115
rect 686 119 692 120
rect 686 115 687 119
rect 691 115 692 119
rect 686 114 692 115
rect 774 119 780 120
rect 774 115 775 119
rect 779 115 780 119
rect 774 114 780 115
rect 862 119 868 120
rect 862 115 863 119
rect 867 115 868 119
rect 862 114 868 115
rect 950 119 956 120
rect 950 115 951 119
rect 955 115 956 119
rect 950 114 956 115
rect 1038 119 1044 120
rect 1038 115 1039 119
rect 1043 115 1044 119
rect 1038 114 1044 115
rect 1126 119 1132 120
rect 1126 115 1127 119
rect 1131 115 1132 119
rect 1126 114 1132 115
rect 1214 119 1220 120
rect 1214 115 1215 119
rect 1219 115 1220 119
rect 1214 114 1220 115
rect 1302 119 1308 120
rect 1302 115 1303 119
rect 1307 115 1308 119
rect 1302 114 1308 115
rect 1390 119 1396 120
rect 1390 115 1391 119
rect 1395 115 1396 119
rect 1390 114 1396 115
rect 1478 119 1484 120
rect 1478 115 1479 119
rect 1483 115 1484 119
rect 1478 114 1484 115
rect 1566 119 1572 120
rect 1566 115 1567 119
rect 1571 115 1572 119
rect 1566 114 1572 115
rect 1654 119 1660 120
rect 1654 115 1655 119
rect 1659 115 1660 119
rect 1654 114 1660 115
rect 1742 119 1748 120
rect 1742 115 1743 119
rect 1747 115 1748 119
rect 1902 119 1903 123
rect 1907 119 1908 123
rect 1902 118 1908 119
rect 1990 123 1996 124
rect 1990 119 1991 123
rect 1995 119 1996 123
rect 1990 118 1996 119
rect 2078 123 2084 124
rect 2078 119 2079 123
rect 2083 119 2084 123
rect 2078 118 2084 119
rect 2166 123 2172 124
rect 2166 119 2167 123
rect 2171 119 2172 123
rect 2166 118 2172 119
rect 2254 123 2260 124
rect 2254 119 2255 123
rect 2259 119 2260 123
rect 2254 118 2260 119
rect 2366 123 2372 124
rect 2366 119 2367 123
rect 2371 119 2372 123
rect 2366 118 2372 119
rect 2374 123 2380 124
rect 2374 119 2375 123
rect 2379 119 2380 123
rect 2374 118 2380 119
rect 2582 123 2588 124
rect 2582 119 2583 123
rect 2587 119 2588 123
rect 2582 118 2588 119
rect 2686 123 2692 124
rect 2686 119 2687 123
rect 2691 119 2692 123
rect 2686 118 2692 119
rect 2790 123 2796 124
rect 2790 119 2791 123
rect 2795 119 2796 123
rect 2790 118 2796 119
rect 2886 123 2892 124
rect 2886 119 2887 123
rect 2891 119 2892 123
rect 2886 118 2892 119
rect 2982 123 2988 124
rect 2982 119 2983 123
rect 2987 119 2988 123
rect 2982 118 2988 119
rect 3078 123 3084 124
rect 3078 119 3079 123
rect 3083 119 3084 123
rect 3078 118 3084 119
rect 3174 123 3180 124
rect 3174 119 3175 123
rect 3179 119 3180 123
rect 3174 118 3180 119
rect 3182 123 3188 124
rect 3182 119 3183 123
rect 3187 119 3188 123
rect 3182 118 3188 119
rect 3358 123 3364 124
rect 3358 119 3359 123
rect 3363 119 3364 123
rect 3358 118 3364 119
rect 1742 114 1748 115
rect 1806 115 1812 116
rect 110 111 116 112
rect 110 107 111 111
rect 115 107 116 111
rect 1766 111 1772 112
rect 110 106 116 107
rect 262 108 268 109
rect 112 87 114 106
rect 262 104 263 108
rect 267 104 268 108
rect 262 103 268 104
rect 350 108 356 109
rect 350 104 351 108
rect 355 104 356 108
rect 350 103 356 104
rect 438 108 444 109
rect 438 104 439 108
rect 443 104 444 108
rect 438 103 444 104
rect 526 108 532 109
rect 526 104 527 108
rect 531 104 532 108
rect 526 103 532 104
rect 614 108 620 109
rect 614 104 615 108
rect 619 104 620 108
rect 614 103 620 104
rect 702 108 708 109
rect 702 104 703 108
rect 707 104 708 108
rect 702 103 708 104
rect 790 108 796 109
rect 790 104 791 108
rect 795 104 796 108
rect 790 103 796 104
rect 878 108 884 109
rect 878 104 879 108
rect 883 104 884 108
rect 878 103 884 104
rect 966 108 972 109
rect 966 104 967 108
rect 971 104 972 108
rect 966 103 972 104
rect 1054 108 1060 109
rect 1054 104 1055 108
rect 1059 104 1060 108
rect 1054 103 1060 104
rect 1142 108 1148 109
rect 1142 104 1143 108
rect 1147 104 1148 108
rect 1142 103 1148 104
rect 1230 108 1236 109
rect 1230 104 1231 108
rect 1235 104 1236 108
rect 1230 103 1236 104
rect 1318 108 1324 109
rect 1318 104 1319 108
rect 1323 104 1324 108
rect 1318 103 1324 104
rect 1406 108 1412 109
rect 1406 104 1407 108
rect 1411 104 1412 108
rect 1406 103 1412 104
rect 1494 108 1500 109
rect 1494 104 1495 108
rect 1499 104 1500 108
rect 1494 103 1500 104
rect 1582 108 1588 109
rect 1582 104 1583 108
rect 1587 104 1588 108
rect 1582 103 1588 104
rect 1670 108 1676 109
rect 1670 104 1671 108
rect 1675 104 1676 108
rect 1766 107 1767 111
rect 1771 107 1772 111
rect 1806 111 1807 115
rect 1811 111 1812 115
rect 3462 115 3468 116
rect 1806 110 1812 111
rect 1830 112 1836 113
rect 1766 106 1772 107
rect 1670 103 1676 104
rect 264 87 266 103
rect 352 87 354 103
rect 440 87 442 103
rect 528 87 530 103
rect 616 87 618 103
rect 704 87 706 103
rect 792 87 794 103
rect 880 87 882 103
rect 968 87 970 103
rect 1056 87 1058 103
rect 1144 87 1146 103
rect 1232 87 1234 103
rect 1320 87 1322 103
rect 1408 87 1410 103
rect 1496 87 1498 103
rect 1584 87 1586 103
rect 1672 87 1674 103
rect 1768 87 1770 106
rect 1808 91 1810 110
rect 1830 108 1831 112
rect 1835 108 1836 112
rect 1830 107 1836 108
rect 1918 112 1924 113
rect 1918 108 1919 112
rect 1923 108 1924 112
rect 1918 107 1924 108
rect 2006 112 2012 113
rect 2006 108 2007 112
rect 2011 108 2012 112
rect 2006 107 2012 108
rect 2094 112 2100 113
rect 2094 108 2095 112
rect 2099 108 2100 112
rect 2094 107 2100 108
rect 2182 112 2188 113
rect 2182 108 2183 112
rect 2187 108 2188 112
rect 2182 107 2188 108
rect 2294 112 2300 113
rect 2294 108 2295 112
rect 2299 108 2300 112
rect 2294 107 2300 108
rect 2406 112 2412 113
rect 2406 108 2407 112
rect 2411 108 2412 112
rect 2406 107 2412 108
rect 2510 112 2516 113
rect 2510 108 2511 112
rect 2515 108 2516 112
rect 2510 107 2516 108
rect 2614 112 2620 113
rect 2614 108 2615 112
rect 2619 108 2620 112
rect 2614 107 2620 108
rect 2718 112 2724 113
rect 2718 108 2719 112
rect 2723 108 2724 112
rect 2718 107 2724 108
rect 2814 112 2820 113
rect 2814 108 2815 112
rect 2819 108 2820 112
rect 2814 107 2820 108
rect 2910 112 2916 113
rect 2910 108 2911 112
rect 2915 108 2916 112
rect 2910 107 2916 108
rect 3006 112 3012 113
rect 3006 108 3007 112
rect 3011 108 3012 112
rect 3006 107 3012 108
rect 3102 112 3108 113
rect 3102 108 3103 112
rect 3107 108 3108 112
rect 3102 107 3108 108
rect 3190 112 3196 113
rect 3190 108 3191 112
rect 3195 108 3196 112
rect 3190 107 3196 108
rect 3278 112 3284 113
rect 3278 108 3279 112
rect 3283 108 3284 112
rect 3278 107 3284 108
rect 3366 112 3372 113
rect 3366 108 3367 112
rect 3371 108 3372 112
rect 3462 111 3463 115
rect 3467 111 3468 115
rect 3462 110 3468 111
rect 3366 107 3372 108
rect 1832 91 1834 107
rect 1920 91 1922 107
rect 2008 91 2010 107
rect 2096 91 2098 107
rect 2184 91 2186 107
rect 2296 91 2298 107
rect 2408 91 2410 107
rect 2512 91 2514 107
rect 2616 91 2618 107
rect 2720 91 2722 107
rect 2816 91 2818 107
rect 2912 91 2914 107
rect 3008 91 3010 107
rect 3104 91 3106 107
rect 3192 91 3194 107
rect 3280 91 3282 107
rect 3368 91 3370 107
rect 3464 91 3466 110
rect 1807 90 1811 91
rect 111 86 115 87
rect 111 81 115 82
rect 263 86 267 87
rect 263 81 267 82
rect 351 86 355 87
rect 351 81 355 82
rect 439 86 443 87
rect 439 81 443 82
rect 527 86 531 87
rect 527 81 531 82
rect 615 86 619 87
rect 615 81 619 82
rect 703 86 707 87
rect 703 81 707 82
rect 791 86 795 87
rect 791 81 795 82
rect 879 86 883 87
rect 879 81 883 82
rect 967 86 971 87
rect 967 81 971 82
rect 1055 86 1059 87
rect 1055 81 1059 82
rect 1143 86 1147 87
rect 1143 81 1147 82
rect 1231 86 1235 87
rect 1231 81 1235 82
rect 1319 86 1323 87
rect 1319 81 1323 82
rect 1407 86 1411 87
rect 1407 81 1411 82
rect 1495 86 1499 87
rect 1495 81 1499 82
rect 1583 86 1587 87
rect 1583 81 1587 82
rect 1671 86 1675 87
rect 1671 81 1675 82
rect 1767 86 1771 87
rect 1807 85 1811 86
rect 1831 90 1835 91
rect 1831 85 1835 86
rect 1919 90 1923 91
rect 1919 85 1923 86
rect 2007 90 2011 91
rect 2007 85 2011 86
rect 2095 90 2099 91
rect 2095 85 2099 86
rect 2183 90 2187 91
rect 2183 85 2187 86
rect 2295 90 2299 91
rect 2295 85 2299 86
rect 2407 90 2411 91
rect 2407 85 2411 86
rect 2511 90 2515 91
rect 2511 85 2515 86
rect 2615 90 2619 91
rect 2615 85 2619 86
rect 2719 90 2723 91
rect 2719 85 2723 86
rect 2815 90 2819 91
rect 2815 85 2819 86
rect 2911 90 2915 91
rect 2911 85 2915 86
rect 3007 90 3011 91
rect 3007 85 3011 86
rect 3103 90 3107 91
rect 3103 85 3107 86
rect 3191 90 3195 91
rect 3191 85 3195 86
rect 3279 90 3283 91
rect 3279 85 3283 86
rect 3367 90 3371 91
rect 3367 85 3371 86
rect 3463 90 3467 91
rect 3463 85 3467 86
rect 1767 81 1771 82
<< m4c >>
rect 111 3502 115 3506
rect 135 3502 139 3506
rect 271 3502 275 3506
rect 439 3502 443 3506
rect 615 3502 619 3506
rect 791 3502 795 3506
rect 959 3502 963 3506
rect 1119 3502 1123 3506
rect 1263 3502 1267 3506
rect 1407 3502 1411 3506
rect 111 3434 115 3438
rect 135 3434 139 3438
rect 255 3434 259 3438
rect 271 3434 275 3438
rect 415 3434 419 3438
rect 439 3434 443 3438
rect 575 3434 579 3438
rect 615 3434 619 3438
rect 735 3434 739 3438
rect 111 3362 115 3366
rect 135 3362 139 3366
rect 255 3362 259 3366
rect 327 3362 331 3366
rect 415 3362 419 3366
rect 791 3434 795 3438
rect 895 3434 899 3438
rect 959 3434 963 3438
rect 1063 3434 1067 3438
rect 1119 3434 1123 3438
rect 1231 3434 1235 3438
rect 1263 3434 1267 3438
rect 1551 3502 1555 3506
rect 1671 3502 1675 3506
rect 1767 3502 1771 3506
rect 1807 3490 1811 3494
rect 1831 3490 1835 3494
rect 1975 3490 1979 3494
rect 2143 3490 2147 3494
rect 2311 3490 2315 3494
rect 2479 3490 2483 3494
rect 2639 3490 2643 3494
rect 2799 3490 2803 3494
rect 2967 3490 2971 3494
rect 3463 3490 3467 3494
rect 1399 3434 1403 3438
rect 1407 3434 1411 3438
rect 1551 3434 1555 3438
rect 1671 3434 1675 3438
rect 1767 3434 1771 3438
rect 1807 3426 1811 3430
rect 1831 3426 1835 3430
rect 1975 3426 1979 3430
rect 2031 3426 2035 3430
rect 2143 3426 2147 3430
rect 2151 3426 2155 3430
rect 535 3362 539 3366
rect 575 3362 579 3366
rect 735 3362 739 3366
rect 743 3362 747 3366
rect 895 3362 899 3366
rect 935 3362 939 3366
rect 1063 3362 1067 3366
rect 1119 3362 1123 3366
rect 1231 3362 1235 3366
rect 1295 3362 1299 3366
rect 1399 3362 1403 3366
rect 1463 3362 1467 3366
rect 1639 3362 1643 3366
rect 1767 3362 1771 3366
rect 2271 3426 2275 3430
rect 2311 3426 2315 3430
rect 2391 3426 2395 3430
rect 2479 3426 2483 3430
rect 2511 3426 2515 3430
rect 2623 3426 2627 3430
rect 2639 3426 2643 3430
rect 2727 3426 2731 3430
rect 2799 3426 2803 3430
rect 2831 3426 2835 3430
rect 111 3290 115 3294
rect 135 3290 139 3294
rect 279 3290 283 3294
rect 327 3290 331 3294
rect 463 3290 467 3294
rect 535 3290 539 3294
rect 647 3290 651 3294
rect 743 3290 747 3294
rect 831 3290 835 3294
rect 935 3290 939 3294
rect 1007 3290 1011 3294
rect 1119 3290 1123 3294
rect 1175 3290 1179 3294
rect 1295 3290 1299 3294
rect 1343 3290 1347 3294
rect 1463 3290 1467 3294
rect 1503 3290 1507 3294
rect 1639 3290 1643 3294
rect 1671 3290 1675 3294
rect 111 3218 115 3222
rect 135 3218 139 3222
rect 183 3218 187 3222
rect 1807 3358 1811 3362
rect 2031 3358 2035 3362
rect 2151 3358 2155 3362
rect 2159 3358 2163 3362
rect 2271 3358 2275 3362
rect 2295 3358 2299 3362
rect 2391 3358 2395 3362
rect 2431 3358 2435 3362
rect 2511 3358 2515 3362
rect 2567 3358 2571 3362
rect 2623 3358 2627 3362
rect 2703 3358 2707 3362
rect 2727 3358 2731 3362
rect 2935 3426 2939 3430
rect 2967 3426 2971 3430
rect 3039 3426 3043 3430
rect 3151 3426 3155 3430
rect 3463 3426 3467 3430
rect 2831 3358 2835 3362
rect 2839 3358 2843 3362
rect 2935 3358 2939 3362
rect 2975 3358 2979 3362
rect 3039 3358 3043 3362
rect 3119 3358 3123 3362
rect 3151 3358 3155 3362
rect 1767 3290 1771 3294
rect 1807 3294 1811 3298
rect 2087 3294 2091 3298
rect 2159 3294 2163 3298
rect 2239 3294 2243 3298
rect 2295 3294 2299 3298
rect 2399 3294 2403 3298
rect 2431 3294 2435 3298
rect 2559 3294 2563 3298
rect 2567 3294 2571 3298
rect 1807 3226 1811 3230
rect 1911 3226 1915 3230
rect 2047 3226 2051 3230
rect 2087 3226 2091 3230
rect 2199 3226 2203 3230
rect 2239 3226 2243 3230
rect 279 3218 283 3222
rect 327 3218 331 3222
rect 463 3218 467 3222
rect 487 3218 491 3222
rect 647 3218 651 3222
rect 807 3218 811 3222
rect 831 3218 835 3222
rect 967 3218 971 3222
rect 1007 3218 1011 3222
rect 1135 3218 1139 3222
rect 1175 3218 1179 3222
rect 1303 3218 1307 3222
rect 111 3154 115 3158
rect 183 3154 187 3158
rect 327 3154 331 3158
rect 367 3154 371 3158
rect 487 3154 491 3158
rect 607 3154 611 3158
rect 647 3154 651 3158
rect 727 3154 731 3158
rect 807 3154 811 3158
rect 847 3154 851 3158
rect 967 3154 971 3158
rect 1079 3154 1083 3158
rect 1135 3154 1139 3158
rect 1199 3154 1203 3158
rect 1343 3218 1347 3222
rect 1471 3218 1475 3222
rect 1503 3218 1507 3222
rect 1671 3218 1675 3222
rect 1767 3218 1771 3222
rect 2703 3294 2707 3298
rect 2719 3294 2723 3298
rect 3463 3358 3467 3362
rect 2839 3294 2843 3298
rect 2879 3294 2883 3298
rect 2359 3226 2363 3230
rect 2399 3226 2403 3230
rect 2527 3226 2531 3230
rect 2559 3226 2563 3230
rect 2687 3226 2691 3230
rect 2719 3226 2723 3230
rect 2975 3294 2979 3298
rect 3039 3294 3043 3298
rect 3119 3294 3123 3298
rect 3199 3294 3203 3298
rect 3463 3294 3467 3298
rect 2847 3226 2851 3230
rect 2879 3226 2883 3230
rect 3007 3226 3011 3230
rect 3039 3226 3043 3230
rect 3167 3226 3171 3230
rect 3199 3226 3203 3230
rect 1807 3162 1811 3166
rect 1831 3162 1835 3166
rect 1911 3162 1915 3166
rect 2007 3162 2011 3166
rect 2047 3162 2051 3166
rect 2199 3162 2203 3166
rect 2207 3162 2211 3166
rect 1303 3154 1307 3158
rect 1319 3154 1323 3158
rect 1471 3154 1475 3158
rect 1767 3154 1771 3158
rect 111 3086 115 3090
rect 367 3086 371 3090
rect 439 3086 443 3090
rect 487 3086 491 3090
rect 527 3086 531 3090
rect 607 3086 611 3090
rect 615 3086 619 3090
rect 703 3086 707 3090
rect 727 3086 731 3090
rect 791 3086 795 3090
rect 847 3086 851 3090
rect 879 3086 883 3090
rect 967 3086 971 3090
rect 1055 3086 1059 3090
rect 1079 3086 1083 3090
rect 1143 3086 1147 3090
rect 111 3014 115 3018
rect 439 3014 443 3018
rect 503 3014 507 3018
rect 527 3014 531 3018
rect 591 3014 595 3018
rect 615 3014 619 3018
rect 679 3014 683 3018
rect 703 3014 707 3018
rect 767 3014 771 3018
rect 791 3014 795 3018
rect 855 3014 859 3018
rect 111 2938 115 2942
rect 327 2938 331 2942
rect 447 2938 451 2942
rect 503 2938 507 2942
rect 575 2938 579 2942
rect 591 2938 595 2942
rect 679 2938 683 2942
rect 711 2938 715 2942
rect 879 3014 883 3018
rect 1199 3086 1203 3090
rect 1319 3086 1323 3090
rect 1767 3086 1771 3090
rect 1807 3090 1811 3094
rect 1831 3090 1835 3094
rect 2359 3162 2363 3166
rect 2399 3162 2403 3166
rect 2527 3162 2531 3166
rect 2583 3162 2587 3166
rect 2687 3162 2691 3166
rect 2759 3162 2763 3166
rect 3335 3226 3339 3230
rect 3463 3226 3467 3230
rect 2847 3162 2851 3166
rect 2919 3162 2923 3166
rect 3007 3162 3011 3166
rect 3079 3162 3083 3166
rect 3167 3162 3171 3166
rect 3231 3162 3235 3166
rect 3335 3162 3339 3166
rect 3367 3162 3371 3166
rect 3463 3162 3467 3166
rect 1959 3090 1963 3094
rect 2007 3090 2011 3094
rect 2119 3090 2123 3094
rect 2207 3090 2211 3094
rect 2295 3090 2299 3094
rect 2399 3090 2403 3094
rect 2487 3090 2491 3094
rect 2583 3090 2587 3094
rect 2695 3090 2699 3094
rect 2759 3090 2763 3094
rect 2919 3090 2923 3094
rect 3079 3090 3083 3094
rect 3151 3090 3155 3094
rect 3231 3090 3235 3094
rect 3367 3090 3371 3094
rect 943 3014 947 3018
rect 967 3014 971 3018
rect 1031 3014 1035 3018
rect 1055 3014 1059 3018
rect 1119 3014 1123 3018
rect 1143 3014 1147 3018
rect 1207 3014 1211 3018
rect 1295 3014 1299 3018
rect 1767 3014 1771 3018
rect 1807 3010 1811 3014
rect 1831 3010 1835 3014
rect 1919 3010 1923 3014
rect 1959 3010 1963 3014
rect 2031 3010 2035 3014
rect 2119 3010 2123 3014
rect 2143 3010 2147 3014
rect 767 2938 771 2942
rect 847 2938 851 2942
rect 855 2938 859 2942
rect 943 2938 947 2942
rect 975 2938 979 2942
rect 1031 2938 1035 2942
rect 1103 2938 1107 2942
rect 1119 2938 1123 2942
rect 1207 2938 1211 2942
rect 1231 2938 1235 2942
rect 1295 2938 1299 2942
rect 1359 2938 1363 2942
rect 1495 2938 1499 2942
rect 1767 2938 1771 2942
rect 111 2866 115 2870
rect 135 2866 139 2870
rect 255 2866 259 2870
rect 327 2866 331 2870
rect 415 2866 419 2870
rect 447 2866 451 2870
rect 575 2866 579 2870
rect 111 2790 115 2794
rect 135 2790 139 2794
rect 711 2866 715 2870
rect 735 2866 739 2870
rect 847 2866 851 2870
rect 895 2866 899 2870
rect 975 2866 979 2870
rect 1047 2866 1051 2870
rect 1103 2866 1107 2870
rect 1191 2866 1195 2870
rect 1231 2866 1235 2870
rect 1343 2866 1347 2870
rect 1359 2866 1363 2870
rect 1495 2866 1499 2870
rect 1807 2934 1811 2938
rect 1831 2934 1835 2938
rect 2247 3010 2251 3014
rect 2295 3010 2299 3014
rect 2359 3010 2363 3014
rect 2479 3010 2483 3014
rect 2487 3010 2491 3014
rect 3463 3090 3467 3094
rect 2623 3010 2627 3014
rect 2695 3010 2699 3014
rect 2791 3010 2795 3014
rect 2919 3010 2923 3014
rect 2983 3010 2987 3014
rect 3151 3010 3155 3014
rect 3183 3010 3187 3014
rect 3367 3010 3371 3014
rect 1919 2934 1923 2938
rect 2015 2934 2019 2938
rect 2031 2934 2035 2938
rect 2143 2934 2147 2938
rect 3463 3010 3467 3014
rect 2215 2934 2219 2938
rect 2247 2934 2251 2938
rect 2359 2934 2363 2938
rect 2407 2934 2411 2938
rect 2479 2934 2483 2938
rect 2591 2934 2595 2938
rect 2623 2934 2627 2938
rect 2759 2934 2763 2938
rect 2791 2934 2795 2938
rect 2911 2934 2915 2938
rect 2983 2934 2987 2938
rect 3063 2934 3067 2938
rect 3183 2934 3187 2938
rect 3207 2934 3211 2938
rect 3359 2934 3363 2938
rect 3367 2934 3371 2938
rect 1767 2866 1771 2870
rect 1807 2870 1811 2874
rect 1831 2870 1835 2874
rect 1999 2870 2003 2874
rect 2015 2870 2019 2874
rect 247 2790 251 2794
rect 255 2790 259 2794
rect 391 2790 395 2794
rect 415 2790 419 2794
rect 543 2790 547 2794
rect 575 2790 579 2794
rect 695 2790 699 2794
rect 735 2790 739 2794
rect 855 2790 859 2794
rect 895 2790 899 2794
rect 1023 2790 1027 2794
rect 1047 2790 1051 2794
rect 1191 2790 1195 2794
rect 111 2718 115 2722
rect 135 2718 139 2722
rect 247 2718 251 2722
rect 359 2718 363 2722
rect 391 2718 395 2722
rect 479 2718 483 2722
rect 543 2718 547 2722
rect 615 2718 619 2722
rect 695 2718 699 2722
rect 759 2718 763 2722
rect 855 2718 859 2722
rect 1807 2802 1811 2806
rect 1831 2802 1835 2806
rect 1343 2790 1347 2794
rect 1359 2790 1363 2794
rect 1495 2790 1499 2794
rect 1527 2790 1531 2794
rect 1671 2790 1675 2794
rect 1767 2790 1771 2794
rect 2191 2870 2195 2874
rect 2215 2870 2219 2874
rect 2383 2870 2387 2874
rect 2407 2870 2411 2874
rect 2567 2870 2571 2874
rect 2591 2870 2595 2874
rect 2735 2870 2739 2874
rect 2759 2870 2763 2874
rect 1999 2802 2003 2806
rect 2015 2802 2019 2806
rect 2903 2870 2907 2874
rect 2911 2870 2915 2874
rect 3063 2870 3067 2874
rect 3207 2870 3211 2874
rect 3223 2870 3227 2874
rect 3359 2870 3363 2874
rect 3367 2870 3371 2874
rect 2191 2802 2195 2806
rect 2215 2802 2219 2806
rect 2383 2802 2387 2806
rect 2407 2802 2411 2806
rect 2567 2802 2571 2806
rect 2583 2802 2587 2806
rect 2735 2802 2739 2806
rect 2751 2802 2755 2806
rect 2903 2802 2907 2806
rect 2911 2802 2915 2806
rect 3063 2802 3067 2806
rect 911 2718 915 2722
rect 1023 2718 1027 2722
rect 1063 2718 1067 2722
rect 1191 2718 1195 2722
rect 1215 2718 1219 2722
rect 1359 2718 1363 2722
rect 1375 2718 1379 2722
rect 1527 2718 1531 2722
rect 1535 2718 1539 2722
rect 111 2646 115 2650
rect 247 2646 251 2650
rect 359 2646 363 2650
rect 463 2646 467 2650
rect 479 2646 483 2650
rect 551 2646 555 2650
rect 615 2646 619 2650
rect 639 2646 643 2650
rect 743 2646 747 2650
rect 759 2646 763 2650
rect 855 2646 859 2650
rect 911 2646 915 2650
rect 983 2646 987 2650
rect 1063 2646 1067 2650
rect 1127 2646 1131 2650
rect 1215 2646 1219 2650
rect 1279 2646 1283 2650
rect 1375 2646 1379 2650
rect 1439 2646 1443 2650
rect 111 2574 115 2578
rect 463 2574 467 2578
rect 503 2574 507 2578
rect 551 2574 555 2578
rect 591 2574 595 2578
rect 639 2574 643 2578
rect 679 2574 683 2578
rect 743 2574 747 2578
rect 775 2574 779 2578
rect 855 2574 859 2578
rect 879 2574 883 2578
rect 983 2574 987 2578
rect 991 2574 995 2578
rect 1103 2574 1107 2578
rect 1127 2574 1131 2578
rect 1223 2574 1227 2578
rect 1279 2574 1283 2578
rect 1671 2718 1675 2722
rect 1767 2718 1771 2722
rect 1807 2722 1811 2726
rect 1831 2722 1835 2726
rect 2015 2722 2019 2726
rect 2039 2722 2043 2726
rect 2159 2722 2163 2726
rect 2215 2722 2219 2726
rect 2279 2722 2283 2726
rect 2407 2722 2411 2726
rect 3071 2802 3075 2806
rect 3223 2802 3227 2806
rect 3231 2802 3235 2806
rect 2543 2722 2547 2726
rect 2583 2722 2587 2726
rect 2687 2722 2691 2726
rect 2751 2722 2755 2726
rect 2847 2722 2851 2726
rect 2911 2722 2915 2726
rect 1535 2646 1539 2650
rect 1607 2646 1611 2650
rect 1671 2646 1675 2650
rect 1767 2646 1771 2650
rect 1807 2646 1811 2650
rect 1871 2646 1875 2650
rect 1967 2646 1971 2650
rect 2039 2646 2043 2650
rect 2071 2646 2075 2650
rect 2159 2646 2163 2650
rect 2183 2646 2187 2650
rect 1351 2574 1355 2578
rect 1439 2574 1443 2578
rect 1479 2574 1483 2578
rect 1607 2574 1611 2578
rect 111 2502 115 2506
rect 503 2502 507 2506
rect 551 2502 555 2506
rect 591 2502 595 2506
rect 679 2502 683 2506
rect 735 2502 739 2506
rect 775 2502 779 2506
rect 879 2502 883 2506
rect 911 2502 915 2506
rect 991 2502 995 2506
rect 1079 2502 1083 2506
rect 1103 2502 1107 2506
rect 1223 2502 1227 2506
rect 1239 2502 1243 2506
rect 1351 2502 1355 2506
rect 1399 2502 1403 2506
rect 111 2438 115 2442
rect 415 2438 419 2442
rect 503 2438 507 2442
rect 551 2438 555 2442
rect 599 2438 603 2442
rect 111 2370 115 2374
rect 319 2370 323 2374
rect 415 2370 419 2374
rect 431 2370 435 2374
rect 503 2370 507 2374
rect 543 2370 547 2374
rect 703 2438 707 2442
rect 735 2438 739 2442
rect 807 2438 811 2442
rect 911 2438 915 2442
rect 919 2438 923 2442
rect 1767 2574 1771 2578
rect 1807 2570 1811 2574
rect 1831 2570 1835 2574
rect 1871 2570 1875 2574
rect 2279 2646 2283 2650
rect 2295 2646 2299 2650
rect 2407 2646 2411 2650
rect 2431 2646 2435 2650
rect 2543 2646 2547 2650
rect 2583 2646 2587 2650
rect 2687 2646 2691 2650
rect 2759 2646 2763 2650
rect 3023 2722 3027 2726
rect 3071 2722 3075 2726
rect 3207 2722 3211 2726
rect 3231 2722 3235 2726
rect 2847 2646 2851 2650
rect 2959 2646 2963 2650
rect 3023 2646 3027 2650
rect 3167 2646 3171 2650
rect 3207 2646 3211 2650
rect 1919 2570 1923 2574
rect 1967 2570 1971 2574
rect 2007 2570 2011 2574
rect 2071 2570 2075 2574
rect 2111 2570 2115 2574
rect 2183 2570 2187 2574
rect 2223 2570 2227 2574
rect 2295 2570 2299 2574
rect 2343 2570 2347 2574
rect 1479 2502 1483 2506
rect 1567 2502 1571 2506
rect 1607 2502 1611 2506
rect 1767 2502 1771 2506
rect 1807 2506 1811 2510
rect 1831 2506 1835 2510
rect 1919 2506 1923 2510
rect 1951 2506 1955 2510
rect 2007 2506 2011 2510
rect 2039 2506 2043 2510
rect 2111 2506 2115 2510
rect 2431 2570 2435 2574
rect 2487 2570 2491 2574
rect 2583 2570 2587 2574
rect 2647 2570 2651 2574
rect 2759 2570 2763 2574
rect 2815 2570 2819 2574
rect 2959 2570 2963 2574
rect 2999 2570 3003 2574
rect 3167 2570 3171 2574
rect 3191 2570 3195 2574
rect 2135 2506 2139 2510
rect 2015 2499 2019 2500
rect 2015 2496 2019 2499
rect 2223 2506 2227 2510
rect 2239 2506 2243 2510
rect 2343 2506 2347 2510
rect 2367 2506 2371 2510
rect 2487 2506 2491 2510
rect 2527 2506 2531 2510
rect 2215 2496 2219 2500
rect 1039 2438 1043 2442
rect 1079 2438 1083 2442
rect 1167 2438 1171 2442
rect 1239 2438 1243 2442
rect 1295 2438 1299 2442
rect 1399 2438 1403 2442
rect 1423 2438 1427 2442
rect 1567 2438 1571 2442
rect 1767 2438 1771 2442
rect 1807 2434 1811 2438
rect 1951 2434 1955 2438
rect 2039 2434 2043 2438
rect 2135 2434 2139 2438
rect 2215 2434 2219 2438
rect 2239 2434 2243 2438
rect 2303 2434 2307 2438
rect 2367 2434 2371 2438
rect 599 2370 603 2374
rect 655 2370 659 2374
rect 703 2370 707 2374
rect 767 2370 771 2374
rect 807 2370 811 2374
rect 879 2370 883 2374
rect 919 2370 923 2374
rect 991 2370 995 2374
rect 1039 2370 1043 2374
rect 111 2298 115 2302
rect 151 2298 155 2302
rect 271 2298 275 2302
rect 319 2298 323 2302
rect 391 2298 395 2302
rect 111 2230 115 2234
rect 135 2230 139 2234
rect 151 2230 155 2234
rect 247 2230 251 2234
rect 271 2230 275 2234
rect 431 2298 435 2302
rect 519 2298 523 2302
rect 543 2298 547 2302
rect 647 2298 651 2302
rect 655 2298 659 2302
rect 767 2298 771 2302
rect 775 2298 779 2302
rect 1103 2370 1107 2374
rect 1167 2370 1171 2374
rect 1215 2370 1219 2374
rect 1295 2370 1299 2374
rect 1335 2370 1339 2374
rect 3367 2802 3371 2806
rect 3463 2934 3467 2938
rect 3463 2870 3467 2874
rect 3463 2802 3467 2806
rect 3367 2722 3371 2726
rect 3367 2646 3371 2650
rect 3463 2722 3467 2726
rect 3463 2646 3467 2650
rect 3367 2570 3371 2574
rect 2647 2506 2651 2510
rect 2711 2506 2715 2510
rect 2815 2506 2819 2510
rect 2919 2506 2923 2510
rect 2999 2506 3003 2510
rect 3143 2506 3147 2510
rect 3191 2506 3195 2510
rect 3367 2506 3371 2510
rect 3463 2570 3467 2574
rect 3463 2506 3467 2510
rect 2391 2434 2395 2438
rect 2479 2434 2483 2438
rect 2527 2434 2531 2438
rect 2567 2434 2571 2438
rect 2655 2434 2659 2438
rect 2711 2434 2715 2438
rect 2743 2434 2747 2438
rect 2839 2434 2843 2438
rect 2919 2434 2923 2438
rect 2935 2434 2939 2438
rect 1423 2370 1427 2374
rect 1767 2370 1771 2374
rect 1807 2370 1811 2374
rect 2167 2370 2171 2374
rect 2215 2370 2219 2374
rect 2263 2370 2267 2374
rect 2303 2370 2307 2374
rect 2367 2370 2371 2374
rect 2391 2370 2395 2374
rect 2471 2370 2475 2374
rect 2479 2370 2483 2374
rect 879 2298 883 2302
rect 895 2298 899 2302
rect 991 2298 995 2302
rect 1015 2298 1019 2302
rect 391 2230 395 2234
rect 407 2230 411 2234
rect 519 2230 523 2234
rect 583 2230 587 2234
rect 647 2230 651 2234
rect 767 2230 771 2234
rect 775 2230 779 2234
rect 895 2230 899 2234
rect 1103 2298 1107 2302
rect 1143 2298 1147 2302
rect 1215 2298 1219 2302
rect 1271 2298 1275 2302
rect 1335 2298 1339 2302
rect 1767 2298 1771 2302
rect 1807 2298 1811 2302
rect 1887 2298 1891 2302
rect 2039 2298 2043 2302
rect 2167 2298 2171 2302
rect 2199 2298 2203 2302
rect 2567 2370 2571 2374
rect 2575 2370 2579 2374
rect 2655 2370 2659 2374
rect 2687 2370 2691 2374
rect 2743 2370 2747 2374
rect 3143 2434 3147 2438
rect 3367 2434 3371 2438
rect 3463 2434 3467 2438
rect 2799 2370 2803 2374
rect 2839 2370 2843 2374
rect 2911 2370 2915 2374
rect 2935 2370 2939 2374
rect 3023 2370 3027 2374
rect 3463 2370 3467 2374
rect 2263 2298 2267 2302
rect 2367 2298 2371 2302
rect 2375 2298 2379 2302
rect 2471 2298 2475 2302
rect 2551 2298 2555 2302
rect 2575 2298 2579 2302
rect 2687 2298 2691 2302
rect 2719 2298 2723 2302
rect 2799 2298 2803 2302
rect 2887 2298 2891 2302
rect 2911 2298 2915 2302
rect 951 2230 955 2234
rect 1015 2230 1019 2234
rect 1135 2230 1139 2234
rect 1143 2230 1147 2234
rect 1271 2230 1275 2234
rect 1319 2230 1323 2234
rect 1503 2230 1507 2234
rect 1671 2230 1675 2234
rect 111 2158 115 2162
rect 135 2158 139 2162
rect 247 2158 251 2162
rect 391 2158 395 2162
rect 407 2158 411 2162
rect 543 2158 547 2162
rect 583 2158 587 2162
rect 695 2158 699 2162
rect 767 2158 771 2162
rect 839 2158 843 2162
rect 951 2158 955 2162
rect 975 2158 979 2162
rect 1103 2158 1107 2162
rect 1135 2158 1139 2162
rect 1231 2158 1235 2162
rect 1767 2230 1771 2234
rect 1807 2234 1811 2238
rect 1831 2234 1835 2238
rect 1887 2234 1891 2238
rect 1967 2234 1971 2238
rect 2039 2234 2043 2238
rect 2135 2234 2139 2238
rect 2199 2234 2203 2238
rect 2311 2234 2315 2238
rect 2375 2234 2379 2238
rect 2487 2234 2491 2238
rect 2551 2234 2555 2238
rect 2655 2234 2659 2238
rect 3023 2298 3027 2302
rect 3055 2298 3059 2302
rect 3223 2298 3227 2302
rect 3367 2298 3371 2302
rect 3463 2298 3467 2302
rect 2719 2234 2723 2238
rect 2815 2234 2819 2238
rect 2887 2234 2891 2238
rect 2959 2234 2963 2238
rect 3055 2234 3059 2238
rect 3103 2234 3107 2238
rect 3223 2234 3227 2238
rect 3247 2234 3251 2238
rect 3367 2234 3371 2238
rect 3463 2234 3467 2238
rect 1807 2170 1811 2174
rect 1831 2170 1835 2174
rect 1967 2170 1971 2174
rect 2135 2170 2139 2174
rect 2311 2170 2315 2174
rect 2487 2170 2491 2174
rect 2655 2170 2659 2174
rect 2815 2170 2819 2174
rect 1319 2158 1323 2162
rect 1351 2158 1355 2162
rect 1463 2158 1467 2162
rect 1503 2158 1507 2162
rect 1575 2158 1579 2162
rect 1671 2158 1675 2162
rect 1767 2158 1771 2162
rect 111 2090 115 2094
rect 135 2090 139 2094
rect 223 2090 227 2094
rect 247 2090 251 2094
rect 343 2090 347 2094
rect 391 2090 395 2094
rect 463 2090 467 2094
rect 543 2090 547 2094
rect 583 2090 587 2094
rect 695 2090 699 2094
rect 703 2090 707 2094
rect 823 2090 827 2094
rect 839 2090 843 2094
rect 935 2090 939 2094
rect 975 2090 979 2094
rect 1047 2090 1051 2094
rect 111 2018 115 2022
rect 135 2018 139 2022
rect 223 2018 227 2022
rect 239 2018 243 2022
rect 343 2018 347 2022
rect 367 2018 371 2022
rect 463 2018 467 2022
rect 503 2018 507 2022
rect 583 2018 587 2022
rect 639 2018 643 2022
rect 703 2018 707 2022
rect 2927 2170 2931 2174
rect 2959 2170 2963 2174
rect 3015 2170 3019 2174
rect 3103 2170 3107 2174
rect 3191 2170 3195 2174
rect 3247 2170 3251 2174
rect 3279 2170 3283 2174
rect 3367 2170 3371 2174
rect 1807 2098 1811 2102
rect 1103 2090 1107 2094
rect 1159 2090 1163 2094
rect 1231 2090 1235 2094
rect 1279 2090 1283 2094
rect 1351 2090 1355 2094
rect 1463 2090 1467 2094
rect 1575 2090 1579 2094
rect 1671 2090 1675 2094
rect 1767 2090 1771 2094
rect 1831 2098 1835 2102
rect 1991 2098 1995 2102
rect 2167 2098 2171 2102
rect 2343 2098 2347 2102
rect 2503 2098 2507 2102
rect 2655 2098 2659 2102
rect 2791 2098 2795 2102
rect 2919 2098 2923 2102
rect 2927 2098 2931 2102
rect 3015 2098 3019 2102
rect 3039 2098 3043 2102
rect 3103 2098 3107 2102
rect 3159 2098 3163 2102
rect 3191 2098 3195 2102
rect 3271 2098 3275 2102
rect 3279 2098 3283 2102
rect 775 2018 779 2022
rect 823 2018 827 2022
rect 911 2018 915 2022
rect 935 2018 939 2022
rect 1047 2018 1051 2022
rect 1159 2018 1163 2022
rect 1183 2018 1187 2022
rect 111 1950 115 1954
rect 135 1950 139 1954
rect 239 1950 243 1954
rect 295 1950 299 1954
rect 367 1950 371 1954
rect 423 1950 427 1954
rect 503 1950 507 1954
rect 559 1950 563 1954
rect 639 1950 643 1954
rect 703 1950 707 1954
rect 775 1950 779 1954
rect 855 1950 859 1954
rect 911 1950 915 1954
rect 111 1886 115 1890
rect 295 1886 299 1890
rect 423 1886 427 1890
rect 431 1886 435 1890
rect 559 1886 563 1890
rect 575 1886 579 1890
rect 703 1886 707 1890
rect 727 1886 731 1890
rect 111 1818 115 1822
rect 431 1818 435 1822
rect 855 1886 859 1890
rect 887 1886 891 1890
rect 1807 2030 1811 2034
rect 1831 2030 1835 2034
rect 1991 2030 1995 2034
rect 2015 2030 2019 2034
rect 2167 2030 2171 2034
rect 2223 2030 2227 2034
rect 2343 2030 2347 2034
rect 1279 2018 1283 2022
rect 1327 2018 1331 2022
rect 1767 2018 1771 2022
rect 2431 2030 2435 2034
rect 2503 2030 2507 2034
rect 1007 1950 1011 1954
rect 1047 1950 1051 1954
rect 1159 1950 1163 1954
rect 1183 1950 1187 1954
rect 1311 1950 1315 1954
rect 1327 1950 1331 1954
rect 1807 1962 1811 1966
rect 1831 1962 1835 1966
rect 1863 1962 1867 1966
rect 1471 1950 1475 1954
rect 1767 1950 1771 1954
rect 2631 2030 2635 2034
rect 2655 2030 2659 2034
rect 2791 2030 2795 2034
rect 2823 2030 2827 2034
rect 2919 2030 2923 2034
rect 3007 2030 3011 2034
rect 3039 2030 3043 2034
rect 3463 2170 3467 2174
rect 3367 2098 3371 2102
rect 3463 2098 3467 2102
rect 3159 2030 3163 2034
rect 3199 2030 3203 2034
rect 3271 2030 3275 2034
rect 3367 2030 3371 2034
rect 1999 1962 2003 1966
rect 2015 1962 2019 1966
rect 2143 1962 2147 1966
rect 2223 1962 2227 1966
rect 2287 1962 2291 1966
rect 2431 1962 2435 1966
rect 1007 1886 1011 1890
rect 1047 1886 1051 1890
rect 1159 1886 1163 1890
rect 1199 1886 1203 1890
rect 511 1818 515 1822
rect 575 1818 579 1822
rect 631 1818 635 1822
rect 727 1818 731 1822
rect 759 1818 763 1822
rect 887 1818 891 1822
rect 1023 1818 1027 1822
rect 1047 1818 1051 1822
rect 111 1750 115 1754
rect 439 1750 443 1754
rect 511 1750 515 1754
rect 535 1750 539 1754
rect 631 1750 635 1754
rect 639 1750 643 1754
rect 111 1682 115 1686
rect 399 1682 403 1686
rect 439 1682 443 1686
rect 487 1682 491 1686
rect 743 1750 747 1754
rect 759 1750 763 1754
rect 1807 1894 1811 1898
rect 1863 1894 1867 1898
rect 1999 1894 2003 1898
rect 2015 1894 2019 1898
rect 2111 1894 2115 1898
rect 2143 1894 2147 1898
rect 2215 1894 2219 1898
rect 2287 1894 2291 1898
rect 1311 1886 1315 1890
rect 1351 1886 1355 1890
rect 1471 1886 1475 1890
rect 1511 1886 1515 1890
rect 1671 1886 1675 1890
rect 1767 1886 1771 1890
rect 2575 1962 2579 1966
rect 2631 1962 2635 1966
rect 2711 1962 2715 1966
rect 2823 1962 2827 1966
rect 2831 1962 2835 1966
rect 2951 1962 2955 1966
rect 3007 1962 3011 1966
rect 3063 1962 3067 1966
rect 3167 1962 3171 1966
rect 3199 1962 3203 1966
rect 3279 1962 3283 1966
rect 3367 1962 3371 1966
rect 3463 2030 3467 2034
rect 3463 1962 3467 1966
rect 2327 1894 2331 1898
rect 2431 1894 2435 1898
rect 2439 1894 2443 1898
rect 2543 1894 2547 1898
rect 2575 1894 2579 1898
rect 1151 1818 1155 1822
rect 1199 1818 1203 1822
rect 1279 1818 1283 1822
rect 1351 1818 1355 1822
rect 1407 1818 1411 1822
rect 1511 1818 1515 1822
rect 1535 1818 1539 1822
rect 1671 1818 1675 1822
rect 1767 1818 1771 1822
rect 1807 1822 1811 1826
rect 2015 1822 2019 1826
rect 2103 1822 2107 1826
rect 2111 1822 2115 1826
rect 2191 1822 2195 1826
rect 2215 1822 2219 1826
rect 2279 1822 2283 1826
rect 2327 1822 2331 1826
rect 2367 1822 2371 1826
rect 2439 1822 2443 1826
rect 2455 1822 2459 1826
rect 847 1750 851 1754
rect 887 1750 891 1754
rect 951 1750 955 1754
rect 1023 1750 1027 1754
rect 1055 1750 1059 1754
rect 1151 1750 1155 1754
rect 1159 1750 1163 1754
rect 1271 1750 1275 1754
rect 1279 1750 1283 1754
rect 535 1682 539 1686
rect 575 1682 579 1686
rect 639 1682 643 1686
rect 663 1682 667 1686
rect 111 1614 115 1618
rect 279 1614 283 1618
rect 383 1614 387 1618
rect 399 1614 403 1618
rect 487 1614 491 1618
rect 495 1614 499 1618
rect 111 1542 115 1546
rect 183 1542 187 1546
rect 279 1542 283 1546
rect 327 1542 331 1546
rect 383 1542 387 1546
rect 575 1614 579 1618
rect 607 1614 611 1618
rect 663 1614 667 1618
rect 743 1682 747 1686
rect 759 1682 763 1686
rect 847 1682 851 1686
rect 855 1682 859 1686
rect 951 1682 955 1686
rect 1047 1682 1051 1686
rect 1055 1682 1059 1686
rect 1383 1750 1387 1754
rect 1407 1750 1411 1754
rect 1535 1750 1539 1754
rect 1671 1750 1675 1754
rect 1767 1750 1771 1754
rect 1807 1746 1811 1750
rect 2103 1746 2107 1750
rect 2143 1746 2147 1750
rect 2191 1746 2195 1750
rect 2647 1894 2651 1898
rect 2711 1894 2715 1898
rect 2759 1894 2763 1898
rect 2831 1894 2835 1898
rect 2871 1894 2875 1898
rect 2951 1894 2955 1898
rect 2983 1894 2987 1898
rect 3063 1894 3067 1898
rect 3167 1894 3171 1898
rect 3279 1894 3283 1898
rect 3367 1894 3371 1898
rect 3463 1894 3467 1898
rect 2543 1822 2547 1826
rect 2631 1822 2635 1826
rect 2647 1822 2651 1826
rect 2719 1822 2723 1826
rect 2759 1822 2763 1826
rect 2807 1822 2811 1826
rect 2871 1822 2875 1826
rect 2895 1822 2899 1826
rect 2983 1822 2987 1826
rect 3463 1822 3467 1826
rect 2231 1746 2235 1750
rect 2279 1746 2283 1750
rect 2319 1746 2323 1750
rect 2367 1746 2371 1750
rect 2407 1746 2411 1750
rect 2455 1746 2459 1750
rect 2495 1746 2499 1750
rect 2543 1746 2547 1750
rect 2583 1746 2587 1750
rect 2631 1746 2635 1750
rect 2671 1746 2675 1750
rect 1143 1682 1147 1686
rect 1159 1682 1163 1686
rect 1271 1682 1275 1686
rect 1383 1682 1387 1686
rect 1767 1682 1771 1686
rect 1807 1678 1811 1682
rect 2103 1678 2107 1682
rect 2143 1678 2147 1682
rect 2191 1678 2195 1682
rect 2231 1678 2235 1682
rect 2279 1678 2283 1682
rect 2319 1678 2323 1682
rect 2367 1678 2371 1682
rect 2407 1678 2411 1682
rect 2455 1678 2459 1682
rect 719 1614 723 1618
rect 759 1614 763 1618
rect 831 1614 835 1618
rect 471 1542 475 1546
rect 495 1542 499 1546
rect 607 1542 611 1546
rect 623 1542 627 1546
rect 855 1614 859 1618
rect 943 1614 947 1618
rect 951 1614 955 1618
rect 1047 1614 1051 1618
rect 1055 1614 1059 1618
rect 1143 1614 1147 1618
rect 1167 1614 1171 1618
rect 1279 1614 1283 1618
rect 1767 1614 1771 1618
rect 1807 1610 1811 1614
rect 2063 1610 2067 1614
rect 2103 1610 2107 1614
rect 2159 1610 2163 1614
rect 2191 1610 2195 1614
rect 2255 1610 2259 1614
rect 2279 1610 2283 1614
rect 2359 1610 2363 1614
rect 2367 1610 2371 1614
rect 2495 1678 2499 1682
rect 2543 1678 2547 1682
rect 2583 1678 2587 1682
rect 2631 1678 2635 1682
rect 2719 1746 2723 1750
rect 2759 1746 2763 1750
rect 2807 1746 2811 1750
rect 2847 1746 2851 1750
rect 2895 1746 2899 1750
rect 3463 1746 3467 1750
rect 2671 1678 2675 1682
rect 2719 1678 2723 1682
rect 2759 1678 2763 1682
rect 2807 1678 2811 1682
rect 2847 1678 2851 1682
rect 2895 1678 2899 1682
rect 3463 1678 3467 1682
rect 2455 1610 2459 1614
rect 2463 1610 2467 1614
rect 2543 1610 2547 1614
rect 2567 1610 2571 1614
rect 2631 1610 2635 1614
rect 2671 1610 2675 1614
rect 2719 1610 2723 1614
rect 2775 1610 2779 1614
rect 2807 1610 2811 1614
rect 2887 1610 2891 1614
rect 2895 1610 2899 1614
rect 3463 1610 3467 1614
rect 719 1542 723 1546
rect 767 1542 771 1546
rect 831 1542 835 1546
rect 911 1542 915 1546
rect 943 1542 947 1546
rect 1047 1542 1051 1546
rect 1055 1542 1059 1546
rect 1167 1542 1171 1546
rect 1175 1542 1179 1546
rect 1279 1542 1283 1546
rect 1311 1542 1315 1546
rect 1447 1542 1451 1546
rect 1767 1542 1771 1546
rect 1807 1546 1811 1550
rect 1919 1546 1923 1550
rect 2039 1546 2043 1550
rect 2063 1546 2067 1550
rect 111 1474 115 1478
rect 159 1474 163 1478
rect 183 1474 187 1478
rect 327 1474 331 1478
rect 375 1474 379 1478
rect 471 1474 475 1478
rect 583 1474 587 1478
rect 623 1474 627 1478
rect 767 1474 771 1478
rect 783 1474 787 1478
rect 911 1474 915 1478
rect 959 1474 963 1478
rect 1047 1474 1051 1478
rect 1127 1474 1131 1478
rect 1175 1474 1179 1478
rect 1279 1474 1283 1478
rect 1311 1474 1315 1478
rect 111 1406 115 1410
rect 135 1406 139 1410
rect 159 1406 163 1410
rect 303 1406 307 1410
rect 375 1406 379 1410
rect 495 1406 499 1410
rect 583 1406 587 1410
rect 679 1406 683 1410
rect 783 1406 787 1410
rect 855 1406 859 1410
rect 959 1406 963 1410
rect 1015 1406 1019 1410
rect 111 1338 115 1342
rect 135 1338 139 1342
rect 247 1338 251 1342
rect 303 1338 307 1342
rect 399 1338 403 1342
rect 495 1338 499 1342
rect 559 1338 563 1342
rect 679 1338 683 1342
rect 727 1338 731 1342
rect 855 1338 859 1342
rect 895 1338 899 1342
rect 1431 1474 1435 1478
rect 1447 1474 1451 1478
rect 1591 1474 1595 1478
rect 1767 1474 1771 1478
rect 1807 1474 1811 1478
rect 1831 1474 1835 1478
rect 1919 1474 1923 1478
rect 1951 1474 1955 1478
rect 2159 1546 2163 1550
rect 2167 1546 2171 1550
rect 2255 1546 2259 1550
rect 2295 1546 2299 1550
rect 2359 1546 2363 1550
rect 2423 1546 2427 1550
rect 2463 1546 2467 1550
rect 2551 1546 2555 1550
rect 2567 1546 2571 1550
rect 2671 1546 2675 1550
rect 2679 1546 2683 1550
rect 2775 1546 2779 1550
rect 2799 1546 2803 1550
rect 2887 1546 2891 1550
rect 2927 1546 2931 1550
rect 3055 1546 3059 1550
rect 3463 1546 3467 1550
rect 2039 1474 2043 1478
rect 2111 1474 2115 1478
rect 2167 1474 2171 1478
rect 2271 1474 2275 1478
rect 2295 1474 2299 1478
rect 2423 1474 2427 1478
rect 2431 1474 2435 1478
rect 2551 1474 2555 1478
rect 2591 1474 2595 1478
rect 2679 1474 2683 1478
rect 2735 1474 2739 1478
rect 2799 1474 2803 1478
rect 2871 1474 2875 1478
rect 2927 1474 2931 1478
rect 3007 1474 3011 1478
rect 1127 1406 1131 1410
rect 1167 1406 1171 1410
rect 1279 1406 1283 1410
rect 1303 1406 1307 1410
rect 1431 1406 1435 1410
rect 1559 1406 1563 1410
rect 1591 1406 1595 1410
rect 1671 1406 1675 1410
rect 1767 1406 1771 1410
rect 1807 1406 1811 1410
rect 1831 1406 1835 1410
rect 1951 1406 1955 1410
rect 2007 1406 2011 1410
rect 2111 1406 2115 1410
rect 2199 1406 2203 1410
rect 2271 1406 2275 1410
rect 2383 1406 2387 1410
rect 1015 1338 1019 1342
rect 1063 1338 1067 1342
rect 1167 1338 1171 1342
rect 1223 1338 1227 1342
rect 1303 1338 1307 1342
rect 1375 1338 1379 1342
rect 1431 1338 1435 1342
rect 187 1280 191 1284
rect 111 1270 115 1274
rect 135 1270 139 1274
rect 499 1280 503 1284
rect 223 1270 227 1274
rect 247 1270 251 1274
rect 319 1270 323 1274
rect 399 1270 403 1274
rect 431 1270 435 1274
rect 551 1270 555 1274
rect 559 1270 563 1274
rect 679 1270 683 1274
rect 727 1270 731 1274
rect 1535 1338 1539 1342
rect 1559 1338 1563 1342
rect 1671 1338 1675 1342
rect 1767 1338 1771 1342
rect 1807 1334 1811 1338
rect 1831 1334 1835 1338
rect 2431 1406 2435 1410
rect 2559 1406 2563 1410
rect 2591 1406 2595 1410
rect 3055 1474 3059 1478
rect 3135 1474 3139 1478
rect 3263 1474 3267 1478
rect 3367 1474 3371 1478
rect 3463 1474 3467 1478
rect 2719 1406 2723 1410
rect 2735 1406 2739 1410
rect 2863 1406 2867 1410
rect 2871 1406 2875 1410
rect 2999 1406 3003 1410
rect 3007 1406 3011 1410
rect 3127 1406 3131 1410
rect 3135 1406 3139 1410
rect 3255 1406 3259 1410
rect 3263 1406 3267 1410
rect 3367 1406 3371 1410
rect 3463 1406 3467 1410
rect 1967 1334 1971 1338
rect 2007 1334 2011 1338
rect 2143 1334 2147 1338
rect 2199 1334 2203 1338
rect 2327 1334 2331 1338
rect 2383 1334 2387 1338
rect 2511 1334 2515 1338
rect 2559 1334 2563 1338
rect 2687 1334 2691 1338
rect 2719 1334 2723 1338
rect 2863 1334 2867 1338
rect 2999 1334 3003 1338
rect 3039 1334 3043 1338
rect 3127 1334 3131 1338
rect 3215 1334 3219 1338
rect 3255 1334 3259 1338
rect 3367 1334 3371 1338
rect 823 1270 827 1274
rect 895 1270 899 1274
rect 975 1270 979 1274
rect 1063 1270 1067 1274
rect 1143 1270 1147 1274
rect 1223 1270 1227 1274
rect 1319 1270 1323 1274
rect 1375 1270 1379 1274
rect 1503 1270 1507 1274
rect 1535 1270 1539 1274
rect 1671 1270 1675 1274
rect 1767 1270 1771 1274
rect 1807 1270 1811 1274
rect 1831 1270 1835 1274
rect 1967 1270 1971 1274
rect 2095 1270 2099 1274
rect 2143 1270 2147 1274
rect 111 1198 115 1202
rect 135 1198 139 1202
rect 223 1198 227 1202
rect 231 1198 235 1202
rect 319 1198 323 1202
rect 359 1198 363 1202
rect 431 1198 435 1202
rect 487 1198 491 1202
rect 551 1198 555 1202
rect 615 1198 619 1202
rect 679 1198 683 1202
rect 743 1198 747 1202
rect 823 1198 827 1202
rect 871 1198 875 1202
rect 975 1198 979 1202
rect 991 1198 995 1202
rect 1119 1198 1123 1202
rect 1143 1198 1147 1202
rect 1247 1198 1251 1202
rect 1319 1198 1323 1202
rect 2327 1270 2331 1274
rect 2359 1270 2363 1274
rect 2511 1270 2515 1274
rect 2599 1270 2603 1274
rect 2687 1270 2691 1274
rect 2807 1270 2811 1274
rect 2863 1270 2867 1274
rect 3007 1270 3011 1274
rect 3039 1270 3043 1274
rect 3199 1270 3203 1274
rect 3215 1270 3219 1274
rect 1503 1198 1507 1202
rect 1671 1198 1675 1202
rect 1767 1198 1771 1202
rect 1807 1198 1811 1202
rect 1831 1198 1835 1202
rect 1935 1198 1939 1202
rect 2039 1198 2043 1202
rect 2095 1198 2099 1202
rect 2159 1198 2163 1202
rect 2287 1198 2291 1202
rect 2359 1198 2363 1202
rect 2423 1198 2427 1202
rect 2567 1198 2571 1202
rect 2599 1198 2603 1202
rect 111 1130 115 1134
rect 135 1130 139 1134
rect 231 1130 235 1134
rect 247 1130 251 1134
rect 359 1130 363 1134
rect 367 1130 371 1134
rect 487 1130 491 1134
rect 495 1130 499 1134
rect 615 1130 619 1134
rect 623 1130 627 1134
rect 743 1130 747 1134
rect 759 1130 763 1134
rect 871 1130 875 1134
rect 887 1130 891 1134
rect 991 1130 995 1134
rect 1015 1130 1019 1134
rect 1119 1130 1123 1134
rect 1143 1130 1147 1134
rect 1247 1130 1251 1134
rect 1271 1130 1275 1134
rect 1399 1130 1403 1134
rect 1767 1130 1771 1134
rect 111 1062 115 1066
rect 247 1062 251 1066
rect 367 1062 371 1066
rect 431 1062 435 1066
rect 495 1062 499 1066
rect 543 1062 547 1066
rect 623 1062 627 1066
rect 663 1062 667 1066
rect 759 1062 763 1066
rect 791 1062 795 1066
rect 887 1062 891 1066
rect 919 1062 923 1066
rect 1015 1062 1019 1066
rect 1039 1062 1043 1066
rect 1143 1062 1147 1066
rect 1159 1062 1163 1066
rect 1271 1062 1275 1066
rect 1279 1062 1283 1066
rect 1807 1126 1811 1130
rect 1935 1126 1939 1130
rect 1943 1126 1947 1130
rect 2039 1126 2043 1130
rect 2063 1126 2067 1130
rect 2159 1126 2163 1130
rect 2191 1126 2195 1130
rect 2287 1126 2291 1130
rect 2319 1126 2323 1130
rect 2423 1126 2427 1130
rect 2455 1126 2459 1130
rect 1399 1062 1403 1066
rect 1407 1062 1411 1066
rect 1535 1062 1539 1066
rect 1767 1062 1771 1066
rect 1807 1058 1811 1062
rect 1847 1058 1851 1062
rect 1943 1058 1947 1062
rect 1983 1058 1987 1062
rect 2063 1058 2067 1062
rect 2119 1058 2123 1062
rect 111 990 115 994
rect 431 990 435 994
rect 543 990 547 994
rect 567 990 571 994
rect 663 990 667 994
rect 679 990 683 994
rect 791 990 795 994
rect 911 990 915 994
rect 919 990 923 994
rect 1031 990 1035 994
rect 1039 990 1043 994
rect 1143 990 1147 994
rect 1159 990 1163 994
rect 1255 990 1259 994
rect 1279 990 1283 994
rect 1359 990 1363 994
rect 1407 990 1411 994
rect 2191 1058 2195 1062
rect 2255 1058 2259 1062
rect 2319 1058 2323 1062
rect 2703 1198 2707 1202
rect 2807 1198 2811 1202
rect 2839 1198 2843 1202
rect 2975 1198 2979 1202
rect 3007 1198 3011 1202
rect 3367 1270 3371 1274
rect 3463 1334 3467 1338
rect 3463 1270 3467 1274
rect 3111 1198 3115 1202
rect 3199 1198 3203 1202
rect 3247 1198 3251 1202
rect 3367 1198 3371 1202
rect 2567 1126 2571 1130
rect 2599 1126 2603 1130
rect 2703 1126 2707 1130
rect 2751 1126 2755 1130
rect 2839 1126 2843 1130
rect 2903 1126 2907 1130
rect 2975 1126 2979 1130
rect 3063 1126 3067 1130
rect 3111 1126 3115 1130
rect 3223 1126 3227 1130
rect 3247 1126 3251 1130
rect 2391 1058 2395 1062
rect 2455 1058 2459 1062
rect 2543 1058 2547 1062
rect 2599 1058 2603 1062
rect 2703 1058 2707 1062
rect 2751 1058 2755 1062
rect 1471 990 1475 994
rect 1535 990 1539 994
rect 1583 990 1587 994
rect 1671 990 1675 994
rect 1767 990 1771 994
rect 1807 990 1811 994
rect 1831 990 1835 994
rect 1847 990 1851 994
rect 1975 990 1979 994
rect 1983 990 1987 994
rect 2119 990 2123 994
rect 2135 990 2139 994
rect 2255 990 2259 994
rect 2295 990 2299 994
rect 111 922 115 926
rect 415 922 419 926
rect 559 922 563 926
rect 567 922 571 926
rect 679 922 683 926
rect 727 922 731 926
rect 791 922 795 926
rect 911 922 915 926
rect 111 854 115 858
rect 135 854 139 858
rect 231 854 235 858
rect 359 854 363 858
rect 415 854 419 858
rect 487 854 491 858
rect 559 854 563 858
rect 623 854 627 858
rect 1031 922 1035 926
rect 1119 922 1123 926
rect 1143 922 1147 926
rect 1255 922 1259 926
rect 1335 922 1339 926
rect 1359 922 1363 926
rect 1471 922 1475 926
rect 2391 990 2395 994
rect 2463 990 2467 994
rect 2543 990 2547 994
rect 2631 990 2635 994
rect 2703 990 2707 994
rect 1559 922 1563 926
rect 1583 922 1587 926
rect 727 854 731 858
rect 751 854 755 858
rect 879 854 883 858
rect 911 854 915 858
rect 1007 854 1011 858
rect 1119 854 1123 858
rect 1135 854 1139 858
rect 1271 854 1275 858
rect 111 786 115 790
rect 135 786 139 790
rect 223 786 227 790
rect 231 786 235 790
rect 343 786 347 790
rect 359 786 363 790
rect 471 786 475 790
rect 487 786 491 790
rect 607 786 611 790
rect 623 786 627 790
rect 743 786 747 790
rect 751 786 755 790
rect 1671 922 1675 926
rect 1767 922 1771 926
rect 1807 926 1811 930
rect 1831 926 1835 930
rect 1975 926 1979 930
rect 2127 926 2131 930
rect 2135 926 2139 930
rect 2215 926 2219 930
rect 2295 926 2299 930
rect 2303 926 2307 930
rect 2391 926 2395 930
rect 2463 926 2467 930
rect 2863 1058 2867 1062
rect 2903 1058 2907 1062
rect 3031 1058 3035 1062
rect 3063 1058 3067 1062
rect 3207 1058 3211 1062
rect 3223 1058 3227 1062
rect 3367 1126 3371 1130
rect 3463 1198 3467 1202
rect 3463 1126 3467 1130
rect 3367 1058 3371 1062
rect 2807 990 2811 994
rect 2863 990 2867 994
rect 2991 990 2995 994
rect 3031 990 3035 994
rect 3183 990 3187 994
rect 3207 990 3211 994
rect 3367 990 3371 994
rect 2479 926 2483 930
rect 2567 926 2571 930
rect 2631 926 2635 930
rect 2655 926 2659 930
rect 2743 926 2747 930
rect 2807 926 2811 930
rect 2831 926 2835 930
rect 2991 926 2995 930
rect 3183 926 3187 930
rect 1335 854 1339 858
rect 1559 854 1563 858
rect 1767 854 1771 858
rect 1807 854 1811 858
rect 2127 854 2131 858
rect 2159 854 2163 858
rect 2215 854 2219 858
rect 2247 854 2251 858
rect 2303 854 2307 858
rect 2335 854 2339 858
rect 2391 854 2395 858
rect 2423 854 2427 858
rect 2479 854 2483 858
rect 879 786 883 790
rect 887 786 891 790
rect 1007 786 1011 790
rect 1039 786 1043 790
rect 1135 786 1139 790
rect 1191 786 1195 790
rect 111 718 115 722
rect 135 718 139 722
rect 167 718 171 722
rect 223 718 227 722
rect 295 718 299 722
rect 343 718 347 722
rect 431 718 435 722
rect 471 718 475 722
rect 575 718 579 722
rect 607 718 611 722
rect 727 718 731 722
rect 743 718 747 722
rect 879 718 883 722
rect 887 718 891 722
rect 1031 718 1035 722
rect 1039 718 1043 722
rect 111 650 115 654
rect 167 650 171 654
rect 295 650 299 654
rect 431 650 435 654
rect 455 650 459 654
rect 559 650 563 654
rect 575 650 579 654
rect 679 650 683 654
rect 727 650 731 654
rect 799 650 803 654
rect 879 650 883 654
rect 927 650 931 654
rect 1271 786 1275 790
rect 1351 786 1355 790
rect 1767 786 1771 790
rect 1807 786 1811 790
rect 2063 786 2067 790
rect 2159 786 2163 790
rect 2175 786 2179 790
rect 2527 854 2531 858
rect 2567 854 2571 858
rect 2639 854 2643 858
rect 2655 854 2659 858
rect 2743 854 2747 858
rect 2767 854 2771 858
rect 2831 854 2835 858
rect 2911 854 2915 858
rect 3063 854 3067 858
rect 3223 854 3227 858
rect 2247 786 2251 790
rect 2295 786 2299 790
rect 2335 786 2339 790
rect 2423 786 2427 790
rect 2527 786 2531 790
rect 2559 786 2563 790
rect 2639 786 2643 790
rect 2711 786 2715 790
rect 2767 786 2771 790
rect 2871 786 2875 790
rect 2911 786 2915 790
rect 1183 718 1187 722
rect 1191 718 1195 722
rect 1343 718 1347 722
rect 1351 718 1355 722
rect 1503 718 1507 722
rect 1767 718 1771 722
rect 1807 722 1811 726
rect 1927 722 1931 726
rect 2063 722 2067 726
rect 3039 786 3043 790
rect 3063 786 3067 790
rect 2071 722 2075 726
rect 1031 650 1035 654
rect 1055 650 1059 654
rect 1183 650 1187 654
rect 111 578 115 582
rect 455 578 459 582
rect 559 578 563 582
rect 599 578 603 582
rect 679 578 683 582
rect 703 578 707 582
rect 799 578 803 582
rect 815 578 819 582
rect 927 578 931 582
rect 2175 722 2179 726
rect 2231 722 2235 726
rect 2295 722 2299 726
rect 2391 722 2395 726
rect 2423 722 2427 726
rect 2551 722 2555 726
rect 2559 722 2563 726
rect 2703 722 2707 726
rect 2711 722 2715 726
rect 2847 722 2851 726
rect 2871 722 2875 726
rect 2983 722 2987 726
rect 3039 722 3043 726
rect 3119 722 3123 726
rect 3463 1058 3467 1062
rect 3463 990 3467 994
rect 3367 926 3371 930
rect 3367 854 3371 858
rect 3463 926 3467 930
rect 3463 854 3467 858
rect 3215 786 3219 790
rect 3223 786 3227 790
rect 3367 786 3371 790
rect 3215 722 3219 726
rect 3255 722 3259 726
rect 3367 722 3371 726
rect 1311 650 1315 654
rect 1343 650 1347 654
rect 1447 650 1451 654
rect 1503 650 1507 654
rect 1583 650 1587 654
rect 1767 650 1771 654
rect 1807 650 1811 654
rect 1831 650 1835 654
rect 1927 650 1931 654
rect 1967 650 1971 654
rect 2071 650 2075 654
rect 2135 650 2139 654
rect 2231 650 2235 654
rect 2311 650 2315 654
rect 2391 650 2395 654
rect 1039 578 1043 582
rect 1055 578 1059 582
rect 1151 578 1155 582
rect 1183 578 1187 582
rect 1255 578 1259 582
rect 1311 578 1315 582
rect 1359 578 1363 582
rect 1447 578 1451 582
rect 1471 578 1475 582
rect 1583 578 1587 582
rect 111 514 115 518
rect 303 514 307 518
rect 431 514 435 518
rect 567 514 571 518
rect 599 514 603 518
rect 703 514 707 518
rect 815 514 819 518
rect 847 514 851 518
rect 111 442 115 446
rect 135 442 139 446
rect 255 442 259 446
rect 303 442 307 446
rect 415 442 419 446
rect 431 442 435 446
rect 567 442 571 446
rect 583 442 587 446
rect 927 514 931 518
rect 983 514 987 518
rect 1039 514 1043 518
rect 1111 514 1115 518
rect 1151 514 1155 518
rect 1807 586 1811 590
rect 1831 586 1835 590
rect 1967 586 1971 590
rect 2127 586 2131 590
rect 2135 586 2139 590
rect 1671 578 1675 582
rect 1767 578 1771 582
rect 1231 514 1235 518
rect 1255 514 1259 518
rect 1351 514 1355 518
rect 1359 514 1363 518
rect 1463 514 1467 518
rect 1471 514 1475 518
rect 1575 514 1579 518
rect 1583 514 1587 518
rect 1671 514 1675 518
rect 2487 650 2491 654
rect 2551 650 2555 654
rect 2655 650 2659 654
rect 2287 586 2291 590
rect 2311 586 2315 590
rect 2455 586 2459 590
rect 2487 586 2491 590
rect 2703 650 2707 654
rect 2815 650 2819 654
rect 2847 650 2851 654
rect 2959 650 2963 654
rect 2983 650 2987 654
rect 3103 650 3107 654
rect 3119 650 3123 654
rect 3247 650 3251 654
rect 3255 650 3259 654
rect 2623 586 2627 590
rect 2655 586 2659 590
rect 2799 586 2803 590
rect 2815 586 2819 590
rect 3463 786 3467 790
rect 3463 722 3467 726
rect 3367 650 3371 654
rect 2959 586 2963 590
rect 2983 586 2987 590
rect 3103 586 3107 590
rect 3167 586 3171 590
rect 3247 586 3251 590
rect 1767 514 1771 518
rect 1807 506 1811 510
rect 1831 506 1835 510
rect 1967 506 1971 510
rect 2127 506 2131 510
rect 2287 506 2291 510
rect 2295 506 2299 510
rect 2455 506 2459 510
rect 2479 506 2483 510
rect 2623 506 2627 510
rect 2679 506 2683 510
rect 2799 506 2803 510
rect 703 442 707 446
rect 743 442 747 446
rect 847 442 851 446
rect 903 442 907 446
rect 983 442 987 446
rect 1047 442 1051 446
rect 1111 442 1115 446
rect 1183 442 1187 446
rect 1231 442 1235 446
rect 1311 442 1315 446
rect 1351 442 1355 446
rect 1439 442 1443 446
rect 1463 442 1467 446
rect 1567 442 1571 446
rect 1575 442 1579 446
rect 1671 442 1675 446
rect 1767 442 1771 446
rect 1807 442 1811 446
rect 1831 442 1835 446
rect 1959 442 1963 446
rect 1967 442 1971 446
rect 111 374 115 378
rect 135 374 139 378
rect 223 374 227 378
rect 255 374 259 378
rect 343 374 347 378
rect 415 374 419 378
rect 471 374 475 378
rect 583 374 587 378
rect 599 374 603 378
rect 719 374 723 378
rect 743 374 747 378
rect 839 374 843 378
rect 903 374 907 378
rect 959 374 963 378
rect 1047 374 1051 378
rect 1079 374 1083 378
rect 1183 374 1187 378
rect 1207 374 1211 378
rect 2111 442 2115 446
rect 2127 442 2131 446
rect 2271 442 2275 446
rect 2295 442 2299 446
rect 1311 374 1315 378
rect 1439 374 1443 378
rect 1567 374 1571 378
rect 1671 374 1675 378
rect 1767 374 1771 378
rect 1807 374 1811 378
rect 1831 374 1835 378
rect 1927 374 1931 378
rect 1959 374 1963 378
rect 2039 374 2043 378
rect 2111 374 2115 378
rect 2887 506 2891 510
rect 2983 506 2987 510
rect 3111 506 3115 510
rect 3167 506 3171 510
rect 3359 586 3363 590
rect 3367 586 3371 590
rect 3463 650 3467 654
rect 3463 586 3467 590
rect 3335 506 3339 510
rect 3359 506 3363 510
rect 3463 506 3467 510
rect 2455 442 2459 446
rect 2479 442 2483 446
rect 2655 442 2659 446
rect 2679 442 2683 446
rect 2871 442 2875 446
rect 2887 442 2891 446
rect 3103 442 3107 446
rect 3111 442 3115 446
rect 3335 442 3339 446
rect 3463 442 3467 446
rect 2159 374 2163 378
rect 2271 374 2275 378
rect 2287 374 2291 378
rect 2423 374 2427 378
rect 2455 374 2459 378
rect 2583 374 2587 378
rect 2655 374 2659 378
rect 2759 374 2763 378
rect 2871 374 2875 378
rect 2951 374 2955 378
rect 111 306 115 310
rect 135 306 139 310
rect 223 306 227 310
rect 263 306 267 310
rect 343 306 347 310
rect 375 306 379 310
rect 471 306 475 310
rect 487 306 491 310
rect 599 306 603 310
rect 711 306 715 310
rect 719 306 723 310
rect 815 306 819 310
rect 839 306 843 310
rect 919 306 923 310
rect 959 306 963 310
rect 1023 306 1027 310
rect 1079 306 1083 310
rect 1127 306 1131 310
rect 1207 306 1211 310
rect 1239 306 1243 310
rect 1767 306 1771 310
rect 1807 310 1811 314
rect 1927 310 1931 314
rect 2039 310 2043 314
rect 111 238 115 242
rect 263 238 267 242
rect 375 238 379 242
rect 447 238 451 242
rect 487 238 491 242
rect 535 238 539 242
rect 111 146 115 150
rect 263 146 267 150
rect 599 238 603 242
rect 623 238 627 242
rect 711 238 715 242
rect 807 238 811 242
rect 815 238 819 242
rect 903 238 907 242
rect 919 238 923 242
rect 2159 310 2163 314
rect 2223 310 2227 314
rect 2287 310 2291 314
rect 2311 310 2315 314
rect 2399 310 2403 314
rect 2423 310 2427 314
rect 999 238 1003 242
rect 1023 238 1027 242
rect 1103 238 1107 242
rect 1127 238 1131 242
rect 1207 238 1211 242
rect 1239 238 1243 242
rect 1311 238 1315 242
rect 351 146 355 150
rect 439 146 443 150
rect 447 146 451 150
rect 527 146 531 150
rect 535 146 539 150
rect 615 146 619 150
rect 623 146 627 150
rect 703 146 707 150
rect 711 146 715 150
rect 791 146 795 150
rect 807 146 811 150
rect 879 146 883 150
rect 903 146 907 150
rect 2487 310 2491 314
rect 2575 310 2579 314
rect 2583 310 2587 314
rect 2679 310 2683 314
rect 1767 238 1771 242
rect 1807 238 1811 242
rect 2143 238 2147 242
rect 2223 238 2227 242
rect 2263 238 2267 242
rect 2311 238 2315 242
rect 2383 238 2387 242
rect 2399 238 2403 242
rect 2487 238 2491 242
rect 2511 238 2515 242
rect 2575 238 2579 242
rect 3103 374 3107 378
rect 3151 374 3155 378
rect 3335 374 3339 378
rect 2759 310 2763 314
rect 2799 310 2803 314
rect 2927 310 2931 314
rect 2951 310 2955 314
rect 3071 310 3075 314
rect 3151 310 3155 314
rect 3223 310 3227 314
rect 2639 238 2643 242
rect 2679 238 2683 242
rect 2767 238 2771 242
rect 2799 238 2803 242
rect 2895 238 2899 242
rect 2927 238 2931 242
rect 3015 238 3019 242
rect 3071 238 3075 242
rect 3135 238 3139 242
rect 967 146 971 150
rect 999 146 1003 150
rect 1055 146 1059 150
rect 1103 146 1107 150
rect 1143 146 1147 150
rect 1207 146 1211 150
rect 1231 146 1235 150
rect 1311 146 1315 150
rect 1319 146 1323 150
rect 1407 146 1411 150
rect 1495 146 1499 150
rect 1583 146 1587 150
rect 1671 146 1675 150
rect 1767 146 1771 150
rect 1807 150 1811 154
rect 1831 150 1835 154
rect 1919 150 1923 154
rect 2007 150 2011 154
rect 2095 150 2099 154
rect 2143 150 2147 154
rect 2183 150 2187 154
rect 2263 150 2267 154
rect 2295 150 2299 154
rect 3223 238 3227 242
rect 3263 238 3267 242
rect 3359 374 3363 378
rect 3463 374 3467 378
rect 3359 310 3363 314
rect 3367 310 3371 314
rect 3463 310 3467 314
rect 3367 238 3371 242
rect 2383 150 2387 154
rect 2407 150 2411 154
rect 2511 150 2515 154
rect 2615 150 2619 154
rect 2639 150 2643 154
rect 2719 150 2723 154
rect 2767 150 2771 154
rect 2815 150 2819 154
rect 2895 150 2899 154
rect 2911 150 2915 154
rect 3007 150 3011 154
rect 3015 150 3019 154
rect 3103 150 3107 154
rect 3135 150 3139 154
rect 3191 150 3195 154
rect 3263 150 3267 154
rect 3279 150 3283 154
rect 3367 150 3371 154
rect 3463 238 3467 242
rect 3463 150 3467 154
rect 111 82 115 86
rect 263 82 267 86
rect 351 82 355 86
rect 439 82 443 86
rect 527 82 531 86
rect 615 82 619 86
rect 703 82 707 86
rect 791 82 795 86
rect 879 82 883 86
rect 967 82 971 86
rect 1055 82 1059 86
rect 1143 82 1147 86
rect 1231 82 1235 86
rect 1319 82 1323 86
rect 1407 82 1411 86
rect 1495 82 1499 86
rect 1583 82 1587 86
rect 1671 82 1675 86
rect 1767 82 1771 86
rect 1807 86 1811 90
rect 1831 86 1835 90
rect 1919 86 1923 90
rect 2007 86 2011 90
rect 2095 86 2099 90
rect 2183 86 2187 90
rect 2295 86 2299 90
rect 2407 86 2411 90
rect 2511 86 2515 90
rect 2615 86 2619 90
rect 2719 86 2723 90
rect 2815 86 2819 90
rect 2911 86 2915 90
rect 3007 86 3011 90
rect 3103 86 3107 90
rect 3191 86 3195 90
rect 3279 86 3283 90
rect 3367 86 3371 90
rect 3463 86 3467 90
<< m4 >>
rect 96 3501 97 3507
rect 103 3506 1791 3507
rect 103 3502 111 3506
rect 115 3502 135 3506
rect 139 3502 271 3506
rect 275 3502 439 3506
rect 443 3502 615 3506
rect 619 3502 791 3506
rect 795 3502 959 3506
rect 963 3502 1119 3506
rect 1123 3502 1263 3506
rect 1267 3502 1407 3506
rect 1411 3502 1551 3506
rect 1555 3502 1671 3506
rect 1675 3502 1767 3506
rect 1771 3502 1791 3506
rect 103 3501 1791 3502
rect 1797 3501 1798 3507
rect 1790 3489 1791 3495
rect 1797 3494 3499 3495
rect 1797 3490 1807 3494
rect 1811 3490 1831 3494
rect 1835 3490 1975 3494
rect 1979 3490 2143 3494
rect 2147 3490 2311 3494
rect 2315 3490 2479 3494
rect 2483 3490 2639 3494
rect 2643 3490 2799 3494
rect 2803 3490 2967 3494
rect 2971 3490 3463 3494
rect 3467 3490 3499 3494
rect 1797 3489 3499 3490
rect 3505 3489 3506 3495
rect 84 3433 85 3439
rect 91 3438 1779 3439
rect 91 3434 111 3438
rect 115 3434 135 3438
rect 139 3434 255 3438
rect 259 3434 271 3438
rect 275 3434 415 3438
rect 419 3434 439 3438
rect 443 3434 575 3438
rect 579 3434 615 3438
rect 619 3434 735 3438
rect 739 3434 791 3438
rect 795 3434 895 3438
rect 899 3434 959 3438
rect 963 3434 1063 3438
rect 1067 3434 1119 3438
rect 1123 3434 1231 3438
rect 1235 3434 1263 3438
rect 1267 3434 1399 3438
rect 1403 3434 1407 3438
rect 1411 3434 1551 3438
rect 1555 3434 1671 3438
rect 1675 3434 1767 3438
rect 1771 3434 1779 3438
rect 91 3433 1779 3434
rect 1785 3433 1786 3439
rect 1778 3431 1786 3433
rect 1778 3425 1779 3431
rect 1785 3430 3487 3431
rect 1785 3426 1807 3430
rect 1811 3426 1831 3430
rect 1835 3426 1975 3430
rect 1979 3426 2031 3430
rect 2035 3426 2143 3430
rect 2147 3426 2151 3430
rect 2155 3426 2271 3430
rect 2275 3426 2311 3430
rect 2315 3426 2391 3430
rect 2395 3426 2479 3430
rect 2483 3426 2511 3430
rect 2515 3426 2623 3430
rect 2627 3426 2639 3430
rect 2643 3426 2727 3430
rect 2731 3426 2799 3430
rect 2803 3426 2831 3430
rect 2835 3426 2935 3430
rect 2939 3426 2967 3430
rect 2971 3426 3039 3430
rect 3043 3426 3151 3430
rect 3155 3426 3463 3430
rect 3467 3426 3487 3430
rect 1785 3425 3487 3426
rect 3493 3425 3494 3431
rect 96 3361 97 3367
rect 103 3366 1791 3367
rect 103 3362 111 3366
rect 115 3362 135 3366
rect 139 3362 255 3366
rect 259 3362 327 3366
rect 331 3362 415 3366
rect 419 3362 535 3366
rect 539 3362 575 3366
rect 579 3362 735 3366
rect 739 3362 743 3366
rect 747 3362 895 3366
rect 899 3362 935 3366
rect 939 3362 1063 3366
rect 1067 3362 1119 3366
rect 1123 3362 1231 3366
rect 1235 3362 1295 3366
rect 1299 3362 1399 3366
rect 1403 3362 1463 3366
rect 1467 3362 1639 3366
rect 1643 3362 1767 3366
rect 1771 3362 1791 3366
rect 103 3361 1791 3362
rect 1797 3363 1798 3367
rect 1797 3362 3506 3363
rect 1797 3361 1807 3362
rect 1790 3358 1807 3361
rect 1811 3358 2031 3362
rect 2035 3358 2151 3362
rect 2155 3358 2159 3362
rect 2163 3358 2271 3362
rect 2275 3358 2295 3362
rect 2299 3358 2391 3362
rect 2395 3358 2431 3362
rect 2435 3358 2511 3362
rect 2515 3358 2567 3362
rect 2571 3358 2623 3362
rect 2627 3358 2703 3362
rect 2707 3358 2727 3362
rect 2731 3358 2831 3362
rect 2835 3358 2839 3362
rect 2843 3358 2935 3362
rect 2939 3358 2975 3362
rect 2979 3358 3039 3362
rect 3043 3358 3119 3362
rect 3123 3358 3151 3362
rect 3155 3358 3463 3362
rect 3467 3358 3506 3362
rect 1790 3357 3506 3358
rect 1778 3298 3494 3299
rect 1778 3295 1807 3298
rect 84 3289 85 3295
rect 91 3294 1779 3295
rect 91 3290 111 3294
rect 115 3290 135 3294
rect 139 3290 279 3294
rect 283 3290 327 3294
rect 331 3290 463 3294
rect 467 3290 535 3294
rect 539 3290 647 3294
rect 651 3290 743 3294
rect 747 3290 831 3294
rect 835 3290 935 3294
rect 939 3290 1007 3294
rect 1011 3290 1119 3294
rect 1123 3290 1175 3294
rect 1179 3290 1295 3294
rect 1299 3290 1343 3294
rect 1347 3290 1463 3294
rect 1467 3290 1503 3294
rect 1507 3290 1639 3294
rect 1643 3290 1671 3294
rect 1675 3290 1767 3294
rect 1771 3290 1779 3294
rect 91 3289 1779 3290
rect 1785 3294 1807 3295
rect 1811 3294 2087 3298
rect 2091 3294 2159 3298
rect 2163 3294 2239 3298
rect 2243 3294 2295 3298
rect 2299 3294 2399 3298
rect 2403 3294 2431 3298
rect 2435 3294 2559 3298
rect 2563 3294 2567 3298
rect 2571 3294 2703 3298
rect 2707 3294 2719 3298
rect 2723 3294 2839 3298
rect 2843 3294 2879 3298
rect 2883 3294 2975 3298
rect 2979 3294 3039 3298
rect 3043 3294 3119 3298
rect 3123 3294 3199 3298
rect 3203 3294 3463 3298
rect 3467 3294 3494 3298
rect 1785 3293 3494 3294
rect 1785 3289 1786 3293
rect 1790 3225 1791 3231
rect 1797 3230 3499 3231
rect 1797 3226 1807 3230
rect 1811 3226 1911 3230
rect 1915 3226 2047 3230
rect 2051 3226 2087 3230
rect 2091 3226 2199 3230
rect 2203 3226 2239 3230
rect 2243 3226 2359 3230
rect 2363 3226 2399 3230
rect 2403 3226 2527 3230
rect 2531 3226 2559 3230
rect 2563 3226 2687 3230
rect 2691 3226 2719 3230
rect 2723 3226 2847 3230
rect 2851 3226 2879 3230
rect 2883 3226 3007 3230
rect 3011 3226 3039 3230
rect 3043 3226 3167 3230
rect 3171 3226 3199 3230
rect 3203 3226 3335 3230
rect 3339 3226 3463 3230
rect 3467 3226 3499 3230
rect 1797 3225 3499 3226
rect 3505 3225 3506 3231
rect 1790 3223 1798 3225
rect 96 3217 97 3223
rect 103 3222 1791 3223
rect 103 3218 111 3222
rect 115 3218 135 3222
rect 139 3218 183 3222
rect 187 3218 279 3222
rect 283 3218 327 3222
rect 331 3218 463 3222
rect 467 3218 487 3222
rect 491 3218 647 3222
rect 651 3218 807 3222
rect 811 3218 831 3222
rect 835 3218 967 3222
rect 971 3218 1007 3222
rect 1011 3218 1135 3222
rect 1139 3218 1175 3222
rect 1179 3218 1303 3222
rect 1307 3218 1343 3222
rect 1347 3218 1471 3222
rect 1475 3218 1503 3222
rect 1507 3218 1671 3222
rect 1675 3218 1767 3222
rect 1771 3218 1791 3222
rect 103 3217 1791 3218
rect 1797 3217 1798 3223
rect 1778 3161 1779 3167
rect 1785 3166 3487 3167
rect 1785 3162 1807 3166
rect 1811 3162 1831 3166
rect 1835 3162 1911 3166
rect 1915 3162 2007 3166
rect 2011 3162 2047 3166
rect 2051 3162 2199 3166
rect 2203 3162 2207 3166
rect 2211 3162 2359 3166
rect 2363 3162 2399 3166
rect 2403 3162 2527 3166
rect 2531 3162 2583 3166
rect 2587 3162 2687 3166
rect 2691 3162 2759 3166
rect 2763 3162 2847 3166
rect 2851 3162 2919 3166
rect 2923 3162 3007 3166
rect 3011 3162 3079 3166
rect 3083 3162 3167 3166
rect 3171 3162 3231 3166
rect 3235 3162 3335 3166
rect 3339 3162 3367 3166
rect 3371 3162 3463 3166
rect 3467 3162 3487 3166
rect 1785 3161 3487 3162
rect 3493 3161 3494 3167
rect 1778 3159 1786 3161
rect 84 3153 85 3159
rect 91 3158 1779 3159
rect 91 3154 111 3158
rect 115 3154 183 3158
rect 187 3154 327 3158
rect 331 3154 367 3158
rect 371 3154 487 3158
rect 491 3154 607 3158
rect 611 3154 647 3158
rect 651 3154 727 3158
rect 731 3154 807 3158
rect 811 3154 847 3158
rect 851 3154 967 3158
rect 971 3154 1079 3158
rect 1083 3154 1135 3158
rect 1139 3154 1199 3158
rect 1203 3154 1303 3158
rect 1307 3154 1319 3158
rect 1323 3154 1471 3158
rect 1475 3154 1767 3158
rect 1771 3154 1779 3158
rect 91 3153 1779 3154
rect 1785 3153 1786 3159
rect 1790 3094 3506 3095
rect 1790 3091 1807 3094
rect 96 3085 97 3091
rect 103 3090 1791 3091
rect 103 3086 111 3090
rect 115 3086 367 3090
rect 371 3086 439 3090
rect 443 3086 487 3090
rect 491 3086 527 3090
rect 531 3086 607 3090
rect 611 3086 615 3090
rect 619 3086 703 3090
rect 707 3086 727 3090
rect 731 3086 791 3090
rect 795 3086 847 3090
rect 851 3086 879 3090
rect 883 3086 967 3090
rect 971 3086 1055 3090
rect 1059 3086 1079 3090
rect 1083 3086 1143 3090
rect 1147 3086 1199 3090
rect 1203 3086 1319 3090
rect 1323 3086 1767 3090
rect 1771 3086 1791 3090
rect 103 3085 1791 3086
rect 1797 3090 1807 3091
rect 1811 3090 1831 3094
rect 1835 3090 1959 3094
rect 1963 3090 2007 3094
rect 2011 3090 2119 3094
rect 2123 3090 2207 3094
rect 2211 3090 2295 3094
rect 2299 3090 2399 3094
rect 2403 3090 2487 3094
rect 2491 3090 2583 3094
rect 2587 3090 2695 3094
rect 2699 3090 2759 3094
rect 2763 3090 2919 3094
rect 2923 3090 3079 3094
rect 3083 3090 3151 3094
rect 3155 3090 3231 3094
rect 3235 3090 3367 3094
rect 3371 3090 3463 3094
rect 3467 3090 3506 3094
rect 1797 3089 3506 3090
rect 1797 3085 1798 3089
rect 84 3013 85 3019
rect 91 3018 1779 3019
rect 91 3014 111 3018
rect 115 3014 439 3018
rect 443 3014 503 3018
rect 507 3014 527 3018
rect 531 3014 591 3018
rect 595 3014 615 3018
rect 619 3014 679 3018
rect 683 3014 703 3018
rect 707 3014 767 3018
rect 771 3014 791 3018
rect 795 3014 855 3018
rect 859 3014 879 3018
rect 883 3014 943 3018
rect 947 3014 967 3018
rect 971 3014 1031 3018
rect 1035 3014 1055 3018
rect 1059 3014 1119 3018
rect 1123 3014 1143 3018
rect 1147 3014 1207 3018
rect 1211 3014 1295 3018
rect 1299 3014 1767 3018
rect 1771 3014 1779 3018
rect 91 3013 1779 3014
rect 1785 3015 1786 3019
rect 1785 3014 3494 3015
rect 1785 3013 1807 3014
rect 1778 3010 1807 3013
rect 1811 3010 1831 3014
rect 1835 3010 1919 3014
rect 1923 3010 1959 3014
rect 1963 3010 2031 3014
rect 2035 3010 2119 3014
rect 2123 3010 2143 3014
rect 2147 3010 2247 3014
rect 2251 3010 2295 3014
rect 2299 3010 2359 3014
rect 2363 3010 2479 3014
rect 2483 3010 2487 3014
rect 2491 3010 2623 3014
rect 2627 3010 2695 3014
rect 2699 3010 2791 3014
rect 2795 3010 2919 3014
rect 2923 3010 2983 3014
rect 2987 3010 3151 3014
rect 3155 3010 3183 3014
rect 3187 3010 3367 3014
rect 3371 3010 3463 3014
rect 3467 3010 3494 3014
rect 1778 3009 3494 3010
rect 96 2937 97 2943
rect 103 2942 1791 2943
rect 103 2938 111 2942
rect 115 2938 327 2942
rect 331 2938 447 2942
rect 451 2938 503 2942
rect 507 2938 575 2942
rect 579 2938 591 2942
rect 595 2938 679 2942
rect 683 2938 711 2942
rect 715 2938 767 2942
rect 771 2938 847 2942
rect 851 2938 855 2942
rect 859 2938 943 2942
rect 947 2938 975 2942
rect 979 2938 1031 2942
rect 1035 2938 1103 2942
rect 1107 2938 1119 2942
rect 1123 2938 1207 2942
rect 1211 2938 1231 2942
rect 1235 2938 1295 2942
rect 1299 2938 1359 2942
rect 1363 2938 1495 2942
rect 1499 2938 1767 2942
rect 1771 2938 1791 2942
rect 103 2937 1791 2938
rect 1797 2939 1798 2943
rect 1797 2938 3506 2939
rect 1797 2937 1807 2938
rect 1790 2934 1807 2937
rect 1811 2934 1831 2938
rect 1835 2934 1919 2938
rect 1923 2934 2015 2938
rect 2019 2934 2031 2938
rect 2035 2934 2143 2938
rect 2147 2934 2215 2938
rect 2219 2934 2247 2938
rect 2251 2934 2359 2938
rect 2363 2934 2407 2938
rect 2411 2934 2479 2938
rect 2483 2934 2591 2938
rect 2595 2934 2623 2938
rect 2627 2934 2759 2938
rect 2763 2934 2791 2938
rect 2795 2934 2911 2938
rect 2915 2934 2983 2938
rect 2987 2934 3063 2938
rect 3067 2934 3183 2938
rect 3187 2934 3207 2938
rect 3211 2934 3359 2938
rect 3363 2934 3367 2938
rect 3371 2934 3463 2938
rect 3467 2934 3506 2938
rect 1790 2933 3506 2934
rect 1778 2874 3494 2875
rect 1778 2871 1807 2874
rect 84 2865 85 2871
rect 91 2870 1779 2871
rect 91 2866 111 2870
rect 115 2866 135 2870
rect 139 2866 255 2870
rect 259 2866 327 2870
rect 331 2866 415 2870
rect 419 2866 447 2870
rect 451 2866 575 2870
rect 579 2866 711 2870
rect 715 2866 735 2870
rect 739 2866 847 2870
rect 851 2866 895 2870
rect 899 2866 975 2870
rect 979 2866 1047 2870
rect 1051 2866 1103 2870
rect 1107 2866 1191 2870
rect 1195 2866 1231 2870
rect 1235 2866 1343 2870
rect 1347 2866 1359 2870
rect 1363 2866 1495 2870
rect 1499 2866 1767 2870
rect 1771 2866 1779 2870
rect 91 2865 1779 2866
rect 1785 2870 1807 2871
rect 1811 2870 1831 2874
rect 1835 2870 1999 2874
rect 2003 2870 2015 2874
rect 2019 2870 2191 2874
rect 2195 2870 2215 2874
rect 2219 2870 2383 2874
rect 2387 2870 2407 2874
rect 2411 2870 2567 2874
rect 2571 2870 2591 2874
rect 2595 2870 2735 2874
rect 2739 2870 2759 2874
rect 2763 2870 2903 2874
rect 2907 2870 2911 2874
rect 2915 2870 3063 2874
rect 3067 2870 3207 2874
rect 3211 2870 3223 2874
rect 3227 2870 3359 2874
rect 3363 2870 3367 2874
rect 3371 2870 3463 2874
rect 3467 2870 3494 2874
rect 1785 2869 3494 2870
rect 1785 2865 1786 2869
rect 1790 2801 1791 2807
rect 1797 2806 3499 2807
rect 1797 2802 1807 2806
rect 1811 2802 1831 2806
rect 1835 2802 1999 2806
rect 2003 2802 2015 2806
rect 2019 2802 2191 2806
rect 2195 2802 2215 2806
rect 2219 2802 2383 2806
rect 2387 2802 2407 2806
rect 2411 2802 2567 2806
rect 2571 2802 2583 2806
rect 2587 2802 2735 2806
rect 2739 2802 2751 2806
rect 2755 2802 2903 2806
rect 2907 2802 2911 2806
rect 2915 2802 3063 2806
rect 3067 2802 3071 2806
rect 3075 2802 3223 2806
rect 3227 2802 3231 2806
rect 3235 2802 3367 2806
rect 3371 2802 3463 2806
rect 3467 2802 3499 2806
rect 1797 2801 3499 2802
rect 3505 2801 3506 2807
rect 96 2789 97 2795
rect 103 2794 1791 2795
rect 103 2790 111 2794
rect 115 2790 135 2794
rect 139 2790 247 2794
rect 251 2790 255 2794
rect 259 2790 391 2794
rect 395 2790 415 2794
rect 419 2790 543 2794
rect 547 2790 575 2794
rect 579 2790 695 2794
rect 699 2790 735 2794
rect 739 2790 855 2794
rect 859 2790 895 2794
rect 899 2790 1023 2794
rect 1027 2790 1047 2794
rect 1051 2790 1191 2794
rect 1195 2790 1343 2794
rect 1347 2790 1359 2794
rect 1363 2790 1495 2794
rect 1499 2790 1527 2794
rect 1531 2790 1671 2794
rect 1675 2790 1767 2794
rect 1771 2790 1791 2794
rect 103 2789 1791 2790
rect 1797 2789 1798 2795
rect 1778 2726 3494 2727
rect 1778 2723 1807 2726
rect 84 2717 85 2723
rect 91 2722 1779 2723
rect 91 2718 111 2722
rect 115 2718 135 2722
rect 139 2718 247 2722
rect 251 2718 359 2722
rect 363 2718 391 2722
rect 395 2718 479 2722
rect 483 2718 543 2722
rect 547 2718 615 2722
rect 619 2718 695 2722
rect 699 2718 759 2722
rect 763 2718 855 2722
rect 859 2718 911 2722
rect 915 2718 1023 2722
rect 1027 2718 1063 2722
rect 1067 2718 1191 2722
rect 1195 2718 1215 2722
rect 1219 2718 1359 2722
rect 1363 2718 1375 2722
rect 1379 2718 1527 2722
rect 1531 2718 1535 2722
rect 1539 2718 1671 2722
rect 1675 2718 1767 2722
rect 1771 2718 1779 2722
rect 91 2717 1779 2718
rect 1785 2722 1807 2723
rect 1811 2722 1831 2726
rect 1835 2722 2015 2726
rect 2019 2722 2039 2726
rect 2043 2722 2159 2726
rect 2163 2722 2215 2726
rect 2219 2722 2279 2726
rect 2283 2722 2407 2726
rect 2411 2722 2543 2726
rect 2547 2722 2583 2726
rect 2587 2722 2687 2726
rect 2691 2722 2751 2726
rect 2755 2722 2847 2726
rect 2851 2722 2911 2726
rect 2915 2722 3023 2726
rect 3027 2722 3071 2726
rect 3075 2722 3207 2726
rect 3211 2722 3231 2726
rect 3235 2722 3367 2726
rect 3371 2722 3463 2726
rect 3467 2722 3494 2726
rect 1785 2721 3494 2722
rect 1785 2717 1786 2721
rect 96 2645 97 2651
rect 103 2650 1791 2651
rect 103 2646 111 2650
rect 115 2646 247 2650
rect 251 2646 359 2650
rect 363 2646 463 2650
rect 467 2646 479 2650
rect 483 2646 551 2650
rect 555 2646 615 2650
rect 619 2646 639 2650
rect 643 2646 743 2650
rect 747 2646 759 2650
rect 763 2646 855 2650
rect 859 2646 911 2650
rect 915 2646 983 2650
rect 987 2646 1063 2650
rect 1067 2646 1127 2650
rect 1131 2646 1215 2650
rect 1219 2646 1279 2650
rect 1283 2646 1375 2650
rect 1379 2646 1439 2650
rect 1443 2646 1535 2650
rect 1539 2646 1607 2650
rect 1611 2646 1671 2650
rect 1675 2646 1767 2650
rect 1771 2646 1791 2650
rect 103 2645 1791 2646
rect 1797 2650 3506 2651
rect 1797 2646 1807 2650
rect 1811 2646 1871 2650
rect 1875 2646 1967 2650
rect 1971 2646 2039 2650
rect 2043 2646 2071 2650
rect 2075 2646 2159 2650
rect 2163 2646 2183 2650
rect 2187 2646 2279 2650
rect 2283 2646 2295 2650
rect 2299 2646 2407 2650
rect 2411 2646 2431 2650
rect 2435 2646 2543 2650
rect 2547 2646 2583 2650
rect 2587 2646 2687 2650
rect 2691 2646 2759 2650
rect 2763 2646 2847 2650
rect 2851 2646 2959 2650
rect 2963 2646 3023 2650
rect 3027 2646 3167 2650
rect 3171 2646 3207 2650
rect 3211 2646 3367 2650
rect 3371 2646 3463 2650
rect 3467 2646 3506 2650
rect 1797 2645 3506 2646
rect 84 2573 85 2579
rect 91 2578 1779 2579
rect 91 2574 111 2578
rect 115 2574 463 2578
rect 467 2574 503 2578
rect 507 2574 551 2578
rect 555 2574 591 2578
rect 595 2574 639 2578
rect 643 2574 679 2578
rect 683 2574 743 2578
rect 747 2574 775 2578
rect 779 2574 855 2578
rect 859 2574 879 2578
rect 883 2574 983 2578
rect 987 2574 991 2578
rect 995 2574 1103 2578
rect 1107 2574 1127 2578
rect 1131 2574 1223 2578
rect 1227 2574 1279 2578
rect 1283 2574 1351 2578
rect 1355 2574 1439 2578
rect 1443 2574 1479 2578
rect 1483 2574 1607 2578
rect 1611 2574 1767 2578
rect 1771 2574 1779 2578
rect 91 2573 1779 2574
rect 1785 2575 1786 2579
rect 1785 2574 3494 2575
rect 1785 2573 1807 2574
rect 1778 2570 1807 2573
rect 1811 2570 1831 2574
rect 1835 2570 1871 2574
rect 1875 2570 1919 2574
rect 1923 2570 1967 2574
rect 1971 2570 2007 2574
rect 2011 2570 2071 2574
rect 2075 2570 2111 2574
rect 2115 2570 2183 2574
rect 2187 2570 2223 2574
rect 2227 2570 2295 2574
rect 2299 2570 2343 2574
rect 2347 2570 2431 2574
rect 2435 2570 2487 2574
rect 2491 2570 2583 2574
rect 2587 2570 2647 2574
rect 2651 2570 2759 2574
rect 2763 2570 2815 2574
rect 2819 2570 2959 2574
rect 2963 2570 2999 2574
rect 3003 2570 3167 2574
rect 3171 2570 3191 2574
rect 3195 2570 3367 2574
rect 3371 2570 3463 2574
rect 3467 2570 3494 2574
rect 1778 2569 3494 2570
rect 1790 2510 3506 2511
rect 1790 2507 1807 2510
rect 96 2501 97 2507
rect 103 2506 1791 2507
rect 103 2502 111 2506
rect 115 2502 503 2506
rect 507 2502 551 2506
rect 555 2502 591 2506
rect 595 2502 679 2506
rect 683 2502 735 2506
rect 739 2502 775 2506
rect 779 2502 879 2506
rect 883 2502 911 2506
rect 915 2502 991 2506
rect 995 2502 1079 2506
rect 1083 2502 1103 2506
rect 1107 2502 1223 2506
rect 1227 2502 1239 2506
rect 1243 2502 1351 2506
rect 1355 2502 1399 2506
rect 1403 2502 1479 2506
rect 1483 2502 1567 2506
rect 1571 2502 1607 2506
rect 1611 2502 1767 2506
rect 1771 2502 1791 2506
rect 103 2501 1791 2502
rect 1797 2506 1807 2507
rect 1811 2506 1831 2510
rect 1835 2506 1919 2510
rect 1923 2506 1951 2510
rect 1955 2506 2007 2510
rect 2011 2506 2039 2510
rect 2043 2506 2111 2510
rect 2115 2506 2135 2510
rect 2139 2506 2223 2510
rect 2227 2506 2239 2510
rect 2243 2506 2343 2510
rect 2347 2506 2367 2510
rect 2371 2506 2487 2510
rect 2491 2506 2527 2510
rect 2531 2506 2647 2510
rect 2651 2506 2711 2510
rect 2715 2506 2815 2510
rect 2819 2506 2919 2510
rect 2923 2506 2999 2510
rect 3003 2506 3143 2510
rect 3147 2506 3191 2510
rect 3195 2506 3367 2510
rect 3371 2506 3463 2510
rect 3467 2506 3506 2510
rect 1797 2505 3506 2506
rect 1797 2501 1798 2505
rect 2014 2500 2020 2501
rect 2214 2500 2220 2501
rect 2014 2496 2015 2500
rect 2019 2496 2215 2500
rect 2219 2496 2220 2500
rect 2014 2495 2020 2496
rect 2214 2495 2220 2496
rect 84 2437 85 2443
rect 91 2442 1779 2443
rect 91 2438 111 2442
rect 115 2438 415 2442
rect 419 2438 503 2442
rect 507 2438 551 2442
rect 555 2438 599 2442
rect 603 2438 703 2442
rect 707 2438 735 2442
rect 739 2438 807 2442
rect 811 2438 911 2442
rect 915 2438 919 2442
rect 923 2438 1039 2442
rect 1043 2438 1079 2442
rect 1083 2438 1167 2442
rect 1171 2438 1239 2442
rect 1243 2438 1295 2442
rect 1299 2438 1399 2442
rect 1403 2438 1423 2442
rect 1427 2438 1567 2442
rect 1571 2438 1767 2442
rect 1771 2438 1779 2442
rect 91 2437 1779 2438
rect 1785 2439 1786 2443
rect 1785 2438 3494 2439
rect 1785 2437 1807 2438
rect 1778 2434 1807 2437
rect 1811 2434 1951 2438
rect 1955 2434 2039 2438
rect 2043 2434 2135 2438
rect 2139 2434 2215 2438
rect 2219 2434 2239 2438
rect 2243 2434 2303 2438
rect 2307 2434 2367 2438
rect 2371 2434 2391 2438
rect 2395 2434 2479 2438
rect 2483 2434 2527 2438
rect 2531 2434 2567 2438
rect 2571 2434 2655 2438
rect 2659 2434 2711 2438
rect 2715 2434 2743 2438
rect 2747 2434 2839 2438
rect 2843 2434 2919 2438
rect 2923 2434 2935 2438
rect 2939 2434 3143 2438
rect 3147 2434 3367 2438
rect 3371 2434 3463 2438
rect 3467 2434 3494 2438
rect 1778 2433 3494 2434
rect 96 2369 97 2375
rect 103 2374 1791 2375
rect 103 2370 111 2374
rect 115 2370 319 2374
rect 323 2370 415 2374
rect 419 2370 431 2374
rect 435 2370 503 2374
rect 507 2370 543 2374
rect 547 2370 599 2374
rect 603 2370 655 2374
rect 659 2370 703 2374
rect 707 2370 767 2374
rect 771 2370 807 2374
rect 811 2370 879 2374
rect 883 2370 919 2374
rect 923 2370 991 2374
rect 995 2370 1039 2374
rect 1043 2370 1103 2374
rect 1107 2370 1167 2374
rect 1171 2370 1215 2374
rect 1219 2370 1295 2374
rect 1299 2370 1335 2374
rect 1339 2370 1423 2374
rect 1427 2370 1767 2374
rect 1771 2370 1791 2374
rect 103 2369 1791 2370
rect 1797 2374 3506 2375
rect 1797 2370 1807 2374
rect 1811 2370 2167 2374
rect 2171 2370 2215 2374
rect 2219 2370 2263 2374
rect 2267 2370 2303 2374
rect 2307 2370 2367 2374
rect 2371 2370 2391 2374
rect 2395 2370 2471 2374
rect 2475 2370 2479 2374
rect 2483 2370 2567 2374
rect 2571 2370 2575 2374
rect 2579 2370 2655 2374
rect 2659 2370 2687 2374
rect 2691 2370 2743 2374
rect 2747 2370 2799 2374
rect 2803 2370 2839 2374
rect 2843 2370 2911 2374
rect 2915 2370 2935 2374
rect 2939 2370 3023 2374
rect 3027 2370 3463 2374
rect 3467 2370 3506 2374
rect 1797 2369 3506 2370
rect 84 2297 85 2303
rect 91 2302 1779 2303
rect 91 2298 111 2302
rect 115 2298 151 2302
rect 155 2298 271 2302
rect 275 2298 319 2302
rect 323 2298 391 2302
rect 395 2298 431 2302
rect 435 2298 519 2302
rect 523 2298 543 2302
rect 547 2298 647 2302
rect 651 2298 655 2302
rect 659 2298 767 2302
rect 771 2298 775 2302
rect 779 2298 879 2302
rect 883 2298 895 2302
rect 899 2298 991 2302
rect 995 2298 1015 2302
rect 1019 2298 1103 2302
rect 1107 2298 1143 2302
rect 1147 2298 1215 2302
rect 1219 2298 1271 2302
rect 1275 2298 1335 2302
rect 1339 2298 1767 2302
rect 1771 2298 1779 2302
rect 91 2297 1779 2298
rect 1785 2302 3494 2303
rect 1785 2298 1807 2302
rect 1811 2298 1887 2302
rect 1891 2298 2039 2302
rect 2043 2298 2167 2302
rect 2171 2298 2199 2302
rect 2203 2298 2263 2302
rect 2267 2298 2367 2302
rect 2371 2298 2375 2302
rect 2379 2298 2471 2302
rect 2475 2298 2551 2302
rect 2555 2298 2575 2302
rect 2579 2298 2687 2302
rect 2691 2298 2719 2302
rect 2723 2298 2799 2302
rect 2803 2298 2887 2302
rect 2891 2298 2911 2302
rect 2915 2298 3023 2302
rect 3027 2298 3055 2302
rect 3059 2298 3223 2302
rect 3227 2298 3367 2302
rect 3371 2298 3463 2302
rect 3467 2298 3494 2302
rect 1785 2297 3494 2298
rect 1790 2238 3506 2239
rect 1790 2235 1807 2238
rect 96 2229 97 2235
rect 103 2234 1791 2235
rect 103 2230 111 2234
rect 115 2230 135 2234
rect 139 2230 151 2234
rect 155 2230 247 2234
rect 251 2230 271 2234
rect 275 2230 391 2234
rect 395 2230 407 2234
rect 411 2230 519 2234
rect 523 2230 583 2234
rect 587 2230 647 2234
rect 651 2230 767 2234
rect 771 2230 775 2234
rect 779 2230 895 2234
rect 899 2230 951 2234
rect 955 2230 1015 2234
rect 1019 2230 1135 2234
rect 1139 2230 1143 2234
rect 1147 2230 1271 2234
rect 1275 2230 1319 2234
rect 1323 2230 1503 2234
rect 1507 2230 1671 2234
rect 1675 2230 1767 2234
rect 1771 2230 1791 2234
rect 103 2229 1791 2230
rect 1797 2234 1807 2235
rect 1811 2234 1831 2238
rect 1835 2234 1887 2238
rect 1891 2234 1967 2238
rect 1971 2234 2039 2238
rect 2043 2234 2135 2238
rect 2139 2234 2199 2238
rect 2203 2234 2311 2238
rect 2315 2234 2375 2238
rect 2379 2234 2487 2238
rect 2491 2234 2551 2238
rect 2555 2234 2655 2238
rect 2659 2234 2719 2238
rect 2723 2234 2815 2238
rect 2819 2234 2887 2238
rect 2891 2234 2959 2238
rect 2963 2234 3055 2238
rect 3059 2234 3103 2238
rect 3107 2234 3223 2238
rect 3227 2234 3247 2238
rect 3251 2234 3367 2238
rect 3371 2234 3463 2238
rect 3467 2234 3506 2238
rect 1797 2233 3506 2234
rect 1797 2229 1798 2233
rect 1778 2169 1779 2175
rect 1785 2174 3487 2175
rect 1785 2170 1807 2174
rect 1811 2170 1831 2174
rect 1835 2170 1967 2174
rect 1971 2170 2135 2174
rect 2139 2170 2311 2174
rect 2315 2170 2487 2174
rect 2491 2170 2655 2174
rect 2659 2170 2815 2174
rect 2819 2170 2927 2174
rect 2931 2170 2959 2174
rect 2963 2170 3015 2174
rect 3019 2170 3103 2174
rect 3107 2170 3191 2174
rect 3195 2170 3247 2174
rect 3251 2170 3279 2174
rect 3283 2170 3367 2174
rect 3371 2170 3463 2174
rect 3467 2170 3487 2174
rect 1785 2169 3487 2170
rect 3493 2169 3494 2175
rect 84 2157 85 2163
rect 91 2162 1779 2163
rect 91 2158 111 2162
rect 115 2158 135 2162
rect 139 2158 247 2162
rect 251 2158 391 2162
rect 395 2158 407 2162
rect 411 2158 543 2162
rect 547 2158 583 2162
rect 587 2158 695 2162
rect 699 2158 767 2162
rect 771 2158 839 2162
rect 843 2158 951 2162
rect 955 2158 975 2162
rect 979 2158 1103 2162
rect 1107 2158 1135 2162
rect 1139 2158 1231 2162
rect 1235 2158 1319 2162
rect 1323 2158 1351 2162
rect 1355 2158 1463 2162
rect 1467 2158 1503 2162
rect 1507 2158 1575 2162
rect 1579 2158 1671 2162
rect 1675 2158 1767 2162
rect 1771 2158 1779 2162
rect 91 2157 1779 2158
rect 1785 2157 1786 2163
rect 1790 2097 1791 2103
rect 1797 2102 3499 2103
rect 1797 2098 1807 2102
rect 1811 2098 1831 2102
rect 1835 2098 1991 2102
rect 1995 2098 2167 2102
rect 2171 2098 2343 2102
rect 2347 2098 2503 2102
rect 2507 2098 2655 2102
rect 2659 2098 2791 2102
rect 2795 2098 2919 2102
rect 2923 2098 2927 2102
rect 2931 2098 3015 2102
rect 3019 2098 3039 2102
rect 3043 2098 3103 2102
rect 3107 2098 3159 2102
rect 3163 2098 3191 2102
rect 3195 2098 3271 2102
rect 3275 2098 3279 2102
rect 3283 2098 3367 2102
rect 3371 2098 3463 2102
rect 3467 2098 3499 2102
rect 1797 2097 3499 2098
rect 3505 2097 3506 2103
rect 1790 2095 1798 2097
rect 96 2089 97 2095
rect 103 2094 1791 2095
rect 103 2090 111 2094
rect 115 2090 135 2094
rect 139 2090 223 2094
rect 227 2090 247 2094
rect 251 2090 343 2094
rect 347 2090 391 2094
rect 395 2090 463 2094
rect 467 2090 543 2094
rect 547 2090 583 2094
rect 587 2090 695 2094
rect 699 2090 703 2094
rect 707 2090 823 2094
rect 827 2090 839 2094
rect 843 2090 935 2094
rect 939 2090 975 2094
rect 979 2090 1047 2094
rect 1051 2090 1103 2094
rect 1107 2090 1159 2094
rect 1163 2090 1231 2094
rect 1235 2090 1279 2094
rect 1283 2090 1351 2094
rect 1355 2090 1463 2094
rect 1467 2090 1575 2094
rect 1579 2090 1671 2094
rect 1675 2090 1767 2094
rect 1771 2090 1791 2094
rect 103 2089 1791 2090
rect 1797 2089 1798 2095
rect 1778 2029 1779 2035
rect 1785 2034 3487 2035
rect 1785 2030 1807 2034
rect 1811 2030 1831 2034
rect 1835 2030 1991 2034
rect 1995 2030 2015 2034
rect 2019 2030 2167 2034
rect 2171 2030 2223 2034
rect 2227 2030 2343 2034
rect 2347 2030 2431 2034
rect 2435 2030 2503 2034
rect 2507 2030 2631 2034
rect 2635 2030 2655 2034
rect 2659 2030 2791 2034
rect 2795 2030 2823 2034
rect 2827 2030 2919 2034
rect 2923 2030 3007 2034
rect 3011 2030 3039 2034
rect 3043 2030 3159 2034
rect 3163 2030 3199 2034
rect 3203 2030 3271 2034
rect 3275 2030 3367 2034
rect 3371 2030 3463 2034
rect 3467 2030 3487 2034
rect 1785 2029 3487 2030
rect 3493 2029 3494 2035
rect 84 2017 85 2023
rect 91 2022 1779 2023
rect 91 2018 111 2022
rect 115 2018 135 2022
rect 139 2018 223 2022
rect 227 2018 239 2022
rect 243 2018 343 2022
rect 347 2018 367 2022
rect 371 2018 463 2022
rect 467 2018 503 2022
rect 507 2018 583 2022
rect 587 2018 639 2022
rect 643 2018 703 2022
rect 707 2018 775 2022
rect 779 2018 823 2022
rect 827 2018 911 2022
rect 915 2018 935 2022
rect 939 2018 1047 2022
rect 1051 2018 1159 2022
rect 1163 2018 1183 2022
rect 1187 2018 1279 2022
rect 1283 2018 1327 2022
rect 1331 2018 1767 2022
rect 1771 2018 1779 2022
rect 91 2017 1779 2018
rect 1785 2017 1786 2023
rect 1790 1961 1791 1967
rect 1797 1966 3499 1967
rect 1797 1962 1807 1966
rect 1811 1962 1831 1966
rect 1835 1962 1863 1966
rect 1867 1962 1999 1966
rect 2003 1962 2015 1966
rect 2019 1962 2143 1966
rect 2147 1962 2223 1966
rect 2227 1962 2287 1966
rect 2291 1962 2431 1966
rect 2435 1962 2575 1966
rect 2579 1962 2631 1966
rect 2635 1962 2711 1966
rect 2715 1962 2823 1966
rect 2827 1962 2831 1966
rect 2835 1962 2951 1966
rect 2955 1962 3007 1966
rect 3011 1962 3063 1966
rect 3067 1962 3167 1966
rect 3171 1962 3199 1966
rect 3203 1962 3279 1966
rect 3283 1962 3367 1966
rect 3371 1962 3463 1966
rect 3467 1962 3499 1966
rect 1797 1961 3499 1962
rect 3505 1961 3506 1967
rect 96 1949 97 1955
rect 103 1954 1791 1955
rect 103 1950 111 1954
rect 115 1950 135 1954
rect 139 1950 239 1954
rect 243 1950 295 1954
rect 299 1950 367 1954
rect 371 1950 423 1954
rect 427 1950 503 1954
rect 507 1950 559 1954
rect 563 1950 639 1954
rect 643 1950 703 1954
rect 707 1950 775 1954
rect 779 1950 855 1954
rect 859 1950 911 1954
rect 915 1950 1007 1954
rect 1011 1950 1047 1954
rect 1051 1950 1159 1954
rect 1163 1950 1183 1954
rect 1187 1950 1311 1954
rect 1315 1950 1327 1954
rect 1331 1950 1471 1954
rect 1475 1950 1767 1954
rect 1771 1950 1791 1954
rect 103 1949 1791 1950
rect 1797 1949 1798 1955
rect 1778 1893 1779 1899
rect 1785 1898 3487 1899
rect 1785 1894 1807 1898
rect 1811 1894 1863 1898
rect 1867 1894 1999 1898
rect 2003 1894 2015 1898
rect 2019 1894 2111 1898
rect 2115 1894 2143 1898
rect 2147 1894 2215 1898
rect 2219 1894 2287 1898
rect 2291 1894 2327 1898
rect 2331 1894 2431 1898
rect 2435 1894 2439 1898
rect 2443 1894 2543 1898
rect 2547 1894 2575 1898
rect 2579 1894 2647 1898
rect 2651 1894 2711 1898
rect 2715 1894 2759 1898
rect 2763 1894 2831 1898
rect 2835 1894 2871 1898
rect 2875 1894 2951 1898
rect 2955 1894 2983 1898
rect 2987 1894 3063 1898
rect 3067 1894 3167 1898
rect 3171 1894 3279 1898
rect 3283 1894 3367 1898
rect 3371 1894 3463 1898
rect 3467 1894 3487 1898
rect 1785 1893 3487 1894
rect 3493 1893 3494 1899
rect 1778 1891 1786 1893
rect 84 1885 85 1891
rect 91 1890 1779 1891
rect 91 1886 111 1890
rect 115 1886 295 1890
rect 299 1886 423 1890
rect 427 1886 431 1890
rect 435 1886 559 1890
rect 563 1886 575 1890
rect 579 1886 703 1890
rect 707 1886 727 1890
rect 731 1886 855 1890
rect 859 1886 887 1890
rect 891 1886 1007 1890
rect 1011 1886 1047 1890
rect 1051 1886 1159 1890
rect 1163 1886 1199 1890
rect 1203 1886 1311 1890
rect 1315 1886 1351 1890
rect 1355 1886 1471 1890
rect 1475 1886 1511 1890
rect 1515 1886 1671 1890
rect 1675 1886 1767 1890
rect 1771 1886 1779 1890
rect 91 1885 1779 1886
rect 1785 1885 1786 1891
rect 1790 1826 3506 1827
rect 1790 1823 1807 1826
rect 96 1817 97 1823
rect 103 1822 1791 1823
rect 103 1818 111 1822
rect 115 1818 431 1822
rect 435 1818 511 1822
rect 515 1818 575 1822
rect 579 1818 631 1822
rect 635 1818 727 1822
rect 731 1818 759 1822
rect 763 1818 887 1822
rect 891 1818 1023 1822
rect 1027 1818 1047 1822
rect 1051 1818 1151 1822
rect 1155 1818 1199 1822
rect 1203 1818 1279 1822
rect 1283 1818 1351 1822
rect 1355 1818 1407 1822
rect 1411 1818 1511 1822
rect 1515 1818 1535 1822
rect 1539 1818 1671 1822
rect 1675 1818 1767 1822
rect 1771 1818 1791 1822
rect 103 1817 1791 1818
rect 1797 1822 1807 1823
rect 1811 1822 2015 1826
rect 2019 1822 2103 1826
rect 2107 1822 2111 1826
rect 2115 1822 2191 1826
rect 2195 1822 2215 1826
rect 2219 1822 2279 1826
rect 2283 1822 2327 1826
rect 2331 1822 2367 1826
rect 2371 1822 2439 1826
rect 2443 1822 2455 1826
rect 2459 1822 2543 1826
rect 2547 1822 2631 1826
rect 2635 1822 2647 1826
rect 2651 1822 2719 1826
rect 2723 1822 2759 1826
rect 2763 1822 2807 1826
rect 2811 1822 2871 1826
rect 2875 1822 2895 1826
rect 2899 1822 2983 1826
rect 2987 1822 3463 1826
rect 3467 1822 3506 1826
rect 1797 1821 3506 1822
rect 1797 1817 1798 1821
rect 84 1749 85 1755
rect 91 1754 1779 1755
rect 91 1750 111 1754
rect 115 1750 439 1754
rect 443 1750 511 1754
rect 515 1750 535 1754
rect 539 1750 631 1754
rect 635 1750 639 1754
rect 643 1750 743 1754
rect 747 1750 759 1754
rect 763 1750 847 1754
rect 851 1750 887 1754
rect 891 1750 951 1754
rect 955 1750 1023 1754
rect 1027 1750 1055 1754
rect 1059 1750 1151 1754
rect 1155 1750 1159 1754
rect 1163 1750 1271 1754
rect 1275 1750 1279 1754
rect 1283 1750 1383 1754
rect 1387 1750 1407 1754
rect 1411 1750 1535 1754
rect 1539 1750 1671 1754
rect 1675 1750 1767 1754
rect 1771 1750 1779 1754
rect 91 1749 1779 1750
rect 1785 1751 1786 1755
rect 1785 1750 3494 1751
rect 1785 1749 1807 1750
rect 1778 1746 1807 1749
rect 1811 1746 2103 1750
rect 2107 1746 2143 1750
rect 2147 1746 2191 1750
rect 2195 1746 2231 1750
rect 2235 1746 2279 1750
rect 2283 1746 2319 1750
rect 2323 1746 2367 1750
rect 2371 1746 2407 1750
rect 2411 1746 2455 1750
rect 2459 1746 2495 1750
rect 2499 1746 2543 1750
rect 2547 1746 2583 1750
rect 2587 1746 2631 1750
rect 2635 1746 2671 1750
rect 2675 1746 2719 1750
rect 2723 1746 2759 1750
rect 2763 1746 2807 1750
rect 2811 1746 2847 1750
rect 2851 1746 2895 1750
rect 2899 1746 3463 1750
rect 3467 1746 3494 1750
rect 1778 1745 3494 1746
rect 96 1681 97 1687
rect 103 1686 1791 1687
rect 103 1682 111 1686
rect 115 1682 399 1686
rect 403 1682 439 1686
rect 443 1682 487 1686
rect 491 1682 535 1686
rect 539 1682 575 1686
rect 579 1682 639 1686
rect 643 1682 663 1686
rect 667 1682 743 1686
rect 747 1682 759 1686
rect 763 1682 847 1686
rect 851 1682 855 1686
rect 859 1682 951 1686
rect 955 1682 1047 1686
rect 1051 1682 1055 1686
rect 1059 1682 1143 1686
rect 1147 1682 1159 1686
rect 1163 1682 1271 1686
rect 1275 1682 1383 1686
rect 1387 1682 1767 1686
rect 1771 1682 1791 1686
rect 103 1681 1791 1682
rect 1797 1683 1798 1687
rect 1797 1682 3506 1683
rect 1797 1681 1807 1682
rect 1790 1678 1807 1681
rect 1811 1678 2103 1682
rect 2107 1678 2143 1682
rect 2147 1678 2191 1682
rect 2195 1678 2231 1682
rect 2235 1678 2279 1682
rect 2283 1678 2319 1682
rect 2323 1678 2367 1682
rect 2371 1678 2407 1682
rect 2411 1678 2455 1682
rect 2459 1678 2495 1682
rect 2499 1678 2543 1682
rect 2547 1678 2583 1682
rect 2587 1678 2631 1682
rect 2635 1678 2671 1682
rect 2675 1678 2719 1682
rect 2723 1678 2759 1682
rect 2763 1678 2807 1682
rect 2811 1678 2847 1682
rect 2851 1678 2895 1682
rect 2899 1678 3463 1682
rect 3467 1678 3506 1682
rect 1790 1677 3506 1678
rect 84 1613 85 1619
rect 91 1618 1779 1619
rect 91 1614 111 1618
rect 115 1614 279 1618
rect 283 1614 383 1618
rect 387 1614 399 1618
rect 403 1614 487 1618
rect 491 1614 495 1618
rect 499 1614 575 1618
rect 579 1614 607 1618
rect 611 1614 663 1618
rect 667 1614 719 1618
rect 723 1614 759 1618
rect 763 1614 831 1618
rect 835 1614 855 1618
rect 859 1614 943 1618
rect 947 1614 951 1618
rect 955 1614 1047 1618
rect 1051 1614 1055 1618
rect 1059 1614 1143 1618
rect 1147 1614 1167 1618
rect 1171 1614 1279 1618
rect 1283 1614 1767 1618
rect 1771 1614 1779 1618
rect 91 1613 1779 1614
rect 1785 1615 1786 1619
rect 1785 1614 3494 1615
rect 1785 1613 1807 1614
rect 1778 1610 1807 1613
rect 1811 1610 2063 1614
rect 2067 1610 2103 1614
rect 2107 1610 2159 1614
rect 2163 1610 2191 1614
rect 2195 1610 2255 1614
rect 2259 1610 2279 1614
rect 2283 1610 2359 1614
rect 2363 1610 2367 1614
rect 2371 1610 2455 1614
rect 2459 1610 2463 1614
rect 2467 1610 2543 1614
rect 2547 1610 2567 1614
rect 2571 1610 2631 1614
rect 2635 1610 2671 1614
rect 2675 1610 2719 1614
rect 2723 1610 2775 1614
rect 2779 1610 2807 1614
rect 2811 1610 2887 1614
rect 2891 1610 2895 1614
rect 2899 1610 3463 1614
rect 3467 1610 3494 1614
rect 1778 1609 3494 1610
rect 1790 1550 3506 1551
rect 1790 1547 1807 1550
rect 96 1541 97 1547
rect 103 1546 1791 1547
rect 103 1542 111 1546
rect 115 1542 183 1546
rect 187 1542 279 1546
rect 283 1542 327 1546
rect 331 1542 383 1546
rect 387 1542 471 1546
rect 475 1542 495 1546
rect 499 1542 607 1546
rect 611 1542 623 1546
rect 627 1542 719 1546
rect 723 1542 767 1546
rect 771 1542 831 1546
rect 835 1542 911 1546
rect 915 1542 943 1546
rect 947 1542 1047 1546
rect 1051 1542 1055 1546
rect 1059 1542 1167 1546
rect 1171 1542 1175 1546
rect 1179 1542 1279 1546
rect 1283 1542 1311 1546
rect 1315 1542 1447 1546
rect 1451 1542 1767 1546
rect 1771 1542 1791 1546
rect 103 1541 1791 1542
rect 1797 1546 1807 1547
rect 1811 1546 1919 1550
rect 1923 1546 2039 1550
rect 2043 1546 2063 1550
rect 2067 1546 2159 1550
rect 2163 1546 2167 1550
rect 2171 1546 2255 1550
rect 2259 1546 2295 1550
rect 2299 1546 2359 1550
rect 2363 1546 2423 1550
rect 2427 1546 2463 1550
rect 2467 1546 2551 1550
rect 2555 1546 2567 1550
rect 2571 1546 2671 1550
rect 2675 1546 2679 1550
rect 2683 1546 2775 1550
rect 2779 1546 2799 1550
rect 2803 1546 2887 1550
rect 2891 1546 2927 1550
rect 2931 1546 3055 1550
rect 3059 1546 3463 1550
rect 3467 1546 3506 1550
rect 1797 1545 3506 1546
rect 1797 1541 1798 1545
rect 84 1473 85 1479
rect 91 1478 1779 1479
rect 91 1474 111 1478
rect 115 1474 159 1478
rect 163 1474 183 1478
rect 187 1474 327 1478
rect 331 1474 375 1478
rect 379 1474 471 1478
rect 475 1474 583 1478
rect 587 1474 623 1478
rect 627 1474 767 1478
rect 771 1474 783 1478
rect 787 1474 911 1478
rect 915 1474 959 1478
rect 963 1474 1047 1478
rect 1051 1474 1127 1478
rect 1131 1474 1175 1478
rect 1179 1474 1279 1478
rect 1283 1474 1311 1478
rect 1315 1474 1431 1478
rect 1435 1474 1447 1478
rect 1451 1474 1591 1478
rect 1595 1474 1767 1478
rect 1771 1474 1779 1478
rect 91 1473 1779 1474
rect 1785 1478 3494 1479
rect 1785 1474 1807 1478
rect 1811 1474 1831 1478
rect 1835 1474 1919 1478
rect 1923 1474 1951 1478
rect 1955 1474 2039 1478
rect 2043 1474 2111 1478
rect 2115 1474 2167 1478
rect 2171 1474 2271 1478
rect 2275 1474 2295 1478
rect 2299 1474 2423 1478
rect 2427 1474 2431 1478
rect 2435 1474 2551 1478
rect 2555 1474 2591 1478
rect 2595 1474 2679 1478
rect 2683 1474 2735 1478
rect 2739 1474 2799 1478
rect 2803 1474 2871 1478
rect 2875 1474 2927 1478
rect 2931 1474 3007 1478
rect 3011 1474 3055 1478
rect 3059 1474 3135 1478
rect 3139 1474 3263 1478
rect 3267 1474 3367 1478
rect 3371 1474 3463 1478
rect 3467 1474 3494 1478
rect 1785 1473 3494 1474
rect 96 1405 97 1411
rect 103 1410 1791 1411
rect 103 1406 111 1410
rect 115 1406 135 1410
rect 139 1406 159 1410
rect 163 1406 303 1410
rect 307 1406 375 1410
rect 379 1406 495 1410
rect 499 1406 583 1410
rect 587 1406 679 1410
rect 683 1406 783 1410
rect 787 1406 855 1410
rect 859 1406 959 1410
rect 963 1406 1015 1410
rect 1019 1406 1127 1410
rect 1131 1406 1167 1410
rect 1171 1406 1279 1410
rect 1283 1406 1303 1410
rect 1307 1406 1431 1410
rect 1435 1406 1559 1410
rect 1563 1406 1591 1410
rect 1595 1406 1671 1410
rect 1675 1406 1767 1410
rect 1771 1406 1791 1410
rect 103 1405 1791 1406
rect 1797 1410 3506 1411
rect 1797 1406 1807 1410
rect 1811 1406 1831 1410
rect 1835 1406 1951 1410
rect 1955 1406 2007 1410
rect 2011 1406 2111 1410
rect 2115 1406 2199 1410
rect 2203 1406 2271 1410
rect 2275 1406 2383 1410
rect 2387 1406 2431 1410
rect 2435 1406 2559 1410
rect 2563 1406 2591 1410
rect 2595 1406 2719 1410
rect 2723 1406 2735 1410
rect 2739 1406 2863 1410
rect 2867 1406 2871 1410
rect 2875 1406 2999 1410
rect 3003 1406 3007 1410
rect 3011 1406 3127 1410
rect 3131 1406 3135 1410
rect 3139 1406 3255 1410
rect 3259 1406 3263 1410
rect 3267 1406 3367 1410
rect 3371 1406 3463 1410
rect 3467 1406 3506 1410
rect 1797 1405 3506 1406
rect 84 1337 85 1343
rect 91 1342 1779 1343
rect 91 1338 111 1342
rect 115 1338 135 1342
rect 139 1338 247 1342
rect 251 1338 303 1342
rect 307 1338 399 1342
rect 403 1338 495 1342
rect 499 1338 559 1342
rect 563 1338 679 1342
rect 683 1338 727 1342
rect 731 1338 855 1342
rect 859 1338 895 1342
rect 899 1338 1015 1342
rect 1019 1338 1063 1342
rect 1067 1338 1167 1342
rect 1171 1338 1223 1342
rect 1227 1338 1303 1342
rect 1307 1338 1375 1342
rect 1379 1338 1431 1342
rect 1435 1338 1535 1342
rect 1539 1338 1559 1342
rect 1563 1338 1671 1342
rect 1675 1338 1767 1342
rect 1771 1338 1779 1342
rect 91 1337 1779 1338
rect 1785 1339 1786 1343
rect 1785 1338 3494 1339
rect 1785 1337 1807 1338
rect 1778 1334 1807 1337
rect 1811 1334 1831 1338
rect 1835 1334 1967 1338
rect 1971 1334 2007 1338
rect 2011 1334 2143 1338
rect 2147 1334 2199 1338
rect 2203 1334 2327 1338
rect 2331 1334 2383 1338
rect 2387 1334 2511 1338
rect 2515 1334 2559 1338
rect 2563 1334 2687 1338
rect 2691 1334 2719 1338
rect 2723 1334 2863 1338
rect 2867 1334 2999 1338
rect 3003 1334 3039 1338
rect 3043 1334 3127 1338
rect 3131 1334 3215 1338
rect 3219 1334 3255 1338
rect 3259 1334 3367 1338
rect 3371 1334 3463 1338
rect 3467 1334 3494 1338
rect 1778 1333 3494 1334
rect 186 1284 192 1285
rect 498 1284 504 1285
rect 186 1280 187 1284
rect 191 1280 499 1284
rect 503 1280 504 1284
rect 186 1279 192 1280
rect 498 1279 504 1280
rect 96 1269 97 1275
rect 103 1274 1791 1275
rect 103 1270 111 1274
rect 115 1270 135 1274
rect 139 1270 223 1274
rect 227 1270 247 1274
rect 251 1270 319 1274
rect 323 1270 399 1274
rect 403 1270 431 1274
rect 435 1270 551 1274
rect 555 1270 559 1274
rect 563 1270 679 1274
rect 683 1270 727 1274
rect 731 1270 823 1274
rect 827 1270 895 1274
rect 899 1270 975 1274
rect 979 1270 1063 1274
rect 1067 1270 1143 1274
rect 1147 1270 1223 1274
rect 1227 1270 1319 1274
rect 1323 1270 1375 1274
rect 1379 1270 1503 1274
rect 1507 1270 1535 1274
rect 1539 1270 1671 1274
rect 1675 1270 1767 1274
rect 1771 1270 1791 1274
rect 103 1269 1791 1270
rect 1797 1274 3506 1275
rect 1797 1270 1807 1274
rect 1811 1270 1831 1274
rect 1835 1270 1967 1274
rect 1971 1270 2095 1274
rect 2099 1270 2143 1274
rect 2147 1270 2327 1274
rect 2331 1270 2359 1274
rect 2363 1270 2511 1274
rect 2515 1270 2599 1274
rect 2603 1270 2687 1274
rect 2691 1270 2807 1274
rect 2811 1270 2863 1274
rect 2867 1270 3007 1274
rect 3011 1270 3039 1274
rect 3043 1270 3199 1274
rect 3203 1270 3215 1274
rect 3219 1270 3367 1274
rect 3371 1270 3463 1274
rect 3467 1270 3506 1274
rect 1797 1269 3506 1270
rect 84 1197 85 1203
rect 91 1202 1779 1203
rect 91 1198 111 1202
rect 115 1198 135 1202
rect 139 1198 223 1202
rect 227 1198 231 1202
rect 235 1198 319 1202
rect 323 1198 359 1202
rect 363 1198 431 1202
rect 435 1198 487 1202
rect 491 1198 551 1202
rect 555 1198 615 1202
rect 619 1198 679 1202
rect 683 1198 743 1202
rect 747 1198 823 1202
rect 827 1198 871 1202
rect 875 1198 975 1202
rect 979 1198 991 1202
rect 995 1198 1119 1202
rect 1123 1198 1143 1202
rect 1147 1198 1247 1202
rect 1251 1198 1319 1202
rect 1323 1198 1503 1202
rect 1507 1198 1671 1202
rect 1675 1198 1767 1202
rect 1771 1198 1779 1202
rect 91 1197 1779 1198
rect 1785 1202 3494 1203
rect 1785 1198 1807 1202
rect 1811 1198 1831 1202
rect 1835 1198 1935 1202
rect 1939 1198 2039 1202
rect 2043 1198 2095 1202
rect 2099 1198 2159 1202
rect 2163 1198 2287 1202
rect 2291 1198 2359 1202
rect 2363 1198 2423 1202
rect 2427 1198 2567 1202
rect 2571 1198 2599 1202
rect 2603 1198 2703 1202
rect 2707 1198 2807 1202
rect 2811 1198 2839 1202
rect 2843 1198 2975 1202
rect 2979 1198 3007 1202
rect 3011 1198 3111 1202
rect 3115 1198 3199 1202
rect 3203 1198 3247 1202
rect 3251 1198 3367 1202
rect 3371 1198 3463 1202
rect 3467 1198 3494 1202
rect 1785 1197 3494 1198
rect 96 1129 97 1135
rect 103 1134 1791 1135
rect 103 1130 111 1134
rect 115 1130 135 1134
rect 139 1130 231 1134
rect 235 1130 247 1134
rect 251 1130 359 1134
rect 363 1130 367 1134
rect 371 1130 487 1134
rect 491 1130 495 1134
rect 499 1130 615 1134
rect 619 1130 623 1134
rect 627 1130 743 1134
rect 747 1130 759 1134
rect 763 1130 871 1134
rect 875 1130 887 1134
rect 891 1130 991 1134
rect 995 1130 1015 1134
rect 1019 1130 1119 1134
rect 1123 1130 1143 1134
rect 1147 1130 1247 1134
rect 1251 1130 1271 1134
rect 1275 1130 1399 1134
rect 1403 1130 1767 1134
rect 1771 1130 1791 1134
rect 103 1129 1791 1130
rect 1797 1131 1798 1135
rect 1797 1130 3506 1131
rect 1797 1129 1807 1130
rect 1790 1126 1807 1129
rect 1811 1126 1935 1130
rect 1939 1126 1943 1130
rect 1947 1126 2039 1130
rect 2043 1126 2063 1130
rect 2067 1126 2159 1130
rect 2163 1126 2191 1130
rect 2195 1126 2287 1130
rect 2291 1126 2319 1130
rect 2323 1126 2423 1130
rect 2427 1126 2455 1130
rect 2459 1126 2567 1130
rect 2571 1126 2599 1130
rect 2603 1126 2703 1130
rect 2707 1126 2751 1130
rect 2755 1126 2839 1130
rect 2843 1126 2903 1130
rect 2907 1126 2975 1130
rect 2979 1126 3063 1130
rect 3067 1126 3111 1130
rect 3115 1126 3223 1130
rect 3227 1126 3247 1130
rect 3251 1126 3367 1130
rect 3371 1126 3463 1130
rect 3467 1126 3506 1130
rect 1790 1125 3506 1126
rect 84 1061 85 1067
rect 91 1066 1779 1067
rect 91 1062 111 1066
rect 115 1062 247 1066
rect 251 1062 367 1066
rect 371 1062 431 1066
rect 435 1062 495 1066
rect 499 1062 543 1066
rect 547 1062 623 1066
rect 627 1062 663 1066
rect 667 1062 759 1066
rect 763 1062 791 1066
rect 795 1062 887 1066
rect 891 1062 919 1066
rect 923 1062 1015 1066
rect 1019 1062 1039 1066
rect 1043 1062 1143 1066
rect 1147 1062 1159 1066
rect 1163 1062 1271 1066
rect 1275 1062 1279 1066
rect 1283 1062 1399 1066
rect 1403 1062 1407 1066
rect 1411 1062 1535 1066
rect 1539 1062 1767 1066
rect 1771 1062 1779 1066
rect 91 1061 1779 1062
rect 1785 1063 1786 1067
rect 1785 1062 3494 1063
rect 1785 1061 1807 1062
rect 1778 1058 1807 1061
rect 1811 1058 1847 1062
rect 1851 1058 1943 1062
rect 1947 1058 1983 1062
rect 1987 1058 2063 1062
rect 2067 1058 2119 1062
rect 2123 1058 2191 1062
rect 2195 1058 2255 1062
rect 2259 1058 2319 1062
rect 2323 1058 2391 1062
rect 2395 1058 2455 1062
rect 2459 1058 2543 1062
rect 2547 1058 2599 1062
rect 2603 1058 2703 1062
rect 2707 1058 2751 1062
rect 2755 1058 2863 1062
rect 2867 1058 2903 1062
rect 2907 1058 3031 1062
rect 3035 1058 3063 1062
rect 3067 1058 3207 1062
rect 3211 1058 3223 1062
rect 3227 1058 3367 1062
rect 3371 1058 3463 1062
rect 3467 1058 3494 1062
rect 1778 1057 3494 1058
rect 96 989 97 995
rect 103 994 1791 995
rect 103 990 111 994
rect 115 990 431 994
rect 435 990 543 994
rect 547 990 567 994
rect 571 990 663 994
rect 667 990 679 994
rect 683 990 791 994
rect 795 990 911 994
rect 915 990 919 994
rect 923 990 1031 994
rect 1035 990 1039 994
rect 1043 990 1143 994
rect 1147 990 1159 994
rect 1163 990 1255 994
rect 1259 990 1279 994
rect 1283 990 1359 994
rect 1363 990 1407 994
rect 1411 990 1471 994
rect 1475 990 1535 994
rect 1539 990 1583 994
rect 1587 990 1671 994
rect 1675 990 1767 994
rect 1771 990 1791 994
rect 103 989 1791 990
rect 1797 994 3506 995
rect 1797 990 1807 994
rect 1811 990 1831 994
rect 1835 990 1847 994
rect 1851 990 1975 994
rect 1979 990 1983 994
rect 1987 990 2119 994
rect 2123 990 2135 994
rect 2139 990 2255 994
rect 2259 990 2295 994
rect 2299 990 2391 994
rect 2395 990 2463 994
rect 2467 990 2543 994
rect 2547 990 2631 994
rect 2635 990 2703 994
rect 2707 990 2807 994
rect 2811 990 2863 994
rect 2867 990 2991 994
rect 2995 990 3031 994
rect 3035 990 3183 994
rect 3187 990 3207 994
rect 3211 990 3367 994
rect 3371 990 3463 994
rect 3467 990 3506 994
rect 1797 989 3506 990
rect 1778 930 3494 931
rect 1778 927 1807 930
rect 84 921 85 927
rect 91 926 1779 927
rect 91 922 111 926
rect 115 922 415 926
rect 419 922 559 926
rect 563 922 567 926
rect 571 922 679 926
rect 683 922 727 926
rect 731 922 791 926
rect 795 922 911 926
rect 915 922 1031 926
rect 1035 922 1119 926
rect 1123 922 1143 926
rect 1147 922 1255 926
rect 1259 922 1335 926
rect 1339 922 1359 926
rect 1363 922 1471 926
rect 1475 922 1559 926
rect 1563 922 1583 926
rect 1587 922 1671 926
rect 1675 922 1767 926
rect 1771 922 1779 926
rect 91 921 1779 922
rect 1785 926 1807 927
rect 1811 926 1831 930
rect 1835 926 1975 930
rect 1979 926 2127 930
rect 2131 926 2135 930
rect 2139 926 2215 930
rect 2219 926 2295 930
rect 2299 926 2303 930
rect 2307 926 2391 930
rect 2395 926 2463 930
rect 2467 926 2479 930
rect 2483 926 2567 930
rect 2571 926 2631 930
rect 2635 926 2655 930
rect 2659 926 2743 930
rect 2747 926 2807 930
rect 2811 926 2831 930
rect 2835 926 2991 930
rect 2995 926 3183 930
rect 3187 926 3367 930
rect 3371 926 3463 930
rect 3467 926 3494 930
rect 1785 925 3494 926
rect 1785 921 1786 925
rect 96 853 97 859
rect 103 858 1791 859
rect 103 854 111 858
rect 115 854 135 858
rect 139 854 231 858
rect 235 854 359 858
rect 363 854 415 858
rect 419 854 487 858
rect 491 854 559 858
rect 563 854 623 858
rect 627 854 727 858
rect 731 854 751 858
rect 755 854 879 858
rect 883 854 911 858
rect 915 854 1007 858
rect 1011 854 1119 858
rect 1123 854 1135 858
rect 1139 854 1271 858
rect 1275 854 1335 858
rect 1339 854 1559 858
rect 1563 854 1767 858
rect 1771 854 1791 858
rect 103 853 1791 854
rect 1797 858 3506 859
rect 1797 854 1807 858
rect 1811 854 2127 858
rect 2131 854 2159 858
rect 2163 854 2215 858
rect 2219 854 2247 858
rect 2251 854 2303 858
rect 2307 854 2335 858
rect 2339 854 2391 858
rect 2395 854 2423 858
rect 2427 854 2479 858
rect 2483 854 2527 858
rect 2531 854 2567 858
rect 2571 854 2639 858
rect 2643 854 2655 858
rect 2659 854 2743 858
rect 2747 854 2767 858
rect 2771 854 2831 858
rect 2835 854 2911 858
rect 2915 854 3063 858
rect 3067 854 3223 858
rect 3227 854 3367 858
rect 3371 854 3463 858
rect 3467 854 3506 858
rect 1797 853 3506 854
rect 84 785 85 791
rect 91 790 1779 791
rect 91 786 111 790
rect 115 786 135 790
rect 139 786 223 790
rect 227 786 231 790
rect 235 786 343 790
rect 347 786 359 790
rect 363 786 471 790
rect 475 786 487 790
rect 491 786 607 790
rect 611 786 623 790
rect 627 786 743 790
rect 747 786 751 790
rect 755 786 879 790
rect 883 786 887 790
rect 891 786 1007 790
rect 1011 786 1039 790
rect 1043 786 1135 790
rect 1139 786 1191 790
rect 1195 786 1271 790
rect 1275 786 1351 790
rect 1355 786 1767 790
rect 1771 786 1779 790
rect 91 785 1779 786
rect 1785 790 3494 791
rect 1785 786 1807 790
rect 1811 786 2063 790
rect 2067 786 2159 790
rect 2163 786 2175 790
rect 2179 786 2247 790
rect 2251 786 2295 790
rect 2299 786 2335 790
rect 2339 786 2423 790
rect 2427 786 2527 790
rect 2531 786 2559 790
rect 2563 786 2639 790
rect 2643 786 2711 790
rect 2715 786 2767 790
rect 2771 786 2871 790
rect 2875 786 2911 790
rect 2915 786 3039 790
rect 3043 786 3063 790
rect 3067 786 3215 790
rect 3219 786 3223 790
rect 3227 786 3367 790
rect 3371 786 3463 790
rect 3467 786 3494 790
rect 1785 785 3494 786
rect 1790 726 3506 727
rect 1790 723 1807 726
rect 96 717 97 723
rect 103 722 1791 723
rect 103 718 111 722
rect 115 718 135 722
rect 139 718 167 722
rect 171 718 223 722
rect 227 718 295 722
rect 299 718 343 722
rect 347 718 431 722
rect 435 718 471 722
rect 475 718 575 722
rect 579 718 607 722
rect 611 718 727 722
rect 731 718 743 722
rect 747 718 879 722
rect 883 718 887 722
rect 891 718 1031 722
rect 1035 718 1039 722
rect 1043 718 1183 722
rect 1187 718 1191 722
rect 1195 718 1343 722
rect 1347 718 1351 722
rect 1355 718 1503 722
rect 1507 718 1767 722
rect 1771 718 1791 722
rect 103 717 1791 718
rect 1797 722 1807 723
rect 1811 722 1927 726
rect 1931 722 2063 726
rect 2067 722 2071 726
rect 2075 722 2175 726
rect 2179 722 2231 726
rect 2235 722 2295 726
rect 2299 722 2391 726
rect 2395 722 2423 726
rect 2427 722 2551 726
rect 2555 722 2559 726
rect 2563 722 2703 726
rect 2707 722 2711 726
rect 2715 722 2847 726
rect 2851 722 2871 726
rect 2875 722 2983 726
rect 2987 722 3039 726
rect 3043 722 3119 726
rect 3123 722 3215 726
rect 3219 722 3255 726
rect 3259 722 3367 726
rect 3371 722 3463 726
rect 3467 722 3506 726
rect 1797 721 3506 722
rect 1797 717 1798 721
rect 84 649 85 655
rect 91 654 1779 655
rect 91 650 111 654
rect 115 650 167 654
rect 171 650 295 654
rect 299 650 431 654
rect 435 650 455 654
rect 459 650 559 654
rect 563 650 575 654
rect 579 650 679 654
rect 683 650 727 654
rect 731 650 799 654
rect 803 650 879 654
rect 883 650 927 654
rect 931 650 1031 654
rect 1035 650 1055 654
rect 1059 650 1183 654
rect 1187 650 1311 654
rect 1315 650 1343 654
rect 1347 650 1447 654
rect 1451 650 1503 654
rect 1507 650 1583 654
rect 1587 650 1767 654
rect 1771 650 1779 654
rect 91 649 1779 650
rect 1785 654 3494 655
rect 1785 650 1807 654
rect 1811 650 1831 654
rect 1835 650 1927 654
rect 1931 650 1967 654
rect 1971 650 2071 654
rect 2075 650 2135 654
rect 2139 650 2231 654
rect 2235 650 2311 654
rect 2315 650 2391 654
rect 2395 650 2487 654
rect 2491 650 2551 654
rect 2555 650 2655 654
rect 2659 650 2703 654
rect 2707 650 2815 654
rect 2819 650 2847 654
rect 2851 650 2959 654
rect 2963 650 2983 654
rect 2987 650 3103 654
rect 3107 650 3119 654
rect 3123 650 3247 654
rect 3251 650 3255 654
rect 3259 650 3367 654
rect 3371 650 3463 654
rect 3467 650 3494 654
rect 1785 649 3494 650
rect 1790 585 1791 591
rect 1797 590 3499 591
rect 1797 586 1807 590
rect 1811 586 1831 590
rect 1835 586 1967 590
rect 1971 586 2127 590
rect 2131 586 2135 590
rect 2139 586 2287 590
rect 2291 586 2311 590
rect 2315 586 2455 590
rect 2459 586 2487 590
rect 2491 586 2623 590
rect 2627 586 2655 590
rect 2659 586 2799 590
rect 2803 586 2815 590
rect 2819 586 2959 590
rect 2963 586 2983 590
rect 2987 586 3103 590
rect 3107 586 3167 590
rect 3171 586 3247 590
rect 3251 586 3359 590
rect 3363 586 3367 590
rect 3371 586 3463 590
rect 3467 586 3499 590
rect 1797 585 3499 586
rect 3505 585 3506 591
rect 1790 583 1798 585
rect 96 577 97 583
rect 103 582 1791 583
rect 103 578 111 582
rect 115 578 455 582
rect 459 578 559 582
rect 563 578 599 582
rect 603 578 679 582
rect 683 578 703 582
rect 707 578 799 582
rect 803 578 815 582
rect 819 578 927 582
rect 931 578 1039 582
rect 1043 578 1055 582
rect 1059 578 1151 582
rect 1155 578 1183 582
rect 1187 578 1255 582
rect 1259 578 1311 582
rect 1315 578 1359 582
rect 1363 578 1447 582
rect 1451 578 1471 582
rect 1475 578 1583 582
rect 1587 578 1671 582
rect 1675 578 1767 582
rect 1771 578 1791 582
rect 103 577 1791 578
rect 1797 577 1798 583
rect 84 513 85 519
rect 91 518 1779 519
rect 91 514 111 518
rect 115 514 303 518
rect 307 514 431 518
rect 435 514 567 518
rect 571 514 599 518
rect 603 514 703 518
rect 707 514 815 518
rect 819 514 847 518
rect 851 514 927 518
rect 931 514 983 518
rect 987 514 1039 518
rect 1043 514 1111 518
rect 1115 514 1151 518
rect 1155 514 1231 518
rect 1235 514 1255 518
rect 1259 514 1351 518
rect 1355 514 1359 518
rect 1363 514 1463 518
rect 1467 514 1471 518
rect 1475 514 1575 518
rect 1579 514 1583 518
rect 1587 514 1671 518
rect 1675 514 1767 518
rect 1771 514 1779 518
rect 91 513 1779 514
rect 1785 513 1786 519
rect 1778 511 1786 513
rect 1778 505 1779 511
rect 1785 510 3487 511
rect 1785 506 1807 510
rect 1811 506 1831 510
rect 1835 506 1967 510
rect 1971 506 2127 510
rect 2131 506 2287 510
rect 2291 506 2295 510
rect 2299 506 2455 510
rect 2459 506 2479 510
rect 2483 506 2623 510
rect 2627 506 2679 510
rect 2683 506 2799 510
rect 2803 506 2887 510
rect 2891 506 2983 510
rect 2987 506 3111 510
rect 3115 506 3167 510
rect 3171 506 3335 510
rect 3339 506 3359 510
rect 3363 506 3463 510
rect 3467 506 3487 510
rect 1785 505 3487 506
rect 3493 505 3494 511
rect 96 441 97 447
rect 103 446 1791 447
rect 103 442 111 446
rect 115 442 135 446
rect 139 442 255 446
rect 259 442 303 446
rect 307 442 415 446
rect 419 442 431 446
rect 435 442 567 446
rect 571 442 583 446
rect 587 442 703 446
rect 707 442 743 446
rect 747 442 847 446
rect 851 442 903 446
rect 907 442 983 446
rect 987 442 1047 446
rect 1051 442 1111 446
rect 1115 442 1183 446
rect 1187 442 1231 446
rect 1235 442 1311 446
rect 1315 442 1351 446
rect 1355 442 1439 446
rect 1443 442 1463 446
rect 1467 442 1567 446
rect 1571 442 1575 446
rect 1579 442 1671 446
rect 1675 442 1767 446
rect 1771 442 1791 446
rect 103 441 1791 442
rect 1797 446 3506 447
rect 1797 442 1807 446
rect 1811 442 1831 446
rect 1835 442 1959 446
rect 1963 442 1967 446
rect 1971 442 2111 446
rect 2115 442 2127 446
rect 2131 442 2271 446
rect 2275 442 2295 446
rect 2299 442 2455 446
rect 2459 442 2479 446
rect 2483 442 2655 446
rect 2659 442 2679 446
rect 2683 442 2871 446
rect 2875 442 2887 446
rect 2891 442 3103 446
rect 3107 442 3111 446
rect 3115 442 3335 446
rect 3339 442 3463 446
rect 3467 442 3506 446
rect 1797 441 3506 442
rect 84 373 85 379
rect 91 378 1779 379
rect 91 374 111 378
rect 115 374 135 378
rect 139 374 223 378
rect 227 374 255 378
rect 259 374 343 378
rect 347 374 415 378
rect 419 374 471 378
rect 475 374 583 378
rect 587 374 599 378
rect 603 374 719 378
rect 723 374 743 378
rect 747 374 839 378
rect 843 374 903 378
rect 907 374 959 378
rect 963 374 1047 378
rect 1051 374 1079 378
rect 1083 374 1183 378
rect 1187 374 1207 378
rect 1211 374 1311 378
rect 1315 374 1439 378
rect 1443 374 1567 378
rect 1571 374 1671 378
rect 1675 374 1767 378
rect 1771 374 1779 378
rect 91 373 1779 374
rect 1785 378 3494 379
rect 1785 374 1807 378
rect 1811 374 1831 378
rect 1835 374 1927 378
rect 1931 374 1959 378
rect 1963 374 2039 378
rect 2043 374 2111 378
rect 2115 374 2159 378
rect 2163 374 2271 378
rect 2275 374 2287 378
rect 2291 374 2423 378
rect 2427 374 2455 378
rect 2459 374 2583 378
rect 2587 374 2655 378
rect 2659 374 2759 378
rect 2763 374 2871 378
rect 2875 374 2951 378
rect 2955 374 3103 378
rect 3107 374 3151 378
rect 3155 374 3335 378
rect 3339 374 3359 378
rect 3363 374 3463 378
rect 3467 374 3494 378
rect 1785 373 3494 374
rect 1790 314 3506 315
rect 1790 311 1807 314
rect 96 305 97 311
rect 103 310 1791 311
rect 103 306 111 310
rect 115 306 135 310
rect 139 306 223 310
rect 227 306 263 310
rect 267 306 343 310
rect 347 306 375 310
rect 379 306 471 310
rect 475 306 487 310
rect 491 306 599 310
rect 603 306 711 310
rect 715 306 719 310
rect 723 306 815 310
rect 819 306 839 310
rect 843 306 919 310
rect 923 306 959 310
rect 963 306 1023 310
rect 1027 306 1079 310
rect 1083 306 1127 310
rect 1131 306 1207 310
rect 1211 306 1239 310
rect 1243 306 1767 310
rect 1771 306 1791 310
rect 103 305 1791 306
rect 1797 310 1807 311
rect 1811 310 1927 314
rect 1931 310 2039 314
rect 2043 310 2159 314
rect 2163 310 2223 314
rect 2227 310 2287 314
rect 2291 310 2311 314
rect 2315 310 2399 314
rect 2403 310 2423 314
rect 2427 310 2487 314
rect 2491 310 2575 314
rect 2579 310 2583 314
rect 2587 310 2679 314
rect 2683 310 2759 314
rect 2763 310 2799 314
rect 2803 310 2927 314
rect 2931 310 2951 314
rect 2955 310 3071 314
rect 3075 310 3151 314
rect 3155 310 3223 314
rect 3227 310 3359 314
rect 3363 310 3367 314
rect 3371 310 3463 314
rect 3467 310 3506 314
rect 1797 309 3506 310
rect 1797 305 1798 309
rect 84 237 85 243
rect 91 242 1779 243
rect 91 238 111 242
rect 115 238 263 242
rect 267 238 375 242
rect 379 238 447 242
rect 451 238 487 242
rect 491 238 535 242
rect 539 238 599 242
rect 603 238 623 242
rect 627 238 711 242
rect 715 238 807 242
rect 811 238 815 242
rect 819 238 903 242
rect 907 238 919 242
rect 923 238 999 242
rect 1003 238 1023 242
rect 1027 238 1103 242
rect 1107 238 1127 242
rect 1131 238 1207 242
rect 1211 238 1239 242
rect 1243 238 1311 242
rect 1315 238 1767 242
rect 1771 238 1779 242
rect 91 237 1779 238
rect 1785 242 3494 243
rect 1785 238 1807 242
rect 1811 238 2143 242
rect 2147 238 2223 242
rect 2227 238 2263 242
rect 2267 238 2311 242
rect 2315 238 2383 242
rect 2387 238 2399 242
rect 2403 238 2487 242
rect 2491 238 2511 242
rect 2515 238 2575 242
rect 2579 238 2639 242
rect 2643 238 2679 242
rect 2683 238 2767 242
rect 2771 238 2799 242
rect 2803 238 2895 242
rect 2899 238 2927 242
rect 2931 238 3015 242
rect 3019 238 3071 242
rect 3075 238 3135 242
rect 3139 238 3223 242
rect 3227 238 3263 242
rect 3267 238 3367 242
rect 3371 238 3463 242
rect 3467 238 3494 242
rect 1785 237 3494 238
rect 1790 154 3506 155
rect 1790 151 1807 154
rect 96 145 97 151
rect 103 150 1791 151
rect 103 146 111 150
rect 115 146 263 150
rect 267 146 351 150
rect 355 146 439 150
rect 443 146 447 150
rect 451 146 527 150
rect 531 146 535 150
rect 539 146 615 150
rect 619 146 623 150
rect 627 146 703 150
rect 707 146 711 150
rect 715 146 791 150
rect 795 146 807 150
rect 811 146 879 150
rect 883 146 903 150
rect 907 146 967 150
rect 971 146 999 150
rect 1003 146 1055 150
rect 1059 146 1103 150
rect 1107 146 1143 150
rect 1147 146 1207 150
rect 1211 146 1231 150
rect 1235 146 1311 150
rect 1315 146 1319 150
rect 1323 146 1407 150
rect 1411 146 1495 150
rect 1499 146 1583 150
rect 1587 146 1671 150
rect 1675 146 1767 150
rect 1771 146 1791 150
rect 103 145 1791 146
rect 1797 150 1807 151
rect 1811 150 1831 154
rect 1835 150 1919 154
rect 1923 150 2007 154
rect 2011 150 2095 154
rect 2099 150 2143 154
rect 2147 150 2183 154
rect 2187 150 2263 154
rect 2267 150 2295 154
rect 2299 150 2383 154
rect 2387 150 2407 154
rect 2411 150 2511 154
rect 2515 150 2615 154
rect 2619 150 2639 154
rect 2643 150 2719 154
rect 2723 150 2767 154
rect 2771 150 2815 154
rect 2819 150 2895 154
rect 2899 150 2911 154
rect 2915 150 3007 154
rect 3011 150 3015 154
rect 3019 150 3103 154
rect 3107 150 3135 154
rect 3139 150 3191 154
rect 3195 150 3263 154
rect 3267 150 3279 154
rect 3283 150 3367 154
rect 3371 150 3463 154
rect 3467 150 3506 154
rect 1797 149 3506 150
rect 1797 145 1798 149
rect 1778 90 3494 91
rect 1778 87 1807 90
rect 84 81 85 87
rect 91 86 1779 87
rect 91 82 111 86
rect 115 82 263 86
rect 267 82 351 86
rect 355 82 439 86
rect 443 82 527 86
rect 531 82 615 86
rect 619 82 703 86
rect 707 82 791 86
rect 795 82 879 86
rect 883 82 967 86
rect 971 82 1055 86
rect 1059 82 1143 86
rect 1147 82 1231 86
rect 1235 82 1319 86
rect 1323 82 1407 86
rect 1411 82 1495 86
rect 1499 82 1583 86
rect 1587 82 1671 86
rect 1675 82 1767 86
rect 1771 82 1779 86
rect 91 81 1779 82
rect 1785 86 1807 87
rect 1811 86 1831 90
rect 1835 86 1919 90
rect 1923 86 2007 90
rect 2011 86 2095 90
rect 2099 86 2183 90
rect 2187 86 2295 90
rect 2299 86 2407 90
rect 2411 86 2511 90
rect 2515 86 2615 90
rect 2619 86 2719 90
rect 2723 86 2815 90
rect 2819 86 2911 90
rect 2915 86 3007 90
rect 3011 86 3103 90
rect 3107 86 3191 90
rect 3195 86 3279 90
rect 3283 86 3367 90
rect 3371 86 3463 90
rect 3467 86 3494 90
rect 1785 85 3494 86
rect 1785 81 1786 85
<< m5c >>
rect 97 3501 103 3507
rect 1791 3501 1797 3507
rect 1791 3489 1797 3495
rect 3499 3489 3505 3495
rect 85 3433 91 3439
rect 1779 3433 1785 3439
rect 1779 3425 1785 3431
rect 3487 3425 3493 3431
rect 97 3361 103 3367
rect 1791 3361 1797 3367
rect 85 3289 91 3295
rect 1779 3289 1785 3295
rect 1791 3225 1797 3231
rect 3499 3225 3505 3231
rect 97 3217 103 3223
rect 1791 3217 1797 3223
rect 1779 3161 1785 3167
rect 3487 3161 3493 3167
rect 85 3153 91 3159
rect 1779 3153 1785 3159
rect 97 3085 103 3091
rect 1791 3085 1797 3091
rect 85 3013 91 3019
rect 1779 3013 1785 3019
rect 97 2937 103 2943
rect 1791 2937 1797 2943
rect 85 2865 91 2871
rect 1779 2865 1785 2871
rect 1791 2801 1797 2807
rect 3499 2801 3505 2807
rect 97 2789 103 2795
rect 1791 2789 1797 2795
rect 85 2717 91 2723
rect 1779 2717 1785 2723
rect 97 2645 103 2651
rect 1791 2645 1797 2651
rect 85 2573 91 2579
rect 1779 2573 1785 2579
rect 97 2501 103 2507
rect 1791 2501 1797 2507
rect 85 2437 91 2443
rect 1779 2437 1785 2443
rect 97 2369 103 2375
rect 1791 2369 1797 2375
rect 85 2297 91 2303
rect 1779 2297 1785 2303
rect 97 2229 103 2235
rect 1791 2229 1797 2235
rect 1779 2169 1785 2175
rect 3487 2169 3493 2175
rect 85 2157 91 2163
rect 1779 2157 1785 2163
rect 1791 2097 1797 2103
rect 3499 2097 3505 2103
rect 97 2089 103 2095
rect 1791 2089 1797 2095
rect 1779 2029 1785 2035
rect 3487 2029 3493 2035
rect 85 2017 91 2023
rect 1779 2017 1785 2023
rect 1791 1961 1797 1967
rect 3499 1961 3505 1967
rect 97 1949 103 1955
rect 1791 1949 1797 1955
rect 1779 1893 1785 1899
rect 3487 1893 3493 1899
rect 85 1885 91 1891
rect 1779 1885 1785 1891
rect 97 1817 103 1823
rect 1791 1817 1797 1823
rect 85 1749 91 1755
rect 1779 1749 1785 1755
rect 97 1681 103 1687
rect 1791 1681 1797 1687
rect 85 1613 91 1619
rect 1779 1613 1785 1619
rect 97 1541 103 1547
rect 1791 1541 1797 1547
rect 85 1473 91 1479
rect 1779 1473 1785 1479
rect 97 1405 103 1411
rect 1791 1405 1797 1411
rect 85 1337 91 1343
rect 1779 1337 1785 1343
rect 97 1269 103 1275
rect 1791 1269 1797 1275
rect 85 1197 91 1203
rect 1779 1197 1785 1203
rect 97 1129 103 1135
rect 1791 1129 1797 1135
rect 85 1061 91 1067
rect 1779 1061 1785 1067
rect 97 989 103 995
rect 1791 989 1797 995
rect 85 921 91 927
rect 1779 921 1785 927
rect 97 853 103 859
rect 1791 853 1797 859
rect 85 785 91 791
rect 1779 785 1785 791
rect 97 717 103 723
rect 1791 717 1797 723
rect 85 649 91 655
rect 1779 649 1785 655
rect 1791 585 1797 591
rect 3499 585 3505 591
rect 97 577 103 583
rect 1791 577 1797 583
rect 85 513 91 519
rect 1779 513 1785 519
rect 1779 505 1785 511
rect 3487 505 3493 511
rect 97 441 103 447
rect 1791 441 1797 447
rect 85 373 91 379
rect 1779 373 1785 379
rect 97 305 103 311
rect 1791 305 1797 311
rect 85 237 91 243
rect 1779 237 1785 243
rect 97 145 103 151
rect 1791 145 1797 151
rect 85 81 91 87
rect 1779 81 1785 87
<< m5 >>
rect 84 3439 92 3528
rect 84 3433 85 3439
rect 91 3433 92 3439
rect 84 3295 92 3433
rect 84 3289 85 3295
rect 91 3289 92 3295
rect 84 3159 92 3289
rect 84 3153 85 3159
rect 91 3153 92 3159
rect 84 3019 92 3153
rect 84 3013 85 3019
rect 91 3013 92 3019
rect 84 2871 92 3013
rect 84 2865 85 2871
rect 91 2865 92 2871
rect 84 2723 92 2865
rect 84 2717 85 2723
rect 91 2717 92 2723
rect 84 2579 92 2717
rect 84 2573 85 2579
rect 91 2573 92 2579
rect 84 2443 92 2573
rect 84 2437 85 2443
rect 91 2437 92 2443
rect 84 2303 92 2437
rect 84 2297 85 2303
rect 91 2297 92 2303
rect 84 2163 92 2297
rect 84 2157 85 2163
rect 91 2157 92 2163
rect 84 2023 92 2157
rect 84 2017 85 2023
rect 91 2017 92 2023
rect 84 1891 92 2017
rect 84 1885 85 1891
rect 91 1885 92 1891
rect 84 1755 92 1885
rect 84 1749 85 1755
rect 91 1749 92 1755
rect 84 1619 92 1749
rect 84 1613 85 1619
rect 91 1613 92 1619
rect 84 1479 92 1613
rect 84 1473 85 1479
rect 91 1473 92 1479
rect 84 1343 92 1473
rect 84 1337 85 1343
rect 91 1337 92 1343
rect 84 1203 92 1337
rect 84 1197 85 1203
rect 91 1197 92 1203
rect 84 1067 92 1197
rect 84 1061 85 1067
rect 91 1061 92 1067
rect 84 927 92 1061
rect 84 921 85 927
rect 91 921 92 927
rect 84 791 92 921
rect 84 785 85 791
rect 91 785 92 791
rect 84 655 92 785
rect 84 649 85 655
rect 91 649 92 655
rect 84 519 92 649
rect 84 513 85 519
rect 91 513 92 519
rect 84 379 92 513
rect 84 373 85 379
rect 91 373 92 379
rect 84 243 92 373
rect 84 237 85 243
rect 91 237 92 243
rect 84 87 92 237
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 3507 104 3528
rect 96 3501 97 3507
rect 103 3501 104 3507
rect 96 3367 104 3501
rect 96 3361 97 3367
rect 103 3361 104 3367
rect 96 3223 104 3361
rect 96 3217 97 3223
rect 103 3217 104 3223
rect 96 3091 104 3217
rect 96 3085 97 3091
rect 103 3085 104 3091
rect 96 2943 104 3085
rect 96 2937 97 2943
rect 103 2937 104 2943
rect 96 2795 104 2937
rect 96 2789 97 2795
rect 103 2789 104 2795
rect 96 2651 104 2789
rect 96 2645 97 2651
rect 103 2645 104 2651
rect 96 2507 104 2645
rect 96 2501 97 2507
rect 103 2501 104 2507
rect 96 2375 104 2501
rect 96 2369 97 2375
rect 103 2369 104 2375
rect 96 2235 104 2369
rect 96 2229 97 2235
rect 103 2229 104 2235
rect 96 2095 104 2229
rect 96 2089 97 2095
rect 103 2089 104 2095
rect 96 1955 104 2089
rect 96 1949 97 1955
rect 103 1949 104 1955
rect 96 1823 104 1949
rect 96 1817 97 1823
rect 103 1817 104 1823
rect 96 1687 104 1817
rect 96 1681 97 1687
rect 103 1681 104 1687
rect 96 1547 104 1681
rect 96 1541 97 1547
rect 103 1541 104 1547
rect 96 1411 104 1541
rect 96 1405 97 1411
rect 103 1405 104 1411
rect 96 1275 104 1405
rect 96 1269 97 1275
rect 103 1269 104 1275
rect 96 1135 104 1269
rect 96 1129 97 1135
rect 103 1129 104 1135
rect 96 995 104 1129
rect 96 989 97 995
rect 103 989 104 995
rect 96 859 104 989
rect 96 853 97 859
rect 103 853 104 859
rect 96 723 104 853
rect 96 717 97 723
rect 103 717 104 723
rect 96 583 104 717
rect 96 577 97 583
rect 103 577 104 583
rect 96 447 104 577
rect 96 441 97 447
rect 103 441 104 447
rect 96 311 104 441
rect 96 305 97 311
rect 103 305 104 311
rect 96 151 104 305
rect 96 145 97 151
rect 103 145 104 151
rect 96 72 104 145
rect 1778 3439 1786 3528
rect 1778 3433 1779 3439
rect 1785 3433 1786 3439
rect 1778 3431 1786 3433
rect 1778 3425 1779 3431
rect 1785 3425 1786 3431
rect 1778 3295 1786 3425
rect 1778 3289 1779 3295
rect 1785 3289 1786 3295
rect 1778 3167 1786 3289
rect 1778 3161 1779 3167
rect 1785 3161 1786 3167
rect 1778 3159 1786 3161
rect 1778 3153 1779 3159
rect 1785 3153 1786 3159
rect 1778 3019 1786 3153
rect 1778 3013 1779 3019
rect 1785 3013 1786 3019
rect 1778 2871 1786 3013
rect 1778 2865 1779 2871
rect 1785 2865 1786 2871
rect 1778 2723 1786 2865
rect 1778 2717 1779 2723
rect 1785 2717 1786 2723
rect 1778 2579 1786 2717
rect 1778 2573 1779 2579
rect 1785 2573 1786 2579
rect 1778 2443 1786 2573
rect 1778 2437 1779 2443
rect 1785 2437 1786 2443
rect 1778 2303 1786 2437
rect 1778 2297 1779 2303
rect 1785 2297 1786 2303
rect 1778 2175 1786 2297
rect 1778 2169 1779 2175
rect 1785 2169 1786 2175
rect 1778 2163 1786 2169
rect 1778 2157 1779 2163
rect 1785 2157 1786 2163
rect 1778 2035 1786 2157
rect 1778 2029 1779 2035
rect 1785 2029 1786 2035
rect 1778 2023 1786 2029
rect 1778 2017 1779 2023
rect 1785 2017 1786 2023
rect 1778 1899 1786 2017
rect 1778 1893 1779 1899
rect 1785 1893 1786 1899
rect 1778 1891 1786 1893
rect 1778 1885 1779 1891
rect 1785 1885 1786 1891
rect 1778 1755 1786 1885
rect 1778 1749 1779 1755
rect 1785 1749 1786 1755
rect 1778 1619 1786 1749
rect 1778 1613 1779 1619
rect 1785 1613 1786 1619
rect 1778 1479 1786 1613
rect 1778 1473 1779 1479
rect 1785 1473 1786 1479
rect 1778 1343 1786 1473
rect 1778 1337 1779 1343
rect 1785 1337 1786 1343
rect 1778 1203 1786 1337
rect 1778 1197 1779 1203
rect 1785 1197 1786 1203
rect 1778 1067 1786 1197
rect 1778 1061 1779 1067
rect 1785 1061 1786 1067
rect 1778 927 1786 1061
rect 1778 921 1779 927
rect 1785 921 1786 927
rect 1778 791 1786 921
rect 1778 785 1779 791
rect 1785 785 1786 791
rect 1778 655 1786 785
rect 1778 649 1779 655
rect 1785 649 1786 655
rect 1778 519 1786 649
rect 1778 513 1779 519
rect 1785 513 1786 519
rect 1778 511 1786 513
rect 1778 505 1779 511
rect 1785 505 1786 511
rect 1778 379 1786 505
rect 1778 373 1779 379
rect 1785 373 1786 379
rect 1778 243 1786 373
rect 1778 237 1779 243
rect 1785 237 1786 243
rect 1778 87 1786 237
rect 1778 81 1779 87
rect 1785 81 1786 87
rect 1778 72 1786 81
rect 1790 3507 1798 3528
rect 1790 3501 1791 3507
rect 1797 3501 1798 3507
rect 1790 3495 1798 3501
rect 1790 3489 1791 3495
rect 1797 3489 1798 3495
rect 1790 3367 1798 3489
rect 1790 3361 1791 3367
rect 1797 3361 1798 3367
rect 1790 3231 1798 3361
rect 1790 3225 1791 3231
rect 1797 3225 1798 3231
rect 1790 3223 1798 3225
rect 1790 3217 1791 3223
rect 1797 3217 1798 3223
rect 1790 3091 1798 3217
rect 1790 3085 1791 3091
rect 1797 3085 1798 3091
rect 1790 2943 1798 3085
rect 1790 2937 1791 2943
rect 1797 2937 1798 2943
rect 1790 2807 1798 2937
rect 1790 2801 1791 2807
rect 1797 2801 1798 2807
rect 1790 2795 1798 2801
rect 1790 2789 1791 2795
rect 1797 2789 1798 2795
rect 1790 2651 1798 2789
rect 1790 2645 1791 2651
rect 1797 2645 1798 2651
rect 1790 2507 1798 2645
rect 1790 2501 1791 2507
rect 1797 2501 1798 2507
rect 1790 2375 1798 2501
rect 1790 2369 1791 2375
rect 1797 2369 1798 2375
rect 1790 2235 1798 2369
rect 1790 2229 1791 2235
rect 1797 2229 1798 2235
rect 1790 2103 1798 2229
rect 1790 2097 1791 2103
rect 1797 2097 1798 2103
rect 1790 2095 1798 2097
rect 1790 2089 1791 2095
rect 1797 2089 1798 2095
rect 1790 1967 1798 2089
rect 1790 1961 1791 1967
rect 1797 1961 1798 1967
rect 1790 1955 1798 1961
rect 1790 1949 1791 1955
rect 1797 1949 1798 1955
rect 1790 1823 1798 1949
rect 1790 1817 1791 1823
rect 1797 1817 1798 1823
rect 1790 1687 1798 1817
rect 1790 1681 1791 1687
rect 1797 1681 1798 1687
rect 1790 1547 1798 1681
rect 1790 1541 1791 1547
rect 1797 1541 1798 1547
rect 1790 1411 1798 1541
rect 1790 1405 1791 1411
rect 1797 1405 1798 1411
rect 1790 1275 1798 1405
rect 1790 1269 1791 1275
rect 1797 1269 1798 1275
rect 1790 1135 1798 1269
rect 1790 1129 1791 1135
rect 1797 1129 1798 1135
rect 1790 995 1798 1129
rect 1790 989 1791 995
rect 1797 989 1798 995
rect 1790 859 1798 989
rect 1790 853 1791 859
rect 1797 853 1798 859
rect 1790 723 1798 853
rect 1790 717 1791 723
rect 1797 717 1798 723
rect 1790 591 1798 717
rect 1790 585 1791 591
rect 1797 585 1798 591
rect 1790 583 1798 585
rect 1790 577 1791 583
rect 1797 577 1798 583
rect 1790 447 1798 577
rect 1790 441 1791 447
rect 1797 441 1798 447
rect 1790 311 1798 441
rect 1790 305 1791 311
rect 1797 305 1798 311
rect 1790 151 1798 305
rect 1790 145 1791 151
rect 1797 145 1798 151
rect 1790 72 1798 145
rect 3486 3431 3494 3528
rect 3486 3425 3487 3431
rect 3493 3425 3494 3431
rect 3486 3167 3494 3425
rect 3486 3161 3487 3167
rect 3493 3161 3494 3167
rect 3486 2175 3494 3161
rect 3486 2169 3487 2175
rect 3493 2169 3494 2175
rect 3486 2035 3494 2169
rect 3486 2029 3487 2035
rect 3493 2029 3494 2035
rect 3486 1899 3494 2029
rect 3486 1893 3487 1899
rect 3493 1893 3494 1899
rect 3486 511 3494 1893
rect 3486 505 3487 511
rect 3493 505 3494 511
rect 3486 72 3494 505
rect 3498 3495 3506 3528
rect 3498 3489 3499 3495
rect 3505 3489 3506 3495
rect 3498 3231 3506 3489
rect 3498 3225 3499 3231
rect 3505 3225 3506 3231
rect 3498 2807 3506 3225
rect 3498 2801 3499 2807
rect 3505 2801 3506 2807
rect 3498 2103 3506 2801
rect 3498 2097 3499 2103
rect 3505 2097 3506 2103
rect 3498 1967 3506 2097
rect 3498 1961 3499 1967
rect 3505 1961 3506 1967
rect 3498 591 3506 1961
rect 3498 585 3499 591
rect 3505 585 3506 591
rect 3498 72 3506 585
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__195
timestamp 1731220337
transform 1 0 3456 0 1 3448
box 7 3 12 24
use welltap_svt  __well_tap__194
timestamp 1731220337
transform 1 0 1800 0 1 3448
box 7 3 12 24
use welltap_svt  __well_tap__193
timestamp 1731220337
transform 1 0 3456 0 -1 3408
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220337
transform 1 0 1800 0 -1 3408
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220337
transform 1 0 3456 0 1 3316
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220337
transform 1 0 1800 0 1 3316
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220337
transform 1 0 3456 0 -1 3276
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220337
transform 1 0 1800 0 -1 3276
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220337
transform 1 0 3456 0 1 3184
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220337
transform 1 0 1800 0 1 3184
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220337
transform 1 0 3456 0 -1 3144
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220337
transform 1 0 1800 0 -1 3144
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220337
transform 1 0 3456 0 1 3048
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220337
transform 1 0 1800 0 1 3048
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220337
transform 1 0 3456 0 -1 2992
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220337
transform 1 0 1800 0 -1 2992
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220337
transform 1 0 3456 0 1 2892
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220337
transform 1 0 1800 0 1 2892
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220337
transform 1 0 3456 0 -1 2852
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220337
transform 1 0 1800 0 -1 2852
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220337
transform 1 0 3456 0 1 2760
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220337
transform 1 0 1800 0 1 2760
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220337
transform 1 0 3456 0 -1 2704
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220337
transform 1 0 1800 0 -1 2704
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220337
transform 1 0 3456 0 1 2604
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220337
transform 1 0 1800 0 1 2604
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220337
transform 1 0 3456 0 -1 2552
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220337
transform 1 0 1800 0 -1 2552
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220337
transform 1 0 3456 0 1 2464
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220337
transform 1 0 1800 0 1 2464
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220337
transform 1 0 3456 0 -1 2416
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220337
transform 1 0 1800 0 -1 2416
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220337
transform 1 0 3456 0 1 2328
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220337
transform 1 0 1800 0 1 2328
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220337
transform 1 0 3456 0 -1 2280
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220337
transform 1 0 1800 0 -1 2280
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220337
transform 1 0 3456 0 1 2192
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220337
transform 1 0 1800 0 1 2192
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220337
transform 1 0 3456 0 -1 2152
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220337
transform 1 0 1800 0 -1 2152
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220337
transform 1 0 3456 0 1 2056
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220337
transform 1 0 1800 0 1 2056
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220337
transform 1 0 3456 0 -1 2012
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220337
transform 1 0 1800 0 -1 2012
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220337
transform 1 0 3456 0 1 1920
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220337
transform 1 0 1800 0 1 1920
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220337
transform 1 0 3456 0 -1 1876
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220337
transform 1 0 1800 0 -1 1876
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220337
transform 1 0 3456 0 1 1780
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220337
transform 1 0 1800 0 1 1780
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220337
transform 1 0 3456 0 -1 1728
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220337
transform 1 0 1800 0 -1 1728
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220337
transform 1 0 3456 0 1 1636
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220337
transform 1 0 1800 0 1 1636
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220337
transform 1 0 3456 0 -1 1592
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220337
transform 1 0 1800 0 -1 1592
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220337
transform 1 0 3456 0 1 1504
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220337
transform 1 0 1800 0 1 1504
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220337
transform 1 0 3456 0 -1 1456
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220337
transform 1 0 1800 0 -1 1456
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220337
transform 1 0 3456 0 1 1364
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220337
transform 1 0 1800 0 1 1364
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220337
transform 1 0 3456 0 -1 1316
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220337
transform 1 0 1800 0 -1 1316
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220337
transform 1 0 3456 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220337
transform 1 0 1800 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220337
transform 1 0 3456 0 -1 1180
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220337
transform 1 0 1800 0 -1 1180
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220337
transform 1 0 3456 0 1 1084
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220337
transform 1 0 1800 0 1 1084
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220337
transform 1 0 3456 0 -1 1040
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220337
transform 1 0 1800 0 -1 1040
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220337
transform 1 0 3456 0 1 948
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220337
transform 1 0 1800 0 1 948
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220337
transform 1 0 3456 0 -1 908
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220337
transform 1 0 1800 0 -1 908
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220337
transform 1 0 3456 0 1 812
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220337
transform 1 0 1800 0 1 812
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220337
transform 1 0 3456 0 -1 768
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220337
transform 1 0 1800 0 -1 768
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220337
transform 1 0 3456 0 1 680
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220337
transform 1 0 1800 0 1 680
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220337
transform 1 0 3456 0 -1 632
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220337
transform 1 0 1800 0 -1 632
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220337
transform 1 0 3456 0 1 544
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220337
transform 1 0 1800 0 1 544
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220337
transform 1 0 3456 0 -1 488
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220337
transform 1 0 1800 0 -1 488
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220337
transform 1 0 3456 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220337
transform 1 0 1800 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220337
transform 1 0 3456 0 -1 356
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220337
transform 1 0 1800 0 -1 356
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220337
transform 1 0 3456 0 1 268
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220337
transform 1 0 1800 0 1 268
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220337
transform 1 0 3456 0 -1 220
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220337
transform 1 0 1800 0 -1 220
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220337
transform 1 0 3456 0 1 108
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220337
transform 1 0 1800 0 1 108
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220337
transform 1 0 1760 0 1 3460
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220337
transform 1 0 104 0 1 3460
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220337
transform 1 0 1760 0 -1 3416
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220337
transform 1 0 104 0 -1 3416
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220337
transform 1 0 1760 0 1 3320
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220337
transform 1 0 104 0 1 3320
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220337
transform 1 0 1760 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220337
transform 1 0 104 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220337
transform 1 0 1760 0 1 3176
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220337
transform 1 0 104 0 1 3176
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220337
transform 1 0 1760 0 -1 3136
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220337
transform 1 0 104 0 -1 3136
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220337
transform 1 0 1760 0 1 3044
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220337
transform 1 0 104 0 1 3044
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220337
transform 1 0 1760 0 -1 2996
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220337
transform 1 0 104 0 -1 2996
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220337
transform 1 0 1760 0 1 2896
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220337
transform 1 0 104 0 1 2896
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220337
transform 1 0 1760 0 -1 2848
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220337
transform 1 0 104 0 -1 2848
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220337
transform 1 0 1760 0 1 2748
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220337
transform 1 0 104 0 1 2748
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220337
transform 1 0 1760 0 -1 2700
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220337
transform 1 0 104 0 -1 2700
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220337
transform 1 0 1760 0 1 2604
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220337
transform 1 0 104 0 1 2604
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220337
transform 1 0 1760 0 -1 2556
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220337
transform 1 0 104 0 -1 2556
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220337
transform 1 0 1760 0 1 2460
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220337
transform 1 0 104 0 1 2460
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220337
transform 1 0 1760 0 -1 2420
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220337
transform 1 0 104 0 -1 2420
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220337
transform 1 0 1760 0 1 2328
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220337
transform 1 0 104 0 1 2328
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220337
transform 1 0 1760 0 -1 2280
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220337
transform 1 0 104 0 -1 2280
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220337
transform 1 0 1760 0 1 2188
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220337
transform 1 0 104 0 1 2188
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220337
transform 1 0 1760 0 -1 2140
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220337
transform 1 0 104 0 -1 2140
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220337
transform 1 0 1760 0 1 2048
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220337
transform 1 0 104 0 1 2048
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220337
transform 1 0 1760 0 -1 2000
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220337
transform 1 0 104 0 -1 2000
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220337
transform 1 0 1760 0 1 1908
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220337
transform 1 0 104 0 1 1908
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220337
transform 1 0 1760 0 -1 1868
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220337
transform 1 0 104 0 -1 1868
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220337
transform 1 0 1760 0 1 1776
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220337
transform 1 0 104 0 1 1776
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220337
transform 1 0 1760 0 -1 1732
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220337
transform 1 0 104 0 -1 1732
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220337
transform 1 0 1760 0 1 1640
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220337
transform 1 0 104 0 1 1640
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220337
transform 1 0 1760 0 -1 1596
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220337
transform 1 0 104 0 -1 1596
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220337
transform 1 0 1760 0 1 1500
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220337
transform 1 0 104 0 1 1500
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220337
transform 1 0 1760 0 -1 1456
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220337
transform 1 0 104 0 -1 1456
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220337
transform 1 0 1760 0 1 1364
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220337
transform 1 0 104 0 1 1364
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220337
transform 1 0 1760 0 -1 1320
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220337
transform 1 0 104 0 -1 1320
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220337
transform 1 0 1760 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220337
transform 1 0 104 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220337
transform 1 0 1760 0 -1 1180
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220337
transform 1 0 104 0 -1 1180
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220337
transform 1 0 1760 0 1 1088
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220337
transform 1 0 104 0 1 1088
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220337
transform 1 0 1760 0 -1 1044
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220337
transform 1 0 104 0 -1 1044
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220337
transform 1 0 1760 0 1 948
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220337
transform 1 0 104 0 1 948
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220337
transform 1 0 1760 0 -1 904
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220337
transform 1 0 104 0 -1 904
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220337
transform 1 0 1760 0 1 812
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220337
transform 1 0 104 0 1 812
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220337
transform 1 0 1760 0 -1 768
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220337
transform 1 0 104 0 -1 768
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220337
transform 1 0 1760 0 1 676
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220337
transform 1 0 104 0 1 676
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220337
transform 1 0 1760 0 -1 632
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220337
transform 1 0 104 0 -1 632
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220337
transform 1 0 1760 0 1 536
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220337
transform 1 0 104 0 1 536
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220337
transform 1 0 1760 0 -1 496
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220337
transform 1 0 104 0 -1 496
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220337
transform 1 0 1760 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220337
transform 1 0 104 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220337
transform 1 0 1760 0 -1 356
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220337
transform 1 0 104 0 -1 356
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220337
transform 1 0 1760 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220337
transform 1 0 104 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220337
transform 1 0 1760 0 -1 220
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220337
transform 1 0 104 0 -1 220
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220337
transform 1 0 1760 0 1 104
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220337
transform 1 0 104 0 1 104
box 7 3 12 24
use _0_0cell_0_0gcelem2x0  tst_5999_6
timestamp 1731220337
transform 1 0 3272 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5998_6
timestamp 1731220337
transform 1 0 3360 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5997_6
timestamp 1731220337
transform 1 0 3360 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5996_6
timestamp 1731220337
transform 1 0 3360 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5995_6
timestamp 1731220337
transform 1 0 3352 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5994_6
timestamp 1731220337
transform 1 0 3328 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5993_6
timestamp 1731220337
transform 1 0 3256 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5992_6
timestamp 1731220337
transform 1 0 3128 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5991_6
timestamp 1731220337
transform 1 0 3184 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5990_6
timestamp 1731220337
transform 1 0 3096 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5989_6
timestamp 1731220337
transform 1 0 3000 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5988_6
timestamp 1731220337
transform 1 0 2904 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5987_6
timestamp 1731220337
transform 1 0 2808 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5986_6
timestamp 1731220337
transform 1 0 2712 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5985_6
timestamp 1731220337
transform 1 0 2608 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5984_6
timestamp 1731220337
transform 1 0 2504 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5983_6
timestamp 1731220337
transform 1 0 2760 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5982_6
timestamp 1731220337
transform 1 0 2888 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5981_6
timestamp 1731220337
transform 1 0 3008 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5980_6
timestamp 1731220337
transform 1 0 3216 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5979_6
timestamp 1731220337
transform 1 0 3064 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5978_6
timestamp 1731220337
transform 1 0 2920 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5977_6
timestamp 1731220337
transform 1 0 2792 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5976_6
timestamp 1731220337
transform 1 0 2672 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5975_6
timestamp 1731220337
transform 1 0 3144 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5974_6
timestamp 1731220337
transform 1 0 2944 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5973_6
timestamp 1731220337
transform 1 0 2752 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5972_6
timestamp 1731220337
transform 1 0 2576 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5971_6
timestamp 1731220337
transform 1 0 3096 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5970_6
timestamp 1731220337
transform 1 0 2864 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5969_6
timestamp 1731220337
transform 1 0 2648 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5968_6
timestamp 1731220337
transform 1 0 2448 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5967_6
timestamp 1731220337
transform 1 0 2264 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5966_6
timestamp 1731220337
transform 1 0 2288 0 -1 508
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5965_6
timestamp 1731220337
transform 1 0 2472 0 -1 508
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5964_6
timestamp 1731220337
transform 1 0 2672 0 -1 508
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5963_6
timestamp 1731220337
transform 1 0 3104 0 -1 508
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5962_6
timestamp 1731220337
transform 1 0 2880 0 -1 508
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5961_6
timestamp 1731220337
transform 1 0 2792 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5960_6
timestamp 1731220337
transform 1 0 2616 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5959_6
timestamp 1731220337
transform 1 0 2448 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5958_6
timestamp 1731220337
transform 1 0 2976 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5957_6
timestamp 1731220337
transform 1 0 3160 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5956_6
timestamp 1731220337
transform 1 0 3096 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5955_6
timestamp 1731220337
transform 1 0 2952 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5954_6
timestamp 1731220337
transform 1 0 2808 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5953_6
timestamp 1731220337
transform 1 0 2648 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5952_6
timestamp 1731220337
transform 1 0 2696 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5951_6
timestamp 1731220337
transform 1 0 2840 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5950_6
timestamp 1731220337
transform 1 0 2976 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5949_6
timestamp 1731220337
transform 1 0 3208 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5948_6
timestamp 1731220337
transform 1 0 3032 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5947_6
timestamp 1731220337
transform 1 0 2864 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5946_6
timestamp 1731220337
transform 1 0 2704 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5945_6
timestamp 1731220337
transform 1 0 3056 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5944_6
timestamp 1731220337
transform 1 0 2904 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5943_6
timestamp 1731220337
transform 1 0 2760 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5942_6
timestamp 1731220337
transform 1 0 2632 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5941_6
timestamp 1731220337
transform 1 0 2824 0 -1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5940_6
timestamp 1731220337
transform 1 0 2736 0 -1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5939_6
timestamp 1731220337
transform 1 0 2648 0 -1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5938_6
timestamp 1731220337
transform 1 0 2560 0 -1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5937_6
timestamp 1731220337
transform 1 0 2384 0 -1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5936_6
timestamp 1731220337
transform 1 0 2296 0 -1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5935_6
timestamp 1731220337
transform 1 0 2208 0 -1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5934_6
timestamp 1731220337
transform 1 0 2120 0 -1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5933_6
timestamp 1731220337
transform 1 0 2128 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5932_6
timestamp 1731220337
transform 1 0 2456 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5931_6
timestamp 1731220337
transform 1 0 2624 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5930_6
timestamp 1731220337
transform 1 0 2984 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5929_6
timestamp 1731220337
transform 1 0 2800 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5928_6
timestamp 1731220337
transform 1 0 2696 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5927_6
timestamp 1731220337
transform 1 0 2536 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5926_6
timestamp 1731220337
transform 1 0 3024 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5925_6
timestamp 1731220337
transform 1 0 2856 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5924_6
timestamp 1731220337
transform 1 0 2744 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5923_6
timestamp 1731220337
transform 1 0 2592 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5922_6
timestamp 1731220337
transform 1 0 2896 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5921_6
timestamp 1731220337
transform 1 0 3056 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5920_6
timestamp 1731220337
transform 1 0 2968 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5919_6
timestamp 1731220337
transform 1 0 2832 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5918_6
timestamp 1731220337
transform 1 0 2696 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5917_6
timestamp 1731220337
transform 1 0 2592 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5916_6
timestamp 1731220337
transform 1 0 2352 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5915_6
timestamp 1731220337
transform 1 0 2800 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5914_6
timestamp 1731220337
transform 1 0 2680 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5913_6
timestamp 1731220337
transform 1 0 2856 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5912_6
timestamp 1731220337
transform 1 0 3032 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5911_6
timestamp 1731220337
transform 1 0 3208 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5910_6
timestamp 1731220337
transform 1 0 3192 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5909_6
timestamp 1731220337
transform 1 0 3000 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5908_6
timestamp 1731220337
transform 1 0 3104 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5907_6
timestamp 1731220337
transform 1 0 3240 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5906_6
timestamp 1731220337
transform 1 0 3216 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5905_6
timestamp 1731220337
transform 1 0 3200 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5904_6
timestamp 1731220337
transform 1 0 3176 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5903_6
timestamp 1731220337
transform 1 0 3216 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5902_6
timestamp 1731220337
transform 1 0 3112 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5901_6
timestamp 1731220337
transform 1 0 3248 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5900_6
timestamp 1731220337
transform 1 0 3240 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5899_6
timestamp 1731220337
transform 1 0 3328 0 -1 508
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5898_6
timestamp 1731220337
transform 1 0 3352 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5897_6
timestamp 1731220337
transform 1 0 3360 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5896_6
timestamp 1731220337
transform 1 0 3360 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5895_6
timestamp 1731220337
transform 1 0 3360 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5894_6
timestamp 1731220337
transform 1 0 3360 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5893_6
timestamp 1731220337
transform 1 0 3360 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5892_6
timestamp 1731220337
transform 1 0 3360 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5891_6
timestamp 1731220337
transform 1 0 3360 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5890_6
timestamp 1731220337
transform 1 0 3360 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5889_6
timestamp 1731220337
transform 1 0 3360 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5888_6
timestamp 1731220337
transform 1 0 3360 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5887_6
timestamp 1731220337
transform 1 0 3360 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5886_6
timestamp 1731220337
transform 1 0 3360 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5885_6
timestamp 1731220337
transform 1 0 3256 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5884_6
timestamp 1731220337
transform 1 0 3248 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5883_6
timestamp 1731220337
transform 1 0 3120 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5882_6
timestamp 1731220337
transform 1 0 2992 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5881_6
timestamp 1731220337
transform 1 0 2856 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5880_6
timestamp 1731220337
transform 1 0 2712 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5879_6
timestamp 1731220337
transform 1 0 2552 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5878_6
timestamp 1731220337
transform 1 0 3128 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5877_6
timestamp 1731220337
transform 1 0 3000 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5876_6
timestamp 1731220337
transform 1 0 2864 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5875_6
timestamp 1731220337
transform 1 0 2728 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5874_6
timestamp 1731220337
transform 1 0 2584 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5873_6
timestamp 1731220337
transform 1 0 3048 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5872_6
timestamp 1731220337
transform 1 0 2920 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5871_6
timestamp 1731220337
transform 1 0 2792 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5870_6
timestamp 1731220337
transform 1 0 2672 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5869_6
timestamp 1731220337
transform 1 0 2544 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5868_6
timestamp 1731220337
transform 1 0 2880 0 -1 1612
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5867_6
timestamp 1731220337
transform 1 0 2768 0 -1 1612
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5866_6
timestamp 1731220337
transform 1 0 2664 0 -1 1612
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5865_6
timestamp 1731220337
transform 1 0 2560 0 -1 1612
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5864_6
timestamp 1731220337
transform 1 0 2888 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5863_6
timestamp 1731220337
transform 1 0 2800 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5862_6
timestamp 1731220337
transform 1 0 2712 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5861_6
timestamp 1731220337
transform 1 0 2624 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5860_6
timestamp 1731220337
transform 1 0 2536 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5859_6
timestamp 1731220337
transform 1 0 2576 0 -1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5858_6
timestamp 1731220337
transform 1 0 2840 0 -1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5857_6
timestamp 1731220337
transform 1 0 2752 0 -1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5856_6
timestamp 1731220337
transform 1 0 2664 0 -1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5855_6
timestamp 1731220337
transform 1 0 2624 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5854_6
timestamp 1731220337
transform 1 0 2536 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5853_6
timestamp 1731220337
transform 1 0 2712 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5852_6
timestamp 1731220337
transform 1 0 2800 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5851_6
timestamp 1731220337
transform 1 0 2888 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5850_6
timestamp 1731220337
transform 1 0 2976 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5849_6
timestamp 1731220337
transform 1 0 2864 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5848_6
timestamp 1731220337
transform 1 0 2752 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5847_6
timestamp 1731220337
transform 1 0 2640 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5846_6
timestamp 1731220337
transform 1 0 2536 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5845_6
timestamp 1731220337
transform 1 0 2568 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5844_6
timestamp 1731220337
transform 1 0 2704 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5843_6
timestamp 1731220337
transform 1 0 2824 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5842_6
timestamp 1731220337
transform 1 0 2944 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5841_6
timestamp 1731220337
transform 1 0 3000 0 -1 2032
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5840_6
timestamp 1731220337
transform 1 0 2816 0 -1 2032
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5839_6
timestamp 1731220337
transform 1 0 2624 0 -1 2032
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5838_6
timestamp 1731220337
transform 1 0 2496 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5837_6
timestamp 1731220337
transform 1 0 2648 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5836_6
timestamp 1731220337
transform 1 0 2784 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5835_6
timestamp 1731220337
transform 1 0 2912 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5834_6
timestamp 1731220337
transform 1 0 3184 0 -1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5833_6
timestamp 1731220337
transform 1 0 3264 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5832_6
timestamp 1731220337
transform 1 0 3152 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5831_6
timestamp 1731220337
transform 1 0 3032 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5830_6
timestamp 1731220337
transform 1 0 3192 0 -1 2032
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5829_6
timestamp 1731220337
transform 1 0 3160 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5828_6
timestamp 1731220337
transform 1 0 3056 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5827_6
timestamp 1731220337
transform 1 0 3272 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5826_6
timestamp 1731220337
transform 1 0 3360 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5825_6
timestamp 1731220337
transform 1 0 3360 0 -1 2032
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5824_6
timestamp 1731220337
transform 1 0 3360 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5823_6
timestamp 1731220337
transform 1 0 3272 0 -1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5822_6
timestamp 1731220337
transform 1 0 3360 0 -1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5821_6
timestamp 1731220337
transform 1 0 3360 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5820_6
timestamp 1731220337
transform 1 0 3360 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5819_6
timestamp 1731220337
transform 1 0 3216 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5818_6
timestamp 1731220337
transform 1 0 3048 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5817_6
timestamp 1731220337
transform 1 0 2952 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5816_6
timestamp 1731220337
transform 1 0 3096 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5815_6
timestamp 1731220337
transform 1 0 3240 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5814_6
timestamp 1731220337
transform 1 0 3096 0 -1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5813_6
timestamp 1731220337
transform 1 0 3008 0 -1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5812_6
timestamp 1731220337
transform 1 0 2920 0 -1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5811_6
timestamp 1731220337
transform 1 0 2808 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5810_6
timestamp 1731220337
transform 1 0 2648 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5809_6
timestamp 1731220337
transform 1 0 2712 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5808_6
timestamp 1731220337
transform 1 0 2880 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5807_6
timestamp 1731220337
transform 1 0 3016 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5806_6
timestamp 1731220337
transform 1 0 2904 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5805_6
timestamp 1731220337
transform 1 0 2792 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5804_6
timestamp 1731220337
transform 1 0 2680 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5803_6
timestamp 1731220337
transform 1 0 2928 0 -1 2436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5802_6
timestamp 1731220337
transform 1 0 2832 0 -1 2436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5801_6
timestamp 1731220337
transform 1 0 2736 0 -1 2436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5800_6
timestamp 1731220337
transform 1 0 2648 0 -1 2436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5799_6
timestamp 1731220337
transform 1 0 2560 0 -1 2436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5798_6
timestamp 1731220337
transform 1 0 3136 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5797_6
timestamp 1731220337
transform 1 0 2912 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5796_6
timestamp 1731220337
transform 1 0 2704 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5795_6
timestamp 1731220337
transform 1 0 2520 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5794_6
timestamp 1731220337
transform 1 0 2992 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5793_6
timestamp 1731220337
transform 1 0 2808 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5792_6
timestamp 1731220337
transform 1 0 2640 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5791_6
timestamp 1731220337
transform 1 0 2480 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5790_6
timestamp 1731220337
transform 1 0 2336 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5789_6
timestamp 1731220337
transform 1 0 2424 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5788_6
timestamp 1731220337
transform 1 0 2576 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5787_6
timestamp 1731220337
transform 1 0 3160 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5786_6
timestamp 1731220337
transform 1 0 2952 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5785_6
timestamp 1731220337
transform 1 0 2752 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5784_6
timestamp 1731220337
transform 1 0 2680 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5783_6
timestamp 1731220337
transform 1 0 2536 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5782_6
timestamp 1731220337
transform 1 0 2840 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5781_6
timestamp 1731220337
transform 1 0 3200 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5780_6
timestamp 1731220337
transform 1 0 3016 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5779_6
timestamp 1731220337
transform 1 0 2904 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5778_6
timestamp 1731220337
transform 1 0 2744 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5777_6
timestamp 1731220337
transform 1 0 2576 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5776_6
timestamp 1731220337
transform 1 0 3064 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5775_6
timestamp 1731220337
transform 1 0 3056 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5774_6
timestamp 1731220337
transform 1 0 2896 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5773_6
timestamp 1731220337
transform 1 0 2728 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5772_6
timestamp 1731220337
transform 1 0 2752 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5771_6
timestamp 1731220337
transform 1 0 2904 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5770_6
timestamp 1731220337
transform 1 0 3056 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5769_6
timestamp 1731220337
transform 1 0 3200 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5768_6
timestamp 1731220337
transform 1 0 3352 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5767_6
timestamp 1731220337
transform 1 0 3216 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5766_6
timestamp 1731220337
transform 1 0 3224 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5765_6
timestamp 1731220337
transform 1 0 3184 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5764_6
timestamp 1731220337
transform 1 0 3360 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5763_6
timestamp 1731220337
transform 1 0 3360 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5762_6
timestamp 1731220337
transform 1 0 3360 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5761_6
timestamp 1731220337
transform 1 0 3360 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5760_6
timestamp 1731220337
transform 1 0 3360 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5759_6
timestamp 1731220337
transform 1 0 3360 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5758_6
timestamp 1731220337
transform 1 0 3360 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5757_6
timestamp 1731220337
transform 1 0 3360 0 1 3028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5756_6
timestamp 1731220337
transform 1 0 3360 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5755_6
timestamp 1731220337
transform 1 0 3328 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5754_6
timestamp 1731220337
transform 1 0 3224 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5753_6
timestamp 1731220337
transform 1 0 3072 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5752_6
timestamp 1731220337
transform 1 0 2912 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5751_6
timestamp 1731220337
transform 1 0 3000 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5750_6
timestamp 1731220337
transform 1 0 3160 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5749_6
timestamp 1731220337
transform 1 0 3192 0 -1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5748_6
timestamp 1731220337
transform 1 0 3032 0 -1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5747_6
timestamp 1731220337
transform 1 0 2872 0 -1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5746_6
timestamp 1731220337
transform 1 0 2832 0 1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5745_6
timestamp 1731220337
transform 1 0 2968 0 1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5744_6
timestamp 1731220337
transform 1 0 3112 0 1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5743_6
timestamp 1731220337
transform 1 0 3144 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5742_6
timestamp 1731220337
transform 1 0 3032 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5741_6
timestamp 1731220337
transform 1 0 2928 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5740_6
timestamp 1731220337
transform 1 0 2824 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5739_6
timestamp 1731220337
transform 1 0 2960 0 1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5738_6
timestamp 1731220337
transform 1 0 2792 0 1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5737_6
timestamp 1731220337
transform 1 0 2632 0 1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5736_6
timestamp 1731220337
transform 1 0 2472 0 1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5735_6
timestamp 1731220337
transform 1 0 2504 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5734_6
timestamp 1731220337
transform 1 0 2616 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5733_6
timestamp 1731220337
transform 1 0 2720 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5732_6
timestamp 1731220337
transform 1 0 2696 0 1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5731_6
timestamp 1731220337
transform 1 0 2712 0 -1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5730_6
timestamp 1731220337
transform 1 0 2680 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5729_6
timestamp 1731220337
transform 1 0 2840 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5728_6
timestamp 1731220337
transform 1 0 2752 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5727_6
timestamp 1731220337
transform 1 0 2576 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5726_6
timestamp 1731220337
transform 1 0 3144 0 1 3028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5725_6
timestamp 1731220337
transform 1 0 2912 0 1 3028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5724_6
timestamp 1731220337
transform 1 0 2688 0 1 3028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5723_6
timestamp 1731220337
transform 1 0 2480 0 1 3028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5722_6
timestamp 1731220337
transform 1 0 3176 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5721_6
timestamp 1731220337
transform 1 0 2976 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5720_6
timestamp 1731220337
transform 1 0 2784 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5719_6
timestamp 1731220337
transform 1 0 2616 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5718_6
timestamp 1731220337
transform 1 0 2472 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5717_6
timestamp 1731220337
transform 1 0 2352 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5716_6
timestamp 1731220337
transform 1 0 2240 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5715_6
timestamp 1731220337
transform 1 0 2136 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5714_6
timestamp 1731220337
transform 1 0 2208 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5713_6
timestamp 1731220337
transform 1 0 2400 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5712_6
timestamp 1731220337
transform 1 0 2584 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5711_6
timestamp 1731220337
transform 1 0 2560 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5710_6
timestamp 1731220337
transform 1 0 2376 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5709_6
timestamp 1731220337
transform 1 0 2184 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5708_6
timestamp 1731220337
transform 1 0 2008 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5707_6
timestamp 1731220337
transform 1 0 2208 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5706_6
timestamp 1731220337
transform 1 0 2400 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5705_6
timestamp 1731220337
transform 1 0 2400 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5704_6
timestamp 1731220337
transform 1 0 2272 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5703_6
timestamp 1731220337
transform 1 0 2152 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5702_6
timestamp 1731220337
transform 1 0 2032 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5701_6
timestamp 1731220337
transform 1 0 2288 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5700_6
timestamp 1731220337
transform 1 0 2176 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5699_6
timestamp 1731220337
transform 1 0 2064 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5698_6
timestamp 1731220337
transform 1 0 1960 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5697_6
timestamp 1731220337
transform 1 0 1864 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5696_6
timestamp 1731220337
transform 1 0 1824 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5695_6
timestamp 1731220337
transform 1 0 1912 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5694_6
timestamp 1731220337
transform 1 0 2000 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5693_6
timestamp 1731220337
transform 1 0 2104 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5692_6
timestamp 1731220337
transform 1 0 2216 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5691_6
timestamp 1731220337
transform 1 0 2128 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5690_6
timestamp 1731220337
transform 1 0 2032 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5689_6
timestamp 1731220337
transform 1 0 1944 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5688_6
timestamp 1731220337
transform 1 0 2232 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5687_6
timestamp 1731220337
transform 1 0 2360 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5686_6
timestamp 1731220337
transform 1 0 2296 0 -1 2436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5685_6
timestamp 1731220337
transform 1 0 2208 0 -1 2436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5684_6
timestamp 1731220337
transform 1 0 2384 0 -1 2436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5683_6
timestamp 1731220337
transform 1 0 2472 0 -1 2436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5682_6
timestamp 1731220337
transform 1 0 2568 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5681_6
timestamp 1731220337
transform 1 0 2464 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5680_6
timestamp 1731220337
transform 1 0 2360 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5679_6
timestamp 1731220337
transform 1 0 2256 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5678_6
timestamp 1731220337
transform 1 0 2160 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5677_6
timestamp 1731220337
transform 1 0 2544 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5676_6
timestamp 1731220337
transform 1 0 2368 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5675_6
timestamp 1731220337
transform 1 0 2192 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5674_6
timestamp 1731220337
transform 1 0 2032 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5673_6
timestamp 1731220337
transform 1 0 1880 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5672_6
timestamp 1731220337
transform 1 0 2480 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5671_6
timestamp 1731220337
transform 1 0 2304 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5670_6
timestamp 1731220337
transform 1 0 2128 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5669_6
timestamp 1731220337
transform 1 0 1960 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5668_6
timestamp 1731220337
transform 1 0 1824 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5667_6
timestamp 1731220337
transform 1 0 1664 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5666_6
timestamp 1731220337
transform 1 0 1496 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5665_6
timestamp 1731220337
transform 1 0 1312 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5664_6
timestamp 1731220337
transform 1 0 1224 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5663_6
timestamp 1731220337
transform 1 0 1096 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5662_6
timestamp 1731220337
transform 1 0 1344 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5661_6
timestamp 1731220337
transform 1 0 1456 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5660_6
timestamp 1731220337
transform 1 0 1568 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5659_6
timestamp 1731220337
transform 1 0 1664 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5658_6
timestamp 1731220337
transform 1 0 1824 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5657_6
timestamp 1731220337
transform 1 0 1984 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5656_6
timestamp 1731220337
transform 1 0 2160 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5655_6
timestamp 1731220337
transform 1 0 2336 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5654_6
timestamp 1731220337
transform 1 0 2424 0 -1 2032
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5653_6
timestamp 1731220337
transform 1 0 2216 0 -1 2032
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5652_6
timestamp 1731220337
transform 1 0 2008 0 -1 2032
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5651_6
timestamp 1731220337
transform 1 0 1824 0 -1 2032
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5650_6
timestamp 1731220337
transform 1 0 1856 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5649_6
timestamp 1731220337
transform 1 0 1992 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5648_6
timestamp 1731220337
transform 1 0 2136 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5647_6
timestamp 1731220337
transform 1 0 2424 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5646_6
timestamp 1731220337
transform 1 0 2280 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5645_6
timestamp 1731220337
transform 1 0 2208 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5644_6
timestamp 1731220337
transform 1 0 2104 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5643_6
timestamp 1731220337
transform 1 0 2008 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5642_6
timestamp 1731220337
transform 1 0 2320 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5641_6
timestamp 1731220337
transform 1 0 2432 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5640_6
timestamp 1731220337
transform 1 0 2448 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5639_6
timestamp 1731220337
transform 1 0 2360 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5638_6
timestamp 1731220337
transform 1 0 2272 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5637_6
timestamp 1731220337
transform 1 0 2184 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5636_6
timestamp 1731220337
transform 1 0 2096 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5635_6
timestamp 1731220337
transform 1 0 2136 0 -1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5634_6
timestamp 1731220337
transform 1 0 2224 0 -1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5633_6
timestamp 1731220337
transform 1 0 2312 0 -1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5632_6
timestamp 1731220337
transform 1 0 2400 0 -1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5631_6
timestamp 1731220337
transform 1 0 2488 0 -1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5630_6
timestamp 1731220337
transform 1 0 2448 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5629_6
timestamp 1731220337
transform 1 0 2360 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5628_6
timestamp 1731220337
transform 1 0 2272 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5627_6
timestamp 1731220337
transform 1 0 2184 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5626_6
timestamp 1731220337
transform 1 0 2096 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5625_6
timestamp 1731220337
transform 1 0 2456 0 -1 1612
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5624_6
timestamp 1731220337
transform 1 0 2352 0 -1 1612
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5623_6
timestamp 1731220337
transform 1 0 2248 0 -1 1612
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5622_6
timestamp 1731220337
transform 1 0 2152 0 -1 1612
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5621_6
timestamp 1731220337
transform 1 0 2056 0 -1 1612
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5620_6
timestamp 1731220337
transform 1 0 2416 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5619_6
timestamp 1731220337
transform 1 0 2288 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5618_6
timestamp 1731220337
transform 1 0 2160 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5617_6
timestamp 1731220337
transform 1 0 2032 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5616_6
timestamp 1731220337
transform 1 0 1912 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5615_6
timestamp 1731220337
transform 1 0 2424 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5614_6
timestamp 1731220337
transform 1 0 2264 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5613_6
timestamp 1731220337
transform 1 0 2104 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5612_6
timestamp 1731220337
transform 1 0 1944 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5611_6
timestamp 1731220337
transform 1 0 1824 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5610_6
timestamp 1731220337
transform 1 0 2376 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5609_6
timestamp 1731220337
transform 1 0 2192 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5608_6
timestamp 1731220337
transform 1 0 2000 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5607_6
timestamp 1731220337
transform 1 0 1664 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5606_6
timestamp 1731220337
transform 1 0 1824 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5605_6
timestamp 1731220337
transform 1 0 1824 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5604_6
timestamp 1731220337
transform 1 0 1960 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5603_6
timestamp 1731220337
transform 1 0 2504 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5602_6
timestamp 1731220337
transform 1 0 2320 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5601_6
timestamp 1731220337
transform 1 0 2136 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5600_6
timestamp 1731220337
transform 1 0 2088 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5599_6
timestamp 1731220337
transform 1 0 1824 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5598_6
timestamp 1731220337
transform 1 0 1664 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5597_6
timestamp 1731220337
transform 1 0 1496 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5596_6
timestamp 1731220337
transform 1 0 1664 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5595_6
timestamp 1731220337
transform 1 0 1528 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5594_6
timestamp 1731220337
transform 1 0 1368 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5593_6
timestamp 1731220337
transform 1 0 1216 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5592_6
timestamp 1731220337
transform 1 0 1552 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5591_6
timestamp 1731220337
transform 1 0 1424 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5590_6
timestamp 1731220337
transform 1 0 1296 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5589_6
timestamp 1731220337
transform 1 0 1160 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5588_6
timestamp 1731220337
transform 1 0 1008 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5587_6
timestamp 1731220337
transform 1 0 1584 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5586_6
timestamp 1731220337
transform 1 0 1424 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5585_6
timestamp 1731220337
transform 1 0 1272 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5584_6
timestamp 1731220337
transform 1 0 1120 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5583_6
timestamp 1731220337
transform 1 0 952 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5582_6
timestamp 1731220337
transform 1 0 1440 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5581_6
timestamp 1731220337
transform 1 0 1304 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5580_6
timestamp 1731220337
transform 1 0 1168 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5579_6
timestamp 1731220337
transform 1 0 1040 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5578_6
timestamp 1731220337
transform 1 0 904 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5577_6
timestamp 1731220337
transform 1 0 1272 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5576_6
timestamp 1731220337
transform 1 0 1160 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5575_6
timestamp 1731220337
transform 1 0 1048 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5574_6
timestamp 1731220337
transform 1 0 936 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5573_6
timestamp 1731220337
transform 1 0 824 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5572_6
timestamp 1731220337
transform 1 0 752 0 1 1620
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5571_6
timestamp 1731220337
transform 1 0 848 0 1 1620
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5570_6
timestamp 1731220337
transform 1 0 944 0 1 1620
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5569_6
timestamp 1731220337
transform 1 0 1136 0 1 1620
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5568_6
timestamp 1731220337
transform 1 0 1040 0 1 1620
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5567_6
timestamp 1731220337
transform 1 0 944 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5566_6
timestamp 1731220337
transform 1 0 1048 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5565_6
timestamp 1731220337
transform 1 0 1152 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5564_6
timestamp 1731220337
transform 1 0 1264 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5563_6
timestamp 1731220337
transform 1 0 1376 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5562_6
timestamp 1731220337
transform 1 0 1272 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5561_6
timestamp 1731220337
transform 1 0 1144 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5560_6
timestamp 1731220337
transform 1 0 1400 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5559_6
timestamp 1731220337
transform 1 0 1528 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5558_6
timestamp 1731220337
transform 1 0 1664 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5557_6
timestamp 1731220337
transform 1 0 1664 0 -1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5556_6
timestamp 1731220337
transform 1 0 1504 0 -1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5555_6
timestamp 1731220337
transform 1 0 1344 0 -1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5554_6
timestamp 1731220337
transform 1 0 1192 0 -1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5553_6
timestamp 1731220337
transform 1 0 1152 0 1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5552_6
timestamp 1731220337
transform 1 0 1304 0 1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5551_6
timestamp 1731220337
transform 1 0 1464 0 1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5550_6
timestamp 1731220337
transform 1 0 1320 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5549_6
timestamp 1731220337
transform 1 0 1176 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5548_6
timestamp 1731220337
transform 1 0 1040 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5547_6
timestamp 1731220337
transform 1 0 1272 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5546_6
timestamp 1731220337
transform 1 0 1152 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5545_6
timestamp 1731220337
transform 1 0 1040 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5544_6
timestamp 1731220337
transform 1 0 968 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5543_6
timestamp 1731220337
transform 1 0 832 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5542_6
timestamp 1731220337
transform 1 0 928 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5541_6
timestamp 1731220337
transform 1 0 816 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5540_6
timestamp 1731220337
transform 1 0 696 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5539_6
timestamp 1731220337
transform 1 0 768 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5538_6
timestamp 1731220337
transform 1 0 904 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5537_6
timestamp 1731220337
transform 1 0 1000 0 1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5536_6
timestamp 1731220337
transform 1 0 848 0 1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5535_6
timestamp 1731220337
transform 1 0 880 0 -1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5534_6
timestamp 1731220337
transform 1 0 1040 0 -1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5533_6
timestamp 1731220337
transform 1 0 1016 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5532_6
timestamp 1731220337
transform 1 0 880 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5531_6
timestamp 1731220337
transform 1 0 752 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5530_6
timestamp 1731220337
transform 1 0 840 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5529_6
timestamp 1731220337
transform 1 0 736 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5528_6
timestamp 1731220337
transform 1 0 656 0 1 1620
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5527_6
timestamp 1731220337
transform 1 0 568 0 1 1620
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5526_6
timestamp 1731220337
transform 1 0 600 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5525_6
timestamp 1731220337
transform 1 0 712 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5524_6
timestamp 1731220337
transform 1 0 616 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5523_6
timestamp 1731220337
transform 1 0 760 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5522_6
timestamp 1731220337
transform 1 0 776 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5521_6
timestamp 1731220337
transform 1 0 576 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5520_6
timestamp 1731220337
transform 1 0 672 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5519_6
timestamp 1731220337
transform 1 0 848 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5518_6
timestamp 1731220337
transform 1 0 1056 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5517_6
timestamp 1731220337
transform 1 0 888 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5516_6
timestamp 1731220337
transform 1 0 720 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5515_6
timestamp 1731220337
transform 1 0 672 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5514_6
timestamp 1731220337
transform 1 0 816 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5513_6
timestamp 1731220337
transform 1 0 968 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5512_6
timestamp 1731220337
transform 1 0 1136 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5511_6
timestamp 1731220337
transform 1 0 1312 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5510_6
timestamp 1731220337
transform 1 0 1240 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5509_6
timestamp 1731220337
transform 1 0 1112 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5508_6
timestamp 1731220337
transform 1 0 984 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5507_6
timestamp 1731220337
transform 1 0 864 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5506_6
timestamp 1731220337
transform 1 0 736 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5505_6
timestamp 1731220337
transform 1 0 880 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5504_6
timestamp 1731220337
transform 1 0 1008 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5503_6
timestamp 1731220337
transform 1 0 1136 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5502_6
timestamp 1731220337
transform 1 0 1264 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5501_6
timestamp 1731220337
transform 1 0 1392 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5500_6
timestamp 1731220337
transform 1 0 1272 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5499_6
timestamp 1731220337
transform 1 0 1152 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5498_6
timestamp 1731220337
transform 1 0 1032 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5497_6
timestamp 1731220337
transform 1 0 1528 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5496_6
timestamp 1731220337
transform 1 0 1400 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5495_6
timestamp 1731220337
transform 1 0 1352 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5494_6
timestamp 1731220337
transform 1 0 1248 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5493_6
timestamp 1731220337
transform 1 0 1136 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5492_6
timestamp 1731220337
transform 1 0 1464 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5491_6
timestamp 1731220337
transform 1 0 1552 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5490_6
timestamp 1731220337
transform 1 0 1576 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5489_6
timestamp 1731220337
transform 1 0 1664 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5488_6
timestamp 1731220337
transform 1 0 1824 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5487_6
timestamp 1731220337
transform 1 0 1968 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5486_6
timestamp 1731220337
transform 1 0 1840 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5485_6
timestamp 1731220337
transform 1 0 1976 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5484_6
timestamp 1731220337
transform 1 0 2112 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5483_6
timestamp 1731220337
transform 1 0 2184 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5482_6
timestamp 1731220337
transform 1 0 2056 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5481_6
timestamp 1731220337
transform 1 0 1936 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5480_6
timestamp 1731220337
transform 1 0 1928 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5479_6
timestamp 1731220337
transform 1 0 2032 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5478_6
timestamp 1731220337
transform 1 0 2152 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5477_6
timestamp 1731220337
transform 1 0 2280 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5476_6
timestamp 1731220337
transform 1 0 2416 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5475_6
timestamp 1731220337
transform 1 0 2560 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5474_6
timestamp 1731220337
transform 1 0 2448 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5473_6
timestamp 1731220337
transform 1 0 2312 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5472_6
timestamp 1731220337
transform 1 0 2384 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5471_6
timestamp 1731220337
transform 1 0 2248 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5470_6
timestamp 1731220337
transform 1 0 2288 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5469_6
timestamp 1731220337
transform 1 0 2472 0 -1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5468_6
timestamp 1731220337
transform 1 0 2520 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5467_6
timestamp 1731220337
transform 1 0 2416 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5466_6
timestamp 1731220337
transform 1 0 2328 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5465_6
timestamp 1731220337
transform 1 0 2240 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5464_6
timestamp 1731220337
transform 1 0 2152 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5463_6
timestamp 1731220337
transform 1 0 2552 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5462_6
timestamp 1731220337
transform 1 0 2416 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5461_6
timestamp 1731220337
transform 1 0 2288 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5460_6
timestamp 1731220337
transform 1 0 2168 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5459_6
timestamp 1731220337
transform 1 0 2056 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5458_6
timestamp 1731220337
transform 1 0 2544 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5457_6
timestamp 1731220337
transform 1 0 2384 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5456_6
timestamp 1731220337
transform 1 0 2224 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5455_6
timestamp 1731220337
transform 1 0 2064 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5454_6
timestamp 1731220337
transform 1 0 1920 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5453_6
timestamp 1731220337
transform 1 0 2480 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5452_6
timestamp 1731220337
transform 1 0 2304 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5451_6
timestamp 1731220337
transform 1 0 2128 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5450_6
timestamp 1731220337
transform 1 0 1960 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5449_6
timestamp 1731220337
transform 1 0 1824 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5448_6
timestamp 1731220337
transform 1 0 2280 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5447_6
timestamp 1731220337
transform 1 0 2120 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5446_6
timestamp 1731220337
transform 1 0 1960 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5445_6
timestamp 1731220337
transform 1 0 1824 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5444_6
timestamp 1731220337
transform 1 0 1664 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5443_6
timestamp 1731220337
transform 1 0 1664 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5442_6
timestamp 1731220337
transform 1 0 1568 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5441_6
timestamp 1731220337
transform 1 0 1824 0 -1 508
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5440_6
timestamp 1731220337
transform 1 0 2120 0 -1 508
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5439_6
timestamp 1731220337
transform 1 0 1960 0 -1 508
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5438_6
timestamp 1731220337
transform 1 0 1952 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5437_6
timestamp 1731220337
transform 1 0 1824 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5436_6
timestamp 1731220337
transform 1 0 1664 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5435_6
timestamp 1731220337
transform 1 0 1560 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5434_6
timestamp 1731220337
transform 1 0 1432 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5433_6
timestamp 1731220337
transform 1 0 1304 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5432_6
timestamp 1731220337
transform 1 0 1224 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5431_6
timestamp 1731220337
transform 1 0 1344 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5430_6
timestamp 1731220337
transform 1 0 1456 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5429_6
timestamp 1731220337
transform 1 0 1352 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5428_6
timestamp 1731220337
transform 1 0 1464 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5427_6
timestamp 1731220337
transform 1 0 1576 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5426_6
timestamp 1731220337
transform 1 0 1576 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5425_6
timestamp 1731220337
transform 1 0 1440 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5424_6
timestamp 1731220337
transform 1 0 1304 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5423_6
timestamp 1731220337
transform 1 0 1176 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5422_6
timestamp 1731220337
transform 1 0 1336 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5421_6
timestamp 1731220337
transform 1 0 1496 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5420_6
timestamp 1731220337
transform 1 0 1344 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5419_6
timestamp 1731220337
transform 1 0 1184 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5418_6
timestamp 1731220337
transform 1 0 1128 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5417_6
timestamp 1731220337
transform 1 0 1000 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5416_6
timestamp 1731220337
transform 1 0 1264 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5415_6
timestamp 1731220337
transform 1 0 1328 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5414_6
timestamp 1731220337
transform 1 0 1112 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5413_6
timestamp 1731220337
transform 1 0 872 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5412_6
timestamp 1731220337
transform 1 0 744 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5411_6
timestamp 1731220337
transform 1 0 736 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5410_6
timestamp 1731220337
transform 1 0 880 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5409_6
timestamp 1731220337
transform 1 0 1032 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5408_6
timestamp 1731220337
transform 1 0 1024 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5407_6
timestamp 1731220337
transform 1 0 872 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5406_6
timestamp 1731220337
transform 1 0 1048 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5405_6
timestamp 1731220337
transform 1 0 1176 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5404_6
timestamp 1731220337
transform 1 0 1248 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5403_6
timestamp 1731220337
transform 1 0 1144 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5402_6
timestamp 1731220337
transform 1 0 1104 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5401_6
timestamp 1731220337
transform 1 0 976 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5400_6
timestamp 1731220337
transform 1 0 896 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5399_6
timestamp 1731220337
transform 1 0 1040 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5398_6
timestamp 1731220337
transform 1 0 1176 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5397_6
timestamp 1731220337
transform 1 0 2104 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5396_6
timestamp 1731220337
transform 1 0 2032 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5395_6
timestamp 1731220337
transform 1 0 1920 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5394_6
timestamp 1731220337
transform 1 0 2152 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5393_6
timestamp 1731220337
transform 1 0 2280 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5392_6
timestamp 1731220337
transform 1 0 2416 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5391_6
timestamp 1731220337
transform 1 0 2392 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5390_6
timestamp 1731220337
transform 1 0 2304 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5389_6
timestamp 1731220337
transform 1 0 2216 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5388_6
timestamp 1731220337
transform 1 0 2480 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5387_6
timestamp 1731220337
transform 1 0 2568 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5386_6
timestamp 1731220337
transform 1 0 2632 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5385_6
timestamp 1731220337
transform 1 0 2504 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5384_6
timestamp 1731220337
transform 1 0 2376 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5383_6
timestamp 1731220337
transform 1 0 2256 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5382_6
timestamp 1731220337
transform 1 0 2136 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5381_6
timestamp 1731220337
transform 1 0 2400 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5380_6
timestamp 1731220337
transform 1 0 2288 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5379_6
timestamp 1731220337
transform 1 0 2176 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5378_6
timestamp 1731220337
transform 1 0 2088 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5377_6
timestamp 1731220337
transform 1 0 2000 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5376_6
timestamp 1731220337
transform 1 0 1912 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5375_6
timestamp 1731220337
transform 1 0 1824 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5374_6
timestamp 1731220337
transform 1 0 1664 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5373_6
timestamp 1731220337
transform 1 0 1576 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5372_6
timestamp 1731220337
transform 1 0 1488 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5371_6
timestamp 1731220337
transform 1 0 1400 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5370_6
timestamp 1731220337
transform 1 0 1312 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5369_6
timestamp 1731220337
transform 1 0 1224 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5368_6
timestamp 1731220337
transform 1 0 1136 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5367_6
timestamp 1731220337
transform 1 0 1048 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5366_6
timestamp 1731220337
transform 1 0 960 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5365_6
timestamp 1731220337
transform 1 0 1096 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5364_6
timestamp 1731220337
transform 1 0 1200 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5363_6
timestamp 1731220337
transform 1 0 1304 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5362_6
timestamp 1731220337
transform 1 0 1232 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5361_6
timestamp 1731220337
transform 1 0 1120 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5360_6
timestamp 1731220337
transform 1 0 1016 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5359_6
timestamp 1731220337
transform 1 0 1200 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5358_6
timestamp 1731220337
transform 1 0 1072 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5357_6
timestamp 1731220337
transform 1 0 952 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5356_6
timestamp 1731220337
transform 1 0 832 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5355_6
timestamp 1731220337
transform 1 0 712 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5354_6
timestamp 1731220337
transform 1 0 808 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5353_6
timestamp 1731220337
transform 1 0 912 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5352_6
timestamp 1731220337
transform 1 0 992 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5351_6
timestamp 1731220337
transform 1 0 800 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5350_6
timestamp 1731220337
transform 1 0 704 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5349_6
timestamp 1731220337
transform 1 0 704 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5348_6
timestamp 1731220337
transform 1 0 616 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5347_6
timestamp 1731220337
transform 1 0 896 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5346_6
timestamp 1731220337
transform 1 0 872 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5345_6
timestamp 1731220337
transform 1 0 784 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5344_6
timestamp 1731220337
transform 1 0 696 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5343_6
timestamp 1731220337
transform 1 0 608 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5342_6
timestamp 1731220337
transform 1 0 520 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5341_6
timestamp 1731220337
transform 1 0 432 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5340_6
timestamp 1731220337
transform 1 0 344 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5339_6
timestamp 1731220337
transform 1 0 256 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5338_6
timestamp 1731220337
transform 1 0 440 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5337_6
timestamp 1731220337
transform 1 0 528 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5336_6
timestamp 1731220337
transform 1 0 592 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5335_6
timestamp 1731220337
transform 1 0 480 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5334_6
timestamp 1731220337
transform 1 0 368 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5333_6
timestamp 1731220337
transform 1 0 256 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5332_6
timestamp 1731220337
transform 1 0 592 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5331_6
timestamp 1731220337
transform 1 0 464 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5330_6
timestamp 1731220337
transform 1 0 336 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5329_6
timestamp 1731220337
transform 1 0 216 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5328_6
timestamp 1731220337
transform 1 0 128 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5327_6
timestamp 1731220337
transform 1 0 128 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5326_6
timestamp 1731220337
transform 1 0 248 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5325_6
timestamp 1731220337
transform 1 0 408 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5324_6
timestamp 1731220337
transform 1 0 736 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5323_6
timestamp 1731220337
transform 1 0 576 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5322_6
timestamp 1731220337
transform 1 0 560 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5321_6
timestamp 1731220337
transform 1 0 424 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5320_6
timestamp 1731220337
transform 1 0 296 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5319_6
timestamp 1731220337
transform 1 0 696 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5318_6
timestamp 1731220337
transform 1 0 840 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5317_6
timestamp 1731220337
transform 1 0 808 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5316_6
timestamp 1731220337
transform 1 0 696 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5315_6
timestamp 1731220337
transform 1 0 592 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5314_6
timestamp 1731220337
transform 1 0 1032 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5313_6
timestamp 1731220337
transform 1 0 920 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5312_6
timestamp 1731220337
transform 1 0 920 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5311_6
timestamp 1731220337
transform 1 0 792 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5310_6
timestamp 1731220337
transform 1 0 672 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5309_6
timestamp 1731220337
transform 1 0 552 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5308_6
timestamp 1731220337
transform 1 0 448 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5307_6
timestamp 1731220337
transform 1 0 720 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5306_6
timestamp 1731220337
transform 1 0 568 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5305_6
timestamp 1731220337
transform 1 0 424 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5304_6
timestamp 1731220337
transform 1 0 288 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5303_6
timestamp 1731220337
transform 1 0 160 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5302_6
timestamp 1731220337
transform 1 0 600 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5301_6
timestamp 1731220337
transform 1 0 464 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5300_6
timestamp 1731220337
transform 1 0 336 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5299_6
timestamp 1731220337
transform 1 0 216 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5298_6
timestamp 1731220337
transform 1 0 128 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5297_6
timestamp 1731220337
transform 1 0 128 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5296_6
timestamp 1731220337
transform 1 0 224 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5295_6
timestamp 1731220337
transform 1 0 352 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5294_6
timestamp 1731220337
transform 1 0 480 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5293_6
timestamp 1731220337
transform 1 0 616 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5292_6
timestamp 1731220337
transform 1 0 552 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5291_6
timestamp 1731220337
transform 1 0 408 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5290_6
timestamp 1731220337
transform 1 0 720 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5289_6
timestamp 1731220337
transform 1 0 904 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5288_6
timestamp 1731220337
transform 1 0 1024 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5287_6
timestamp 1731220337
transform 1 0 904 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5286_6
timestamp 1731220337
transform 1 0 784 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5285_6
timestamp 1731220337
transform 1 0 672 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5284_6
timestamp 1731220337
transform 1 0 560 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5283_6
timestamp 1731220337
transform 1 0 912 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5282_6
timestamp 1731220337
transform 1 0 784 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5281_6
timestamp 1731220337
transform 1 0 656 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5280_6
timestamp 1731220337
transform 1 0 536 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5279_6
timestamp 1731220337
transform 1 0 424 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5278_6
timestamp 1731220337
transform 1 0 752 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5277_6
timestamp 1731220337
transform 1 0 616 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5276_6
timestamp 1731220337
transform 1 0 488 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5275_6
timestamp 1731220337
transform 1 0 360 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5274_6
timestamp 1731220337
transform 1 0 240 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5273_6
timestamp 1731220337
transform 1 0 608 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5272_6
timestamp 1731220337
transform 1 0 480 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5271_6
timestamp 1731220337
transform 1 0 352 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5270_6
timestamp 1731220337
transform 1 0 224 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5269_6
timestamp 1731220337
transform 1 0 128 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5268_6
timestamp 1731220337
transform 1 0 544 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5267_6
timestamp 1731220337
transform 1 0 424 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5266_6
timestamp 1731220337
transform 1 0 312 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5265_6
timestamp 1731220337
transform 1 0 216 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5264_6
timestamp 1731220337
transform 1 0 128 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5263_6
timestamp 1731220337
transform 1 0 552 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5262_6
timestamp 1731220337
transform 1 0 392 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5261_6
timestamp 1731220337
transform 1 0 240 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5260_6
timestamp 1731220337
transform 1 0 128 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5259_6
timestamp 1731220337
transform 1 0 128 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5258_6
timestamp 1731220337
transform 1 0 296 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5257_6
timestamp 1731220337
transform 1 0 488 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5256_6
timestamp 1731220337
transform 1 0 368 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5255_6
timestamp 1731220337
transform 1 0 152 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5254_6
timestamp 1731220337
transform 1 0 176 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5253_6
timestamp 1731220337
transform 1 0 320 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5252_6
timestamp 1731220337
transform 1 0 464 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5251_6
timestamp 1731220337
transform 1 0 376 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5250_6
timestamp 1731220337
transform 1 0 272 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5249_6
timestamp 1731220337
transform 1 0 488 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5248_6
timestamp 1731220337
transform 1 0 480 0 1 1620
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5247_6
timestamp 1731220337
transform 1 0 392 0 1 1620
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5246_6
timestamp 1731220337
transform 1 0 432 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5245_6
timestamp 1731220337
transform 1 0 528 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5244_6
timestamp 1731220337
transform 1 0 632 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5243_6
timestamp 1731220337
transform 1 0 624 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5242_6
timestamp 1731220337
transform 1 0 504 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5241_6
timestamp 1731220337
transform 1 0 424 0 -1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5240_6
timestamp 1731220337
transform 1 0 568 0 -1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5239_6
timestamp 1731220337
transform 1 0 720 0 -1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5238_6
timestamp 1731220337
transform 1 0 696 0 1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5237_6
timestamp 1731220337
transform 1 0 552 0 1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5236_6
timestamp 1731220337
transform 1 0 416 0 1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5235_6
timestamp 1731220337
transform 1 0 288 0 1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5234_6
timestamp 1731220337
transform 1 0 632 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5233_6
timestamp 1731220337
transform 1 0 496 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5232_6
timestamp 1731220337
transform 1 0 360 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5231_6
timestamp 1731220337
transform 1 0 232 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5230_6
timestamp 1731220337
transform 1 0 128 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5229_6
timestamp 1731220337
transform 1 0 576 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5228_6
timestamp 1731220337
transform 1 0 456 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5227_6
timestamp 1731220337
transform 1 0 336 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5226_6
timestamp 1731220337
transform 1 0 216 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5225_6
timestamp 1731220337
transform 1 0 128 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5224_6
timestamp 1731220337
transform 1 0 688 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5223_6
timestamp 1731220337
transform 1 0 536 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5222_6
timestamp 1731220337
transform 1 0 384 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5221_6
timestamp 1731220337
transform 1 0 240 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5220_6
timestamp 1731220337
transform 1 0 128 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5219_6
timestamp 1731220337
transform 1 0 128 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5218_6
timestamp 1731220337
transform 1 0 240 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5217_6
timestamp 1731220337
transform 1 0 760 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5216_6
timestamp 1731220337
transform 1 0 576 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5215_6
timestamp 1731220337
transform 1 0 400 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5214_6
timestamp 1731220337
transform 1 0 264 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5213_6
timestamp 1731220337
transform 1 0 144 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5212_6
timestamp 1731220337
transform 1 0 640 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5211_6
timestamp 1731220337
transform 1 0 512 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5210_6
timestamp 1731220337
transform 1 0 384 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5209_6
timestamp 1731220337
transform 1 0 312 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5208_6
timestamp 1731220337
transform 1 0 424 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5207_6
timestamp 1731220337
transform 1 0 648 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5206_6
timestamp 1731220337
transform 1 0 536 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5205_6
timestamp 1731220337
transform 1 0 496 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5204_6
timestamp 1731220337
transform 1 0 408 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5203_6
timestamp 1731220337
transform 1 0 592 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5202_6
timestamp 1731220337
transform 1 0 544 0 1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5201_6
timestamp 1731220337
transform 1 0 728 0 1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5200_6
timestamp 1731220337
transform 1 0 904 0 1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5199_6
timestamp 1731220337
transform 1 0 912 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5198_6
timestamp 1731220337
transform 1 0 800 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5197_6
timestamp 1731220337
transform 1 0 696 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5196_6
timestamp 1731220337
transform 1 0 1032 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5195_6
timestamp 1731220337
transform 1 0 984 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5194_6
timestamp 1731220337
transform 1 0 872 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5193_6
timestamp 1731220337
transform 1 0 760 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5192_6
timestamp 1731220337
transform 1 0 768 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5191_6
timestamp 1731220337
transform 1 0 888 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5190_6
timestamp 1731220337
transform 1 0 944 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5189_6
timestamp 1731220337
transform 1 0 1128 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5188_6
timestamp 1731220337
transform 1 0 1264 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5187_6
timestamp 1731220337
transform 1 0 1136 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5186_6
timestamp 1731220337
transform 1 0 1008 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5185_6
timestamp 1731220337
transform 1 0 1096 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5184_6
timestamp 1731220337
transform 1 0 1208 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5183_6
timestamp 1731220337
transform 1 0 1328 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5182_6
timestamp 1731220337
transform 1 0 1416 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5181_6
timestamp 1731220337
transform 1 0 1288 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5180_6
timestamp 1731220337
transform 1 0 1160 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5179_6
timestamp 1731220337
transform 1 0 1072 0 1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5178_6
timestamp 1731220337
transform 1 0 1232 0 1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5177_6
timestamp 1731220337
transform 1 0 1560 0 1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5176_6
timestamp 1731220337
transform 1 0 1392 0 1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5175_6
timestamp 1731220337
transform 1 0 1344 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5174_6
timestamp 1731220337
transform 1 0 1472 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5173_6
timestamp 1731220337
transform 1 0 1600 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5172_6
timestamp 1731220337
transform 1 0 1600 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5171_6
timestamp 1731220337
transform 1 0 1432 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5170_6
timestamp 1731220337
transform 1 0 1368 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5169_6
timestamp 1731220337
transform 1 0 1664 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5168_6
timestamp 1731220337
transform 1 0 1528 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5167_6
timestamp 1731220337
transform 1 0 1520 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5166_6
timestamp 1731220337
transform 1 0 1664 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5165_6
timestamp 1731220337
transform 1 0 1824 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5164_6
timestamp 1731220337
transform 1 0 1824 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5163_6
timestamp 1731220337
transform 1 0 1992 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5162_6
timestamp 1731220337
transform 1 0 2008 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5161_6
timestamp 1731220337
transform 1 0 1824 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5160_6
timestamp 1731220337
transform 1 0 1824 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5159_6
timestamp 1731220337
transform 1 0 1912 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5158_6
timestamp 1731220337
transform 1 0 2024 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5157_6
timestamp 1731220337
transform 1 0 2288 0 1 3028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5156_6
timestamp 1731220337
transform 1 0 2112 0 1 3028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5155_6
timestamp 1731220337
transform 1 0 1952 0 1 3028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5154_6
timestamp 1731220337
transform 1 0 1824 0 1 3028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5153_6
timestamp 1731220337
transform 1 0 1824 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5152_6
timestamp 1731220337
transform 1 0 2000 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5151_6
timestamp 1731220337
transform 1 0 2392 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5150_6
timestamp 1731220337
transform 1 0 2200 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5149_6
timestamp 1731220337
transform 1 0 2192 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5148_6
timestamp 1731220337
transform 1 0 2040 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5147_6
timestamp 1731220337
transform 1 0 1904 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5146_6
timestamp 1731220337
transform 1 0 2520 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5145_6
timestamp 1731220337
transform 1 0 2352 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5144_6
timestamp 1731220337
transform 1 0 2232 0 -1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5143_6
timestamp 1731220337
transform 1 0 2080 0 -1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5142_6
timestamp 1731220337
transform 1 0 2392 0 -1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5141_6
timestamp 1731220337
transform 1 0 2552 0 -1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5140_6
timestamp 1731220337
transform 1 0 2560 0 1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5139_6
timestamp 1731220337
transform 1 0 2424 0 1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5138_6
timestamp 1731220337
transform 1 0 2288 0 1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5137_6
timestamp 1731220337
transform 1 0 2152 0 1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5136_6
timestamp 1731220337
transform 1 0 2384 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5135_6
timestamp 1731220337
transform 1 0 2264 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5134_6
timestamp 1731220337
transform 1 0 2144 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5133_6
timestamp 1731220337
transform 1 0 2024 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5132_6
timestamp 1731220337
transform 1 0 2304 0 1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5131_6
timestamp 1731220337
transform 1 0 2136 0 1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5130_6
timestamp 1731220337
transform 1 0 1968 0 1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5129_6
timestamp 1731220337
transform 1 0 1824 0 1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5128_6
timestamp 1731220337
transform 1 0 1664 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5127_6
timestamp 1731220337
transform 1 0 1544 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5126_6
timestamp 1731220337
transform 1 0 1400 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5125_6
timestamp 1731220337
transform 1 0 1256 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5124_6
timestamp 1731220337
transform 1 0 1112 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5123_6
timestamp 1731220337
transform 1 0 952 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5122_6
timestamp 1731220337
transform 1 0 1392 0 -1 3436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5121_6
timestamp 1731220337
transform 1 0 1224 0 -1 3436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5120_6
timestamp 1731220337
transform 1 0 1056 0 -1 3436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5119_6
timestamp 1731220337
transform 1 0 888 0 -1 3436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5118_6
timestamp 1731220337
transform 1 0 928 0 1 3300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5117_6
timestamp 1731220337
transform 1 0 1112 0 1 3300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5116_6
timestamp 1731220337
transform 1 0 1288 0 1 3300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5115_6
timestamp 1731220337
transform 1 0 1456 0 1 3300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5114_6
timestamp 1731220337
transform 1 0 1632 0 1 3300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5113_6
timestamp 1731220337
transform 1 0 1664 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5112_6
timestamp 1731220337
transform 1 0 1496 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5111_6
timestamp 1731220337
transform 1 0 1336 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5110_6
timestamp 1731220337
transform 1 0 1168 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5109_6
timestamp 1731220337
transform 1 0 1000 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5108_6
timestamp 1731220337
transform 1 0 1464 0 1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5107_6
timestamp 1731220337
transform 1 0 1296 0 1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5106_6
timestamp 1731220337
transform 1 0 1128 0 1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5105_6
timestamp 1731220337
transform 1 0 960 0 1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5104_6
timestamp 1731220337
transform 1 0 1312 0 -1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5103_6
timestamp 1731220337
transform 1 0 1192 0 -1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5102_6
timestamp 1731220337
transform 1 0 1072 0 -1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5101_6
timestamp 1731220337
transform 1 0 960 0 -1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5100_6
timestamp 1731220337
transform 1 0 840 0 -1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_599_6
timestamp 1731220337
transform 1 0 1136 0 1 3024
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_598_6
timestamp 1731220337
transform 1 0 1048 0 1 3024
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_597_6
timestamp 1731220337
transform 1 0 960 0 1 3024
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_596_6
timestamp 1731220337
transform 1 0 872 0 1 3024
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_595_6
timestamp 1731220337
transform 1 0 936 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_594_6
timestamp 1731220337
transform 1 0 1024 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_593_6
timestamp 1731220337
transform 1 0 1288 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_592_6
timestamp 1731220337
transform 1 0 1200 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_591_6
timestamp 1731220337
transform 1 0 1112 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_590_6
timestamp 1731220337
transform 1 0 1096 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_589_6
timestamp 1731220337
transform 1 0 968 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_588_6
timestamp 1731220337
transform 1 0 1224 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_587_6
timestamp 1731220337
transform 1 0 1352 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_586_6
timestamp 1731220337
transform 1 0 1488 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_585_6
timestamp 1731220337
transform 1 0 1488 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_584_6
timestamp 1731220337
transform 1 0 1336 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_583_6
timestamp 1731220337
transform 1 0 1184 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_582_6
timestamp 1731220337
transform 1 0 1040 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_581_6
timestamp 1731220337
transform 1 0 888 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_580_6
timestamp 1731220337
transform 1 0 1352 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_579_6
timestamp 1731220337
transform 1 0 1184 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_578_6
timestamp 1731220337
transform 1 0 1016 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_577_6
timestamp 1731220337
transform 1 0 848 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_576_6
timestamp 1731220337
transform 1 0 904 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_575_6
timestamp 1731220337
transform 1 0 1208 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_574_6
timestamp 1731220337
transform 1 0 1056 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_573_6
timestamp 1731220337
transform 1 0 976 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_572_6
timestamp 1731220337
transform 1 0 1120 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_571_6
timestamp 1731220337
transform 1 0 1272 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_570_6
timestamp 1731220337
transform 1 0 1216 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_569_6
timestamp 1731220337
transform 1 0 1096 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_568_6
timestamp 1731220337
transform 1 0 984 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_567_6
timestamp 1731220337
transform 1 0 872 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_566_6
timestamp 1731220337
transform 1 0 768 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_565_6
timestamp 1731220337
transform 1 0 672 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_564_6
timestamp 1731220337
transform 1 0 584 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_563_6
timestamp 1731220337
transform 1 0 496 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_562_6
timestamp 1731220337
transform 1 0 848 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_561_6
timestamp 1731220337
transform 1 0 736 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_560_6
timestamp 1731220337
transform 1 0 632 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_559_6
timestamp 1731220337
transform 1 0 544 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_558_6
timestamp 1731220337
transform 1 0 456 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_557_6
timestamp 1731220337
transform 1 0 752 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_556_6
timestamp 1731220337
transform 1 0 608 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_555_6
timestamp 1731220337
transform 1 0 472 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_554_6
timestamp 1731220337
transform 1 0 352 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_553_6
timestamp 1731220337
transform 1 0 240 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_552_6
timestamp 1731220337
transform 1 0 688 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_551_6
timestamp 1731220337
transform 1 0 536 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_550_6
timestamp 1731220337
transform 1 0 384 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_549_6
timestamp 1731220337
transform 1 0 240 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_548_6
timestamp 1731220337
transform 1 0 128 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_547_6
timestamp 1731220337
transform 1 0 128 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_546_6
timestamp 1731220337
transform 1 0 248 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_545_6
timestamp 1731220337
transform 1 0 408 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_544_6
timestamp 1731220337
transform 1 0 728 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_543_6
timestamp 1731220337
transform 1 0 568 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_542_6
timestamp 1731220337
transform 1 0 568 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_541_6
timestamp 1731220337
transform 1 0 440 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_540_6
timestamp 1731220337
transform 1 0 320 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_539_6
timestamp 1731220337
transform 1 0 840 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_538_6
timestamp 1731220337
transform 1 0 704 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_537_6
timestamp 1731220337
transform 1 0 672 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_536_6
timestamp 1731220337
transform 1 0 584 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_535_6
timestamp 1731220337
transform 1 0 496 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_534_6
timestamp 1731220337
transform 1 0 760 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_533_6
timestamp 1731220337
transform 1 0 848 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_532_6
timestamp 1731220337
transform 1 0 784 0 1 3024
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_531_6
timestamp 1731220337
transform 1 0 696 0 1 3024
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_530_6
timestamp 1731220337
transform 1 0 608 0 1 3024
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_529_6
timestamp 1731220337
transform 1 0 520 0 1 3024
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_528_6
timestamp 1731220337
transform 1 0 432 0 1 3024
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_527_6
timestamp 1731220337
transform 1 0 720 0 -1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_526_6
timestamp 1731220337
transform 1 0 600 0 -1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_525_6
timestamp 1731220337
transform 1 0 480 0 -1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_524_6
timestamp 1731220337
transform 1 0 360 0 -1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_523_6
timestamp 1731220337
transform 1 0 800 0 1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_522_6
timestamp 1731220337
transform 1 0 640 0 1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_521_6
timestamp 1731220337
transform 1 0 480 0 1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_520_6
timestamp 1731220337
transform 1 0 320 0 1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_519_6
timestamp 1731220337
transform 1 0 176 0 1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_518_6
timestamp 1731220337
transform 1 0 824 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_517_6
timestamp 1731220337
transform 1 0 640 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_516_6
timestamp 1731220337
transform 1 0 456 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_515_6
timestamp 1731220337
transform 1 0 272 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_514_6
timestamp 1731220337
transform 1 0 128 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_513_6
timestamp 1731220337
transform 1 0 128 0 1 3300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_512_6
timestamp 1731220337
transform 1 0 320 0 1 3300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_511_6
timestamp 1731220337
transform 1 0 736 0 1 3300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_510_6
timestamp 1731220337
transform 1 0 528 0 1 3300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_59_6
timestamp 1731220337
transform 1 0 408 0 -1 3436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_58_6
timestamp 1731220337
transform 1 0 248 0 -1 3436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_57_6
timestamp 1731220337
transform 1 0 128 0 -1 3436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_56_6
timestamp 1731220337
transform 1 0 568 0 -1 3436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_55_6
timestamp 1731220337
transform 1 0 728 0 -1 3436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_54_6
timestamp 1731220337
transform 1 0 784 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_53_6
timestamp 1731220337
transform 1 0 608 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_52_6
timestamp 1731220337
transform 1 0 432 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_51_6
timestamp 1731220337
transform 1 0 264 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_50_6
timestamp 1731220337
transform 1 0 128 0 1 3440
box 8 4 84 60
<< end >>
