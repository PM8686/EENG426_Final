magic
tech sky130l
timestamp 1729066705
<< ndiffusion >>
rect 8 19 13 24
rect 8 16 9 19
rect 12 16 13 19
rect 8 14 13 16
rect 15 18 22 24
rect 15 15 17 18
rect 20 15 22 18
rect 15 14 22 15
rect 24 14 29 24
rect 31 22 36 24
rect 31 19 32 22
rect 35 19 36 22
rect 31 14 36 19
rect 38 19 43 24
rect 38 16 39 19
rect 42 16 43 19
rect 38 14 43 16
rect 45 22 52 24
rect 45 19 47 22
rect 50 19 52 22
rect 45 14 52 19
rect 48 4 52 14
rect 54 16 59 24
rect 54 13 55 16
rect 58 13 59 16
rect 54 4 59 13
rect 61 22 68 24
rect 61 19 63 22
rect 66 19 68 22
rect 61 4 68 19
rect 70 16 75 24
rect 70 13 71 16
rect 74 13 75 16
rect 70 4 75 13
rect 77 15 84 24
rect 77 12 80 15
rect 83 12 84 15
rect 77 4 84 12
rect 86 4 89 24
rect 91 4 94 24
rect 96 22 101 24
rect 96 19 97 22
rect 100 19 101 22
rect 96 18 101 19
rect 103 23 108 24
rect 103 20 104 23
rect 107 20 108 23
rect 103 18 108 20
rect 114 22 119 24
rect 114 19 115 22
rect 118 19 119 22
rect 114 18 119 19
rect 121 23 126 24
rect 121 20 122 23
rect 125 20 126 23
rect 121 18 126 20
rect 96 4 100 18
<< ndc >>
rect 9 16 12 19
rect 17 15 20 18
rect 32 19 35 22
rect 39 16 42 19
rect 47 19 50 22
rect 55 13 58 16
rect 63 19 66 22
rect 71 13 74 16
rect 80 12 83 15
rect 97 19 100 22
rect 104 20 107 23
rect 115 19 118 22
rect 122 20 125 23
<< ntransistor >>
rect 13 14 15 24
rect 22 14 24 24
rect 29 14 31 24
rect 36 14 38 24
rect 43 14 45 24
rect 52 4 54 24
rect 59 4 61 24
rect 68 4 70 24
rect 75 4 77 24
rect 84 4 86 24
rect 89 4 91 24
rect 94 4 96 24
rect 101 18 103 24
rect 119 18 121 24
<< pdiffusion >>
rect 64 67 68 71
rect 48 54 52 67
rect 18 42 22 54
rect 8 36 13 42
rect 8 33 9 36
rect 12 33 13 36
rect 8 31 13 33
rect 15 41 22 42
rect 15 38 16 41
rect 19 38 22 41
rect 15 31 22 38
rect 24 35 29 54
rect 24 32 25 35
rect 28 32 29 35
rect 24 31 29 32
rect 31 41 36 54
rect 31 38 32 41
rect 35 38 36 41
rect 31 31 36 38
rect 38 31 43 54
rect 45 36 52 54
rect 45 33 47 36
rect 50 33 52 36
rect 45 31 52 33
rect 54 42 59 67
rect 54 39 55 42
rect 58 39 59 42
rect 54 31 59 39
rect 61 36 68 67
rect 61 33 63 36
rect 66 33 68 36
rect 61 31 68 33
rect 70 67 74 71
rect 80 67 84 79
rect 70 42 75 67
rect 70 39 71 42
rect 74 39 75 42
rect 70 31 75 39
rect 77 35 84 67
rect 77 32 80 35
rect 83 32 84 35
rect 77 31 84 32
rect 86 31 89 79
rect 91 31 94 79
rect 96 39 100 79
rect 96 36 101 39
rect 96 33 97 36
rect 100 33 101 36
rect 96 31 101 33
rect 103 38 108 39
rect 103 35 104 38
rect 107 35 108 38
rect 103 31 108 35
rect 114 38 119 39
rect 114 35 115 38
rect 118 35 119 38
rect 114 31 119 35
rect 121 36 126 39
rect 121 33 122 36
rect 125 33 126 36
rect 121 31 126 33
<< pdc >>
rect 9 33 12 36
rect 16 38 19 41
rect 25 32 28 35
rect 32 38 35 41
rect 47 33 50 36
rect 55 39 58 42
rect 63 33 66 36
rect 71 39 74 42
rect 80 32 83 35
rect 97 33 100 36
rect 104 35 107 38
rect 115 35 118 38
rect 122 33 125 36
<< ptransistor >>
rect 13 31 15 42
rect 22 31 24 54
rect 29 31 31 54
rect 36 31 38 54
rect 43 31 45 54
rect 52 31 54 67
rect 59 31 61 67
rect 68 31 70 71
rect 75 31 77 67
rect 84 31 86 79
rect 89 31 91 79
rect 94 31 96 79
rect 101 31 103 39
rect 119 31 121 39
<< polysilicon >>
rect 29 89 34 90
rect 29 86 30 89
rect 33 86 34 89
rect 29 85 34 86
rect 43 89 48 90
rect 43 86 44 89
rect 47 86 48 89
rect 43 85 48 86
rect 68 89 73 90
rect 68 86 69 89
rect 72 86 73 89
rect 68 85 73 86
rect 80 89 85 90
rect 80 86 81 89
rect 84 86 85 89
rect 21 81 26 82
rect 21 78 22 81
rect 25 78 26 81
rect 21 77 26 78
rect 13 73 19 74
rect 13 70 15 73
rect 18 70 19 73
rect 13 69 19 70
rect 13 42 15 69
rect 22 54 24 77
rect 29 54 31 85
rect 35 81 40 82
rect 35 78 36 81
rect 39 78 40 81
rect 35 77 40 78
rect 36 54 38 77
rect 43 54 45 85
rect 49 81 54 82
rect 49 78 50 81
rect 53 78 54 81
rect 49 77 54 78
rect 52 67 54 77
rect 57 78 62 79
rect 57 75 58 78
rect 61 75 62 78
rect 57 74 62 75
rect 59 67 61 74
rect 68 71 70 85
rect 80 82 85 86
rect 88 89 93 90
rect 88 86 89 89
rect 92 86 93 89
rect 88 85 93 86
rect 96 89 101 90
rect 96 86 97 89
rect 100 86 101 89
rect 80 80 86 82
rect 84 79 86 80
rect 89 79 91 85
rect 96 82 101 86
rect 94 80 101 82
rect 94 79 96 80
rect 75 67 77 69
rect 101 39 103 41
rect 119 39 121 41
rect 13 24 15 31
rect 22 24 24 31
rect 29 24 31 31
rect 36 24 38 31
rect 43 24 45 31
rect 52 24 54 31
rect 59 24 61 31
rect 68 24 70 31
rect 75 24 77 31
rect 84 24 86 31
rect 89 24 91 31
rect 94 24 96 31
rect 101 24 103 31
rect 119 24 121 31
rect 13 12 15 14
rect 22 12 24 14
rect 29 12 31 14
rect 36 12 38 14
rect 43 12 45 14
rect 52 2 54 4
rect 59 2 61 4
rect 68 2 70 4
rect 75 2 77 4
rect 84 2 86 4
rect 89 2 91 4
rect 94 2 96 4
rect 101 2 103 18
rect 119 16 121 18
rect 116 15 121 16
rect 116 12 117 15
rect 120 12 121 15
rect 116 11 121 12
rect 75 1 80 2
rect 75 -2 76 1
rect 79 -2 80 1
rect 75 -3 80 -2
rect 101 1 106 2
rect 101 -2 102 1
rect 105 -2 106 1
rect 101 -3 106 -2
<< pc >>
rect 30 86 33 89
rect 44 86 47 89
rect 69 86 72 89
rect 81 86 84 89
rect 22 78 25 81
rect 15 70 18 73
rect 36 78 39 81
rect 50 78 53 81
rect 58 75 61 78
rect 89 86 92 89
rect 97 86 100 89
rect 117 12 120 15
rect 76 -2 79 1
rect 102 -2 105 1
<< m1 >>
rect 8 89 12 90
rect 8 86 9 89
rect 8 64 12 86
rect 30 89 33 90
rect 30 85 33 86
rect 44 89 47 90
rect 44 85 47 86
rect 69 89 72 90
rect 69 85 72 86
rect 81 89 84 90
rect 22 81 25 82
rect 22 77 25 78
rect 36 81 39 82
rect 36 77 39 78
rect 50 81 53 82
rect 64 81 68 82
rect 50 77 53 78
rect 58 78 61 79
rect 15 73 18 74
rect 15 69 18 70
rect 58 73 61 75
rect 58 69 61 70
rect 67 78 68 81
rect 64 64 68 78
rect 72 73 76 74
rect 75 70 76 73
rect 72 64 76 70
rect 81 73 84 86
rect 89 89 92 90
rect 89 81 92 86
rect 97 89 100 90
rect 97 85 100 86
rect 81 69 84 70
rect 8 36 12 44
rect 15 38 16 41
rect 19 38 32 41
rect 35 38 36 41
rect 54 39 55 42
rect 58 39 71 42
rect 74 39 75 42
rect 104 38 108 44
rect 8 33 9 36
rect 47 36 50 37
rect 97 36 100 37
rect 8 32 12 33
rect 24 32 25 35
rect 28 32 29 35
rect 62 33 63 36
rect 66 33 67 36
rect 80 35 83 36
rect 47 32 50 33
rect 97 32 100 33
rect 107 35 108 38
rect 9 19 12 20
rect 9 15 12 16
rect 9 11 12 12
rect 17 18 20 19
rect 17 1 20 15
rect 17 -3 20 -2
rect 24 1 29 32
rect 32 22 35 23
rect 47 22 50 23
rect 32 8 35 19
rect 39 19 42 20
rect 62 19 63 22
rect 66 19 67 22
rect 47 18 50 19
rect 39 15 42 16
rect 54 13 55 16
rect 58 13 71 16
rect 74 13 75 16
rect 80 15 83 32
rect 104 23 108 35
rect 112 38 118 44
rect 112 35 115 38
rect 112 29 118 35
rect 122 36 125 37
rect 122 32 125 33
rect 112 26 125 29
rect 122 23 125 26
rect 97 22 100 23
rect 107 20 108 23
rect 104 19 108 20
rect 115 22 118 23
rect 122 19 125 20
rect 97 18 100 19
rect 115 18 118 19
rect 39 11 42 12
rect 116 12 117 15
rect 120 12 121 15
rect 80 11 83 12
rect 32 4 36 8
rect 24 -2 25 1
rect 28 -2 29 1
rect 75 -2 76 1
rect 79 -2 80 1
rect 101 -2 102 1
rect 105 -2 106 1
rect 24 -3 29 -2
<< m2c >>
rect 9 86 12 89
rect 30 86 33 89
rect 44 86 47 89
rect 69 86 72 89
rect 22 78 25 81
rect 36 78 39 81
rect 50 78 53 81
rect 15 70 18 73
rect 58 70 61 73
rect 64 78 67 81
rect 72 70 75 73
rect 97 86 100 89
rect 89 78 92 81
rect 81 70 84 73
rect 9 33 12 36
rect 47 33 50 36
rect 63 33 66 36
rect 97 33 100 36
rect 9 12 12 15
rect 17 -2 20 1
rect 32 19 35 22
rect 47 19 50 22
rect 63 19 66 22
rect 39 12 42 15
rect 122 33 125 36
rect 97 19 100 22
rect 115 19 118 22
rect 80 12 83 15
rect 117 12 120 15
rect 25 -2 28 1
rect 76 -2 79 1
rect 102 -2 105 1
<< m2 >>
rect 8 89 101 90
rect 8 86 9 89
rect 12 86 30 89
rect 33 86 44 89
rect 47 86 69 89
rect 72 86 97 89
rect 100 86 101 89
rect 8 85 101 86
rect 21 81 93 82
rect 21 78 22 81
rect 25 78 36 81
rect 39 78 50 81
rect 53 78 64 81
rect 67 78 89 81
rect 92 78 93 81
rect 21 77 93 78
rect 14 73 85 74
rect 14 70 15 73
rect 18 70 58 73
rect 61 70 72 73
rect 75 70 81 73
rect 84 70 85 73
rect 14 69 85 70
rect 8 36 126 37
rect 8 33 9 36
rect 12 33 47 36
rect 50 33 63 36
rect 66 33 97 36
rect 100 33 122 36
rect 125 33 126 36
rect 8 32 126 33
rect 31 22 119 23
rect 31 19 32 22
rect 35 19 47 22
rect 50 19 63 22
rect 66 19 97 22
rect 100 19 115 22
rect 118 19 119 22
rect 31 18 119 19
rect 8 15 43 16
rect 8 12 9 15
rect 12 12 39 15
rect 42 12 43 15
rect 8 11 43 12
rect 79 15 121 16
rect 79 12 80 15
rect 83 12 117 15
rect 120 12 121 15
rect 79 11 121 12
rect 16 1 106 2
rect 16 -2 17 1
rect 20 -2 25 1
rect 28 -2 76 1
rect 79 -2 102 1
rect 105 -2 106 1
rect 16 -3 106 -2
<< labels >>
rlabel pdiffusion 104 32 104 32 3 YC
rlabel pdiffusion 97 32 97 32 3 Vdd
rlabel polysilicon 102 25 102 25 3 _YC
rlabel polysilicon 102 30 102 30 3 _YC
rlabel polysilicon 95 25 95 25 3 A
rlabel polysilicon 95 30 95 30 3 A
rlabel polysilicon 90 25 90 25 3 B
rlabel polysilicon 90 30 90 30 3 B
rlabel pdiffusion 78 32 78 32 3 _YS
rlabel polysilicon 85 25 85 25 3 C
rlabel polysilicon 85 30 85 30 3 C
rlabel ndiffusion 104 19 104 19 3 YC
rlabel pdiffusion 71 32 71 32 3 #12
rlabel polysilicon 76 25 76 25 3 _YC
rlabel polysilicon 76 30 76 30 3 _YC
rlabel ndiffusion 97 5 97 5 3 GND
rlabel polysilicon 69 25 69 25 3 A
rlabel polysilicon 69 30 69 30 3 A
rlabel pdiffusion 62 32 62 32 3 Vdd
rlabel polysilicon 60 25 60 25 3 C
rlabel polysilicon 60 30 60 30 3 C
rlabel pdiffusion 55 32 55 32 3 #12
rlabel polysilicon 53 25 53 25 3 B
rlabel polysilicon 53 30 53 30 3 B
rlabel pdiffusion 46 32 46 32 3 Vdd
rlabel ndiffusion 78 5 78 5 3 _YS
rlabel ndiffusion 46 15 46 15 3 GND
rlabel polysilicon 44 25 44 25 3 A
rlabel polysilicon 44 30 44 30 3 A
rlabel ndiffusion 71 5 71 5 3 #15
rlabel ndiffusion 39 15 39 15 3 #3
rlabel polysilicon 37 25 37 25 3 B
rlabel polysilicon 37 30 37 30 3 B
rlabel pdiffusion 32 32 32 32 3 #8
rlabel ndiffusion 62 5 62 5 3 GND
rlabel ndiffusion 32 15 32 15 3 GND
rlabel polysilicon 30 25 30 25 3 A
rlabel polysilicon 30 30 30 30 3 A
rlabel pdiffusion 25 32 25 32 3 _YC
rlabel ndiffusion 55 5 55 5 3 #15
rlabel polysilicon 23 25 23 25 3 B
rlabel polysilicon 23 30 23 30 3 B
rlabel ndiffusion 16 15 16 15 3 _YC
rlabel pdiffusion 16 32 16 32 3 #8
rlabel polysilicon 14 25 14 25 3 C
rlabel polysilicon 14 30 14 30 3 C
rlabel ndiffusion 9 15 9 15 3 #3
rlabel ndiffusion 122 19 122 19 3 YS
rlabel pdiffusion 122 32 122 32 3 Vdd
rlabel polysilicon 120 25 120 25 3 _YS
rlabel polysilicon 120 30 120 30 3 _YS
rlabel ndiffusion 115 19 115 19 3 GND
rlabel pdiffusion 115 32 115 32 3 YS
rlabel m2 9 32 9 32 3 Vdd
rlabel m1 33 5 33 5 3 GND
rlabel m2 32 19 32 19 3 GND
rlabel m1 9 41 9 41 3 Vdd
rlabel m1 113 41 113 41 3 YS
rlabel m1 105 41 105 41 3 YC
rlabel m1 73 65 73 65 3 C
rlabel m1 65 65 65 65 3 B
rlabel m1 9 65 9 65 3 A
<< end >>
