magic
tech sky130l
timestamp 1731220596
<< m1 >>
rect 216 3607 220 3631
rect 208 3571 212 3591
rect 296 3571 300 3591
rect 384 3571 388 3591
rect 472 3571 476 3591
rect 1968 3531 1972 3555
rect 2056 3531 2060 3555
rect 2144 3531 2148 3555
rect 2232 3531 2236 3555
rect 2312 3531 2316 3555
rect 2424 3531 2428 3555
rect 2528 3531 2532 3555
rect 2720 3531 2724 3555
rect 2816 3531 2820 3555
rect 2912 3531 2916 3555
rect 3008 3531 3012 3555
rect 3112 3531 3116 3555
rect 368 3471 372 3495
rect 496 3471 500 3495
rect 856 3471 860 3495
rect 1072 3471 1076 3495
rect 1168 3471 1172 3495
rect 1264 3471 1268 3495
rect 1360 3471 1364 3495
rect 1464 3471 1468 3495
rect 1568 3471 1572 3495
rect 2168 3495 2172 3515
rect 2440 3495 2444 3515
rect 2640 3491 2644 3527
rect 824 3431 828 3467
rect 1024 3379 1028 3455
rect 2016 3387 2020 3411
rect 2536 3387 2540 3459
rect 3024 3387 3028 3411
rect 3184 3387 3188 3411
rect 3352 3387 3356 3411
rect 256 3335 260 3359
rect 400 3335 404 3359
rect 560 3335 564 3359
rect 720 3335 724 3359
rect 1040 3335 1044 3359
rect 1360 3335 1364 3359
rect 1512 3335 1516 3359
rect 272 3295 276 3315
rect 408 3295 412 3315
rect 552 3295 556 3315
rect 720 3295 724 3315
rect 896 3291 900 3331
rect 1520 3319 1524 3359
rect 1880 3287 1884 3363
rect 2112 3343 2116 3363
rect 2264 3343 2268 3363
rect 2464 3343 2468 3363
rect 2800 3339 2804 3363
rect 3104 3343 3108 3363
rect 3264 3343 3268 3363
rect 3416 3343 3420 3363
rect 488 3191 492 3259
rect 496 3191 500 3215
rect 632 3191 636 3215
rect 776 3191 780 3215
rect 1088 3191 1092 3215
rect 1408 3191 1412 3259
rect 2456 3243 2460 3267
rect 2624 3243 2628 3267
rect 3472 3243 3476 3267
rect 1568 3191 1572 3215
rect 2808 3199 2812 3219
rect 512 3147 516 3167
rect 648 3147 652 3167
rect 752 3147 756 3167
rect 896 3147 900 3167
rect 1200 3147 1204 3187
rect 1208 3143 1212 3167
rect 656 3039 660 3063
rect 776 3039 780 3063
rect 896 3039 900 3063
rect 1024 3039 1028 3063
rect 1104 3023 1108 3063
rect 1280 3039 1284 3063
rect 1416 3039 1420 3063
rect 1552 3039 1556 3127
rect 2040 3095 2044 3119
rect 2344 3095 2348 3119
rect 2504 3095 2508 3119
rect 2672 3095 2676 3119
rect 3176 3095 3180 3119
rect 3472 3095 3476 3179
rect 1688 3039 1692 3063
rect 1896 3047 1900 3091
rect 664 2995 668 3019
rect 1040 2995 1044 3019
rect 1568 2995 1572 3019
rect 2264 2991 2268 3071
rect 2848 3051 2852 3071
rect 2152 2947 2156 2971
rect 2280 2947 2284 2971
rect 2528 2947 2532 2971
rect 2656 2947 2660 2971
rect 2800 2947 2804 2971
rect 2960 2947 2964 2971
rect 3064 2947 3068 2971
rect 3312 2947 3316 2971
rect 3472 2947 3476 3031
rect 776 2899 780 2923
rect 872 2883 876 2939
rect 912 2899 916 2923
rect 1176 2899 1180 2923
rect 1296 2899 1300 2923
rect 1408 2899 1412 2923
rect 1520 2899 1524 2923
rect 1720 2899 1724 2923
rect 2032 2899 2036 2943
rect 1072 2859 1076 2879
rect 1208 2859 1212 2879
rect 1344 2859 1348 2879
rect 288 2751 292 2775
rect 416 2751 420 2839
rect 1880 2803 1884 2883
rect 2664 2847 2668 2923
rect 3152 2847 3156 2923
rect 2016 2803 2020 2827
rect 2352 2803 2356 2827
rect 2512 2803 2516 2827
rect 2800 2803 2804 2827
rect 2928 2803 2932 2827
rect 552 2751 556 2775
rect 944 2751 948 2775
rect 1072 2751 1076 2775
rect 1200 2751 1204 2775
rect 1336 2751 1340 2775
rect 1968 2763 1972 2787
rect 2200 2763 2204 2799
rect 3048 2791 3052 2827
rect 3472 2803 3476 2883
rect 2856 2767 2860 2787
rect 3176 2767 3180 2787
rect 416 2707 420 2727
rect 544 2707 548 2727
rect 552 2703 556 2735
rect 128 2603 132 2687
rect 688 2647 692 2727
rect 832 2707 836 2727
rect 976 2707 980 2727
rect 984 2703 988 2739
rect 1880 2643 1884 2687
rect 2040 2663 2044 2747
rect 3184 2727 3188 2747
rect 2352 2663 2356 2687
rect 2488 2663 2492 2687
rect 3096 2663 3100 2687
rect 224 2603 228 2627
rect 344 2603 348 2627
rect 464 2603 468 2627
rect 792 2603 796 2627
rect 896 2603 900 2627
rect 992 2603 996 2627
rect 1096 2603 1100 2627
rect 1200 2603 1204 2627
rect 1304 2603 1308 2627
rect 1960 2619 1964 2639
rect 128 2463 132 2543
rect 1880 2499 1884 2539
rect 1984 2515 1988 2599
rect 2104 2559 2108 2639
rect 2184 2619 2188 2639
rect 2720 2619 2724 2639
rect 2824 2619 2828 2639
rect 2832 2615 2836 2647
rect 2584 2515 2588 2539
rect 2704 2515 2708 2539
rect 2824 2515 2828 2539
rect 272 2463 276 2487
rect 424 2463 428 2487
rect 432 2451 436 2487
rect 1000 2463 1004 2487
rect 1136 2463 1140 2487
rect 1272 2463 1276 2487
rect 1960 2475 1964 2495
rect 1064 2427 1068 2447
rect 1200 2427 1204 2447
rect 1336 2427 1340 2447
rect 2168 2419 2172 2495
rect 2256 2475 2260 2495
rect 2552 2475 2556 2495
rect 2688 2475 2692 2495
rect 2816 2475 2820 2495
rect 2944 2475 2948 2495
rect 2792 2375 2796 2399
rect 2944 2375 2948 2399
rect 3104 2375 3108 2399
rect 512 2315 516 2339
rect 1280 2315 1284 2339
rect 2008 2335 2012 2355
rect 2328 2335 2332 2355
rect 2472 2335 2476 2371
rect 2768 2335 2772 2355
rect 2896 2335 2900 2355
rect 3016 2335 3020 2355
rect 3136 2335 3140 2355
rect 776 2271 780 2291
rect 928 2271 932 2311
rect 1248 2271 1252 2291
rect 1392 2271 1396 2291
rect 1528 2271 1532 2291
rect 1664 2271 1668 2291
rect 2136 2231 2140 2299
rect 3264 2275 3268 2355
rect 3384 2335 3388 2355
rect 3464 2335 3468 2355
rect 2472 2231 2476 2255
rect 2632 2231 2636 2255
rect 2912 2231 2916 2255
rect 3032 2231 3036 2255
rect 3472 2231 3476 2315
rect 2088 2195 2092 2215
rect 2240 2195 2244 2215
rect 2808 2191 2812 2215
rect 3288 2195 3292 2215
rect 3368 2195 3372 2227
rect 712 2163 716 2187
rect 888 2163 892 2187
rect 1064 2163 1068 2187
rect 1400 2163 1404 2187
rect 1568 2163 1572 2187
rect 1720 2163 1724 2187
rect 560 2127 564 2147
rect 688 2127 692 2147
rect 824 2127 828 2147
rect 968 2127 972 2147
rect 1256 2127 1260 2147
rect 1400 2095 1404 2119
rect 1984 2071 1988 2111
rect 2464 2087 2468 2111
rect 2608 2087 2612 2111
rect 2752 2087 2756 2111
rect 3472 2087 3476 2175
rect 424 2023 428 2047
rect 544 2023 548 2047
rect 672 2023 676 2047
rect 792 2023 796 2047
rect 1032 2023 1036 2047
rect 1136 2015 1140 2047
rect 2064 2047 2068 2067
rect 2392 2043 2396 2067
rect 2552 2043 2556 2067
rect 2840 2047 2844 2067
rect 3104 2047 3108 2067
rect 3224 2047 3228 2083
rect 3232 2043 3236 2075
rect 248 1983 252 2003
rect 360 1983 364 2003
rect 480 1983 484 2003
rect 600 1983 604 2003
rect 608 1979 612 2011
rect 1200 1983 1204 2003
rect 2192 1947 2196 2011
rect 2536 1947 2540 1971
rect 2864 1947 2868 1971
rect 3024 1947 3028 2027
rect 216 1879 220 1903
rect 344 1879 348 1903
rect 488 1879 492 1903
rect 648 1879 652 1903
rect 832 1879 836 1947
rect 1008 1879 1012 1903
rect 1240 1879 1244 1903
rect 1256 1867 1260 1875
rect 1248 1863 1260 1867
rect 648 1831 652 1855
rect 1120 1835 1124 1855
rect 1248 1835 1252 1863
rect 1456 1859 1460 1903
rect 2056 1903 2060 1923
rect 2064 1899 2068 1931
rect 1328 1835 1332 1855
rect 2352 1795 2356 1819
rect 2616 1795 2620 1819
rect 2736 1795 2740 1819
rect 2856 1795 2860 1819
rect 2984 1795 2988 1819
rect 296 1723 300 1747
rect 568 1723 572 1747
rect 840 1707 844 1763
rect 2632 1751 2636 1775
rect 2824 1755 2828 1775
rect 2928 1755 2932 1775
rect 3032 1755 3036 1775
rect 3152 1755 3156 1775
rect 864 1723 868 1747
rect 1208 1723 1212 1747
rect 1520 1715 1524 1747
rect 1528 1707 1532 1747
rect 1696 1707 1700 1747
rect 128 1619 132 1703
rect 600 1679 604 1703
rect 1264 1679 1268 1703
rect 2360 1651 2364 1675
rect 2488 1651 2492 1675
rect 2616 1651 2620 1675
rect 2752 1651 2756 1675
rect 3008 1651 3012 1675
rect 3240 1651 3244 1675
rect 440 1575 444 1599
rect 624 1575 628 1599
rect 768 1563 772 1615
rect 808 1575 812 1599
rect 1264 1563 1268 1615
rect 1296 1575 1300 1599
rect 1592 1575 1596 1599
rect 1720 1575 1724 1647
rect 2216 1611 2220 1631
rect 2432 1611 2436 1631
rect 2616 1611 2620 1631
rect 2624 1607 2628 1639
rect 3352 1635 3356 1691
rect 3360 1651 3364 1675
rect 3472 1635 3476 1675
rect 2952 1611 2956 1631
rect 3272 1607 3276 1631
rect 2448 1511 2452 1535
rect 2784 1511 2788 1535
rect 2944 1511 2948 1535
rect 3104 1511 3108 1591
rect 3264 1511 3268 1535
rect 464 1435 468 1459
rect 600 1435 604 1459
rect 704 1415 708 1475
rect 1960 1467 1964 1487
rect 2336 1463 2340 1487
rect 2616 1467 2620 1487
rect 3192 1467 3196 1487
rect 736 1435 740 1459
rect 1224 1415 1228 1459
rect 528 1391 532 1411
rect 880 1391 884 1411
rect 984 1391 988 1411
rect 1080 1391 1084 1411
rect 1288 1391 1292 1411
rect 320 1287 324 1311
rect 688 1287 692 1371
rect 1880 1347 1884 1387
rect 2064 1363 2068 1447
rect 2800 1363 2804 1447
rect 3024 1363 3028 1387
rect 1960 1323 1964 1343
rect 2048 1323 2052 1343
rect 2168 1323 2172 1343
rect 2192 1319 2196 1359
rect 2432 1323 2436 1343
rect 2600 1323 2604 1343
rect 2776 1323 2780 1343
rect 2968 1323 2972 1343
rect 3368 1323 3372 1507
rect 3472 1363 3476 1447
rect 1000 1275 1004 1311
rect 288 1251 292 1271
rect 440 1251 444 1271
rect 584 1251 588 1271
rect 760 1251 764 1271
rect 1072 1251 1076 1271
rect 1224 1251 1228 1271
rect 1368 1251 1372 1271
rect 1576 1251 1580 1271
rect 2136 1195 2140 1235
rect 2328 1211 2332 1235
rect 2680 1211 2684 1235
rect 2848 1211 2852 1235
rect 3032 1211 3036 1235
rect 3224 1211 3228 1235
rect 2216 1171 2220 1191
rect 680 1143 684 1167
rect 2224 1167 2228 1199
rect 128 1051 132 1127
rect 216 1107 220 1127
rect 360 1107 364 1139
rect 1392 1131 1396 1167
rect 752 1107 756 1127
rect 1120 1107 1124 1127
rect 1496 1107 1500 1127
rect 1656 1107 1660 1127
rect 3312 1103 3316 1191
rect 424 1007 428 1031
rect 576 1007 580 1031
rect 728 1007 732 1031
rect 1376 1007 1380 1031
rect 1656 1007 1660 1031
rect 1720 1007 1724 1087
rect 2080 1059 2084 1083
rect 2224 1059 2228 1083
rect 2528 1059 2532 1083
rect 2832 1059 2836 1083
rect 2984 1059 2988 1083
rect 3144 1059 3148 1083
rect 3472 1059 3476 1151
rect 2392 1011 2396 1055
rect 2424 1007 2428 1031
rect 2776 1011 2780 1031
rect 2944 1011 2948 1031
rect 3088 1011 3092 1031
rect 3328 1007 3332 1055
rect 128 903 132 987
rect 216 967 220 987
rect 224 963 228 1003
rect 536 963 540 987
rect 728 963 732 987
rect 1080 967 1084 987
rect 1400 967 1404 987
rect 600 859 604 947
rect 768 859 772 883
rect 1392 859 1396 883
rect 128 763 132 843
rect 208 823 212 855
rect 376 823 380 843
rect 544 823 548 843
rect 720 823 724 843
rect 1048 823 1052 855
rect 1480 847 1484 883
rect 1544 859 1548 931
rect 2064 907 2068 931
rect 2448 907 2452 931
rect 2624 907 2628 931
rect 2944 907 2948 931
rect 3088 907 3092 931
rect 3224 907 3228 931
rect 3360 907 3364 931
rect 3472 907 3476 991
rect 2104 859 2108 883
rect 2288 859 2292 903
rect 1408 819 1412 843
rect 1880 755 1884 843
rect 3352 799 3356 883
rect 2064 755 2068 779
rect 2440 755 2444 779
rect 2616 755 2620 779
rect 2936 755 2940 779
rect 3080 755 3084 779
rect 3352 755 3356 779
rect 432 703 436 743
rect 1080 719 1084 743
rect 1384 719 1388 743
rect 1544 719 1548 743
rect 1984 719 1988 739
rect 2712 719 2716 739
rect 3240 719 3244 739
rect 128 615 132 699
rect 944 675 948 715
rect 1104 615 1108 699
rect 136 467 140 551
rect 232 531 236 551
rect 296 527 300 567
rect 448 555 452 595
rect 1112 571 1116 595
rect 1264 571 1268 659
rect 1880 599 1884 639
rect 2344 615 2348 639
rect 2472 615 2476 639
rect 2760 615 2764 639
rect 2928 615 2932 699
rect 3112 615 3116 639
rect 1408 571 1412 595
rect 1552 571 1556 595
rect 1704 571 1708 595
rect 2128 575 2132 595
rect 2488 571 2492 595
rect 2912 575 2916 595
rect 3088 575 3092 595
rect 3176 571 3180 603
rect 3464 571 3468 751
rect 3472 743 3476 843
rect 3472 615 3476 699
rect 552 531 556 551
rect 704 531 708 551
rect 1256 531 1260 551
rect 1376 531 1380 551
rect 2272 467 2276 491
rect 2480 467 2484 555
rect 2624 467 2628 491
rect 2800 467 2804 491
rect 2984 467 2988 491
rect 3176 467 3180 491
rect 248 423 252 447
rect 552 423 556 447
rect 1000 423 1004 447
rect 1232 423 1236 447
rect 1336 423 1340 447
rect 1536 423 1540 447
rect 1632 423 1636 447
rect 1712 423 1716 447
rect 2120 423 2124 463
rect 2128 419 2132 443
rect 2480 423 2484 443
rect 2680 423 2684 443
rect 2896 423 2900 443
rect 3080 423 3084 443
rect 216 387 220 407
rect 392 315 396 407
rect 800 387 804 407
rect 1152 387 1156 407
rect 1536 387 1540 407
rect 216 271 220 295
rect 304 271 308 295
rect 392 271 396 295
rect 568 271 572 295
rect 656 271 660 295
rect 744 255 748 295
rect 1008 271 1012 295
rect 1376 271 1380 295
rect 1472 271 1476 295
rect 824 231 828 251
rect 912 231 916 251
rect 920 227 924 259
rect 1552 255 1556 295
rect 1664 271 1668 351
rect 1880 323 1884 403
rect 3424 367 3428 463
rect 1968 323 1972 347
rect 2056 323 2060 347
rect 2144 323 2148 347
rect 2352 323 2356 347
rect 2840 323 2844 347
rect 3024 323 3028 347
rect 1960 287 1964 307
rect 2048 287 2052 307
rect 2136 287 2140 307
rect 2224 287 2228 307
rect 2424 287 2428 307
rect 2760 287 2764 307
rect 2872 287 2876 307
rect 2984 287 2988 307
rect 3104 287 3108 307
rect 1088 231 1092 251
rect 1176 231 1180 251
rect 1616 231 1620 251
rect 1968 187 1972 211
rect 2056 187 2060 211
rect 2144 187 2148 211
rect 2256 187 2260 211
rect 2392 187 2396 211
rect 2528 187 2532 211
rect 2672 187 2676 211
rect 2944 187 2948 211
rect 3080 187 3084 211
rect 3216 187 3220 211
rect 3472 143 3476 211
rect 2848 119 2852 139
rect 2936 119 2940 139
rect 3024 119 3028 139
rect 3112 119 3116 139
rect 3200 119 3204 139
rect 3288 119 3292 139
<< m2c >>
rect 216 3631 220 3635
rect 216 3603 220 3607
rect 224 3603 228 3607
rect 136 3591 140 3595
rect 208 3591 212 3595
rect 224 3591 228 3595
rect 296 3591 300 3595
rect 312 3591 316 3595
rect 384 3591 388 3595
rect 400 3591 404 3595
rect 472 3591 476 3595
rect 488 3591 492 3595
rect 208 3567 212 3571
rect 296 3567 300 3571
rect 384 3567 388 3571
rect 472 3567 476 3571
rect 1968 3555 1972 3559
rect 2056 3555 2060 3559
rect 2144 3555 2148 3559
rect 2232 3555 2236 3559
rect 2312 3555 2316 3559
rect 2424 3555 2428 3559
rect 2528 3555 2532 3559
rect 2720 3555 2724 3559
rect 2816 3555 2820 3559
rect 2912 3555 2916 3559
rect 3008 3555 3012 3559
rect 3112 3555 3116 3559
rect 1888 3527 1892 3531
rect 1968 3527 1972 3531
rect 1976 3527 1980 3531
rect 2056 3527 2060 3531
rect 2064 3527 2068 3531
rect 2144 3527 2148 3531
rect 2152 3527 2156 3531
rect 2232 3527 2236 3531
rect 2240 3527 2244 3531
rect 2312 3527 2316 3531
rect 2328 3527 2332 3531
rect 2424 3527 2428 3531
rect 2432 3527 2436 3531
rect 2528 3527 2532 3531
rect 2536 3527 2540 3531
rect 2632 3527 2636 3531
rect 2640 3527 2644 3531
rect 2720 3527 2724 3531
rect 2728 3527 2732 3531
rect 2816 3527 2820 3531
rect 2824 3527 2828 3531
rect 2912 3527 2916 3531
rect 2920 3527 2924 3531
rect 3008 3527 3012 3531
rect 3016 3527 3020 3531
rect 3112 3527 3116 3531
rect 3120 3527 3124 3531
rect 3224 3527 3228 3531
rect 1888 3515 1892 3519
rect 1976 3515 1980 3519
rect 2096 3515 2100 3519
rect 2168 3515 2172 3519
rect 2224 3515 2228 3519
rect 2360 3515 2364 3519
rect 2440 3515 2444 3519
rect 2504 3515 2508 3519
rect 368 3495 372 3499
rect 496 3495 500 3499
rect 856 3495 860 3499
rect 1072 3495 1076 3499
rect 1168 3495 1172 3499
rect 1264 3495 1268 3499
rect 1360 3495 1364 3499
rect 1464 3495 1468 3499
rect 1568 3495 1572 3499
rect 2168 3491 2172 3495
rect 2440 3491 2444 3495
rect 2648 3515 2652 3519
rect 2784 3515 2788 3519
rect 2928 3515 2932 3519
rect 3072 3515 3076 3519
rect 3216 3515 3220 3519
rect 2640 3487 2644 3491
rect 248 3467 252 3471
rect 368 3467 372 3471
rect 376 3467 380 3471
rect 496 3467 500 3471
rect 504 3467 508 3471
rect 624 3467 628 3471
rect 744 3467 748 3471
rect 824 3467 828 3471
rect 856 3467 860 3471
rect 864 3467 868 3471
rect 976 3467 980 3471
rect 1072 3467 1076 3471
rect 1080 3467 1084 3471
rect 1168 3467 1172 3471
rect 1176 3467 1180 3471
rect 1264 3467 1268 3471
rect 1272 3467 1276 3471
rect 1360 3467 1364 3471
rect 1368 3467 1372 3471
rect 1464 3467 1468 3471
rect 1472 3467 1476 3471
rect 1568 3467 1572 3471
rect 1576 3467 1580 3471
rect 168 3455 172 3459
rect 296 3455 300 3459
rect 440 3455 444 3459
rect 584 3455 588 3459
rect 736 3455 740 3459
rect 2536 3459 2540 3463
rect 2552 3459 2556 3463
rect 888 3455 892 3459
rect 1024 3455 1028 3459
rect 1032 3455 1036 3459
rect 1176 3455 1180 3459
rect 1320 3455 1324 3459
rect 1472 3455 1476 3459
rect 824 3427 828 3431
rect 2016 3411 2020 3415
rect 1224 3399 1228 3403
rect 3024 3411 3028 3415
rect 3184 3411 3188 3415
rect 3352 3411 3356 3415
rect 1888 3383 1892 3387
rect 2016 3383 2020 3387
rect 2024 3383 2028 3387
rect 2192 3383 2196 3387
rect 2368 3383 2372 3387
rect 2536 3383 2540 3387
rect 2544 3383 2548 3387
rect 2712 3383 2716 3387
rect 2872 3383 2876 3387
rect 3024 3383 3028 3387
rect 3032 3383 3036 3387
rect 3184 3383 3188 3387
rect 3192 3383 3196 3387
rect 3352 3383 3356 3387
rect 3360 3383 3364 3387
rect 1024 3375 1028 3379
rect 1880 3363 1884 3367
rect 1888 3363 1892 3367
rect 2024 3363 2028 3367
rect 2112 3363 2116 3367
rect 2192 3363 2196 3367
rect 2264 3363 2268 3367
rect 2368 3363 2372 3367
rect 2464 3363 2468 3367
rect 2544 3363 2548 3367
rect 2712 3363 2716 3367
rect 2800 3363 2804 3367
rect 2872 3363 2876 3367
rect 3032 3363 3036 3367
rect 3104 3363 3108 3367
rect 3184 3363 3188 3367
rect 3264 3363 3268 3367
rect 3336 3363 3340 3367
rect 3416 3363 3420 3367
rect 3480 3363 3484 3367
rect 256 3359 260 3363
rect 400 3359 404 3363
rect 560 3359 564 3363
rect 720 3359 724 3363
rect 1040 3359 1044 3363
rect 1360 3359 1364 3363
rect 1512 3359 1516 3363
rect 136 3331 140 3335
rect 256 3331 260 3335
rect 264 3331 268 3335
rect 400 3331 404 3335
rect 408 3331 412 3335
rect 560 3331 564 3335
rect 568 3331 572 3335
rect 720 3331 724 3335
rect 728 3331 732 3335
rect 888 3331 892 3335
rect 896 3331 900 3335
rect 1040 3331 1044 3335
rect 1048 3331 1052 3335
rect 1208 3331 1212 3335
rect 1360 3331 1364 3335
rect 1368 3331 1372 3335
rect 1512 3331 1516 3335
rect 1520 3359 1524 3363
rect 200 3315 204 3319
rect 272 3315 276 3319
rect 328 3315 332 3319
rect 408 3315 412 3319
rect 472 3315 476 3319
rect 552 3315 556 3319
rect 632 3315 636 3319
rect 720 3315 724 3319
rect 800 3315 804 3319
rect 272 3291 276 3295
rect 408 3291 412 3295
rect 552 3291 556 3295
rect 720 3291 724 3295
rect 1528 3331 1532 3335
rect 976 3315 980 3319
rect 1160 3315 1164 3319
rect 1344 3315 1348 3319
rect 1520 3315 1524 3319
rect 1536 3315 1540 3319
rect 896 3287 900 3291
rect 2112 3339 2116 3343
rect 2264 3339 2268 3343
rect 2464 3339 2468 3343
rect 3104 3339 3108 3343
rect 3264 3339 3268 3343
rect 3416 3339 3420 3343
rect 2800 3335 2804 3339
rect 1880 3283 1884 3287
rect 2456 3267 2460 3271
rect 488 3259 492 3263
rect 1392 3259 1396 3263
rect 1408 3259 1412 3263
rect 368 3187 372 3191
rect 488 3187 492 3191
rect 496 3215 500 3219
rect 632 3215 636 3219
rect 776 3215 780 3219
rect 1088 3215 1092 3219
rect 2624 3267 2628 3271
rect 3472 3267 3476 3271
rect 1888 3239 1892 3243
rect 2008 3239 2012 3243
rect 2152 3239 2156 3243
rect 2304 3239 2308 3243
rect 2456 3239 2460 3243
rect 2464 3239 2468 3243
rect 2624 3239 2628 3243
rect 2632 3239 2636 3243
rect 2800 3239 2804 3243
rect 2968 3239 2972 3243
rect 3136 3239 3140 3243
rect 3312 3239 3316 3243
rect 3472 3239 3476 3243
rect 3480 3239 3484 3243
rect 1888 3219 1892 3223
rect 2016 3219 2020 3223
rect 2168 3219 2172 3223
rect 2320 3219 2324 3223
rect 2456 3219 2460 3223
rect 2592 3219 2596 3223
rect 2728 3219 2732 3223
rect 2808 3219 2812 3223
rect 2864 3219 2868 3223
rect 3008 3219 3012 3223
rect 3160 3219 3164 3223
rect 3320 3219 3324 3223
rect 3480 3219 3484 3223
rect 1568 3215 1572 3219
rect 2808 3195 2812 3199
rect 496 3187 500 3191
rect 504 3187 508 3191
rect 632 3187 636 3191
rect 640 3187 644 3191
rect 776 3187 780 3191
rect 784 3187 788 3191
rect 936 3187 940 3191
rect 1088 3187 1092 3191
rect 1096 3187 1100 3191
rect 1200 3187 1204 3191
rect 1256 3187 1260 3191
rect 1408 3187 1412 3191
rect 1416 3187 1420 3191
rect 1568 3187 1572 3191
rect 1576 3187 1580 3191
rect 440 3167 444 3171
rect 512 3167 516 3171
rect 552 3167 556 3171
rect 648 3167 652 3171
rect 680 3167 684 3171
rect 752 3167 756 3171
rect 816 3167 820 3171
rect 896 3167 900 3171
rect 968 3167 972 3171
rect 1128 3167 1132 3171
rect 512 3143 516 3147
rect 648 3143 652 3147
rect 752 3143 756 3147
rect 896 3143 900 3147
rect 3472 3179 3476 3183
rect 1200 3143 1204 3147
rect 1208 3167 1212 3171
rect 1288 3167 1292 3171
rect 1456 3167 1460 3171
rect 1632 3167 1636 3171
rect 1208 3139 1212 3143
rect 1552 3127 1556 3131
rect 656 3063 660 3067
rect 776 3063 780 3067
rect 896 3063 900 3067
rect 1024 3063 1028 3067
rect 1104 3063 1108 3067
rect 552 3035 556 3039
rect 656 3035 660 3039
rect 664 3035 668 3039
rect 776 3035 780 3039
rect 784 3035 788 3039
rect 896 3035 900 3039
rect 904 3035 908 3039
rect 1024 3035 1028 3039
rect 1032 3035 1036 3039
rect 1280 3063 1284 3067
rect 1416 3063 1420 3067
rect 2040 3119 2044 3123
rect 2344 3119 2348 3123
rect 2504 3119 2508 3123
rect 2672 3119 2676 3123
rect 3176 3119 3180 3123
rect 1888 3091 1892 3095
rect 1896 3091 1900 3095
rect 2040 3091 2044 3095
rect 2048 3091 2052 3095
rect 2200 3091 2204 3095
rect 2344 3091 2348 3095
rect 2352 3091 2356 3095
rect 2504 3091 2508 3095
rect 2512 3091 2516 3095
rect 2672 3091 2676 3095
rect 2680 3091 2684 3095
rect 2872 3091 2876 3095
rect 3072 3091 3076 3095
rect 3176 3091 3180 3095
rect 3288 3091 3292 3095
rect 3472 3091 3476 3095
rect 3480 3091 3484 3095
rect 1688 3063 1692 3067
rect 1912 3071 1916 3075
rect 2080 3071 2084 3075
rect 2264 3071 2268 3075
rect 2272 3071 2276 3075
rect 2480 3071 2484 3075
rect 2712 3071 2716 3075
rect 2848 3071 2852 3075
rect 2968 3071 2972 3075
rect 3232 3071 3236 3075
rect 3480 3071 3484 3075
rect 1896 3043 1900 3047
rect 1160 3035 1164 3039
rect 1280 3035 1284 3039
rect 1288 3035 1292 3039
rect 1416 3035 1420 3039
rect 1424 3035 1428 3039
rect 1552 3035 1556 3039
rect 1560 3035 1564 3039
rect 1688 3035 1692 3039
rect 1696 3035 1700 3039
rect 568 3019 572 3023
rect 664 3019 668 3023
rect 696 3019 700 3023
rect 824 3019 828 3023
rect 960 3019 964 3023
rect 1040 3019 1044 3023
rect 1096 3019 1100 3023
rect 1104 3019 1108 3023
rect 1232 3019 1236 3023
rect 1360 3019 1364 3023
rect 1488 3019 1492 3023
rect 1568 3019 1572 3023
rect 1616 3019 1620 3023
rect 1728 3019 1732 3023
rect 664 2991 668 2995
rect 1040 2991 1044 2995
rect 1568 2991 1572 2995
rect 2848 3047 2852 3051
rect 2264 2987 2268 2991
rect 3472 3031 3476 3035
rect 2152 2971 2156 2975
rect 2280 2971 2284 2975
rect 2528 2971 2532 2975
rect 2656 2971 2660 2975
rect 2800 2971 2804 2975
rect 2960 2971 2964 2975
rect 3064 2971 3068 2975
rect 3312 2971 3316 2975
rect 2024 2943 2028 2947
rect 2032 2943 2036 2947
rect 2152 2943 2156 2947
rect 2160 2943 2164 2947
rect 2280 2943 2284 2947
rect 2288 2943 2292 2947
rect 2416 2943 2420 2947
rect 2528 2943 2532 2947
rect 2536 2943 2540 2947
rect 2656 2943 2660 2947
rect 2664 2943 2668 2947
rect 2800 2943 2804 2947
rect 2808 2943 2812 2947
rect 2960 2943 2964 2947
rect 2968 2943 2972 2947
rect 3064 2943 3068 2947
rect 3144 2943 3148 2947
rect 3312 2943 3316 2947
rect 3320 2943 3324 2947
rect 3472 2943 3476 2947
rect 3480 2943 3484 2947
rect 872 2939 876 2943
rect 776 2923 780 2927
rect 496 2895 500 2899
rect 640 2895 644 2899
rect 776 2895 780 2899
rect 784 2895 788 2899
rect 912 2923 916 2927
rect 1176 2923 1180 2927
rect 1296 2923 1300 2927
rect 1408 2923 1412 2927
rect 1520 2923 1524 2927
rect 1720 2923 1724 2927
rect 1888 2923 1892 2927
rect 2168 2923 2172 2927
rect 2488 2923 2492 2927
rect 2664 2923 2668 2927
rect 2816 2923 2820 2927
rect 3152 2923 3156 2927
rect 3160 2923 3164 2927
rect 3480 2923 3484 2927
rect 912 2895 916 2899
rect 920 2895 924 2899
rect 1056 2895 1060 2899
rect 1176 2895 1180 2899
rect 1184 2895 1188 2899
rect 1296 2895 1300 2899
rect 1304 2895 1308 2899
rect 1408 2895 1412 2899
rect 1416 2895 1420 2899
rect 1520 2895 1524 2899
rect 1528 2895 1532 2899
rect 1640 2895 1644 2899
rect 1720 2895 1724 2899
rect 1728 2895 1732 2899
rect 2032 2895 2036 2899
rect 1880 2883 1884 2887
rect 320 2879 324 2883
rect 448 2879 452 2883
rect 584 2879 588 2883
rect 720 2879 724 2883
rect 864 2879 868 2883
rect 872 2879 876 2883
rect 1000 2879 1004 2883
rect 1072 2879 1076 2883
rect 1136 2879 1140 2883
rect 1208 2879 1212 2883
rect 1272 2879 1276 2883
rect 1344 2879 1348 2883
rect 1408 2879 1412 2883
rect 1544 2879 1548 2883
rect 1072 2855 1076 2859
rect 1208 2855 1212 2859
rect 1344 2855 1348 2859
rect 416 2839 420 2843
rect 288 2775 292 2779
rect 2664 2843 2668 2847
rect 3152 2843 3156 2847
rect 3472 2883 3476 2887
rect 2016 2827 2020 2831
rect 2352 2827 2356 2831
rect 2512 2827 2516 2831
rect 2800 2827 2804 2831
rect 2928 2827 2932 2831
rect 3048 2827 3052 2831
rect 1880 2799 1884 2803
rect 1888 2799 1892 2803
rect 2016 2799 2020 2803
rect 2024 2799 2028 2803
rect 2192 2799 2196 2803
rect 2200 2799 2204 2803
rect 2352 2799 2356 2803
rect 2360 2799 2364 2803
rect 2512 2799 2516 2803
rect 2520 2799 2524 2803
rect 2672 2799 2676 2803
rect 2800 2799 2804 2803
rect 2808 2799 2812 2803
rect 2928 2799 2932 2803
rect 2936 2799 2940 2803
rect 1888 2787 1892 2791
rect 1968 2787 1972 2791
rect 2056 2787 2060 2791
rect 552 2775 556 2779
rect 944 2775 948 2779
rect 1072 2775 1076 2779
rect 1200 2775 1204 2779
rect 1336 2775 1340 2779
rect 1968 2759 1972 2763
rect 3056 2799 3060 2803
rect 3168 2799 3172 2803
rect 3280 2799 3284 2803
rect 3392 2799 3396 2803
rect 3472 2799 3476 2803
rect 3480 2799 3484 2803
rect 2248 2787 2252 2791
rect 2432 2787 2436 2791
rect 2608 2787 2612 2791
rect 2776 2787 2780 2791
rect 2856 2787 2860 2791
rect 2928 2787 2932 2791
rect 3048 2787 3052 2791
rect 3072 2787 3076 2791
rect 3176 2787 3180 2791
rect 3216 2787 3220 2791
rect 3360 2787 3364 2791
rect 3480 2787 3484 2791
rect 2856 2763 2860 2767
rect 3176 2763 3180 2767
rect 2200 2759 2204 2763
rect 168 2747 172 2751
rect 288 2747 292 2751
rect 296 2747 300 2751
rect 416 2747 420 2751
rect 424 2747 428 2751
rect 552 2747 556 2751
rect 560 2747 564 2751
rect 696 2747 700 2751
rect 824 2747 828 2751
rect 944 2747 948 2751
rect 952 2747 956 2751
rect 1072 2747 1076 2751
rect 1080 2747 1084 2751
rect 1200 2747 1204 2751
rect 1208 2747 1212 2751
rect 1336 2747 1340 2751
rect 1344 2747 1348 2751
rect 2040 2747 2044 2751
rect 984 2739 988 2743
rect 552 2735 556 2739
rect 136 2727 140 2731
rect 224 2727 228 2731
rect 344 2727 348 2731
rect 416 2727 420 2731
rect 472 2727 476 2731
rect 544 2727 548 2731
rect 416 2703 420 2707
rect 544 2703 548 2707
rect 608 2727 612 2731
rect 688 2727 692 2731
rect 752 2727 756 2731
rect 832 2727 836 2731
rect 896 2727 900 2731
rect 976 2727 980 2731
rect 552 2699 556 2703
rect 128 2687 132 2691
rect 832 2703 836 2707
rect 976 2703 980 2707
rect 1040 2727 1044 2731
rect 984 2699 988 2703
rect 688 2643 692 2647
rect 1880 2687 1884 2691
rect 3184 2747 3188 2751
rect 2976 2731 2980 2735
rect 3184 2723 3188 2727
rect 2352 2687 2356 2691
rect 2488 2687 2492 2691
rect 3096 2687 3100 2691
rect 1888 2659 1892 2663
rect 2040 2659 2044 2663
rect 2048 2659 2052 2663
rect 2208 2659 2212 2663
rect 2352 2659 2356 2663
rect 2360 2659 2364 2663
rect 2488 2659 2492 2663
rect 2496 2659 2500 2663
rect 2624 2659 2628 2663
rect 2744 2659 2748 2663
rect 2864 2659 2868 2663
rect 2984 2659 2988 2663
rect 3096 2659 3100 2663
rect 3104 2659 3108 2663
rect 2832 2647 2836 2651
rect 1880 2639 1884 2643
rect 1888 2639 1892 2643
rect 1960 2639 1964 2643
rect 1992 2639 1996 2643
rect 2104 2639 2108 2643
rect 2112 2639 2116 2643
rect 2184 2639 2188 2643
rect 2232 2639 2236 2643
rect 2344 2639 2348 2643
rect 2448 2639 2452 2643
rect 2544 2639 2548 2643
rect 2648 2639 2652 2643
rect 2720 2639 2724 2643
rect 2752 2639 2756 2643
rect 2824 2639 2828 2643
rect 224 2627 228 2631
rect 344 2627 348 2631
rect 464 2627 468 2631
rect 792 2627 796 2631
rect 896 2627 900 2631
rect 992 2627 996 2631
rect 1096 2627 1100 2631
rect 1200 2627 1204 2631
rect 1304 2627 1308 2631
rect 1960 2615 1964 2619
rect 128 2599 132 2603
rect 136 2599 140 2603
rect 224 2599 228 2603
rect 232 2599 236 2603
rect 344 2599 348 2603
rect 352 2599 356 2603
rect 464 2599 468 2603
rect 472 2599 476 2603
rect 584 2599 588 2603
rect 696 2599 700 2603
rect 792 2599 796 2603
rect 800 2599 804 2603
rect 896 2599 900 2603
rect 904 2599 908 2603
rect 992 2599 996 2603
rect 1000 2599 1004 2603
rect 1096 2599 1100 2603
rect 1104 2599 1108 2603
rect 1200 2599 1204 2603
rect 1208 2599 1212 2603
rect 1304 2599 1308 2603
rect 1312 2599 1316 2603
rect 1984 2599 1988 2603
rect 136 2583 140 2587
rect 264 2583 268 2587
rect 408 2583 412 2587
rect 544 2583 548 2587
rect 672 2583 676 2587
rect 800 2583 804 2587
rect 920 2583 924 2587
rect 1040 2583 1044 2587
rect 1168 2583 1172 2587
rect 128 2543 132 2547
rect 1880 2539 1884 2543
rect 2184 2615 2188 2619
rect 2720 2615 2724 2619
rect 2824 2615 2828 2619
rect 2856 2639 2860 2643
rect 2832 2611 2836 2615
rect 2496 2583 2500 2587
rect 2104 2555 2108 2559
rect 2584 2539 2588 2543
rect 2704 2539 2708 2543
rect 2824 2539 2828 2543
rect 1888 2511 1892 2515
rect 1984 2511 1988 2515
rect 1992 2511 1996 2515
rect 2112 2511 2116 2515
rect 2232 2511 2236 2515
rect 2352 2511 2356 2515
rect 2472 2511 2476 2515
rect 2584 2511 2588 2515
rect 2592 2511 2596 2515
rect 2704 2511 2708 2515
rect 2712 2511 2716 2515
rect 2824 2511 2828 2515
rect 2832 2511 2836 2515
rect 1880 2495 1884 2499
rect 1888 2495 1892 2499
rect 1960 2495 1964 2499
rect 2024 2495 2028 2499
rect 2168 2495 2172 2499
rect 2184 2495 2188 2499
rect 2256 2495 2260 2499
rect 2336 2495 2340 2499
rect 2480 2495 2484 2499
rect 2552 2495 2556 2499
rect 2616 2495 2620 2499
rect 2688 2495 2692 2499
rect 2744 2495 2748 2499
rect 2816 2495 2820 2499
rect 2872 2495 2876 2499
rect 2944 2495 2948 2499
rect 3008 2495 3012 2499
rect 272 2487 276 2491
rect 424 2487 428 2491
rect 128 2459 132 2463
rect 136 2459 140 2463
rect 272 2459 276 2463
rect 280 2459 284 2463
rect 424 2459 428 2463
rect 432 2487 436 2491
rect 1000 2487 1004 2491
rect 1136 2487 1140 2491
rect 1272 2487 1276 2491
rect 1960 2471 1964 2475
rect 440 2459 444 2463
rect 592 2459 596 2463
rect 736 2459 740 2463
rect 872 2459 876 2463
rect 1000 2459 1004 2463
rect 1008 2459 1012 2463
rect 1136 2459 1140 2463
rect 1144 2459 1148 2463
rect 1272 2459 1276 2463
rect 1280 2459 1284 2463
rect 184 2447 188 2451
rect 312 2447 316 2451
rect 432 2447 436 2451
rect 448 2447 452 2451
rect 584 2447 588 2451
rect 720 2447 724 2451
rect 856 2447 860 2451
rect 992 2447 996 2451
rect 1064 2447 1068 2451
rect 1128 2447 1132 2451
rect 1200 2447 1204 2451
rect 1264 2447 1268 2451
rect 1336 2447 1340 2451
rect 1400 2447 1404 2451
rect 1064 2423 1068 2427
rect 1200 2423 1204 2427
rect 1336 2423 1340 2427
rect 2256 2471 2260 2475
rect 2552 2471 2556 2475
rect 2688 2471 2692 2475
rect 2816 2471 2820 2475
rect 2944 2471 2948 2475
rect 2168 2415 2172 2419
rect 2792 2399 2796 2403
rect 2944 2399 2948 2403
rect 3104 2399 3108 2403
rect 1888 2371 1892 2375
rect 2016 2371 2020 2375
rect 2176 2371 2180 2375
rect 2336 2371 2340 2375
rect 2472 2371 2476 2375
rect 2496 2371 2500 2375
rect 2648 2371 2652 2375
rect 2792 2371 2796 2375
rect 2800 2371 2804 2375
rect 2944 2371 2948 2375
rect 2952 2371 2956 2375
rect 3104 2371 3108 2375
rect 3112 2371 3116 2375
rect 1920 2355 1924 2359
rect 2008 2355 2012 2359
rect 2080 2355 2084 2359
rect 2240 2355 2244 2359
rect 2328 2355 2332 2359
rect 2400 2355 2404 2359
rect 512 2339 516 2343
rect 1280 2339 1284 2343
rect 2008 2331 2012 2335
rect 2328 2331 2332 2335
rect 2552 2355 2556 2359
rect 2696 2355 2700 2359
rect 2768 2355 2772 2359
rect 2824 2355 2828 2359
rect 2896 2355 2900 2359
rect 2944 2355 2948 2359
rect 3016 2355 3020 2359
rect 3064 2355 3068 2359
rect 3136 2355 3140 2359
rect 3176 2355 3180 2359
rect 3264 2355 3268 2359
rect 3280 2355 3284 2359
rect 3384 2355 3388 2359
rect 3392 2355 3396 2359
rect 3464 2355 3468 2359
rect 3480 2355 3484 2359
rect 2472 2331 2476 2335
rect 2768 2331 2772 2335
rect 2896 2331 2900 2335
rect 3016 2331 3020 2335
rect 3136 2331 3140 2335
rect 160 2311 164 2315
rect 248 2311 252 2315
rect 336 2311 340 2315
rect 440 2311 444 2315
rect 512 2311 516 2315
rect 560 2311 564 2315
rect 688 2311 692 2315
rect 816 2311 820 2315
rect 928 2311 932 2315
rect 952 2311 956 2315
rect 1080 2311 1084 2315
rect 1208 2311 1212 2315
rect 1280 2311 1284 2315
rect 1328 2311 1332 2315
rect 1456 2311 1460 2315
rect 1584 2311 1588 2315
rect 688 2291 692 2295
rect 776 2291 780 2295
rect 856 2291 860 2295
rect 776 2267 780 2271
rect 2128 2299 2132 2303
rect 2136 2299 2140 2303
rect 1016 2291 1020 2295
rect 1168 2291 1172 2295
rect 1248 2291 1252 2295
rect 1312 2291 1316 2295
rect 1392 2291 1396 2295
rect 1456 2291 1460 2295
rect 1528 2291 1532 2295
rect 1592 2291 1596 2295
rect 1664 2291 1668 2295
rect 1728 2291 1732 2295
rect 928 2267 932 2271
rect 1248 2267 1252 2271
rect 1392 2267 1396 2271
rect 1528 2267 1532 2271
rect 1664 2267 1668 2271
rect 3384 2331 3388 2335
rect 3464 2331 3468 2335
rect 3264 2271 3268 2275
rect 3472 2315 3476 2319
rect 2472 2255 2476 2259
rect 2632 2255 2636 2259
rect 2912 2255 2916 2259
rect 3032 2255 3036 2259
rect 1976 2227 1980 2231
rect 2136 2227 2140 2231
rect 2144 2227 2148 2231
rect 2312 2227 2316 2231
rect 2472 2227 2476 2231
rect 2480 2227 2484 2231
rect 2632 2227 2636 2231
rect 2640 2227 2644 2231
rect 2784 2227 2788 2231
rect 2912 2227 2916 2231
rect 2920 2227 2924 2231
rect 3032 2227 3036 2231
rect 3040 2227 3044 2231
rect 3160 2227 3164 2231
rect 3272 2227 3276 2231
rect 3368 2227 3372 2231
rect 3384 2227 3388 2231
rect 3472 2227 3476 2231
rect 3480 2227 3484 2231
rect 2000 2215 2004 2219
rect 2088 2215 2092 2219
rect 2160 2215 2164 2219
rect 2240 2215 2244 2219
rect 2328 2215 2332 2219
rect 2512 2215 2516 2219
rect 2704 2215 2708 2219
rect 2808 2215 2812 2219
rect 2896 2215 2900 2219
rect 3096 2215 3100 2219
rect 3288 2215 3292 2219
rect 3296 2215 3300 2219
rect 2088 2191 2092 2195
rect 2240 2191 2244 2195
rect 3288 2191 3292 2195
rect 3480 2215 3484 2219
rect 3368 2191 3372 2195
rect 712 2187 716 2191
rect 888 2187 892 2191
rect 1064 2187 1068 2191
rect 1400 2187 1404 2191
rect 1568 2187 1572 2191
rect 1720 2187 1724 2191
rect 2808 2187 2812 2191
rect 3472 2175 3476 2179
rect 536 2159 540 2163
rect 712 2159 716 2163
rect 720 2159 724 2163
rect 888 2159 892 2163
rect 896 2159 900 2163
rect 1064 2159 1068 2163
rect 1072 2159 1076 2163
rect 1240 2159 1244 2163
rect 1400 2159 1404 2163
rect 1408 2159 1412 2163
rect 1568 2159 1572 2163
rect 1576 2159 1580 2163
rect 1720 2159 1724 2163
rect 1728 2159 1732 2163
rect 488 2147 492 2151
rect 560 2147 564 2151
rect 616 2147 620 2151
rect 688 2147 692 2151
rect 752 2147 756 2151
rect 824 2147 828 2151
rect 888 2147 892 2151
rect 968 2147 972 2151
rect 1032 2147 1036 2151
rect 1176 2147 1180 2151
rect 1256 2147 1260 2151
rect 1320 2147 1324 2151
rect 1464 2147 1468 2151
rect 1616 2147 1620 2151
rect 560 2123 564 2127
rect 688 2123 692 2127
rect 824 2123 828 2127
rect 968 2123 972 2127
rect 1256 2123 1260 2127
rect 1400 2119 1404 2123
rect 1400 2091 1404 2095
rect 1984 2111 1988 2115
rect 2464 2111 2468 2115
rect 2608 2111 2612 2115
rect 2752 2111 2756 2115
rect 2024 2083 2028 2087
rect 2168 2083 2172 2087
rect 2320 2083 2324 2087
rect 2464 2083 2468 2087
rect 2472 2083 2476 2087
rect 2608 2083 2612 2087
rect 2616 2083 2620 2087
rect 2752 2083 2756 2087
rect 2760 2083 2764 2087
rect 2896 2083 2900 2087
rect 3024 2083 3028 2087
rect 3144 2083 3148 2087
rect 3224 2083 3228 2087
rect 3264 2083 3268 2087
rect 3384 2083 3388 2087
rect 3472 2083 3476 2087
rect 3480 2083 3484 2087
rect 1976 2067 1980 2071
rect 1984 2067 1988 2071
rect 2064 2067 2068 2071
rect 2136 2067 2140 2071
rect 2304 2067 2308 2071
rect 2392 2067 2396 2071
rect 2464 2067 2468 2071
rect 2552 2067 2556 2071
rect 2624 2067 2628 2071
rect 2768 2067 2772 2071
rect 2840 2067 2844 2071
rect 2904 2067 2908 2071
rect 3032 2067 3036 2071
rect 3104 2067 3108 2071
rect 3152 2067 3156 2071
rect 424 2047 428 2051
rect 544 2047 548 2051
rect 672 2047 676 2051
rect 792 2047 796 2051
rect 1032 2047 1036 2051
rect 1136 2047 1140 2051
rect 320 2019 324 2023
rect 424 2019 428 2023
rect 432 2019 436 2023
rect 544 2019 548 2023
rect 552 2019 556 2023
rect 672 2019 676 2023
rect 680 2019 684 2023
rect 792 2019 796 2023
rect 800 2019 804 2023
rect 920 2019 924 2023
rect 1032 2019 1036 2023
rect 1040 2019 1044 2023
rect 2064 2043 2068 2047
rect 2392 2039 2396 2043
rect 2840 2043 2844 2047
rect 3104 2043 3108 2047
rect 3224 2043 3228 2047
rect 3232 2075 3236 2079
rect 3272 2067 3276 2071
rect 3384 2067 3388 2071
rect 3480 2067 3484 2071
rect 2552 2039 2556 2043
rect 3232 2039 3236 2043
rect 3024 2027 3028 2031
rect 1160 2019 1164 2023
rect 1280 2019 1284 2023
rect 1408 2019 1412 2023
rect 608 2011 612 2015
rect 1136 2011 1140 2015
rect 2184 2011 2188 2015
rect 2192 2011 2196 2015
rect 176 2003 180 2007
rect 248 2003 252 2007
rect 288 2003 292 2007
rect 360 2003 364 2007
rect 408 2003 412 2007
rect 480 2003 484 2007
rect 528 2003 532 2007
rect 600 2003 604 2007
rect 248 1979 252 1983
rect 360 1979 364 1983
rect 480 1979 484 1983
rect 600 1979 604 1983
rect 648 2003 652 2007
rect 768 2003 772 2007
rect 888 2003 892 2007
rect 1008 2003 1012 2007
rect 1128 2003 1132 2007
rect 1200 2003 1204 2007
rect 1248 2003 1252 2007
rect 1200 1979 1204 1983
rect 608 1975 612 1979
rect 816 1947 820 1951
rect 832 1947 836 1951
rect 2536 1971 2540 1975
rect 2864 1971 2868 1975
rect 216 1903 220 1907
rect 344 1903 348 1907
rect 488 1903 492 1907
rect 648 1903 652 1907
rect 1888 1943 1892 1947
rect 2032 1943 2036 1947
rect 2192 1943 2196 1947
rect 2200 1943 2204 1947
rect 2376 1943 2380 1947
rect 2536 1943 2540 1947
rect 2544 1943 2548 1947
rect 2712 1943 2716 1947
rect 2864 1943 2868 1947
rect 2872 1943 2876 1947
rect 3024 1943 3028 1947
rect 3040 1943 3044 1947
rect 3208 1943 3212 1947
rect 2064 1931 2068 1935
rect 1888 1923 1892 1927
rect 1984 1923 1988 1927
rect 2056 1923 2060 1927
rect 1008 1903 1012 1907
rect 1240 1903 1244 1907
rect 1456 1903 1460 1907
rect 136 1875 140 1879
rect 216 1875 220 1879
rect 224 1875 228 1879
rect 344 1875 348 1879
rect 352 1875 356 1879
rect 488 1875 492 1879
rect 496 1875 500 1879
rect 648 1875 652 1879
rect 656 1875 660 1879
rect 832 1875 836 1879
rect 840 1875 844 1879
rect 1008 1875 1012 1879
rect 1040 1875 1044 1879
rect 1240 1875 1244 1879
rect 1248 1875 1252 1879
rect 1256 1875 1260 1879
rect 136 1855 140 1859
rect 264 1855 268 1859
rect 408 1855 412 1859
rect 552 1855 556 1859
rect 648 1855 652 1859
rect 688 1855 692 1859
rect 816 1855 820 1859
rect 936 1855 940 1859
rect 1048 1855 1052 1859
rect 1120 1855 1124 1859
rect 1152 1855 1156 1859
rect 1120 1831 1124 1835
rect 2056 1899 2060 1903
rect 2112 1923 2116 1927
rect 2248 1923 2252 1927
rect 2376 1923 2380 1927
rect 2504 1923 2508 1927
rect 2624 1923 2628 1927
rect 2744 1923 2748 1927
rect 2872 1923 2876 1927
rect 3000 1923 3004 1927
rect 2064 1895 2068 1899
rect 1464 1875 1468 1879
rect 1256 1855 1260 1859
rect 1328 1855 1332 1859
rect 1352 1855 1356 1859
rect 1448 1855 1452 1859
rect 1456 1855 1460 1859
rect 1544 1855 1548 1859
rect 1640 1855 1644 1859
rect 1728 1855 1732 1859
rect 1248 1831 1252 1835
rect 1328 1831 1332 1835
rect 648 1827 652 1831
rect 2352 1819 2356 1823
rect 1400 1799 1404 1803
rect 2616 1819 2620 1823
rect 2736 1819 2740 1823
rect 2856 1819 2860 1823
rect 2984 1819 2988 1823
rect 2224 1791 2228 1795
rect 2352 1791 2356 1795
rect 2360 1791 2364 1795
rect 2496 1791 2500 1795
rect 2616 1791 2620 1795
rect 2624 1791 2628 1795
rect 2736 1791 2740 1795
rect 2744 1791 2748 1795
rect 2856 1791 2860 1795
rect 2864 1791 2868 1795
rect 2984 1791 2988 1795
rect 2992 1791 2996 1795
rect 2264 1775 2268 1779
rect 2352 1775 2356 1779
rect 2448 1775 2452 1779
rect 2552 1775 2556 1779
rect 2632 1775 2636 1779
rect 2656 1775 2660 1779
rect 2752 1775 2756 1779
rect 2824 1775 2828 1779
rect 2856 1775 2860 1779
rect 2928 1775 2932 1779
rect 2960 1775 2964 1779
rect 3032 1775 3036 1779
rect 3064 1775 3068 1779
rect 3152 1775 3156 1779
rect 3168 1775 3172 1779
rect 840 1763 844 1767
rect 296 1747 300 1751
rect 568 1747 572 1751
rect 136 1719 140 1723
rect 296 1719 300 1723
rect 304 1719 308 1723
rect 496 1719 500 1723
rect 568 1719 572 1723
rect 688 1719 692 1723
rect 2824 1751 2828 1755
rect 2928 1751 2932 1755
rect 3032 1751 3036 1755
rect 3152 1751 3156 1755
rect 864 1747 868 1751
rect 1208 1747 1212 1751
rect 1520 1747 1524 1751
rect 864 1719 868 1723
rect 872 1719 876 1723
rect 1048 1719 1052 1723
rect 1208 1719 1212 1723
rect 1216 1719 1220 1723
rect 1376 1719 1380 1723
rect 1520 1711 1524 1715
rect 1528 1747 1532 1751
rect 1696 1747 1700 1751
rect 2632 1747 2636 1751
rect 1536 1719 1540 1723
rect 1704 1719 1708 1723
rect 128 1703 132 1707
rect 136 1703 140 1707
rect 280 1703 284 1707
rect 464 1703 468 1707
rect 600 1703 604 1707
rect 648 1703 652 1707
rect 832 1703 836 1707
rect 840 1703 844 1707
rect 1016 1703 1020 1707
rect 1184 1703 1188 1707
rect 1264 1703 1268 1707
rect 1352 1703 1356 1707
rect 1520 1703 1524 1707
rect 1528 1703 1532 1707
rect 1688 1703 1692 1707
rect 1696 1703 1700 1707
rect 600 1675 604 1679
rect 3352 1691 3356 1695
rect 1264 1675 1268 1679
rect 2360 1675 2364 1679
rect 2488 1675 2492 1679
rect 2616 1675 2620 1679
rect 2752 1675 2756 1679
rect 3008 1675 3012 1679
rect 3240 1675 3244 1679
rect 1720 1647 1724 1651
rect 1736 1647 1740 1651
rect 2248 1647 2252 1651
rect 2360 1647 2364 1651
rect 2368 1647 2372 1651
rect 2488 1647 2492 1651
rect 2496 1647 2500 1651
rect 2616 1647 2620 1651
rect 2624 1647 2628 1651
rect 2752 1647 2756 1651
rect 2760 1647 2764 1651
rect 2888 1647 2892 1651
rect 3008 1647 3012 1651
rect 3016 1647 3020 1651
rect 3136 1647 3140 1651
rect 3240 1647 3244 1651
rect 3248 1647 3252 1651
rect 128 1615 132 1619
rect 768 1615 772 1619
rect 440 1599 444 1603
rect 624 1599 628 1603
rect 136 1571 140 1575
rect 272 1571 276 1575
rect 440 1571 444 1575
rect 448 1571 452 1575
rect 624 1571 628 1575
rect 632 1571 636 1575
rect 1264 1615 1268 1619
rect 808 1599 812 1603
rect 808 1571 812 1575
rect 816 1571 820 1575
rect 992 1571 996 1575
rect 1152 1571 1156 1575
rect 1296 1599 1300 1603
rect 1592 1599 1596 1603
rect 2624 1639 2628 1643
rect 2144 1631 2148 1635
rect 2216 1631 2220 1635
rect 2336 1631 2340 1635
rect 2432 1631 2436 1635
rect 2520 1631 2524 1635
rect 2616 1631 2620 1635
rect 2216 1607 2220 1611
rect 2432 1607 2436 1611
rect 2616 1607 2620 1611
rect 3360 1675 3364 1679
rect 3472 1675 3476 1679
rect 3360 1647 3364 1651
rect 3368 1647 3372 1651
rect 2696 1631 2700 1635
rect 2864 1631 2868 1635
rect 2952 1631 2956 1635
rect 3024 1631 3028 1635
rect 3184 1631 3188 1635
rect 3272 1631 3276 1635
rect 3344 1631 3348 1635
rect 3352 1631 3356 1635
rect 3480 1647 3484 1651
rect 3472 1631 3476 1635
rect 3480 1631 3484 1635
rect 2952 1607 2956 1611
rect 2624 1603 2628 1607
rect 3272 1603 3276 1607
rect 3104 1591 3108 1595
rect 1296 1571 1300 1575
rect 1304 1571 1308 1575
rect 1456 1571 1460 1575
rect 1592 1571 1596 1575
rect 1600 1571 1604 1575
rect 1720 1571 1724 1575
rect 1728 1571 1732 1575
rect 136 1559 140 1563
rect 264 1559 268 1563
rect 424 1559 428 1563
rect 592 1559 596 1563
rect 760 1559 764 1563
rect 768 1559 772 1563
rect 928 1559 932 1563
rect 1096 1559 1100 1563
rect 1256 1559 1260 1563
rect 1264 1559 1268 1563
rect 1416 1559 1420 1563
rect 1584 1559 1588 1563
rect 1728 1559 1732 1563
rect 2448 1535 2452 1539
rect 2784 1535 2788 1539
rect 2944 1535 2948 1539
rect 3264 1535 3268 1539
rect 2088 1507 2092 1511
rect 2280 1507 2284 1511
rect 2448 1507 2452 1511
rect 2456 1507 2460 1511
rect 2624 1507 2628 1511
rect 2784 1507 2788 1511
rect 2792 1507 2796 1511
rect 2944 1507 2948 1511
rect 2952 1507 2956 1511
rect 3104 1507 3108 1511
rect 3112 1507 3116 1511
rect 3264 1507 3268 1511
rect 3272 1507 3276 1511
rect 3368 1507 3372 1511
rect 3432 1507 3436 1511
rect 1888 1487 1892 1491
rect 1960 1487 1964 1491
rect 1984 1487 1988 1491
rect 2112 1487 2116 1491
rect 2240 1487 2244 1491
rect 2336 1487 2340 1491
rect 2376 1487 2380 1491
rect 2528 1487 2532 1491
rect 2616 1487 2620 1491
rect 2696 1487 2700 1491
rect 2880 1487 2884 1491
rect 3080 1487 3084 1491
rect 3192 1487 3196 1491
rect 3288 1487 3292 1491
rect 704 1475 708 1479
rect 464 1459 468 1463
rect 600 1459 604 1463
rect 184 1431 188 1435
rect 328 1431 332 1435
rect 464 1431 468 1435
rect 472 1431 476 1435
rect 600 1431 604 1435
rect 608 1431 612 1435
rect 1960 1463 1964 1467
rect 2616 1463 2620 1467
rect 3192 1463 3196 1467
rect 736 1459 740 1463
rect 1224 1459 1228 1463
rect 2336 1459 2340 1463
rect 736 1431 740 1435
rect 744 1431 748 1435
rect 872 1431 876 1435
rect 992 1431 996 1435
rect 1120 1431 1124 1435
rect 2064 1447 2068 1451
rect 1248 1431 1252 1435
rect 1376 1431 1380 1435
rect 192 1411 196 1415
rect 328 1411 332 1415
rect 456 1411 460 1415
rect 528 1411 532 1415
rect 576 1411 580 1415
rect 696 1411 700 1415
rect 704 1411 708 1415
rect 808 1411 812 1415
rect 880 1411 884 1415
rect 912 1411 916 1415
rect 984 1411 988 1415
rect 1008 1411 1012 1415
rect 1080 1411 1084 1415
rect 1112 1411 1116 1415
rect 1216 1411 1220 1415
rect 1224 1411 1228 1415
rect 1288 1411 1292 1415
rect 1320 1411 1324 1415
rect 528 1387 532 1391
rect 880 1387 884 1391
rect 984 1387 988 1391
rect 1080 1387 1084 1391
rect 1288 1387 1292 1391
rect 1880 1387 1884 1391
rect 688 1371 692 1375
rect 320 1311 324 1315
rect 1368 1355 1372 1359
rect 2800 1447 2804 1451
rect 3024 1387 3028 1391
rect 1888 1359 1892 1363
rect 1976 1359 1980 1363
rect 2064 1359 2068 1363
rect 2072 1359 2076 1363
rect 2184 1359 2188 1363
rect 2192 1359 2196 1363
rect 2304 1359 2308 1363
rect 2440 1359 2444 1363
rect 2608 1359 2612 1363
rect 2800 1359 2804 1363
rect 2808 1359 2812 1363
rect 3024 1359 3028 1363
rect 3032 1359 3036 1363
rect 3264 1359 3268 1363
rect 1880 1343 1884 1347
rect 1888 1343 1892 1347
rect 1960 1343 1964 1347
rect 1976 1343 1980 1347
rect 2048 1343 2052 1347
rect 2096 1343 2100 1347
rect 2168 1343 2172 1347
rect 1960 1319 1964 1323
rect 2048 1319 2052 1323
rect 2168 1319 2172 1323
rect 2216 1343 2220 1347
rect 2352 1343 2356 1347
rect 2432 1343 2436 1347
rect 2504 1343 2508 1347
rect 2600 1343 2604 1347
rect 2680 1343 2684 1347
rect 2776 1343 2780 1347
rect 2864 1343 2868 1347
rect 2968 1343 2972 1347
rect 3064 1343 3068 1347
rect 3272 1343 3276 1347
rect 2432 1319 2436 1323
rect 2600 1319 2604 1323
rect 2776 1319 2780 1323
rect 2968 1319 2972 1323
rect 3480 1487 3484 1491
rect 3472 1447 3476 1451
rect 3472 1359 3476 1363
rect 3480 1359 3484 1363
rect 3480 1343 3484 1347
rect 3368 1319 3372 1323
rect 2192 1315 2196 1319
rect 1000 1311 1004 1315
rect 232 1283 236 1287
rect 320 1283 324 1287
rect 384 1283 388 1287
rect 544 1283 548 1287
rect 688 1283 692 1287
rect 704 1283 708 1287
rect 872 1283 876 1287
rect 1040 1283 1044 1287
rect 1208 1283 1212 1287
rect 1376 1283 1380 1287
rect 208 1271 212 1275
rect 288 1271 292 1275
rect 352 1271 356 1275
rect 440 1271 444 1275
rect 512 1271 516 1275
rect 584 1271 588 1275
rect 672 1271 676 1275
rect 760 1271 764 1275
rect 832 1271 836 1275
rect 992 1271 996 1275
rect 1000 1271 1004 1275
rect 1072 1271 1076 1275
rect 1144 1271 1148 1275
rect 1224 1271 1228 1275
rect 1288 1271 1292 1275
rect 1368 1271 1372 1275
rect 1432 1271 1436 1275
rect 1576 1271 1580 1275
rect 1584 1271 1588 1275
rect 288 1247 292 1251
rect 440 1247 444 1251
rect 584 1247 588 1251
rect 760 1247 764 1251
rect 1072 1247 1076 1251
rect 1224 1247 1228 1251
rect 1368 1247 1372 1251
rect 1576 1247 1580 1251
rect 2136 1235 2140 1239
rect 2056 1207 2060 1211
rect 2328 1235 2332 1239
rect 2680 1235 2684 1239
rect 2848 1235 2852 1239
rect 3032 1235 3036 1239
rect 3224 1235 3228 1239
rect 2144 1207 2148 1211
rect 2240 1207 2244 1211
rect 2328 1207 2332 1211
rect 2336 1207 2340 1211
rect 2432 1207 2436 1211
rect 2552 1207 2556 1211
rect 2680 1207 2684 1211
rect 2688 1207 2692 1211
rect 2848 1207 2852 1211
rect 2856 1207 2860 1211
rect 3032 1207 3036 1211
rect 3040 1207 3044 1211
rect 3224 1207 3228 1211
rect 3232 1207 3236 1211
rect 3432 1207 3436 1211
rect 2224 1199 2228 1203
rect 2032 1191 2036 1195
rect 2136 1191 2140 1195
rect 2144 1191 2148 1195
rect 2216 1191 2220 1195
rect 680 1167 684 1171
rect 1392 1167 1396 1171
rect 2216 1167 2220 1171
rect 2272 1191 2276 1195
rect 2408 1191 2412 1195
rect 2552 1191 2556 1195
rect 2704 1191 2708 1195
rect 2856 1191 2860 1195
rect 3008 1191 3012 1195
rect 3160 1191 3164 1195
rect 3312 1191 3316 1195
rect 3320 1191 3324 1195
rect 3480 1191 3484 1195
rect 136 1139 140 1143
rect 272 1139 276 1143
rect 360 1139 364 1143
rect 424 1139 428 1143
rect 576 1139 580 1143
rect 680 1139 684 1143
rect 728 1139 732 1143
rect 888 1139 892 1143
rect 1056 1139 1060 1143
rect 1232 1139 1236 1143
rect 128 1127 132 1131
rect 136 1127 140 1131
rect 216 1127 220 1131
rect 288 1127 292 1131
rect 216 1103 220 1107
rect 2224 1163 2228 1167
rect 1416 1139 1420 1143
rect 1600 1139 1604 1143
rect 472 1127 476 1131
rect 656 1127 660 1131
rect 752 1127 756 1131
rect 840 1127 844 1131
rect 1024 1127 1028 1131
rect 1120 1127 1124 1131
rect 1200 1127 1204 1131
rect 1384 1127 1388 1131
rect 1392 1127 1396 1131
rect 1496 1127 1500 1131
rect 1568 1127 1572 1131
rect 1656 1127 1660 1131
rect 1728 1127 1732 1131
rect 360 1103 364 1107
rect 752 1103 756 1107
rect 1120 1103 1124 1107
rect 1496 1103 1500 1107
rect 1656 1103 1660 1107
rect 3312 1099 3316 1103
rect 3472 1151 3476 1155
rect 128 1047 132 1051
rect 1720 1087 1724 1091
rect 424 1031 428 1035
rect 576 1031 580 1035
rect 728 1031 732 1035
rect 1376 1031 1380 1035
rect 1656 1031 1660 1035
rect 136 1003 140 1007
rect 224 1003 228 1007
rect 272 1003 276 1007
rect 424 1003 428 1007
rect 432 1003 436 1007
rect 576 1003 580 1007
rect 584 1003 588 1007
rect 728 1003 732 1007
rect 736 1003 740 1007
rect 888 1003 892 1007
rect 1048 1003 1052 1007
rect 1216 1003 1220 1007
rect 1376 1003 1380 1007
rect 1384 1003 1388 1007
rect 1560 1003 1564 1007
rect 1656 1003 1660 1007
rect 2080 1083 2084 1087
rect 2224 1083 2228 1087
rect 2528 1083 2532 1087
rect 2832 1083 2836 1087
rect 2984 1083 2988 1087
rect 3144 1083 3148 1087
rect 1944 1055 1948 1059
rect 2080 1055 2084 1059
rect 2088 1055 2092 1059
rect 2224 1055 2228 1059
rect 2232 1055 2236 1059
rect 2384 1055 2388 1059
rect 2392 1055 2396 1059
rect 2528 1055 2532 1059
rect 2536 1055 2540 1059
rect 2688 1055 2692 1059
rect 2832 1055 2836 1059
rect 2840 1055 2844 1059
rect 2984 1055 2988 1059
rect 2992 1055 2996 1059
rect 3144 1055 3148 1059
rect 3152 1055 3156 1059
rect 3320 1055 3324 1059
rect 3328 1055 3332 1059
rect 3472 1055 3476 1059
rect 3480 1055 3484 1059
rect 1912 1031 1916 1035
rect 2120 1031 2124 1035
rect 2320 1031 2324 1035
rect 2392 1007 2396 1011
rect 2424 1031 2428 1035
rect 2512 1031 2516 1035
rect 2688 1031 2692 1035
rect 2776 1031 2780 1035
rect 2856 1031 2860 1035
rect 2944 1031 2948 1035
rect 3016 1031 3020 1035
rect 3088 1031 3092 1035
rect 3176 1031 3180 1035
rect 2776 1007 2780 1011
rect 2944 1007 2948 1011
rect 3088 1007 3092 1011
rect 3336 1031 3340 1035
rect 3480 1031 3484 1035
rect 1720 1003 1724 1007
rect 1728 1003 1732 1007
rect 2424 1003 2428 1007
rect 3328 1003 3332 1007
rect 128 987 132 991
rect 136 987 140 991
rect 216 987 220 991
rect 216 963 220 967
rect 3472 991 3476 995
rect 280 987 284 991
rect 456 987 460 991
rect 536 987 540 991
rect 640 987 644 991
rect 728 987 732 991
rect 816 987 820 991
rect 992 987 996 991
rect 1080 987 1084 991
rect 1160 987 1164 991
rect 1320 987 1324 991
rect 1400 987 1404 991
rect 1480 987 1484 991
rect 1648 987 1652 991
rect 224 959 228 963
rect 536 959 540 963
rect 1080 963 1084 967
rect 1400 963 1404 967
rect 728 959 732 963
rect 128 899 132 903
rect 600 947 604 951
rect 1528 931 1532 935
rect 1544 931 1548 935
rect 768 883 772 887
rect 1392 883 1396 887
rect 1480 883 1484 887
rect 136 855 140 859
rect 208 855 212 859
rect 272 855 276 859
rect 440 855 444 859
rect 600 855 604 859
rect 608 855 612 859
rect 768 855 772 859
rect 776 855 780 859
rect 936 855 940 859
rect 1048 855 1052 859
rect 1096 855 1100 859
rect 1248 855 1252 859
rect 1392 855 1396 859
rect 1400 855 1404 859
rect 128 843 132 847
rect 136 843 140 847
rect 280 843 284 847
rect 376 843 380 847
rect 456 843 460 847
rect 544 843 548 847
rect 632 843 636 847
rect 720 843 724 847
rect 800 843 804 847
rect 976 843 980 847
rect 208 819 212 823
rect 376 819 380 823
rect 544 819 548 823
rect 720 819 724 823
rect 2064 931 2068 935
rect 2448 931 2452 935
rect 2624 931 2628 935
rect 2944 931 2948 935
rect 3088 931 3092 935
rect 3224 931 3228 935
rect 3360 931 3364 935
rect 1888 903 1892 907
rect 2064 903 2068 907
rect 2072 903 2076 907
rect 2264 903 2268 907
rect 2288 903 2292 907
rect 2448 903 2452 907
rect 2456 903 2460 907
rect 2624 903 2628 907
rect 2632 903 2636 907
rect 2800 903 2804 907
rect 2944 903 2948 907
rect 2952 903 2956 907
rect 3088 903 3092 907
rect 3096 903 3100 907
rect 3224 903 3228 907
rect 3232 903 3236 907
rect 3360 903 3364 907
rect 3368 903 3372 907
rect 3472 903 3476 907
rect 3480 903 3484 907
rect 1888 883 1892 887
rect 2016 883 2020 887
rect 2104 883 2108 887
rect 2176 883 2180 887
rect 1544 855 1548 859
rect 1552 855 1556 859
rect 2104 855 2108 859
rect 2344 883 2348 887
rect 2512 883 2516 887
rect 2680 883 2684 887
rect 2832 883 2836 887
rect 2976 883 2980 887
rect 3112 883 3116 887
rect 3240 883 3244 887
rect 3352 883 3356 887
rect 3368 883 3372 887
rect 3480 883 3484 887
rect 2288 855 2292 859
rect 1152 843 1156 847
rect 1328 843 1332 847
rect 1408 843 1412 847
rect 1480 843 1484 847
rect 1504 843 1508 847
rect 1880 843 1884 847
rect 1048 819 1052 823
rect 1408 815 1412 819
rect 128 759 132 763
rect 3352 795 3356 799
rect 3472 843 3476 847
rect 2064 779 2068 783
rect 2440 779 2444 783
rect 2616 779 2620 783
rect 2936 779 2940 783
rect 3080 779 3084 783
rect 3352 779 3356 783
rect 1880 751 1884 755
rect 1888 751 1892 755
rect 2064 751 2068 755
rect 2072 751 2076 755
rect 2264 751 2268 755
rect 2440 751 2444 755
rect 2448 751 2452 755
rect 2616 751 2620 755
rect 2624 751 2628 755
rect 2792 751 2796 755
rect 2936 751 2940 755
rect 2944 751 2948 755
rect 3080 751 3084 755
rect 3088 751 3092 755
rect 3224 751 3228 755
rect 3352 751 3356 755
rect 3360 751 3364 755
rect 3464 751 3468 755
rect 432 743 436 747
rect 136 715 140 719
rect 272 715 276 719
rect 1080 743 1084 747
rect 1384 743 1388 747
rect 1544 743 1548 747
rect 1888 739 1892 743
rect 1984 739 1988 743
rect 2064 739 2068 743
rect 2256 739 2260 743
rect 2440 739 2444 743
rect 2616 739 2620 743
rect 2712 739 2716 743
rect 2792 739 2796 743
rect 2968 739 2972 743
rect 3144 739 3148 743
rect 3240 739 3244 743
rect 3320 739 3324 743
rect 440 715 444 719
rect 608 715 612 719
rect 776 715 780 719
rect 936 715 940 719
rect 944 715 948 719
rect 1080 715 1084 719
rect 1088 715 1092 719
rect 1240 715 1244 719
rect 1384 715 1388 719
rect 1392 715 1396 719
rect 1544 715 1548 719
rect 1552 715 1556 719
rect 1984 715 1988 719
rect 2712 715 2716 719
rect 3240 715 3244 719
rect 128 699 132 703
rect 136 699 140 703
rect 280 699 284 703
rect 432 699 436 703
rect 448 699 452 703
rect 616 699 620 703
rect 784 699 788 703
rect 952 699 956 703
rect 1104 699 1108 703
rect 1112 699 1116 703
rect 1272 699 1276 703
rect 1432 699 1436 703
rect 1592 699 1596 703
rect 2928 699 2932 703
rect 944 671 948 675
rect 128 611 132 615
rect 2112 683 2116 687
rect 1104 611 1108 615
rect 1264 659 1268 663
rect 448 595 452 599
rect 136 567 140 571
rect 288 567 292 571
rect 296 567 300 571
rect 136 551 140 555
rect 144 551 148 555
rect 232 551 236 555
rect 232 527 236 531
rect 1112 595 1116 599
rect 1880 639 1884 643
rect 2344 639 2348 643
rect 2472 639 2476 643
rect 2760 639 2764 643
rect 3112 639 3116 643
rect 1888 611 1892 615
rect 1976 611 1980 615
rect 2096 611 2100 615
rect 2224 611 2228 615
rect 2344 611 2348 615
rect 2352 611 2356 615
rect 2472 611 2476 615
rect 2480 611 2484 615
rect 2616 611 2620 615
rect 2760 611 2764 615
rect 2768 611 2772 615
rect 2928 611 2932 615
rect 2936 611 2940 615
rect 3112 611 3116 615
rect 3120 611 3124 615
rect 3312 611 3316 615
rect 3176 603 3180 607
rect 1408 595 1412 599
rect 1552 595 1556 599
rect 1704 595 1708 599
rect 1880 595 1884 599
rect 1888 595 1892 599
rect 2040 595 2044 599
rect 2128 595 2132 599
rect 2208 595 2212 599
rect 2384 595 2388 599
rect 2488 595 2492 599
rect 2576 595 2580 599
rect 2792 595 2796 599
rect 2912 595 2916 599
rect 3016 595 3020 599
rect 3088 595 3092 599
rect 2128 571 2132 575
rect 2912 571 2916 575
rect 3088 571 3092 575
rect 3248 595 3252 599
rect 456 567 460 571
rect 632 567 636 571
rect 800 567 804 571
rect 968 567 972 571
rect 1112 567 1116 571
rect 1120 567 1124 571
rect 1264 567 1268 571
rect 1272 567 1276 571
rect 1408 567 1412 571
rect 1416 567 1420 571
rect 1552 567 1556 571
rect 1560 567 1564 571
rect 1704 567 1708 571
rect 1712 567 1716 571
rect 2488 567 2492 571
rect 3176 567 3180 571
rect 3480 751 3484 755
rect 3472 739 3476 743
rect 3480 739 3484 743
rect 3472 699 3476 703
rect 3472 611 3476 615
rect 3480 611 3484 615
rect 3480 595 3484 599
rect 3464 567 3468 571
rect 2480 555 2484 559
rect 304 551 308 555
rect 448 551 452 555
rect 464 551 468 555
rect 552 551 556 555
rect 624 551 628 555
rect 704 551 708 555
rect 776 551 780 555
rect 920 551 924 555
rect 1056 551 1060 555
rect 1184 551 1188 555
rect 1256 551 1260 555
rect 1304 551 1308 555
rect 1376 551 1380 555
rect 1416 551 1420 555
rect 1528 551 1532 555
rect 1640 551 1644 555
rect 1728 551 1732 555
rect 552 527 556 531
rect 704 527 708 531
rect 1256 527 1260 531
rect 1376 527 1380 531
rect 296 523 300 527
rect 1464 495 1468 499
rect 2272 491 2276 495
rect 2624 491 2628 495
rect 2800 491 2804 495
rect 2984 491 2988 495
rect 3176 491 3180 495
rect 136 463 140 467
rect 2120 463 2124 467
rect 2192 463 2196 467
rect 2272 463 2276 467
rect 2280 463 2284 467
rect 2376 463 2380 467
rect 2480 463 2484 467
rect 2488 463 2492 467
rect 2624 463 2628 467
rect 2632 463 2636 467
rect 2800 463 2804 467
rect 2808 463 2812 467
rect 2984 463 2988 467
rect 3008 463 3012 467
rect 3176 463 3180 467
rect 3216 463 3220 467
rect 3424 463 3428 467
rect 3432 463 3436 467
rect 248 447 252 451
rect 552 447 556 451
rect 1000 447 1004 451
rect 1232 447 1236 451
rect 1336 447 1340 451
rect 1536 447 1540 451
rect 1632 447 1636 451
rect 1712 447 1716 451
rect 1888 443 1892 447
rect 2032 443 2036 447
rect 160 419 164 423
rect 248 419 252 423
rect 312 419 316 423
rect 464 419 468 423
rect 552 419 556 423
rect 616 419 620 423
rect 760 419 764 423
rect 888 419 892 423
rect 1000 419 1004 423
rect 1008 419 1012 423
rect 1128 419 1132 423
rect 1232 419 1236 423
rect 1240 419 1244 423
rect 1336 419 1340 423
rect 1344 419 1348 423
rect 1440 419 1444 423
rect 1536 419 1540 423
rect 1544 419 1548 423
rect 1632 419 1636 423
rect 1640 419 1644 423
rect 1712 419 1716 423
rect 1728 419 1732 423
rect 2120 419 2124 423
rect 2128 443 2132 447
rect 2200 443 2204 447
rect 2376 443 2380 447
rect 2480 443 2484 447
rect 2568 443 2572 447
rect 2680 443 2684 447
rect 2776 443 2780 447
rect 2896 443 2900 447
rect 3000 443 3004 447
rect 3080 443 3084 447
rect 3232 443 3236 447
rect 2480 419 2484 423
rect 2680 419 2684 423
rect 2896 419 2900 423
rect 3080 419 3084 423
rect 2128 415 2132 419
rect 144 407 148 411
rect 216 407 220 411
rect 264 407 268 411
rect 392 407 396 411
rect 400 407 404 411
rect 544 407 548 411
rect 704 407 708 411
rect 800 407 804 411
rect 880 407 884 411
rect 1056 407 1060 411
rect 1152 407 1156 411
rect 1240 407 1244 411
rect 1432 407 1436 411
rect 1536 407 1540 411
rect 1632 407 1636 411
rect 216 383 220 387
rect 800 383 804 387
rect 1152 383 1156 387
rect 1536 383 1540 387
rect 1880 403 1884 407
rect 392 311 396 315
rect 1664 351 1668 355
rect 1680 351 1684 355
rect 216 295 220 299
rect 304 295 308 299
rect 392 295 396 299
rect 568 295 572 299
rect 656 295 660 299
rect 744 295 748 299
rect 136 267 140 271
rect 216 267 220 271
rect 224 267 228 271
rect 304 267 308 271
rect 312 267 316 271
rect 392 267 396 271
rect 400 267 404 271
rect 488 267 492 271
rect 568 267 572 271
rect 576 267 580 271
rect 656 267 660 271
rect 664 267 668 271
rect 1008 295 1012 299
rect 1376 295 1380 299
rect 1472 295 1476 299
rect 1552 295 1556 299
rect 752 267 756 271
rect 840 267 844 271
rect 928 267 932 271
rect 1008 267 1012 271
rect 1016 267 1020 271
rect 1104 267 1108 271
rect 1192 267 1196 271
rect 1288 267 1292 271
rect 1376 267 1380 271
rect 1384 267 1388 271
rect 1472 267 1476 271
rect 1480 267 1484 271
rect 920 259 924 263
rect 136 251 140 255
rect 224 251 228 255
rect 312 251 316 255
rect 400 251 404 255
rect 488 251 492 255
rect 576 251 580 255
rect 664 251 668 255
rect 744 251 748 255
rect 752 251 756 255
rect 824 251 828 255
rect 840 251 844 255
rect 912 251 916 255
rect 824 227 828 231
rect 912 227 916 231
rect 3464 443 3468 447
rect 3424 363 3428 367
rect 1968 347 1972 351
rect 2056 347 2060 351
rect 2144 347 2148 351
rect 2352 347 2356 351
rect 2840 347 2844 351
rect 3024 347 3028 351
rect 1880 319 1884 323
rect 1888 319 1892 323
rect 1968 319 1972 323
rect 1976 319 1980 323
rect 2056 319 2060 323
rect 2064 319 2068 323
rect 2144 319 2148 323
rect 2152 319 2156 323
rect 2264 319 2268 323
rect 2352 319 2356 323
rect 2384 319 2388 323
rect 2520 319 2524 323
rect 2672 319 2676 323
rect 2840 319 2844 323
rect 2848 319 2852 323
rect 3024 319 3028 323
rect 3032 319 3036 323
rect 3232 319 3236 323
rect 3432 319 3436 323
rect 1888 307 1892 311
rect 1960 307 1964 311
rect 1976 307 1980 311
rect 2048 307 2052 311
rect 2064 307 2068 311
rect 2136 307 2140 311
rect 2152 307 2156 311
rect 2224 307 2228 311
rect 2240 307 2244 311
rect 2352 307 2356 311
rect 2424 307 2428 311
rect 2464 307 2468 311
rect 2576 307 2580 311
rect 2688 307 2692 311
rect 2760 307 2764 311
rect 2800 307 2804 311
rect 2872 307 2876 311
rect 2912 307 2916 311
rect 2984 307 2988 311
rect 3032 307 3036 311
rect 3104 307 3108 311
rect 3152 307 3156 311
rect 1960 283 1964 287
rect 2048 283 2052 287
rect 2136 283 2140 287
rect 2224 283 2228 287
rect 2424 283 2428 287
rect 2760 283 2764 287
rect 2872 283 2876 287
rect 2984 283 2988 287
rect 3104 283 3108 287
rect 1576 267 1580 271
rect 1664 267 1668 271
rect 1672 267 1676 271
rect 928 251 932 255
rect 1016 251 1020 255
rect 1088 251 1092 255
rect 1104 251 1108 255
rect 1176 251 1180 255
rect 1192 251 1196 255
rect 1280 251 1284 255
rect 1368 251 1372 255
rect 1456 251 1460 255
rect 1544 251 1548 255
rect 1552 251 1556 255
rect 1616 251 1620 255
rect 1632 251 1636 255
rect 1720 251 1724 255
rect 1088 227 1092 231
rect 1176 227 1180 231
rect 1616 227 1620 231
rect 920 223 924 227
rect 1968 211 1972 215
rect 2056 211 2060 215
rect 2144 211 2148 215
rect 2256 211 2260 215
rect 2392 211 2396 215
rect 2528 211 2532 215
rect 2672 211 2676 215
rect 2944 211 2948 215
rect 3080 211 3084 215
rect 3216 211 3220 215
rect 3472 211 3476 215
rect 1888 183 1892 187
rect 1968 183 1972 187
rect 1976 183 1980 187
rect 2056 183 2060 187
rect 2064 183 2068 187
rect 2144 183 2148 187
rect 2152 183 2156 187
rect 2256 183 2260 187
rect 2264 183 2268 187
rect 2392 183 2396 187
rect 2400 183 2404 187
rect 2528 183 2532 187
rect 2536 183 2540 187
rect 2672 183 2676 187
rect 2680 183 2684 187
rect 2816 183 2820 187
rect 2944 183 2948 187
rect 2952 183 2956 187
rect 3080 183 3084 187
rect 3088 183 3092 187
rect 3216 183 3220 187
rect 3224 183 3228 187
rect 3360 183 3364 187
rect 3480 183 3484 187
rect 2776 139 2780 143
rect 2848 139 2852 143
rect 2864 139 2868 143
rect 2936 139 2940 143
rect 2952 139 2956 143
rect 3024 139 3028 143
rect 3040 139 3044 143
rect 3112 139 3116 143
rect 3128 139 3132 143
rect 3200 139 3204 143
rect 3216 139 3220 143
rect 3288 139 3292 143
rect 3304 139 3308 143
rect 3392 139 3396 143
rect 3472 139 3476 143
rect 3480 139 3484 143
rect 2848 115 2852 119
rect 2936 115 2940 119
rect 3024 115 3028 119
rect 3112 115 3116 119
rect 3200 115 3204 119
rect 3288 115 3292 119
<< m2 >>
rect 134 3659 140 3660
rect 134 3655 135 3659
rect 139 3655 140 3659
rect 134 3654 140 3655
rect 222 3659 228 3660
rect 222 3655 223 3659
rect 227 3655 228 3659
rect 222 3654 228 3655
rect 202 3651 208 3652
rect 110 3649 116 3650
rect 110 3645 111 3649
rect 115 3645 116 3649
rect 202 3647 203 3651
rect 207 3650 208 3651
rect 207 3648 241 3650
rect 1822 3649 1828 3650
rect 207 3647 208 3648
rect 202 3646 208 3647
rect 110 3644 116 3645
rect 1822 3645 1823 3649
rect 1827 3645 1828 3649
rect 1822 3644 1828 3645
rect 215 3635 221 3636
rect 215 3634 216 3635
rect 110 3632 116 3633
rect 197 3632 216 3634
rect 110 3628 111 3632
rect 115 3628 116 3632
rect 215 3631 216 3632
rect 220 3631 221 3635
rect 215 3630 221 3631
rect 1822 3632 1828 3633
rect 110 3627 116 3628
rect 1822 3628 1823 3632
rect 1827 3628 1828 3632
rect 1822 3627 1828 3628
rect 142 3619 148 3620
rect 142 3615 143 3619
rect 147 3615 148 3619
rect 142 3614 148 3615
rect 230 3619 236 3620
rect 230 3615 231 3619
rect 235 3615 236 3619
rect 230 3614 236 3615
rect 215 3607 221 3608
rect 215 3603 216 3607
rect 220 3606 221 3607
rect 223 3607 229 3608
rect 223 3606 224 3607
rect 220 3604 224 3606
rect 220 3603 221 3604
rect 215 3602 221 3603
rect 223 3603 224 3604
rect 228 3603 229 3607
rect 223 3602 229 3603
rect 135 3595 141 3596
rect 135 3591 136 3595
rect 140 3594 141 3595
rect 198 3595 204 3596
rect 198 3594 199 3595
rect 140 3592 199 3594
rect 140 3591 141 3592
rect 135 3590 141 3591
rect 198 3591 199 3592
rect 203 3591 204 3595
rect 198 3590 204 3591
rect 207 3595 213 3596
rect 207 3591 208 3595
rect 212 3594 213 3595
rect 223 3595 229 3596
rect 223 3594 224 3595
rect 212 3592 224 3594
rect 212 3591 213 3592
rect 207 3590 213 3591
rect 223 3591 224 3592
rect 228 3591 229 3595
rect 223 3590 229 3591
rect 295 3595 301 3596
rect 295 3591 296 3595
rect 300 3594 301 3595
rect 311 3595 317 3596
rect 311 3594 312 3595
rect 300 3592 312 3594
rect 300 3591 301 3592
rect 295 3590 301 3591
rect 311 3591 312 3592
rect 316 3591 317 3595
rect 311 3590 317 3591
rect 383 3595 389 3596
rect 383 3591 384 3595
rect 388 3594 389 3595
rect 399 3595 405 3596
rect 399 3594 400 3595
rect 388 3592 400 3594
rect 388 3591 389 3592
rect 383 3590 389 3591
rect 399 3591 400 3592
rect 404 3591 405 3595
rect 399 3590 405 3591
rect 471 3595 477 3596
rect 471 3591 472 3595
rect 476 3594 477 3595
rect 487 3595 493 3596
rect 487 3594 488 3595
rect 476 3592 488 3594
rect 476 3591 477 3592
rect 471 3590 477 3591
rect 487 3591 488 3592
rect 492 3591 493 3595
rect 487 3590 493 3591
rect 142 3585 148 3586
rect 142 3581 143 3585
rect 147 3581 148 3585
rect 142 3580 148 3581
rect 230 3585 236 3586
rect 230 3581 231 3585
rect 235 3581 236 3585
rect 230 3580 236 3581
rect 318 3585 324 3586
rect 318 3581 319 3585
rect 323 3581 324 3585
rect 318 3580 324 3581
rect 406 3585 412 3586
rect 406 3581 407 3585
rect 411 3581 412 3585
rect 406 3580 412 3581
rect 494 3585 500 3586
rect 494 3581 495 3585
rect 499 3581 500 3585
rect 494 3580 500 3581
rect 1886 3583 1892 3584
rect 1886 3579 1887 3583
rect 1891 3579 1892 3583
rect 1886 3578 1892 3579
rect 1974 3583 1980 3584
rect 1974 3579 1975 3583
rect 1979 3579 1980 3583
rect 1974 3578 1980 3579
rect 2062 3583 2068 3584
rect 2062 3579 2063 3583
rect 2067 3579 2068 3583
rect 2062 3578 2068 3579
rect 2150 3583 2156 3584
rect 2150 3579 2151 3583
rect 2155 3579 2156 3583
rect 2150 3578 2156 3579
rect 2238 3583 2244 3584
rect 2238 3579 2239 3583
rect 2243 3579 2244 3583
rect 2238 3578 2244 3579
rect 2326 3583 2332 3584
rect 2326 3579 2327 3583
rect 2331 3579 2332 3583
rect 2326 3578 2332 3579
rect 2430 3583 2436 3584
rect 2430 3579 2431 3583
rect 2435 3579 2436 3583
rect 2430 3578 2436 3579
rect 2534 3583 2540 3584
rect 2534 3579 2535 3583
rect 2539 3579 2540 3583
rect 2534 3578 2540 3579
rect 2630 3583 2636 3584
rect 2630 3579 2631 3583
rect 2635 3579 2636 3583
rect 2630 3578 2636 3579
rect 2726 3583 2732 3584
rect 2726 3579 2727 3583
rect 2731 3579 2732 3583
rect 2726 3578 2732 3579
rect 2822 3583 2828 3584
rect 2822 3579 2823 3583
rect 2827 3579 2828 3583
rect 2822 3578 2828 3579
rect 2918 3583 2924 3584
rect 2918 3579 2919 3583
rect 2923 3579 2924 3583
rect 2918 3578 2924 3579
rect 3014 3583 3020 3584
rect 3014 3579 3015 3583
rect 3019 3579 3020 3583
rect 3014 3578 3020 3579
rect 3118 3583 3124 3584
rect 3118 3579 3119 3583
rect 3123 3579 3124 3583
rect 3118 3578 3124 3579
rect 3222 3583 3228 3584
rect 3222 3579 3223 3583
rect 3227 3579 3228 3583
rect 3222 3578 3228 3579
rect 2498 3575 2504 3576
rect 1862 3573 1868 3574
rect 110 3572 116 3573
rect 1822 3572 1828 3573
rect 110 3568 111 3572
rect 115 3568 116 3572
rect 207 3571 213 3572
rect 207 3570 208 3571
rect 197 3568 208 3570
rect 110 3567 116 3568
rect 207 3567 208 3568
rect 212 3567 213 3571
rect 295 3571 301 3572
rect 295 3570 296 3571
rect 285 3568 296 3570
rect 207 3566 213 3567
rect 295 3567 296 3568
rect 300 3567 301 3571
rect 383 3571 389 3572
rect 383 3570 384 3571
rect 373 3568 384 3570
rect 295 3566 301 3567
rect 383 3567 384 3568
rect 388 3567 389 3571
rect 471 3571 477 3572
rect 471 3570 472 3571
rect 461 3568 472 3570
rect 383 3566 389 3567
rect 471 3567 472 3568
rect 476 3567 477 3571
rect 1822 3568 1823 3572
rect 1827 3568 1828 3572
rect 1862 3569 1863 3573
rect 1867 3569 1868 3573
rect 2498 3571 2499 3575
rect 2503 3574 2504 3575
rect 2503 3572 2553 3574
rect 3574 3573 3580 3574
rect 2503 3571 2504 3572
rect 2498 3570 2504 3571
rect 1862 3568 1868 3569
rect 3574 3569 3575 3573
rect 3579 3569 3580 3573
rect 3574 3568 3580 3569
rect 1822 3567 1828 3568
rect 471 3566 477 3567
rect 1967 3559 1973 3560
rect 1967 3558 1968 3559
rect 1862 3556 1868 3557
rect 1949 3556 1968 3558
rect 110 3555 116 3556
rect 110 3551 111 3555
rect 115 3551 116 3555
rect 1822 3555 1828 3556
rect 110 3550 116 3551
rect 468 3552 505 3554
rect 134 3545 140 3546
rect 134 3541 135 3545
rect 139 3541 140 3545
rect 134 3540 140 3541
rect 222 3545 228 3546
rect 222 3541 223 3545
rect 227 3541 228 3545
rect 222 3540 228 3541
rect 310 3545 316 3546
rect 310 3541 311 3545
rect 315 3541 316 3545
rect 310 3540 316 3541
rect 398 3545 404 3546
rect 398 3541 399 3545
rect 403 3541 404 3545
rect 398 3540 404 3541
rect 266 3539 272 3540
rect 266 3535 267 3539
rect 271 3538 272 3539
rect 468 3538 470 3552
rect 1822 3551 1823 3555
rect 1827 3551 1828 3555
rect 1862 3552 1863 3556
rect 1867 3552 1868 3556
rect 1967 3555 1968 3556
rect 1972 3555 1973 3559
rect 2055 3559 2061 3560
rect 2055 3558 2056 3559
rect 2037 3556 2056 3558
rect 1967 3554 1973 3555
rect 2055 3555 2056 3556
rect 2060 3555 2061 3559
rect 2143 3559 2149 3560
rect 2143 3558 2144 3559
rect 2125 3556 2144 3558
rect 2055 3554 2061 3555
rect 2143 3555 2144 3556
rect 2148 3555 2149 3559
rect 2231 3559 2237 3560
rect 2231 3558 2232 3559
rect 2213 3556 2232 3558
rect 2143 3554 2149 3555
rect 2231 3555 2232 3556
rect 2236 3555 2237 3559
rect 2311 3559 2317 3560
rect 2311 3558 2312 3559
rect 2301 3556 2312 3558
rect 2231 3554 2237 3555
rect 2311 3555 2312 3556
rect 2316 3555 2317 3559
rect 2423 3559 2429 3560
rect 2423 3558 2424 3559
rect 2389 3556 2424 3558
rect 2311 3554 2317 3555
rect 2423 3555 2424 3556
rect 2428 3555 2429 3559
rect 2527 3559 2533 3560
rect 2527 3558 2528 3559
rect 2493 3556 2528 3558
rect 2423 3554 2429 3555
rect 2527 3555 2528 3556
rect 2532 3555 2533 3559
rect 2719 3559 2725 3560
rect 2719 3558 2720 3559
rect 2693 3556 2720 3558
rect 2527 3554 2533 3555
rect 2719 3555 2720 3556
rect 2724 3555 2725 3559
rect 2815 3559 2821 3560
rect 2815 3558 2816 3559
rect 2789 3556 2816 3558
rect 2719 3554 2725 3555
rect 2815 3555 2816 3556
rect 2820 3555 2821 3559
rect 2911 3559 2917 3560
rect 2911 3558 2912 3559
rect 2885 3556 2912 3558
rect 2815 3554 2821 3555
rect 2911 3555 2912 3556
rect 2916 3555 2917 3559
rect 3007 3559 3013 3560
rect 3007 3558 3008 3559
rect 2981 3556 3008 3558
rect 2911 3554 2917 3555
rect 3007 3555 3008 3556
rect 3012 3555 3013 3559
rect 3111 3559 3117 3560
rect 3111 3558 3112 3559
rect 3077 3556 3112 3558
rect 3007 3554 3013 3555
rect 3111 3555 3112 3556
rect 3116 3555 3117 3559
rect 3186 3559 3192 3560
rect 3186 3558 3187 3559
rect 3181 3556 3187 3558
rect 3111 3554 3117 3555
rect 3186 3555 3187 3556
rect 3191 3555 3192 3559
rect 3186 3554 3192 3555
rect 3214 3559 3220 3560
rect 3214 3555 3215 3559
rect 3219 3558 3220 3559
rect 3219 3556 3249 3558
rect 3574 3556 3580 3557
rect 3219 3555 3220 3556
rect 3214 3554 3220 3555
rect 1862 3551 1868 3552
rect 3574 3552 3575 3556
rect 3579 3552 3580 3556
rect 3574 3551 3580 3552
rect 1822 3550 1828 3551
rect 486 3545 492 3546
rect 486 3541 487 3545
rect 491 3541 492 3545
rect 486 3540 492 3541
rect 1894 3543 1900 3544
rect 1894 3539 1895 3543
rect 1899 3539 1900 3543
rect 1894 3538 1900 3539
rect 1982 3543 1988 3544
rect 1982 3539 1983 3543
rect 1987 3539 1988 3543
rect 1982 3538 1988 3539
rect 2070 3543 2076 3544
rect 2070 3539 2071 3543
rect 2075 3539 2076 3543
rect 2070 3538 2076 3539
rect 2158 3543 2164 3544
rect 2158 3539 2159 3543
rect 2163 3539 2164 3543
rect 2158 3538 2164 3539
rect 2246 3543 2252 3544
rect 2246 3539 2247 3543
rect 2251 3539 2252 3543
rect 2246 3538 2252 3539
rect 2334 3543 2340 3544
rect 2334 3539 2335 3543
rect 2339 3539 2340 3543
rect 2334 3538 2340 3539
rect 2438 3543 2444 3544
rect 2438 3539 2439 3543
rect 2443 3539 2444 3543
rect 2438 3538 2444 3539
rect 2542 3543 2548 3544
rect 2542 3539 2543 3543
rect 2547 3539 2548 3543
rect 2542 3538 2548 3539
rect 2638 3543 2644 3544
rect 2638 3539 2639 3543
rect 2643 3539 2644 3543
rect 2638 3538 2644 3539
rect 2734 3543 2740 3544
rect 2734 3539 2735 3543
rect 2739 3539 2740 3543
rect 2734 3538 2740 3539
rect 2830 3543 2836 3544
rect 2830 3539 2831 3543
rect 2835 3539 2836 3543
rect 2830 3538 2836 3539
rect 2926 3543 2932 3544
rect 2926 3539 2927 3543
rect 2931 3539 2932 3543
rect 2926 3538 2932 3539
rect 3022 3543 3028 3544
rect 3022 3539 3023 3543
rect 3027 3539 3028 3543
rect 3022 3538 3028 3539
rect 3126 3543 3132 3544
rect 3126 3539 3127 3543
rect 3131 3539 3132 3543
rect 3126 3538 3132 3539
rect 3230 3543 3236 3544
rect 3230 3539 3231 3543
rect 3235 3539 3236 3543
rect 3230 3538 3236 3539
rect 271 3536 470 3538
rect 271 3535 272 3536
rect 266 3534 272 3535
rect 1886 3531 1893 3532
rect 1886 3527 1887 3531
rect 1892 3527 1893 3531
rect 1886 3526 1893 3527
rect 1967 3531 1973 3532
rect 1967 3527 1968 3531
rect 1972 3530 1973 3531
rect 1975 3531 1981 3532
rect 1975 3530 1976 3531
rect 1972 3528 1976 3530
rect 1972 3527 1973 3528
rect 1967 3526 1973 3527
rect 1975 3527 1976 3528
rect 1980 3527 1981 3531
rect 1975 3526 1981 3527
rect 2055 3531 2061 3532
rect 2055 3527 2056 3531
rect 2060 3530 2061 3531
rect 2063 3531 2069 3532
rect 2063 3530 2064 3531
rect 2060 3528 2064 3530
rect 2060 3527 2061 3528
rect 2055 3526 2061 3527
rect 2063 3527 2064 3528
rect 2068 3527 2069 3531
rect 2063 3526 2069 3527
rect 2143 3531 2149 3532
rect 2143 3527 2144 3531
rect 2148 3530 2149 3531
rect 2151 3531 2157 3532
rect 2151 3530 2152 3531
rect 2148 3528 2152 3530
rect 2148 3527 2149 3528
rect 2143 3526 2149 3527
rect 2151 3527 2152 3528
rect 2156 3527 2157 3531
rect 2151 3526 2157 3527
rect 2231 3531 2237 3532
rect 2231 3527 2232 3531
rect 2236 3530 2237 3531
rect 2239 3531 2245 3532
rect 2239 3530 2240 3531
rect 2236 3528 2240 3530
rect 2236 3527 2237 3528
rect 2231 3526 2237 3527
rect 2239 3527 2240 3528
rect 2244 3527 2245 3531
rect 2239 3526 2245 3527
rect 2311 3531 2317 3532
rect 2311 3527 2312 3531
rect 2316 3530 2317 3531
rect 2327 3531 2333 3532
rect 2327 3530 2328 3531
rect 2316 3528 2328 3530
rect 2316 3527 2317 3528
rect 2311 3526 2317 3527
rect 2327 3527 2328 3528
rect 2332 3527 2333 3531
rect 2327 3526 2333 3527
rect 2423 3531 2429 3532
rect 2423 3527 2424 3531
rect 2428 3530 2429 3531
rect 2431 3531 2437 3532
rect 2431 3530 2432 3531
rect 2428 3528 2432 3530
rect 2428 3527 2429 3528
rect 2423 3526 2429 3527
rect 2431 3527 2432 3528
rect 2436 3527 2437 3531
rect 2431 3526 2437 3527
rect 2527 3531 2533 3532
rect 2527 3527 2528 3531
rect 2532 3530 2533 3531
rect 2535 3531 2541 3532
rect 2535 3530 2536 3531
rect 2532 3528 2536 3530
rect 2532 3527 2533 3528
rect 2527 3526 2533 3527
rect 2535 3527 2536 3528
rect 2540 3527 2541 3531
rect 2535 3526 2541 3527
rect 2631 3531 2637 3532
rect 2631 3527 2632 3531
rect 2636 3530 2637 3531
rect 2639 3531 2645 3532
rect 2639 3530 2640 3531
rect 2636 3528 2640 3530
rect 2636 3527 2637 3528
rect 2631 3526 2637 3527
rect 2639 3527 2640 3528
rect 2644 3527 2645 3531
rect 2639 3526 2645 3527
rect 2719 3531 2725 3532
rect 2719 3527 2720 3531
rect 2724 3530 2725 3531
rect 2727 3531 2733 3532
rect 2727 3530 2728 3531
rect 2724 3528 2728 3530
rect 2724 3527 2725 3528
rect 2719 3526 2725 3527
rect 2727 3527 2728 3528
rect 2732 3527 2733 3531
rect 2727 3526 2733 3527
rect 2815 3531 2821 3532
rect 2815 3527 2816 3531
rect 2820 3530 2821 3531
rect 2823 3531 2829 3532
rect 2823 3530 2824 3531
rect 2820 3528 2824 3530
rect 2820 3527 2821 3528
rect 2815 3526 2821 3527
rect 2823 3527 2824 3528
rect 2828 3527 2829 3531
rect 2823 3526 2829 3527
rect 2911 3531 2917 3532
rect 2911 3527 2912 3531
rect 2916 3530 2917 3531
rect 2919 3531 2925 3532
rect 2919 3530 2920 3531
rect 2916 3528 2920 3530
rect 2916 3527 2917 3528
rect 2911 3526 2917 3527
rect 2919 3527 2920 3528
rect 2924 3527 2925 3531
rect 2919 3526 2925 3527
rect 3007 3531 3013 3532
rect 3007 3527 3008 3531
rect 3012 3530 3013 3531
rect 3015 3531 3021 3532
rect 3015 3530 3016 3531
rect 3012 3528 3016 3530
rect 3012 3527 3013 3528
rect 3007 3526 3013 3527
rect 3015 3527 3016 3528
rect 3020 3527 3021 3531
rect 3015 3526 3021 3527
rect 3111 3531 3117 3532
rect 3111 3527 3112 3531
rect 3116 3530 3117 3531
rect 3119 3531 3125 3532
rect 3119 3530 3120 3531
rect 3116 3528 3120 3530
rect 3116 3527 3117 3528
rect 3111 3526 3117 3527
rect 3119 3527 3120 3528
rect 3124 3527 3125 3531
rect 3119 3526 3125 3527
rect 3186 3531 3192 3532
rect 3186 3527 3187 3531
rect 3191 3530 3192 3531
rect 3223 3531 3229 3532
rect 3223 3530 3224 3531
rect 3191 3528 3224 3530
rect 3191 3527 3192 3528
rect 3186 3526 3192 3527
rect 3223 3527 3224 3528
rect 3228 3527 3229 3531
rect 3223 3526 3229 3527
rect 246 3523 252 3524
rect 246 3519 247 3523
rect 251 3519 252 3523
rect 246 3518 252 3519
rect 374 3523 380 3524
rect 374 3519 375 3523
rect 379 3519 380 3523
rect 374 3518 380 3519
rect 502 3523 508 3524
rect 502 3519 503 3523
rect 507 3519 508 3523
rect 502 3518 508 3519
rect 622 3523 628 3524
rect 622 3519 623 3523
rect 627 3519 628 3523
rect 622 3518 628 3519
rect 742 3523 748 3524
rect 742 3519 743 3523
rect 747 3519 748 3523
rect 742 3518 748 3519
rect 862 3523 868 3524
rect 862 3519 863 3523
rect 867 3519 868 3523
rect 862 3518 868 3519
rect 974 3523 980 3524
rect 974 3519 975 3523
rect 979 3519 980 3523
rect 974 3518 980 3519
rect 1078 3523 1084 3524
rect 1078 3519 1079 3523
rect 1083 3519 1084 3523
rect 1078 3518 1084 3519
rect 1174 3523 1180 3524
rect 1174 3519 1175 3523
rect 1179 3519 1180 3523
rect 1174 3518 1180 3519
rect 1270 3523 1276 3524
rect 1270 3519 1271 3523
rect 1275 3519 1276 3523
rect 1270 3518 1276 3519
rect 1366 3523 1372 3524
rect 1366 3519 1367 3523
rect 1371 3519 1372 3523
rect 1366 3518 1372 3519
rect 1470 3523 1476 3524
rect 1470 3519 1471 3523
rect 1475 3519 1476 3523
rect 1470 3518 1476 3519
rect 1574 3523 1580 3524
rect 1574 3519 1575 3523
rect 1579 3519 1580 3523
rect 1574 3518 1580 3519
rect 1887 3519 1893 3520
rect 1538 3515 1544 3516
rect 110 3513 116 3514
rect 110 3509 111 3513
rect 115 3509 116 3513
rect 1538 3511 1539 3515
rect 1543 3514 1544 3515
rect 1887 3515 1888 3519
rect 1892 3518 1893 3519
rect 1962 3519 1968 3520
rect 1962 3518 1963 3519
rect 1892 3516 1963 3518
rect 1892 3515 1893 3516
rect 1887 3514 1893 3515
rect 1962 3515 1963 3516
rect 1967 3515 1968 3519
rect 1962 3514 1968 3515
rect 1975 3519 1981 3520
rect 1975 3515 1976 3519
rect 1980 3518 1981 3519
rect 1990 3519 1996 3520
rect 1990 3518 1991 3519
rect 1980 3516 1991 3518
rect 1980 3515 1981 3516
rect 1975 3514 1981 3515
rect 1990 3515 1991 3516
rect 1995 3515 1996 3519
rect 1990 3514 1996 3515
rect 2095 3519 2101 3520
rect 2095 3515 2096 3519
rect 2100 3518 2101 3519
rect 2110 3519 2116 3520
rect 2110 3518 2111 3519
rect 2100 3516 2111 3518
rect 2100 3515 2101 3516
rect 2095 3514 2101 3515
rect 2110 3515 2111 3516
rect 2115 3515 2116 3519
rect 2110 3514 2116 3515
rect 2167 3519 2173 3520
rect 2167 3515 2168 3519
rect 2172 3518 2173 3519
rect 2223 3519 2229 3520
rect 2223 3518 2224 3519
rect 2172 3516 2224 3518
rect 2172 3515 2173 3516
rect 2167 3514 2173 3515
rect 2223 3515 2224 3516
rect 2228 3515 2229 3519
rect 2223 3514 2229 3515
rect 2290 3519 2296 3520
rect 2290 3515 2291 3519
rect 2295 3518 2296 3519
rect 2359 3519 2365 3520
rect 2359 3518 2360 3519
rect 2295 3516 2360 3518
rect 2295 3515 2296 3516
rect 2290 3514 2296 3515
rect 2359 3515 2360 3516
rect 2364 3515 2365 3519
rect 2359 3514 2365 3515
rect 2439 3519 2445 3520
rect 2439 3515 2440 3519
rect 2444 3518 2445 3519
rect 2503 3519 2509 3520
rect 2503 3518 2504 3519
rect 2444 3516 2504 3518
rect 2444 3515 2445 3516
rect 2439 3514 2445 3515
rect 2503 3515 2504 3516
rect 2508 3515 2509 3519
rect 2503 3514 2509 3515
rect 2647 3519 2653 3520
rect 2647 3515 2648 3519
rect 2652 3518 2653 3519
rect 2722 3519 2728 3520
rect 2722 3518 2723 3519
rect 2652 3516 2723 3518
rect 2652 3515 2653 3516
rect 2647 3514 2653 3515
rect 2722 3515 2723 3516
rect 2727 3515 2728 3519
rect 2722 3514 2728 3515
rect 2783 3519 2789 3520
rect 2783 3515 2784 3519
rect 2788 3518 2789 3519
rect 2798 3519 2804 3520
rect 2798 3518 2799 3519
rect 2788 3516 2799 3518
rect 2788 3515 2789 3516
rect 2783 3514 2789 3515
rect 2798 3515 2799 3516
rect 2803 3515 2804 3519
rect 2798 3514 2804 3515
rect 2927 3519 2933 3520
rect 2927 3515 2928 3519
rect 2932 3518 2933 3519
rect 3002 3519 3008 3520
rect 3002 3518 3003 3519
rect 2932 3516 3003 3518
rect 2932 3515 2933 3516
rect 2927 3514 2933 3515
rect 3002 3515 3003 3516
rect 3007 3515 3008 3519
rect 3002 3514 3008 3515
rect 3071 3519 3077 3520
rect 3071 3515 3072 3519
rect 3076 3518 3077 3519
rect 3182 3519 3188 3520
rect 3182 3518 3183 3519
rect 3076 3516 3183 3518
rect 3076 3515 3077 3516
rect 3071 3514 3077 3515
rect 3182 3515 3183 3516
rect 3187 3515 3188 3519
rect 3182 3514 3188 3515
rect 3214 3519 3221 3520
rect 3214 3515 3215 3519
rect 3220 3515 3221 3519
rect 3214 3514 3221 3515
rect 1543 3512 1593 3514
rect 1822 3513 1828 3514
rect 1543 3511 1544 3512
rect 1538 3510 1544 3511
rect 110 3508 116 3509
rect 1822 3509 1823 3513
rect 1827 3509 1828 3513
rect 1822 3508 1828 3509
rect 1894 3509 1900 3510
rect 1894 3505 1895 3509
rect 1899 3505 1900 3509
rect 1894 3504 1900 3505
rect 1982 3509 1988 3510
rect 1982 3505 1983 3509
rect 1987 3505 1988 3509
rect 1982 3504 1988 3505
rect 2102 3509 2108 3510
rect 2102 3505 2103 3509
rect 2107 3505 2108 3509
rect 2102 3504 2108 3505
rect 2230 3509 2236 3510
rect 2230 3505 2231 3509
rect 2235 3505 2236 3509
rect 2230 3504 2236 3505
rect 2366 3509 2372 3510
rect 2366 3505 2367 3509
rect 2371 3505 2372 3509
rect 2366 3504 2372 3505
rect 2510 3509 2516 3510
rect 2510 3505 2511 3509
rect 2515 3505 2516 3509
rect 2510 3504 2516 3505
rect 2654 3509 2660 3510
rect 2654 3505 2655 3509
rect 2659 3505 2660 3509
rect 2654 3504 2660 3505
rect 2790 3509 2796 3510
rect 2790 3505 2791 3509
rect 2795 3505 2796 3509
rect 2790 3504 2796 3505
rect 2934 3509 2940 3510
rect 2934 3505 2935 3509
rect 2939 3505 2940 3509
rect 2934 3504 2940 3505
rect 3078 3509 3084 3510
rect 3078 3505 3079 3509
rect 3083 3505 3084 3509
rect 3078 3504 3084 3505
rect 3222 3509 3228 3510
rect 3222 3505 3223 3509
rect 3227 3505 3228 3509
rect 3222 3504 3228 3505
rect 367 3499 373 3500
rect 367 3498 368 3499
rect 110 3496 116 3497
rect 309 3496 368 3498
rect 110 3492 111 3496
rect 115 3492 116 3496
rect 367 3495 368 3496
rect 372 3495 373 3499
rect 495 3499 501 3500
rect 495 3498 496 3499
rect 437 3496 496 3498
rect 367 3494 373 3495
rect 495 3495 496 3496
rect 500 3495 501 3499
rect 570 3499 576 3500
rect 570 3498 571 3499
rect 565 3496 571 3498
rect 495 3494 501 3495
rect 570 3495 571 3496
rect 575 3495 576 3499
rect 734 3499 740 3500
rect 734 3498 735 3499
rect 685 3496 735 3498
rect 570 3494 576 3495
rect 734 3495 735 3496
rect 739 3495 740 3499
rect 855 3499 861 3500
rect 855 3498 856 3499
rect 805 3496 856 3498
rect 734 3494 740 3495
rect 855 3495 856 3496
rect 860 3495 861 3499
rect 966 3499 972 3500
rect 966 3498 967 3499
rect 925 3496 967 3498
rect 855 3494 861 3495
rect 966 3495 967 3496
rect 971 3495 972 3499
rect 1071 3499 1077 3500
rect 1071 3498 1072 3499
rect 1037 3496 1072 3498
rect 966 3494 972 3495
rect 1071 3495 1072 3496
rect 1076 3495 1077 3499
rect 1167 3499 1173 3500
rect 1167 3498 1168 3499
rect 1141 3496 1168 3498
rect 1071 3494 1077 3495
rect 1167 3495 1168 3496
rect 1172 3495 1173 3499
rect 1263 3499 1269 3500
rect 1263 3498 1264 3499
rect 1237 3496 1264 3498
rect 1167 3494 1173 3495
rect 1263 3495 1264 3496
rect 1268 3495 1269 3499
rect 1359 3499 1365 3500
rect 1359 3498 1360 3499
rect 1333 3496 1360 3498
rect 1263 3494 1269 3495
rect 1359 3495 1360 3496
rect 1364 3495 1365 3499
rect 1463 3499 1469 3500
rect 1463 3498 1464 3499
rect 1429 3496 1464 3498
rect 1359 3494 1365 3495
rect 1463 3495 1464 3496
rect 1468 3495 1469 3499
rect 1567 3499 1573 3500
rect 1567 3498 1568 3499
rect 1533 3496 1568 3498
rect 1463 3494 1469 3495
rect 1567 3495 1568 3496
rect 1572 3495 1573 3499
rect 1567 3494 1573 3495
rect 1822 3496 1828 3497
rect 110 3491 116 3492
rect 1822 3492 1823 3496
rect 1827 3492 1828 3496
rect 1822 3491 1828 3492
rect 1862 3496 1868 3497
rect 3574 3496 3580 3497
rect 1862 3492 1863 3496
rect 1867 3492 1868 3496
rect 2167 3495 2173 3496
rect 2167 3494 2168 3495
rect 2157 3492 2168 3494
rect 1862 3491 1868 3492
rect 1886 3491 1892 3492
rect 1886 3487 1887 3491
rect 1891 3490 1892 3491
rect 1962 3491 1968 3492
rect 1891 3488 1913 3490
rect 1891 3487 1892 3488
rect 1886 3486 1892 3487
rect 1962 3487 1963 3491
rect 1967 3490 1968 3491
rect 2167 3491 2168 3492
rect 2172 3491 2173 3495
rect 2290 3495 2296 3496
rect 2290 3494 2291 3495
rect 2285 3492 2291 3494
rect 2167 3490 2173 3491
rect 2290 3491 2291 3492
rect 2295 3491 2296 3495
rect 2439 3495 2445 3496
rect 2439 3494 2440 3495
rect 2421 3492 2440 3494
rect 2290 3490 2296 3491
rect 2439 3491 2440 3492
rect 2444 3491 2445 3495
rect 3574 3492 3575 3496
rect 3579 3492 3580 3496
rect 2439 3490 2445 3491
rect 2639 3491 2645 3492
rect 1967 3488 2001 3490
rect 1967 3487 1968 3488
rect 1962 3486 1968 3487
rect 2639 3487 2640 3491
rect 2644 3490 2645 3491
rect 2722 3491 2728 3492
rect 2644 3488 2673 3490
rect 2644 3487 2645 3488
rect 2639 3486 2645 3487
rect 2722 3487 2723 3491
rect 2727 3490 2728 3491
rect 3002 3491 3008 3492
rect 2727 3488 2809 3490
rect 2727 3487 2728 3488
rect 2722 3486 2728 3487
rect 3002 3487 3003 3491
rect 3007 3490 3008 3491
rect 3182 3491 3188 3492
rect 3574 3491 3580 3492
rect 3007 3488 3097 3490
rect 3007 3487 3008 3488
rect 3002 3486 3008 3487
rect 3182 3487 3183 3491
rect 3187 3490 3188 3491
rect 3187 3488 3241 3490
rect 3187 3487 3188 3488
rect 3182 3486 3188 3487
rect 254 3483 260 3484
rect 254 3479 255 3483
rect 259 3479 260 3483
rect 254 3478 260 3479
rect 382 3483 388 3484
rect 382 3479 383 3483
rect 387 3479 388 3483
rect 382 3478 388 3479
rect 510 3483 516 3484
rect 510 3479 511 3483
rect 515 3479 516 3483
rect 510 3478 516 3479
rect 630 3483 636 3484
rect 630 3479 631 3483
rect 635 3479 636 3483
rect 630 3478 636 3479
rect 750 3483 756 3484
rect 750 3479 751 3483
rect 755 3479 756 3483
rect 750 3478 756 3479
rect 870 3483 876 3484
rect 870 3479 871 3483
rect 875 3479 876 3483
rect 870 3478 876 3479
rect 982 3483 988 3484
rect 982 3479 983 3483
rect 987 3479 988 3483
rect 982 3478 988 3479
rect 1086 3483 1092 3484
rect 1086 3479 1087 3483
rect 1091 3479 1092 3483
rect 1086 3478 1092 3479
rect 1182 3483 1188 3484
rect 1182 3479 1183 3483
rect 1187 3479 1188 3483
rect 1182 3478 1188 3479
rect 1278 3483 1284 3484
rect 1278 3479 1279 3483
rect 1283 3479 1284 3483
rect 1278 3478 1284 3479
rect 1374 3483 1380 3484
rect 1374 3479 1375 3483
rect 1379 3479 1380 3483
rect 1374 3478 1380 3479
rect 1478 3483 1484 3484
rect 1478 3479 1479 3483
rect 1483 3479 1484 3483
rect 1478 3478 1484 3479
rect 1582 3483 1588 3484
rect 1582 3479 1583 3483
rect 1587 3479 1588 3483
rect 1582 3478 1588 3479
rect 1862 3479 1868 3480
rect 570 3475 576 3476
rect 247 3471 253 3472
rect 247 3467 248 3471
rect 252 3470 253 3471
rect 266 3471 272 3472
rect 266 3470 267 3471
rect 252 3468 267 3470
rect 252 3467 253 3468
rect 247 3466 253 3467
rect 266 3467 267 3468
rect 271 3467 272 3471
rect 266 3466 272 3467
rect 367 3471 373 3472
rect 367 3467 368 3471
rect 372 3470 373 3471
rect 375 3471 381 3472
rect 375 3470 376 3471
rect 372 3468 376 3470
rect 372 3467 373 3468
rect 367 3466 373 3467
rect 375 3467 376 3468
rect 380 3467 381 3471
rect 375 3466 381 3467
rect 495 3471 501 3472
rect 495 3467 496 3471
rect 500 3470 501 3471
rect 503 3471 509 3472
rect 503 3470 504 3471
rect 500 3468 504 3470
rect 500 3467 501 3468
rect 495 3466 501 3467
rect 503 3467 504 3468
rect 508 3467 509 3471
rect 570 3471 571 3475
rect 575 3474 576 3475
rect 1862 3475 1863 3479
rect 1867 3475 1868 3479
rect 1862 3474 1868 3475
rect 2886 3479 2892 3480
rect 2886 3475 2887 3479
rect 2891 3478 2892 3479
rect 3574 3479 3580 3480
rect 2891 3476 2945 3478
rect 2891 3475 2892 3476
rect 2886 3474 2892 3475
rect 3574 3475 3575 3479
rect 3579 3475 3580 3479
rect 3574 3474 3580 3475
rect 575 3472 627 3474
rect 575 3471 576 3472
rect 570 3470 576 3471
rect 623 3471 629 3472
rect 503 3466 509 3467
rect 623 3467 624 3471
rect 628 3467 629 3471
rect 623 3466 629 3467
rect 743 3471 749 3472
rect 743 3467 744 3471
rect 748 3470 749 3471
rect 823 3471 829 3472
rect 823 3470 824 3471
rect 748 3468 824 3470
rect 748 3467 749 3468
rect 743 3466 749 3467
rect 823 3467 824 3468
rect 828 3467 829 3471
rect 823 3466 829 3467
rect 855 3471 861 3472
rect 855 3467 856 3471
rect 860 3470 861 3471
rect 863 3471 869 3472
rect 863 3470 864 3471
rect 860 3468 864 3470
rect 860 3467 861 3468
rect 855 3466 861 3467
rect 863 3467 864 3468
rect 868 3467 869 3471
rect 863 3466 869 3467
rect 966 3471 972 3472
rect 966 3467 967 3471
rect 971 3470 972 3471
rect 975 3471 981 3472
rect 975 3470 976 3471
rect 971 3468 976 3470
rect 971 3467 972 3468
rect 966 3466 972 3467
rect 975 3467 976 3468
rect 980 3467 981 3471
rect 975 3466 981 3467
rect 1071 3471 1077 3472
rect 1071 3467 1072 3471
rect 1076 3470 1077 3471
rect 1079 3471 1085 3472
rect 1079 3470 1080 3471
rect 1076 3468 1080 3470
rect 1076 3467 1077 3468
rect 1071 3466 1077 3467
rect 1079 3467 1080 3468
rect 1084 3467 1085 3471
rect 1079 3466 1085 3467
rect 1167 3471 1173 3472
rect 1167 3467 1168 3471
rect 1172 3470 1173 3471
rect 1175 3471 1181 3472
rect 1175 3470 1176 3471
rect 1172 3468 1176 3470
rect 1172 3467 1173 3468
rect 1167 3466 1173 3467
rect 1175 3467 1176 3468
rect 1180 3467 1181 3471
rect 1175 3466 1181 3467
rect 1263 3471 1269 3472
rect 1263 3467 1264 3471
rect 1268 3470 1269 3471
rect 1271 3471 1277 3472
rect 1271 3470 1272 3471
rect 1268 3468 1272 3470
rect 1268 3467 1269 3468
rect 1263 3466 1269 3467
rect 1271 3467 1272 3468
rect 1276 3467 1277 3471
rect 1271 3466 1277 3467
rect 1359 3471 1365 3472
rect 1359 3467 1360 3471
rect 1364 3470 1365 3471
rect 1367 3471 1373 3472
rect 1367 3470 1368 3471
rect 1364 3468 1368 3470
rect 1364 3467 1365 3468
rect 1359 3466 1365 3467
rect 1367 3467 1368 3468
rect 1372 3467 1373 3471
rect 1367 3466 1373 3467
rect 1463 3471 1469 3472
rect 1463 3467 1464 3471
rect 1468 3470 1469 3471
rect 1471 3471 1477 3472
rect 1471 3470 1472 3471
rect 1468 3468 1472 3470
rect 1468 3467 1469 3468
rect 1463 3466 1469 3467
rect 1471 3467 1472 3468
rect 1476 3467 1477 3471
rect 1471 3466 1477 3467
rect 1567 3471 1573 3472
rect 1567 3467 1568 3471
rect 1572 3470 1573 3471
rect 1575 3471 1581 3472
rect 1575 3470 1576 3471
rect 1572 3468 1576 3470
rect 1572 3467 1573 3468
rect 1567 3466 1573 3467
rect 1575 3467 1576 3468
rect 1580 3467 1581 3471
rect 1575 3466 1581 3467
rect 1886 3469 1892 3470
rect 576 3464 621 3466
rect 1886 3465 1887 3469
rect 1891 3465 1892 3469
rect 1886 3464 1892 3465
rect 1974 3469 1980 3470
rect 1974 3465 1975 3469
rect 1979 3465 1980 3469
rect 1974 3464 1980 3465
rect 2094 3469 2100 3470
rect 2094 3465 2095 3469
rect 2099 3465 2100 3469
rect 2094 3464 2100 3465
rect 2222 3469 2228 3470
rect 2222 3465 2223 3469
rect 2227 3465 2228 3469
rect 2222 3464 2228 3465
rect 2358 3469 2364 3470
rect 2358 3465 2359 3469
rect 2363 3465 2364 3469
rect 2358 3464 2364 3465
rect 2502 3469 2508 3470
rect 2502 3465 2503 3469
rect 2507 3465 2508 3469
rect 2502 3464 2508 3465
rect 2646 3469 2652 3470
rect 2646 3465 2647 3469
rect 2651 3465 2652 3469
rect 2646 3464 2652 3465
rect 2782 3469 2788 3470
rect 2782 3465 2783 3469
rect 2787 3465 2788 3469
rect 2782 3464 2788 3465
rect 2926 3469 2932 3470
rect 2926 3465 2927 3469
rect 2931 3465 2932 3469
rect 2926 3464 2932 3465
rect 3070 3469 3076 3470
rect 3070 3465 3071 3469
rect 3075 3465 3076 3469
rect 3070 3464 3076 3465
rect 3214 3469 3220 3470
rect 3214 3465 3215 3469
rect 3219 3465 3220 3469
rect 3214 3464 3220 3465
rect 167 3459 173 3460
rect 167 3455 168 3459
rect 172 3458 173 3459
rect 242 3459 248 3460
rect 242 3458 243 3459
rect 172 3456 243 3458
rect 172 3455 173 3456
rect 167 3454 173 3455
rect 242 3455 243 3456
rect 247 3455 248 3459
rect 242 3454 248 3455
rect 295 3459 301 3460
rect 295 3455 296 3459
rect 300 3458 301 3459
rect 370 3459 376 3460
rect 370 3458 371 3459
rect 300 3456 371 3458
rect 300 3455 301 3456
rect 295 3454 301 3455
rect 370 3455 371 3456
rect 375 3455 376 3459
rect 370 3454 376 3455
rect 439 3459 445 3460
rect 439 3455 440 3459
rect 444 3458 445 3459
rect 576 3458 578 3464
rect 619 3462 621 3464
rect 650 3463 656 3464
rect 650 3462 651 3463
rect 619 3460 651 3462
rect 444 3456 578 3458
rect 583 3459 589 3460
rect 444 3455 445 3456
rect 439 3454 445 3455
rect 583 3455 584 3459
rect 588 3458 589 3459
rect 650 3459 651 3460
rect 655 3459 656 3463
rect 2535 3463 2541 3464
rect 650 3458 656 3459
rect 734 3459 741 3460
rect 588 3456 621 3458
rect 588 3455 589 3456
rect 583 3454 589 3455
rect 619 3454 621 3456
rect 682 3455 688 3456
rect 682 3454 683 3455
rect 619 3452 683 3454
rect 682 3451 683 3452
rect 687 3451 688 3455
rect 734 3455 735 3459
rect 740 3455 741 3459
rect 734 3454 741 3455
rect 887 3459 893 3460
rect 887 3455 888 3459
rect 892 3458 893 3459
rect 962 3459 968 3460
rect 962 3458 963 3459
rect 892 3456 963 3458
rect 892 3455 893 3456
rect 887 3454 893 3455
rect 962 3455 963 3456
rect 967 3455 968 3459
rect 962 3454 968 3455
rect 1023 3459 1029 3460
rect 1023 3455 1024 3459
rect 1028 3458 1029 3459
rect 1031 3459 1037 3460
rect 1031 3458 1032 3459
rect 1028 3456 1032 3458
rect 1028 3455 1029 3456
rect 1023 3454 1029 3455
rect 1031 3455 1032 3456
rect 1036 3455 1037 3459
rect 1031 3454 1037 3455
rect 1175 3459 1181 3460
rect 1175 3455 1176 3459
rect 1180 3458 1181 3459
rect 1250 3459 1256 3460
rect 1250 3458 1251 3459
rect 1180 3456 1251 3458
rect 1180 3455 1181 3456
rect 1175 3454 1181 3455
rect 1250 3455 1251 3456
rect 1255 3455 1256 3459
rect 1250 3454 1256 3455
rect 1319 3459 1325 3460
rect 1319 3455 1320 3459
rect 1324 3458 1325 3459
rect 1438 3459 1444 3460
rect 1438 3458 1439 3459
rect 1324 3456 1439 3458
rect 1324 3455 1325 3456
rect 1319 3454 1325 3455
rect 1438 3455 1439 3456
rect 1443 3455 1444 3459
rect 1438 3454 1444 3455
rect 1471 3459 1477 3460
rect 1471 3455 1472 3459
rect 1476 3458 1477 3459
rect 1538 3459 1544 3460
rect 1538 3458 1539 3459
rect 1476 3456 1539 3458
rect 1476 3455 1477 3456
rect 1471 3454 1477 3455
rect 1538 3455 1539 3456
rect 1543 3455 1544 3459
rect 2535 3459 2536 3463
rect 2540 3462 2541 3463
rect 2551 3463 2557 3464
rect 2551 3462 2552 3463
rect 2540 3460 2552 3462
rect 2540 3459 2541 3460
rect 2535 3458 2541 3459
rect 2551 3459 2552 3460
rect 2556 3459 2557 3463
rect 2551 3458 2557 3459
rect 1538 3454 1544 3455
rect 682 3450 688 3451
rect 174 3449 180 3450
rect 174 3445 175 3449
rect 179 3445 180 3449
rect 174 3444 180 3445
rect 302 3449 308 3450
rect 302 3445 303 3449
rect 307 3445 308 3449
rect 302 3444 308 3445
rect 446 3449 452 3450
rect 446 3445 447 3449
rect 451 3445 452 3449
rect 446 3444 452 3445
rect 590 3449 596 3450
rect 590 3445 591 3449
rect 595 3445 596 3449
rect 590 3444 596 3445
rect 742 3449 748 3450
rect 742 3445 743 3449
rect 747 3445 748 3449
rect 742 3444 748 3445
rect 894 3449 900 3450
rect 894 3445 895 3449
rect 899 3445 900 3449
rect 894 3444 900 3445
rect 1038 3449 1044 3450
rect 1038 3445 1039 3449
rect 1043 3445 1044 3449
rect 1038 3444 1044 3445
rect 1182 3449 1188 3450
rect 1182 3445 1183 3449
rect 1187 3445 1188 3449
rect 1182 3444 1188 3445
rect 1326 3449 1332 3450
rect 1326 3445 1327 3449
rect 1331 3445 1332 3449
rect 1326 3444 1332 3445
rect 1478 3449 1484 3450
rect 1478 3445 1479 3449
rect 1483 3445 1484 3449
rect 1478 3444 1484 3445
rect 1886 3439 1892 3440
rect 110 3436 116 3437
rect 1822 3436 1828 3437
rect 110 3432 111 3436
rect 115 3432 116 3436
rect 650 3435 656 3436
rect 650 3434 651 3435
rect 645 3432 651 3434
rect 110 3431 116 3432
rect 242 3431 248 3432
rect 242 3427 243 3431
rect 247 3430 248 3431
rect 370 3431 376 3432
rect 247 3428 321 3430
rect 247 3427 248 3428
rect 242 3426 248 3427
rect 370 3427 371 3431
rect 375 3430 376 3431
rect 650 3431 651 3432
rect 655 3431 656 3435
rect 1822 3432 1823 3436
rect 1827 3432 1828 3436
rect 1886 3435 1887 3439
rect 1891 3435 1892 3439
rect 1886 3434 1892 3435
rect 2022 3439 2028 3440
rect 2022 3435 2023 3439
rect 2027 3435 2028 3439
rect 2022 3434 2028 3435
rect 2190 3439 2196 3440
rect 2190 3435 2191 3439
rect 2195 3435 2196 3439
rect 2190 3434 2196 3435
rect 2366 3439 2372 3440
rect 2366 3435 2367 3439
rect 2371 3435 2372 3439
rect 2366 3434 2372 3435
rect 2542 3439 2548 3440
rect 2542 3435 2543 3439
rect 2547 3435 2548 3439
rect 2542 3434 2548 3435
rect 2710 3439 2716 3440
rect 2710 3435 2711 3439
rect 2715 3435 2716 3439
rect 2710 3434 2716 3435
rect 2870 3439 2876 3440
rect 2870 3435 2871 3439
rect 2875 3435 2876 3439
rect 2870 3434 2876 3435
rect 3030 3439 3036 3440
rect 3030 3435 3031 3439
rect 3035 3435 3036 3439
rect 3030 3434 3036 3435
rect 3190 3439 3196 3440
rect 3190 3435 3191 3439
rect 3195 3435 3196 3439
rect 3190 3434 3196 3435
rect 3358 3439 3364 3440
rect 3358 3435 3359 3439
rect 3363 3435 3364 3439
rect 3358 3434 3364 3435
rect 650 3430 656 3431
rect 682 3431 688 3432
rect 375 3428 465 3430
rect 375 3427 376 3428
rect 370 3426 376 3427
rect 682 3427 683 3431
rect 687 3430 688 3431
rect 823 3431 829 3432
rect 687 3428 761 3430
rect 687 3427 688 3428
rect 682 3426 688 3427
rect 823 3427 824 3431
rect 828 3430 829 3431
rect 962 3431 968 3432
rect 828 3428 913 3430
rect 828 3427 829 3428
rect 823 3426 829 3427
rect 962 3427 963 3431
rect 967 3430 968 3431
rect 1250 3431 1256 3432
rect 967 3428 1057 3430
rect 967 3427 968 3428
rect 962 3426 968 3427
rect 1250 3427 1251 3431
rect 1255 3430 1256 3431
rect 1470 3431 1476 3432
rect 1822 3431 1828 3432
rect 1990 3431 1996 3432
rect 1255 3428 1345 3430
rect 1255 3427 1256 3428
rect 1250 3426 1256 3427
rect 1470 3427 1471 3431
rect 1475 3430 1476 3431
rect 1475 3428 1497 3430
rect 1862 3429 1868 3430
rect 1475 3427 1476 3428
rect 1470 3426 1476 3427
rect 1862 3425 1863 3429
rect 1867 3425 1868 3429
rect 1990 3427 1991 3431
rect 1995 3430 1996 3431
rect 2798 3431 2804 3432
rect 2798 3430 2799 3431
rect 1995 3428 2041 3430
rect 2769 3428 2799 3430
rect 1995 3427 1996 3428
rect 1990 3426 1996 3427
rect 2798 3427 2799 3428
rect 2803 3427 2804 3431
rect 2798 3426 2804 3427
rect 3258 3431 3264 3432
rect 3258 3427 3259 3431
rect 3263 3430 3264 3431
rect 3263 3428 3377 3430
rect 3574 3429 3580 3430
rect 3263 3427 3264 3428
rect 3258 3426 3264 3427
rect 1862 3424 1868 3425
rect 3574 3425 3575 3429
rect 3579 3425 3580 3429
rect 3574 3424 3580 3425
rect 110 3419 116 3420
rect 110 3415 111 3419
rect 115 3415 116 3419
rect 110 3414 116 3415
rect 150 3419 156 3420
rect 150 3415 151 3419
rect 155 3418 156 3419
rect 1822 3419 1828 3420
rect 155 3416 185 3418
rect 155 3415 156 3416
rect 150 3414 156 3415
rect 1822 3415 1823 3419
rect 1827 3415 1828 3419
rect 1822 3414 1828 3415
rect 2015 3415 2021 3416
rect 2015 3414 2016 3415
rect 1862 3412 1868 3413
rect 1949 3412 2016 3414
rect 166 3409 172 3410
rect 166 3405 167 3409
rect 171 3405 172 3409
rect 166 3404 172 3405
rect 294 3409 300 3410
rect 294 3405 295 3409
rect 299 3405 300 3409
rect 294 3404 300 3405
rect 438 3409 444 3410
rect 438 3405 439 3409
rect 443 3405 444 3409
rect 438 3404 444 3405
rect 582 3409 588 3410
rect 582 3405 583 3409
rect 587 3405 588 3409
rect 582 3404 588 3405
rect 734 3409 740 3410
rect 734 3405 735 3409
rect 739 3405 740 3409
rect 734 3404 740 3405
rect 886 3409 892 3410
rect 886 3405 887 3409
rect 891 3405 892 3409
rect 886 3404 892 3405
rect 1030 3409 1036 3410
rect 1030 3405 1031 3409
rect 1035 3405 1036 3409
rect 1030 3404 1036 3405
rect 1174 3409 1180 3410
rect 1174 3405 1175 3409
rect 1179 3405 1180 3409
rect 1174 3404 1180 3405
rect 1318 3409 1324 3410
rect 1318 3405 1319 3409
rect 1323 3405 1324 3409
rect 1318 3404 1324 3405
rect 1470 3409 1476 3410
rect 1470 3405 1471 3409
rect 1475 3405 1476 3409
rect 1862 3408 1863 3412
rect 1867 3408 1868 3412
rect 2015 3411 2016 3412
rect 2020 3411 2021 3415
rect 2015 3410 2021 3411
rect 2090 3415 2096 3416
rect 2090 3411 2091 3415
rect 2095 3414 2096 3415
rect 2258 3415 2264 3416
rect 2095 3412 2217 3414
rect 2095 3411 2096 3412
rect 2090 3410 2096 3411
rect 2258 3411 2259 3415
rect 2263 3414 2264 3415
rect 2434 3415 2440 3416
rect 2263 3412 2393 3414
rect 2263 3411 2264 3412
rect 2258 3410 2264 3411
rect 2434 3411 2435 3415
rect 2439 3414 2440 3415
rect 3023 3415 3029 3416
rect 3023 3414 3024 3415
rect 2439 3412 2569 3414
rect 2933 3412 3024 3414
rect 2439 3411 2440 3412
rect 2434 3410 2440 3411
rect 3023 3411 3024 3412
rect 3028 3411 3029 3415
rect 3183 3415 3189 3416
rect 3183 3414 3184 3415
rect 3093 3412 3184 3414
rect 3023 3410 3029 3411
rect 3183 3411 3184 3412
rect 3188 3411 3189 3415
rect 3351 3415 3357 3416
rect 3351 3414 3352 3415
rect 3253 3412 3352 3414
rect 3183 3410 3189 3411
rect 3351 3411 3352 3412
rect 3356 3411 3357 3415
rect 3351 3410 3357 3411
rect 3574 3412 3580 3413
rect 1862 3407 1868 3408
rect 3574 3408 3575 3412
rect 3579 3408 3580 3412
rect 3574 3407 3580 3408
rect 1470 3404 1476 3405
rect 1222 3403 1229 3404
rect 1222 3399 1223 3403
rect 1228 3399 1229 3403
rect 1222 3398 1229 3399
rect 1894 3399 1900 3400
rect 1894 3395 1895 3399
rect 1899 3395 1900 3399
rect 1894 3394 1900 3395
rect 2030 3399 2036 3400
rect 2030 3395 2031 3399
rect 2035 3395 2036 3399
rect 2030 3394 2036 3395
rect 2198 3399 2204 3400
rect 2198 3395 2199 3399
rect 2203 3395 2204 3399
rect 2198 3394 2204 3395
rect 2374 3399 2380 3400
rect 2374 3395 2375 3399
rect 2379 3395 2380 3399
rect 2374 3394 2380 3395
rect 2550 3399 2556 3400
rect 2550 3395 2551 3399
rect 2555 3395 2556 3399
rect 2550 3394 2556 3395
rect 2718 3399 2724 3400
rect 2718 3395 2719 3399
rect 2723 3395 2724 3399
rect 2718 3394 2724 3395
rect 2878 3399 2884 3400
rect 2878 3395 2879 3399
rect 2883 3395 2884 3399
rect 2878 3394 2884 3395
rect 3038 3399 3044 3400
rect 3038 3395 3039 3399
rect 3043 3395 3044 3399
rect 3038 3394 3044 3395
rect 3198 3399 3204 3400
rect 3198 3395 3199 3399
rect 3203 3395 3204 3399
rect 3198 3394 3204 3395
rect 3366 3399 3372 3400
rect 3366 3395 3367 3399
rect 3371 3395 3372 3399
rect 3366 3394 3372 3395
rect 134 3387 140 3388
rect 134 3383 135 3387
rect 139 3383 140 3387
rect 134 3382 140 3383
rect 262 3387 268 3388
rect 262 3383 263 3387
rect 267 3383 268 3387
rect 262 3382 268 3383
rect 406 3387 412 3388
rect 406 3383 407 3387
rect 411 3383 412 3387
rect 406 3382 412 3383
rect 566 3387 572 3388
rect 566 3383 567 3387
rect 571 3383 572 3387
rect 566 3382 572 3383
rect 726 3387 732 3388
rect 726 3383 727 3387
rect 731 3383 732 3387
rect 726 3382 732 3383
rect 886 3387 892 3388
rect 886 3383 887 3387
rect 891 3383 892 3387
rect 886 3382 892 3383
rect 1046 3387 1052 3388
rect 1046 3383 1047 3387
rect 1051 3383 1052 3387
rect 1046 3382 1052 3383
rect 1206 3387 1212 3388
rect 1206 3383 1207 3387
rect 1211 3383 1212 3387
rect 1206 3382 1212 3383
rect 1366 3387 1372 3388
rect 1366 3383 1367 3387
rect 1371 3383 1372 3387
rect 1366 3382 1372 3383
rect 1526 3387 1532 3388
rect 1526 3383 1527 3387
rect 1531 3383 1532 3387
rect 1526 3382 1532 3383
rect 1886 3387 1893 3388
rect 1886 3383 1887 3387
rect 1892 3383 1893 3387
rect 1886 3382 1893 3383
rect 2015 3387 2021 3388
rect 2015 3383 2016 3387
rect 2020 3386 2021 3387
rect 2023 3387 2029 3388
rect 2023 3386 2024 3387
rect 2020 3384 2024 3386
rect 2020 3383 2021 3384
rect 2015 3382 2021 3383
rect 2023 3383 2024 3384
rect 2028 3383 2029 3387
rect 2023 3382 2029 3383
rect 2191 3387 2197 3388
rect 2191 3383 2192 3387
rect 2196 3386 2197 3387
rect 2258 3387 2264 3388
rect 2258 3386 2259 3387
rect 2196 3384 2259 3386
rect 2196 3383 2197 3384
rect 2191 3382 2197 3383
rect 2258 3383 2259 3384
rect 2263 3383 2264 3387
rect 2258 3382 2264 3383
rect 2367 3387 2373 3388
rect 2367 3383 2368 3387
rect 2372 3386 2373 3387
rect 2434 3387 2440 3388
rect 2434 3386 2435 3387
rect 2372 3384 2435 3386
rect 2372 3383 2373 3384
rect 2367 3382 2373 3383
rect 2434 3383 2435 3384
rect 2439 3383 2440 3387
rect 2434 3382 2440 3383
rect 2535 3387 2541 3388
rect 2535 3383 2536 3387
rect 2540 3386 2541 3387
rect 2543 3387 2549 3388
rect 2543 3386 2544 3387
rect 2540 3384 2544 3386
rect 2540 3383 2541 3384
rect 2535 3382 2541 3383
rect 2543 3383 2544 3384
rect 2548 3383 2549 3387
rect 2543 3382 2549 3383
rect 2710 3387 2717 3388
rect 2710 3383 2711 3387
rect 2716 3383 2717 3387
rect 2710 3382 2717 3383
rect 2871 3387 2877 3388
rect 2871 3383 2872 3387
rect 2876 3386 2877 3387
rect 2886 3387 2892 3388
rect 2886 3386 2887 3387
rect 2876 3384 2887 3386
rect 2876 3383 2877 3384
rect 2871 3382 2877 3383
rect 2886 3383 2887 3384
rect 2891 3383 2892 3387
rect 2886 3382 2892 3383
rect 3023 3387 3029 3388
rect 3023 3383 3024 3387
rect 3028 3386 3029 3387
rect 3031 3387 3037 3388
rect 3031 3386 3032 3387
rect 3028 3384 3032 3386
rect 3028 3383 3029 3384
rect 3023 3382 3029 3383
rect 3031 3383 3032 3384
rect 3036 3383 3037 3387
rect 3031 3382 3037 3383
rect 3183 3387 3189 3388
rect 3183 3383 3184 3387
rect 3188 3386 3189 3387
rect 3191 3387 3197 3388
rect 3191 3386 3192 3387
rect 3188 3384 3192 3386
rect 3188 3383 3189 3384
rect 3183 3382 3189 3383
rect 3191 3383 3192 3384
rect 3196 3383 3197 3387
rect 3191 3382 3197 3383
rect 3351 3387 3357 3388
rect 3351 3383 3352 3387
rect 3356 3386 3357 3387
rect 3359 3387 3365 3388
rect 3359 3386 3360 3387
rect 3356 3384 3360 3386
rect 3356 3383 3357 3384
rect 3351 3382 3357 3383
rect 3359 3383 3360 3384
rect 3364 3383 3365 3387
rect 3359 3382 3365 3383
rect 682 3379 688 3380
rect 110 3377 116 3378
rect 110 3373 111 3377
rect 115 3373 116 3377
rect 682 3375 683 3379
rect 687 3378 688 3379
rect 1023 3379 1029 3380
rect 687 3376 745 3378
rect 687 3375 688 3376
rect 682 3374 688 3375
rect 1023 3375 1024 3379
rect 1028 3378 1029 3379
rect 1028 3376 1065 3378
rect 1822 3377 1828 3378
rect 1028 3375 1029 3376
rect 1023 3374 1029 3375
rect 110 3372 116 3373
rect 1822 3373 1823 3377
rect 1827 3373 1828 3377
rect 1822 3372 1828 3373
rect 1879 3367 1885 3368
rect 255 3363 261 3364
rect 255 3362 256 3363
rect 110 3360 116 3361
rect 197 3360 256 3362
rect 110 3356 111 3360
rect 115 3356 116 3360
rect 255 3359 256 3360
rect 260 3359 261 3363
rect 399 3363 405 3364
rect 399 3362 400 3363
rect 325 3360 400 3362
rect 255 3358 261 3359
rect 399 3359 400 3360
rect 404 3359 405 3363
rect 559 3363 565 3364
rect 559 3362 560 3363
rect 469 3360 560 3362
rect 399 3358 405 3359
rect 559 3359 560 3360
rect 564 3359 565 3363
rect 719 3363 725 3364
rect 719 3362 720 3363
rect 629 3360 720 3362
rect 559 3358 565 3359
rect 719 3359 720 3360
rect 724 3359 725 3363
rect 1039 3363 1045 3364
rect 1039 3362 1040 3363
rect 949 3360 1040 3362
rect 719 3358 725 3359
rect 1039 3359 1040 3360
rect 1044 3359 1045 3363
rect 1359 3363 1365 3364
rect 1359 3362 1360 3363
rect 1269 3360 1360 3362
rect 1039 3358 1045 3359
rect 1359 3359 1360 3360
rect 1364 3359 1365 3363
rect 1511 3363 1517 3364
rect 1511 3362 1512 3363
rect 1429 3360 1512 3362
rect 1359 3358 1365 3359
rect 1511 3359 1512 3360
rect 1516 3359 1517 3363
rect 1511 3358 1517 3359
rect 1519 3363 1525 3364
rect 1519 3359 1520 3363
rect 1524 3362 1525 3363
rect 1879 3363 1880 3367
rect 1884 3366 1885 3367
rect 1887 3367 1893 3368
rect 1887 3366 1888 3367
rect 1884 3364 1888 3366
rect 1884 3363 1885 3364
rect 1879 3362 1885 3363
rect 1887 3363 1888 3364
rect 1892 3363 1893 3367
rect 1887 3362 1893 3363
rect 2023 3367 2029 3368
rect 2023 3363 2024 3367
rect 2028 3366 2029 3367
rect 2090 3367 2096 3368
rect 2090 3366 2091 3367
rect 2028 3364 2091 3366
rect 2028 3363 2029 3364
rect 2023 3362 2029 3363
rect 2090 3363 2091 3364
rect 2095 3363 2096 3367
rect 2090 3362 2096 3363
rect 2111 3367 2117 3368
rect 2111 3363 2112 3367
rect 2116 3366 2117 3367
rect 2191 3367 2197 3368
rect 2191 3366 2192 3367
rect 2116 3364 2192 3366
rect 2116 3363 2117 3364
rect 2111 3362 2117 3363
rect 2191 3363 2192 3364
rect 2196 3363 2197 3367
rect 2191 3362 2197 3363
rect 2263 3367 2269 3368
rect 2263 3363 2264 3367
rect 2268 3366 2269 3367
rect 2367 3367 2373 3368
rect 2367 3366 2368 3367
rect 2268 3364 2368 3366
rect 2268 3363 2269 3364
rect 2263 3362 2269 3363
rect 2367 3363 2368 3364
rect 2372 3363 2373 3367
rect 2367 3362 2373 3363
rect 2463 3367 2469 3368
rect 2463 3363 2464 3367
rect 2468 3366 2469 3367
rect 2543 3367 2549 3368
rect 2543 3366 2544 3367
rect 2468 3364 2544 3366
rect 2468 3363 2469 3364
rect 2463 3362 2469 3363
rect 2543 3363 2544 3364
rect 2548 3363 2549 3367
rect 2543 3362 2549 3363
rect 2711 3367 2717 3368
rect 2711 3363 2712 3367
rect 2716 3366 2717 3367
rect 2799 3367 2805 3368
rect 2799 3366 2800 3367
rect 2716 3364 2800 3366
rect 2716 3363 2717 3364
rect 2711 3362 2717 3363
rect 2799 3363 2800 3364
rect 2804 3363 2805 3367
rect 2799 3362 2805 3363
rect 2871 3367 2877 3368
rect 2871 3363 2872 3367
rect 2876 3366 2877 3367
rect 2886 3367 2892 3368
rect 2886 3366 2887 3367
rect 2876 3364 2887 3366
rect 2876 3363 2877 3364
rect 2871 3362 2877 3363
rect 2886 3363 2887 3364
rect 2891 3363 2892 3367
rect 2886 3362 2892 3363
rect 3031 3367 3037 3368
rect 3031 3363 3032 3367
rect 3036 3366 3037 3367
rect 3046 3367 3052 3368
rect 3046 3366 3047 3367
rect 3036 3364 3047 3366
rect 3036 3363 3037 3364
rect 3031 3362 3037 3363
rect 3046 3363 3047 3364
rect 3051 3363 3052 3367
rect 3046 3362 3052 3363
rect 3103 3367 3109 3368
rect 3103 3363 3104 3367
rect 3108 3366 3109 3367
rect 3183 3367 3189 3368
rect 3183 3366 3184 3367
rect 3108 3364 3184 3366
rect 3108 3363 3109 3364
rect 3103 3362 3109 3363
rect 3183 3363 3184 3364
rect 3188 3363 3189 3367
rect 3183 3362 3189 3363
rect 3263 3367 3269 3368
rect 3263 3363 3264 3367
rect 3268 3366 3269 3367
rect 3335 3367 3341 3368
rect 3335 3366 3336 3367
rect 3268 3364 3336 3366
rect 3268 3363 3269 3364
rect 3263 3362 3269 3363
rect 3335 3363 3336 3364
rect 3340 3363 3341 3367
rect 3335 3362 3341 3363
rect 3415 3367 3421 3368
rect 3415 3363 3416 3367
rect 3420 3366 3421 3367
rect 3479 3367 3485 3368
rect 3479 3366 3480 3367
rect 3420 3364 3480 3366
rect 3420 3363 3421 3364
rect 3415 3362 3421 3363
rect 3479 3363 3480 3364
rect 3484 3363 3485 3367
rect 3479 3362 3485 3363
rect 1524 3360 1553 3362
rect 1822 3360 1828 3361
rect 1524 3359 1525 3360
rect 1519 3358 1525 3359
rect 110 3355 116 3356
rect 1822 3356 1823 3360
rect 1827 3356 1828 3360
rect 1822 3355 1828 3356
rect 1894 3357 1900 3358
rect 1894 3353 1895 3357
rect 1899 3353 1900 3357
rect 1894 3352 1900 3353
rect 2030 3357 2036 3358
rect 2030 3353 2031 3357
rect 2035 3353 2036 3357
rect 2030 3352 2036 3353
rect 2198 3357 2204 3358
rect 2198 3353 2199 3357
rect 2203 3353 2204 3357
rect 2198 3352 2204 3353
rect 2374 3357 2380 3358
rect 2374 3353 2375 3357
rect 2379 3353 2380 3357
rect 2374 3352 2380 3353
rect 2550 3357 2556 3358
rect 2550 3353 2551 3357
rect 2555 3353 2556 3357
rect 2550 3352 2556 3353
rect 2718 3357 2724 3358
rect 2718 3353 2719 3357
rect 2723 3353 2724 3357
rect 2718 3352 2724 3353
rect 2878 3357 2884 3358
rect 2878 3353 2879 3357
rect 2883 3353 2884 3357
rect 2878 3352 2884 3353
rect 3038 3357 3044 3358
rect 3038 3353 3039 3357
rect 3043 3353 3044 3357
rect 3038 3352 3044 3353
rect 3190 3357 3196 3358
rect 3190 3353 3191 3357
rect 3195 3353 3196 3357
rect 3190 3352 3196 3353
rect 3342 3357 3348 3358
rect 3342 3353 3343 3357
rect 3347 3353 3348 3357
rect 3342 3352 3348 3353
rect 3486 3357 3492 3358
rect 3486 3353 3487 3357
rect 3491 3353 3492 3357
rect 3486 3352 3492 3353
rect 142 3347 148 3348
rect 142 3343 143 3347
rect 147 3343 148 3347
rect 142 3342 148 3343
rect 270 3347 276 3348
rect 270 3343 271 3347
rect 275 3343 276 3347
rect 270 3342 276 3343
rect 414 3347 420 3348
rect 414 3343 415 3347
rect 419 3343 420 3347
rect 414 3342 420 3343
rect 574 3347 580 3348
rect 574 3343 575 3347
rect 579 3343 580 3347
rect 574 3342 580 3343
rect 734 3347 740 3348
rect 734 3343 735 3347
rect 739 3343 740 3347
rect 734 3342 740 3343
rect 894 3347 900 3348
rect 894 3343 895 3347
rect 899 3343 900 3347
rect 894 3342 900 3343
rect 1054 3347 1060 3348
rect 1054 3343 1055 3347
rect 1059 3343 1060 3347
rect 1054 3342 1060 3343
rect 1214 3347 1220 3348
rect 1214 3343 1215 3347
rect 1219 3343 1220 3347
rect 1214 3342 1220 3343
rect 1374 3347 1380 3348
rect 1374 3343 1375 3347
rect 1379 3343 1380 3347
rect 1374 3342 1380 3343
rect 1534 3347 1540 3348
rect 1534 3343 1535 3347
rect 1539 3343 1540 3347
rect 1534 3342 1540 3343
rect 1862 3344 1868 3345
rect 3574 3344 3580 3345
rect 1862 3340 1863 3344
rect 1867 3340 1868 3344
rect 2111 3343 2117 3344
rect 2111 3342 2112 3343
rect 2085 3340 2112 3342
rect 1862 3339 1868 3340
rect 1886 3339 1892 3340
rect 135 3335 141 3336
rect 135 3331 136 3335
rect 140 3334 141 3335
rect 150 3335 156 3336
rect 150 3334 151 3335
rect 140 3332 151 3334
rect 140 3331 141 3332
rect 135 3330 141 3331
rect 150 3331 151 3332
rect 155 3331 156 3335
rect 150 3330 156 3331
rect 255 3335 261 3336
rect 255 3331 256 3335
rect 260 3334 261 3335
rect 263 3335 269 3336
rect 263 3334 264 3335
rect 260 3332 264 3334
rect 260 3331 261 3332
rect 255 3330 261 3331
rect 263 3331 264 3332
rect 268 3331 269 3335
rect 263 3330 269 3331
rect 399 3335 405 3336
rect 399 3331 400 3335
rect 404 3334 405 3335
rect 407 3335 413 3336
rect 407 3334 408 3335
rect 404 3332 408 3334
rect 404 3331 405 3332
rect 399 3330 405 3331
rect 407 3331 408 3332
rect 412 3331 413 3335
rect 407 3330 413 3331
rect 559 3335 565 3336
rect 559 3331 560 3335
rect 564 3334 565 3335
rect 567 3335 573 3336
rect 567 3334 568 3335
rect 564 3332 568 3334
rect 564 3331 565 3332
rect 559 3330 565 3331
rect 567 3331 568 3332
rect 572 3331 573 3335
rect 567 3330 573 3331
rect 719 3335 725 3336
rect 719 3331 720 3335
rect 724 3334 725 3335
rect 727 3335 733 3336
rect 727 3334 728 3335
rect 724 3332 728 3334
rect 724 3331 725 3332
rect 719 3330 725 3331
rect 727 3331 728 3332
rect 732 3331 733 3335
rect 727 3330 733 3331
rect 887 3335 893 3336
rect 887 3331 888 3335
rect 892 3334 893 3335
rect 895 3335 901 3336
rect 895 3334 896 3335
rect 892 3332 896 3334
rect 892 3331 893 3332
rect 887 3330 893 3331
rect 895 3331 896 3332
rect 900 3331 901 3335
rect 895 3330 901 3331
rect 1039 3335 1045 3336
rect 1039 3331 1040 3335
rect 1044 3334 1045 3335
rect 1047 3335 1053 3336
rect 1047 3334 1048 3335
rect 1044 3332 1048 3334
rect 1044 3331 1045 3332
rect 1039 3330 1045 3331
rect 1047 3331 1048 3332
rect 1052 3331 1053 3335
rect 1047 3330 1053 3331
rect 1207 3335 1213 3336
rect 1207 3331 1208 3335
rect 1212 3334 1213 3335
rect 1222 3335 1228 3336
rect 1222 3334 1223 3335
rect 1212 3332 1223 3334
rect 1212 3331 1213 3332
rect 1207 3330 1213 3331
rect 1222 3331 1223 3332
rect 1227 3331 1228 3335
rect 1222 3330 1228 3331
rect 1359 3335 1365 3336
rect 1359 3331 1360 3335
rect 1364 3334 1365 3335
rect 1367 3335 1373 3336
rect 1367 3334 1368 3335
rect 1364 3332 1368 3334
rect 1364 3331 1365 3332
rect 1359 3330 1365 3331
rect 1367 3331 1368 3332
rect 1372 3331 1373 3335
rect 1367 3330 1373 3331
rect 1511 3335 1517 3336
rect 1511 3331 1512 3335
rect 1516 3334 1517 3335
rect 1527 3335 1533 3336
rect 1527 3334 1528 3335
rect 1516 3332 1528 3334
rect 1516 3331 1517 3332
rect 1511 3330 1517 3331
rect 1527 3331 1528 3332
rect 1532 3331 1533 3335
rect 1886 3335 1887 3339
rect 1891 3338 1892 3339
rect 2111 3339 2112 3340
rect 2116 3339 2117 3343
rect 2263 3343 2269 3344
rect 2263 3342 2264 3343
rect 2253 3340 2264 3342
rect 2111 3338 2117 3339
rect 2263 3339 2264 3340
rect 2268 3339 2269 3343
rect 2463 3343 2469 3344
rect 2463 3342 2464 3343
rect 2429 3340 2464 3342
rect 2263 3338 2269 3339
rect 2463 3339 2464 3340
rect 2468 3339 2469 3343
rect 3103 3343 3109 3344
rect 3103 3342 3104 3343
rect 3093 3340 3104 3342
rect 2463 3338 2469 3339
rect 2710 3339 2716 3340
rect 1891 3336 1913 3338
rect 1891 3335 1892 3336
rect 1886 3334 1892 3335
rect 2710 3335 2711 3339
rect 2715 3338 2716 3339
rect 2799 3339 2805 3340
rect 2715 3336 2737 3338
rect 2715 3335 2716 3336
rect 2710 3334 2716 3335
rect 2799 3335 2800 3339
rect 2804 3338 2805 3339
rect 3103 3339 3104 3340
rect 3108 3339 3109 3343
rect 3263 3343 3269 3344
rect 3263 3342 3264 3343
rect 3245 3340 3264 3342
rect 3103 3338 3109 3339
rect 3263 3339 3264 3340
rect 3268 3339 3269 3343
rect 3415 3343 3421 3344
rect 3415 3342 3416 3343
rect 3397 3340 3416 3342
rect 3263 3338 3269 3339
rect 3415 3339 3416 3340
rect 3420 3339 3421 3343
rect 3574 3340 3575 3344
rect 3579 3340 3580 3344
rect 3574 3339 3580 3340
rect 3415 3338 3421 3339
rect 2804 3336 2897 3338
rect 2804 3335 2805 3336
rect 2799 3334 2805 3335
rect 1527 3330 1533 3331
rect 1862 3327 1868 3328
rect 1862 3323 1863 3327
rect 1867 3323 1868 3327
rect 1862 3322 1868 3323
rect 2478 3327 2484 3328
rect 2478 3323 2479 3327
rect 2483 3326 2484 3327
rect 3410 3327 3416 3328
rect 2483 3324 2561 3326
rect 2483 3323 2484 3324
rect 2478 3322 2484 3323
rect 3410 3323 3411 3327
rect 3415 3326 3416 3327
rect 3574 3327 3580 3328
rect 3415 3324 3497 3326
rect 3415 3323 3416 3324
rect 3410 3322 3416 3323
rect 3574 3323 3575 3327
rect 3579 3323 3580 3327
rect 3574 3322 3580 3323
rect 199 3319 205 3320
rect 199 3315 200 3319
rect 204 3318 205 3319
rect 214 3319 220 3320
rect 214 3318 215 3319
rect 204 3316 215 3318
rect 204 3315 205 3316
rect 199 3314 205 3315
rect 214 3315 215 3316
rect 219 3315 220 3319
rect 214 3314 220 3315
rect 271 3319 277 3320
rect 271 3315 272 3319
rect 276 3318 277 3319
rect 327 3319 333 3320
rect 327 3318 328 3319
rect 276 3316 328 3318
rect 276 3315 277 3316
rect 271 3314 277 3315
rect 327 3315 328 3316
rect 332 3315 333 3319
rect 327 3314 333 3315
rect 407 3319 413 3320
rect 407 3315 408 3319
rect 412 3318 413 3319
rect 471 3319 477 3320
rect 471 3318 472 3319
rect 412 3316 472 3318
rect 412 3315 413 3316
rect 407 3314 413 3315
rect 471 3315 472 3316
rect 476 3315 477 3319
rect 471 3314 477 3315
rect 551 3319 557 3320
rect 551 3315 552 3319
rect 556 3318 557 3319
rect 631 3319 637 3320
rect 631 3318 632 3319
rect 556 3316 632 3318
rect 556 3315 557 3316
rect 551 3314 557 3315
rect 631 3315 632 3316
rect 636 3315 637 3319
rect 631 3314 637 3315
rect 719 3319 725 3320
rect 719 3315 720 3319
rect 724 3318 725 3319
rect 799 3319 805 3320
rect 799 3318 800 3319
rect 724 3316 800 3318
rect 724 3315 725 3316
rect 719 3314 725 3315
rect 799 3315 800 3316
rect 804 3315 805 3319
rect 799 3314 805 3315
rect 975 3319 981 3320
rect 975 3315 976 3319
rect 980 3318 981 3319
rect 1078 3319 1084 3320
rect 1078 3318 1079 3319
rect 980 3316 1079 3318
rect 980 3315 981 3316
rect 975 3314 981 3315
rect 1078 3315 1079 3316
rect 1083 3315 1084 3319
rect 1078 3314 1084 3315
rect 1159 3319 1165 3320
rect 1159 3315 1160 3319
rect 1164 3318 1165 3319
rect 1174 3319 1180 3320
rect 1174 3318 1175 3319
rect 1164 3316 1175 3318
rect 1164 3315 1165 3316
rect 1159 3314 1165 3315
rect 1174 3315 1175 3316
rect 1179 3315 1180 3319
rect 1174 3314 1180 3315
rect 1343 3319 1349 3320
rect 1343 3315 1344 3319
rect 1348 3318 1349 3319
rect 1426 3319 1432 3320
rect 1426 3318 1427 3319
rect 1348 3316 1427 3318
rect 1348 3315 1349 3316
rect 1343 3314 1349 3315
rect 1426 3315 1427 3316
rect 1431 3315 1432 3319
rect 1426 3314 1432 3315
rect 1519 3319 1525 3320
rect 1519 3315 1520 3319
rect 1524 3318 1525 3319
rect 1535 3319 1541 3320
rect 1535 3318 1536 3319
rect 1524 3316 1536 3318
rect 1524 3315 1525 3316
rect 1519 3314 1525 3315
rect 1535 3315 1536 3316
rect 1540 3315 1541 3319
rect 1535 3314 1541 3315
rect 1886 3317 1892 3318
rect 1886 3313 1887 3317
rect 1891 3313 1892 3317
rect 1886 3312 1892 3313
rect 2022 3317 2028 3318
rect 2022 3313 2023 3317
rect 2027 3313 2028 3317
rect 2022 3312 2028 3313
rect 2190 3317 2196 3318
rect 2190 3313 2191 3317
rect 2195 3313 2196 3317
rect 2190 3312 2196 3313
rect 2366 3317 2372 3318
rect 2366 3313 2367 3317
rect 2371 3313 2372 3317
rect 2366 3312 2372 3313
rect 2542 3317 2548 3318
rect 2542 3313 2543 3317
rect 2547 3313 2548 3317
rect 2542 3312 2548 3313
rect 2710 3317 2716 3318
rect 2710 3313 2711 3317
rect 2715 3313 2716 3317
rect 2710 3312 2716 3313
rect 2870 3317 2876 3318
rect 2870 3313 2871 3317
rect 2875 3313 2876 3317
rect 2870 3312 2876 3313
rect 3030 3317 3036 3318
rect 3030 3313 3031 3317
rect 3035 3313 3036 3317
rect 3030 3312 3036 3313
rect 3182 3317 3188 3318
rect 3182 3313 3183 3317
rect 3187 3313 3188 3317
rect 3182 3312 3188 3313
rect 3334 3317 3340 3318
rect 3334 3313 3335 3317
rect 3339 3313 3340 3317
rect 3334 3312 3340 3313
rect 3478 3317 3484 3318
rect 3478 3313 3479 3317
rect 3483 3313 3484 3317
rect 3478 3312 3484 3313
rect 206 3309 212 3310
rect 206 3305 207 3309
rect 211 3305 212 3309
rect 206 3304 212 3305
rect 334 3309 340 3310
rect 334 3305 335 3309
rect 339 3305 340 3309
rect 334 3304 340 3305
rect 478 3309 484 3310
rect 478 3305 479 3309
rect 483 3305 484 3309
rect 478 3304 484 3305
rect 638 3309 644 3310
rect 638 3305 639 3309
rect 643 3305 644 3309
rect 638 3304 644 3305
rect 806 3309 812 3310
rect 806 3305 807 3309
rect 811 3305 812 3309
rect 806 3304 812 3305
rect 982 3309 988 3310
rect 982 3305 983 3309
rect 987 3305 988 3309
rect 982 3304 988 3305
rect 1166 3309 1172 3310
rect 1166 3305 1167 3309
rect 1171 3305 1172 3309
rect 1166 3304 1172 3305
rect 1350 3309 1356 3310
rect 1350 3305 1351 3309
rect 1355 3305 1356 3309
rect 1350 3304 1356 3305
rect 1542 3309 1548 3310
rect 1542 3305 1543 3309
rect 1547 3305 1548 3309
rect 1542 3304 1548 3305
rect 110 3296 116 3297
rect 1822 3296 1828 3297
rect 110 3292 111 3296
rect 115 3292 116 3296
rect 271 3295 277 3296
rect 271 3294 272 3295
rect 261 3292 272 3294
rect 110 3291 116 3292
rect 271 3291 272 3292
rect 276 3291 277 3295
rect 407 3295 413 3296
rect 407 3294 408 3295
rect 389 3292 408 3294
rect 271 3290 277 3291
rect 407 3291 408 3292
rect 412 3291 413 3295
rect 551 3295 557 3296
rect 551 3294 552 3295
rect 533 3292 552 3294
rect 407 3290 413 3291
rect 551 3291 552 3292
rect 556 3291 557 3295
rect 719 3295 725 3296
rect 719 3294 720 3295
rect 693 3292 720 3294
rect 551 3290 557 3291
rect 719 3291 720 3292
rect 724 3291 725 3295
rect 1822 3292 1823 3296
rect 1827 3292 1828 3296
rect 719 3290 725 3291
rect 895 3291 901 3292
rect 895 3287 896 3291
rect 900 3290 901 3291
rect 1078 3291 1084 3292
rect 900 3288 1001 3290
rect 900 3287 901 3288
rect 895 3286 901 3287
rect 1078 3287 1079 3291
rect 1083 3290 1084 3291
rect 1426 3291 1432 3292
rect 1822 3291 1828 3292
rect 1886 3295 1892 3296
rect 1886 3291 1887 3295
rect 1891 3291 1892 3295
rect 1083 3288 1185 3290
rect 1083 3287 1084 3288
rect 1078 3286 1084 3287
rect 1426 3287 1427 3291
rect 1431 3290 1432 3291
rect 1886 3290 1892 3291
rect 2006 3295 2012 3296
rect 2006 3291 2007 3295
rect 2011 3291 2012 3295
rect 2006 3290 2012 3291
rect 2150 3295 2156 3296
rect 2150 3291 2151 3295
rect 2155 3291 2156 3295
rect 2150 3290 2156 3291
rect 2302 3295 2308 3296
rect 2302 3291 2303 3295
rect 2307 3291 2308 3295
rect 2302 3290 2308 3291
rect 2462 3295 2468 3296
rect 2462 3291 2463 3295
rect 2467 3291 2468 3295
rect 2462 3290 2468 3291
rect 2630 3295 2636 3296
rect 2630 3291 2631 3295
rect 2635 3291 2636 3295
rect 2630 3290 2636 3291
rect 2798 3295 2804 3296
rect 2798 3291 2799 3295
rect 2803 3291 2804 3295
rect 2798 3290 2804 3291
rect 2966 3295 2972 3296
rect 2966 3291 2967 3295
rect 2971 3291 2972 3295
rect 2966 3290 2972 3291
rect 3134 3295 3140 3296
rect 3134 3291 3135 3295
rect 3139 3291 3140 3295
rect 3134 3290 3140 3291
rect 3310 3295 3316 3296
rect 3310 3291 3311 3295
rect 3315 3291 3316 3295
rect 3310 3290 3316 3291
rect 3478 3295 3484 3296
rect 3478 3291 3479 3295
rect 3483 3291 3484 3295
rect 3478 3290 3484 3291
rect 1431 3288 1561 3290
rect 1431 3287 1432 3288
rect 1426 3286 1432 3287
rect 1879 3287 1885 3288
rect 1862 3285 1868 3286
rect 1862 3281 1863 3285
rect 1867 3281 1868 3285
rect 1879 3283 1880 3287
rect 1884 3286 1885 3287
rect 2538 3287 2544 3288
rect 1884 3284 1905 3286
rect 1884 3283 1885 3284
rect 1879 3282 1885 3283
rect 2538 3283 2539 3287
rect 2543 3286 2544 3287
rect 2886 3287 2892 3288
rect 2886 3286 2887 3287
rect 2543 3284 2649 3286
rect 2857 3284 2887 3286
rect 2543 3283 2544 3284
rect 2538 3282 2544 3283
rect 2886 3283 2887 3284
rect 2891 3283 2892 3287
rect 3480 3284 3497 3286
rect 3574 3285 3580 3286
rect 2886 3282 2892 3283
rect 3478 3283 3484 3284
rect 1862 3280 1868 3281
rect 110 3279 116 3280
rect 110 3275 111 3279
rect 115 3275 116 3279
rect 1822 3279 1828 3280
rect 110 3274 116 3275
rect 744 3276 817 3278
rect 198 3269 204 3270
rect 198 3265 199 3269
rect 203 3265 204 3269
rect 198 3264 204 3265
rect 326 3269 332 3270
rect 326 3265 327 3269
rect 331 3265 332 3269
rect 326 3264 332 3265
rect 470 3269 476 3270
rect 470 3265 471 3269
rect 475 3265 476 3269
rect 470 3264 476 3265
rect 630 3269 636 3270
rect 630 3265 631 3269
rect 635 3265 636 3269
rect 630 3264 636 3265
rect 487 3263 493 3264
rect 487 3259 488 3263
rect 492 3262 493 3263
rect 744 3262 746 3276
rect 1822 3275 1823 3279
rect 1827 3275 1828 3279
rect 3478 3279 3479 3283
rect 3483 3279 3484 3283
rect 3574 3281 3575 3285
rect 3579 3281 3580 3285
rect 3574 3280 3580 3281
rect 3478 3278 3484 3279
rect 1822 3274 1828 3275
rect 1954 3271 1960 3272
rect 798 3269 804 3270
rect 798 3265 799 3269
rect 803 3265 804 3269
rect 798 3264 804 3265
rect 974 3269 980 3270
rect 974 3265 975 3269
rect 979 3265 980 3269
rect 974 3264 980 3265
rect 1158 3269 1164 3270
rect 1158 3265 1159 3269
rect 1163 3265 1164 3269
rect 1158 3264 1164 3265
rect 1342 3269 1348 3270
rect 1342 3265 1343 3269
rect 1347 3265 1348 3269
rect 1342 3264 1348 3265
rect 1534 3269 1540 3270
rect 1534 3265 1535 3269
rect 1539 3265 1540 3269
rect 1534 3264 1540 3265
rect 1862 3268 1868 3269
rect 1862 3264 1863 3268
rect 1867 3264 1868 3268
rect 1954 3267 1955 3271
rect 1959 3270 1960 3271
rect 2234 3271 2240 3272
rect 2234 3270 2235 3271
rect 1959 3268 2033 3270
rect 2213 3268 2235 3270
rect 1959 3267 1960 3268
rect 1954 3266 1960 3267
rect 2234 3267 2235 3268
rect 2239 3267 2240 3271
rect 2455 3271 2461 3272
rect 2455 3270 2456 3271
rect 2365 3268 2456 3270
rect 2234 3266 2240 3267
rect 2455 3267 2456 3268
rect 2460 3267 2461 3271
rect 2623 3271 2629 3272
rect 2623 3270 2624 3271
rect 2525 3268 2624 3270
rect 2455 3266 2461 3267
rect 2623 3267 2624 3268
rect 2628 3267 2629 3271
rect 2623 3266 2629 3267
rect 2866 3271 2872 3272
rect 2866 3267 2867 3271
rect 2871 3270 2872 3271
rect 3054 3271 3060 3272
rect 2871 3268 2993 3270
rect 2871 3267 2872 3268
rect 2866 3266 2872 3267
rect 3054 3267 3055 3271
rect 3059 3270 3060 3271
rect 3471 3271 3477 3272
rect 3471 3270 3472 3271
rect 3059 3268 3161 3270
rect 3373 3268 3472 3270
rect 3059 3267 3060 3268
rect 3054 3266 3060 3267
rect 3471 3267 3472 3268
rect 3476 3267 3477 3271
rect 3471 3266 3477 3267
rect 3574 3268 3580 3269
rect 492 3260 746 3262
rect 1391 3263 1397 3264
rect 492 3259 493 3260
rect 487 3258 493 3259
rect 1391 3259 1392 3263
rect 1396 3262 1397 3263
rect 1407 3263 1413 3264
rect 1862 3263 1868 3264
rect 3574 3264 3575 3268
rect 3579 3264 3580 3268
rect 3574 3263 3580 3264
rect 1407 3262 1408 3263
rect 1396 3260 1408 3262
rect 1396 3259 1397 3260
rect 1391 3258 1397 3259
rect 1407 3259 1408 3260
rect 1412 3259 1413 3263
rect 1407 3258 1413 3259
rect 1894 3255 1900 3256
rect 1894 3251 1895 3255
rect 1899 3251 1900 3255
rect 1894 3250 1900 3251
rect 2014 3255 2020 3256
rect 2014 3251 2015 3255
rect 2019 3251 2020 3255
rect 2014 3250 2020 3251
rect 2158 3255 2164 3256
rect 2158 3251 2159 3255
rect 2163 3251 2164 3255
rect 2158 3250 2164 3251
rect 2310 3255 2316 3256
rect 2310 3251 2311 3255
rect 2315 3251 2316 3255
rect 2310 3250 2316 3251
rect 2470 3255 2476 3256
rect 2470 3251 2471 3255
rect 2475 3251 2476 3255
rect 2470 3250 2476 3251
rect 2638 3255 2644 3256
rect 2638 3251 2639 3255
rect 2643 3251 2644 3255
rect 2638 3250 2644 3251
rect 2806 3255 2812 3256
rect 2806 3251 2807 3255
rect 2811 3251 2812 3255
rect 2806 3250 2812 3251
rect 2974 3255 2980 3256
rect 2974 3251 2975 3255
rect 2979 3251 2980 3255
rect 2974 3250 2980 3251
rect 3142 3255 3148 3256
rect 3142 3251 3143 3255
rect 3147 3251 3148 3255
rect 3142 3250 3148 3251
rect 3318 3255 3324 3256
rect 3318 3251 3319 3255
rect 3323 3251 3324 3255
rect 3318 3250 3324 3251
rect 3486 3255 3492 3256
rect 3486 3251 3487 3255
rect 3491 3251 3492 3255
rect 3486 3250 3492 3251
rect 366 3243 372 3244
rect 366 3239 367 3243
rect 371 3239 372 3243
rect 366 3238 372 3239
rect 502 3243 508 3244
rect 502 3239 503 3243
rect 507 3239 508 3243
rect 502 3238 508 3239
rect 638 3243 644 3244
rect 638 3239 639 3243
rect 643 3239 644 3243
rect 638 3238 644 3239
rect 782 3243 788 3244
rect 782 3239 783 3243
rect 787 3239 788 3243
rect 782 3238 788 3239
rect 934 3243 940 3244
rect 934 3239 935 3243
rect 939 3239 940 3243
rect 934 3238 940 3239
rect 1094 3243 1100 3244
rect 1094 3239 1095 3243
rect 1099 3239 1100 3243
rect 1094 3238 1100 3239
rect 1254 3243 1260 3244
rect 1254 3239 1255 3243
rect 1259 3239 1260 3243
rect 1254 3238 1260 3239
rect 1414 3243 1420 3244
rect 1414 3239 1415 3243
rect 1419 3239 1420 3243
rect 1414 3238 1420 3239
rect 1574 3243 1580 3244
rect 1574 3239 1575 3243
rect 1579 3239 1580 3243
rect 1574 3238 1580 3239
rect 1887 3243 1893 3244
rect 1887 3239 1888 3243
rect 1892 3242 1893 3243
rect 1950 3243 1956 3244
rect 1950 3242 1951 3243
rect 1892 3240 1951 3242
rect 1892 3239 1893 3240
rect 1887 3238 1893 3239
rect 1950 3239 1951 3240
rect 1955 3239 1956 3243
rect 1950 3238 1956 3239
rect 1958 3243 1964 3244
rect 1958 3239 1959 3243
rect 1963 3242 1964 3243
rect 2007 3243 2013 3244
rect 2007 3242 2008 3243
rect 1963 3240 2008 3242
rect 1963 3239 1964 3240
rect 1958 3238 1964 3239
rect 2007 3239 2008 3240
rect 2012 3239 2013 3243
rect 2007 3238 2013 3239
rect 2151 3243 2157 3244
rect 2151 3239 2152 3243
rect 2156 3242 2157 3243
rect 2166 3243 2172 3244
rect 2166 3242 2167 3243
rect 2156 3240 2167 3242
rect 2156 3239 2157 3240
rect 2151 3238 2157 3239
rect 2166 3239 2167 3240
rect 2171 3239 2172 3243
rect 2166 3238 2172 3239
rect 2234 3243 2240 3244
rect 2234 3239 2235 3243
rect 2239 3242 2240 3243
rect 2303 3243 2309 3244
rect 2303 3242 2304 3243
rect 2239 3240 2304 3242
rect 2239 3239 2240 3240
rect 2234 3238 2240 3239
rect 2303 3239 2304 3240
rect 2308 3239 2309 3243
rect 2303 3238 2309 3239
rect 2455 3243 2461 3244
rect 2455 3239 2456 3243
rect 2460 3242 2461 3243
rect 2463 3243 2469 3244
rect 2463 3242 2464 3243
rect 2460 3240 2464 3242
rect 2460 3239 2461 3240
rect 2455 3238 2461 3239
rect 2463 3239 2464 3240
rect 2468 3239 2469 3243
rect 2463 3238 2469 3239
rect 2623 3243 2629 3244
rect 2623 3239 2624 3243
rect 2628 3242 2629 3243
rect 2631 3243 2637 3244
rect 2631 3242 2632 3243
rect 2628 3240 2632 3242
rect 2628 3239 2629 3240
rect 2623 3238 2629 3239
rect 2631 3239 2632 3240
rect 2636 3239 2637 3243
rect 2631 3238 2637 3239
rect 2799 3243 2805 3244
rect 2799 3239 2800 3243
rect 2804 3242 2805 3243
rect 2866 3243 2872 3244
rect 2866 3242 2867 3243
rect 2804 3240 2867 3242
rect 2804 3239 2805 3240
rect 2799 3238 2805 3239
rect 2866 3239 2867 3240
rect 2871 3239 2872 3243
rect 2866 3238 2872 3239
rect 2967 3243 2973 3244
rect 2967 3239 2968 3243
rect 2972 3242 2973 3243
rect 3054 3243 3060 3244
rect 3054 3242 3055 3243
rect 2972 3240 3055 3242
rect 2972 3239 2973 3240
rect 2967 3238 2973 3239
rect 3054 3239 3055 3240
rect 3059 3239 3060 3243
rect 3054 3238 3060 3239
rect 3135 3243 3141 3244
rect 3135 3239 3136 3243
rect 3140 3242 3141 3243
rect 3258 3243 3264 3244
rect 3258 3242 3259 3243
rect 3140 3240 3259 3242
rect 3140 3239 3141 3240
rect 3135 3238 3141 3239
rect 3258 3239 3259 3240
rect 3263 3239 3264 3243
rect 3258 3238 3264 3239
rect 3311 3243 3317 3244
rect 3311 3239 3312 3243
rect 3316 3242 3317 3243
rect 3410 3243 3416 3244
rect 3410 3242 3411 3243
rect 3316 3240 3411 3242
rect 3316 3239 3317 3240
rect 3311 3238 3317 3239
rect 3410 3239 3411 3240
rect 3415 3239 3416 3243
rect 3410 3238 3416 3239
rect 3471 3243 3477 3244
rect 3471 3239 3472 3243
rect 3476 3242 3477 3243
rect 3479 3243 3485 3244
rect 3479 3242 3480 3243
rect 3476 3240 3480 3242
rect 3476 3239 3477 3240
rect 3471 3238 3477 3239
rect 3479 3239 3480 3240
rect 3484 3239 3485 3243
rect 3479 3238 3485 3239
rect 710 3235 716 3236
rect 110 3233 116 3234
rect 110 3229 111 3233
rect 115 3229 116 3233
rect 710 3231 711 3235
rect 715 3234 716 3235
rect 1174 3235 1180 3236
rect 1174 3234 1175 3235
rect 715 3232 801 3234
rect 1153 3232 1175 3234
rect 715 3231 716 3232
rect 710 3230 716 3231
rect 1174 3231 1175 3232
rect 1179 3231 1180 3235
rect 1174 3230 1180 3231
rect 1822 3233 1828 3234
rect 110 3228 116 3229
rect 1822 3229 1823 3233
rect 1827 3229 1828 3233
rect 1822 3228 1828 3229
rect 1887 3223 1893 3224
rect 495 3219 501 3220
rect 495 3218 496 3219
rect 110 3216 116 3217
rect 429 3216 496 3218
rect 110 3212 111 3216
rect 115 3212 116 3216
rect 495 3215 496 3216
rect 500 3215 501 3219
rect 631 3219 637 3220
rect 631 3218 632 3219
rect 565 3216 632 3218
rect 495 3214 501 3215
rect 631 3215 632 3216
rect 636 3215 637 3219
rect 775 3219 781 3220
rect 775 3218 776 3219
rect 701 3216 776 3218
rect 631 3214 637 3215
rect 775 3215 776 3216
rect 780 3215 781 3219
rect 1087 3219 1093 3220
rect 1087 3218 1088 3219
rect 997 3216 1088 3218
rect 775 3214 781 3215
rect 1087 3215 1088 3216
rect 1092 3215 1093 3219
rect 1087 3214 1093 3215
rect 1162 3219 1168 3220
rect 1162 3215 1163 3219
rect 1167 3218 1168 3219
rect 1567 3219 1573 3220
rect 1567 3218 1568 3219
rect 1167 3216 1281 3218
rect 1477 3216 1568 3218
rect 1167 3215 1168 3216
rect 1162 3214 1168 3215
rect 1567 3215 1568 3216
rect 1572 3215 1573 3219
rect 1646 3219 1652 3220
rect 1646 3218 1647 3219
rect 1637 3216 1647 3218
rect 1567 3214 1573 3215
rect 1646 3215 1647 3216
rect 1651 3215 1652 3219
rect 1887 3219 1888 3223
rect 1892 3222 1893 3223
rect 1966 3223 1972 3224
rect 1966 3222 1967 3223
rect 1892 3220 1967 3222
rect 1892 3219 1893 3220
rect 1887 3218 1893 3219
rect 1966 3219 1967 3220
rect 1971 3219 1972 3223
rect 1966 3218 1972 3219
rect 2015 3223 2021 3224
rect 2015 3219 2016 3223
rect 2020 3222 2021 3223
rect 2030 3223 2036 3224
rect 2030 3222 2031 3223
rect 2020 3220 2031 3222
rect 2020 3219 2021 3220
rect 2015 3218 2021 3219
rect 2030 3219 2031 3220
rect 2035 3219 2036 3223
rect 2030 3218 2036 3219
rect 2167 3223 2173 3224
rect 2167 3219 2168 3223
rect 2172 3222 2173 3223
rect 2182 3223 2188 3224
rect 2182 3222 2183 3223
rect 2172 3220 2183 3222
rect 2172 3219 2173 3220
rect 2167 3218 2173 3219
rect 2182 3219 2183 3220
rect 2187 3219 2188 3223
rect 2182 3218 2188 3219
rect 2242 3223 2248 3224
rect 2242 3219 2243 3223
rect 2247 3222 2248 3223
rect 2319 3223 2325 3224
rect 2319 3222 2320 3223
rect 2247 3220 2320 3222
rect 2247 3219 2248 3220
rect 2242 3218 2248 3219
rect 2319 3219 2320 3220
rect 2324 3219 2325 3223
rect 2319 3218 2325 3219
rect 2398 3223 2404 3224
rect 2398 3219 2399 3223
rect 2403 3222 2404 3223
rect 2455 3223 2461 3224
rect 2455 3222 2456 3223
rect 2403 3220 2456 3222
rect 2403 3219 2404 3220
rect 2398 3218 2404 3219
rect 2455 3219 2456 3220
rect 2460 3219 2461 3223
rect 2455 3218 2461 3219
rect 2526 3223 2532 3224
rect 2526 3219 2527 3223
rect 2531 3222 2532 3223
rect 2591 3223 2597 3224
rect 2591 3222 2592 3223
rect 2531 3220 2592 3222
rect 2531 3219 2532 3220
rect 2526 3218 2532 3219
rect 2591 3219 2592 3220
rect 2596 3219 2597 3223
rect 2591 3218 2597 3219
rect 2727 3223 2733 3224
rect 2727 3219 2728 3223
rect 2732 3222 2733 3223
rect 2790 3223 2796 3224
rect 2790 3222 2791 3223
rect 2732 3220 2791 3222
rect 2732 3219 2733 3220
rect 2727 3218 2733 3219
rect 2790 3219 2791 3220
rect 2795 3219 2796 3223
rect 2790 3218 2796 3219
rect 2807 3223 2813 3224
rect 2807 3219 2808 3223
rect 2812 3222 2813 3223
rect 2863 3223 2869 3224
rect 2863 3222 2864 3223
rect 2812 3220 2864 3222
rect 2812 3219 2813 3220
rect 2807 3218 2813 3219
rect 2863 3219 2864 3220
rect 2868 3219 2869 3223
rect 2863 3218 2869 3219
rect 2942 3223 2948 3224
rect 2942 3219 2943 3223
rect 2947 3222 2948 3223
rect 3007 3223 3013 3224
rect 3007 3222 3008 3223
rect 2947 3220 3008 3222
rect 2947 3219 2948 3220
rect 2942 3218 2948 3219
rect 3007 3219 3008 3220
rect 3012 3219 3013 3223
rect 3007 3218 3013 3219
rect 3082 3223 3088 3224
rect 3082 3219 3083 3223
rect 3087 3222 3088 3223
rect 3159 3223 3165 3224
rect 3159 3222 3160 3223
rect 3087 3220 3160 3222
rect 3087 3219 3088 3220
rect 3082 3218 3088 3219
rect 3159 3219 3160 3220
rect 3164 3219 3165 3223
rect 3159 3218 3165 3219
rect 3250 3223 3256 3224
rect 3250 3219 3251 3223
rect 3255 3222 3256 3223
rect 3319 3223 3325 3224
rect 3319 3222 3320 3223
rect 3255 3220 3320 3222
rect 3255 3219 3256 3220
rect 3250 3218 3256 3219
rect 3319 3219 3320 3220
rect 3324 3219 3325 3223
rect 3319 3218 3325 3219
rect 3478 3223 3485 3224
rect 3478 3219 3479 3223
rect 3484 3219 3485 3223
rect 3478 3218 3485 3219
rect 1646 3214 1652 3215
rect 1822 3216 1828 3217
rect 110 3211 116 3212
rect 1822 3212 1823 3216
rect 1827 3212 1828 3216
rect 1822 3211 1828 3212
rect 1894 3213 1900 3214
rect 1894 3209 1895 3213
rect 1899 3209 1900 3213
rect 1894 3208 1900 3209
rect 2022 3213 2028 3214
rect 2022 3209 2023 3213
rect 2027 3209 2028 3213
rect 2022 3208 2028 3209
rect 2174 3213 2180 3214
rect 2174 3209 2175 3213
rect 2179 3209 2180 3213
rect 2174 3208 2180 3209
rect 2326 3213 2332 3214
rect 2326 3209 2327 3213
rect 2331 3209 2332 3213
rect 2326 3208 2332 3209
rect 2462 3213 2468 3214
rect 2462 3209 2463 3213
rect 2467 3209 2468 3213
rect 2462 3208 2468 3209
rect 2598 3213 2604 3214
rect 2598 3209 2599 3213
rect 2603 3209 2604 3213
rect 2598 3208 2604 3209
rect 2734 3213 2740 3214
rect 2734 3209 2735 3213
rect 2739 3209 2740 3213
rect 2734 3208 2740 3209
rect 2870 3213 2876 3214
rect 2870 3209 2871 3213
rect 2875 3209 2876 3213
rect 2870 3208 2876 3209
rect 3014 3213 3020 3214
rect 3014 3209 3015 3213
rect 3019 3209 3020 3213
rect 3014 3208 3020 3209
rect 3166 3213 3172 3214
rect 3166 3209 3167 3213
rect 3171 3209 3172 3213
rect 3166 3208 3172 3209
rect 3326 3213 3332 3214
rect 3326 3209 3327 3213
rect 3331 3209 3332 3213
rect 3326 3208 3332 3209
rect 3486 3213 3492 3214
rect 3486 3209 3487 3213
rect 3491 3209 3492 3213
rect 3486 3208 3492 3209
rect 374 3203 380 3204
rect 374 3199 375 3203
rect 379 3199 380 3203
rect 374 3198 380 3199
rect 510 3203 516 3204
rect 510 3199 511 3203
rect 515 3199 516 3203
rect 510 3198 516 3199
rect 646 3203 652 3204
rect 646 3199 647 3203
rect 651 3199 652 3203
rect 646 3198 652 3199
rect 790 3203 796 3204
rect 790 3199 791 3203
rect 795 3199 796 3203
rect 790 3198 796 3199
rect 942 3203 948 3204
rect 942 3199 943 3203
rect 947 3199 948 3203
rect 942 3198 948 3199
rect 1102 3203 1108 3204
rect 1102 3199 1103 3203
rect 1107 3199 1108 3203
rect 1102 3198 1108 3199
rect 1262 3203 1268 3204
rect 1262 3199 1263 3203
rect 1267 3199 1268 3203
rect 1262 3198 1268 3199
rect 1422 3203 1428 3204
rect 1422 3199 1423 3203
rect 1427 3199 1428 3203
rect 1422 3198 1428 3199
rect 1582 3203 1588 3204
rect 1582 3199 1583 3203
rect 1587 3199 1588 3203
rect 1582 3198 1588 3199
rect 1862 3200 1868 3201
rect 3574 3200 3580 3201
rect 1862 3196 1863 3200
rect 1867 3196 1868 3200
rect 1958 3199 1964 3200
rect 1958 3198 1959 3199
rect 1949 3196 1959 3198
rect 1862 3195 1868 3196
rect 1958 3195 1959 3196
rect 1963 3195 1964 3199
rect 2242 3199 2248 3200
rect 2242 3198 2243 3199
rect 2229 3196 2243 3198
rect 1958 3194 1964 3195
rect 1966 3195 1972 3196
rect 367 3191 373 3192
rect 367 3187 368 3191
rect 372 3190 373 3191
rect 487 3191 493 3192
rect 487 3190 488 3191
rect 372 3188 488 3190
rect 372 3187 373 3188
rect 367 3186 373 3187
rect 487 3187 488 3188
rect 492 3187 493 3191
rect 487 3186 493 3187
rect 495 3191 501 3192
rect 495 3187 496 3191
rect 500 3190 501 3191
rect 503 3191 509 3192
rect 503 3190 504 3191
rect 500 3188 504 3190
rect 500 3187 501 3188
rect 495 3186 501 3187
rect 503 3187 504 3188
rect 508 3187 509 3191
rect 503 3186 509 3187
rect 631 3191 637 3192
rect 631 3187 632 3191
rect 636 3190 637 3191
rect 639 3191 645 3192
rect 639 3190 640 3191
rect 636 3188 640 3190
rect 636 3187 637 3188
rect 631 3186 637 3187
rect 639 3187 640 3188
rect 644 3187 645 3191
rect 639 3186 645 3187
rect 775 3191 781 3192
rect 775 3187 776 3191
rect 780 3190 781 3191
rect 783 3191 789 3192
rect 783 3190 784 3191
rect 780 3188 784 3190
rect 780 3187 781 3188
rect 775 3186 781 3187
rect 783 3187 784 3188
rect 788 3187 789 3191
rect 783 3186 789 3187
rect 935 3191 941 3192
rect 935 3187 936 3191
rect 940 3190 941 3191
rect 950 3191 956 3192
rect 950 3190 951 3191
rect 940 3188 951 3190
rect 940 3187 941 3188
rect 935 3186 941 3187
rect 950 3187 951 3188
rect 955 3187 956 3191
rect 950 3186 956 3187
rect 1087 3191 1093 3192
rect 1087 3187 1088 3191
rect 1092 3190 1093 3191
rect 1095 3191 1101 3192
rect 1095 3190 1096 3191
rect 1092 3188 1096 3190
rect 1092 3187 1093 3188
rect 1087 3186 1093 3187
rect 1095 3187 1096 3188
rect 1100 3187 1101 3191
rect 1095 3186 1101 3187
rect 1199 3191 1205 3192
rect 1199 3187 1200 3191
rect 1204 3190 1205 3191
rect 1255 3191 1261 3192
rect 1255 3190 1256 3191
rect 1204 3188 1256 3190
rect 1204 3187 1205 3188
rect 1199 3186 1205 3187
rect 1255 3187 1256 3188
rect 1260 3187 1261 3191
rect 1255 3186 1261 3187
rect 1407 3191 1413 3192
rect 1407 3187 1408 3191
rect 1412 3190 1413 3191
rect 1415 3191 1421 3192
rect 1415 3190 1416 3191
rect 1412 3188 1416 3190
rect 1412 3187 1413 3188
rect 1407 3186 1413 3187
rect 1415 3187 1416 3188
rect 1420 3187 1421 3191
rect 1415 3186 1421 3187
rect 1567 3191 1573 3192
rect 1567 3187 1568 3191
rect 1572 3190 1573 3191
rect 1575 3191 1581 3192
rect 1575 3190 1576 3191
rect 1572 3188 1576 3190
rect 1572 3187 1573 3188
rect 1567 3186 1573 3187
rect 1575 3187 1576 3188
rect 1580 3187 1581 3191
rect 1966 3191 1967 3195
rect 1971 3194 1972 3195
rect 2242 3195 2243 3196
rect 2247 3195 2248 3199
rect 2398 3199 2404 3200
rect 2398 3198 2399 3199
rect 2381 3196 2399 3198
rect 2242 3194 2248 3195
rect 2398 3195 2399 3196
rect 2403 3195 2404 3199
rect 2526 3199 2532 3200
rect 2526 3198 2527 3199
rect 2517 3196 2527 3198
rect 2398 3194 2404 3195
rect 2526 3195 2527 3196
rect 2531 3195 2532 3199
rect 2807 3199 2813 3200
rect 2807 3198 2808 3199
rect 2789 3196 2808 3198
rect 2526 3194 2532 3195
rect 2807 3195 2808 3196
rect 2812 3195 2813 3199
rect 2942 3199 2948 3200
rect 2942 3198 2943 3199
rect 2925 3196 2943 3198
rect 2807 3194 2813 3195
rect 2942 3195 2943 3196
rect 2947 3195 2948 3199
rect 3082 3199 3088 3200
rect 3082 3198 3083 3199
rect 3069 3196 3083 3198
rect 2942 3194 2948 3195
rect 3082 3195 3083 3196
rect 3087 3195 3088 3199
rect 3250 3199 3256 3200
rect 3250 3198 3251 3199
rect 3221 3196 3251 3198
rect 3082 3194 3088 3195
rect 3250 3195 3251 3196
rect 3255 3195 3256 3199
rect 3574 3196 3575 3200
rect 3579 3196 3580 3200
rect 3250 3194 3256 3195
rect 3258 3195 3264 3196
rect 3574 3195 3580 3196
rect 1971 3192 2041 3194
rect 1971 3191 1972 3192
rect 1966 3190 1972 3191
rect 3258 3191 3259 3195
rect 3263 3194 3264 3195
rect 3263 3192 3345 3194
rect 3263 3191 3264 3192
rect 3258 3190 3264 3191
rect 1575 3186 1581 3187
rect 1862 3183 1868 3184
rect 1862 3179 1863 3183
rect 1867 3179 1868 3183
rect 1862 3178 1868 3179
rect 2530 3183 2536 3184
rect 2530 3179 2531 3183
rect 2535 3182 2536 3183
rect 3471 3183 3477 3184
rect 2535 3180 2609 3182
rect 2535 3179 2536 3180
rect 2530 3178 2536 3179
rect 3471 3179 3472 3183
rect 3476 3182 3477 3183
rect 3574 3183 3580 3184
rect 3476 3180 3497 3182
rect 3476 3179 3477 3180
rect 3471 3178 3477 3179
rect 3574 3179 3575 3183
rect 3579 3179 3580 3183
rect 3574 3178 3580 3179
rect 1886 3173 1892 3174
rect 439 3171 445 3172
rect 439 3167 440 3171
rect 444 3170 445 3171
rect 486 3171 492 3172
rect 486 3170 487 3171
rect 444 3168 487 3170
rect 444 3167 445 3168
rect 439 3166 445 3167
rect 486 3167 487 3168
rect 491 3167 492 3171
rect 486 3166 492 3167
rect 511 3171 517 3172
rect 511 3167 512 3171
rect 516 3170 517 3171
rect 551 3171 557 3172
rect 551 3170 552 3171
rect 516 3168 552 3170
rect 516 3167 517 3168
rect 511 3166 517 3167
rect 551 3167 552 3168
rect 556 3167 557 3171
rect 551 3166 557 3167
rect 647 3171 653 3172
rect 647 3167 648 3171
rect 652 3170 653 3171
rect 679 3171 685 3172
rect 679 3170 680 3171
rect 652 3168 680 3170
rect 652 3167 653 3168
rect 647 3166 653 3167
rect 679 3167 680 3168
rect 684 3167 685 3171
rect 679 3166 685 3167
rect 751 3171 757 3172
rect 751 3167 752 3171
rect 756 3170 757 3171
rect 815 3171 821 3172
rect 815 3170 816 3171
rect 756 3168 816 3170
rect 756 3167 757 3168
rect 751 3166 757 3167
rect 815 3167 816 3168
rect 820 3167 821 3171
rect 815 3166 821 3167
rect 895 3171 901 3172
rect 895 3167 896 3171
rect 900 3170 901 3171
rect 967 3171 973 3172
rect 967 3170 968 3171
rect 900 3168 968 3170
rect 900 3167 901 3168
rect 895 3166 901 3167
rect 967 3167 968 3168
rect 972 3167 973 3171
rect 967 3166 973 3167
rect 1127 3171 1133 3172
rect 1127 3167 1128 3171
rect 1132 3170 1133 3171
rect 1207 3171 1213 3172
rect 1207 3170 1208 3171
rect 1132 3168 1208 3170
rect 1132 3167 1133 3168
rect 1127 3166 1133 3167
rect 1207 3167 1208 3168
rect 1212 3167 1213 3171
rect 1207 3166 1213 3167
rect 1287 3171 1293 3172
rect 1287 3167 1288 3171
rect 1292 3170 1293 3171
rect 1366 3171 1372 3172
rect 1366 3170 1367 3171
rect 1292 3168 1367 3170
rect 1292 3167 1293 3168
rect 1287 3166 1293 3167
rect 1366 3167 1367 3168
rect 1371 3167 1372 3171
rect 1366 3166 1372 3167
rect 1455 3171 1461 3172
rect 1455 3167 1456 3171
rect 1460 3170 1461 3171
rect 1538 3171 1544 3172
rect 1538 3170 1539 3171
rect 1460 3168 1539 3170
rect 1460 3167 1461 3168
rect 1455 3166 1461 3167
rect 1538 3167 1539 3168
rect 1543 3167 1544 3171
rect 1538 3166 1544 3167
rect 1631 3171 1637 3172
rect 1631 3167 1632 3171
rect 1636 3170 1637 3171
rect 1646 3171 1652 3172
rect 1646 3170 1647 3171
rect 1636 3168 1647 3170
rect 1636 3167 1637 3168
rect 1631 3166 1637 3167
rect 1646 3167 1647 3168
rect 1651 3167 1652 3171
rect 1886 3169 1887 3173
rect 1891 3169 1892 3173
rect 1886 3168 1892 3169
rect 2014 3173 2020 3174
rect 2014 3169 2015 3173
rect 2019 3169 2020 3173
rect 2014 3168 2020 3169
rect 2166 3173 2172 3174
rect 2166 3169 2167 3173
rect 2171 3169 2172 3173
rect 2166 3168 2172 3169
rect 2318 3173 2324 3174
rect 2318 3169 2319 3173
rect 2323 3169 2324 3173
rect 2318 3168 2324 3169
rect 2454 3173 2460 3174
rect 2454 3169 2455 3173
rect 2459 3169 2460 3173
rect 2454 3168 2460 3169
rect 2590 3173 2596 3174
rect 2590 3169 2591 3173
rect 2595 3169 2596 3173
rect 2590 3168 2596 3169
rect 2726 3173 2732 3174
rect 2726 3169 2727 3173
rect 2731 3169 2732 3173
rect 2726 3168 2732 3169
rect 2862 3173 2868 3174
rect 2862 3169 2863 3173
rect 2867 3169 2868 3173
rect 2862 3168 2868 3169
rect 3006 3173 3012 3174
rect 3006 3169 3007 3173
rect 3011 3169 3012 3173
rect 3006 3168 3012 3169
rect 3158 3173 3164 3174
rect 3158 3169 3159 3173
rect 3163 3169 3164 3173
rect 3158 3168 3164 3169
rect 3318 3173 3324 3174
rect 3318 3169 3319 3173
rect 3323 3169 3324 3173
rect 3318 3168 3324 3169
rect 3478 3173 3484 3174
rect 3478 3169 3479 3173
rect 3483 3169 3484 3173
rect 3478 3168 3484 3169
rect 1646 3166 1652 3167
rect 446 3161 452 3162
rect 446 3157 447 3161
rect 451 3157 452 3161
rect 446 3156 452 3157
rect 558 3161 564 3162
rect 558 3157 559 3161
rect 563 3157 564 3161
rect 558 3156 564 3157
rect 686 3161 692 3162
rect 686 3157 687 3161
rect 691 3157 692 3161
rect 686 3156 692 3157
rect 822 3161 828 3162
rect 822 3157 823 3161
rect 827 3157 828 3161
rect 822 3156 828 3157
rect 974 3161 980 3162
rect 974 3157 975 3161
rect 979 3157 980 3161
rect 974 3156 980 3157
rect 1134 3161 1140 3162
rect 1134 3157 1135 3161
rect 1139 3157 1140 3161
rect 1134 3156 1140 3157
rect 1294 3161 1300 3162
rect 1294 3157 1295 3161
rect 1299 3157 1300 3161
rect 1294 3156 1300 3157
rect 1462 3161 1468 3162
rect 1462 3157 1463 3161
rect 1467 3157 1468 3161
rect 1462 3156 1468 3157
rect 1638 3161 1644 3162
rect 1638 3157 1639 3161
rect 1643 3157 1644 3161
rect 1638 3156 1644 3157
rect 110 3148 116 3149
rect 1822 3148 1828 3149
rect 110 3144 111 3148
rect 115 3144 116 3148
rect 511 3147 517 3148
rect 511 3146 512 3147
rect 501 3144 512 3146
rect 110 3143 116 3144
rect 511 3143 512 3144
rect 516 3143 517 3147
rect 647 3147 653 3148
rect 647 3146 648 3147
rect 613 3144 648 3146
rect 511 3142 517 3143
rect 647 3143 648 3144
rect 652 3143 653 3147
rect 751 3147 757 3148
rect 751 3146 752 3147
rect 741 3144 752 3146
rect 647 3142 653 3143
rect 751 3143 752 3144
rect 756 3143 757 3147
rect 895 3147 901 3148
rect 895 3146 896 3147
rect 877 3144 896 3146
rect 751 3142 757 3143
rect 895 3143 896 3144
rect 900 3143 901 3147
rect 1199 3147 1205 3148
rect 1199 3146 1200 3147
rect 1189 3144 1200 3146
rect 895 3142 901 3143
rect 1199 3143 1200 3144
rect 1204 3143 1205 3147
rect 1822 3144 1823 3148
rect 1827 3144 1828 3148
rect 1199 3142 1205 3143
rect 1207 3143 1213 3144
rect 1207 3139 1208 3143
rect 1212 3142 1213 3143
rect 1538 3143 1544 3144
rect 1822 3143 1828 3144
rect 1886 3147 1892 3148
rect 1886 3143 1887 3147
rect 1891 3143 1892 3147
rect 1212 3140 1313 3142
rect 1212 3139 1213 3140
rect 1207 3138 1213 3139
rect 1538 3139 1539 3143
rect 1543 3142 1544 3143
rect 1886 3142 1892 3143
rect 2046 3147 2052 3148
rect 2046 3143 2047 3147
rect 2051 3143 2052 3147
rect 2046 3142 2052 3143
rect 2198 3147 2204 3148
rect 2198 3143 2199 3147
rect 2203 3143 2204 3147
rect 2198 3142 2204 3143
rect 2350 3147 2356 3148
rect 2350 3143 2351 3147
rect 2355 3143 2356 3147
rect 2350 3142 2356 3143
rect 2510 3147 2516 3148
rect 2510 3143 2511 3147
rect 2515 3143 2516 3147
rect 2510 3142 2516 3143
rect 2678 3147 2684 3148
rect 2678 3143 2679 3147
rect 2683 3143 2684 3147
rect 2678 3142 2684 3143
rect 2870 3147 2876 3148
rect 2870 3143 2871 3147
rect 2875 3143 2876 3147
rect 2870 3142 2876 3143
rect 3070 3147 3076 3148
rect 3070 3143 3071 3147
rect 3075 3143 3076 3147
rect 3070 3142 3076 3143
rect 3286 3147 3292 3148
rect 3286 3143 3287 3147
rect 3291 3143 3292 3147
rect 3286 3142 3292 3143
rect 3478 3147 3484 3148
rect 3478 3143 3479 3147
rect 3483 3143 3484 3147
rect 3478 3142 3484 3143
rect 1543 3140 1657 3142
rect 1543 3139 1544 3140
rect 1538 3138 1544 3139
rect 2030 3139 2036 3140
rect 1862 3137 1868 3138
rect 1862 3133 1863 3137
rect 1867 3133 1868 3137
rect 2030 3135 2031 3139
rect 2035 3138 2036 3139
rect 2790 3139 2796 3140
rect 2035 3136 2065 3138
rect 2035 3135 2036 3136
rect 2030 3134 2036 3135
rect 2790 3135 2791 3139
rect 2795 3138 2796 3139
rect 2795 3136 2889 3138
rect 3574 3137 3580 3138
rect 2795 3135 2796 3136
rect 2790 3134 2796 3135
rect 1862 3132 1868 3133
rect 3574 3133 3575 3137
rect 3579 3133 3580 3137
rect 3574 3132 3580 3133
rect 110 3131 116 3132
rect 110 3127 111 3131
rect 115 3127 116 3131
rect 110 3126 116 3127
rect 890 3131 896 3132
rect 890 3127 891 3131
rect 895 3130 896 3131
rect 1551 3131 1557 3132
rect 1551 3130 1552 3131
rect 895 3128 985 3130
rect 1513 3128 1552 3130
rect 895 3127 896 3128
rect 890 3126 896 3127
rect 1551 3127 1552 3128
rect 1556 3127 1557 3131
rect 1551 3126 1557 3127
rect 1822 3131 1828 3132
rect 1822 3127 1823 3131
rect 1827 3127 1828 3131
rect 1822 3126 1828 3127
rect 2039 3123 2045 3124
rect 2039 3122 2040 3123
rect 438 3121 444 3122
rect 438 3117 439 3121
rect 443 3117 444 3121
rect 438 3116 444 3117
rect 550 3121 556 3122
rect 550 3117 551 3121
rect 555 3117 556 3121
rect 550 3116 556 3117
rect 678 3121 684 3122
rect 678 3117 679 3121
rect 683 3117 684 3121
rect 678 3116 684 3117
rect 814 3121 820 3122
rect 814 3117 815 3121
rect 819 3117 820 3121
rect 814 3116 820 3117
rect 966 3121 972 3122
rect 966 3117 967 3121
rect 971 3117 972 3121
rect 966 3116 972 3117
rect 1126 3121 1132 3122
rect 1126 3117 1127 3121
rect 1131 3117 1132 3121
rect 1126 3116 1132 3117
rect 1286 3121 1292 3122
rect 1286 3117 1287 3121
rect 1291 3117 1292 3121
rect 1286 3116 1292 3117
rect 1454 3121 1460 3122
rect 1454 3117 1455 3121
rect 1459 3117 1460 3121
rect 1454 3116 1460 3117
rect 1630 3121 1636 3122
rect 1630 3117 1631 3121
rect 1635 3117 1636 3121
rect 1630 3116 1636 3117
rect 1862 3120 1868 3121
rect 1949 3120 2040 3122
rect 1862 3116 1863 3120
rect 1867 3116 1868 3120
rect 2039 3119 2040 3120
rect 2044 3119 2045 3123
rect 2343 3123 2349 3124
rect 2343 3122 2344 3123
rect 2261 3120 2344 3122
rect 2039 3118 2045 3119
rect 2343 3119 2344 3120
rect 2348 3119 2349 3123
rect 2503 3123 2509 3124
rect 2503 3122 2504 3123
rect 2413 3120 2504 3122
rect 2343 3118 2349 3119
rect 2503 3119 2504 3120
rect 2508 3119 2509 3123
rect 2671 3123 2677 3124
rect 2671 3122 2672 3123
rect 2573 3120 2672 3122
rect 2503 3118 2509 3119
rect 2671 3119 2672 3120
rect 2676 3119 2677 3123
rect 2746 3123 2752 3124
rect 2746 3122 2747 3123
rect 2741 3120 2747 3122
rect 2671 3118 2677 3119
rect 2746 3119 2747 3120
rect 2751 3119 2752 3123
rect 2746 3118 2752 3119
rect 2938 3123 2944 3124
rect 2938 3119 2939 3123
rect 2943 3122 2944 3123
rect 3175 3123 3181 3124
rect 2943 3120 3097 3122
rect 2943 3119 2944 3120
rect 2938 3118 2944 3119
rect 3175 3119 3176 3123
rect 3180 3122 3181 3123
rect 3470 3123 3476 3124
rect 3180 3120 3313 3122
rect 3180 3119 3181 3120
rect 3175 3118 3181 3119
rect 3470 3119 3471 3123
rect 3475 3122 3476 3123
rect 3475 3120 3505 3122
rect 3574 3120 3580 3121
rect 3475 3119 3476 3120
rect 3470 3118 3476 3119
rect 1862 3115 1868 3116
rect 3574 3116 3575 3120
rect 3579 3116 3580 3120
rect 3574 3115 3580 3116
rect 1894 3107 1900 3108
rect 1894 3103 1895 3107
rect 1899 3103 1900 3107
rect 1894 3102 1900 3103
rect 2054 3107 2060 3108
rect 2054 3103 2055 3107
rect 2059 3103 2060 3107
rect 2054 3102 2060 3103
rect 2206 3107 2212 3108
rect 2206 3103 2207 3107
rect 2211 3103 2212 3107
rect 2206 3102 2212 3103
rect 2358 3107 2364 3108
rect 2358 3103 2359 3107
rect 2363 3103 2364 3107
rect 2358 3102 2364 3103
rect 2518 3107 2524 3108
rect 2518 3103 2519 3107
rect 2523 3103 2524 3107
rect 2518 3102 2524 3103
rect 2686 3107 2692 3108
rect 2686 3103 2687 3107
rect 2691 3103 2692 3107
rect 2686 3102 2692 3103
rect 2878 3107 2884 3108
rect 2878 3103 2879 3107
rect 2883 3103 2884 3107
rect 2878 3102 2884 3103
rect 3078 3107 3084 3108
rect 3078 3103 3079 3107
rect 3083 3103 3084 3107
rect 3078 3102 3084 3103
rect 3294 3107 3300 3108
rect 3294 3103 3295 3107
rect 3299 3103 3300 3107
rect 3294 3102 3300 3103
rect 3486 3107 3492 3108
rect 3486 3103 3487 3107
rect 3491 3103 3492 3107
rect 3486 3102 3492 3103
rect 1887 3095 1893 3096
rect 550 3091 556 3092
rect 550 3087 551 3091
rect 555 3087 556 3091
rect 550 3086 556 3087
rect 662 3091 668 3092
rect 662 3087 663 3091
rect 667 3087 668 3091
rect 662 3086 668 3087
rect 782 3091 788 3092
rect 782 3087 783 3091
rect 787 3087 788 3091
rect 782 3086 788 3087
rect 902 3091 908 3092
rect 902 3087 903 3091
rect 907 3087 908 3091
rect 902 3086 908 3087
rect 1030 3091 1036 3092
rect 1030 3087 1031 3091
rect 1035 3087 1036 3091
rect 1030 3086 1036 3087
rect 1158 3091 1164 3092
rect 1158 3087 1159 3091
rect 1163 3087 1164 3091
rect 1158 3086 1164 3087
rect 1286 3091 1292 3092
rect 1286 3087 1287 3091
rect 1291 3087 1292 3091
rect 1286 3086 1292 3087
rect 1422 3091 1428 3092
rect 1422 3087 1423 3091
rect 1427 3087 1428 3091
rect 1422 3086 1428 3087
rect 1558 3091 1564 3092
rect 1558 3087 1559 3091
rect 1563 3087 1564 3091
rect 1558 3086 1564 3087
rect 1694 3091 1700 3092
rect 1694 3087 1695 3091
rect 1699 3087 1700 3091
rect 1887 3091 1888 3095
rect 1892 3094 1893 3095
rect 1895 3095 1901 3096
rect 1895 3094 1896 3095
rect 1892 3092 1896 3094
rect 1892 3091 1893 3092
rect 1887 3090 1893 3091
rect 1895 3091 1896 3092
rect 1900 3091 1901 3095
rect 1895 3090 1901 3091
rect 2039 3095 2045 3096
rect 2039 3091 2040 3095
rect 2044 3094 2045 3095
rect 2047 3095 2053 3096
rect 2047 3094 2048 3095
rect 2044 3092 2048 3094
rect 2044 3091 2045 3092
rect 2039 3090 2045 3091
rect 2047 3091 2048 3092
rect 2052 3091 2053 3095
rect 2047 3090 2053 3091
rect 2199 3095 2205 3096
rect 2199 3091 2200 3095
rect 2204 3094 2205 3095
rect 2214 3095 2220 3096
rect 2214 3094 2215 3095
rect 2204 3092 2215 3094
rect 2204 3091 2205 3092
rect 2199 3090 2205 3091
rect 2214 3091 2215 3092
rect 2219 3091 2220 3095
rect 2214 3090 2220 3091
rect 2343 3095 2349 3096
rect 2343 3091 2344 3095
rect 2348 3094 2349 3095
rect 2351 3095 2357 3096
rect 2351 3094 2352 3095
rect 2348 3092 2352 3094
rect 2348 3091 2349 3092
rect 2343 3090 2349 3091
rect 2351 3091 2352 3092
rect 2356 3091 2357 3095
rect 2351 3090 2357 3091
rect 2503 3095 2509 3096
rect 2503 3091 2504 3095
rect 2508 3094 2509 3095
rect 2511 3095 2517 3096
rect 2511 3094 2512 3095
rect 2508 3092 2512 3094
rect 2508 3091 2509 3092
rect 2503 3090 2509 3091
rect 2511 3091 2512 3092
rect 2516 3091 2517 3095
rect 2511 3090 2517 3091
rect 2671 3095 2677 3096
rect 2671 3091 2672 3095
rect 2676 3094 2677 3095
rect 2679 3095 2685 3096
rect 2679 3094 2680 3095
rect 2676 3092 2680 3094
rect 2676 3091 2677 3092
rect 2671 3090 2677 3091
rect 2679 3091 2680 3092
rect 2684 3091 2685 3095
rect 2679 3090 2685 3091
rect 2871 3095 2877 3096
rect 2871 3091 2872 3095
rect 2876 3094 2877 3095
rect 2938 3095 2944 3096
rect 2938 3094 2939 3095
rect 2876 3092 2939 3094
rect 2876 3091 2877 3092
rect 2871 3090 2877 3091
rect 2938 3091 2939 3092
rect 2943 3091 2944 3095
rect 2938 3090 2944 3091
rect 3071 3095 3077 3096
rect 3071 3091 3072 3095
rect 3076 3094 3077 3095
rect 3175 3095 3181 3096
rect 3175 3094 3176 3095
rect 3076 3092 3176 3094
rect 3076 3091 3077 3092
rect 3071 3090 3077 3091
rect 3175 3091 3176 3092
rect 3180 3091 3181 3095
rect 3175 3090 3181 3091
rect 3287 3095 3293 3096
rect 3287 3091 3288 3095
rect 3292 3094 3293 3095
rect 3302 3095 3308 3096
rect 3302 3094 3303 3095
rect 3292 3092 3303 3094
rect 3292 3091 3293 3092
rect 3287 3090 3293 3091
rect 3302 3091 3303 3092
rect 3307 3091 3308 3095
rect 3302 3090 3308 3091
rect 3471 3095 3477 3096
rect 3471 3091 3472 3095
rect 3476 3094 3477 3095
rect 3479 3095 3485 3096
rect 3479 3094 3480 3095
rect 3476 3092 3480 3094
rect 3476 3091 3477 3092
rect 3471 3090 3477 3091
rect 3479 3091 3480 3092
rect 3484 3091 3485 3095
rect 3479 3090 3485 3091
rect 1694 3086 1700 3087
rect 1366 3083 1372 3084
rect 110 3081 116 3082
rect 110 3077 111 3081
rect 115 3077 116 3081
rect 1366 3079 1367 3083
rect 1371 3082 1372 3083
rect 1371 3080 1441 3082
rect 1822 3081 1828 3082
rect 1371 3079 1372 3080
rect 1366 3078 1372 3079
rect 110 3076 116 3077
rect 1822 3077 1823 3081
rect 1827 3077 1828 3081
rect 1822 3076 1828 3077
rect 1911 3075 1917 3076
rect 1911 3071 1912 3075
rect 1916 3074 1917 3075
rect 2006 3075 2012 3076
rect 2006 3074 2007 3075
rect 1916 3072 2007 3074
rect 1916 3071 1917 3072
rect 1911 3070 1917 3071
rect 2006 3071 2007 3072
rect 2011 3071 2012 3075
rect 2006 3070 2012 3071
rect 2079 3075 2085 3076
rect 2079 3071 2080 3075
rect 2084 3074 2085 3075
rect 2182 3075 2188 3076
rect 2182 3074 2183 3075
rect 2084 3072 2183 3074
rect 2084 3071 2085 3072
rect 2079 3070 2085 3071
rect 2182 3071 2183 3072
rect 2187 3071 2188 3075
rect 2182 3070 2188 3071
rect 2263 3075 2269 3076
rect 2263 3071 2264 3075
rect 2268 3074 2269 3075
rect 2271 3075 2277 3076
rect 2271 3074 2272 3075
rect 2268 3072 2272 3074
rect 2268 3071 2269 3072
rect 2263 3070 2269 3071
rect 2271 3071 2272 3072
rect 2276 3071 2277 3075
rect 2271 3070 2277 3071
rect 2479 3075 2485 3076
rect 2479 3071 2480 3075
rect 2484 3074 2485 3075
rect 2502 3075 2508 3076
rect 2502 3074 2503 3075
rect 2484 3072 2503 3074
rect 2484 3071 2485 3072
rect 2479 3070 2485 3071
rect 2502 3071 2503 3072
rect 2507 3071 2508 3075
rect 2502 3070 2508 3071
rect 2711 3075 2717 3076
rect 2711 3071 2712 3075
rect 2716 3074 2717 3075
rect 2746 3075 2752 3076
rect 2746 3074 2747 3075
rect 2716 3072 2747 3074
rect 2716 3071 2717 3072
rect 2711 3070 2717 3071
rect 2746 3071 2747 3072
rect 2751 3071 2752 3075
rect 2746 3070 2752 3071
rect 2847 3075 2853 3076
rect 2847 3071 2848 3075
rect 2852 3074 2853 3075
rect 2967 3075 2973 3076
rect 2967 3074 2968 3075
rect 2852 3072 2968 3074
rect 2852 3071 2853 3072
rect 2847 3070 2853 3071
rect 2967 3071 2968 3072
rect 2972 3071 2973 3075
rect 2967 3070 2973 3071
rect 3231 3075 3237 3076
rect 3231 3071 3232 3075
rect 3236 3074 3237 3075
rect 3246 3075 3252 3076
rect 3246 3074 3247 3075
rect 3236 3072 3247 3074
rect 3236 3071 3237 3072
rect 3231 3070 3237 3071
rect 3246 3071 3247 3072
rect 3251 3071 3252 3075
rect 3246 3070 3252 3071
rect 3470 3075 3476 3076
rect 3470 3071 3471 3075
rect 3475 3074 3476 3075
rect 3479 3075 3485 3076
rect 3479 3074 3480 3075
rect 3475 3072 3480 3074
rect 3475 3071 3476 3072
rect 3470 3070 3476 3071
rect 3479 3071 3480 3072
rect 3484 3071 3485 3075
rect 3479 3070 3485 3071
rect 655 3067 661 3068
rect 655 3066 656 3067
rect 110 3064 116 3065
rect 613 3064 656 3066
rect 110 3060 111 3064
rect 115 3060 116 3064
rect 655 3063 656 3064
rect 660 3063 661 3067
rect 775 3067 781 3068
rect 775 3066 776 3067
rect 725 3064 776 3066
rect 655 3062 661 3063
rect 775 3063 776 3064
rect 780 3063 781 3067
rect 895 3067 901 3068
rect 895 3066 896 3067
rect 845 3064 896 3066
rect 775 3062 781 3063
rect 895 3063 896 3064
rect 900 3063 901 3067
rect 1023 3067 1029 3068
rect 1023 3066 1024 3067
rect 965 3064 1024 3066
rect 895 3062 901 3063
rect 1023 3063 1024 3064
rect 1028 3063 1029 3067
rect 1103 3067 1109 3068
rect 1103 3066 1104 3067
rect 1093 3064 1104 3066
rect 1023 3062 1029 3063
rect 1103 3063 1104 3064
rect 1108 3063 1109 3067
rect 1279 3067 1285 3068
rect 1279 3066 1280 3067
rect 1221 3064 1280 3066
rect 1103 3062 1109 3063
rect 1279 3063 1280 3064
rect 1284 3063 1285 3067
rect 1415 3067 1421 3068
rect 1415 3066 1416 3067
rect 1349 3064 1416 3066
rect 1279 3062 1285 3063
rect 1415 3063 1416 3064
rect 1420 3063 1421 3067
rect 1687 3067 1693 3068
rect 1687 3066 1688 3067
rect 1621 3064 1688 3066
rect 1415 3062 1421 3063
rect 1687 3063 1688 3064
rect 1692 3063 1693 3067
rect 1762 3067 1768 3068
rect 1762 3066 1763 3067
rect 1757 3064 1763 3066
rect 1687 3062 1693 3063
rect 1762 3063 1763 3064
rect 1767 3063 1768 3067
rect 1918 3065 1924 3066
rect 1762 3062 1768 3063
rect 1822 3064 1828 3065
rect 110 3059 116 3060
rect 1822 3060 1823 3064
rect 1827 3060 1828 3064
rect 1918 3061 1919 3065
rect 1923 3061 1924 3065
rect 1918 3060 1924 3061
rect 2086 3065 2092 3066
rect 2086 3061 2087 3065
rect 2091 3061 2092 3065
rect 2086 3060 2092 3061
rect 2278 3065 2284 3066
rect 2278 3061 2279 3065
rect 2283 3061 2284 3065
rect 2278 3060 2284 3061
rect 2486 3065 2492 3066
rect 2486 3061 2487 3065
rect 2491 3061 2492 3065
rect 2486 3060 2492 3061
rect 2718 3065 2724 3066
rect 2718 3061 2719 3065
rect 2723 3061 2724 3065
rect 2718 3060 2724 3061
rect 2974 3065 2980 3066
rect 2974 3061 2975 3065
rect 2979 3061 2980 3065
rect 2974 3060 2980 3061
rect 3238 3065 3244 3066
rect 3238 3061 3239 3065
rect 3243 3061 3244 3065
rect 3238 3060 3244 3061
rect 3486 3065 3492 3066
rect 3486 3061 3487 3065
rect 3491 3061 3492 3065
rect 3486 3060 3492 3061
rect 1822 3059 1828 3060
rect 1862 3052 1868 3053
rect 3574 3052 3580 3053
rect 558 3051 564 3052
rect 558 3047 559 3051
rect 563 3047 564 3051
rect 558 3046 564 3047
rect 670 3051 676 3052
rect 670 3047 671 3051
rect 675 3047 676 3051
rect 670 3046 676 3047
rect 790 3051 796 3052
rect 790 3047 791 3051
rect 795 3047 796 3051
rect 790 3046 796 3047
rect 910 3051 916 3052
rect 910 3047 911 3051
rect 915 3047 916 3051
rect 910 3046 916 3047
rect 1038 3051 1044 3052
rect 1038 3047 1039 3051
rect 1043 3047 1044 3051
rect 1038 3046 1044 3047
rect 1166 3051 1172 3052
rect 1166 3047 1167 3051
rect 1171 3047 1172 3051
rect 1166 3046 1172 3047
rect 1294 3051 1300 3052
rect 1294 3047 1295 3051
rect 1299 3047 1300 3051
rect 1294 3046 1300 3047
rect 1430 3051 1436 3052
rect 1430 3047 1431 3051
rect 1435 3047 1436 3051
rect 1430 3046 1436 3047
rect 1566 3051 1572 3052
rect 1566 3047 1567 3051
rect 1571 3047 1572 3051
rect 1566 3046 1572 3047
rect 1702 3051 1708 3052
rect 1702 3047 1703 3051
rect 1707 3047 1708 3051
rect 1862 3048 1863 3052
rect 1867 3048 1868 3052
rect 2847 3051 2853 3052
rect 2847 3050 2848 3051
rect 2773 3048 2848 3050
rect 1862 3047 1868 3048
rect 1895 3047 1901 3048
rect 1702 3046 1708 3047
rect 1895 3043 1896 3047
rect 1900 3046 1901 3047
rect 2006 3047 2012 3048
rect 1900 3044 1937 3046
rect 1900 3043 1901 3044
rect 1895 3042 1901 3043
rect 2006 3043 2007 3047
rect 2011 3046 2012 3047
rect 2182 3047 2188 3048
rect 2011 3044 2105 3046
rect 2011 3043 2012 3044
rect 2006 3042 2012 3043
rect 2182 3043 2183 3047
rect 2187 3046 2188 3047
rect 2847 3047 2848 3048
rect 2852 3047 2853 3051
rect 3302 3051 3308 3052
rect 3302 3050 3303 3051
rect 3293 3048 3303 3050
rect 2847 3046 2853 3047
rect 2898 3047 2904 3048
rect 2187 3044 2297 3046
rect 2187 3043 2188 3044
rect 2182 3042 2188 3043
rect 2898 3043 2899 3047
rect 2903 3046 2904 3047
rect 3302 3047 3303 3048
rect 3307 3047 3308 3051
rect 3574 3048 3575 3052
rect 3579 3048 3580 3052
rect 3574 3047 3580 3048
rect 3302 3046 3308 3047
rect 2903 3044 2993 3046
rect 2903 3043 2904 3044
rect 2898 3042 2904 3043
rect 551 3039 557 3040
rect 551 3035 552 3039
rect 556 3038 557 3039
rect 566 3039 572 3040
rect 566 3038 567 3039
rect 556 3036 567 3038
rect 556 3035 557 3036
rect 551 3034 557 3035
rect 566 3035 567 3036
rect 571 3035 572 3039
rect 566 3034 572 3035
rect 655 3039 661 3040
rect 655 3035 656 3039
rect 660 3038 661 3039
rect 663 3039 669 3040
rect 663 3038 664 3039
rect 660 3036 664 3038
rect 660 3035 661 3036
rect 655 3034 661 3035
rect 663 3035 664 3036
rect 668 3035 669 3039
rect 663 3034 669 3035
rect 775 3039 781 3040
rect 775 3035 776 3039
rect 780 3038 781 3039
rect 783 3039 789 3040
rect 783 3038 784 3039
rect 780 3036 784 3038
rect 780 3035 781 3036
rect 775 3034 781 3035
rect 783 3035 784 3036
rect 788 3035 789 3039
rect 783 3034 789 3035
rect 895 3039 901 3040
rect 895 3035 896 3039
rect 900 3038 901 3039
rect 903 3039 909 3040
rect 903 3038 904 3039
rect 900 3036 904 3038
rect 900 3035 901 3036
rect 895 3034 901 3035
rect 903 3035 904 3036
rect 908 3035 909 3039
rect 903 3034 909 3035
rect 1023 3039 1029 3040
rect 1023 3035 1024 3039
rect 1028 3038 1029 3039
rect 1031 3039 1037 3040
rect 1031 3038 1032 3039
rect 1028 3036 1032 3038
rect 1028 3035 1029 3036
rect 1023 3034 1029 3035
rect 1031 3035 1032 3036
rect 1036 3035 1037 3039
rect 1031 3034 1037 3035
rect 1159 3039 1165 3040
rect 1159 3035 1160 3039
rect 1164 3038 1165 3039
rect 1174 3039 1180 3040
rect 1174 3038 1175 3039
rect 1164 3036 1175 3038
rect 1164 3035 1165 3036
rect 1159 3034 1165 3035
rect 1174 3035 1175 3036
rect 1179 3035 1180 3039
rect 1174 3034 1180 3035
rect 1279 3039 1285 3040
rect 1279 3035 1280 3039
rect 1284 3038 1285 3039
rect 1287 3039 1293 3040
rect 1287 3038 1288 3039
rect 1284 3036 1288 3038
rect 1284 3035 1285 3036
rect 1279 3034 1285 3035
rect 1287 3035 1288 3036
rect 1292 3035 1293 3039
rect 1287 3034 1293 3035
rect 1415 3039 1421 3040
rect 1415 3035 1416 3039
rect 1420 3038 1421 3039
rect 1423 3039 1429 3040
rect 1423 3038 1424 3039
rect 1420 3036 1424 3038
rect 1420 3035 1421 3036
rect 1415 3034 1421 3035
rect 1423 3035 1424 3036
rect 1428 3035 1429 3039
rect 1423 3034 1429 3035
rect 1551 3039 1557 3040
rect 1551 3035 1552 3039
rect 1556 3038 1557 3039
rect 1559 3039 1565 3040
rect 1559 3038 1560 3039
rect 1556 3036 1560 3038
rect 1556 3035 1557 3036
rect 1551 3034 1557 3035
rect 1559 3035 1560 3036
rect 1564 3035 1565 3039
rect 1559 3034 1565 3035
rect 1687 3039 1693 3040
rect 1687 3035 1688 3039
rect 1692 3038 1693 3039
rect 1695 3039 1701 3040
rect 1695 3038 1696 3039
rect 1692 3036 1696 3038
rect 1692 3035 1693 3036
rect 1687 3034 1693 3035
rect 1695 3035 1696 3036
rect 1700 3035 1701 3039
rect 1695 3034 1701 3035
rect 1862 3035 1868 3036
rect 1862 3031 1863 3035
rect 1867 3031 1868 3035
rect 1862 3030 1868 3031
rect 2430 3035 2436 3036
rect 2430 3031 2431 3035
rect 2435 3034 2436 3035
rect 3471 3035 3477 3036
rect 2435 3032 2497 3034
rect 2435 3031 2436 3032
rect 2430 3030 2436 3031
rect 3471 3031 3472 3035
rect 3476 3034 3477 3035
rect 3574 3035 3580 3036
rect 3476 3032 3497 3034
rect 3476 3031 3477 3032
rect 3471 3030 3477 3031
rect 3574 3031 3575 3035
rect 3579 3031 3580 3035
rect 3574 3030 3580 3031
rect 1910 3025 1916 3026
rect 567 3023 573 3024
rect 567 3019 568 3023
rect 572 3022 573 3023
rect 663 3023 669 3024
rect 663 3022 664 3023
rect 572 3020 664 3022
rect 572 3019 573 3020
rect 567 3018 573 3019
rect 663 3019 664 3020
rect 668 3019 669 3023
rect 663 3018 669 3019
rect 695 3023 701 3024
rect 695 3019 696 3023
rect 700 3022 701 3023
rect 770 3023 776 3024
rect 770 3022 771 3023
rect 700 3020 771 3022
rect 700 3019 701 3020
rect 695 3018 701 3019
rect 770 3019 771 3020
rect 775 3019 776 3023
rect 770 3018 776 3019
rect 823 3023 829 3024
rect 823 3019 824 3023
rect 828 3022 829 3023
rect 898 3023 904 3024
rect 898 3022 899 3023
rect 828 3020 899 3022
rect 828 3019 829 3020
rect 823 3018 829 3019
rect 898 3019 899 3020
rect 903 3019 904 3023
rect 898 3018 904 3019
rect 959 3023 965 3024
rect 959 3019 960 3023
rect 964 3022 965 3023
rect 1039 3023 1045 3024
rect 1039 3022 1040 3023
rect 964 3020 1040 3022
rect 964 3019 965 3020
rect 959 3018 965 3019
rect 1039 3019 1040 3020
rect 1044 3019 1045 3023
rect 1039 3018 1045 3019
rect 1095 3023 1101 3024
rect 1095 3019 1096 3023
rect 1100 3022 1101 3023
rect 1103 3023 1109 3024
rect 1103 3022 1104 3023
rect 1100 3020 1104 3022
rect 1100 3019 1101 3020
rect 1095 3018 1101 3019
rect 1103 3019 1104 3020
rect 1108 3019 1109 3023
rect 1103 3018 1109 3019
rect 1231 3023 1237 3024
rect 1231 3019 1232 3023
rect 1236 3022 1237 3023
rect 1306 3023 1312 3024
rect 1306 3022 1307 3023
rect 1236 3020 1307 3022
rect 1236 3019 1237 3020
rect 1231 3018 1237 3019
rect 1306 3019 1307 3020
rect 1311 3019 1312 3023
rect 1306 3018 1312 3019
rect 1359 3023 1365 3024
rect 1359 3019 1360 3023
rect 1364 3022 1365 3023
rect 1438 3023 1444 3024
rect 1438 3022 1439 3023
rect 1364 3020 1439 3022
rect 1364 3019 1365 3020
rect 1359 3018 1365 3019
rect 1438 3019 1439 3020
rect 1443 3019 1444 3023
rect 1438 3018 1444 3019
rect 1487 3023 1493 3024
rect 1487 3019 1488 3023
rect 1492 3022 1493 3023
rect 1567 3023 1573 3024
rect 1567 3022 1568 3023
rect 1492 3020 1568 3022
rect 1492 3019 1493 3020
rect 1487 3018 1493 3019
rect 1567 3019 1568 3020
rect 1572 3019 1573 3023
rect 1567 3018 1573 3019
rect 1594 3023 1600 3024
rect 1594 3019 1595 3023
rect 1599 3022 1600 3023
rect 1615 3023 1621 3024
rect 1615 3022 1616 3023
rect 1599 3020 1616 3022
rect 1599 3019 1600 3020
rect 1594 3018 1600 3019
rect 1615 3019 1616 3020
rect 1620 3019 1621 3023
rect 1615 3018 1621 3019
rect 1727 3023 1733 3024
rect 1727 3019 1728 3023
rect 1732 3022 1733 3023
rect 1762 3023 1768 3024
rect 1762 3022 1763 3023
rect 1732 3020 1763 3022
rect 1732 3019 1733 3020
rect 1727 3018 1733 3019
rect 1762 3019 1763 3020
rect 1767 3019 1768 3023
rect 1910 3021 1911 3025
rect 1915 3021 1916 3025
rect 1910 3020 1916 3021
rect 2078 3025 2084 3026
rect 2078 3021 2079 3025
rect 2083 3021 2084 3025
rect 2078 3020 2084 3021
rect 2270 3025 2276 3026
rect 2270 3021 2271 3025
rect 2275 3021 2276 3025
rect 2270 3020 2276 3021
rect 2478 3025 2484 3026
rect 2478 3021 2479 3025
rect 2483 3021 2484 3025
rect 2478 3020 2484 3021
rect 2710 3025 2716 3026
rect 2710 3021 2711 3025
rect 2715 3021 2716 3025
rect 2710 3020 2716 3021
rect 2966 3025 2972 3026
rect 2966 3021 2967 3025
rect 2971 3021 2972 3025
rect 2966 3020 2972 3021
rect 3230 3025 3236 3026
rect 3230 3021 3231 3025
rect 3235 3021 3236 3025
rect 3230 3020 3236 3021
rect 3478 3025 3484 3026
rect 3478 3021 3479 3025
rect 3483 3021 3484 3025
rect 3478 3020 3484 3021
rect 1762 3018 1768 3019
rect 574 3013 580 3014
rect 574 3009 575 3013
rect 579 3009 580 3013
rect 574 3008 580 3009
rect 702 3013 708 3014
rect 702 3009 703 3013
rect 707 3009 708 3013
rect 702 3008 708 3009
rect 830 3013 836 3014
rect 830 3009 831 3013
rect 835 3009 836 3013
rect 830 3008 836 3009
rect 966 3013 972 3014
rect 966 3009 967 3013
rect 971 3009 972 3013
rect 966 3008 972 3009
rect 1102 3013 1108 3014
rect 1102 3009 1103 3013
rect 1107 3009 1108 3013
rect 1102 3008 1108 3009
rect 1238 3013 1244 3014
rect 1238 3009 1239 3013
rect 1243 3009 1244 3013
rect 1238 3008 1244 3009
rect 1366 3013 1372 3014
rect 1366 3009 1367 3013
rect 1371 3009 1372 3013
rect 1366 3008 1372 3009
rect 1494 3013 1500 3014
rect 1494 3009 1495 3013
rect 1499 3009 1500 3013
rect 1494 3008 1500 3009
rect 1622 3013 1628 3014
rect 1622 3009 1623 3013
rect 1627 3009 1628 3013
rect 1622 3008 1628 3009
rect 1734 3013 1740 3014
rect 1734 3009 1735 3013
rect 1739 3009 1740 3013
rect 1734 3008 1740 3009
rect 110 3000 116 3001
rect 110 2996 111 3000
rect 115 2996 116 3000
rect 1822 3000 1828 3001
rect 1822 2996 1823 3000
rect 1827 2996 1828 3000
rect 110 2995 116 2996
rect 663 2995 669 2996
rect 663 2991 664 2995
rect 668 2994 669 2995
rect 770 2995 776 2996
rect 668 2992 721 2994
rect 668 2991 669 2992
rect 663 2990 669 2991
rect 770 2991 771 2995
rect 775 2994 776 2995
rect 898 2995 904 2996
rect 775 2992 849 2994
rect 775 2991 776 2992
rect 770 2990 776 2991
rect 898 2991 899 2995
rect 903 2994 904 2995
rect 1039 2995 1045 2996
rect 903 2992 985 2994
rect 903 2991 904 2992
rect 898 2990 904 2991
rect 1039 2991 1040 2995
rect 1044 2994 1045 2995
rect 1174 2995 1180 2996
rect 1044 2992 1121 2994
rect 1044 2991 1045 2992
rect 1039 2990 1045 2991
rect 1174 2991 1175 2995
rect 1179 2994 1180 2995
rect 1306 2995 1312 2996
rect 1179 2992 1257 2994
rect 1179 2991 1180 2992
rect 1174 2990 1180 2991
rect 1306 2991 1307 2995
rect 1311 2994 1312 2995
rect 1438 2995 1444 2996
rect 1311 2992 1385 2994
rect 1311 2991 1312 2992
rect 1306 2990 1312 2991
rect 1438 2991 1439 2995
rect 1443 2994 1444 2995
rect 1567 2995 1573 2996
rect 1822 2995 1828 2996
rect 2022 2999 2028 3000
rect 2022 2995 2023 2999
rect 2027 2995 2028 2999
rect 1443 2992 1513 2994
rect 1443 2991 1444 2992
rect 1438 2990 1444 2991
rect 1567 2991 1568 2995
rect 1572 2994 1573 2995
rect 2022 2994 2028 2995
rect 2158 2999 2164 3000
rect 2158 2995 2159 2999
rect 2163 2995 2164 2999
rect 2158 2994 2164 2995
rect 2286 2999 2292 3000
rect 2286 2995 2287 2999
rect 2291 2995 2292 2999
rect 2286 2994 2292 2995
rect 2414 2999 2420 3000
rect 2414 2995 2415 2999
rect 2419 2995 2420 2999
rect 2414 2994 2420 2995
rect 2534 2999 2540 3000
rect 2534 2995 2535 2999
rect 2539 2995 2540 2999
rect 2534 2994 2540 2995
rect 2662 2999 2668 3000
rect 2662 2995 2663 2999
rect 2667 2995 2668 2999
rect 2662 2994 2668 2995
rect 2806 2999 2812 3000
rect 2806 2995 2807 2999
rect 2811 2995 2812 2999
rect 2806 2994 2812 2995
rect 2966 2999 2972 3000
rect 2966 2995 2967 2999
rect 2971 2995 2972 2999
rect 2966 2994 2972 2995
rect 3142 2999 3148 3000
rect 3142 2995 3143 2999
rect 3147 2995 3148 2999
rect 3142 2994 3148 2995
rect 3318 2999 3324 3000
rect 3318 2995 3319 2999
rect 3323 2995 3324 2999
rect 3318 2994 3324 2995
rect 3478 2999 3484 3000
rect 3478 2995 3479 2999
rect 3483 2995 3484 2999
rect 3478 2994 3484 2995
rect 1572 2992 1641 2994
rect 1572 2991 1573 2992
rect 1567 2990 1573 2991
rect 2263 2991 2269 2992
rect 1862 2989 1868 2990
rect 1862 2985 1863 2989
rect 1867 2985 1868 2989
rect 2263 2987 2264 2991
rect 2268 2990 2269 2991
rect 3246 2991 3252 2992
rect 2268 2988 2305 2990
rect 2268 2987 2269 2988
rect 2263 2986 2269 2987
rect 3246 2987 3247 2991
rect 3251 2990 3252 2991
rect 3251 2988 3337 2990
rect 3574 2989 3580 2990
rect 3251 2987 3252 2988
rect 3246 2986 3252 2987
rect 1862 2984 1868 2985
rect 3574 2985 3575 2989
rect 3579 2985 3580 2989
rect 3574 2984 3580 2985
rect 110 2983 116 2984
rect 110 2979 111 2983
rect 115 2979 116 2983
rect 110 2978 116 2979
rect 510 2983 516 2984
rect 510 2979 511 2983
rect 515 2982 516 2983
rect 1690 2983 1696 2984
rect 515 2980 585 2982
rect 515 2979 516 2980
rect 510 2978 516 2979
rect 1690 2979 1691 2983
rect 1695 2982 1696 2983
rect 1822 2983 1828 2984
rect 1695 2980 1745 2982
rect 1695 2979 1696 2980
rect 1690 2978 1696 2979
rect 1822 2979 1823 2983
rect 1827 2979 1828 2983
rect 1822 2978 1828 2979
rect 2151 2975 2157 2976
rect 2151 2974 2152 2975
rect 566 2973 572 2974
rect 566 2969 567 2973
rect 571 2969 572 2973
rect 566 2968 572 2969
rect 694 2973 700 2974
rect 694 2969 695 2973
rect 699 2969 700 2973
rect 694 2968 700 2969
rect 822 2973 828 2974
rect 822 2969 823 2973
rect 827 2969 828 2973
rect 822 2968 828 2969
rect 958 2973 964 2974
rect 958 2969 959 2973
rect 963 2969 964 2973
rect 958 2968 964 2969
rect 1094 2973 1100 2974
rect 1094 2969 1095 2973
rect 1099 2969 1100 2973
rect 1094 2968 1100 2969
rect 1230 2973 1236 2974
rect 1230 2969 1231 2973
rect 1235 2969 1236 2973
rect 1230 2968 1236 2969
rect 1358 2973 1364 2974
rect 1358 2969 1359 2973
rect 1363 2969 1364 2973
rect 1358 2968 1364 2969
rect 1486 2973 1492 2974
rect 1486 2969 1487 2973
rect 1491 2969 1492 2973
rect 1486 2968 1492 2969
rect 1614 2973 1620 2974
rect 1614 2969 1615 2973
rect 1619 2969 1620 2973
rect 1614 2968 1620 2969
rect 1726 2973 1732 2974
rect 1726 2969 1727 2973
rect 1731 2969 1732 2973
rect 1726 2968 1732 2969
rect 1862 2972 1868 2973
rect 2085 2972 2152 2974
rect 1862 2968 1863 2972
rect 1867 2968 1868 2972
rect 2151 2971 2152 2972
rect 2156 2971 2157 2975
rect 2279 2975 2285 2976
rect 2279 2974 2280 2975
rect 2221 2972 2280 2974
rect 2151 2970 2157 2971
rect 2279 2971 2280 2972
rect 2284 2971 2285 2975
rect 2527 2975 2533 2976
rect 2527 2974 2528 2975
rect 2477 2972 2528 2974
rect 2279 2970 2285 2971
rect 2527 2971 2528 2972
rect 2532 2971 2533 2975
rect 2655 2975 2661 2976
rect 2655 2974 2656 2975
rect 2597 2972 2656 2974
rect 2527 2970 2533 2971
rect 2655 2971 2656 2972
rect 2660 2971 2661 2975
rect 2799 2975 2805 2976
rect 2799 2974 2800 2975
rect 2725 2972 2800 2974
rect 2655 2970 2661 2971
rect 2799 2971 2800 2972
rect 2804 2971 2805 2975
rect 2959 2975 2965 2976
rect 2959 2974 2960 2975
rect 2869 2972 2960 2974
rect 2799 2970 2805 2971
rect 2959 2971 2960 2972
rect 2964 2971 2965 2975
rect 3063 2975 3069 2976
rect 3063 2974 3064 2975
rect 3029 2972 3064 2974
rect 2959 2970 2965 2971
rect 3063 2971 3064 2972
rect 3068 2971 3069 2975
rect 3311 2975 3317 2976
rect 3311 2974 3312 2975
rect 3205 2972 3312 2974
rect 3063 2970 3069 2971
rect 3311 2971 3312 2972
rect 3316 2971 3317 2975
rect 3311 2970 3317 2971
rect 3470 2975 3476 2976
rect 3470 2971 3471 2975
rect 3475 2974 3476 2975
rect 3475 2972 3505 2974
rect 3574 2972 3580 2973
rect 3475 2971 3476 2972
rect 3470 2970 3476 2971
rect 1862 2967 1868 2968
rect 3574 2968 3575 2972
rect 3579 2968 3580 2972
rect 3574 2967 3580 2968
rect 2030 2959 2036 2960
rect 2030 2955 2031 2959
rect 2035 2955 2036 2959
rect 2030 2954 2036 2955
rect 2166 2959 2172 2960
rect 2166 2955 2167 2959
rect 2171 2955 2172 2959
rect 2166 2954 2172 2955
rect 2294 2959 2300 2960
rect 2294 2955 2295 2959
rect 2299 2955 2300 2959
rect 2294 2954 2300 2955
rect 2422 2959 2428 2960
rect 2422 2955 2423 2959
rect 2427 2955 2428 2959
rect 2422 2954 2428 2955
rect 2542 2959 2548 2960
rect 2542 2955 2543 2959
rect 2547 2955 2548 2959
rect 2542 2954 2548 2955
rect 2670 2959 2676 2960
rect 2670 2955 2671 2959
rect 2675 2955 2676 2959
rect 2670 2954 2676 2955
rect 2814 2959 2820 2960
rect 2814 2955 2815 2959
rect 2819 2955 2820 2959
rect 2814 2954 2820 2955
rect 2974 2959 2980 2960
rect 2974 2955 2975 2959
rect 2979 2955 2980 2959
rect 2974 2954 2980 2955
rect 3150 2959 3156 2960
rect 3150 2955 3151 2959
rect 3155 2955 3156 2959
rect 3150 2954 3156 2955
rect 3326 2959 3332 2960
rect 3326 2955 3327 2959
rect 3331 2955 3332 2959
rect 3326 2954 3332 2955
rect 3486 2959 3492 2960
rect 3486 2955 3487 2959
rect 3491 2955 3492 2959
rect 3486 2954 3492 2955
rect 494 2951 500 2952
rect 494 2947 495 2951
rect 499 2947 500 2951
rect 494 2946 500 2947
rect 638 2951 644 2952
rect 638 2947 639 2951
rect 643 2947 644 2951
rect 638 2946 644 2947
rect 782 2951 788 2952
rect 782 2947 783 2951
rect 787 2947 788 2951
rect 782 2946 788 2947
rect 918 2951 924 2952
rect 918 2947 919 2951
rect 923 2947 924 2951
rect 918 2946 924 2947
rect 1054 2951 1060 2952
rect 1054 2947 1055 2951
rect 1059 2947 1060 2951
rect 1054 2946 1060 2947
rect 1182 2951 1188 2952
rect 1182 2947 1183 2951
rect 1187 2947 1188 2951
rect 1182 2946 1188 2947
rect 1302 2951 1308 2952
rect 1302 2947 1303 2951
rect 1307 2947 1308 2951
rect 1302 2946 1308 2947
rect 1414 2951 1420 2952
rect 1414 2947 1415 2951
rect 1419 2947 1420 2951
rect 1414 2946 1420 2947
rect 1526 2951 1532 2952
rect 1526 2947 1527 2951
rect 1531 2947 1532 2951
rect 1526 2946 1532 2947
rect 1638 2951 1644 2952
rect 1638 2947 1639 2951
rect 1643 2947 1644 2951
rect 1638 2946 1644 2947
rect 1726 2951 1732 2952
rect 1726 2947 1727 2951
rect 1731 2947 1732 2951
rect 1726 2946 1732 2947
rect 2023 2947 2029 2948
rect 871 2943 877 2944
rect 110 2941 116 2942
rect 110 2937 111 2941
rect 115 2937 116 2941
rect 871 2939 872 2943
rect 876 2942 877 2943
rect 1594 2943 1600 2944
rect 1594 2942 1595 2943
rect 876 2940 937 2942
rect 1585 2940 1595 2942
rect 876 2939 877 2940
rect 871 2938 877 2939
rect 1594 2939 1595 2940
rect 1599 2939 1600 2943
rect 2023 2943 2024 2947
rect 2028 2946 2029 2947
rect 2031 2947 2037 2948
rect 2031 2946 2032 2947
rect 2028 2944 2032 2946
rect 2028 2943 2029 2944
rect 2023 2942 2029 2943
rect 2031 2943 2032 2944
rect 2036 2943 2037 2947
rect 2031 2942 2037 2943
rect 2151 2947 2157 2948
rect 2151 2943 2152 2947
rect 2156 2946 2157 2947
rect 2159 2947 2165 2948
rect 2159 2946 2160 2947
rect 2156 2944 2160 2946
rect 2156 2943 2157 2944
rect 2151 2942 2157 2943
rect 2159 2943 2160 2944
rect 2164 2943 2165 2947
rect 2159 2942 2165 2943
rect 2279 2947 2285 2948
rect 2279 2943 2280 2947
rect 2284 2946 2285 2947
rect 2287 2947 2293 2948
rect 2287 2946 2288 2947
rect 2284 2944 2288 2946
rect 2284 2943 2285 2944
rect 2279 2942 2285 2943
rect 2287 2943 2288 2944
rect 2292 2943 2293 2947
rect 2287 2942 2293 2943
rect 2415 2947 2421 2948
rect 2415 2943 2416 2947
rect 2420 2946 2421 2947
rect 2430 2947 2436 2948
rect 2430 2946 2431 2947
rect 2420 2944 2431 2946
rect 2420 2943 2421 2944
rect 2415 2942 2421 2943
rect 2430 2943 2431 2944
rect 2435 2943 2436 2947
rect 2430 2942 2436 2943
rect 2527 2947 2533 2948
rect 2527 2943 2528 2947
rect 2532 2946 2533 2947
rect 2535 2947 2541 2948
rect 2535 2946 2536 2947
rect 2532 2944 2536 2946
rect 2532 2943 2533 2944
rect 2527 2942 2533 2943
rect 2535 2943 2536 2944
rect 2540 2943 2541 2947
rect 2535 2942 2541 2943
rect 2655 2947 2661 2948
rect 2655 2943 2656 2947
rect 2660 2946 2661 2947
rect 2663 2947 2669 2948
rect 2663 2946 2664 2947
rect 2660 2944 2664 2946
rect 2660 2943 2661 2944
rect 2655 2942 2661 2943
rect 2663 2943 2664 2944
rect 2668 2943 2669 2947
rect 2663 2942 2669 2943
rect 2799 2947 2805 2948
rect 2799 2943 2800 2947
rect 2804 2946 2805 2947
rect 2807 2947 2813 2948
rect 2807 2946 2808 2947
rect 2804 2944 2808 2946
rect 2804 2943 2805 2944
rect 2799 2942 2805 2943
rect 2807 2943 2808 2944
rect 2812 2943 2813 2947
rect 2807 2942 2813 2943
rect 2959 2947 2965 2948
rect 2959 2943 2960 2947
rect 2964 2946 2965 2947
rect 2967 2947 2973 2948
rect 2967 2946 2968 2947
rect 2964 2944 2968 2946
rect 2964 2943 2965 2944
rect 2959 2942 2965 2943
rect 2967 2943 2968 2944
rect 2972 2943 2973 2947
rect 2967 2942 2973 2943
rect 3063 2947 3069 2948
rect 3063 2943 3064 2947
rect 3068 2946 3069 2947
rect 3143 2947 3149 2948
rect 3143 2946 3144 2947
rect 3068 2944 3144 2946
rect 3068 2943 3069 2944
rect 3063 2942 3069 2943
rect 3143 2943 3144 2944
rect 3148 2943 3149 2947
rect 3143 2942 3149 2943
rect 3311 2947 3317 2948
rect 3311 2943 3312 2947
rect 3316 2946 3317 2947
rect 3319 2947 3325 2948
rect 3319 2946 3320 2947
rect 3316 2944 3320 2946
rect 3316 2943 3317 2944
rect 3311 2942 3317 2943
rect 3319 2943 3320 2944
rect 3324 2943 3325 2947
rect 3319 2942 3325 2943
rect 3471 2947 3477 2948
rect 3471 2943 3472 2947
rect 3476 2946 3477 2947
rect 3479 2947 3485 2948
rect 3479 2946 3480 2947
rect 3476 2944 3480 2946
rect 3476 2943 3477 2944
rect 3471 2942 3477 2943
rect 3479 2943 3480 2944
rect 3484 2943 3485 2947
rect 3479 2942 3485 2943
rect 1594 2938 1600 2939
rect 1822 2941 1828 2942
rect 110 2936 116 2937
rect 1822 2937 1823 2941
rect 1827 2937 1828 2941
rect 1822 2936 1828 2937
rect 1816 2928 1834 2930
rect 630 2927 636 2928
rect 630 2926 631 2927
rect 110 2924 116 2925
rect 557 2924 631 2926
rect 110 2920 111 2924
rect 115 2920 116 2924
rect 630 2923 631 2924
rect 635 2923 636 2927
rect 775 2927 781 2928
rect 775 2926 776 2927
rect 701 2924 776 2926
rect 630 2922 636 2923
rect 775 2923 776 2924
rect 780 2923 781 2927
rect 911 2927 917 2928
rect 911 2926 912 2927
rect 845 2924 912 2926
rect 775 2922 781 2923
rect 911 2923 912 2924
rect 916 2923 917 2927
rect 1175 2927 1181 2928
rect 1175 2926 1176 2927
rect 1117 2924 1176 2926
rect 911 2922 917 2923
rect 1175 2923 1176 2924
rect 1180 2923 1181 2927
rect 1295 2927 1301 2928
rect 1295 2926 1296 2927
rect 1245 2924 1296 2926
rect 1175 2922 1181 2923
rect 1295 2923 1296 2924
rect 1300 2923 1301 2927
rect 1407 2927 1413 2928
rect 1407 2926 1408 2927
rect 1365 2924 1408 2926
rect 1295 2922 1301 2923
rect 1407 2923 1408 2924
rect 1412 2923 1413 2927
rect 1519 2927 1525 2928
rect 1519 2926 1520 2927
rect 1477 2924 1520 2926
rect 1407 2922 1413 2923
rect 1519 2923 1520 2924
rect 1524 2923 1525 2927
rect 1719 2927 1725 2928
rect 1719 2926 1720 2927
rect 1701 2924 1720 2926
rect 1519 2922 1525 2923
rect 1719 2923 1720 2924
rect 1724 2923 1725 2927
rect 1816 2926 1818 2928
rect 1789 2924 1818 2926
rect 1832 2926 1834 2928
rect 1887 2927 1893 2928
rect 1887 2926 1888 2927
rect 1822 2924 1828 2925
rect 1832 2924 1888 2926
rect 1719 2922 1725 2923
rect 110 2919 116 2920
rect 1822 2920 1823 2924
rect 1827 2920 1828 2924
rect 1887 2923 1888 2924
rect 1892 2923 1893 2927
rect 1887 2922 1893 2923
rect 2167 2927 2173 2928
rect 2167 2923 2168 2927
rect 2172 2926 2173 2927
rect 2318 2927 2324 2928
rect 2318 2926 2319 2927
rect 2172 2924 2319 2926
rect 2172 2923 2173 2924
rect 2167 2922 2173 2923
rect 2318 2923 2319 2924
rect 2323 2923 2324 2927
rect 2318 2922 2324 2923
rect 2487 2927 2493 2928
rect 2487 2923 2488 2927
rect 2492 2926 2493 2927
rect 2562 2927 2568 2928
rect 2562 2926 2563 2927
rect 2492 2924 2563 2926
rect 2492 2923 2493 2924
rect 2487 2922 2493 2923
rect 2562 2923 2563 2924
rect 2567 2923 2568 2927
rect 2562 2922 2568 2923
rect 2663 2927 2669 2928
rect 2663 2923 2664 2927
rect 2668 2926 2669 2927
rect 2815 2927 2821 2928
rect 2815 2926 2816 2927
rect 2668 2924 2816 2926
rect 2668 2923 2669 2924
rect 2663 2922 2669 2923
rect 2815 2923 2816 2924
rect 2820 2923 2821 2927
rect 2815 2922 2821 2923
rect 3151 2927 3157 2928
rect 3151 2923 3152 2927
rect 3156 2926 3157 2927
rect 3159 2927 3165 2928
rect 3159 2926 3160 2927
rect 3156 2924 3160 2926
rect 3156 2923 3157 2924
rect 3151 2922 3157 2923
rect 3159 2923 3160 2924
rect 3164 2923 3165 2927
rect 3159 2922 3165 2923
rect 3470 2927 3476 2928
rect 3470 2923 3471 2927
rect 3475 2926 3476 2927
rect 3479 2927 3485 2928
rect 3479 2926 3480 2927
rect 3475 2924 3480 2926
rect 3475 2923 3476 2924
rect 3470 2922 3476 2923
rect 3479 2923 3480 2924
rect 3484 2923 3485 2927
rect 3479 2922 3485 2923
rect 1822 2919 1828 2920
rect 1894 2917 1900 2918
rect 1894 2913 1895 2917
rect 1899 2913 1900 2917
rect 1894 2912 1900 2913
rect 2174 2917 2180 2918
rect 2174 2913 2175 2917
rect 2179 2913 2180 2917
rect 2174 2912 2180 2913
rect 2494 2917 2500 2918
rect 2494 2913 2495 2917
rect 2499 2913 2500 2917
rect 2494 2912 2500 2913
rect 2822 2917 2828 2918
rect 2822 2913 2823 2917
rect 2827 2913 2828 2917
rect 2822 2912 2828 2913
rect 3166 2917 3172 2918
rect 3166 2913 3167 2917
rect 3171 2913 3172 2917
rect 3166 2912 3172 2913
rect 3486 2917 3492 2918
rect 3486 2913 3487 2917
rect 3491 2913 3492 2917
rect 3486 2912 3492 2913
rect 502 2911 508 2912
rect 502 2907 503 2911
rect 507 2907 508 2911
rect 502 2906 508 2907
rect 646 2911 652 2912
rect 646 2907 647 2911
rect 651 2907 652 2911
rect 646 2906 652 2907
rect 790 2911 796 2912
rect 790 2907 791 2911
rect 795 2907 796 2911
rect 790 2906 796 2907
rect 926 2911 932 2912
rect 926 2907 927 2911
rect 931 2907 932 2911
rect 926 2906 932 2907
rect 1062 2911 1068 2912
rect 1062 2907 1063 2911
rect 1067 2907 1068 2911
rect 1062 2906 1068 2907
rect 1190 2911 1196 2912
rect 1190 2907 1191 2911
rect 1195 2907 1196 2911
rect 1190 2906 1196 2907
rect 1310 2911 1316 2912
rect 1310 2907 1311 2911
rect 1315 2907 1316 2911
rect 1310 2906 1316 2907
rect 1422 2911 1428 2912
rect 1422 2907 1423 2911
rect 1427 2907 1428 2911
rect 1422 2906 1428 2907
rect 1534 2911 1540 2912
rect 1534 2907 1535 2911
rect 1539 2907 1540 2911
rect 1534 2906 1540 2907
rect 1646 2911 1652 2912
rect 1646 2907 1647 2911
rect 1651 2907 1652 2911
rect 1646 2906 1652 2907
rect 1734 2911 1740 2912
rect 1734 2907 1735 2911
rect 1739 2907 1740 2911
rect 1734 2906 1740 2907
rect 1862 2904 1868 2905
rect 1862 2900 1863 2904
rect 1867 2900 1868 2904
rect 3574 2904 3580 2905
rect 3574 2900 3575 2904
rect 3579 2900 3580 2904
rect 495 2899 501 2900
rect 495 2895 496 2899
rect 500 2898 501 2899
rect 510 2899 516 2900
rect 510 2898 511 2899
rect 500 2896 511 2898
rect 500 2895 501 2896
rect 495 2894 501 2895
rect 510 2895 511 2896
rect 515 2895 516 2899
rect 510 2894 516 2895
rect 630 2899 636 2900
rect 630 2895 631 2899
rect 635 2898 636 2899
rect 639 2899 645 2900
rect 639 2898 640 2899
rect 635 2896 640 2898
rect 635 2895 636 2896
rect 630 2894 636 2895
rect 639 2895 640 2896
rect 644 2895 645 2899
rect 639 2894 645 2895
rect 775 2899 781 2900
rect 775 2895 776 2899
rect 780 2898 781 2899
rect 783 2899 789 2900
rect 783 2898 784 2899
rect 780 2896 784 2898
rect 780 2895 781 2896
rect 775 2894 781 2895
rect 783 2895 784 2896
rect 788 2895 789 2899
rect 783 2894 789 2895
rect 911 2899 917 2900
rect 911 2895 912 2899
rect 916 2898 917 2899
rect 919 2899 925 2900
rect 919 2898 920 2899
rect 916 2896 920 2898
rect 916 2895 917 2896
rect 911 2894 917 2895
rect 919 2895 920 2896
rect 924 2895 925 2899
rect 919 2894 925 2895
rect 1055 2899 1061 2900
rect 1055 2895 1056 2899
rect 1060 2898 1061 2899
rect 1166 2899 1172 2900
rect 1166 2898 1167 2899
rect 1060 2896 1167 2898
rect 1060 2895 1061 2896
rect 1055 2894 1061 2895
rect 1166 2895 1167 2896
rect 1171 2895 1172 2899
rect 1166 2894 1172 2895
rect 1175 2899 1181 2900
rect 1175 2895 1176 2899
rect 1180 2898 1181 2899
rect 1183 2899 1189 2900
rect 1183 2898 1184 2899
rect 1180 2896 1184 2898
rect 1180 2895 1181 2896
rect 1175 2894 1181 2895
rect 1183 2895 1184 2896
rect 1188 2895 1189 2899
rect 1183 2894 1189 2895
rect 1295 2899 1301 2900
rect 1295 2895 1296 2899
rect 1300 2898 1301 2899
rect 1303 2899 1309 2900
rect 1303 2898 1304 2899
rect 1300 2896 1304 2898
rect 1300 2895 1301 2896
rect 1295 2894 1301 2895
rect 1303 2895 1304 2896
rect 1308 2895 1309 2899
rect 1303 2894 1309 2895
rect 1407 2899 1413 2900
rect 1407 2895 1408 2899
rect 1412 2898 1413 2899
rect 1415 2899 1421 2900
rect 1415 2898 1416 2899
rect 1412 2896 1416 2898
rect 1412 2895 1413 2896
rect 1407 2894 1413 2895
rect 1415 2895 1416 2896
rect 1420 2895 1421 2899
rect 1415 2894 1421 2895
rect 1519 2899 1525 2900
rect 1519 2895 1520 2899
rect 1524 2898 1525 2899
rect 1527 2899 1533 2900
rect 1527 2898 1528 2899
rect 1524 2896 1528 2898
rect 1524 2895 1525 2896
rect 1519 2894 1525 2895
rect 1527 2895 1528 2896
rect 1532 2895 1533 2899
rect 1527 2894 1533 2895
rect 1639 2899 1645 2900
rect 1639 2895 1640 2899
rect 1644 2898 1645 2899
rect 1690 2899 1696 2900
rect 1690 2898 1691 2899
rect 1644 2896 1691 2898
rect 1644 2895 1645 2896
rect 1639 2894 1645 2895
rect 1690 2895 1691 2896
rect 1695 2895 1696 2899
rect 1690 2894 1696 2895
rect 1719 2899 1725 2900
rect 1719 2895 1720 2899
rect 1724 2898 1725 2899
rect 1727 2899 1733 2900
rect 1862 2899 1868 2900
rect 2031 2899 2037 2900
rect 1727 2898 1728 2899
rect 1724 2896 1728 2898
rect 1724 2895 1725 2896
rect 1719 2894 1725 2895
rect 1727 2895 1728 2896
rect 1732 2895 1733 2899
rect 1727 2894 1733 2895
rect 2031 2895 2032 2899
rect 2036 2898 2037 2899
rect 2318 2899 2324 2900
rect 2036 2896 2193 2898
rect 2036 2895 2037 2896
rect 2031 2894 2037 2895
rect 2318 2895 2319 2899
rect 2323 2898 2324 2899
rect 2562 2899 2568 2900
rect 3574 2899 3580 2900
rect 2323 2896 2513 2898
rect 2323 2895 2324 2896
rect 2318 2894 2324 2895
rect 2562 2895 2563 2899
rect 2567 2898 2568 2899
rect 2567 2896 2841 2898
rect 2567 2895 2568 2896
rect 2562 2894 2568 2895
rect 1862 2887 1868 2888
rect 319 2883 325 2884
rect 319 2879 320 2883
rect 324 2882 325 2883
rect 394 2883 400 2884
rect 394 2882 395 2883
rect 324 2880 395 2882
rect 324 2879 325 2880
rect 319 2878 325 2879
rect 394 2879 395 2880
rect 399 2879 400 2883
rect 394 2878 400 2879
rect 447 2883 453 2884
rect 447 2879 448 2883
rect 452 2882 453 2883
rect 522 2883 528 2884
rect 522 2882 523 2883
rect 452 2880 523 2882
rect 452 2879 453 2880
rect 447 2878 453 2879
rect 522 2879 523 2880
rect 527 2879 528 2883
rect 522 2878 528 2879
rect 583 2883 589 2884
rect 583 2879 584 2883
rect 588 2882 589 2883
rect 670 2883 676 2884
rect 670 2882 671 2883
rect 588 2880 671 2882
rect 588 2879 589 2880
rect 583 2878 589 2879
rect 670 2879 671 2880
rect 675 2879 676 2883
rect 670 2878 676 2879
rect 719 2883 725 2884
rect 719 2879 720 2883
rect 724 2882 725 2883
rect 798 2883 804 2884
rect 798 2882 799 2883
rect 724 2880 799 2882
rect 724 2879 725 2880
rect 719 2878 725 2879
rect 798 2879 799 2880
rect 803 2879 804 2883
rect 798 2878 804 2879
rect 863 2883 869 2884
rect 863 2879 864 2883
rect 868 2882 869 2883
rect 871 2883 877 2884
rect 871 2882 872 2883
rect 868 2880 872 2882
rect 868 2879 869 2880
rect 863 2878 869 2879
rect 871 2879 872 2880
rect 876 2879 877 2883
rect 871 2878 877 2879
rect 999 2883 1005 2884
rect 999 2879 1000 2883
rect 1004 2882 1005 2883
rect 1014 2883 1020 2884
rect 1014 2882 1015 2883
rect 1004 2880 1015 2882
rect 1004 2879 1005 2880
rect 999 2878 1005 2879
rect 1014 2879 1015 2880
rect 1019 2879 1020 2883
rect 1014 2878 1020 2879
rect 1071 2883 1077 2884
rect 1071 2879 1072 2883
rect 1076 2882 1077 2883
rect 1135 2883 1141 2884
rect 1135 2882 1136 2883
rect 1076 2880 1136 2882
rect 1076 2879 1077 2880
rect 1071 2878 1077 2879
rect 1135 2879 1136 2880
rect 1140 2879 1141 2883
rect 1135 2878 1141 2879
rect 1207 2883 1213 2884
rect 1207 2879 1208 2883
rect 1212 2882 1213 2883
rect 1271 2883 1277 2884
rect 1271 2882 1272 2883
rect 1212 2880 1272 2882
rect 1212 2879 1213 2880
rect 1207 2878 1213 2879
rect 1271 2879 1272 2880
rect 1276 2879 1277 2883
rect 1271 2878 1277 2879
rect 1343 2883 1349 2884
rect 1343 2879 1344 2883
rect 1348 2882 1349 2883
rect 1407 2883 1413 2884
rect 1407 2882 1408 2883
rect 1348 2880 1408 2882
rect 1348 2879 1349 2880
rect 1343 2878 1349 2879
rect 1407 2879 1408 2880
rect 1412 2879 1413 2883
rect 1407 2878 1413 2879
rect 1502 2883 1508 2884
rect 1502 2879 1503 2883
rect 1507 2882 1508 2883
rect 1543 2883 1549 2884
rect 1543 2882 1544 2883
rect 1507 2880 1544 2882
rect 1507 2879 1508 2880
rect 1502 2878 1508 2879
rect 1543 2879 1544 2880
rect 1548 2879 1549 2883
rect 1862 2883 1863 2887
rect 1867 2883 1868 2887
rect 1862 2882 1868 2883
rect 1879 2887 1885 2888
rect 1879 2883 1880 2887
rect 1884 2886 1885 2887
rect 3070 2887 3076 2888
rect 1884 2884 1905 2886
rect 1884 2883 1885 2884
rect 1879 2882 1885 2883
rect 3070 2883 3071 2887
rect 3075 2886 3076 2887
rect 3471 2887 3477 2888
rect 3075 2884 3177 2886
rect 3075 2883 3076 2884
rect 3070 2882 3076 2883
rect 3471 2883 3472 2887
rect 3476 2886 3477 2887
rect 3574 2887 3580 2888
rect 3476 2884 3497 2886
rect 3476 2883 3477 2884
rect 3471 2882 3477 2883
rect 3574 2883 3575 2887
rect 3579 2883 3580 2887
rect 3574 2882 3580 2883
rect 1543 2878 1549 2879
rect 1886 2877 1892 2878
rect 326 2873 332 2874
rect 326 2869 327 2873
rect 331 2869 332 2873
rect 326 2868 332 2869
rect 454 2873 460 2874
rect 454 2869 455 2873
rect 459 2869 460 2873
rect 454 2868 460 2869
rect 590 2873 596 2874
rect 590 2869 591 2873
rect 595 2869 596 2873
rect 590 2868 596 2869
rect 726 2873 732 2874
rect 726 2869 727 2873
rect 731 2869 732 2873
rect 726 2868 732 2869
rect 870 2873 876 2874
rect 870 2869 871 2873
rect 875 2869 876 2873
rect 870 2868 876 2869
rect 1006 2873 1012 2874
rect 1006 2869 1007 2873
rect 1011 2869 1012 2873
rect 1006 2868 1012 2869
rect 1142 2873 1148 2874
rect 1142 2869 1143 2873
rect 1147 2869 1148 2873
rect 1142 2868 1148 2869
rect 1278 2873 1284 2874
rect 1278 2869 1279 2873
rect 1283 2869 1284 2873
rect 1278 2868 1284 2869
rect 1414 2873 1420 2874
rect 1414 2869 1415 2873
rect 1419 2869 1420 2873
rect 1414 2868 1420 2869
rect 1550 2873 1556 2874
rect 1550 2869 1551 2873
rect 1555 2869 1556 2873
rect 1886 2873 1887 2877
rect 1891 2873 1892 2877
rect 1886 2872 1892 2873
rect 2166 2877 2172 2878
rect 2166 2873 2167 2877
rect 2171 2873 2172 2877
rect 2166 2872 2172 2873
rect 2486 2877 2492 2878
rect 2486 2873 2487 2877
rect 2491 2873 2492 2877
rect 2486 2872 2492 2873
rect 2814 2877 2820 2878
rect 2814 2873 2815 2877
rect 2819 2873 2820 2877
rect 2814 2872 2820 2873
rect 3158 2877 3164 2878
rect 3158 2873 3159 2877
rect 3163 2873 3164 2877
rect 3158 2872 3164 2873
rect 3478 2877 3484 2878
rect 3478 2873 3479 2877
rect 3483 2873 3484 2877
rect 3478 2872 3484 2873
rect 1550 2868 1556 2869
rect 2686 2863 2692 2864
rect 110 2860 116 2861
rect 1822 2860 1828 2861
rect 110 2856 111 2860
rect 115 2856 116 2860
rect 1071 2859 1077 2860
rect 1071 2858 1072 2859
rect 1061 2856 1072 2858
rect 110 2855 116 2856
rect 394 2855 400 2856
rect 394 2851 395 2855
rect 399 2854 400 2855
rect 522 2855 528 2856
rect 399 2852 473 2854
rect 399 2851 400 2852
rect 394 2850 400 2851
rect 522 2851 523 2855
rect 527 2854 528 2855
rect 670 2855 676 2856
rect 527 2852 609 2854
rect 527 2851 528 2852
rect 522 2850 528 2851
rect 670 2851 671 2855
rect 675 2854 676 2855
rect 798 2855 804 2856
rect 675 2852 745 2854
rect 675 2851 676 2852
rect 670 2850 676 2851
rect 798 2851 799 2855
rect 803 2854 804 2855
rect 1071 2855 1072 2856
rect 1076 2855 1077 2859
rect 1207 2859 1213 2860
rect 1207 2858 1208 2859
rect 1197 2856 1208 2858
rect 1071 2854 1077 2855
rect 1207 2855 1208 2856
rect 1212 2855 1213 2859
rect 1343 2859 1349 2860
rect 1343 2858 1344 2859
rect 1333 2856 1344 2858
rect 1207 2854 1213 2855
rect 1343 2855 1344 2856
rect 1348 2855 1349 2859
rect 1502 2859 1508 2860
rect 1502 2858 1503 2859
rect 1469 2856 1503 2858
rect 1343 2854 1349 2855
rect 1502 2855 1503 2856
rect 1507 2855 1508 2859
rect 1822 2856 1823 2860
rect 1827 2856 1828 2860
rect 2686 2859 2687 2863
rect 2691 2862 2692 2863
rect 2691 2860 3006 2862
rect 2691 2859 2692 2860
rect 2686 2858 2692 2859
rect 1502 2854 1508 2855
rect 1510 2855 1516 2856
rect 1822 2855 1828 2856
rect 1886 2855 1892 2856
rect 803 2852 889 2854
rect 803 2851 804 2852
rect 798 2850 804 2851
rect 1510 2851 1511 2855
rect 1515 2854 1516 2855
rect 1515 2852 1569 2854
rect 1515 2851 1516 2852
rect 1510 2850 1516 2851
rect 1886 2851 1887 2855
rect 1891 2851 1892 2855
rect 1886 2850 1892 2851
rect 2022 2855 2028 2856
rect 2022 2851 2023 2855
rect 2027 2851 2028 2855
rect 2022 2850 2028 2851
rect 2190 2855 2196 2856
rect 2190 2851 2191 2855
rect 2195 2851 2196 2855
rect 2190 2850 2196 2851
rect 2358 2855 2364 2856
rect 2358 2851 2359 2855
rect 2363 2851 2364 2855
rect 2358 2850 2364 2851
rect 2518 2855 2524 2856
rect 2518 2851 2519 2855
rect 2523 2851 2524 2855
rect 2518 2850 2524 2851
rect 2670 2855 2676 2856
rect 2670 2851 2671 2855
rect 2675 2851 2676 2855
rect 2670 2850 2676 2851
rect 2806 2855 2812 2856
rect 2806 2851 2807 2855
rect 2811 2851 2812 2855
rect 2806 2850 2812 2851
rect 2934 2855 2940 2856
rect 2934 2851 2935 2855
rect 2939 2851 2940 2855
rect 2934 2850 2940 2851
rect 2663 2847 2669 2848
rect 2663 2846 2664 2847
rect 1862 2845 1868 2846
rect 110 2843 116 2844
rect 110 2839 111 2843
rect 115 2839 116 2843
rect 415 2843 421 2844
rect 415 2842 416 2843
rect 377 2840 416 2842
rect 110 2838 116 2839
rect 415 2839 416 2840
rect 420 2839 421 2843
rect 415 2838 421 2839
rect 1822 2843 1828 2844
rect 1822 2839 1823 2843
rect 1827 2839 1828 2843
rect 1862 2841 1863 2845
rect 1867 2841 1868 2845
rect 2577 2844 2664 2846
rect 2663 2843 2664 2844
rect 2668 2843 2669 2847
rect 3004 2846 3006 2860
rect 3054 2855 3060 2856
rect 3054 2851 3055 2855
rect 3059 2851 3060 2855
rect 3054 2850 3060 2851
rect 3166 2855 3172 2856
rect 3166 2851 3167 2855
rect 3171 2851 3172 2855
rect 3166 2850 3172 2851
rect 3278 2855 3284 2856
rect 3278 2851 3279 2855
rect 3283 2851 3284 2855
rect 3278 2850 3284 2851
rect 3390 2855 3396 2856
rect 3390 2851 3391 2855
rect 3395 2851 3396 2855
rect 3390 2850 3396 2851
rect 3478 2855 3484 2856
rect 3478 2851 3479 2855
rect 3483 2851 3484 2855
rect 3478 2850 3484 2851
rect 3151 2847 3157 2848
rect 3004 2844 3073 2846
rect 2663 2842 2669 2843
rect 3151 2843 3152 2847
rect 3156 2846 3157 2847
rect 3156 2844 3185 2846
rect 3574 2845 3580 2846
rect 3156 2843 3157 2844
rect 3151 2842 3157 2843
rect 1862 2840 1868 2841
rect 3574 2841 3575 2845
rect 3579 2841 3580 2845
rect 3574 2840 3580 2841
rect 1822 2838 1828 2839
rect 318 2833 324 2834
rect 318 2829 319 2833
rect 323 2829 324 2833
rect 318 2828 324 2829
rect 446 2833 452 2834
rect 446 2829 447 2833
rect 451 2829 452 2833
rect 446 2828 452 2829
rect 582 2833 588 2834
rect 582 2829 583 2833
rect 587 2829 588 2833
rect 582 2828 588 2829
rect 718 2833 724 2834
rect 718 2829 719 2833
rect 723 2829 724 2833
rect 718 2828 724 2829
rect 862 2833 868 2834
rect 862 2829 863 2833
rect 867 2829 868 2833
rect 862 2828 868 2829
rect 998 2833 1004 2834
rect 998 2829 999 2833
rect 1003 2829 1004 2833
rect 998 2828 1004 2829
rect 1134 2833 1140 2834
rect 1134 2829 1135 2833
rect 1139 2829 1140 2833
rect 1134 2828 1140 2829
rect 1270 2833 1276 2834
rect 1270 2829 1271 2833
rect 1275 2829 1276 2833
rect 1270 2828 1276 2829
rect 1406 2833 1412 2834
rect 1406 2829 1407 2833
rect 1411 2829 1412 2833
rect 1406 2828 1412 2829
rect 1542 2833 1548 2834
rect 1542 2829 1543 2833
rect 1547 2829 1548 2833
rect 2015 2831 2021 2832
rect 2015 2830 2016 2831
rect 1542 2828 1548 2829
rect 1862 2828 1868 2829
rect 1949 2828 2016 2830
rect 1862 2824 1863 2828
rect 1867 2824 1868 2828
rect 2015 2827 2016 2828
rect 2020 2827 2021 2831
rect 2090 2831 2096 2832
rect 2090 2830 2091 2831
rect 2085 2828 2091 2830
rect 2015 2826 2021 2827
rect 2090 2827 2091 2828
rect 2095 2827 2096 2831
rect 2351 2831 2357 2832
rect 2351 2830 2352 2831
rect 2253 2828 2352 2830
rect 2090 2826 2096 2827
rect 2351 2827 2352 2828
rect 2356 2827 2357 2831
rect 2511 2831 2517 2832
rect 2511 2830 2512 2831
rect 2421 2828 2512 2830
rect 2351 2826 2357 2827
rect 2511 2827 2512 2828
rect 2516 2827 2517 2831
rect 2799 2831 2805 2832
rect 2799 2830 2800 2831
rect 2733 2828 2800 2830
rect 2511 2826 2517 2827
rect 2799 2827 2800 2828
rect 2804 2827 2805 2831
rect 2927 2831 2933 2832
rect 2927 2830 2928 2831
rect 2869 2828 2928 2830
rect 2799 2826 2805 2827
rect 2927 2827 2928 2828
rect 2932 2827 2933 2831
rect 3047 2831 3053 2832
rect 3047 2830 3048 2831
rect 2997 2828 3048 2830
rect 2927 2826 2933 2827
rect 3047 2827 3048 2828
rect 3052 2827 3053 2831
rect 3047 2826 3053 2827
rect 3234 2831 3240 2832
rect 3234 2827 3235 2831
rect 3239 2830 3240 2831
rect 3346 2831 3352 2832
rect 3239 2828 3305 2830
rect 3239 2827 3240 2828
rect 3234 2826 3240 2827
rect 3346 2827 3347 2831
rect 3351 2830 3352 2831
rect 3470 2831 3476 2832
rect 3351 2828 3417 2830
rect 3351 2827 3352 2828
rect 3346 2826 3352 2827
rect 3470 2827 3471 2831
rect 3475 2830 3476 2831
rect 3475 2828 3505 2830
rect 3574 2828 3580 2829
rect 3475 2827 3476 2828
rect 3470 2826 3476 2827
rect 1862 2823 1868 2824
rect 3574 2824 3575 2828
rect 3579 2824 3580 2828
rect 3574 2823 3580 2824
rect 1894 2815 1900 2816
rect 1014 2811 1020 2812
rect 1014 2807 1015 2811
rect 1019 2810 1020 2811
rect 1894 2811 1895 2815
rect 1899 2811 1900 2815
rect 1894 2810 1900 2811
rect 2030 2815 2036 2816
rect 2030 2811 2031 2815
rect 2035 2811 2036 2815
rect 2030 2810 2036 2811
rect 2198 2815 2204 2816
rect 2198 2811 2199 2815
rect 2203 2811 2204 2815
rect 2198 2810 2204 2811
rect 2366 2815 2372 2816
rect 2366 2811 2367 2815
rect 2371 2811 2372 2815
rect 2366 2810 2372 2811
rect 2526 2815 2532 2816
rect 2526 2811 2527 2815
rect 2531 2811 2532 2815
rect 2526 2810 2532 2811
rect 2678 2815 2684 2816
rect 2678 2811 2679 2815
rect 2683 2811 2684 2815
rect 2678 2810 2684 2811
rect 2814 2815 2820 2816
rect 2814 2811 2815 2815
rect 2819 2811 2820 2815
rect 2814 2810 2820 2811
rect 2942 2815 2948 2816
rect 2942 2811 2943 2815
rect 2947 2811 2948 2815
rect 2942 2810 2948 2811
rect 3062 2815 3068 2816
rect 3062 2811 3063 2815
rect 3067 2811 3068 2815
rect 3062 2810 3068 2811
rect 3174 2815 3180 2816
rect 3174 2811 3175 2815
rect 3179 2811 3180 2815
rect 3174 2810 3180 2811
rect 3286 2815 3292 2816
rect 3286 2811 3287 2815
rect 3291 2811 3292 2815
rect 3286 2810 3292 2811
rect 3398 2815 3404 2816
rect 3398 2811 3399 2815
rect 3403 2811 3404 2815
rect 3398 2810 3404 2811
rect 3486 2815 3492 2816
rect 3486 2811 3487 2815
rect 3491 2811 3492 2815
rect 3486 2810 3492 2811
rect 1019 2808 1278 2810
rect 1019 2807 1020 2808
rect 1014 2806 1020 2807
rect 166 2803 172 2804
rect 166 2799 167 2803
rect 171 2799 172 2803
rect 166 2798 172 2799
rect 294 2803 300 2804
rect 294 2799 295 2803
rect 299 2799 300 2803
rect 294 2798 300 2799
rect 422 2803 428 2804
rect 422 2799 423 2803
rect 427 2799 428 2803
rect 422 2798 428 2799
rect 558 2803 564 2804
rect 558 2799 559 2803
rect 563 2799 564 2803
rect 558 2798 564 2799
rect 694 2803 700 2804
rect 694 2799 695 2803
rect 699 2799 700 2803
rect 694 2798 700 2799
rect 822 2803 828 2804
rect 822 2799 823 2803
rect 827 2799 828 2803
rect 822 2798 828 2799
rect 950 2803 956 2804
rect 950 2799 951 2803
rect 955 2799 956 2803
rect 950 2798 956 2799
rect 1078 2803 1084 2804
rect 1078 2799 1079 2803
rect 1083 2799 1084 2803
rect 1078 2798 1084 2799
rect 1206 2803 1212 2804
rect 1206 2799 1207 2803
rect 1211 2799 1212 2803
rect 1206 2798 1212 2799
rect 1276 2794 1278 2808
rect 1342 2803 1348 2804
rect 1342 2799 1343 2803
rect 1347 2799 1348 2803
rect 1342 2798 1348 2799
rect 1879 2803 1885 2804
rect 1879 2799 1880 2803
rect 1884 2802 1885 2803
rect 1887 2803 1893 2804
rect 1887 2802 1888 2803
rect 1884 2800 1888 2802
rect 1884 2799 1885 2800
rect 1879 2798 1885 2799
rect 1887 2799 1888 2800
rect 1892 2799 1893 2803
rect 1887 2798 1893 2799
rect 2015 2803 2021 2804
rect 2015 2799 2016 2803
rect 2020 2802 2021 2803
rect 2023 2803 2029 2804
rect 2023 2802 2024 2803
rect 2020 2800 2024 2802
rect 2020 2799 2021 2800
rect 2015 2798 2021 2799
rect 2023 2799 2024 2800
rect 2028 2799 2029 2803
rect 2023 2798 2029 2799
rect 2191 2803 2197 2804
rect 2191 2799 2192 2803
rect 2196 2802 2197 2803
rect 2199 2803 2205 2804
rect 2199 2802 2200 2803
rect 2196 2800 2200 2802
rect 2196 2799 2197 2800
rect 2191 2798 2197 2799
rect 2199 2799 2200 2800
rect 2204 2799 2205 2803
rect 2199 2798 2205 2799
rect 2351 2803 2357 2804
rect 2351 2799 2352 2803
rect 2356 2802 2357 2803
rect 2359 2803 2365 2804
rect 2359 2802 2360 2803
rect 2356 2800 2360 2802
rect 2356 2799 2357 2800
rect 2351 2798 2357 2799
rect 2359 2799 2360 2800
rect 2364 2799 2365 2803
rect 2359 2798 2365 2799
rect 2511 2803 2517 2804
rect 2511 2799 2512 2803
rect 2516 2802 2517 2803
rect 2519 2803 2525 2804
rect 2519 2802 2520 2803
rect 2516 2800 2520 2802
rect 2516 2799 2517 2800
rect 2511 2798 2517 2799
rect 2519 2799 2520 2800
rect 2524 2799 2525 2803
rect 2519 2798 2525 2799
rect 2671 2803 2677 2804
rect 2671 2799 2672 2803
rect 2676 2802 2677 2803
rect 2686 2803 2692 2804
rect 2686 2802 2687 2803
rect 2676 2800 2687 2802
rect 2676 2799 2677 2800
rect 2671 2798 2677 2799
rect 2686 2799 2687 2800
rect 2691 2799 2692 2803
rect 2686 2798 2692 2799
rect 2799 2803 2805 2804
rect 2799 2799 2800 2803
rect 2804 2802 2805 2803
rect 2807 2803 2813 2804
rect 2807 2802 2808 2803
rect 2804 2800 2808 2802
rect 2804 2799 2805 2800
rect 2799 2798 2805 2799
rect 2807 2799 2808 2800
rect 2812 2799 2813 2803
rect 2807 2798 2813 2799
rect 2927 2803 2933 2804
rect 2927 2799 2928 2803
rect 2932 2802 2933 2803
rect 2935 2803 2941 2804
rect 2935 2802 2936 2803
rect 2932 2800 2936 2802
rect 2932 2799 2933 2800
rect 2927 2798 2933 2799
rect 2935 2799 2936 2800
rect 2940 2799 2941 2803
rect 2935 2798 2941 2799
rect 3055 2803 3061 2804
rect 3055 2799 3056 2803
rect 3060 2802 3061 2803
rect 3070 2803 3076 2804
rect 3070 2802 3071 2803
rect 3060 2800 3071 2802
rect 3060 2799 3061 2800
rect 3055 2798 3061 2799
rect 3070 2799 3071 2800
rect 3075 2799 3076 2803
rect 3070 2798 3076 2799
rect 3167 2803 3173 2804
rect 3167 2799 3168 2803
rect 3172 2802 3173 2803
rect 3234 2803 3240 2804
rect 3234 2802 3235 2803
rect 3172 2800 3235 2802
rect 3172 2799 3173 2800
rect 3167 2798 3173 2799
rect 3234 2799 3235 2800
rect 3239 2799 3240 2803
rect 3234 2798 3240 2799
rect 3279 2803 3285 2804
rect 3279 2799 3280 2803
rect 3284 2802 3285 2803
rect 3346 2803 3352 2804
rect 3346 2802 3347 2803
rect 3284 2800 3347 2802
rect 3284 2799 3285 2800
rect 3279 2798 3285 2799
rect 3346 2799 3347 2800
rect 3351 2799 3352 2803
rect 3346 2798 3352 2799
rect 3391 2803 3397 2804
rect 3391 2799 3392 2803
rect 3396 2802 3397 2803
rect 3426 2803 3432 2804
rect 3426 2802 3427 2803
rect 3396 2800 3427 2802
rect 3396 2799 3397 2800
rect 3391 2798 3397 2799
rect 3426 2799 3427 2800
rect 3431 2799 3432 2803
rect 3426 2798 3432 2799
rect 3471 2803 3477 2804
rect 3471 2799 3472 2803
rect 3476 2802 3477 2803
rect 3479 2803 3485 2804
rect 3479 2802 3480 2803
rect 3476 2800 3480 2802
rect 3476 2799 3477 2800
rect 3471 2798 3477 2799
rect 3479 2799 3480 2800
rect 3484 2799 3485 2803
rect 3479 2798 3485 2799
rect 110 2793 116 2794
rect 110 2789 111 2793
rect 115 2789 116 2793
rect 1276 2792 1361 2794
rect 1822 2793 1828 2794
rect 110 2788 116 2789
rect 1822 2789 1823 2793
rect 1827 2789 1828 2793
rect 1822 2788 1828 2789
rect 1887 2791 1893 2792
rect 1887 2787 1888 2791
rect 1892 2790 1893 2791
rect 1967 2791 1973 2792
rect 1967 2790 1968 2791
rect 1892 2788 1968 2790
rect 1892 2787 1893 2788
rect 1887 2786 1893 2787
rect 1967 2787 1968 2788
rect 1972 2787 1973 2791
rect 1967 2786 1973 2787
rect 2055 2791 2061 2792
rect 2055 2787 2056 2791
rect 2060 2790 2061 2791
rect 2090 2791 2096 2792
rect 2090 2790 2091 2791
rect 2060 2788 2091 2790
rect 2060 2787 2061 2788
rect 2055 2786 2061 2787
rect 2090 2787 2091 2788
rect 2095 2787 2096 2791
rect 2090 2786 2096 2787
rect 2247 2791 2253 2792
rect 2247 2787 2248 2791
rect 2252 2790 2253 2791
rect 2338 2791 2344 2792
rect 2338 2790 2339 2791
rect 2252 2788 2339 2790
rect 2252 2787 2253 2788
rect 2247 2786 2253 2787
rect 2338 2787 2339 2788
rect 2343 2787 2344 2791
rect 2338 2786 2344 2787
rect 2431 2791 2437 2792
rect 2431 2787 2432 2791
rect 2436 2790 2437 2791
rect 2506 2791 2512 2792
rect 2506 2790 2507 2791
rect 2436 2788 2507 2790
rect 2436 2787 2437 2788
rect 2431 2786 2437 2787
rect 2506 2787 2507 2788
rect 2511 2787 2512 2791
rect 2506 2786 2512 2787
rect 2562 2791 2568 2792
rect 2562 2787 2563 2791
rect 2567 2790 2568 2791
rect 2607 2791 2613 2792
rect 2607 2790 2608 2791
rect 2567 2788 2608 2790
rect 2567 2787 2568 2788
rect 2562 2786 2568 2787
rect 2607 2787 2608 2788
rect 2612 2787 2613 2791
rect 2607 2786 2613 2787
rect 2775 2791 2781 2792
rect 2775 2787 2776 2791
rect 2780 2790 2781 2791
rect 2846 2791 2852 2792
rect 2846 2790 2847 2791
rect 2780 2788 2847 2790
rect 2780 2787 2781 2788
rect 2775 2786 2781 2787
rect 2846 2787 2847 2788
rect 2851 2787 2852 2791
rect 2846 2786 2852 2787
rect 2855 2791 2861 2792
rect 2855 2787 2856 2791
rect 2860 2790 2861 2791
rect 2927 2791 2933 2792
rect 2927 2790 2928 2791
rect 2860 2788 2928 2790
rect 2860 2787 2861 2788
rect 2855 2786 2861 2787
rect 2927 2787 2928 2788
rect 2932 2787 2933 2791
rect 2927 2786 2933 2787
rect 3047 2791 3053 2792
rect 3047 2787 3048 2791
rect 3052 2790 3053 2791
rect 3071 2791 3077 2792
rect 3071 2790 3072 2791
rect 3052 2788 3072 2790
rect 3052 2787 3053 2788
rect 3047 2786 3053 2787
rect 3071 2787 3072 2788
rect 3076 2787 3077 2791
rect 3071 2786 3077 2787
rect 3175 2791 3181 2792
rect 3175 2787 3176 2791
rect 3180 2790 3181 2791
rect 3215 2791 3221 2792
rect 3215 2790 3216 2791
rect 3180 2788 3216 2790
rect 3180 2787 3181 2788
rect 3175 2786 3181 2787
rect 3215 2787 3216 2788
rect 3220 2787 3221 2791
rect 3215 2786 3221 2787
rect 3359 2791 3365 2792
rect 3359 2787 3360 2791
rect 3364 2790 3365 2791
rect 3434 2791 3440 2792
rect 3434 2790 3435 2791
rect 3364 2788 3435 2790
rect 3364 2787 3365 2788
rect 3359 2786 3365 2787
rect 3434 2787 3435 2788
rect 3439 2787 3440 2791
rect 3434 2786 3440 2787
rect 3470 2791 3476 2792
rect 3470 2787 3471 2791
rect 3475 2790 3476 2791
rect 3479 2791 3485 2792
rect 3479 2790 3480 2791
rect 3475 2788 3480 2790
rect 3475 2787 3476 2788
rect 3470 2786 3476 2787
rect 3479 2787 3480 2788
rect 3484 2787 3485 2791
rect 3479 2786 3485 2787
rect 1894 2781 1900 2782
rect 287 2779 293 2780
rect 287 2778 288 2779
rect 110 2776 116 2777
rect 229 2776 288 2778
rect 110 2772 111 2776
rect 115 2772 116 2776
rect 287 2775 288 2776
rect 292 2775 293 2779
rect 362 2779 368 2780
rect 362 2778 363 2779
rect 357 2776 363 2778
rect 287 2774 293 2775
rect 362 2775 363 2776
rect 367 2775 368 2779
rect 551 2779 557 2780
rect 551 2778 552 2779
rect 485 2776 552 2778
rect 362 2774 368 2775
rect 551 2775 552 2776
rect 556 2775 557 2779
rect 626 2779 632 2780
rect 626 2778 627 2779
rect 621 2776 627 2778
rect 551 2774 557 2775
rect 626 2775 627 2776
rect 631 2775 632 2779
rect 626 2774 632 2775
rect 646 2779 652 2780
rect 646 2775 647 2779
rect 651 2778 652 2779
rect 943 2779 949 2780
rect 943 2778 944 2779
rect 651 2776 721 2778
rect 885 2776 944 2778
rect 651 2775 652 2776
rect 646 2774 652 2775
rect 943 2775 944 2776
rect 948 2775 949 2779
rect 1071 2779 1077 2780
rect 1071 2778 1072 2779
rect 1013 2776 1072 2778
rect 943 2774 949 2775
rect 1071 2775 1072 2776
rect 1076 2775 1077 2779
rect 1199 2779 1205 2780
rect 1199 2778 1200 2779
rect 1141 2776 1200 2778
rect 1071 2774 1077 2775
rect 1199 2775 1200 2776
rect 1204 2775 1205 2779
rect 1335 2779 1341 2780
rect 1335 2778 1336 2779
rect 1269 2776 1336 2778
rect 1199 2774 1205 2775
rect 1335 2775 1336 2776
rect 1340 2775 1341 2779
rect 1894 2777 1895 2781
rect 1899 2777 1900 2781
rect 1335 2774 1341 2775
rect 1822 2776 1828 2777
rect 1894 2776 1900 2777
rect 2062 2781 2068 2782
rect 2062 2777 2063 2781
rect 2067 2777 2068 2781
rect 2062 2776 2068 2777
rect 2254 2781 2260 2782
rect 2254 2777 2255 2781
rect 2259 2777 2260 2781
rect 2254 2776 2260 2777
rect 2438 2781 2444 2782
rect 2438 2777 2439 2781
rect 2443 2777 2444 2781
rect 2438 2776 2444 2777
rect 2614 2781 2620 2782
rect 2614 2777 2615 2781
rect 2619 2777 2620 2781
rect 2614 2776 2620 2777
rect 2782 2781 2788 2782
rect 2782 2777 2783 2781
rect 2787 2777 2788 2781
rect 2782 2776 2788 2777
rect 2934 2781 2940 2782
rect 2934 2777 2935 2781
rect 2939 2777 2940 2781
rect 2934 2776 2940 2777
rect 3078 2781 3084 2782
rect 3078 2777 3079 2781
rect 3083 2777 3084 2781
rect 3078 2776 3084 2777
rect 3222 2781 3228 2782
rect 3222 2777 3223 2781
rect 3227 2777 3228 2781
rect 3222 2776 3228 2777
rect 3366 2781 3372 2782
rect 3366 2777 3367 2781
rect 3371 2777 3372 2781
rect 3366 2776 3372 2777
rect 3486 2781 3492 2782
rect 3486 2777 3487 2781
rect 3491 2777 3492 2781
rect 3486 2776 3492 2777
rect 110 2771 116 2772
rect 1822 2772 1823 2776
rect 1827 2772 1828 2776
rect 1822 2771 1828 2772
rect 1862 2768 1868 2769
rect 3574 2768 3580 2769
rect 1862 2764 1863 2768
rect 1867 2764 1868 2768
rect 2855 2767 2861 2768
rect 2855 2766 2856 2767
rect 2837 2764 2856 2766
rect 174 2763 180 2764
rect 174 2759 175 2763
rect 179 2759 180 2763
rect 174 2758 180 2759
rect 302 2763 308 2764
rect 302 2759 303 2763
rect 307 2759 308 2763
rect 302 2758 308 2759
rect 430 2763 436 2764
rect 430 2759 431 2763
rect 435 2759 436 2763
rect 430 2758 436 2759
rect 566 2763 572 2764
rect 566 2759 567 2763
rect 571 2759 572 2763
rect 566 2758 572 2759
rect 702 2763 708 2764
rect 702 2759 703 2763
rect 707 2759 708 2763
rect 702 2758 708 2759
rect 830 2763 836 2764
rect 830 2759 831 2763
rect 835 2759 836 2763
rect 830 2758 836 2759
rect 958 2763 964 2764
rect 958 2759 959 2763
rect 963 2759 964 2763
rect 958 2758 964 2759
rect 1086 2763 1092 2764
rect 1086 2759 1087 2763
rect 1091 2759 1092 2763
rect 1086 2758 1092 2759
rect 1214 2763 1220 2764
rect 1214 2759 1215 2763
rect 1219 2759 1220 2763
rect 1214 2758 1220 2759
rect 1350 2763 1356 2764
rect 1862 2763 1868 2764
rect 1967 2763 1973 2764
rect 1350 2759 1351 2763
rect 1355 2759 1356 2763
rect 1350 2758 1356 2759
rect 1967 2759 1968 2763
rect 1972 2762 1973 2763
rect 2199 2763 2205 2764
rect 1972 2760 2081 2762
rect 1972 2759 1973 2760
rect 1967 2758 1973 2759
rect 2199 2759 2200 2763
rect 2204 2762 2205 2763
rect 2338 2763 2344 2764
rect 2204 2760 2273 2762
rect 2204 2759 2205 2760
rect 2199 2758 2205 2759
rect 2338 2759 2339 2763
rect 2343 2762 2344 2763
rect 2506 2763 2512 2764
rect 2343 2760 2457 2762
rect 2343 2759 2344 2760
rect 2338 2758 2344 2759
rect 2506 2759 2507 2763
rect 2511 2762 2512 2763
rect 2855 2763 2856 2764
rect 2860 2763 2861 2767
rect 3175 2767 3181 2768
rect 3175 2766 3176 2767
rect 3133 2764 3176 2766
rect 2855 2762 2861 2763
rect 3175 2763 3176 2764
rect 3180 2763 3181 2767
rect 3426 2767 3432 2768
rect 3426 2766 3427 2767
rect 3421 2764 3427 2766
rect 3175 2762 3181 2763
rect 3426 2763 3427 2764
rect 3431 2763 3432 2767
rect 3574 2764 3575 2768
rect 3579 2764 3580 2768
rect 3426 2762 3432 2763
rect 3434 2763 3440 2764
rect 3574 2763 3580 2764
rect 2511 2760 2633 2762
rect 2511 2759 2512 2760
rect 2506 2758 2512 2759
rect 3434 2759 3435 2763
rect 3439 2762 3440 2763
rect 3439 2760 3505 2762
rect 3439 2759 3440 2760
rect 3434 2758 3440 2759
rect 167 2751 173 2752
rect 167 2747 168 2751
rect 172 2750 173 2751
rect 182 2751 188 2752
rect 182 2750 183 2751
rect 172 2748 183 2750
rect 172 2747 173 2748
rect 167 2746 173 2747
rect 182 2747 183 2748
rect 187 2747 188 2751
rect 182 2746 188 2747
rect 287 2751 293 2752
rect 287 2747 288 2751
rect 292 2750 293 2751
rect 295 2751 301 2752
rect 295 2750 296 2751
rect 292 2748 296 2750
rect 292 2747 293 2748
rect 287 2746 293 2747
rect 295 2747 296 2748
rect 300 2747 301 2751
rect 295 2746 301 2747
rect 415 2751 421 2752
rect 415 2747 416 2751
rect 420 2750 421 2751
rect 423 2751 429 2752
rect 423 2750 424 2751
rect 420 2748 424 2750
rect 420 2747 421 2748
rect 415 2746 421 2747
rect 423 2747 424 2748
rect 428 2747 429 2751
rect 423 2746 429 2747
rect 551 2751 557 2752
rect 551 2747 552 2751
rect 556 2750 557 2751
rect 559 2751 565 2752
rect 559 2750 560 2751
rect 556 2748 560 2750
rect 556 2747 557 2748
rect 551 2746 557 2747
rect 559 2747 560 2748
rect 564 2747 565 2751
rect 559 2746 565 2747
rect 626 2751 632 2752
rect 626 2747 627 2751
rect 631 2750 632 2751
rect 695 2751 701 2752
rect 695 2750 696 2751
rect 631 2748 696 2750
rect 631 2747 632 2748
rect 626 2746 632 2747
rect 695 2747 696 2748
rect 700 2747 701 2751
rect 695 2746 701 2747
rect 823 2751 829 2752
rect 823 2747 824 2751
rect 828 2750 829 2751
rect 943 2751 949 2752
rect 828 2748 938 2750
rect 828 2747 829 2748
rect 823 2746 829 2747
rect 936 2742 938 2748
rect 943 2747 944 2751
rect 948 2750 949 2751
rect 951 2751 957 2752
rect 951 2750 952 2751
rect 948 2748 952 2750
rect 948 2747 949 2748
rect 943 2746 949 2747
rect 951 2747 952 2748
rect 956 2747 957 2751
rect 951 2746 957 2747
rect 1071 2751 1077 2752
rect 1071 2747 1072 2751
rect 1076 2750 1077 2751
rect 1079 2751 1085 2752
rect 1079 2750 1080 2751
rect 1076 2748 1080 2750
rect 1076 2747 1077 2748
rect 1071 2746 1077 2747
rect 1079 2747 1080 2748
rect 1084 2747 1085 2751
rect 1079 2746 1085 2747
rect 1199 2751 1205 2752
rect 1199 2747 1200 2751
rect 1204 2750 1205 2751
rect 1207 2751 1213 2752
rect 1207 2750 1208 2751
rect 1204 2748 1208 2750
rect 1204 2747 1205 2748
rect 1199 2746 1205 2747
rect 1207 2747 1208 2748
rect 1212 2747 1213 2751
rect 1207 2746 1213 2747
rect 1335 2751 1341 2752
rect 1335 2747 1336 2751
rect 1340 2750 1341 2751
rect 1343 2751 1349 2752
rect 1343 2750 1344 2751
rect 1340 2748 1344 2750
rect 1340 2747 1341 2748
rect 1335 2746 1341 2747
rect 1343 2747 1344 2748
rect 1348 2747 1349 2751
rect 1343 2746 1349 2747
rect 1862 2751 1868 2752
rect 1862 2747 1863 2751
rect 1867 2747 1868 2751
rect 2039 2751 2045 2752
rect 2039 2750 2040 2751
rect 1945 2748 2040 2750
rect 1862 2746 1868 2747
rect 2039 2747 2040 2748
rect 2044 2747 2045 2751
rect 2039 2746 2045 2747
rect 3183 2751 3189 2752
rect 3183 2747 3184 2751
rect 3188 2750 3189 2751
rect 3574 2751 3580 2752
rect 3188 2748 3233 2750
rect 3188 2747 3189 2748
rect 3183 2746 3189 2747
rect 3574 2747 3575 2751
rect 3579 2747 3580 2751
rect 3574 2746 3580 2747
rect 983 2743 989 2744
rect 983 2742 984 2743
rect 936 2740 984 2742
rect 551 2739 557 2740
rect 551 2738 552 2739
rect 336 2736 552 2738
rect 135 2731 141 2732
rect 135 2727 136 2731
rect 140 2730 141 2731
rect 210 2731 216 2732
rect 210 2730 211 2731
rect 140 2728 211 2730
rect 140 2727 141 2728
rect 135 2726 141 2727
rect 210 2727 211 2728
rect 215 2727 216 2731
rect 210 2726 216 2727
rect 223 2731 229 2732
rect 223 2727 224 2731
rect 228 2730 229 2731
rect 336 2730 338 2736
rect 551 2735 552 2736
rect 556 2735 557 2739
rect 983 2739 984 2740
rect 988 2739 989 2743
rect 983 2738 989 2739
rect 1886 2741 1892 2742
rect 1886 2737 1887 2741
rect 1891 2737 1892 2741
rect 1886 2736 1892 2737
rect 2054 2741 2060 2742
rect 2054 2737 2055 2741
rect 2059 2737 2060 2741
rect 2054 2736 2060 2737
rect 2246 2741 2252 2742
rect 2246 2737 2247 2741
rect 2251 2737 2252 2741
rect 2246 2736 2252 2737
rect 2430 2741 2436 2742
rect 2430 2737 2431 2741
rect 2435 2737 2436 2741
rect 2430 2736 2436 2737
rect 2606 2741 2612 2742
rect 2606 2737 2607 2741
rect 2611 2737 2612 2741
rect 2606 2736 2612 2737
rect 2774 2741 2780 2742
rect 2774 2737 2775 2741
rect 2779 2737 2780 2741
rect 2774 2736 2780 2737
rect 2926 2741 2932 2742
rect 2926 2737 2927 2741
rect 2931 2737 2932 2741
rect 2926 2736 2932 2737
rect 3070 2741 3076 2742
rect 3070 2737 3071 2741
rect 3075 2737 3076 2741
rect 3070 2736 3076 2737
rect 3214 2741 3220 2742
rect 3214 2737 3215 2741
rect 3219 2737 3220 2741
rect 3214 2736 3220 2737
rect 3358 2741 3364 2742
rect 3358 2737 3359 2741
rect 3363 2737 3364 2741
rect 3358 2736 3364 2737
rect 3478 2741 3484 2742
rect 3478 2737 3479 2741
rect 3483 2737 3484 2741
rect 3478 2736 3484 2737
rect 551 2734 557 2735
rect 2974 2735 2981 2736
rect 228 2728 338 2730
rect 343 2731 349 2732
rect 228 2727 229 2728
rect 223 2726 229 2727
rect 343 2727 344 2731
rect 348 2730 349 2731
rect 362 2731 368 2732
rect 362 2730 363 2731
rect 348 2728 363 2730
rect 348 2727 349 2728
rect 343 2726 349 2727
rect 362 2727 363 2728
rect 367 2727 368 2731
rect 362 2726 368 2727
rect 415 2731 421 2732
rect 415 2727 416 2731
rect 420 2730 421 2731
rect 471 2731 477 2732
rect 471 2730 472 2731
rect 420 2728 472 2730
rect 420 2727 421 2728
rect 415 2726 421 2727
rect 471 2727 472 2728
rect 476 2727 477 2731
rect 471 2726 477 2727
rect 543 2731 549 2732
rect 543 2727 544 2731
rect 548 2730 549 2731
rect 607 2731 613 2732
rect 607 2730 608 2731
rect 548 2728 608 2730
rect 548 2727 549 2728
rect 543 2726 549 2727
rect 607 2727 608 2728
rect 612 2727 613 2731
rect 607 2726 613 2727
rect 687 2731 693 2732
rect 687 2727 688 2731
rect 692 2730 693 2731
rect 751 2731 757 2732
rect 751 2730 752 2731
rect 692 2728 752 2730
rect 692 2727 693 2728
rect 687 2726 693 2727
rect 751 2727 752 2728
rect 756 2727 757 2731
rect 751 2726 757 2727
rect 831 2731 837 2732
rect 831 2727 832 2731
rect 836 2730 837 2731
rect 895 2731 901 2732
rect 895 2730 896 2731
rect 836 2728 896 2730
rect 836 2727 837 2728
rect 831 2726 837 2727
rect 895 2727 896 2728
rect 900 2727 901 2731
rect 895 2726 901 2727
rect 975 2731 981 2732
rect 975 2727 976 2731
rect 980 2730 981 2731
rect 1039 2731 1045 2732
rect 1039 2730 1040 2731
rect 980 2728 1040 2730
rect 980 2727 981 2728
rect 975 2726 981 2727
rect 1039 2727 1040 2728
rect 1044 2727 1045 2731
rect 2974 2731 2975 2735
rect 2980 2731 2981 2735
rect 2974 2730 2981 2731
rect 1039 2726 1045 2727
rect 2846 2727 2852 2728
rect 2846 2723 2847 2727
rect 2851 2726 2852 2727
rect 3183 2727 3189 2728
rect 3183 2726 3184 2727
rect 2851 2724 3184 2726
rect 2851 2723 2852 2724
rect 2846 2722 2852 2723
rect 3183 2723 3184 2724
rect 3188 2723 3189 2727
rect 3183 2722 3189 2723
rect 142 2721 148 2722
rect 142 2717 143 2721
rect 147 2717 148 2721
rect 142 2716 148 2717
rect 230 2721 236 2722
rect 230 2717 231 2721
rect 235 2717 236 2721
rect 230 2716 236 2717
rect 350 2721 356 2722
rect 350 2717 351 2721
rect 355 2717 356 2721
rect 350 2716 356 2717
rect 478 2721 484 2722
rect 478 2717 479 2721
rect 483 2717 484 2721
rect 478 2716 484 2717
rect 614 2721 620 2722
rect 614 2717 615 2721
rect 619 2717 620 2721
rect 614 2716 620 2717
rect 758 2721 764 2722
rect 758 2717 759 2721
rect 763 2717 764 2721
rect 758 2716 764 2717
rect 902 2721 908 2722
rect 902 2717 903 2721
rect 907 2717 908 2721
rect 902 2716 908 2717
rect 1046 2721 1052 2722
rect 1046 2717 1047 2721
rect 1051 2717 1052 2721
rect 1046 2716 1052 2717
rect 1886 2715 1892 2716
rect 1886 2711 1887 2715
rect 1891 2711 1892 2715
rect 1886 2710 1892 2711
rect 2046 2715 2052 2716
rect 2046 2711 2047 2715
rect 2051 2711 2052 2715
rect 2046 2710 2052 2711
rect 2206 2715 2212 2716
rect 2206 2711 2207 2715
rect 2211 2711 2212 2715
rect 2206 2710 2212 2711
rect 2358 2715 2364 2716
rect 2358 2711 2359 2715
rect 2363 2711 2364 2715
rect 2358 2710 2364 2711
rect 2494 2715 2500 2716
rect 2494 2711 2495 2715
rect 2499 2711 2500 2715
rect 2494 2710 2500 2711
rect 2622 2715 2628 2716
rect 2622 2711 2623 2715
rect 2627 2711 2628 2715
rect 2622 2710 2628 2711
rect 2742 2715 2748 2716
rect 2742 2711 2743 2715
rect 2747 2711 2748 2715
rect 2742 2710 2748 2711
rect 2862 2715 2868 2716
rect 2862 2711 2863 2715
rect 2867 2711 2868 2715
rect 2862 2710 2868 2711
rect 2982 2715 2988 2716
rect 2982 2711 2983 2715
rect 2987 2711 2988 2715
rect 2982 2710 2988 2711
rect 3102 2715 3108 2716
rect 3102 2711 3103 2715
rect 3107 2711 3108 2715
rect 3102 2710 3108 2711
rect 110 2708 116 2709
rect 1822 2708 1828 2709
rect 110 2704 111 2708
rect 115 2704 116 2708
rect 415 2707 421 2708
rect 415 2706 416 2707
rect 405 2704 416 2706
rect 110 2703 116 2704
rect 210 2703 216 2704
rect 210 2699 211 2703
rect 215 2702 216 2703
rect 415 2703 416 2704
rect 420 2703 421 2707
rect 543 2707 549 2708
rect 543 2706 544 2707
rect 533 2704 544 2706
rect 415 2702 421 2703
rect 543 2703 544 2704
rect 548 2703 549 2707
rect 831 2707 837 2708
rect 831 2706 832 2707
rect 813 2704 832 2706
rect 543 2702 549 2703
rect 551 2703 557 2704
rect 215 2700 249 2702
rect 215 2699 216 2700
rect 210 2698 216 2699
rect 551 2699 552 2703
rect 556 2702 557 2703
rect 831 2703 832 2704
rect 836 2703 837 2707
rect 975 2707 981 2708
rect 975 2706 976 2707
rect 957 2704 976 2706
rect 831 2702 837 2703
rect 975 2703 976 2704
rect 980 2703 981 2707
rect 1822 2704 1823 2708
rect 1827 2704 1828 2708
rect 2562 2707 2568 2708
rect 2562 2706 2563 2707
rect 975 2702 981 2703
rect 983 2703 989 2704
rect 1822 2703 1828 2704
rect 1862 2705 1868 2706
rect 556 2700 633 2702
rect 556 2699 557 2700
rect 551 2698 557 2699
rect 983 2699 984 2703
rect 988 2702 989 2703
rect 988 2700 1065 2702
rect 1862 2701 1863 2705
rect 1867 2701 1868 2705
rect 2553 2704 2563 2706
rect 2562 2703 2563 2704
rect 2567 2703 2568 2707
rect 2562 2702 2568 2703
rect 3050 2707 3056 2708
rect 3050 2703 3051 2707
rect 3055 2706 3056 2707
rect 3055 2704 3121 2706
rect 3574 2705 3580 2706
rect 3055 2703 3056 2704
rect 3050 2702 3056 2703
rect 1862 2700 1868 2701
rect 3574 2701 3575 2705
rect 3579 2701 3580 2705
rect 3574 2700 3580 2701
rect 988 2699 989 2700
rect 983 2698 989 2699
rect 110 2691 116 2692
rect 110 2687 111 2691
rect 115 2687 116 2691
rect 110 2686 116 2687
rect 127 2691 133 2692
rect 127 2687 128 2691
rect 132 2690 133 2691
rect 1822 2691 1828 2692
rect 132 2688 153 2690
rect 132 2687 133 2688
rect 127 2686 133 2687
rect 1822 2687 1823 2691
rect 1827 2687 1828 2691
rect 1879 2691 1885 2692
rect 1822 2686 1828 2687
rect 1862 2688 1868 2689
rect 1862 2684 1863 2688
rect 1867 2684 1868 2688
rect 1879 2687 1880 2691
rect 1884 2690 1885 2691
rect 1954 2691 1960 2692
rect 1884 2688 1913 2690
rect 1884 2687 1885 2688
rect 1879 2686 1885 2687
rect 1954 2687 1955 2691
rect 1959 2690 1960 2691
rect 2351 2691 2357 2692
rect 2351 2690 2352 2691
rect 1959 2688 2073 2690
rect 2269 2688 2352 2690
rect 1959 2687 1960 2688
rect 1954 2686 1960 2687
rect 2351 2687 2352 2688
rect 2356 2687 2357 2691
rect 2487 2691 2493 2692
rect 2487 2690 2488 2691
rect 2421 2688 2488 2690
rect 2351 2686 2357 2687
rect 2487 2687 2488 2688
rect 2492 2687 2493 2691
rect 2690 2691 2696 2692
rect 2690 2690 2691 2691
rect 2685 2688 2691 2690
rect 2487 2686 2493 2687
rect 2690 2687 2691 2688
rect 2695 2687 2696 2691
rect 2690 2686 2696 2687
rect 2698 2691 2704 2692
rect 2698 2687 2699 2691
rect 2703 2690 2704 2691
rect 2810 2691 2816 2692
rect 2703 2688 2769 2690
rect 2703 2687 2704 2688
rect 2698 2686 2704 2687
rect 2810 2687 2811 2691
rect 2815 2690 2816 2691
rect 3095 2691 3101 2692
rect 3095 2690 3096 2691
rect 2815 2688 2889 2690
rect 3045 2688 3096 2690
rect 2815 2687 2816 2688
rect 2810 2686 2816 2687
rect 3095 2687 3096 2688
rect 3100 2687 3101 2691
rect 3095 2686 3101 2687
rect 3574 2688 3580 2689
rect 1862 2683 1868 2684
rect 3574 2684 3575 2688
rect 3579 2684 3580 2688
rect 3574 2683 3580 2684
rect 134 2681 140 2682
rect 134 2677 135 2681
rect 139 2677 140 2681
rect 134 2676 140 2677
rect 222 2681 228 2682
rect 222 2677 223 2681
rect 227 2677 228 2681
rect 222 2676 228 2677
rect 342 2681 348 2682
rect 342 2677 343 2681
rect 347 2677 348 2681
rect 342 2676 348 2677
rect 470 2681 476 2682
rect 470 2677 471 2681
rect 475 2677 476 2681
rect 470 2676 476 2677
rect 606 2681 612 2682
rect 606 2677 607 2681
rect 611 2677 612 2681
rect 606 2676 612 2677
rect 750 2681 756 2682
rect 750 2677 751 2681
rect 755 2677 756 2681
rect 750 2676 756 2677
rect 894 2681 900 2682
rect 894 2677 895 2681
rect 899 2677 900 2681
rect 894 2676 900 2677
rect 1038 2681 1044 2682
rect 1038 2677 1039 2681
rect 1043 2677 1044 2681
rect 1038 2676 1044 2677
rect 1894 2675 1900 2676
rect 1894 2671 1895 2675
rect 1899 2671 1900 2675
rect 1894 2670 1900 2671
rect 2054 2675 2060 2676
rect 2054 2671 2055 2675
rect 2059 2671 2060 2675
rect 2054 2670 2060 2671
rect 2214 2675 2220 2676
rect 2214 2671 2215 2675
rect 2219 2671 2220 2675
rect 2214 2670 2220 2671
rect 2366 2675 2372 2676
rect 2366 2671 2367 2675
rect 2371 2671 2372 2675
rect 2366 2670 2372 2671
rect 2502 2675 2508 2676
rect 2502 2671 2503 2675
rect 2507 2671 2508 2675
rect 2502 2670 2508 2671
rect 2630 2675 2636 2676
rect 2630 2671 2631 2675
rect 2635 2671 2636 2675
rect 2630 2670 2636 2671
rect 2750 2675 2756 2676
rect 2750 2671 2751 2675
rect 2755 2671 2756 2675
rect 2750 2670 2756 2671
rect 2870 2675 2876 2676
rect 2870 2671 2871 2675
rect 2875 2671 2876 2675
rect 2870 2670 2876 2671
rect 2990 2675 2996 2676
rect 2990 2671 2991 2675
rect 2995 2671 2996 2675
rect 2990 2670 2996 2671
rect 3110 2675 3116 2676
rect 3110 2671 3111 2675
rect 3115 2671 3116 2675
rect 3110 2670 3116 2671
rect 1887 2663 1893 2664
rect 1887 2659 1888 2663
rect 1892 2662 1893 2663
rect 1954 2663 1960 2664
rect 1954 2662 1955 2663
rect 1892 2660 1955 2662
rect 1892 2659 1893 2660
rect 1887 2658 1893 2659
rect 1954 2659 1955 2660
rect 1959 2659 1960 2663
rect 1954 2658 1960 2659
rect 2039 2663 2045 2664
rect 2039 2659 2040 2663
rect 2044 2662 2045 2663
rect 2047 2663 2053 2664
rect 2047 2662 2048 2663
rect 2044 2660 2048 2662
rect 2044 2659 2045 2660
rect 2039 2658 2045 2659
rect 2047 2659 2048 2660
rect 2052 2659 2053 2663
rect 2047 2658 2053 2659
rect 2207 2663 2213 2664
rect 2207 2659 2208 2663
rect 2212 2662 2213 2663
rect 2326 2663 2332 2664
rect 2326 2662 2327 2663
rect 2212 2660 2327 2662
rect 2212 2659 2213 2660
rect 2207 2658 2213 2659
rect 2326 2659 2327 2660
rect 2331 2659 2332 2663
rect 2326 2658 2332 2659
rect 2351 2663 2357 2664
rect 2351 2659 2352 2663
rect 2356 2662 2357 2663
rect 2359 2663 2365 2664
rect 2359 2662 2360 2663
rect 2356 2660 2360 2662
rect 2356 2659 2357 2660
rect 2351 2658 2357 2659
rect 2359 2659 2360 2660
rect 2364 2659 2365 2663
rect 2359 2658 2365 2659
rect 2487 2663 2493 2664
rect 2487 2659 2488 2663
rect 2492 2662 2493 2663
rect 2495 2663 2501 2664
rect 2495 2662 2496 2663
rect 2492 2660 2496 2662
rect 2492 2659 2493 2660
rect 2487 2658 2493 2659
rect 2495 2659 2496 2660
rect 2500 2659 2501 2663
rect 2495 2658 2501 2659
rect 2623 2663 2629 2664
rect 2623 2659 2624 2663
rect 2628 2662 2629 2663
rect 2698 2663 2704 2664
rect 2698 2662 2699 2663
rect 2628 2660 2699 2662
rect 2628 2659 2629 2660
rect 2623 2658 2629 2659
rect 2698 2659 2699 2660
rect 2703 2659 2704 2663
rect 2698 2658 2704 2659
rect 2743 2663 2749 2664
rect 2743 2659 2744 2663
rect 2748 2662 2749 2663
rect 2810 2663 2816 2664
rect 2810 2662 2811 2663
rect 2748 2660 2811 2662
rect 2748 2659 2749 2660
rect 2743 2658 2749 2659
rect 2810 2659 2811 2660
rect 2815 2659 2816 2663
rect 2810 2658 2816 2659
rect 2863 2663 2869 2664
rect 2863 2659 2864 2663
rect 2868 2662 2869 2663
rect 2974 2663 2980 2664
rect 2868 2660 2970 2662
rect 2868 2659 2869 2660
rect 2863 2658 2869 2659
rect 134 2655 140 2656
rect 134 2651 135 2655
rect 139 2651 140 2655
rect 134 2650 140 2651
rect 230 2655 236 2656
rect 230 2651 231 2655
rect 235 2651 236 2655
rect 230 2650 236 2651
rect 350 2655 356 2656
rect 350 2651 351 2655
rect 355 2651 356 2655
rect 350 2650 356 2651
rect 470 2655 476 2656
rect 470 2651 471 2655
rect 475 2651 476 2655
rect 470 2650 476 2651
rect 582 2655 588 2656
rect 582 2651 583 2655
rect 587 2651 588 2655
rect 582 2650 588 2651
rect 694 2655 700 2656
rect 694 2651 695 2655
rect 699 2651 700 2655
rect 694 2650 700 2651
rect 798 2655 804 2656
rect 798 2651 799 2655
rect 803 2651 804 2655
rect 798 2650 804 2651
rect 902 2655 908 2656
rect 902 2651 903 2655
rect 907 2651 908 2655
rect 902 2650 908 2651
rect 998 2655 1004 2656
rect 998 2651 999 2655
rect 1003 2651 1004 2655
rect 998 2650 1004 2651
rect 1102 2655 1108 2656
rect 1102 2651 1103 2655
rect 1107 2651 1108 2655
rect 1102 2650 1108 2651
rect 1206 2655 1212 2656
rect 1206 2651 1207 2655
rect 1211 2651 1212 2655
rect 1206 2650 1212 2651
rect 1310 2655 1316 2656
rect 1310 2651 1311 2655
rect 1315 2651 1316 2655
rect 2968 2654 2970 2660
rect 2974 2659 2975 2663
rect 2979 2662 2980 2663
rect 2983 2663 2989 2664
rect 2983 2662 2984 2663
rect 2979 2660 2984 2662
rect 2979 2659 2980 2660
rect 2974 2658 2980 2659
rect 2983 2659 2984 2660
rect 2988 2659 2989 2663
rect 2983 2658 2989 2659
rect 3095 2663 3101 2664
rect 3095 2659 3096 2663
rect 3100 2662 3101 2663
rect 3103 2663 3109 2664
rect 3103 2662 3104 2663
rect 3100 2660 3104 2662
rect 3100 2659 3101 2660
rect 3095 2658 3101 2659
rect 3103 2659 3104 2660
rect 3108 2659 3109 2663
rect 3103 2658 3109 2659
rect 3050 2655 3056 2656
rect 3050 2654 3051 2655
rect 2968 2652 3051 2654
rect 1310 2650 1316 2651
rect 2831 2651 2837 2652
rect 2831 2650 2832 2651
rect 2640 2648 2832 2650
rect 422 2647 428 2648
rect 110 2645 116 2646
rect 110 2641 111 2645
rect 115 2641 116 2645
rect 422 2643 423 2647
rect 427 2646 428 2647
rect 687 2647 693 2648
rect 687 2646 688 2647
rect 427 2644 489 2646
rect 641 2644 688 2646
rect 427 2643 428 2644
rect 422 2642 428 2643
rect 687 2643 688 2644
rect 692 2643 693 2647
rect 687 2642 693 2643
rect 1274 2647 1280 2648
rect 1274 2643 1275 2647
rect 1279 2646 1280 2647
rect 1279 2644 1329 2646
rect 1822 2645 1828 2646
rect 1279 2643 1280 2644
rect 1274 2642 1280 2643
rect 110 2640 116 2641
rect 1822 2641 1823 2645
rect 1827 2641 1828 2645
rect 1822 2640 1828 2641
rect 1879 2643 1885 2644
rect 1879 2639 1880 2643
rect 1884 2642 1885 2643
rect 1887 2643 1893 2644
rect 1887 2642 1888 2643
rect 1884 2640 1888 2642
rect 1884 2639 1885 2640
rect 1879 2638 1885 2639
rect 1887 2639 1888 2640
rect 1892 2639 1893 2643
rect 1887 2638 1893 2639
rect 1959 2643 1965 2644
rect 1959 2639 1960 2643
rect 1964 2642 1965 2643
rect 1991 2643 1997 2644
rect 1991 2642 1992 2643
rect 1964 2640 1992 2642
rect 1964 2639 1965 2640
rect 1959 2638 1965 2639
rect 1991 2639 1992 2640
rect 1996 2639 1997 2643
rect 1991 2638 1997 2639
rect 2103 2643 2109 2644
rect 2103 2639 2104 2643
rect 2108 2642 2109 2643
rect 2111 2643 2117 2644
rect 2111 2642 2112 2643
rect 2108 2640 2112 2642
rect 2108 2639 2109 2640
rect 2103 2638 2109 2639
rect 2111 2639 2112 2640
rect 2116 2639 2117 2643
rect 2111 2638 2117 2639
rect 2183 2643 2189 2644
rect 2183 2639 2184 2643
rect 2188 2642 2189 2643
rect 2231 2643 2237 2644
rect 2231 2642 2232 2643
rect 2188 2640 2232 2642
rect 2188 2639 2189 2640
rect 2183 2638 2189 2639
rect 2231 2639 2232 2640
rect 2236 2639 2237 2643
rect 2231 2638 2237 2639
rect 2314 2643 2320 2644
rect 2314 2639 2315 2643
rect 2319 2642 2320 2643
rect 2343 2643 2349 2644
rect 2343 2642 2344 2643
rect 2319 2640 2344 2642
rect 2319 2639 2320 2640
rect 2314 2638 2320 2639
rect 2343 2639 2344 2640
rect 2348 2639 2349 2643
rect 2343 2638 2349 2639
rect 2447 2643 2453 2644
rect 2447 2639 2448 2643
rect 2452 2642 2453 2643
rect 2522 2643 2528 2644
rect 2522 2642 2523 2643
rect 2452 2640 2523 2642
rect 2452 2639 2453 2640
rect 2447 2638 2453 2639
rect 2522 2639 2523 2640
rect 2527 2639 2528 2643
rect 2522 2638 2528 2639
rect 2543 2643 2549 2644
rect 2543 2639 2544 2643
rect 2548 2642 2549 2643
rect 2640 2642 2642 2648
rect 2831 2647 2832 2648
rect 2836 2647 2837 2651
rect 3050 2651 3051 2652
rect 3055 2651 3056 2655
rect 3050 2650 3056 2651
rect 2831 2646 2837 2647
rect 2548 2640 2642 2642
rect 2647 2643 2653 2644
rect 2548 2639 2549 2640
rect 2543 2638 2549 2639
rect 2647 2639 2648 2643
rect 2652 2642 2653 2643
rect 2690 2643 2696 2644
rect 2690 2642 2691 2643
rect 2652 2640 2691 2642
rect 2652 2639 2653 2640
rect 2647 2638 2653 2639
rect 2690 2639 2691 2640
rect 2695 2639 2696 2643
rect 2690 2638 2696 2639
rect 2719 2643 2725 2644
rect 2719 2639 2720 2643
rect 2724 2642 2725 2643
rect 2751 2643 2757 2644
rect 2751 2642 2752 2643
rect 2724 2640 2752 2642
rect 2724 2639 2725 2640
rect 2719 2638 2725 2639
rect 2751 2639 2752 2640
rect 2756 2639 2757 2643
rect 2751 2638 2757 2639
rect 2823 2643 2829 2644
rect 2823 2639 2824 2643
rect 2828 2642 2829 2643
rect 2855 2643 2861 2644
rect 2855 2642 2856 2643
rect 2828 2640 2856 2642
rect 2828 2639 2829 2640
rect 2823 2638 2829 2639
rect 2855 2639 2856 2640
rect 2860 2639 2861 2643
rect 2855 2638 2861 2639
rect 1894 2633 1900 2634
rect 223 2631 229 2632
rect 223 2630 224 2631
rect 110 2628 116 2629
rect 197 2628 224 2630
rect 110 2624 111 2628
rect 115 2624 116 2628
rect 223 2627 224 2628
rect 228 2627 229 2631
rect 343 2631 349 2632
rect 343 2630 344 2631
rect 293 2628 344 2630
rect 223 2626 229 2627
rect 343 2627 344 2628
rect 348 2627 349 2631
rect 463 2631 469 2632
rect 463 2630 464 2631
rect 413 2628 464 2630
rect 343 2626 349 2627
rect 463 2627 464 2628
rect 468 2627 469 2631
rect 791 2631 797 2632
rect 791 2630 792 2631
rect 757 2628 792 2630
rect 463 2626 469 2627
rect 791 2627 792 2628
rect 796 2627 797 2631
rect 895 2631 901 2632
rect 895 2630 896 2631
rect 861 2628 896 2630
rect 791 2626 797 2627
rect 895 2627 896 2628
rect 900 2627 901 2631
rect 991 2631 997 2632
rect 991 2630 992 2631
rect 965 2628 992 2630
rect 895 2626 901 2627
rect 991 2627 992 2628
rect 996 2627 997 2631
rect 1095 2631 1101 2632
rect 1095 2630 1096 2631
rect 1061 2628 1096 2630
rect 991 2626 997 2627
rect 1095 2627 1096 2628
rect 1100 2627 1101 2631
rect 1199 2631 1205 2632
rect 1199 2630 1200 2631
rect 1165 2628 1200 2630
rect 1095 2626 1101 2627
rect 1199 2627 1200 2628
rect 1204 2627 1205 2631
rect 1303 2631 1309 2632
rect 1303 2630 1304 2631
rect 1269 2628 1304 2630
rect 1199 2626 1205 2627
rect 1303 2627 1304 2628
rect 1308 2627 1309 2631
rect 1894 2629 1895 2633
rect 1899 2629 1900 2633
rect 1303 2626 1309 2627
rect 1822 2628 1828 2629
rect 1894 2628 1900 2629
rect 1998 2633 2004 2634
rect 1998 2629 1999 2633
rect 2003 2629 2004 2633
rect 1998 2628 2004 2629
rect 2118 2633 2124 2634
rect 2118 2629 2119 2633
rect 2123 2629 2124 2633
rect 2118 2628 2124 2629
rect 2238 2633 2244 2634
rect 2238 2629 2239 2633
rect 2243 2629 2244 2633
rect 2238 2628 2244 2629
rect 2350 2633 2356 2634
rect 2350 2629 2351 2633
rect 2355 2629 2356 2633
rect 2350 2628 2356 2629
rect 2454 2633 2460 2634
rect 2454 2629 2455 2633
rect 2459 2629 2460 2633
rect 2454 2628 2460 2629
rect 2550 2633 2556 2634
rect 2550 2629 2551 2633
rect 2555 2629 2556 2633
rect 2550 2628 2556 2629
rect 2654 2633 2660 2634
rect 2654 2629 2655 2633
rect 2659 2629 2660 2633
rect 2654 2628 2660 2629
rect 2758 2633 2764 2634
rect 2758 2629 2759 2633
rect 2763 2629 2764 2633
rect 2758 2628 2764 2629
rect 2862 2633 2868 2634
rect 2862 2629 2863 2633
rect 2867 2629 2868 2633
rect 2862 2628 2868 2629
rect 110 2623 116 2624
rect 1822 2624 1823 2628
rect 1827 2624 1828 2628
rect 1822 2623 1828 2624
rect 1862 2620 1868 2621
rect 3574 2620 3580 2621
rect 1862 2616 1863 2620
rect 1867 2616 1868 2620
rect 1959 2619 1965 2620
rect 1959 2618 1960 2619
rect 1949 2616 1960 2618
rect 142 2615 148 2616
rect 142 2611 143 2615
rect 147 2611 148 2615
rect 142 2610 148 2611
rect 238 2615 244 2616
rect 238 2611 239 2615
rect 243 2611 244 2615
rect 238 2610 244 2611
rect 358 2615 364 2616
rect 358 2611 359 2615
rect 363 2611 364 2615
rect 358 2610 364 2611
rect 478 2615 484 2616
rect 478 2611 479 2615
rect 483 2611 484 2615
rect 478 2610 484 2611
rect 590 2615 596 2616
rect 590 2611 591 2615
rect 595 2611 596 2615
rect 590 2610 596 2611
rect 702 2615 708 2616
rect 702 2611 703 2615
rect 707 2611 708 2615
rect 702 2610 708 2611
rect 806 2615 812 2616
rect 806 2611 807 2615
rect 811 2611 812 2615
rect 806 2610 812 2611
rect 910 2615 916 2616
rect 910 2611 911 2615
rect 915 2611 916 2615
rect 910 2610 916 2611
rect 1006 2615 1012 2616
rect 1006 2611 1007 2615
rect 1011 2611 1012 2615
rect 1006 2610 1012 2611
rect 1110 2615 1116 2616
rect 1110 2611 1111 2615
rect 1115 2611 1116 2615
rect 1110 2610 1116 2611
rect 1214 2615 1220 2616
rect 1214 2611 1215 2615
rect 1219 2611 1220 2615
rect 1214 2610 1220 2611
rect 1318 2615 1324 2616
rect 1862 2615 1868 2616
rect 1959 2615 1960 2616
rect 1964 2615 1965 2619
rect 2183 2619 2189 2620
rect 2183 2618 2184 2619
rect 2173 2616 2184 2618
rect 1318 2611 1319 2615
rect 1323 2611 1324 2615
rect 1959 2614 1965 2615
rect 2183 2615 2184 2616
rect 2188 2615 2189 2619
rect 2314 2619 2320 2620
rect 2314 2618 2315 2619
rect 2293 2616 2315 2618
rect 2183 2614 2189 2615
rect 2314 2615 2315 2616
rect 2319 2615 2320 2619
rect 2719 2619 2725 2620
rect 2719 2618 2720 2619
rect 2709 2616 2720 2618
rect 2314 2614 2320 2615
rect 2326 2615 2332 2616
rect 1318 2610 1324 2611
rect 2326 2611 2327 2615
rect 2331 2614 2332 2615
rect 2522 2615 2528 2616
rect 2331 2612 2369 2614
rect 2331 2611 2332 2612
rect 2326 2610 2332 2611
rect 2522 2611 2523 2615
rect 2527 2614 2528 2615
rect 2719 2615 2720 2616
rect 2724 2615 2725 2619
rect 2823 2619 2829 2620
rect 2823 2618 2824 2619
rect 2813 2616 2824 2618
rect 2719 2614 2725 2615
rect 2823 2615 2824 2616
rect 2828 2615 2829 2619
rect 3574 2616 3575 2620
rect 3579 2616 3580 2620
rect 2823 2614 2829 2615
rect 2831 2615 2837 2616
rect 3574 2615 3580 2616
rect 2527 2612 2569 2614
rect 2527 2611 2528 2612
rect 2522 2610 2528 2611
rect 2831 2611 2832 2615
rect 2836 2614 2837 2615
rect 2836 2612 2881 2614
rect 2836 2611 2837 2612
rect 2831 2610 2837 2611
rect 127 2603 133 2604
rect 127 2599 128 2603
rect 132 2602 133 2603
rect 135 2603 141 2604
rect 135 2602 136 2603
rect 132 2600 136 2602
rect 132 2599 133 2600
rect 127 2598 133 2599
rect 135 2599 136 2600
rect 140 2599 141 2603
rect 135 2598 141 2599
rect 223 2603 229 2604
rect 223 2599 224 2603
rect 228 2602 229 2603
rect 231 2603 237 2604
rect 231 2602 232 2603
rect 228 2600 232 2602
rect 228 2599 229 2600
rect 223 2598 229 2599
rect 231 2599 232 2600
rect 236 2599 237 2603
rect 231 2598 237 2599
rect 343 2603 349 2604
rect 343 2599 344 2603
rect 348 2602 349 2603
rect 351 2603 357 2604
rect 351 2602 352 2603
rect 348 2600 352 2602
rect 348 2599 349 2600
rect 343 2598 349 2599
rect 351 2599 352 2600
rect 356 2599 357 2603
rect 351 2598 357 2599
rect 463 2603 469 2604
rect 463 2599 464 2603
rect 468 2602 469 2603
rect 471 2603 477 2604
rect 471 2602 472 2603
rect 468 2600 472 2602
rect 468 2599 469 2600
rect 463 2598 469 2599
rect 471 2599 472 2600
rect 476 2599 477 2603
rect 471 2598 477 2599
rect 583 2603 589 2604
rect 583 2599 584 2603
rect 588 2602 589 2603
rect 618 2603 624 2604
rect 618 2602 619 2603
rect 588 2600 619 2602
rect 588 2599 589 2600
rect 583 2598 589 2599
rect 618 2599 619 2600
rect 623 2599 624 2603
rect 618 2598 624 2599
rect 695 2603 701 2604
rect 695 2599 696 2603
rect 700 2602 701 2603
rect 746 2603 752 2604
rect 746 2602 747 2603
rect 700 2600 747 2602
rect 700 2599 701 2600
rect 695 2598 701 2599
rect 746 2599 747 2600
rect 751 2599 752 2603
rect 746 2598 752 2599
rect 791 2603 797 2604
rect 791 2599 792 2603
rect 796 2602 797 2603
rect 799 2603 805 2604
rect 799 2602 800 2603
rect 796 2600 800 2602
rect 796 2599 797 2600
rect 791 2598 797 2599
rect 799 2599 800 2600
rect 804 2599 805 2603
rect 799 2598 805 2599
rect 895 2603 901 2604
rect 895 2599 896 2603
rect 900 2602 901 2603
rect 903 2603 909 2604
rect 903 2602 904 2603
rect 900 2600 904 2602
rect 900 2599 901 2600
rect 895 2598 901 2599
rect 903 2599 904 2600
rect 908 2599 909 2603
rect 903 2598 909 2599
rect 991 2603 997 2604
rect 991 2599 992 2603
rect 996 2602 997 2603
rect 999 2603 1005 2604
rect 999 2602 1000 2603
rect 996 2600 1000 2602
rect 996 2599 997 2600
rect 991 2598 997 2599
rect 999 2599 1000 2600
rect 1004 2599 1005 2603
rect 999 2598 1005 2599
rect 1095 2603 1101 2604
rect 1095 2599 1096 2603
rect 1100 2602 1101 2603
rect 1103 2603 1109 2604
rect 1103 2602 1104 2603
rect 1100 2600 1104 2602
rect 1100 2599 1101 2600
rect 1095 2598 1101 2599
rect 1103 2599 1104 2600
rect 1108 2599 1109 2603
rect 1103 2598 1109 2599
rect 1199 2603 1205 2604
rect 1199 2599 1200 2603
rect 1204 2602 1205 2603
rect 1207 2603 1213 2604
rect 1207 2602 1208 2603
rect 1204 2600 1208 2602
rect 1204 2599 1205 2600
rect 1199 2598 1205 2599
rect 1207 2599 1208 2600
rect 1212 2599 1213 2603
rect 1207 2598 1213 2599
rect 1303 2603 1309 2604
rect 1303 2599 1304 2603
rect 1308 2602 1309 2603
rect 1311 2603 1317 2604
rect 1311 2602 1312 2603
rect 1308 2600 1312 2602
rect 1308 2599 1309 2600
rect 1303 2598 1309 2599
rect 1311 2599 1312 2600
rect 1316 2599 1317 2603
rect 1311 2598 1317 2599
rect 1862 2603 1868 2604
rect 1862 2599 1863 2603
rect 1867 2599 1868 2603
rect 1862 2598 1868 2599
rect 1983 2603 1989 2604
rect 1983 2599 1984 2603
rect 1988 2602 1989 2603
rect 3574 2603 3580 2604
rect 1988 2600 2009 2602
rect 1988 2599 1989 2600
rect 1983 2598 1989 2599
rect 3574 2599 3575 2603
rect 3579 2599 3580 2603
rect 3574 2598 3580 2599
rect 1886 2593 1892 2594
rect 1886 2589 1887 2593
rect 1891 2589 1892 2593
rect 1886 2588 1892 2589
rect 1990 2593 1996 2594
rect 1990 2589 1991 2593
rect 1995 2589 1996 2593
rect 1990 2588 1996 2589
rect 2110 2593 2116 2594
rect 2110 2589 2111 2593
rect 2115 2589 2116 2593
rect 2110 2588 2116 2589
rect 2230 2593 2236 2594
rect 2230 2589 2231 2593
rect 2235 2589 2236 2593
rect 2230 2588 2236 2589
rect 2342 2593 2348 2594
rect 2342 2589 2343 2593
rect 2347 2589 2348 2593
rect 2342 2588 2348 2589
rect 2446 2593 2452 2594
rect 2446 2589 2447 2593
rect 2451 2589 2452 2593
rect 2446 2588 2452 2589
rect 2542 2593 2548 2594
rect 2542 2589 2543 2593
rect 2547 2589 2548 2593
rect 2542 2588 2548 2589
rect 2646 2593 2652 2594
rect 2646 2589 2647 2593
rect 2651 2589 2652 2593
rect 2646 2588 2652 2589
rect 2750 2593 2756 2594
rect 2750 2589 2751 2593
rect 2755 2589 2756 2593
rect 2750 2588 2756 2589
rect 2854 2593 2860 2594
rect 2854 2589 2855 2593
rect 2859 2589 2860 2593
rect 2854 2588 2860 2589
rect 135 2587 141 2588
rect 135 2583 136 2587
rect 140 2586 141 2587
rect 210 2587 216 2588
rect 210 2586 211 2587
rect 140 2584 211 2586
rect 140 2583 141 2584
rect 135 2582 141 2583
rect 210 2583 211 2584
rect 215 2583 216 2587
rect 210 2582 216 2583
rect 263 2587 269 2588
rect 263 2583 264 2587
rect 268 2586 269 2587
rect 338 2587 344 2588
rect 338 2586 339 2587
rect 268 2584 339 2586
rect 268 2583 269 2584
rect 263 2582 269 2583
rect 338 2583 339 2584
rect 343 2583 344 2587
rect 338 2582 344 2583
rect 407 2587 413 2588
rect 407 2583 408 2587
rect 412 2586 413 2587
rect 422 2587 428 2588
rect 422 2586 423 2587
rect 412 2584 423 2586
rect 412 2583 413 2584
rect 407 2582 413 2583
rect 422 2583 423 2584
rect 427 2583 428 2587
rect 422 2582 428 2583
rect 543 2587 549 2588
rect 543 2583 544 2587
rect 548 2586 549 2587
rect 650 2587 656 2588
rect 650 2586 651 2587
rect 548 2584 651 2586
rect 548 2583 549 2584
rect 543 2582 549 2583
rect 650 2583 651 2584
rect 655 2583 656 2587
rect 650 2582 656 2583
rect 662 2587 668 2588
rect 662 2583 663 2587
rect 667 2586 668 2587
rect 671 2587 677 2588
rect 671 2586 672 2587
rect 667 2584 672 2586
rect 667 2583 668 2584
rect 662 2582 668 2583
rect 671 2583 672 2584
rect 676 2583 677 2587
rect 671 2582 677 2583
rect 799 2587 805 2588
rect 799 2583 800 2587
rect 804 2586 805 2587
rect 814 2587 820 2588
rect 814 2586 815 2587
rect 804 2584 815 2586
rect 804 2583 805 2584
rect 799 2582 805 2583
rect 814 2583 815 2584
rect 819 2583 820 2587
rect 814 2582 820 2583
rect 919 2587 925 2588
rect 919 2583 920 2587
rect 924 2586 925 2587
rect 994 2587 1000 2588
rect 994 2586 995 2587
rect 924 2584 995 2586
rect 924 2583 925 2584
rect 919 2582 925 2583
rect 994 2583 995 2584
rect 999 2583 1000 2587
rect 994 2582 1000 2583
rect 1039 2587 1045 2588
rect 1039 2583 1040 2587
rect 1044 2586 1045 2587
rect 1118 2587 1124 2588
rect 1118 2586 1119 2587
rect 1044 2584 1119 2586
rect 1044 2583 1045 2584
rect 1039 2582 1045 2583
rect 1118 2583 1119 2584
rect 1123 2583 1124 2587
rect 1118 2582 1124 2583
rect 1167 2587 1173 2588
rect 1167 2583 1168 2587
rect 1172 2586 1173 2587
rect 1274 2587 1280 2588
rect 1274 2586 1275 2587
rect 1172 2584 1275 2586
rect 1172 2583 1173 2584
rect 1167 2582 1173 2583
rect 1274 2583 1275 2584
rect 1279 2583 1280 2587
rect 1274 2582 1280 2583
rect 2486 2587 2492 2588
rect 2486 2583 2487 2587
rect 2491 2586 2492 2587
rect 2495 2587 2501 2588
rect 2495 2586 2496 2587
rect 2491 2584 2496 2586
rect 2491 2583 2492 2584
rect 2486 2582 2492 2583
rect 2495 2583 2496 2584
rect 2500 2583 2501 2587
rect 2495 2582 2501 2583
rect 142 2577 148 2578
rect 142 2573 143 2577
rect 147 2573 148 2577
rect 142 2572 148 2573
rect 270 2577 276 2578
rect 270 2573 271 2577
rect 275 2573 276 2577
rect 270 2572 276 2573
rect 414 2577 420 2578
rect 414 2573 415 2577
rect 419 2573 420 2577
rect 414 2572 420 2573
rect 550 2577 556 2578
rect 550 2573 551 2577
rect 555 2573 556 2577
rect 550 2572 556 2573
rect 678 2577 684 2578
rect 678 2573 679 2577
rect 683 2573 684 2577
rect 678 2572 684 2573
rect 806 2577 812 2578
rect 806 2573 807 2577
rect 811 2573 812 2577
rect 806 2572 812 2573
rect 926 2577 932 2578
rect 926 2573 927 2577
rect 931 2573 932 2577
rect 926 2572 932 2573
rect 1046 2577 1052 2578
rect 1046 2573 1047 2577
rect 1051 2573 1052 2577
rect 1046 2572 1052 2573
rect 1174 2577 1180 2578
rect 1174 2573 1175 2577
rect 1179 2573 1180 2577
rect 1174 2572 1180 2573
rect 1886 2567 1892 2568
rect 110 2564 116 2565
rect 1822 2564 1828 2565
rect 110 2560 111 2564
rect 115 2560 116 2564
rect 618 2563 624 2564
rect 618 2562 619 2563
rect 605 2560 619 2562
rect 110 2559 116 2560
rect 210 2559 216 2560
rect 210 2555 211 2559
rect 215 2558 216 2559
rect 338 2559 344 2560
rect 215 2556 289 2558
rect 215 2555 216 2556
rect 210 2554 216 2555
rect 338 2555 339 2559
rect 343 2558 344 2559
rect 618 2559 619 2560
rect 623 2559 624 2563
rect 1822 2560 1823 2564
rect 1827 2560 1828 2564
rect 1886 2563 1887 2567
rect 1891 2563 1892 2567
rect 1886 2562 1892 2563
rect 1990 2567 1996 2568
rect 1990 2563 1991 2567
rect 1995 2563 1996 2567
rect 1990 2562 1996 2563
rect 2110 2567 2116 2568
rect 2110 2563 2111 2567
rect 2115 2563 2116 2567
rect 2110 2562 2116 2563
rect 2230 2567 2236 2568
rect 2230 2563 2231 2567
rect 2235 2563 2236 2567
rect 2230 2562 2236 2563
rect 2350 2567 2356 2568
rect 2350 2563 2351 2567
rect 2355 2563 2356 2567
rect 2350 2562 2356 2563
rect 2470 2567 2476 2568
rect 2470 2563 2471 2567
rect 2475 2563 2476 2567
rect 2470 2562 2476 2563
rect 2590 2567 2596 2568
rect 2590 2563 2591 2567
rect 2595 2563 2596 2567
rect 2590 2562 2596 2563
rect 2710 2567 2716 2568
rect 2710 2563 2711 2567
rect 2715 2563 2716 2567
rect 2710 2562 2716 2563
rect 2830 2567 2836 2568
rect 2830 2563 2831 2567
rect 2835 2563 2836 2567
rect 2830 2562 2836 2563
rect 618 2558 624 2559
rect 650 2559 656 2560
rect 343 2556 433 2558
rect 343 2555 344 2556
rect 338 2554 344 2555
rect 650 2555 651 2559
rect 655 2558 656 2559
rect 746 2559 752 2560
rect 655 2556 697 2558
rect 655 2555 656 2556
rect 650 2554 656 2555
rect 746 2555 747 2559
rect 751 2558 752 2559
rect 994 2559 1000 2560
rect 751 2556 825 2558
rect 751 2555 752 2556
rect 746 2554 752 2555
rect 994 2555 995 2559
rect 999 2558 1000 2559
rect 1118 2559 1124 2560
rect 1822 2559 1828 2560
rect 2103 2559 2109 2560
rect 999 2556 1065 2558
rect 999 2555 1000 2556
rect 994 2554 1000 2555
rect 1118 2555 1119 2559
rect 1123 2558 1124 2559
rect 1123 2556 1193 2558
rect 1862 2557 1868 2558
rect 1123 2555 1124 2556
rect 1118 2554 1124 2555
rect 1862 2553 1863 2557
rect 1867 2553 1868 2557
rect 2103 2555 2104 2559
rect 2108 2558 2109 2559
rect 2778 2559 2784 2560
rect 2108 2556 2129 2558
rect 2108 2555 2109 2556
rect 2103 2554 2109 2555
rect 2778 2555 2779 2559
rect 2783 2558 2784 2559
rect 2783 2556 2849 2558
rect 3574 2557 3580 2558
rect 2783 2555 2784 2556
rect 2778 2554 2784 2555
rect 1862 2552 1868 2553
rect 3574 2553 3575 2557
rect 3579 2553 3580 2557
rect 3574 2552 3580 2553
rect 110 2547 116 2548
rect 110 2543 111 2547
rect 115 2543 116 2547
rect 110 2542 116 2543
rect 127 2547 133 2548
rect 127 2543 128 2547
rect 132 2546 133 2547
rect 886 2547 892 2548
rect 132 2544 153 2546
rect 132 2543 133 2544
rect 127 2542 133 2543
rect 886 2543 887 2547
rect 891 2546 892 2547
rect 1822 2547 1828 2548
rect 891 2544 937 2546
rect 891 2543 892 2544
rect 886 2542 892 2543
rect 1822 2543 1823 2547
rect 1827 2543 1828 2547
rect 1822 2542 1828 2543
rect 1879 2543 1885 2544
rect 1862 2540 1868 2541
rect 134 2537 140 2538
rect 134 2533 135 2537
rect 139 2533 140 2537
rect 134 2532 140 2533
rect 262 2537 268 2538
rect 262 2533 263 2537
rect 267 2533 268 2537
rect 262 2532 268 2533
rect 406 2537 412 2538
rect 406 2533 407 2537
rect 411 2533 412 2537
rect 406 2532 412 2533
rect 542 2537 548 2538
rect 542 2533 543 2537
rect 547 2533 548 2537
rect 542 2532 548 2533
rect 670 2537 676 2538
rect 670 2533 671 2537
rect 675 2533 676 2537
rect 670 2532 676 2533
rect 798 2537 804 2538
rect 798 2533 799 2537
rect 803 2533 804 2537
rect 798 2532 804 2533
rect 918 2537 924 2538
rect 918 2533 919 2537
rect 923 2533 924 2537
rect 918 2532 924 2533
rect 1038 2537 1044 2538
rect 1038 2533 1039 2537
rect 1043 2533 1044 2537
rect 1038 2532 1044 2533
rect 1166 2537 1172 2538
rect 1166 2533 1167 2537
rect 1171 2533 1172 2537
rect 1862 2536 1863 2540
rect 1867 2536 1868 2540
rect 1879 2539 1880 2543
rect 1884 2542 1885 2543
rect 1954 2543 1960 2544
rect 1884 2540 1913 2542
rect 1884 2539 1885 2540
rect 1879 2538 1885 2539
rect 1954 2539 1955 2543
rect 1959 2542 1960 2543
rect 2178 2543 2184 2544
rect 1959 2540 2017 2542
rect 1959 2539 1960 2540
rect 1954 2538 1960 2539
rect 2178 2539 2179 2543
rect 2183 2542 2184 2543
rect 2326 2543 2332 2544
rect 2183 2540 2257 2542
rect 2183 2539 2184 2540
rect 2178 2538 2184 2539
rect 2326 2539 2327 2543
rect 2331 2542 2332 2543
rect 2583 2543 2589 2544
rect 2583 2542 2584 2543
rect 2331 2540 2377 2542
rect 2533 2540 2584 2542
rect 2331 2539 2332 2540
rect 2326 2538 2332 2539
rect 2583 2539 2584 2540
rect 2588 2539 2589 2543
rect 2703 2543 2709 2544
rect 2703 2542 2704 2543
rect 2653 2540 2704 2542
rect 2583 2538 2589 2539
rect 2703 2539 2704 2540
rect 2708 2539 2709 2543
rect 2823 2543 2829 2544
rect 2823 2542 2824 2543
rect 2773 2540 2824 2542
rect 2703 2538 2709 2539
rect 2823 2539 2824 2540
rect 2828 2539 2829 2543
rect 2823 2538 2829 2539
rect 3574 2540 3580 2541
rect 1862 2535 1868 2536
rect 3574 2536 3575 2540
rect 3579 2536 3580 2540
rect 3574 2535 3580 2536
rect 1166 2532 1172 2533
rect 1894 2527 1900 2528
rect 1894 2523 1895 2527
rect 1899 2523 1900 2527
rect 1894 2522 1900 2523
rect 1998 2527 2004 2528
rect 1998 2523 1999 2527
rect 2003 2523 2004 2527
rect 1998 2522 2004 2523
rect 2118 2527 2124 2528
rect 2118 2523 2119 2527
rect 2123 2523 2124 2527
rect 2118 2522 2124 2523
rect 2238 2527 2244 2528
rect 2238 2523 2239 2527
rect 2243 2523 2244 2527
rect 2238 2522 2244 2523
rect 2358 2527 2364 2528
rect 2358 2523 2359 2527
rect 2363 2523 2364 2527
rect 2358 2522 2364 2523
rect 2478 2527 2484 2528
rect 2478 2523 2479 2527
rect 2483 2523 2484 2527
rect 2478 2522 2484 2523
rect 2598 2527 2604 2528
rect 2598 2523 2599 2527
rect 2603 2523 2604 2527
rect 2598 2522 2604 2523
rect 2718 2527 2724 2528
rect 2718 2523 2719 2527
rect 2723 2523 2724 2527
rect 2718 2522 2724 2523
rect 2838 2527 2844 2528
rect 2838 2523 2839 2527
rect 2843 2523 2844 2527
rect 2838 2522 2844 2523
rect 134 2515 140 2516
rect 134 2511 135 2515
rect 139 2511 140 2515
rect 134 2510 140 2511
rect 278 2515 284 2516
rect 278 2511 279 2515
rect 283 2511 284 2515
rect 278 2510 284 2511
rect 438 2515 444 2516
rect 438 2511 439 2515
rect 443 2511 444 2515
rect 438 2510 444 2511
rect 590 2515 596 2516
rect 590 2511 591 2515
rect 595 2511 596 2515
rect 590 2510 596 2511
rect 734 2515 740 2516
rect 734 2511 735 2515
rect 739 2511 740 2515
rect 734 2510 740 2511
rect 870 2515 876 2516
rect 870 2511 871 2515
rect 875 2511 876 2515
rect 870 2510 876 2511
rect 1006 2515 1012 2516
rect 1006 2511 1007 2515
rect 1011 2511 1012 2515
rect 1006 2510 1012 2511
rect 1142 2515 1148 2516
rect 1142 2511 1143 2515
rect 1147 2511 1148 2515
rect 1142 2510 1148 2511
rect 1278 2515 1284 2516
rect 1278 2511 1279 2515
rect 1283 2511 1284 2515
rect 1278 2510 1284 2511
rect 1887 2515 1893 2516
rect 1887 2511 1888 2515
rect 1892 2514 1893 2515
rect 1954 2515 1960 2516
rect 1954 2514 1955 2515
rect 1892 2512 1955 2514
rect 1892 2511 1893 2512
rect 1887 2510 1893 2511
rect 1954 2511 1955 2512
rect 1959 2511 1960 2515
rect 1954 2510 1960 2511
rect 1983 2515 1989 2516
rect 1983 2511 1984 2515
rect 1988 2514 1989 2515
rect 1991 2515 1997 2516
rect 1991 2514 1992 2515
rect 1988 2512 1992 2514
rect 1988 2511 1989 2512
rect 1983 2510 1989 2511
rect 1991 2511 1992 2512
rect 1996 2511 1997 2515
rect 1991 2510 1997 2511
rect 2111 2515 2117 2516
rect 2111 2511 2112 2515
rect 2116 2514 2117 2515
rect 2178 2515 2184 2516
rect 2178 2514 2179 2515
rect 2116 2512 2179 2514
rect 2116 2511 2117 2512
rect 2111 2510 2117 2511
rect 2178 2511 2179 2512
rect 2183 2511 2184 2515
rect 2178 2510 2184 2511
rect 2231 2515 2237 2516
rect 2231 2511 2232 2515
rect 2236 2514 2237 2515
rect 2326 2515 2332 2516
rect 2326 2514 2327 2515
rect 2236 2512 2327 2514
rect 2236 2511 2237 2512
rect 2231 2510 2237 2511
rect 2326 2511 2327 2512
rect 2331 2511 2332 2515
rect 2326 2510 2332 2511
rect 2334 2515 2340 2516
rect 2334 2511 2335 2515
rect 2339 2514 2340 2515
rect 2351 2515 2357 2516
rect 2351 2514 2352 2515
rect 2339 2512 2352 2514
rect 2339 2511 2340 2512
rect 2334 2510 2340 2511
rect 2351 2511 2352 2512
rect 2356 2511 2357 2515
rect 2351 2510 2357 2511
rect 2471 2515 2477 2516
rect 2471 2511 2472 2515
rect 2476 2514 2477 2515
rect 2486 2515 2492 2516
rect 2486 2514 2487 2515
rect 2476 2512 2487 2514
rect 2476 2511 2477 2512
rect 2471 2510 2477 2511
rect 2486 2511 2487 2512
rect 2491 2511 2492 2515
rect 2486 2510 2492 2511
rect 2583 2515 2589 2516
rect 2583 2511 2584 2515
rect 2588 2514 2589 2515
rect 2591 2515 2597 2516
rect 2591 2514 2592 2515
rect 2588 2512 2592 2514
rect 2588 2511 2589 2512
rect 2583 2510 2589 2511
rect 2591 2511 2592 2512
rect 2596 2511 2597 2515
rect 2591 2510 2597 2511
rect 2703 2515 2709 2516
rect 2703 2511 2704 2515
rect 2708 2514 2709 2515
rect 2711 2515 2717 2516
rect 2711 2514 2712 2515
rect 2708 2512 2712 2514
rect 2708 2511 2709 2512
rect 2703 2510 2709 2511
rect 2711 2511 2712 2512
rect 2716 2511 2717 2515
rect 2711 2510 2717 2511
rect 2823 2515 2829 2516
rect 2823 2511 2824 2515
rect 2828 2514 2829 2515
rect 2831 2515 2837 2516
rect 2831 2514 2832 2515
rect 2828 2512 2832 2514
rect 2828 2511 2829 2512
rect 2823 2510 2829 2511
rect 2831 2511 2832 2512
rect 2836 2511 2837 2515
rect 2831 2510 2837 2511
rect 662 2507 668 2508
rect 662 2506 663 2507
rect 110 2505 116 2506
rect 110 2501 111 2505
rect 115 2501 116 2505
rect 649 2504 663 2506
rect 662 2503 663 2504
rect 667 2503 668 2507
rect 814 2507 820 2508
rect 814 2506 815 2507
rect 793 2504 815 2506
rect 662 2502 668 2503
rect 814 2503 815 2504
rect 819 2503 820 2507
rect 814 2502 820 2503
rect 1218 2507 1224 2508
rect 1218 2503 1219 2507
rect 1223 2506 1224 2507
rect 1223 2504 1297 2506
rect 1822 2505 1828 2506
rect 1223 2503 1224 2504
rect 1218 2502 1224 2503
rect 110 2500 116 2501
rect 1822 2501 1823 2505
rect 1827 2501 1828 2505
rect 1822 2500 1828 2501
rect 1879 2499 1885 2500
rect 1879 2495 1880 2499
rect 1884 2498 1885 2499
rect 1887 2499 1893 2500
rect 1887 2498 1888 2499
rect 1884 2496 1888 2498
rect 1884 2495 1885 2496
rect 1879 2494 1885 2495
rect 1887 2495 1888 2496
rect 1892 2495 1893 2499
rect 1887 2494 1893 2495
rect 1959 2499 1965 2500
rect 1959 2495 1960 2499
rect 1964 2498 1965 2499
rect 2023 2499 2029 2500
rect 2023 2498 2024 2499
rect 1964 2496 2024 2498
rect 1964 2495 1965 2496
rect 1959 2494 1965 2495
rect 2023 2495 2024 2496
rect 2028 2495 2029 2499
rect 2023 2494 2029 2495
rect 2167 2499 2173 2500
rect 2167 2495 2168 2499
rect 2172 2498 2173 2499
rect 2183 2499 2189 2500
rect 2183 2498 2184 2499
rect 2172 2496 2184 2498
rect 2172 2495 2173 2496
rect 2167 2494 2173 2495
rect 2183 2495 2184 2496
rect 2188 2495 2189 2499
rect 2183 2494 2189 2495
rect 2255 2499 2261 2500
rect 2255 2495 2256 2499
rect 2260 2498 2261 2499
rect 2335 2499 2341 2500
rect 2335 2498 2336 2499
rect 2260 2496 2336 2498
rect 2260 2495 2261 2496
rect 2255 2494 2261 2495
rect 2335 2495 2336 2496
rect 2340 2495 2341 2499
rect 2335 2494 2341 2495
rect 2479 2499 2485 2500
rect 2479 2495 2480 2499
rect 2484 2498 2485 2499
rect 2494 2499 2500 2500
rect 2494 2498 2495 2499
rect 2484 2496 2495 2498
rect 2484 2495 2485 2496
rect 2479 2494 2485 2495
rect 2494 2495 2495 2496
rect 2499 2495 2500 2499
rect 2494 2494 2500 2495
rect 2551 2499 2557 2500
rect 2551 2495 2552 2499
rect 2556 2498 2557 2499
rect 2615 2499 2621 2500
rect 2615 2498 2616 2499
rect 2556 2496 2616 2498
rect 2556 2495 2557 2496
rect 2551 2494 2557 2495
rect 2615 2495 2616 2496
rect 2620 2495 2621 2499
rect 2615 2494 2621 2495
rect 2687 2499 2693 2500
rect 2687 2495 2688 2499
rect 2692 2498 2693 2499
rect 2743 2499 2749 2500
rect 2743 2498 2744 2499
rect 2692 2496 2744 2498
rect 2692 2495 2693 2496
rect 2687 2494 2693 2495
rect 2743 2495 2744 2496
rect 2748 2495 2749 2499
rect 2743 2494 2749 2495
rect 2815 2499 2821 2500
rect 2815 2495 2816 2499
rect 2820 2498 2821 2499
rect 2871 2499 2877 2500
rect 2871 2498 2872 2499
rect 2820 2496 2872 2498
rect 2820 2495 2821 2496
rect 2815 2494 2821 2495
rect 2871 2495 2872 2496
rect 2876 2495 2877 2499
rect 2871 2494 2877 2495
rect 2943 2499 2949 2500
rect 2943 2495 2944 2499
rect 2948 2498 2949 2499
rect 3007 2499 3013 2500
rect 3007 2498 3008 2499
rect 2948 2496 3008 2498
rect 2948 2495 2949 2496
rect 2943 2494 2949 2495
rect 3007 2495 3008 2496
rect 3012 2495 3013 2499
rect 3007 2494 3013 2495
rect 271 2491 277 2492
rect 271 2490 272 2491
rect 110 2488 116 2489
rect 197 2488 272 2490
rect 110 2484 111 2488
rect 115 2484 116 2488
rect 271 2487 272 2488
rect 276 2487 277 2491
rect 423 2491 429 2492
rect 423 2490 424 2491
rect 341 2488 424 2490
rect 271 2486 277 2487
rect 423 2487 424 2488
rect 428 2487 429 2491
rect 423 2486 429 2487
rect 431 2491 437 2492
rect 431 2487 432 2491
rect 436 2490 437 2491
rect 999 2491 1005 2492
rect 999 2490 1000 2491
rect 436 2488 465 2490
rect 933 2488 1000 2490
rect 436 2487 437 2488
rect 431 2486 437 2487
rect 999 2487 1000 2488
rect 1004 2487 1005 2491
rect 1135 2491 1141 2492
rect 1135 2490 1136 2491
rect 1069 2488 1136 2490
rect 999 2486 1005 2487
rect 1135 2487 1136 2488
rect 1140 2487 1141 2491
rect 1271 2491 1277 2492
rect 1271 2490 1272 2491
rect 1205 2488 1272 2490
rect 1135 2486 1141 2487
rect 1271 2487 1272 2488
rect 1276 2487 1277 2491
rect 1894 2489 1900 2490
rect 1271 2486 1277 2487
rect 1822 2488 1828 2489
rect 110 2483 116 2484
rect 1822 2484 1823 2488
rect 1827 2484 1828 2488
rect 1894 2485 1895 2489
rect 1899 2485 1900 2489
rect 1894 2484 1900 2485
rect 2030 2489 2036 2490
rect 2030 2485 2031 2489
rect 2035 2485 2036 2489
rect 2030 2484 2036 2485
rect 2190 2489 2196 2490
rect 2190 2485 2191 2489
rect 2195 2485 2196 2489
rect 2190 2484 2196 2485
rect 2342 2489 2348 2490
rect 2342 2485 2343 2489
rect 2347 2485 2348 2489
rect 2342 2484 2348 2485
rect 2486 2489 2492 2490
rect 2486 2485 2487 2489
rect 2491 2485 2492 2489
rect 2486 2484 2492 2485
rect 2622 2489 2628 2490
rect 2622 2485 2623 2489
rect 2627 2485 2628 2489
rect 2622 2484 2628 2485
rect 2750 2489 2756 2490
rect 2750 2485 2751 2489
rect 2755 2485 2756 2489
rect 2750 2484 2756 2485
rect 2878 2489 2884 2490
rect 2878 2485 2879 2489
rect 2883 2485 2884 2489
rect 2878 2484 2884 2485
rect 3014 2489 3020 2490
rect 3014 2485 3015 2489
rect 3019 2485 3020 2489
rect 3014 2484 3020 2485
rect 1822 2483 1828 2484
rect 1862 2476 1868 2477
rect 3574 2476 3580 2477
rect 142 2475 148 2476
rect 142 2471 143 2475
rect 147 2471 148 2475
rect 142 2470 148 2471
rect 286 2475 292 2476
rect 286 2471 287 2475
rect 291 2471 292 2475
rect 286 2470 292 2471
rect 446 2475 452 2476
rect 446 2471 447 2475
rect 451 2471 452 2475
rect 446 2470 452 2471
rect 598 2475 604 2476
rect 598 2471 599 2475
rect 603 2471 604 2475
rect 598 2470 604 2471
rect 742 2475 748 2476
rect 742 2471 743 2475
rect 747 2471 748 2475
rect 742 2470 748 2471
rect 878 2475 884 2476
rect 878 2471 879 2475
rect 883 2471 884 2475
rect 878 2470 884 2471
rect 1014 2475 1020 2476
rect 1014 2471 1015 2475
rect 1019 2471 1020 2475
rect 1014 2470 1020 2471
rect 1150 2475 1156 2476
rect 1150 2471 1151 2475
rect 1155 2471 1156 2475
rect 1150 2470 1156 2471
rect 1286 2475 1292 2476
rect 1286 2471 1287 2475
rect 1291 2471 1292 2475
rect 1862 2472 1863 2476
rect 1867 2472 1868 2476
rect 1959 2475 1965 2476
rect 1959 2474 1960 2475
rect 1949 2472 1960 2474
rect 1862 2471 1868 2472
rect 1959 2471 1960 2472
rect 1964 2471 1965 2475
rect 2255 2475 2261 2476
rect 2255 2474 2256 2475
rect 2245 2472 2256 2474
rect 1286 2470 1292 2471
rect 1959 2470 1965 2471
rect 2255 2471 2256 2472
rect 2260 2471 2261 2475
rect 2551 2475 2557 2476
rect 2551 2474 2552 2475
rect 2541 2472 2552 2474
rect 2255 2470 2261 2471
rect 2334 2471 2340 2472
rect 2334 2467 2335 2471
rect 2339 2470 2340 2471
rect 2551 2471 2552 2472
rect 2556 2471 2557 2475
rect 2687 2475 2693 2476
rect 2687 2474 2688 2475
rect 2677 2472 2688 2474
rect 2551 2470 2557 2471
rect 2687 2471 2688 2472
rect 2692 2471 2693 2475
rect 2815 2475 2821 2476
rect 2815 2474 2816 2475
rect 2805 2472 2816 2474
rect 2687 2470 2693 2471
rect 2815 2471 2816 2472
rect 2820 2471 2821 2475
rect 2943 2475 2949 2476
rect 2943 2474 2944 2475
rect 2933 2472 2944 2474
rect 2815 2470 2821 2471
rect 2943 2471 2944 2472
rect 2948 2471 2949 2475
rect 3574 2472 3575 2476
rect 3579 2472 3580 2476
rect 3574 2471 3580 2472
rect 2943 2470 2949 2471
rect 2339 2468 2361 2470
rect 2339 2467 2340 2468
rect 2334 2466 2340 2467
rect 127 2463 133 2464
rect 127 2459 128 2463
rect 132 2462 133 2463
rect 135 2463 141 2464
rect 135 2462 136 2463
rect 132 2460 136 2462
rect 132 2459 133 2460
rect 127 2458 133 2459
rect 135 2459 136 2460
rect 140 2459 141 2463
rect 135 2458 141 2459
rect 271 2463 277 2464
rect 271 2459 272 2463
rect 276 2462 277 2463
rect 279 2463 285 2464
rect 279 2462 280 2463
rect 276 2460 280 2462
rect 276 2459 277 2460
rect 271 2458 277 2459
rect 279 2459 280 2460
rect 284 2459 285 2463
rect 279 2458 285 2459
rect 423 2463 429 2464
rect 423 2459 424 2463
rect 428 2462 429 2463
rect 439 2463 445 2464
rect 439 2462 440 2463
rect 428 2460 440 2462
rect 428 2459 429 2460
rect 423 2458 429 2459
rect 439 2459 440 2460
rect 444 2459 445 2463
rect 439 2458 445 2459
rect 582 2463 588 2464
rect 582 2459 583 2463
rect 587 2462 588 2463
rect 591 2463 597 2464
rect 591 2462 592 2463
rect 587 2460 592 2462
rect 587 2459 588 2460
rect 582 2458 588 2459
rect 591 2459 592 2460
rect 596 2459 597 2463
rect 591 2458 597 2459
rect 735 2463 741 2464
rect 735 2459 736 2463
rect 740 2462 741 2463
rect 794 2463 800 2464
rect 794 2462 795 2463
rect 740 2460 795 2462
rect 740 2459 741 2460
rect 735 2458 741 2459
rect 794 2459 795 2460
rect 799 2459 800 2463
rect 794 2458 800 2459
rect 871 2463 877 2464
rect 871 2459 872 2463
rect 876 2462 877 2463
rect 886 2463 892 2464
rect 886 2462 887 2463
rect 876 2460 887 2462
rect 876 2459 877 2460
rect 871 2458 877 2459
rect 886 2459 887 2460
rect 891 2459 892 2463
rect 886 2458 892 2459
rect 999 2463 1005 2464
rect 999 2459 1000 2463
rect 1004 2462 1005 2463
rect 1007 2463 1013 2464
rect 1007 2462 1008 2463
rect 1004 2460 1008 2462
rect 1004 2459 1005 2460
rect 999 2458 1005 2459
rect 1007 2459 1008 2460
rect 1012 2459 1013 2463
rect 1007 2458 1013 2459
rect 1135 2463 1141 2464
rect 1135 2459 1136 2463
rect 1140 2462 1141 2463
rect 1143 2463 1149 2464
rect 1143 2462 1144 2463
rect 1140 2460 1144 2462
rect 1140 2459 1141 2460
rect 1135 2458 1141 2459
rect 1143 2459 1144 2460
rect 1148 2459 1149 2463
rect 1143 2458 1149 2459
rect 1271 2463 1277 2464
rect 1271 2459 1272 2463
rect 1276 2462 1277 2463
rect 1279 2463 1285 2464
rect 1279 2462 1280 2463
rect 1276 2460 1280 2462
rect 1276 2459 1277 2460
rect 1271 2458 1277 2459
rect 1279 2459 1280 2460
rect 1284 2459 1285 2463
rect 1279 2458 1285 2459
rect 1862 2459 1868 2460
rect 1862 2455 1863 2459
rect 1867 2455 1868 2459
rect 1862 2454 1868 2455
rect 2030 2459 2036 2460
rect 2030 2455 2031 2459
rect 2035 2458 2036 2459
rect 2966 2459 2972 2460
rect 2035 2456 2041 2458
rect 2035 2455 2036 2456
rect 2030 2454 2036 2455
rect 2966 2455 2967 2459
rect 2971 2458 2972 2459
rect 3574 2459 3580 2460
rect 2971 2456 3025 2458
rect 2971 2455 2972 2456
rect 2966 2454 2972 2455
rect 3574 2455 3575 2459
rect 3579 2455 3580 2459
rect 3574 2454 3580 2455
rect 183 2451 189 2452
rect 183 2447 184 2451
rect 188 2450 189 2451
rect 258 2451 264 2452
rect 258 2450 259 2451
rect 188 2448 259 2450
rect 188 2447 189 2448
rect 183 2446 189 2447
rect 258 2447 259 2448
rect 263 2447 264 2451
rect 258 2446 264 2447
rect 311 2451 317 2452
rect 311 2447 312 2451
rect 316 2450 317 2451
rect 390 2451 396 2452
rect 390 2450 391 2451
rect 316 2448 391 2450
rect 316 2447 317 2448
rect 311 2446 317 2447
rect 390 2447 391 2448
rect 395 2447 396 2451
rect 390 2446 396 2447
rect 431 2451 437 2452
rect 431 2447 432 2451
rect 436 2450 437 2451
rect 447 2451 453 2452
rect 447 2450 448 2451
rect 436 2448 448 2450
rect 436 2447 437 2448
rect 431 2446 437 2447
rect 447 2447 448 2448
rect 452 2447 453 2451
rect 447 2446 453 2447
rect 583 2451 589 2452
rect 583 2447 584 2451
rect 588 2450 589 2451
rect 678 2451 684 2452
rect 678 2450 679 2451
rect 588 2448 679 2450
rect 588 2447 589 2448
rect 583 2446 589 2447
rect 678 2447 679 2448
rect 683 2447 684 2451
rect 678 2446 684 2447
rect 719 2451 725 2452
rect 719 2447 720 2451
rect 724 2450 725 2451
rect 766 2451 772 2452
rect 766 2450 767 2451
rect 724 2448 767 2450
rect 724 2447 725 2448
rect 719 2446 725 2447
rect 766 2447 767 2448
rect 771 2447 772 2451
rect 766 2446 772 2447
rect 855 2451 861 2452
rect 855 2447 856 2451
rect 860 2450 861 2451
rect 886 2451 892 2452
rect 886 2450 887 2451
rect 860 2448 887 2450
rect 860 2447 861 2448
rect 855 2446 861 2447
rect 886 2447 887 2448
rect 891 2447 892 2451
rect 886 2446 892 2447
rect 991 2451 997 2452
rect 991 2447 992 2451
rect 996 2450 997 2451
rect 1006 2451 1012 2452
rect 1006 2450 1007 2451
rect 996 2448 1007 2450
rect 996 2447 997 2448
rect 991 2446 997 2447
rect 1006 2447 1007 2448
rect 1011 2447 1012 2451
rect 1006 2446 1012 2447
rect 1063 2451 1069 2452
rect 1063 2447 1064 2451
rect 1068 2450 1069 2451
rect 1127 2451 1133 2452
rect 1127 2450 1128 2451
rect 1068 2448 1128 2450
rect 1068 2447 1069 2448
rect 1063 2446 1069 2447
rect 1127 2447 1128 2448
rect 1132 2447 1133 2451
rect 1127 2446 1133 2447
rect 1199 2451 1205 2452
rect 1199 2447 1200 2451
rect 1204 2450 1205 2451
rect 1263 2451 1269 2452
rect 1263 2450 1264 2451
rect 1204 2448 1264 2450
rect 1204 2447 1205 2448
rect 1199 2446 1205 2447
rect 1263 2447 1264 2448
rect 1268 2447 1269 2451
rect 1263 2446 1269 2447
rect 1335 2451 1341 2452
rect 1335 2447 1336 2451
rect 1340 2450 1341 2451
rect 1399 2451 1405 2452
rect 1399 2450 1400 2451
rect 1340 2448 1400 2450
rect 1340 2447 1341 2448
rect 1335 2446 1341 2447
rect 1399 2447 1400 2448
rect 1404 2447 1405 2451
rect 1399 2446 1405 2447
rect 1886 2449 1892 2450
rect 1886 2445 1887 2449
rect 1891 2445 1892 2449
rect 1886 2444 1892 2445
rect 2022 2449 2028 2450
rect 2022 2445 2023 2449
rect 2027 2445 2028 2449
rect 2022 2444 2028 2445
rect 2182 2449 2188 2450
rect 2182 2445 2183 2449
rect 2187 2445 2188 2449
rect 2182 2444 2188 2445
rect 2334 2449 2340 2450
rect 2334 2445 2335 2449
rect 2339 2445 2340 2449
rect 2334 2444 2340 2445
rect 2478 2449 2484 2450
rect 2478 2445 2479 2449
rect 2483 2445 2484 2449
rect 2478 2444 2484 2445
rect 2614 2449 2620 2450
rect 2614 2445 2615 2449
rect 2619 2445 2620 2449
rect 2614 2444 2620 2445
rect 2742 2449 2748 2450
rect 2742 2445 2743 2449
rect 2747 2445 2748 2449
rect 2742 2444 2748 2445
rect 2870 2449 2876 2450
rect 2870 2445 2871 2449
rect 2875 2445 2876 2449
rect 2870 2444 2876 2445
rect 3006 2449 3012 2450
rect 3006 2445 3007 2449
rect 3011 2445 3012 2449
rect 3006 2444 3012 2445
rect 190 2441 196 2442
rect 190 2437 191 2441
rect 195 2437 196 2441
rect 190 2436 196 2437
rect 318 2441 324 2442
rect 318 2437 319 2441
rect 323 2437 324 2441
rect 318 2436 324 2437
rect 454 2441 460 2442
rect 454 2437 455 2441
rect 459 2437 460 2441
rect 454 2436 460 2437
rect 590 2441 596 2442
rect 590 2437 591 2441
rect 595 2437 596 2441
rect 590 2436 596 2437
rect 726 2441 732 2442
rect 726 2437 727 2441
rect 731 2437 732 2441
rect 726 2436 732 2437
rect 862 2441 868 2442
rect 862 2437 863 2441
rect 867 2437 868 2441
rect 862 2436 868 2437
rect 998 2441 1004 2442
rect 998 2437 999 2441
rect 1003 2437 1004 2441
rect 998 2436 1004 2437
rect 1134 2441 1140 2442
rect 1134 2437 1135 2441
rect 1139 2437 1140 2441
rect 1134 2436 1140 2437
rect 1270 2441 1276 2442
rect 1270 2437 1271 2441
rect 1275 2437 1276 2441
rect 1270 2436 1276 2437
rect 1406 2441 1412 2442
rect 1406 2437 1407 2441
rect 1411 2437 1412 2441
rect 1406 2436 1412 2437
rect 110 2428 116 2429
rect 1822 2428 1828 2429
rect 110 2424 111 2428
rect 115 2424 116 2428
rect 1063 2427 1069 2428
rect 1063 2426 1064 2427
rect 1053 2424 1064 2426
rect 110 2423 116 2424
rect 258 2423 264 2424
rect 258 2419 259 2423
rect 263 2422 264 2423
rect 390 2423 396 2424
rect 263 2420 337 2422
rect 263 2419 264 2420
rect 258 2418 264 2419
rect 390 2419 391 2423
rect 395 2422 396 2423
rect 582 2423 588 2424
rect 395 2420 473 2422
rect 395 2419 396 2420
rect 390 2418 396 2419
rect 582 2419 583 2423
rect 587 2422 588 2423
rect 678 2423 684 2424
rect 587 2420 609 2422
rect 587 2419 588 2420
rect 582 2418 588 2419
rect 678 2419 679 2423
rect 683 2422 684 2423
rect 794 2423 800 2424
rect 683 2420 745 2422
rect 683 2419 684 2420
rect 678 2418 684 2419
rect 794 2419 795 2423
rect 799 2422 800 2423
rect 1063 2423 1064 2424
rect 1068 2423 1069 2427
rect 1199 2427 1205 2428
rect 1199 2426 1200 2427
rect 1189 2424 1200 2426
rect 1063 2422 1069 2423
rect 1199 2423 1200 2424
rect 1204 2423 1205 2427
rect 1335 2427 1341 2428
rect 1335 2426 1336 2427
rect 1325 2424 1336 2426
rect 1199 2422 1205 2423
rect 1335 2423 1336 2424
rect 1340 2423 1341 2427
rect 1822 2424 1823 2428
rect 1827 2424 1828 2428
rect 1822 2423 1828 2424
rect 1886 2427 1892 2428
rect 1886 2423 1887 2427
rect 1891 2423 1892 2427
rect 1335 2422 1341 2423
rect 1886 2422 1892 2423
rect 2014 2427 2020 2428
rect 2014 2423 2015 2427
rect 2019 2423 2020 2427
rect 2014 2422 2020 2423
rect 2174 2427 2180 2428
rect 2174 2423 2175 2427
rect 2179 2423 2180 2427
rect 2174 2422 2180 2423
rect 2334 2427 2340 2428
rect 2334 2423 2335 2427
rect 2339 2423 2340 2427
rect 2334 2422 2340 2423
rect 2494 2427 2500 2428
rect 2494 2423 2495 2427
rect 2499 2423 2500 2427
rect 2494 2422 2500 2423
rect 2646 2427 2652 2428
rect 2646 2423 2647 2427
rect 2651 2423 2652 2427
rect 2646 2422 2652 2423
rect 2798 2427 2804 2428
rect 2798 2423 2799 2427
rect 2803 2423 2804 2427
rect 2798 2422 2804 2423
rect 2950 2427 2956 2428
rect 2950 2423 2951 2427
rect 2955 2423 2956 2427
rect 2950 2422 2956 2423
rect 3110 2427 3116 2428
rect 3110 2423 3111 2427
rect 3115 2423 3116 2427
rect 3110 2422 3116 2423
rect 799 2420 881 2422
rect 799 2419 800 2420
rect 794 2418 800 2419
rect 2167 2419 2173 2420
rect 1862 2417 1868 2418
rect 1862 2413 1863 2417
rect 1867 2413 1868 2417
rect 2167 2415 2168 2419
rect 2172 2418 2173 2419
rect 3018 2419 3024 2420
rect 2172 2416 2193 2418
rect 2172 2415 2173 2416
rect 2167 2414 2173 2415
rect 3018 2415 3019 2419
rect 3023 2418 3024 2419
rect 3023 2416 3129 2418
rect 3574 2417 3580 2418
rect 3023 2415 3024 2416
rect 3018 2414 3024 2415
rect 1862 2412 1868 2413
rect 3574 2413 3575 2417
rect 3579 2413 3580 2417
rect 3574 2412 3580 2413
rect 110 2411 116 2412
rect 110 2407 111 2411
rect 115 2407 116 2411
rect 110 2406 116 2407
rect 174 2411 180 2412
rect 174 2407 175 2411
rect 179 2410 180 2411
rect 1338 2411 1344 2412
rect 179 2408 201 2410
rect 179 2407 180 2408
rect 174 2406 180 2407
rect 1338 2407 1339 2411
rect 1343 2410 1344 2411
rect 1822 2411 1828 2412
rect 1343 2408 1417 2410
rect 1343 2407 1344 2408
rect 1338 2406 1344 2407
rect 1822 2407 1823 2411
rect 1827 2407 1828 2411
rect 1822 2406 1828 2407
rect 1954 2403 1960 2404
rect 1954 2402 1955 2403
rect 182 2401 188 2402
rect 182 2397 183 2401
rect 187 2397 188 2401
rect 182 2396 188 2397
rect 310 2401 316 2402
rect 310 2397 311 2401
rect 315 2397 316 2401
rect 310 2396 316 2397
rect 446 2401 452 2402
rect 446 2397 447 2401
rect 451 2397 452 2401
rect 446 2396 452 2397
rect 582 2401 588 2402
rect 582 2397 583 2401
rect 587 2397 588 2401
rect 582 2396 588 2397
rect 718 2401 724 2402
rect 718 2397 719 2401
rect 723 2397 724 2401
rect 718 2396 724 2397
rect 854 2401 860 2402
rect 854 2397 855 2401
rect 859 2397 860 2401
rect 854 2396 860 2397
rect 990 2401 996 2402
rect 990 2397 991 2401
rect 995 2397 996 2401
rect 990 2396 996 2397
rect 1126 2401 1132 2402
rect 1126 2397 1127 2401
rect 1131 2397 1132 2401
rect 1126 2396 1132 2397
rect 1262 2401 1268 2402
rect 1262 2397 1263 2401
rect 1267 2397 1268 2401
rect 1262 2396 1268 2397
rect 1398 2401 1404 2402
rect 1398 2397 1399 2401
rect 1403 2397 1404 2401
rect 1398 2396 1404 2397
rect 1862 2400 1868 2401
rect 1949 2400 1955 2402
rect 1862 2396 1863 2400
rect 1867 2396 1868 2400
rect 1954 2399 1955 2400
rect 1959 2399 1960 2403
rect 1954 2398 1960 2399
rect 1962 2403 1968 2404
rect 1962 2399 1963 2403
rect 1967 2402 1968 2403
rect 2242 2403 2248 2404
rect 1967 2400 2041 2402
rect 1967 2399 1968 2400
rect 1962 2398 1968 2399
rect 2242 2399 2243 2403
rect 2247 2402 2248 2403
rect 2402 2403 2408 2404
rect 2247 2400 2361 2402
rect 2247 2399 2248 2400
rect 2242 2398 2248 2399
rect 2402 2399 2403 2403
rect 2407 2402 2408 2403
rect 2791 2403 2797 2404
rect 2791 2402 2792 2403
rect 2407 2400 2521 2402
rect 2709 2400 2792 2402
rect 2407 2399 2408 2400
rect 2402 2398 2408 2399
rect 2791 2399 2792 2400
rect 2796 2399 2797 2403
rect 2943 2403 2949 2404
rect 2943 2402 2944 2403
rect 2861 2400 2944 2402
rect 2791 2398 2797 2399
rect 2943 2399 2944 2400
rect 2948 2399 2949 2403
rect 3103 2403 3109 2404
rect 3103 2402 3104 2403
rect 3013 2400 3104 2402
rect 2943 2398 2949 2399
rect 3103 2399 3104 2400
rect 3108 2399 3109 2403
rect 3103 2398 3109 2399
rect 3574 2400 3580 2401
rect 1862 2395 1868 2396
rect 3574 2396 3575 2400
rect 3579 2396 3580 2400
rect 3574 2395 3580 2396
rect 1894 2387 1900 2388
rect 1894 2383 1895 2387
rect 1899 2383 1900 2387
rect 1894 2382 1900 2383
rect 2022 2387 2028 2388
rect 2022 2383 2023 2387
rect 2027 2383 2028 2387
rect 2022 2382 2028 2383
rect 2182 2387 2188 2388
rect 2182 2383 2183 2387
rect 2187 2383 2188 2387
rect 2182 2382 2188 2383
rect 2342 2387 2348 2388
rect 2342 2383 2343 2387
rect 2347 2383 2348 2387
rect 2342 2382 2348 2383
rect 2502 2387 2508 2388
rect 2502 2383 2503 2387
rect 2507 2383 2508 2387
rect 2502 2382 2508 2383
rect 2654 2387 2660 2388
rect 2654 2383 2655 2387
rect 2659 2383 2660 2387
rect 2654 2382 2660 2383
rect 2806 2387 2812 2388
rect 2806 2383 2807 2387
rect 2811 2383 2812 2387
rect 2806 2382 2812 2383
rect 2958 2387 2964 2388
rect 2958 2383 2959 2387
rect 2963 2383 2964 2387
rect 2958 2382 2964 2383
rect 3118 2387 3124 2388
rect 3118 2383 3119 2387
rect 3123 2383 3124 2387
rect 3118 2382 3124 2383
rect 1887 2375 1893 2376
rect 1887 2371 1888 2375
rect 1892 2374 1893 2375
rect 1962 2375 1968 2376
rect 1962 2374 1963 2375
rect 1892 2372 1963 2374
rect 1892 2371 1893 2372
rect 1887 2370 1893 2371
rect 1962 2371 1963 2372
rect 1967 2371 1968 2375
rect 1962 2370 1968 2371
rect 2015 2375 2021 2376
rect 2015 2371 2016 2375
rect 2020 2374 2021 2375
rect 2030 2375 2036 2376
rect 2030 2374 2031 2375
rect 2020 2372 2031 2374
rect 2020 2371 2021 2372
rect 2015 2370 2021 2371
rect 2030 2371 2031 2372
rect 2035 2371 2036 2375
rect 2030 2370 2036 2371
rect 2175 2375 2181 2376
rect 2175 2371 2176 2375
rect 2180 2374 2181 2375
rect 2242 2375 2248 2376
rect 2242 2374 2243 2375
rect 2180 2372 2243 2374
rect 2180 2371 2181 2372
rect 2175 2370 2181 2371
rect 2242 2371 2243 2372
rect 2247 2371 2248 2375
rect 2242 2370 2248 2371
rect 2335 2375 2341 2376
rect 2335 2371 2336 2375
rect 2340 2374 2341 2375
rect 2402 2375 2408 2376
rect 2402 2374 2403 2375
rect 2340 2372 2403 2374
rect 2340 2371 2341 2372
rect 2335 2370 2341 2371
rect 2402 2371 2403 2372
rect 2407 2371 2408 2375
rect 2402 2370 2408 2371
rect 2471 2375 2477 2376
rect 2471 2371 2472 2375
rect 2476 2374 2477 2375
rect 2495 2375 2501 2376
rect 2495 2374 2496 2375
rect 2476 2372 2496 2374
rect 2476 2371 2477 2372
rect 2471 2370 2477 2371
rect 2495 2371 2496 2372
rect 2500 2371 2501 2375
rect 2495 2370 2501 2371
rect 2647 2375 2653 2376
rect 2647 2371 2648 2375
rect 2652 2374 2653 2375
rect 2662 2375 2668 2376
rect 2662 2374 2663 2375
rect 2652 2372 2663 2374
rect 2652 2371 2653 2372
rect 2647 2370 2653 2371
rect 2662 2371 2663 2372
rect 2667 2371 2668 2375
rect 2662 2370 2668 2371
rect 2791 2375 2797 2376
rect 2791 2371 2792 2375
rect 2796 2374 2797 2375
rect 2799 2375 2805 2376
rect 2799 2374 2800 2375
rect 2796 2372 2800 2374
rect 2796 2371 2797 2372
rect 2791 2370 2797 2371
rect 2799 2371 2800 2372
rect 2804 2371 2805 2375
rect 2799 2370 2805 2371
rect 2943 2375 2949 2376
rect 2943 2371 2944 2375
rect 2948 2374 2949 2375
rect 2951 2375 2957 2376
rect 2951 2374 2952 2375
rect 2948 2372 2952 2374
rect 2948 2371 2949 2372
rect 2943 2370 2949 2371
rect 2951 2371 2952 2372
rect 2956 2371 2957 2375
rect 2951 2370 2957 2371
rect 3103 2375 3109 2376
rect 3103 2371 3104 2375
rect 3108 2374 3109 2375
rect 3111 2375 3117 2376
rect 3111 2374 3112 2375
rect 3108 2372 3112 2374
rect 3108 2371 3109 2372
rect 3103 2370 3109 2371
rect 3111 2371 3112 2372
rect 3116 2371 3117 2375
rect 3111 2370 3117 2371
rect 158 2367 164 2368
rect 158 2363 159 2367
rect 163 2363 164 2367
rect 158 2362 164 2363
rect 246 2367 252 2368
rect 246 2363 247 2367
rect 251 2363 252 2367
rect 246 2362 252 2363
rect 334 2367 340 2368
rect 334 2363 335 2367
rect 339 2363 340 2367
rect 334 2362 340 2363
rect 438 2367 444 2368
rect 438 2363 439 2367
rect 443 2363 444 2367
rect 438 2362 444 2363
rect 558 2367 564 2368
rect 558 2363 559 2367
rect 563 2363 564 2367
rect 558 2362 564 2363
rect 686 2367 692 2368
rect 686 2363 687 2367
rect 691 2363 692 2367
rect 686 2362 692 2363
rect 814 2367 820 2368
rect 814 2363 815 2367
rect 819 2363 820 2367
rect 814 2362 820 2363
rect 950 2367 956 2368
rect 950 2363 951 2367
rect 955 2363 956 2367
rect 950 2362 956 2363
rect 1078 2367 1084 2368
rect 1078 2363 1079 2367
rect 1083 2363 1084 2367
rect 1078 2362 1084 2363
rect 1206 2367 1212 2368
rect 1206 2363 1207 2367
rect 1211 2363 1212 2367
rect 1206 2362 1212 2363
rect 1326 2367 1332 2368
rect 1326 2363 1327 2367
rect 1331 2363 1332 2367
rect 1326 2362 1332 2363
rect 1454 2367 1460 2368
rect 1454 2363 1455 2367
rect 1459 2363 1460 2367
rect 1454 2362 1460 2363
rect 1582 2367 1588 2368
rect 1582 2363 1583 2367
rect 1587 2363 1588 2367
rect 2478 2367 2484 2368
rect 2478 2366 2479 2367
rect 1582 2362 1588 2363
rect 2299 2364 2479 2366
rect 766 2359 772 2360
rect 110 2357 116 2358
rect 110 2353 111 2357
rect 115 2353 116 2357
rect 766 2355 767 2359
rect 771 2358 772 2359
rect 886 2359 892 2360
rect 771 2356 833 2358
rect 771 2355 772 2356
rect 766 2354 772 2355
rect 886 2355 887 2359
rect 891 2358 892 2359
rect 1522 2359 1528 2360
rect 891 2356 969 2358
rect 891 2355 892 2356
rect 886 2354 892 2355
rect 1522 2355 1523 2359
rect 1527 2358 1528 2359
rect 1919 2359 1925 2360
rect 1527 2356 1601 2358
rect 1822 2357 1828 2358
rect 1527 2355 1528 2356
rect 1522 2354 1528 2355
rect 110 2352 116 2353
rect 1822 2353 1823 2357
rect 1827 2353 1828 2357
rect 1919 2355 1920 2359
rect 1924 2358 1925 2359
rect 1954 2359 1960 2360
rect 1954 2358 1955 2359
rect 1924 2356 1955 2358
rect 1924 2355 1925 2356
rect 1919 2354 1925 2355
rect 1954 2355 1955 2356
rect 1959 2355 1960 2359
rect 1954 2354 1960 2355
rect 2007 2359 2013 2360
rect 2007 2355 2008 2359
rect 2012 2358 2013 2359
rect 2079 2359 2085 2360
rect 2079 2358 2080 2359
rect 2012 2356 2080 2358
rect 2012 2355 2013 2356
rect 2007 2354 2013 2355
rect 2079 2355 2080 2356
rect 2084 2355 2085 2359
rect 2079 2354 2085 2355
rect 2239 2359 2245 2360
rect 2239 2355 2240 2359
rect 2244 2358 2245 2359
rect 2299 2358 2301 2364
rect 2478 2363 2479 2364
rect 2483 2363 2484 2367
rect 2478 2362 2484 2363
rect 2244 2356 2301 2358
rect 2327 2359 2333 2360
rect 2244 2355 2245 2356
rect 2239 2354 2245 2355
rect 2327 2355 2328 2359
rect 2332 2358 2333 2359
rect 2399 2359 2405 2360
rect 2399 2358 2400 2359
rect 2332 2356 2400 2358
rect 2332 2355 2333 2356
rect 2327 2354 2333 2355
rect 2399 2355 2400 2356
rect 2404 2355 2405 2359
rect 2399 2354 2405 2355
rect 2551 2359 2557 2360
rect 2551 2355 2552 2359
rect 2556 2358 2557 2359
rect 2566 2359 2572 2360
rect 2566 2358 2567 2359
rect 2556 2356 2567 2358
rect 2556 2355 2557 2356
rect 2551 2354 2557 2355
rect 2566 2355 2567 2356
rect 2571 2355 2572 2359
rect 2566 2354 2572 2355
rect 2695 2359 2701 2360
rect 2695 2355 2696 2359
rect 2700 2358 2701 2359
rect 2710 2359 2716 2360
rect 2710 2358 2711 2359
rect 2700 2356 2711 2358
rect 2700 2355 2701 2356
rect 2695 2354 2701 2355
rect 2710 2355 2711 2356
rect 2715 2355 2716 2359
rect 2710 2354 2716 2355
rect 2767 2359 2773 2360
rect 2767 2355 2768 2359
rect 2772 2358 2773 2359
rect 2823 2359 2829 2360
rect 2823 2358 2824 2359
rect 2772 2356 2824 2358
rect 2772 2355 2773 2356
rect 2767 2354 2773 2355
rect 2823 2355 2824 2356
rect 2828 2355 2829 2359
rect 2823 2354 2829 2355
rect 2895 2359 2901 2360
rect 2895 2355 2896 2359
rect 2900 2358 2901 2359
rect 2943 2359 2949 2360
rect 2943 2358 2944 2359
rect 2900 2356 2944 2358
rect 2900 2355 2901 2356
rect 2895 2354 2901 2355
rect 2943 2355 2944 2356
rect 2948 2355 2949 2359
rect 2943 2354 2949 2355
rect 3015 2359 3021 2360
rect 3015 2355 3016 2359
rect 3020 2358 3021 2359
rect 3063 2359 3069 2360
rect 3063 2358 3064 2359
rect 3020 2356 3064 2358
rect 3020 2355 3021 2356
rect 3015 2354 3021 2355
rect 3063 2355 3064 2356
rect 3068 2355 3069 2359
rect 3063 2354 3069 2355
rect 3135 2359 3141 2360
rect 3135 2355 3136 2359
rect 3140 2358 3141 2359
rect 3175 2359 3181 2360
rect 3175 2358 3176 2359
rect 3140 2356 3176 2358
rect 3140 2355 3141 2356
rect 3135 2354 3141 2355
rect 3175 2355 3176 2356
rect 3180 2355 3181 2359
rect 3175 2354 3181 2355
rect 3263 2359 3269 2360
rect 3263 2355 3264 2359
rect 3268 2358 3269 2359
rect 3279 2359 3285 2360
rect 3279 2358 3280 2359
rect 3268 2356 3280 2358
rect 3268 2355 3269 2356
rect 3263 2354 3269 2355
rect 3279 2355 3280 2356
rect 3284 2355 3285 2359
rect 3279 2354 3285 2355
rect 3383 2359 3389 2360
rect 3383 2355 3384 2359
rect 3388 2358 3389 2359
rect 3391 2359 3397 2360
rect 3391 2358 3392 2359
rect 3388 2356 3392 2358
rect 3388 2355 3389 2356
rect 3383 2354 3389 2355
rect 3391 2355 3392 2356
rect 3396 2355 3397 2359
rect 3391 2354 3397 2355
rect 3463 2359 3469 2360
rect 3463 2355 3464 2359
rect 3468 2358 3469 2359
rect 3479 2359 3485 2360
rect 3479 2358 3480 2359
rect 3468 2356 3480 2358
rect 3468 2355 3469 2356
rect 3463 2354 3469 2355
rect 3479 2355 3480 2356
rect 3484 2355 3485 2359
rect 3479 2354 3485 2355
rect 1822 2352 1828 2353
rect 1926 2349 1932 2350
rect 1926 2345 1927 2349
rect 1931 2345 1932 2349
rect 1926 2344 1932 2345
rect 2086 2349 2092 2350
rect 2086 2345 2087 2349
rect 2091 2345 2092 2349
rect 2086 2344 2092 2345
rect 2246 2349 2252 2350
rect 2246 2345 2247 2349
rect 2251 2345 2252 2349
rect 2246 2344 2252 2345
rect 2406 2349 2412 2350
rect 2406 2345 2407 2349
rect 2411 2345 2412 2349
rect 2406 2344 2412 2345
rect 2558 2349 2564 2350
rect 2558 2345 2559 2349
rect 2563 2345 2564 2349
rect 2558 2344 2564 2345
rect 2702 2349 2708 2350
rect 2702 2345 2703 2349
rect 2707 2345 2708 2349
rect 2702 2344 2708 2345
rect 2830 2349 2836 2350
rect 2830 2345 2831 2349
rect 2835 2345 2836 2349
rect 2830 2344 2836 2345
rect 2950 2349 2956 2350
rect 2950 2345 2951 2349
rect 2955 2345 2956 2349
rect 2950 2344 2956 2345
rect 3070 2349 3076 2350
rect 3070 2345 3071 2349
rect 3075 2345 3076 2349
rect 3070 2344 3076 2345
rect 3182 2349 3188 2350
rect 3182 2345 3183 2349
rect 3187 2345 3188 2349
rect 3182 2344 3188 2345
rect 3286 2349 3292 2350
rect 3286 2345 3287 2349
rect 3291 2345 3292 2349
rect 3286 2344 3292 2345
rect 3398 2349 3404 2350
rect 3398 2345 3399 2349
rect 3403 2345 3404 2349
rect 3398 2344 3404 2345
rect 3486 2349 3492 2350
rect 3486 2345 3487 2349
rect 3491 2345 3492 2349
rect 3486 2344 3492 2345
rect 226 2343 232 2344
rect 226 2342 227 2343
rect 110 2340 116 2341
rect 221 2340 227 2342
rect 110 2336 111 2340
rect 115 2336 116 2340
rect 226 2339 227 2340
rect 231 2339 232 2343
rect 314 2343 320 2344
rect 314 2342 315 2343
rect 309 2340 315 2342
rect 226 2338 232 2339
rect 314 2339 315 2340
rect 319 2339 320 2343
rect 402 2343 408 2344
rect 402 2342 403 2343
rect 397 2340 403 2342
rect 314 2338 320 2339
rect 402 2339 403 2340
rect 407 2339 408 2343
rect 511 2343 517 2344
rect 511 2342 512 2343
rect 501 2340 512 2342
rect 402 2338 408 2339
rect 511 2339 512 2340
rect 516 2339 517 2343
rect 654 2343 660 2344
rect 654 2342 655 2343
rect 621 2340 655 2342
rect 511 2338 517 2339
rect 654 2339 655 2340
rect 659 2339 660 2343
rect 762 2343 768 2344
rect 762 2342 763 2343
rect 749 2340 763 2342
rect 654 2338 660 2339
rect 762 2339 763 2340
rect 767 2339 768 2343
rect 1154 2343 1160 2344
rect 1154 2342 1155 2343
rect 1141 2340 1155 2342
rect 762 2338 768 2339
rect 1154 2339 1155 2340
rect 1159 2339 1160 2343
rect 1279 2343 1285 2344
rect 1279 2342 1280 2343
rect 1269 2340 1280 2342
rect 1154 2338 1160 2339
rect 1279 2339 1280 2340
rect 1284 2339 1285 2343
rect 1402 2343 1408 2344
rect 1402 2342 1403 2343
rect 1389 2340 1403 2342
rect 1279 2338 1285 2339
rect 1402 2339 1403 2340
rect 1407 2339 1408 2343
rect 1530 2343 1536 2344
rect 1530 2342 1531 2343
rect 1517 2340 1531 2342
rect 1402 2338 1408 2339
rect 1530 2339 1531 2340
rect 1535 2339 1536 2343
rect 1530 2338 1536 2339
rect 1822 2340 1828 2341
rect 110 2335 116 2336
rect 1822 2336 1823 2340
rect 1827 2336 1828 2340
rect 1822 2335 1828 2336
rect 1862 2336 1868 2337
rect 3574 2336 3580 2337
rect 1862 2332 1863 2336
rect 1867 2332 1868 2336
rect 2007 2335 2013 2336
rect 2007 2334 2008 2335
rect 1981 2332 2008 2334
rect 1862 2331 1868 2332
rect 2007 2331 2008 2332
rect 2012 2331 2013 2335
rect 2327 2335 2333 2336
rect 2327 2334 2328 2335
rect 2301 2332 2328 2334
rect 2007 2330 2013 2331
rect 2327 2331 2328 2332
rect 2332 2331 2333 2335
rect 2471 2335 2477 2336
rect 2471 2334 2472 2335
rect 2461 2332 2472 2334
rect 2327 2330 2333 2331
rect 2471 2331 2472 2332
rect 2476 2331 2477 2335
rect 2767 2335 2773 2336
rect 2767 2334 2768 2335
rect 2757 2332 2768 2334
rect 2471 2330 2477 2331
rect 2767 2331 2768 2332
rect 2772 2331 2773 2335
rect 2895 2335 2901 2336
rect 2895 2334 2896 2335
rect 2885 2332 2896 2334
rect 2767 2330 2773 2331
rect 2895 2331 2896 2332
rect 2900 2331 2901 2335
rect 3015 2335 3021 2336
rect 3015 2334 3016 2335
rect 3005 2332 3016 2334
rect 2895 2330 2901 2331
rect 3015 2331 3016 2332
rect 3020 2331 3021 2335
rect 3135 2335 3141 2336
rect 3135 2334 3136 2335
rect 3125 2332 3136 2334
rect 3015 2330 3021 2331
rect 3135 2331 3136 2332
rect 3140 2331 3141 2335
rect 3383 2335 3389 2336
rect 3383 2334 3384 2335
rect 3341 2332 3384 2334
rect 3135 2330 3141 2331
rect 3383 2331 3384 2332
rect 3388 2331 3389 2335
rect 3463 2335 3469 2336
rect 3463 2334 3464 2335
rect 3453 2332 3464 2334
rect 3383 2330 3389 2331
rect 3463 2331 3464 2332
rect 3468 2331 3469 2335
rect 3574 2332 3575 2336
rect 3579 2332 3580 2336
rect 3574 2331 3580 2332
rect 3463 2330 3469 2331
rect 166 2327 172 2328
rect 166 2323 167 2327
rect 171 2323 172 2327
rect 166 2322 172 2323
rect 254 2327 260 2328
rect 254 2323 255 2327
rect 259 2323 260 2327
rect 254 2322 260 2323
rect 342 2327 348 2328
rect 342 2323 343 2327
rect 347 2323 348 2327
rect 342 2322 348 2323
rect 446 2327 452 2328
rect 446 2323 447 2327
rect 451 2323 452 2327
rect 446 2322 452 2323
rect 566 2327 572 2328
rect 566 2323 567 2327
rect 571 2323 572 2327
rect 566 2322 572 2323
rect 694 2327 700 2328
rect 694 2323 695 2327
rect 699 2323 700 2327
rect 694 2322 700 2323
rect 822 2327 828 2328
rect 822 2323 823 2327
rect 827 2323 828 2327
rect 822 2322 828 2323
rect 958 2327 964 2328
rect 958 2323 959 2327
rect 963 2323 964 2327
rect 958 2322 964 2323
rect 1086 2327 1092 2328
rect 1086 2323 1087 2327
rect 1091 2323 1092 2327
rect 1086 2322 1092 2323
rect 1214 2327 1220 2328
rect 1214 2323 1215 2327
rect 1219 2323 1220 2327
rect 1214 2322 1220 2323
rect 1334 2327 1340 2328
rect 1334 2323 1335 2327
rect 1339 2323 1340 2327
rect 1334 2322 1340 2323
rect 1462 2327 1468 2328
rect 1462 2323 1463 2327
rect 1467 2323 1468 2327
rect 1462 2322 1468 2323
rect 1590 2327 1596 2328
rect 1590 2323 1591 2327
rect 1595 2323 1596 2327
rect 1590 2322 1596 2323
rect 1862 2319 1868 2320
rect 159 2315 165 2316
rect 159 2311 160 2315
rect 164 2314 165 2315
rect 174 2315 180 2316
rect 174 2314 175 2315
rect 164 2312 175 2314
rect 164 2311 165 2312
rect 159 2310 165 2311
rect 174 2311 175 2312
rect 179 2311 180 2315
rect 174 2310 180 2311
rect 226 2315 232 2316
rect 226 2311 227 2315
rect 231 2314 232 2315
rect 247 2315 253 2316
rect 247 2314 248 2315
rect 231 2312 248 2314
rect 231 2311 232 2312
rect 226 2310 232 2311
rect 247 2311 248 2312
rect 252 2311 253 2315
rect 247 2310 253 2311
rect 314 2315 320 2316
rect 314 2311 315 2315
rect 319 2314 320 2315
rect 335 2315 341 2316
rect 335 2314 336 2315
rect 319 2312 336 2314
rect 319 2311 320 2312
rect 314 2310 320 2311
rect 335 2311 336 2312
rect 340 2311 341 2315
rect 335 2310 341 2311
rect 402 2315 408 2316
rect 402 2311 403 2315
rect 407 2314 408 2315
rect 439 2315 445 2316
rect 439 2314 440 2315
rect 407 2312 440 2314
rect 407 2311 408 2312
rect 402 2310 408 2311
rect 439 2311 440 2312
rect 444 2311 445 2315
rect 439 2310 445 2311
rect 511 2315 517 2316
rect 511 2311 512 2315
rect 516 2314 517 2315
rect 559 2315 565 2316
rect 559 2314 560 2315
rect 516 2312 560 2314
rect 516 2311 517 2312
rect 511 2310 517 2311
rect 559 2311 560 2312
rect 564 2311 565 2315
rect 559 2310 565 2311
rect 654 2315 660 2316
rect 654 2311 655 2315
rect 659 2314 660 2315
rect 687 2315 693 2316
rect 687 2314 688 2315
rect 659 2312 688 2314
rect 659 2311 660 2312
rect 654 2310 660 2311
rect 687 2311 688 2312
rect 692 2311 693 2315
rect 687 2310 693 2311
rect 762 2315 768 2316
rect 762 2311 763 2315
rect 767 2314 768 2315
rect 815 2315 821 2316
rect 815 2314 816 2315
rect 767 2312 816 2314
rect 767 2311 768 2312
rect 762 2310 768 2311
rect 815 2311 816 2312
rect 820 2311 821 2315
rect 815 2310 821 2311
rect 927 2315 933 2316
rect 927 2311 928 2315
rect 932 2314 933 2315
rect 951 2315 957 2316
rect 951 2314 952 2315
rect 932 2312 952 2314
rect 932 2311 933 2312
rect 927 2310 933 2311
rect 951 2311 952 2312
rect 956 2311 957 2315
rect 951 2310 957 2311
rect 1079 2315 1085 2316
rect 1079 2311 1080 2315
rect 1084 2314 1085 2315
rect 1134 2315 1140 2316
rect 1134 2314 1135 2315
rect 1084 2312 1135 2314
rect 1084 2311 1085 2312
rect 1079 2310 1085 2311
rect 1134 2311 1135 2312
rect 1139 2311 1140 2315
rect 1134 2310 1140 2311
rect 1154 2315 1160 2316
rect 1154 2311 1155 2315
rect 1159 2314 1160 2315
rect 1207 2315 1213 2316
rect 1207 2314 1208 2315
rect 1159 2312 1208 2314
rect 1159 2311 1160 2312
rect 1154 2310 1160 2311
rect 1207 2311 1208 2312
rect 1212 2311 1213 2315
rect 1207 2310 1213 2311
rect 1279 2315 1285 2316
rect 1279 2311 1280 2315
rect 1284 2314 1285 2315
rect 1327 2315 1333 2316
rect 1327 2314 1328 2315
rect 1284 2312 1328 2314
rect 1284 2311 1285 2312
rect 1279 2310 1285 2311
rect 1327 2311 1328 2312
rect 1332 2311 1333 2315
rect 1327 2310 1333 2311
rect 1402 2315 1408 2316
rect 1402 2311 1403 2315
rect 1407 2314 1408 2315
rect 1455 2315 1461 2316
rect 1455 2314 1456 2315
rect 1407 2312 1456 2314
rect 1407 2311 1408 2312
rect 1402 2310 1408 2311
rect 1455 2311 1456 2312
rect 1460 2311 1461 2315
rect 1455 2310 1461 2311
rect 1530 2315 1536 2316
rect 1530 2311 1531 2315
rect 1535 2314 1536 2315
rect 1583 2315 1589 2316
rect 1583 2314 1584 2315
rect 1535 2312 1584 2314
rect 1535 2311 1536 2312
rect 1530 2310 1536 2311
rect 1583 2311 1584 2312
rect 1588 2311 1589 2315
rect 1862 2315 1863 2319
rect 1867 2315 1868 2319
rect 1862 2314 1868 2315
rect 2478 2319 2484 2320
rect 2478 2315 2479 2319
rect 2483 2318 2484 2319
rect 3182 2319 3188 2320
rect 2483 2316 2569 2318
rect 2483 2315 2484 2316
rect 2478 2314 2484 2315
rect 3182 2315 3183 2319
rect 3187 2318 3188 2319
rect 3471 2319 3477 2320
rect 3187 2316 3193 2318
rect 3187 2315 3188 2316
rect 3182 2314 3188 2315
rect 3471 2315 3472 2319
rect 3476 2318 3477 2319
rect 3574 2319 3580 2320
rect 3476 2316 3497 2318
rect 3476 2315 3477 2316
rect 3471 2314 3477 2315
rect 3574 2315 3575 2319
rect 3579 2315 3580 2319
rect 3574 2314 3580 2315
rect 1583 2310 1589 2311
rect 1918 2309 1924 2310
rect 1918 2305 1919 2309
rect 1923 2305 1924 2309
rect 1918 2304 1924 2305
rect 2078 2309 2084 2310
rect 2078 2305 2079 2309
rect 2083 2305 2084 2309
rect 2078 2304 2084 2305
rect 2238 2309 2244 2310
rect 2238 2305 2239 2309
rect 2243 2305 2244 2309
rect 2238 2304 2244 2305
rect 2398 2309 2404 2310
rect 2398 2305 2399 2309
rect 2403 2305 2404 2309
rect 2398 2304 2404 2305
rect 2550 2309 2556 2310
rect 2550 2305 2551 2309
rect 2555 2305 2556 2309
rect 2550 2304 2556 2305
rect 2694 2309 2700 2310
rect 2694 2305 2695 2309
rect 2699 2305 2700 2309
rect 2694 2304 2700 2305
rect 2822 2309 2828 2310
rect 2822 2305 2823 2309
rect 2827 2305 2828 2309
rect 2822 2304 2828 2305
rect 2942 2309 2948 2310
rect 2942 2305 2943 2309
rect 2947 2305 2948 2309
rect 2942 2304 2948 2305
rect 3062 2309 3068 2310
rect 3062 2305 3063 2309
rect 3067 2305 3068 2309
rect 3062 2304 3068 2305
rect 3174 2309 3180 2310
rect 3174 2305 3175 2309
rect 3179 2305 3180 2309
rect 3174 2304 3180 2305
rect 3278 2309 3284 2310
rect 3278 2305 3279 2309
rect 3283 2305 3284 2309
rect 3278 2304 3284 2305
rect 3390 2309 3396 2310
rect 3390 2305 3391 2309
rect 3395 2305 3396 2309
rect 3390 2304 3396 2305
rect 3478 2309 3484 2310
rect 3478 2305 3479 2309
rect 3483 2305 3484 2309
rect 3478 2304 3484 2305
rect 2127 2303 2133 2304
rect 2127 2299 2128 2303
rect 2132 2302 2133 2303
rect 2135 2303 2141 2304
rect 2135 2302 2136 2303
rect 2132 2300 2136 2302
rect 2132 2299 2133 2300
rect 2127 2298 2133 2299
rect 2135 2299 2136 2300
rect 2140 2299 2141 2303
rect 2135 2298 2141 2299
rect 687 2295 693 2296
rect 687 2291 688 2295
rect 692 2294 693 2295
rect 702 2295 708 2296
rect 702 2294 703 2295
rect 692 2292 703 2294
rect 692 2291 693 2292
rect 687 2290 693 2291
rect 702 2291 703 2292
rect 707 2291 708 2295
rect 702 2290 708 2291
rect 775 2295 781 2296
rect 775 2291 776 2295
rect 780 2294 781 2295
rect 855 2295 861 2296
rect 855 2294 856 2295
rect 780 2292 856 2294
rect 780 2291 781 2292
rect 775 2290 781 2291
rect 855 2291 856 2292
rect 860 2291 861 2295
rect 855 2290 861 2291
rect 1015 2295 1021 2296
rect 1015 2291 1016 2295
rect 1020 2294 1021 2295
rect 1030 2295 1036 2296
rect 1030 2294 1031 2295
rect 1020 2292 1031 2294
rect 1020 2291 1021 2292
rect 1015 2290 1021 2291
rect 1030 2291 1031 2292
rect 1035 2291 1036 2295
rect 1030 2290 1036 2291
rect 1167 2295 1173 2296
rect 1167 2291 1168 2295
rect 1172 2294 1173 2295
rect 1182 2295 1188 2296
rect 1182 2294 1183 2295
rect 1172 2292 1183 2294
rect 1172 2291 1173 2292
rect 1167 2290 1173 2291
rect 1182 2291 1183 2292
rect 1187 2291 1188 2295
rect 1182 2290 1188 2291
rect 1247 2295 1253 2296
rect 1247 2291 1248 2295
rect 1252 2294 1253 2295
rect 1311 2295 1317 2296
rect 1311 2294 1312 2295
rect 1252 2292 1312 2294
rect 1252 2291 1253 2292
rect 1247 2290 1253 2291
rect 1311 2291 1312 2292
rect 1316 2291 1317 2295
rect 1311 2290 1317 2291
rect 1391 2295 1397 2296
rect 1391 2291 1392 2295
rect 1396 2294 1397 2295
rect 1455 2295 1461 2296
rect 1455 2294 1456 2295
rect 1396 2292 1456 2294
rect 1396 2291 1397 2292
rect 1391 2290 1397 2291
rect 1455 2291 1456 2292
rect 1460 2291 1461 2295
rect 1455 2290 1461 2291
rect 1527 2295 1533 2296
rect 1527 2291 1528 2295
rect 1532 2294 1533 2295
rect 1591 2295 1597 2296
rect 1591 2294 1592 2295
rect 1532 2292 1592 2294
rect 1532 2291 1533 2292
rect 1527 2290 1533 2291
rect 1591 2291 1592 2292
rect 1596 2291 1597 2295
rect 1591 2290 1597 2291
rect 1663 2295 1669 2296
rect 1663 2291 1664 2295
rect 1668 2294 1669 2295
rect 1727 2295 1733 2296
rect 1727 2294 1728 2295
rect 1668 2292 1728 2294
rect 1668 2291 1669 2292
rect 1663 2290 1669 2291
rect 1727 2291 1728 2292
rect 1732 2291 1733 2295
rect 1727 2290 1733 2291
rect 694 2285 700 2286
rect 694 2281 695 2285
rect 699 2281 700 2285
rect 694 2280 700 2281
rect 862 2285 868 2286
rect 862 2281 863 2285
rect 867 2281 868 2285
rect 862 2280 868 2281
rect 1022 2285 1028 2286
rect 1022 2281 1023 2285
rect 1027 2281 1028 2285
rect 1022 2280 1028 2281
rect 1174 2285 1180 2286
rect 1174 2281 1175 2285
rect 1179 2281 1180 2285
rect 1174 2280 1180 2281
rect 1318 2285 1324 2286
rect 1318 2281 1319 2285
rect 1323 2281 1324 2285
rect 1318 2280 1324 2281
rect 1462 2285 1468 2286
rect 1462 2281 1463 2285
rect 1467 2281 1468 2285
rect 1462 2280 1468 2281
rect 1598 2285 1604 2286
rect 1598 2281 1599 2285
rect 1603 2281 1604 2285
rect 1598 2280 1604 2281
rect 1734 2285 1740 2286
rect 1734 2281 1735 2285
rect 1739 2281 1740 2285
rect 1734 2280 1740 2281
rect 1974 2283 1980 2284
rect 1974 2279 1975 2283
rect 1979 2279 1980 2283
rect 1974 2278 1980 2279
rect 2142 2283 2148 2284
rect 2142 2279 2143 2283
rect 2147 2279 2148 2283
rect 2142 2278 2148 2279
rect 2310 2283 2316 2284
rect 2310 2279 2311 2283
rect 2315 2279 2316 2283
rect 2310 2278 2316 2279
rect 2478 2283 2484 2284
rect 2478 2279 2479 2283
rect 2483 2279 2484 2283
rect 2478 2278 2484 2279
rect 2638 2283 2644 2284
rect 2638 2279 2639 2283
rect 2643 2279 2644 2283
rect 2638 2278 2644 2279
rect 2782 2283 2788 2284
rect 2782 2279 2783 2283
rect 2787 2279 2788 2283
rect 2782 2278 2788 2279
rect 2918 2283 2924 2284
rect 2918 2279 2919 2283
rect 2923 2279 2924 2283
rect 2918 2278 2924 2279
rect 3038 2283 3044 2284
rect 3038 2279 3039 2283
rect 3043 2279 3044 2283
rect 3038 2278 3044 2279
rect 3158 2283 3164 2284
rect 3158 2279 3159 2283
rect 3163 2279 3164 2283
rect 3158 2278 3164 2279
rect 3270 2283 3276 2284
rect 3270 2279 3271 2283
rect 3275 2279 3276 2283
rect 3270 2278 3276 2279
rect 3382 2283 3388 2284
rect 3382 2279 3383 2283
rect 3387 2279 3388 2283
rect 3382 2278 3388 2279
rect 3478 2283 3484 2284
rect 3478 2279 3479 2283
rect 3483 2279 3484 2283
rect 3478 2278 3484 2279
rect 2566 2275 2572 2276
rect 1862 2273 1868 2274
rect 110 2272 116 2273
rect 1822 2272 1828 2273
rect 110 2268 111 2272
rect 115 2268 116 2272
rect 775 2271 781 2272
rect 775 2270 776 2271
rect 749 2268 776 2270
rect 110 2267 116 2268
rect 775 2267 776 2268
rect 780 2267 781 2271
rect 927 2271 933 2272
rect 927 2270 928 2271
rect 917 2268 928 2270
rect 775 2266 781 2267
rect 927 2267 928 2268
rect 932 2267 933 2271
rect 1247 2271 1253 2272
rect 1247 2270 1248 2271
rect 1229 2268 1248 2270
rect 927 2266 933 2267
rect 938 2267 944 2268
rect 938 2263 939 2267
rect 943 2266 944 2267
rect 1247 2267 1248 2268
rect 1252 2267 1253 2271
rect 1391 2271 1397 2272
rect 1391 2270 1392 2271
rect 1373 2268 1392 2270
rect 1247 2266 1253 2267
rect 1391 2267 1392 2268
rect 1396 2267 1397 2271
rect 1527 2271 1533 2272
rect 1527 2270 1528 2271
rect 1517 2268 1528 2270
rect 1391 2266 1397 2267
rect 1527 2267 1528 2268
rect 1532 2267 1533 2271
rect 1663 2271 1669 2272
rect 1663 2270 1664 2271
rect 1653 2268 1664 2270
rect 1527 2266 1533 2267
rect 1663 2267 1664 2268
rect 1668 2267 1669 2271
rect 1822 2268 1823 2272
rect 1827 2268 1828 2272
rect 1862 2269 1863 2273
rect 1867 2269 1868 2273
rect 2566 2271 2567 2275
rect 2571 2274 2572 2275
rect 3110 2275 3116 2276
rect 2571 2272 2657 2274
rect 2571 2271 2572 2272
rect 2566 2270 2572 2271
rect 3110 2271 3111 2275
rect 3115 2274 3116 2275
rect 3263 2275 3269 2276
rect 3115 2272 3177 2274
rect 3115 2271 3116 2272
rect 3110 2270 3116 2271
rect 3263 2271 3264 2275
rect 3268 2274 3269 2275
rect 3268 2272 3289 2274
rect 3574 2273 3580 2274
rect 3268 2271 3269 2272
rect 3263 2270 3269 2271
rect 1862 2268 1868 2269
rect 3574 2269 3575 2273
rect 3579 2269 3580 2273
rect 3574 2268 3580 2269
rect 1822 2267 1828 2268
rect 1663 2266 1669 2267
rect 943 2264 1041 2266
rect 943 2263 944 2264
rect 938 2262 944 2263
rect 2042 2259 2048 2260
rect 2042 2258 2043 2259
rect 1862 2256 1868 2257
rect 2037 2256 2043 2258
rect 110 2255 116 2256
rect 110 2251 111 2255
rect 115 2251 116 2255
rect 110 2250 116 2251
rect 1666 2255 1672 2256
rect 1666 2251 1667 2255
rect 1671 2254 1672 2255
rect 1822 2255 1828 2256
rect 1671 2252 1745 2254
rect 1671 2251 1672 2252
rect 1666 2250 1672 2251
rect 1822 2251 1823 2255
rect 1827 2251 1828 2255
rect 1862 2252 1863 2256
rect 1867 2252 1868 2256
rect 2042 2255 2043 2256
rect 2047 2255 2048 2259
rect 2042 2254 2048 2255
rect 2050 2259 2056 2260
rect 2050 2255 2051 2259
rect 2055 2258 2056 2259
rect 2471 2259 2477 2260
rect 2471 2258 2472 2259
rect 2055 2256 2169 2258
rect 2373 2256 2472 2258
rect 2055 2255 2056 2256
rect 2050 2254 2056 2255
rect 2471 2255 2472 2256
rect 2476 2255 2477 2259
rect 2631 2259 2637 2260
rect 2631 2258 2632 2259
rect 2541 2256 2632 2258
rect 2471 2254 2477 2255
rect 2631 2255 2632 2256
rect 2636 2255 2637 2259
rect 2911 2259 2917 2260
rect 2911 2258 2912 2259
rect 2845 2256 2912 2258
rect 2631 2254 2637 2255
rect 2911 2255 2912 2256
rect 2916 2255 2917 2259
rect 3031 2259 3037 2260
rect 3031 2258 3032 2259
rect 2981 2256 3032 2258
rect 2911 2254 2917 2255
rect 3031 2255 3032 2256
rect 3036 2255 3037 2259
rect 3150 2259 3156 2260
rect 3150 2258 3151 2259
rect 3101 2256 3151 2258
rect 3031 2254 3037 2255
rect 3150 2255 3151 2256
rect 3155 2255 3156 2259
rect 3150 2254 3156 2255
rect 3338 2259 3344 2260
rect 3338 2255 3339 2259
rect 3343 2258 3344 2259
rect 3470 2259 3476 2260
rect 3343 2256 3409 2258
rect 3343 2255 3344 2256
rect 3338 2254 3344 2255
rect 3470 2255 3471 2259
rect 3475 2258 3476 2259
rect 3475 2256 3505 2258
rect 3574 2256 3580 2257
rect 3475 2255 3476 2256
rect 3470 2254 3476 2255
rect 1862 2251 1868 2252
rect 3574 2252 3575 2256
rect 3579 2252 3580 2256
rect 3574 2251 3580 2252
rect 1822 2250 1828 2251
rect 686 2245 692 2246
rect 686 2241 687 2245
rect 691 2241 692 2245
rect 686 2240 692 2241
rect 854 2245 860 2246
rect 854 2241 855 2245
rect 859 2241 860 2245
rect 854 2240 860 2241
rect 1014 2245 1020 2246
rect 1014 2241 1015 2245
rect 1019 2241 1020 2245
rect 1014 2240 1020 2241
rect 1166 2245 1172 2246
rect 1166 2241 1167 2245
rect 1171 2241 1172 2245
rect 1166 2240 1172 2241
rect 1310 2245 1316 2246
rect 1310 2241 1311 2245
rect 1315 2241 1316 2245
rect 1310 2240 1316 2241
rect 1454 2245 1460 2246
rect 1454 2241 1455 2245
rect 1459 2241 1460 2245
rect 1454 2240 1460 2241
rect 1590 2245 1596 2246
rect 1590 2241 1591 2245
rect 1595 2241 1596 2245
rect 1590 2240 1596 2241
rect 1726 2245 1732 2246
rect 1726 2241 1727 2245
rect 1731 2241 1732 2245
rect 1726 2240 1732 2241
rect 1982 2243 1988 2244
rect 1982 2239 1983 2243
rect 1987 2239 1988 2243
rect 1982 2238 1988 2239
rect 2150 2243 2156 2244
rect 2150 2239 2151 2243
rect 2155 2239 2156 2243
rect 2150 2238 2156 2239
rect 2318 2243 2324 2244
rect 2318 2239 2319 2243
rect 2323 2239 2324 2243
rect 2318 2238 2324 2239
rect 2486 2243 2492 2244
rect 2486 2239 2487 2243
rect 2491 2239 2492 2243
rect 2486 2238 2492 2239
rect 2646 2243 2652 2244
rect 2646 2239 2647 2243
rect 2651 2239 2652 2243
rect 2646 2238 2652 2239
rect 2790 2243 2796 2244
rect 2790 2239 2791 2243
rect 2795 2239 2796 2243
rect 2790 2238 2796 2239
rect 2926 2243 2932 2244
rect 2926 2239 2927 2243
rect 2931 2239 2932 2243
rect 2926 2238 2932 2239
rect 3046 2243 3052 2244
rect 3046 2239 3047 2243
rect 3051 2239 3052 2243
rect 3046 2238 3052 2239
rect 3166 2243 3172 2244
rect 3166 2239 3167 2243
rect 3171 2239 3172 2243
rect 3166 2238 3172 2239
rect 3278 2243 3284 2244
rect 3278 2239 3279 2243
rect 3283 2239 3284 2243
rect 3278 2238 3284 2239
rect 3390 2243 3396 2244
rect 3390 2239 3391 2243
rect 3395 2239 3396 2243
rect 3390 2238 3396 2239
rect 3486 2243 3492 2244
rect 3486 2239 3487 2243
rect 3491 2239 3492 2243
rect 3486 2238 3492 2239
rect 1975 2231 1981 2232
rect 1975 2227 1976 2231
rect 1980 2230 1981 2231
rect 2050 2231 2056 2232
rect 2050 2230 2051 2231
rect 1980 2228 2051 2230
rect 1980 2227 1981 2228
rect 1975 2226 1981 2227
rect 2050 2227 2051 2228
rect 2055 2227 2056 2231
rect 2050 2226 2056 2227
rect 2135 2231 2141 2232
rect 2135 2227 2136 2231
rect 2140 2230 2141 2231
rect 2143 2231 2149 2232
rect 2143 2230 2144 2231
rect 2140 2228 2144 2230
rect 2140 2227 2141 2228
rect 2135 2226 2141 2227
rect 2143 2227 2144 2228
rect 2148 2227 2149 2231
rect 2143 2226 2149 2227
rect 2311 2231 2317 2232
rect 2311 2227 2312 2231
rect 2316 2230 2317 2231
rect 2402 2231 2408 2232
rect 2402 2230 2403 2231
rect 2316 2228 2403 2230
rect 2316 2227 2317 2228
rect 2311 2226 2317 2227
rect 2402 2227 2403 2228
rect 2407 2227 2408 2231
rect 2402 2226 2408 2227
rect 2471 2231 2477 2232
rect 2471 2227 2472 2231
rect 2476 2230 2477 2231
rect 2479 2231 2485 2232
rect 2479 2230 2480 2231
rect 2476 2228 2480 2230
rect 2476 2227 2477 2228
rect 2471 2226 2477 2227
rect 2479 2227 2480 2228
rect 2484 2227 2485 2231
rect 2479 2226 2485 2227
rect 2631 2231 2637 2232
rect 2631 2227 2632 2231
rect 2636 2230 2637 2231
rect 2639 2231 2645 2232
rect 2639 2230 2640 2231
rect 2636 2228 2640 2230
rect 2636 2227 2637 2228
rect 2631 2226 2637 2227
rect 2639 2227 2640 2228
rect 2644 2227 2645 2231
rect 2639 2226 2645 2227
rect 2783 2231 2789 2232
rect 2783 2227 2784 2231
rect 2788 2230 2789 2231
rect 2798 2231 2804 2232
rect 2798 2230 2799 2231
rect 2788 2228 2799 2230
rect 2788 2227 2789 2228
rect 2783 2226 2789 2227
rect 2798 2227 2799 2228
rect 2803 2227 2804 2231
rect 2798 2226 2804 2227
rect 2911 2231 2917 2232
rect 2911 2227 2912 2231
rect 2916 2230 2917 2231
rect 2919 2231 2925 2232
rect 2919 2230 2920 2231
rect 2916 2228 2920 2230
rect 2916 2227 2917 2228
rect 2911 2226 2917 2227
rect 2919 2227 2920 2228
rect 2924 2227 2925 2231
rect 2919 2226 2925 2227
rect 3031 2231 3037 2232
rect 3031 2227 3032 2231
rect 3036 2230 3037 2231
rect 3039 2231 3045 2232
rect 3039 2230 3040 2231
rect 3036 2228 3040 2230
rect 3036 2227 3037 2228
rect 3031 2226 3037 2227
rect 3039 2227 3040 2228
rect 3044 2227 3045 2231
rect 3039 2226 3045 2227
rect 3150 2231 3156 2232
rect 3150 2227 3151 2231
rect 3155 2230 3156 2231
rect 3159 2231 3165 2232
rect 3159 2230 3160 2231
rect 3155 2228 3160 2230
rect 3155 2227 3156 2228
rect 3150 2226 3156 2227
rect 3159 2227 3160 2228
rect 3164 2227 3165 2231
rect 3159 2226 3165 2227
rect 3271 2231 3277 2232
rect 3271 2227 3272 2231
rect 3276 2230 3277 2231
rect 3338 2231 3344 2232
rect 3338 2230 3339 2231
rect 3276 2228 3339 2230
rect 3276 2227 3277 2228
rect 3271 2226 3277 2227
rect 3338 2227 3339 2228
rect 3343 2227 3344 2231
rect 3338 2226 3344 2227
rect 3367 2231 3373 2232
rect 3367 2227 3368 2231
rect 3372 2230 3373 2231
rect 3383 2231 3389 2232
rect 3383 2230 3384 2231
rect 3372 2228 3384 2230
rect 3372 2227 3373 2228
rect 3367 2226 3373 2227
rect 3383 2227 3384 2228
rect 3388 2227 3389 2231
rect 3383 2226 3389 2227
rect 3471 2231 3477 2232
rect 3471 2227 3472 2231
rect 3476 2230 3477 2231
rect 3479 2231 3485 2232
rect 3479 2230 3480 2231
rect 3476 2228 3480 2230
rect 3476 2227 3477 2228
rect 3471 2226 3477 2227
rect 3479 2227 3480 2228
rect 3484 2227 3485 2231
rect 3479 2226 3485 2227
rect 1999 2219 2005 2220
rect 534 2215 540 2216
rect 534 2211 535 2215
rect 539 2211 540 2215
rect 534 2210 540 2211
rect 718 2215 724 2216
rect 718 2211 719 2215
rect 723 2211 724 2215
rect 718 2210 724 2211
rect 894 2215 900 2216
rect 894 2211 895 2215
rect 899 2211 900 2215
rect 894 2210 900 2211
rect 1070 2215 1076 2216
rect 1070 2211 1071 2215
rect 1075 2211 1076 2215
rect 1070 2210 1076 2211
rect 1238 2215 1244 2216
rect 1238 2211 1239 2215
rect 1243 2211 1244 2215
rect 1238 2210 1244 2211
rect 1406 2215 1412 2216
rect 1406 2211 1407 2215
rect 1411 2211 1412 2215
rect 1406 2210 1412 2211
rect 1574 2215 1580 2216
rect 1574 2211 1575 2215
rect 1579 2211 1580 2215
rect 1574 2210 1580 2211
rect 1726 2215 1732 2216
rect 1726 2211 1727 2215
rect 1731 2211 1732 2215
rect 1999 2215 2000 2219
rect 2004 2218 2005 2219
rect 2042 2219 2048 2220
rect 2042 2218 2043 2219
rect 2004 2216 2043 2218
rect 2004 2215 2005 2216
rect 1999 2214 2005 2215
rect 2042 2215 2043 2216
rect 2047 2215 2048 2219
rect 2042 2214 2048 2215
rect 2087 2219 2093 2220
rect 2087 2215 2088 2219
rect 2092 2218 2093 2219
rect 2159 2219 2165 2220
rect 2159 2218 2160 2219
rect 2092 2216 2160 2218
rect 2092 2215 2093 2216
rect 2087 2214 2093 2215
rect 2159 2215 2160 2216
rect 2164 2215 2165 2219
rect 2159 2214 2165 2215
rect 2239 2219 2245 2220
rect 2239 2215 2240 2219
rect 2244 2218 2245 2219
rect 2327 2219 2333 2220
rect 2327 2218 2328 2219
rect 2244 2216 2328 2218
rect 2244 2215 2245 2216
rect 2239 2214 2245 2215
rect 2327 2215 2328 2216
rect 2332 2215 2333 2219
rect 2327 2214 2333 2215
rect 2511 2219 2517 2220
rect 2511 2215 2512 2219
rect 2516 2218 2517 2219
rect 2586 2219 2592 2220
rect 2586 2218 2587 2219
rect 2516 2216 2587 2218
rect 2516 2215 2517 2216
rect 2511 2214 2517 2215
rect 2586 2215 2587 2216
rect 2591 2215 2592 2219
rect 2586 2214 2592 2215
rect 2703 2219 2709 2220
rect 2703 2215 2704 2219
rect 2708 2218 2709 2219
rect 2807 2219 2813 2220
rect 2807 2218 2808 2219
rect 2708 2216 2808 2218
rect 2708 2215 2709 2216
rect 2703 2214 2709 2215
rect 2807 2215 2808 2216
rect 2812 2215 2813 2219
rect 2807 2214 2813 2215
rect 2838 2219 2844 2220
rect 2838 2215 2839 2219
rect 2843 2218 2844 2219
rect 2895 2219 2901 2220
rect 2895 2218 2896 2219
rect 2843 2216 2896 2218
rect 2843 2215 2844 2216
rect 2838 2214 2844 2215
rect 2895 2215 2896 2216
rect 2900 2215 2901 2219
rect 2895 2214 2901 2215
rect 3095 2219 3101 2220
rect 3095 2215 3096 2219
rect 3100 2218 3101 2219
rect 3110 2219 3116 2220
rect 3110 2218 3111 2219
rect 3100 2216 3111 2218
rect 3100 2215 3101 2216
rect 3095 2214 3101 2215
rect 3110 2215 3111 2216
rect 3115 2215 3116 2219
rect 3110 2214 3116 2215
rect 3287 2219 3293 2220
rect 3287 2215 3288 2219
rect 3292 2218 3293 2219
rect 3295 2219 3301 2220
rect 3295 2218 3296 2219
rect 3292 2216 3296 2218
rect 3292 2215 3293 2216
rect 3287 2214 3293 2215
rect 3295 2215 3296 2216
rect 3300 2215 3301 2219
rect 3295 2214 3301 2215
rect 3470 2219 3476 2220
rect 3470 2215 3471 2219
rect 3475 2218 3476 2219
rect 3479 2219 3485 2220
rect 3479 2218 3480 2219
rect 3475 2216 3480 2218
rect 3475 2215 3476 2216
rect 3470 2214 3476 2215
rect 3479 2215 3480 2216
rect 3484 2215 3485 2219
rect 3479 2214 3485 2215
rect 1726 2210 1732 2211
rect 2006 2209 2012 2210
rect 1030 2207 1036 2208
rect 110 2205 116 2206
rect 110 2201 111 2205
rect 115 2201 116 2205
rect 1030 2203 1031 2207
rect 1035 2206 1036 2207
rect 1642 2207 1648 2208
rect 1035 2204 1089 2206
rect 1035 2203 1036 2204
rect 1030 2202 1036 2203
rect 1642 2203 1643 2207
rect 1647 2206 1648 2207
rect 1647 2204 1745 2206
rect 1822 2205 1828 2206
rect 1647 2203 1648 2204
rect 1642 2202 1648 2203
rect 110 2200 116 2201
rect 1822 2201 1823 2205
rect 1827 2201 1828 2205
rect 2006 2205 2007 2209
rect 2011 2205 2012 2209
rect 2006 2204 2012 2205
rect 2166 2209 2172 2210
rect 2166 2205 2167 2209
rect 2171 2205 2172 2209
rect 2166 2204 2172 2205
rect 2334 2209 2340 2210
rect 2334 2205 2335 2209
rect 2339 2205 2340 2209
rect 2334 2204 2340 2205
rect 2518 2209 2524 2210
rect 2518 2205 2519 2209
rect 2523 2205 2524 2209
rect 2518 2204 2524 2205
rect 2710 2209 2716 2210
rect 2710 2205 2711 2209
rect 2715 2205 2716 2209
rect 2710 2204 2716 2205
rect 2902 2209 2908 2210
rect 2902 2205 2903 2209
rect 2907 2205 2908 2209
rect 2902 2204 2908 2205
rect 3102 2209 3108 2210
rect 3102 2205 3103 2209
rect 3107 2205 3108 2209
rect 3102 2204 3108 2205
rect 3302 2209 3308 2210
rect 3302 2205 3303 2209
rect 3307 2205 3308 2209
rect 3302 2204 3308 2205
rect 3486 2209 3492 2210
rect 3486 2205 3487 2209
rect 3491 2205 3492 2209
rect 3486 2204 3492 2205
rect 1822 2200 1828 2201
rect 1862 2196 1868 2197
rect 3574 2196 3580 2197
rect 1862 2192 1863 2196
rect 1867 2192 1868 2196
rect 2087 2195 2093 2196
rect 2087 2194 2088 2195
rect 2061 2192 2088 2194
rect 711 2191 717 2192
rect 711 2190 712 2191
rect 110 2188 116 2189
rect 597 2188 712 2190
rect 110 2184 111 2188
rect 115 2184 116 2188
rect 711 2187 712 2188
rect 716 2187 717 2191
rect 887 2191 893 2192
rect 887 2190 888 2191
rect 781 2188 888 2190
rect 711 2186 717 2187
rect 887 2187 888 2188
rect 892 2187 893 2191
rect 1063 2191 1069 2192
rect 1063 2190 1064 2191
rect 957 2188 1064 2190
rect 887 2186 893 2187
rect 1063 2187 1064 2188
rect 1068 2187 1069 2191
rect 1399 2191 1405 2192
rect 1399 2190 1400 2191
rect 1301 2188 1400 2190
rect 1063 2186 1069 2187
rect 1399 2187 1400 2188
rect 1404 2187 1405 2191
rect 1567 2191 1573 2192
rect 1567 2190 1568 2191
rect 1469 2188 1568 2190
rect 1399 2186 1405 2187
rect 1567 2187 1568 2188
rect 1572 2187 1573 2191
rect 1719 2191 1725 2192
rect 1862 2191 1868 2192
rect 2087 2191 2088 2192
rect 2092 2191 2093 2195
rect 2239 2195 2245 2196
rect 2239 2194 2240 2195
rect 2221 2192 2240 2194
rect 1719 2190 1720 2191
rect 1637 2188 1720 2190
rect 1567 2186 1573 2187
rect 1719 2187 1720 2188
rect 1724 2187 1725 2191
rect 2087 2190 2093 2191
rect 2239 2191 2240 2192
rect 2244 2191 2245 2195
rect 3287 2195 3293 2196
rect 3287 2194 3288 2195
rect 3157 2192 3288 2194
rect 2239 2190 2245 2191
rect 2402 2191 2408 2192
rect 1719 2186 1725 2187
rect 1822 2188 1828 2189
rect 110 2183 116 2184
rect 1822 2184 1823 2188
rect 1827 2184 1828 2188
rect 2402 2187 2403 2191
rect 2407 2190 2408 2191
rect 2586 2191 2592 2192
rect 2407 2188 2537 2190
rect 2407 2187 2408 2188
rect 2402 2186 2408 2187
rect 2586 2187 2587 2191
rect 2591 2190 2592 2191
rect 2807 2191 2813 2192
rect 2591 2188 2729 2190
rect 2591 2187 2592 2188
rect 2586 2186 2592 2187
rect 2807 2187 2808 2191
rect 2812 2190 2813 2191
rect 3287 2191 3288 2192
rect 3292 2191 3293 2195
rect 3367 2195 3373 2196
rect 3367 2194 3368 2195
rect 3357 2192 3368 2194
rect 3287 2190 3293 2191
rect 3367 2191 3368 2192
rect 3372 2191 3373 2195
rect 3574 2192 3575 2196
rect 3579 2192 3580 2196
rect 3574 2191 3580 2192
rect 3367 2190 3373 2191
rect 2812 2188 2921 2190
rect 2812 2187 2813 2188
rect 2807 2186 2813 2187
rect 1822 2183 1828 2184
rect 1862 2179 1868 2180
rect 542 2175 548 2176
rect 542 2171 543 2175
rect 547 2171 548 2175
rect 542 2170 548 2171
rect 726 2175 732 2176
rect 726 2171 727 2175
rect 731 2171 732 2175
rect 726 2170 732 2171
rect 902 2175 908 2176
rect 902 2171 903 2175
rect 907 2171 908 2175
rect 902 2170 908 2171
rect 1078 2175 1084 2176
rect 1078 2171 1079 2175
rect 1083 2171 1084 2175
rect 1078 2170 1084 2171
rect 1246 2175 1252 2176
rect 1246 2171 1247 2175
rect 1251 2171 1252 2175
rect 1246 2170 1252 2171
rect 1414 2175 1420 2176
rect 1414 2171 1415 2175
rect 1419 2171 1420 2175
rect 1414 2170 1420 2171
rect 1582 2175 1588 2176
rect 1582 2171 1583 2175
rect 1587 2171 1588 2175
rect 1582 2170 1588 2171
rect 1734 2175 1740 2176
rect 1734 2171 1735 2175
rect 1739 2171 1740 2175
rect 1862 2175 1863 2179
rect 1867 2175 1868 2179
rect 1862 2174 1868 2175
rect 2234 2179 2240 2180
rect 2234 2175 2235 2179
rect 2239 2178 2240 2179
rect 3471 2179 3477 2180
rect 2239 2176 2345 2178
rect 2239 2175 2240 2176
rect 2234 2174 2240 2175
rect 3471 2175 3472 2179
rect 3476 2178 3477 2179
rect 3574 2179 3580 2180
rect 3476 2176 3497 2178
rect 3476 2175 3477 2176
rect 3471 2174 3477 2175
rect 3574 2175 3575 2179
rect 3579 2175 3580 2179
rect 3574 2174 3580 2175
rect 1734 2170 1740 2171
rect 1998 2169 2004 2170
rect 1998 2165 1999 2169
rect 2003 2165 2004 2169
rect 1998 2164 2004 2165
rect 2158 2169 2164 2170
rect 2158 2165 2159 2169
rect 2163 2165 2164 2169
rect 2158 2164 2164 2165
rect 2326 2169 2332 2170
rect 2326 2165 2327 2169
rect 2331 2165 2332 2169
rect 2326 2164 2332 2165
rect 2510 2169 2516 2170
rect 2510 2165 2511 2169
rect 2515 2165 2516 2169
rect 2510 2164 2516 2165
rect 2702 2169 2708 2170
rect 2702 2165 2703 2169
rect 2707 2165 2708 2169
rect 2702 2164 2708 2165
rect 2894 2169 2900 2170
rect 2894 2165 2895 2169
rect 2899 2165 2900 2169
rect 2894 2164 2900 2165
rect 3094 2169 3100 2170
rect 3094 2165 3095 2169
rect 3099 2165 3100 2169
rect 3094 2164 3100 2165
rect 3294 2169 3300 2170
rect 3294 2165 3295 2169
rect 3299 2165 3300 2169
rect 3294 2164 3300 2165
rect 3478 2169 3484 2170
rect 3478 2165 3479 2169
rect 3483 2165 3484 2169
rect 3478 2164 3484 2165
rect 535 2163 541 2164
rect 535 2159 536 2163
rect 540 2162 541 2163
rect 574 2163 580 2164
rect 574 2162 575 2163
rect 540 2160 575 2162
rect 540 2159 541 2160
rect 535 2158 541 2159
rect 574 2159 575 2160
rect 579 2159 580 2163
rect 574 2158 580 2159
rect 711 2163 717 2164
rect 711 2159 712 2163
rect 716 2162 717 2163
rect 719 2163 725 2164
rect 719 2162 720 2163
rect 716 2160 720 2162
rect 716 2159 717 2160
rect 711 2158 717 2159
rect 719 2159 720 2160
rect 724 2159 725 2163
rect 719 2158 725 2159
rect 887 2163 893 2164
rect 887 2159 888 2163
rect 892 2162 893 2163
rect 895 2163 901 2164
rect 895 2162 896 2163
rect 892 2160 896 2162
rect 892 2159 893 2160
rect 887 2158 893 2159
rect 895 2159 896 2160
rect 900 2159 901 2163
rect 895 2158 901 2159
rect 1063 2163 1069 2164
rect 1063 2159 1064 2163
rect 1068 2162 1069 2163
rect 1071 2163 1077 2164
rect 1071 2162 1072 2163
rect 1068 2160 1072 2162
rect 1068 2159 1069 2160
rect 1063 2158 1069 2159
rect 1071 2159 1072 2160
rect 1076 2159 1077 2163
rect 1071 2158 1077 2159
rect 1239 2163 1245 2164
rect 1239 2159 1240 2163
rect 1244 2162 1245 2163
rect 1254 2163 1260 2164
rect 1254 2162 1255 2163
rect 1244 2160 1255 2162
rect 1244 2159 1245 2160
rect 1239 2158 1245 2159
rect 1254 2159 1255 2160
rect 1259 2159 1260 2163
rect 1254 2158 1260 2159
rect 1399 2163 1405 2164
rect 1399 2159 1400 2163
rect 1404 2162 1405 2163
rect 1407 2163 1413 2164
rect 1407 2162 1408 2163
rect 1404 2160 1408 2162
rect 1404 2159 1405 2160
rect 1399 2158 1405 2159
rect 1407 2159 1408 2160
rect 1412 2159 1413 2163
rect 1407 2158 1413 2159
rect 1567 2163 1573 2164
rect 1567 2159 1568 2163
rect 1572 2162 1573 2163
rect 1575 2163 1581 2164
rect 1575 2162 1576 2163
rect 1572 2160 1576 2162
rect 1572 2159 1573 2160
rect 1567 2158 1573 2159
rect 1575 2159 1576 2160
rect 1580 2159 1581 2163
rect 1575 2158 1581 2159
rect 1719 2163 1725 2164
rect 1719 2159 1720 2163
rect 1724 2162 1725 2163
rect 1727 2163 1733 2164
rect 1727 2162 1728 2163
rect 1724 2160 1728 2162
rect 1724 2159 1725 2160
rect 1719 2158 1725 2159
rect 1727 2159 1728 2160
rect 1732 2159 1733 2163
rect 1727 2158 1733 2159
rect 487 2151 493 2152
rect 487 2147 488 2151
rect 492 2150 493 2151
rect 550 2151 556 2152
rect 550 2150 551 2151
rect 492 2148 551 2150
rect 492 2147 493 2148
rect 487 2146 493 2147
rect 550 2147 551 2148
rect 555 2147 556 2151
rect 550 2146 556 2147
rect 559 2151 565 2152
rect 559 2147 560 2151
rect 564 2150 565 2151
rect 615 2151 621 2152
rect 615 2150 616 2151
rect 564 2148 616 2150
rect 564 2147 565 2148
rect 559 2146 565 2147
rect 615 2147 616 2148
rect 620 2147 621 2151
rect 615 2146 621 2147
rect 687 2151 693 2152
rect 687 2147 688 2151
rect 692 2150 693 2151
rect 751 2151 757 2152
rect 751 2150 752 2151
rect 692 2148 752 2150
rect 692 2147 693 2148
rect 687 2146 693 2147
rect 751 2147 752 2148
rect 756 2147 757 2151
rect 751 2146 757 2147
rect 823 2151 829 2152
rect 823 2147 824 2151
rect 828 2150 829 2151
rect 887 2151 893 2152
rect 887 2150 888 2151
rect 828 2148 888 2150
rect 828 2147 829 2148
rect 823 2146 829 2147
rect 887 2147 888 2148
rect 892 2147 893 2151
rect 887 2146 893 2147
rect 967 2151 973 2152
rect 967 2147 968 2151
rect 972 2150 973 2151
rect 1031 2151 1037 2152
rect 1031 2150 1032 2151
rect 972 2148 1032 2150
rect 972 2147 973 2148
rect 967 2146 973 2147
rect 1031 2147 1032 2148
rect 1036 2147 1037 2151
rect 1031 2146 1037 2147
rect 1175 2151 1181 2152
rect 1175 2147 1176 2151
rect 1180 2150 1181 2151
rect 1238 2151 1244 2152
rect 1238 2150 1239 2151
rect 1180 2148 1239 2150
rect 1180 2147 1181 2148
rect 1175 2146 1181 2147
rect 1238 2147 1239 2148
rect 1243 2147 1244 2151
rect 1238 2146 1244 2147
rect 1255 2151 1261 2152
rect 1255 2147 1256 2151
rect 1260 2150 1261 2151
rect 1319 2151 1325 2152
rect 1319 2150 1320 2151
rect 1260 2148 1320 2150
rect 1260 2147 1261 2148
rect 1255 2146 1261 2147
rect 1319 2147 1320 2148
rect 1324 2147 1325 2151
rect 1319 2146 1325 2147
rect 1463 2151 1469 2152
rect 1463 2147 1464 2151
rect 1468 2150 1469 2151
rect 1538 2151 1544 2152
rect 1538 2150 1539 2151
rect 1468 2148 1539 2150
rect 1468 2147 1469 2148
rect 1463 2146 1469 2147
rect 1538 2147 1539 2148
rect 1543 2147 1544 2151
rect 1538 2146 1544 2147
rect 1615 2151 1621 2152
rect 1615 2147 1616 2151
rect 1620 2150 1621 2151
rect 1642 2151 1648 2152
rect 1642 2150 1643 2151
rect 1620 2148 1643 2150
rect 1620 2147 1621 2148
rect 1615 2146 1621 2147
rect 1642 2147 1643 2148
rect 1647 2147 1648 2151
rect 1642 2146 1648 2147
rect 494 2141 500 2142
rect 494 2137 495 2141
rect 499 2137 500 2141
rect 494 2136 500 2137
rect 622 2141 628 2142
rect 622 2137 623 2141
rect 627 2137 628 2141
rect 622 2136 628 2137
rect 758 2141 764 2142
rect 758 2137 759 2141
rect 763 2137 764 2141
rect 758 2136 764 2137
rect 894 2141 900 2142
rect 894 2137 895 2141
rect 899 2137 900 2141
rect 894 2136 900 2137
rect 1038 2141 1044 2142
rect 1038 2137 1039 2141
rect 1043 2137 1044 2141
rect 1038 2136 1044 2137
rect 1182 2141 1188 2142
rect 1182 2137 1183 2141
rect 1187 2137 1188 2141
rect 1182 2136 1188 2137
rect 1326 2141 1332 2142
rect 1326 2137 1327 2141
rect 1331 2137 1332 2141
rect 1326 2136 1332 2137
rect 1470 2141 1476 2142
rect 1470 2137 1471 2141
rect 1475 2137 1476 2141
rect 1470 2136 1476 2137
rect 1622 2141 1628 2142
rect 1622 2137 1623 2141
rect 1627 2137 1628 2141
rect 1622 2136 1628 2137
rect 2022 2139 2028 2140
rect 2022 2135 2023 2139
rect 2027 2135 2028 2139
rect 2022 2134 2028 2135
rect 2166 2139 2172 2140
rect 2166 2135 2167 2139
rect 2171 2135 2172 2139
rect 2166 2134 2172 2135
rect 2318 2139 2324 2140
rect 2318 2135 2319 2139
rect 2323 2135 2324 2139
rect 2318 2134 2324 2135
rect 2470 2139 2476 2140
rect 2470 2135 2471 2139
rect 2475 2135 2476 2139
rect 2470 2134 2476 2135
rect 2614 2139 2620 2140
rect 2614 2135 2615 2139
rect 2619 2135 2620 2139
rect 2614 2134 2620 2135
rect 2758 2139 2764 2140
rect 2758 2135 2759 2139
rect 2763 2135 2764 2139
rect 2758 2134 2764 2135
rect 2894 2139 2900 2140
rect 2894 2135 2895 2139
rect 2899 2135 2900 2139
rect 2894 2134 2900 2135
rect 3022 2139 3028 2140
rect 3022 2135 3023 2139
rect 3027 2135 3028 2139
rect 3022 2134 3028 2135
rect 3142 2139 3148 2140
rect 3142 2135 3143 2139
rect 3147 2135 3148 2139
rect 3142 2134 3148 2135
rect 3262 2139 3268 2140
rect 3262 2135 3263 2139
rect 3267 2135 3268 2139
rect 3262 2134 3268 2135
rect 3382 2139 3388 2140
rect 3382 2135 3383 2139
rect 3387 2135 3388 2139
rect 3382 2134 3388 2135
rect 3478 2139 3484 2140
rect 3478 2135 3479 2139
rect 3483 2135 3484 2139
rect 3478 2134 3484 2135
rect 2838 2131 2844 2132
rect 2838 2130 2839 2131
rect 1862 2129 1868 2130
rect 110 2128 116 2129
rect 1822 2128 1828 2129
rect 110 2124 111 2128
rect 115 2124 116 2128
rect 559 2127 565 2128
rect 559 2126 560 2127
rect 549 2124 560 2126
rect 110 2123 116 2124
rect 559 2123 560 2124
rect 564 2123 565 2127
rect 687 2127 693 2128
rect 687 2126 688 2127
rect 677 2124 688 2126
rect 559 2122 565 2123
rect 687 2123 688 2124
rect 692 2123 693 2127
rect 823 2127 829 2128
rect 823 2126 824 2127
rect 813 2124 824 2126
rect 687 2122 693 2123
rect 823 2123 824 2124
rect 828 2123 829 2127
rect 967 2127 973 2128
rect 967 2126 968 2127
rect 949 2124 968 2126
rect 823 2122 829 2123
rect 967 2123 968 2124
rect 972 2123 973 2127
rect 1255 2127 1261 2128
rect 1255 2126 1256 2127
rect 1237 2124 1256 2126
rect 967 2122 973 2123
rect 1255 2123 1256 2124
rect 1260 2123 1261 2127
rect 1822 2124 1823 2128
rect 1827 2124 1828 2128
rect 1862 2125 1863 2129
rect 1867 2125 1868 2129
rect 2817 2128 2839 2130
rect 2838 2127 2839 2128
rect 2843 2127 2844 2131
rect 2838 2126 2844 2127
rect 3450 2131 3456 2132
rect 3450 2127 3451 2131
rect 3455 2130 3456 2131
rect 3455 2128 3497 2130
rect 3574 2129 3580 2130
rect 3455 2127 3456 2128
rect 3450 2126 3456 2127
rect 1862 2124 1868 2125
rect 3574 2125 3575 2129
rect 3579 2125 3580 2129
rect 3574 2124 3580 2125
rect 1255 2122 1261 2123
rect 1399 2123 1405 2124
rect 1399 2119 1400 2123
rect 1404 2122 1405 2123
rect 1538 2123 1544 2124
rect 1822 2123 1828 2124
rect 1404 2120 1489 2122
rect 1404 2119 1405 2120
rect 1399 2118 1405 2119
rect 1538 2119 1539 2123
rect 1543 2122 1544 2123
rect 1543 2120 1641 2122
rect 1543 2119 1544 2120
rect 1538 2118 1544 2119
rect 1983 2115 1989 2116
rect 1862 2112 1868 2113
rect 110 2111 116 2112
rect 110 2107 111 2111
rect 115 2107 116 2111
rect 110 2106 116 2107
rect 1038 2111 1044 2112
rect 1038 2107 1039 2111
rect 1043 2110 1044 2111
rect 1398 2111 1404 2112
rect 1398 2110 1399 2111
rect 1043 2108 1049 2110
rect 1377 2108 1399 2110
rect 1043 2107 1044 2108
rect 1038 2106 1044 2107
rect 1398 2107 1399 2108
rect 1403 2107 1404 2111
rect 1398 2106 1404 2107
rect 1822 2111 1828 2112
rect 1822 2107 1823 2111
rect 1827 2107 1828 2111
rect 1862 2108 1863 2112
rect 1867 2108 1868 2112
rect 1983 2111 1984 2115
rect 1988 2114 1989 2115
rect 2106 2115 2112 2116
rect 1988 2112 2049 2114
rect 1988 2111 1989 2112
rect 1983 2110 1989 2111
rect 2106 2111 2107 2115
rect 2111 2114 2112 2115
rect 2463 2115 2469 2116
rect 2463 2114 2464 2115
rect 2111 2112 2193 2114
rect 2381 2112 2464 2114
rect 2111 2111 2112 2112
rect 2106 2110 2112 2111
rect 2463 2111 2464 2112
rect 2468 2111 2469 2115
rect 2607 2115 2613 2116
rect 2607 2114 2608 2115
rect 2533 2112 2608 2114
rect 2463 2110 2469 2111
rect 2607 2111 2608 2112
rect 2612 2111 2613 2115
rect 2751 2115 2757 2116
rect 2751 2114 2752 2115
rect 2677 2112 2752 2114
rect 2607 2110 2613 2111
rect 2751 2111 2752 2112
rect 2756 2111 2757 2115
rect 2751 2110 2757 2111
rect 2826 2115 2832 2116
rect 2826 2111 2827 2115
rect 2831 2114 2832 2115
rect 2962 2115 2968 2116
rect 2831 2112 2921 2114
rect 2831 2111 2832 2112
rect 2826 2110 2832 2111
rect 2962 2111 2963 2115
rect 2967 2114 2968 2115
rect 3090 2115 3096 2116
rect 2967 2112 3049 2114
rect 2967 2111 2968 2112
rect 2962 2110 2968 2111
rect 3090 2111 3091 2115
rect 3095 2114 3096 2115
rect 3210 2115 3216 2116
rect 3095 2112 3169 2114
rect 3095 2111 3096 2112
rect 3090 2110 3096 2111
rect 3210 2111 3211 2115
rect 3215 2114 3216 2115
rect 3470 2115 3476 2116
rect 3470 2114 3471 2115
rect 3215 2112 3289 2114
rect 3445 2112 3471 2114
rect 3215 2111 3216 2112
rect 3210 2110 3216 2111
rect 3470 2111 3471 2112
rect 3475 2111 3476 2115
rect 3470 2110 3476 2111
rect 3574 2112 3580 2113
rect 1862 2107 1868 2108
rect 3574 2108 3575 2112
rect 3579 2108 3580 2112
rect 3574 2107 3580 2108
rect 1822 2106 1828 2107
rect 486 2101 492 2102
rect 486 2097 487 2101
rect 491 2097 492 2101
rect 486 2096 492 2097
rect 614 2101 620 2102
rect 614 2097 615 2101
rect 619 2097 620 2101
rect 614 2096 620 2097
rect 750 2101 756 2102
rect 750 2097 751 2101
rect 755 2097 756 2101
rect 750 2096 756 2097
rect 886 2101 892 2102
rect 886 2097 887 2101
rect 891 2097 892 2101
rect 886 2096 892 2097
rect 1030 2101 1036 2102
rect 1030 2097 1031 2101
rect 1035 2097 1036 2101
rect 1030 2096 1036 2097
rect 1174 2101 1180 2102
rect 1174 2097 1175 2101
rect 1179 2097 1180 2101
rect 1174 2096 1180 2097
rect 1318 2101 1324 2102
rect 1318 2097 1319 2101
rect 1323 2097 1324 2101
rect 1318 2096 1324 2097
rect 1462 2101 1468 2102
rect 1462 2097 1463 2101
rect 1467 2097 1468 2101
rect 1462 2096 1468 2097
rect 1614 2101 1620 2102
rect 1614 2097 1615 2101
rect 1619 2097 1620 2101
rect 1614 2096 1620 2097
rect 2030 2099 2036 2100
rect 1238 2095 1244 2096
rect 1238 2091 1239 2095
rect 1243 2094 1244 2095
rect 1399 2095 1405 2096
rect 1399 2094 1400 2095
rect 1243 2092 1400 2094
rect 1243 2091 1244 2092
rect 1238 2090 1244 2091
rect 1399 2091 1400 2092
rect 1404 2091 1405 2095
rect 2030 2095 2031 2099
rect 2035 2095 2036 2099
rect 2030 2094 2036 2095
rect 2174 2099 2180 2100
rect 2174 2095 2175 2099
rect 2179 2095 2180 2099
rect 2174 2094 2180 2095
rect 2326 2099 2332 2100
rect 2326 2095 2327 2099
rect 2331 2095 2332 2099
rect 2326 2094 2332 2095
rect 2478 2099 2484 2100
rect 2478 2095 2479 2099
rect 2483 2095 2484 2099
rect 2478 2094 2484 2095
rect 2622 2099 2628 2100
rect 2622 2095 2623 2099
rect 2627 2095 2628 2099
rect 2622 2094 2628 2095
rect 2766 2099 2772 2100
rect 2766 2095 2767 2099
rect 2771 2095 2772 2099
rect 2766 2094 2772 2095
rect 2902 2099 2908 2100
rect 2902 2095 2903 2099
rect 2907 2095 2908 2099
rect 2902 2094 2908 2095
rect 3030 2099 3036 2100
rect 3030 2095 3031 2099
rect 3035 2095 3036 2099
rect 3030 2094 3036 2095
rect 3150 2099 3156 2100
rect 3150 2095 3151 2099
rect 3155 2095 3156 2099
rect 3150 2094 3156 2095
rect 3270 2099 3276 2100
rect 3270 2095 3271 2099
rect 3275 2095 3276 2099
rect 3270 2094 3276 2095
rect 3390 2099 3396 2100
rect 3390 2095 3391 2099
rect 3395 2095 3396 2099
rect 3390 2094 3396 2095
rect 3486 2099 3492 2100
rect 3486 2095 3487 2099
rect 3491 2095 3492 2099
rect 3486 2094 3492 2095
rect 1399 2090 1405 2091
rect 2023 2087 2029 2088
rect 2023 2083 2024 2087
rect 2028 2086 2029 2087
rect 2106 2087 2112 2088
rect 2106 2086 2107 2087
rect 2028 2084 2107 2086
rect 2028 2083 2029 2084
rect 2023 2082 2029 2083
rect 2106 2083 2107 2084
rect 2111 2083 2112 2087
rect 2106 2082 2112 2083
rect 2167 2087 2173 2088
rect 2167 2083 2168 2087
rect 2172 2086 2173 2087
rect 2234 2087 2240 2088
rect 2234 2086 2235 2087
rect 2172 2084 2235 2086
rect 2172 2083 2173 2084
rect 2167 2082 2173 2083
rect 2234 2083 2235 2084
rect 2239 2083 2240 2087
rect 2234 2082 2240 2083
rect 2302 2087 2308 2088
rect 2302 2083 2303 2087
rect 2307 2086 2308 2087
rect 2319 2087 2325 2088
rect 2319 2086 2320 2087
rect 2307 2084 2320 2086
rect 2307 2083 2308 2084
rect 2302 2082 2308 2083
rect 2319 2083 2320 2084
rect 2324 2083 2325 2087
rect 2319 2082 2325 2083
rect 2463 2087 2469 2088
rect 2463 2083 2464 2087
rect 2468 2086 2469 2087
rect 2471 2087 2477 2088
rect 2471 2086 2472 2087
rect 2468 2084 2472 2086
rect 2468 2083 2469 2084
rect 2463 2082 2469 2083
rect 2471 2083 2472 2084
rect 2476 2083 2477 2087
rect 2471 2082 2477 2083
rect 2607 2087 2613 2088
rect 2607 2083 2608 2087
rect 2612 2086 2613 2087
rect 2615 2087 2621 2088
rect 2615 2086 2616 2087
rect 2612 2084 2616 2086
rect 2612 2083 2613 2084
rect 2607 2082 2613 2083
rect 2615 2083 2616 2084
rect 2620 2083 2621 2087
rect 2615 2082 2621 2083
rect 2751 2087 2757 2088
rect 2751 2083 2752 2087
rect 2756 2086 2757 2087
rect 2759 2087 2765 2088
rect 2759 2086 2760 2087
rect 2756 2084 2760 2086
rect 2756 2083 2757 2084
rect 2751 2082 2757 2083
rect 2759 2083 2760 2084
rect 2764 2083 2765 2087
rect 2759 2082 2765 2083
rect 2895 2087 2901 2088
rect 2895 2083 2896 2087
rect 2900 2086 2901 2087
rect 2962 2087 2968 2088
rect 2962 2086 2963 2087
rect 2900 2084 2963 2086
rect 2900 2083 2901 2084
rect 2895 2082 2901 2083
rect 2962 2083 2963 2084
rect 2967 2083 2968 2087
rect 2962 2082 2968 2083
rect 3023 2087 3029 2088
rect 3023 2083 3024 2087
rect 3028 2086 3029 2087
rect 3090 2087 3096 2088
rect 3090 2086 3091 2087
rect 3028 2084 3091 2086
rect 3028 2083 3029 2084
rect 3023 2082 3029 2083
rect 3090 2083 3091 2084
rect 3095 2083 3096 2087
rect 3090 2082 3096 2083
rect 3143 2087 3149 2088
rect 3143 2083 3144 2087
rect 3148 2086 3149 2087
rect 3210 2087 3216 2088
rect 3210 2086 3211 2087
rect 3148 2084 3211 2086
rect 3148 2083 3149 2084
rect 3143 2082 3149 2083
rect 3210 2083 3211 2084
rect 3215 2083 3216 2087
rect 3210 2082 3216 2083
rect 3223 2087 3229 2088
rect 3223 2083 3224 2087
rect 3228 2086 3229 2087
rect 3263 2087 3269 2088
rect 3263 2086 3264 2087
rect 3228 2084 3264 2086
rect 3228 2083 3229 2084
rect 3223 2082 3229 2083
rect 3263 2083 3264 2084
rect 3268 2083 3269 2087
rect 3263 2082 3269 2083
rect 3383 2087 3389 2088
rect 3383 2083 3384 2087
rect 3388 2086 3389 2087
rect 3450 2087 3456 2088
rect 3450 2086 3451 2087
rect 3388 2084 3451 2086
rect 3388 2083 3389 2084
rect 3383 2082 3389 2083
rect 3450 2083 3451 2084
rect 3455 2083 3456 2087
rect 3450 2082 3456 2083
rect 3471 2087 3477 2088
rect 3471 2083 3472 2087
rect 3476 2086 3477 2087
rect 3479 2087 3485 2088
rect 3479 2086 3480 2087
rect 3476 2084 3480 2086
rect 3476 2083 3477 2084
rect 3471 2082 3477 2083
rect 3479 2083 3480 2084
rect 3484 2083 3485 2087
rect 3479 2082 3485 2083
rect 3231 2079 3237 2080
rect 3231 2078 3232 2079
rect 3088 2076 3232 2078
rect 318 2075 324 2076
rect 318 2071 319 2075
rect 323 2071 324 2075
rect 318 2070 324 2071
rect 430 2075 436 2076
rect 430 2071 431 2075
rect 435 2071 436 2075
rect 430 2070 436 2071
rect 550 2075 556 2076
rect 550 2071 551 2075
rect 555 2071 556 2075
rect 550 2070 556 2071
rect 678 2075 684 2076
rect 678 2071 679 2075
rect 683 2071 684 2075
rect 678 2070 684 2071
rect 798 2075 804 2076
rect 798 2071 799 2075
rect 803 2071 804 2075
rect 798 2070 804 2071
rect 918 2075 924 2076
rect 918 2071 919 2075
rect 923 2071 924 2075
rect 918 2070 924 2071
rect 1038 2075 1044 2076
rect 1038 2071 1039 2075
rect 1043 2071 1044 2075
rect 1038 2070 1044 2071
rect 1158 2075 1164 2076
rect 1158 2071 1159 2075
rect 1163 2071 1164 2075
rect 1158 2070 1164 2071
rect 1278 2075 1284 2076
rect 1278 2071 1279 2075
rect 1283 2071 1284 2075
rect 1278 2070 1284 2071
rect 1406 2075 1412 2076
rect 1406 2071 1407 2075
rect 1411 2071 1412 2075
rect 1406 2070 1412 2071
rect 1975 2071 1981 2072
rect 766 2067 772 2068
rect 110 2065 116 2066
rect 110 2061 111 2065
rect 115 2061 116 2065
rect 766 2063 767 2067
rect 771 2066 772 2067
rect 1975 2067 1976 2071
rect 1980 2070 1981 2071
rect 1983 2071 1989 2072
rect 1983 2070 1984 2071
rect 1980 2068 1984 2070
rect 1980 2067 1981 2068
rect 1975 2066 1981 2067
rect 1983 2067 1984 2068
rect 1988 2067 1989 2071
rect 1983 2066 1989 2067
rect 2063 2071 2069 2072
rect 2063 2067 2064 2071
rect 2068 2070 2069 2071
rect 2135 2071 2141 2072
rect 2135 2070 2136 2071
rect 2068 2068 2136 2070
rect 2068 2067 2069 2068
rect 2063 2066 2069 2067
rect 2135 2067 2136 2068
rect 2140 2067 2141 2071
rect 2135 2066 2141 2067
rect 2303 2071 2309 2072
rect 2303 2067 2304 2071
rect 2308 2070 2309 2071
rect 2391 2071 2397 2072
rect 2391 2070 2392 2071
rect 2308 2068 2392 2070
rect 2308 2067 2309 2068
rect 2303 2066 2309 2067
rect 2391 2067 2392 2068
rect 2396 2067 2397 2071
rect 2391 2066 2397 2067
rect 2463 2071 2469 2072
rect 2463 2067 2464 2071
rect 2468 2070 2469 2071
rect 2551 2071 2557 2072
rect 2551 2070 2552 2071
rect 2468 2068 2552 2070
rect 2468 2067 2469 2068
rect 2463 2066 2469 2067
rect 2551 2067 2552 2068
rect 2556 2067 2557 2071
rect 2551 2066 2557 2067
rect 2610 2071 2616 2072
rect 2610 2067 2611 2071
rect 2615 2070 2616 2071
rect 2623 2071 2629 2072
rect 2623 2070 2624 2071
rect 2615 2068 2624 2070
rect 2615 2067 2616 2068
rect 2610 2066 2616 2067
rect 2623 2067 2624 2068
rect 2628 2067 2629 2071
rect 2623 2066 2629 2067
rect 2767 2071 2773 2072
rect 2767 2067 2768 2071
rect 2772 2070 2773 2071
rect 2826 2071 2832 2072
rect 2826 2070 2827 2071
rect 2772 2068 2827 2070
rect 2772 2067 2773 2068
rect 2767 2066 2773 2067
rect 2826 2067 2827 2068
rect 2831 2067 2832 2071
rect 2826 2066 2832 2067
rect 2839 2071 2845 2072
rect 2839 2067 2840 2071
rect 2844 2070 2845 2071
rect 2903 2071 2909 2072
rect 2903 2070 2904 2071
rect 2844 2068 2904 2070
rect 2844 2067 2845 2068
rect 2839 2066 2845 2067
rect 2903 2067 2904 2068
rect 2908 2067 2909 2071
rect 2903 2066 2909 2067
rect 3031 2071 3037 2072
rect 3031 2067 3032 2071
rect 3036 2070 3037 2071
rect 3088 2070 3090 2076
rect 3231 2075 3232 2076
rect 3236 2075 3237 2079
rect 3231 2074 3237 2075
rect 3036 2068 3090 2070
rect 3103 2071 3109 2072
rect 3036 2067 3037 2068
rect 3031 2066 3037 2067
rect 3103 2067 3104 2071
rect 3108 2070 3109 2071
rect 3151 2071 3157 2072
rect 3151 2070 3152 2071
rect 3108 2068 3152 2070
rect 3108 2067 3109 2068
rect 3103 2066 3109 2067
rect 3151 2067 3152 2068
rect 3156 2067 3157 2071
rect 3151 2066 3157 2067
rect 3271 2071 3277 2072
rect 3271 2067 3272 2071
rect 3276 2070 3277 2071
rect 3346 2071 3352 2072
rect 3346 2070 3347 2071
rect 3276 2068 3347 2070
rect 3276 2067 3277 2068
rect 3271 2066 3277 2067
rect 3346 2067 3347 2068
rect 3351 2067 3352 2071
rect 3346 2066 3352 2067
rect 3383 2071 3389 2072
rect 3383 2067 3384 2071
rect 3388 2070 3389 2071
rect 3458 2071 3464 2072
rect 3458 2070 3459 2071
rect 3388 2068 3459 2070
rect 3388 2067 3389 2068
rect 3383 2066 3389 2067
rect 3458 2067 3459 2068
rect 3463 2067 3464 2071
rect 3458 2066 3464 2067
rect 3470 2071 3476 2072
rect 3470 2067 3471 2071
rect 3475 2070 3476 2071
rect 3479 2071 3485 2072
rect 3479 2070 3480 2071
rect 3475 2068 3480 2070
rect 3475 2067 3476 2068
rect 3470 2066 3476 2067
rect 3479 2067 3480 2068
rect 3484 2067 3485 2071
rect 3479 2066 3485 2067
rect 771 2064 817 2066
rect 1822 2065 1828 2066
rect 771 2063 772 2064
rect 766 2062 772 2063
rect 110 2060 116 2061
rect 1822 2061 1823 2065
rect 1827 2061 1828 2065
rect 1822 2060 1828 2061
rect 1982 2061 1988 2062
rect 1982 2057 1983 2061
rect 1987 2057 1988 2061
rect 1982 2056 1988 2057
rect 2142 2061 2148 2062
rect 2142 2057 2143 2061
rect 2147 2057 2148 2061
rect 2142 2056 2148 2057
rect 2310 2061 2316 2062
rect 2310 2057 2311 2061
rect 2315 2057 2316 2061
rect 2310 2056 2316 2057
rect 2470 2061 2476 2062
rect 2470 2057 2471 2061
rect 2475 2057 2476 2061
rect 2470 2056 2476 2057
rect 2630 2061 2636 2062
rect 2630 2057 2631 2061
rect 2635 2057 2636 2061
rect 2630 2056 2636 2057
rect 2774 2061 2780 2062
rect 2774 2057 2775 2061
rect 2779 2057 2780 2061
rect 2774 2056 2780 2057
rect 2910 2061 2916 2062
rect 2910 2057 2911 2061
rect 2915 2057 2916 2061
rect 2910 2056 2916 2057
rect 3038 2061 3044 2062
rect 3038 2057 3039 2061
rect 3043 2057 3044 2061
rect 3038 2056 3044 2057
rect 3158 2061 3164 2062
rect 3158 2057 3159 2061
rect 3163 2057 3164 2061
rect 3158 2056 3164 2057
rect 3278 2061 3284 2062
rect 3278 2057 3279 2061
rect 3283 2057 3284 2061
rect 3278 2056 3284 2057
rect 3390 2061 3396 2062
rect 3390 2057 3391 2061
rect 3395 2057 3396 2061
rect 3390 2056 3396 2057
rect 3486 2061 3492 2062
rect 3486 2057 3487 2061
rect 3491 2057 3492 2061
rect 3486 2056 3492 2057
rect 423 2051 429 2052
rect 423 2050 424 2051
rect 110 2048 116 2049
rect 381 2048 424 2050
rect 110 2044 111 2048
rect 115 2044 116 2048
rect 423 2047 424 2048
rect 428 2047 429 2051
rect 543 2051 549 2052
rect 543 2050 544 2051
rect 493 2048 544 2050
rect 423 2046 429 2047
rect 543 2047 544 2048
rect 548 2047 549 2051
rect 671 2051 677 2052
rect 671 2050 672 2051
rect 613 2048 672 2050
rect 543 2046 549 2047
rect 671 2047 672 2048
rect 676 2047 677 2051
rect 791 2051 797 2052
rect 791 2050 792 2051
rect 741 2048 792 2050
rect 671 2046 677 2047
rect 791 2047 792 2048
rect 796 2047 797 2051
rect 1031 2051 1037 2052
rect 1031 2050 1032 2051
rect 981 2048 1032 2050
rect 791 2046 797 2047
rect 1031 2047 1032 2048
rect 1036 2047 1037 2051
rect 1126 2051 1132 2052
rect 1126 2050 1127 2051
rect 1101 2048 1127 2050
rect 1031 2046 1037 2047
rect 1126 2047 1127 2048
rect 1131 2047 1132 2051
rect 1126 2046 1132 2047
rect 1135 2051 1141 2052
rect 1135 2047 1136 2051
rect 1140 2050 1141 2051
rect 1226 2051 1232 2052
rect 1140 2048 1185 2050
rect 1140 2047 1141 2048
rect 1135 2046 1141 2047
rect 1226 2047 1227 2051
rect 1231 2050 1232 2051
rect 1346 2051 1352 2052
rect 1231 2048 1305 2050
rect 1231 2047 1232 2048
rect 1226 2046 1232 2047
rect 1346 2047 1347 2051
rect 1351 2050 1352 2051
rect 1351 2048 1433 2050
rect 1822 2048 1828 2049
rect 1351 2047 1352 2048
rect 1346 2046 1352 2047
rect 110 2043 116 2044
rect 1822 2044 1823 2048
rect 1827 2044 1828 2048
rect 1822 2043 1828 2044
rect 1862 2048 1868 2049
rect 3574 2048 3580 2049
rect 1862 2044 1863 2048
rect 1867 2044 1868 2048
rect 2063 2047 2069 2048
rect 2063 2046 2064 2047
rect 2037 2044 2064 2046
rect 1862 2043 1868 2044
rect 2063 2043 2064 2044
rect 2068 2043 2069 2047
rect 2839 2047 2845 2048
rect 2839 2046 2840 2047
rect 2829 2044 2840 2046
rect 2063 2042 2069 2043
rect 2302 2043 2308 2044
rect 2302 2039 2303 2043
rect 2307 2042 2308 2043
rect 2391 2043 2397 2044
rect 2307 2040 2329 2042
rect 2307 2039 2308 2040
rect 2302 2038 2308 2039
rect 2391 2039 2392 2043
rect 2396 2042 2397 2043
rect 2551 2043 2557 2044
rect 2396 2040 2489 2042
rect 2396 2039 2397 2040
rect 2391 2038 2397 2039
rect 2551 2039 2552 2043
rect 2556 2042 2557 2043
rect 2839 2043 2840 2044
rect 2844 2043 2845 2047
rect 3103 2047 3109 2048
rect 3103 2046 3104 2047
rect 3093 2044 3104 2046
rect 2839 2042 2845 2043
rect 3103 2043 3104 2044
rect 3108 2043 3109 2047
rect 3223 2047 3229 2048
rect 3223 2046 3224 2047
rect 3213 2044 3224 2046
rect 3103 2042 3109 2043
rect 3223 2043 3224 2044
rect 3228 2043 3229 2047
rect 3574 2044 3575 2048
rect 3579 2044 3580 2048
rect 3223 2042 3229 2043
rect 3231 2043 3237 2044
rect 2556 2040 2649 2042
rect 2556 2039 2557 2040
rect 2551 2038 2557 2039
rect 3231 2039 3232 2043
rect 3236 2042 3237 2043
rect 3346 2043 3352 2044
rect 3236 2040 3297 2042
rect 3236 2039 3237 2040
rect 3231 2038 3237 2039
rect 3346 2039 3347 2043
rect 3351 2042 3352 2043
rect 3458 2043 3464 2044
rect 3574 2043 3580 2044
rect 3351 2040 3409 2042
rect 3351 2039 3352 2040
rect 3346 2038 3352 2039
rect 3458 2039 3459 2043
rect 3463 2042 3464 2043
rect 3463 2040 3505 2042
rect 3463 2039 3464 2040
rect 3458 2038 3464 2039
rect 326 2035 332 2036
rect 326 2031 327 2035
rect 331 2031 332 2035
rect 326 2030 332 2031
rect 438 2035 444 2036
rect 438 2031 439 2035
rect 443 2031 444 2035
rect 438 2030 444 2031
rect 558 2035 564 2036
rect 558 2031 559 2035
rect 563 2031 564 2035
rect 558 2030 564 2031
rect 686 2035 692 2036
rect 686 2031 687 2035
rect 691 2031 692 2035
rect 686 2030 692 2031
rect 806 2035 812 2036
rect 806 2031 807 2035
rect 811 2031 812 2035
rect 806 2030 812 2031
rect 926 2035 932 2036
rect 926 2031 927 2035
rect 931 2031 932 2035
rect 926 2030 932 2031
rect 1046 2035 1052 2036
rect 1046 2031 1047 2035
rect 1051 2031 1052 2035
rect 1046 2030 1052 2031
rect 1166 2035 1172 2036
rect 1166 2031 1167 2035
rect 1171 2031 1172 2035
rect 1166 2030 1172 2031
rect 1286 2035 1292 2036
rect 1286 2031 1287 2035
rect 1291 2031 1292 2035
rect 1286 2030 1292 2031
rect 1414 2035 1420 2036
rect 1414 2031 1415 2035
rect 1419 2031 1420 2035
rect 1414 2030 1420 2031
rect 1862 2031 1868 2032
rect 1862 2027 1863 2031
rect 1867 2027 1868 2031
rect 3023 2031 3029 2032
rect 3023 2030 3024 2031
rect 2961 2028 3024 2030
rect 1862 2026 1868 2027
rect 3023 2027 3024 2028
rect 3028 2027 3029 2031
rect 3023 2026 3029 2027
rect 3574 2031 3580 2032
rect 3574 2027 3575 2031
rect 3579 2027 3580 2031
rect 3574 2026 3580 2027
rect 319 2023 325 2024
rect 319 2019 320 2023
rect 324 2022 325 2023
rect 423 2023 429 2024
rect 324 2020 418 2022
rect 324 2019 325 2020
rect 319 2018 325 2019
rect 416 2014 418 2020
rect 423 2019 424 2023
rect 428 2022 429 2023
rect 431 2023 437 2024
rect 431 2022 432 2023
rect 428 2020 432 2022
rect 428 2019 429 2020
rect 423 2018 429 2019
rect 431 2019 432 2020
rect 436 2019 437 2023
rect 431 2018 437 2019
rect 543 2023 549 2024
rect 543 2019 544 2023
rect 548 2022 549 2023
rect 551 2023 557 2024
rect 551 2022 552 2023
rect 548 2020 552 2022
rect 548 2019 549 2020
rect 543 2018 549 2019
rect 551 2019 552 2020
rect 556 2019 557 2023
rect 551 2018 557 2019
rect 671 2023 677 2024
rect 671 2019 672 2023
rect 676 2022 677 2023
rect 679 2023 685 2024
rect 679 2022 680 2023
rect 676 2020 680 2022
rect 676 2019 677 2020
rect 671 2018 677 2019
rect 679 2019 680 2020
rect 684 2019 685 2023
rect 679 2018 685 2019
rect 791 2023 797 2024
rect 791 2019 792 2023
rect 796 2022 797 2023
rect 799 2023 805 2024
rect 799 2022 800 2023
rect 796 2020 800 2022
rect 796 2019 797 2020
rect 791 2018 797 2019
rect 799 2019 800 2020
rect 804 2019 805 2023
rect 799 2018 805 2019
rect 919 2023 925 2024
rect 919 2019 920 2023
rect 924 2022 925 2023
rect 1031 2023 1037 2024
rect 924 2020 1026 2022
rect 924 2019 925 2020
rect 919 2018 925 2019
rect 607 2015 613 2016
rect 607 2014 608 2015
rect 416 2012 608 2014
rect 607 2011 608 2012
rect 612 2011 613 2015
rect 1024 2014 1026 2020
rect 1031 2019 1032 2023
rect 1036 2022 1037 2023
rect 1039 2023 1045 2024
rect 1039 2022 1040 2023
rect 1036 2020 1040 2022
rect 1036 2019 1037 2020
rect 1031 2018 1037 2019
rect 1039 2019 1040 2020
rect 1044 2019 1045 2023
rect 1039 2018 1045 2019
rect 1159 2023 1165 2024
rect 1159 2019 1160 2023
rect 1164 2022 1165 2023
rect 1226 2023 1232 2024
rect 1226 2022 1227 2023
rect 1164 2020 1227 2022
rect 1164 2019 1165 2020
rect 1159 2018 1165 2019
rect 1226 2019 1227 2020
rect 1231 2019 1232 2023
rect 1226 2018 1232 2019
rect 1279 2023 1285 2024
rect 1279 2019 1280 2023
rect 1284 2022 1285 2023
rect 1346 2023 1352 2024
rect 1346 2022 1347 2023
rect 1284 2020 1347 2022
rect 1284 2019 1285 2020
rect 1279 2018 1285 2019
rect 1346 2019 1347 2020
rect 1351 2019 1352 2023
rect 1346 2018 1352 2019
rect 1398 2023 1404 2024
rect 1398 2019 1399 2023
rect 1403 2022 1404 2023
rect 1407 2023 1413 2024
rect 1407 2022 1408 2023
rect 1403 2020 1408 2022
rect 1403 2019 1404 2020
rect 1398 2018 1404 2019
rect 1407 2019 1408 2020
rect 1412 2019 1413 2023
rect 1407 2018 1413 2019
rect 1974 2021 1980 2022
rect 1974 2017 1975 2021
rect 1979 2017 1980 2021
rect 1974 2016 1980 2017
rect 2134 2021 2140 2022
rect 2134 2017 2135 2021
rect 2139 2017 2140 2021
rect 2134 2016 2140 2017
rect 2302 2021 2308 2022
rect 2302 2017 2303 2021
rect 2307 2017 2308 2021
rect 2302 2016 2308 2017
rect 2462 2021 2468 2022
rect 2462 2017 2463 2021
rect 2467 2017 2468 2021
rect 2462 2016 2468 2017
rect 2622 2021 2628 2022
rect 2622 2017 2623 2021
rect 2627 2017 2628 2021
rect 2622 2016 2628 2017
rect 2766 2021 2772 2022
rect 2766 2017 2767 2021
rect 2771 2017 2772 2021
rect 2766 2016 2772 2017
rect 2902 2021 2908 2022
rect 2902 2017 2903 2021
rect 2907 2017 2908 2021
rect 2902 2016 2908 2017
rect 3030 2021 3036 2022
rect 3030 2017 3031 2021
rect 3035 2017 3036 2021
rect 3030 2016 3036 2017
rect 3150 2021 3156 2022
rect 3150 2017 3151 2021
rect 3155 2017 3156 2021
rect 3150 2016 3156 2017
rect 3270 2021 3276 2022
rect 3270 2017 3271 2021
rect 3275 2017 3276 2021
rect 3270 2016 3276 2017
rect 3382 2021 3388 2022
rect 3382 2017 3383 2021
rect 3387 2017 3388 2021
rect 3382 2016 3388 2017
rect 3478 2021 3484 2022
rect 3478 2017 3479 2021
rect 3483 2017 3484 2021
rect 3478 2016 3484 2017
rect 1135 2015 1141 2016
rect 1135 2014 1136 2015
rect 1024 2012 1136 2014
rect 607 2010 613 2011
rect 1135 2011 1136 2012
rect 1140 2011 1141 2015
rect 1135 2010 1141 2011
rect 2183 2015 2189 2016
rect 2183 2011 2184 2015
rect 2188 2014 2189 2015
rect 2191 2015 2197 2016
rect 2191 2014 2192 2015
rect 2188 2012 2192 2014
rect 2188 2011 2189 2012
rect 2183 2010 2189 2011
rect 2191 2011 2192 2012
rect 2196 2011 2197 2015
rect 2191 2010 2197 2011
rect 175 2007 181 2008
rect 175 2003 176 2007
rect 180 2006 181 2007
rect 238 2007 244 2008
rect 238 2006 239 2007
rect 180 2004 239 2006
rect 180 2003 181 2004
rect 175 2002 181 2003
rect 238 2003 239 2004
rect 243 2003 244 2007
rect 238 2002 244 2003
rect 247 2007 253 2008
rect 247 2003 248 2007
rect 252 2006 253 2007
rect 287 2007 293 2008
rect 287 2006 288 2007
rect 252 2004 288 2006
rect 252 2003 253 2004
rect 247 2002 253 2003
rect 287 2003 288 2004
rect 292 2003 293 2007
rect 287 2002 293 2003
rect 359 2007 365 2008
rect 359 2003 360 2007
rect 364 2006 365 2007
rect 407 2007 413 2008
rect 407 2006 408 2007
rect 364 2004 408 2006
rect 364 2003 365 2004
rect 359 2002 365 2003
rect 407 2003 408 2004
rect 412 2003 413 2007
rect 407 2002 413 2003
rect 479 2007 485 2008
rect 479 2003 480 2007
rect 484 2006 485 2007
rect 527 2007 533 2008
rect 527 2006 528 2007
rect 484 2004 528 2006
rect 484 2003 485 2004
rect 479 2002 485 2003
rect 527 2003 528 2004
rect 532 2003 533 2007
rect 527 2002 533 2003
rect 599 2007 605 2008
rect 599 2003 600 2007
rect 604 2006 605 2007
rect 647 2007 653 2008
rect 647 2006 648 2007
rect 604 2004 648 2006
rect 604 2003 605 2004
rect 599 2002 605 2003
rect 647 2003 648 2004
rect 652 2003 653 2007
rect 647 2002 653 2003
rect 767 2007 773 2008
rect 767 2003 768 2007
rect 772 2006 773 2007
rect 842 2007 848 2008
rect 842 2006 843 2007
rect 772 2004 843 2006
rect 772 2003 773 2004
rect 767 2002 773 2003
rect 842 2003 843 2004
rect 847 2003 848 2007
rect 842 2002 848 2003
rect 887 2007 893 2008
rect 887 2003 888 2007
rect 892 2006 893 2007
rect 962 2007 968 2008
rect 962 2006 963 2007
rect 892 2004 963 2006
rect 892 2003 893 2004
rect 887 2002 893 2003
rect 962 2003 963 2004
rect 967 2003 968 2007
rect 962 2002 968 2003
rect 1007 2007 1013 2008
rect 1007 2003 1008 2007
rect 1012 2006 1013 2007
rect 1118 2007 1124 2008
rect 1118 2006 1119 2007
rect 1012 2004 1119 2006
rect 1012 2003 1013 2004
rect 1007 2002 1013 2003
rect 1118 2003 1119 2004
rect 1123 2003 1124 2007
rect 1118 2002 1124 2003
rect 1126 2007 1133 2008
rect 1126 2003 1127 2007
rect 1132 2003 1133 2007
rect 1126 2002 1133 2003
rect 1199 2007 1205 2008
rect 1199 2003 1200 2007
rect 1204 2006 1205 2007
rect 1247 2007 1253 2008
rect 1247 2006 1248 2007
rect 1204 2004 1248 2006
rect 1204 2003 1205 2004
rect 1199 2002 1205 2003
rect 1247 2003 1248 2004
rect 1252 2003 1253 2007
rect 1247 2002 1253 2003
rect 1886 1999 1892 2000
rect 182 1997 188 1998
rect 182 1993 183 1997
rect 187 1993 188 1997
rect 182 1992 188 1993
rect 294 1997 300 1998
rect 294 1993 295 1997
rect 299 1993 300 1997
rect 294 1992 300 1993
rect 414 1997 420 1998
rect 414 1993 415 1997
rect 419 1993 420 1997
rect 414 1992 420 1993
rect 534 1997 540 1998
rect 534 1993 535 1997
rect 539 1993 540 1997
rect 534 1992 540 1993
rect 654 1997 660 1998
rect 654 1993 655 1997
rect 659 1993 660 1997
rect 654 1992 660 1993
rect 774 1997 780 1998
rect 774 1993 775 1997
rect 779 1993 780 1997
rect 774 1992 780 1993
rect 894 1997 900 1998
rect 894 1993 895 1997
rect 899 1993 900 1997
rect 894 1992 900 1993
rect 1014 1997 1020 1998
rect 1014 1993 1015 1997
rect 1019 1993 1020 1997
rect 1014 1992 1020 1993
rect 1134 1997 1140 1998
rect 1134 1993 1135 1997
rect 1139 1993 1140 1997
rect 1134 1992 1140 1993
rect 1254 1997 1260 1998
rect 1254 1993 1255 1997
rect 1259 1993 1260 1997
rect 1886 1995 1887 1999
rect 1891 1995 1892 1999
rect 1886 1994 1892 1995
rect 2030 1999 2036 2000
rect 2030 1995 2031 1999
rect 2035 1995 2036 1999
rect 2030 1994 2036 1995
rect 2198 1999 2204 2000
rect 2198 1995 2199 1999
rect 2203 1995 2204 1999
rect 2198 1994 2204 1995
rect 2374 1999 2380 2000
rect 2374 1995 2375 1999
rect 2379 1995 2380 1999
rect 2374 1994 2380 1995
rect 2542 1999 2548 2000
rect 2542 1995 2543 1999
rect 2547 1995 2548 1999
rect 2542 1994 2548 1995
rect 2710 1999 2716 2000
rect 2710 1995 2711 1999
rect 2715 1995 2716 1999
rect 2710 1994 2716 1995
rect 2870 1999 2876 2000
rect 2870 1995 2871 1999
rect 2875 1995 2876 1999
rect 2870 1994 2876 1995
rect 3038 1999 3044 2000
rect 3038 1995 3039 1999
rect 3043 1995 3044 1999
rect 3038 1994 3044 1995
rect 3206 1999 3212 2000
rect 3206 1995 3207 1999
rect 3211 1995 3212 1999
rect 3206 1994 3212 1995
rect 1254 1992 1260 1993
rect 2610 1991 2616 1992
rect 2610 1990 2611 1991
rect 1862 1989 1868 1990
rect 1862 1985 1863 1989
rect 1867 1985 1868 1989
rect 2601 1988 2611 1990
rect 2610 1987 2611 1988
rect 2615 1987 2616 1991
rect 2610 1986 2616 1987
rect 3574 1989 3580 1990
rect 110 1984 116 1985
rect 1822 1984 1828 1985
rect 1862 1984 1868 1985
rect 3574 1985 3575 1989
rect 3579 1985 3580 1989
rect 3574 1984 3580 1985
rect 110 1980 111 1984
rect 115 1980 116 1984
rect 247 1983 253 1984
rect 247 1982 248 1983
rect 237 1980 248 1982
rect 110 1979 116 1980
rect 247 1979 248 1980
rect 252 1979 253 1983
rect 359 1983 365 1984
rect 359 1982 360 1983
rect 349 1980 360 1982
rect 247 1978 253 1979
rect 359 1979 360 1980
rect 364 1979 365 1983
rect 479 1983 485 1984
rect 479 1982 480 1983
rect 469 1980 480 1982
rect 359 1978 365 1979
rect 479 1979 480 1980
rect 484 1979 485 1983
rect 599 1983 605 1984
rect 599 1982 600 1983
rect 589 1980 600 1982
rect 479 1978 485 1979
rect 599 1979 600 1980
rect 604 1979 605 1983
rect 1199 1983 1205 1984
rect 1199 1982 1200 1983
rect 1189 1980 1200 1982
rect 599 1978 605 1979
rect 607 1979 613 1980
rect 607 1975 608 1979
rect 612 1978 613 1979
rect 842 1979 848 1980
rect 612 1976 673 1978
rect 612 1975 613 1976
rect 607 1974 613 1975
rect 842 1975 843 1979
rect 847 1978 848 1979
rect 962 1979 968 1980
rect 847 1976 913 1978
rect 847 1975 848 1976
rect 842 1974 848 1975
rect 962 1975 963 1979
rect 967 1978 968 1979
rect 1199 1979 1200 1980
rect 1204 1979 1205 1983
rect 1822 1980 1823 1984
rect 1827 1980 1828 1984
rect 1822 1979 1828 1980
rect 1199 1978 1205 1979
rect 967 1976 1033 1978
rect 967 1975 968 1976
rect 962 1974 968 1975
rect 1982 1975 1988 1976
rect 1982 1974 1983 1975
rect 1862 1972 1868 1973
rect 1949 1972 1983 1974
rect 1862 1968 1863 1972
rect 1867 1968 1868 1972
rect 1982 1971 1983 1972
rect 1987 1971 1988 1975
rect 1982 1970 1988 1971
rect 1990 1975 1996 1976
rect 1990 1971 1991 1975
rect 1995 1974 1996 1975
rect 2098 1975 2104 1976
rect 1995 1972 2057 1974
rect 1995 1971 1996 1972
rect 1990 1970 1996 1971
rect 2098 1971 2099 1975
rect 2103 1974 2104 1975
rect 2535 1975 2541 1976
rect 2535 1974 2536 1975
rect 2103 1972 2225 1974
rect 2437 1972 2536 1974
rect 2103 1971 2104 1972
rect 2098 1970 2104 1971
rect 2535 1971 2536 1972
rect 2540 1971 2541 1975
rect 2863 1975 2869 1976
rect 2863 1974 2864 1975
rect 2773 1972 2864 1974
rect 2535 1970 2541 1971
rect 2863 1971 2864 1972
rect 2868 1971 2869 1975
rect 2998 1975 3004 1976
rect 2998 1974 2999 1975
rect 2933 1972 2999 1974
rect 2863 1970 2869 1971
rect 2998 1971 2999 1972
rect 3003 1971 3004 1975
rect 3150 1975 3156 1976
rect 3150 1974 3151 1975
rect 3101 1972 3151 1974
rect 2998 1970 3004 1971
rect 3150 1971 3151 1972
rect 3155 1971 3156 1975
rect 3150 1970 3156 1971
rect 3158 1975 3164 1976
rect 3158 1971 3159 1975
rect 3163 1974 3164 1975
rect 3163 1972 3233 1974
rect 3574 1972 3580 1973
rect 3163 1971 3164 1972
rect 3158 1970 3164 1971
rect 110 1967 116 1968
rect 110 1963 111 1967
rect 115 1963 116 1967
rect 1822 1967 1828 1968
rect 1862 1967 1868 1968
rect 3574 1968 3575 1972
rect 3579 1968 3580 1972
rect 3574 1967 3580 1968
rect 110 1962 116 1963
rect 1196 1964 1265 1966
rect 174 1957 180 1958
rect 174 1953 175 1957
rect 179 1953 180 1957
rect 174 1952 180 1953
rect 286 1957 292 1958
rect 286 1953 287 1957
rect 291 1953 292 1957
rect 286 1952 292 1953
rect 406 1957 412 1958
rect 406 1953 407 1957
rect 411 1953 412 1957
rect 406 1952 412 1953
rect 526 1957 532 1958
rect 526 1953 527 1957
rect 531 1953 532 1957
rect 526 1952 532 1953
rect 646 1957 652 1958
rect 646 1953 647 1957
rect 651 1953 652 1957
rect 646 1952 652 1953
rect 766 1957 772 1958
rect 766 1953 767 1957
rect 771 1953 772 1957
rect 766 1952 772 1953
rect 886 1957 892 1958
rect 886 1953 887 1957
rect 891 1953 892 1957
rect 886 1952 892 1953
rect 1006 1957 1012 1958
rect 1006 1953 1007 1957
rect 1011 1953 1012 1957
rect 1006 1952 1012 1953
rect 1126 1957 1132 1958
rect 1126 1953 1127 1957
rect 1131 1953 1132 1957
rect 1126 1952 1132 1953
rect 815 1951 821 1952
rect 815 1947 816 1951
rect 820 1950 821 1951
rect 831 1951 837 1952
rect 831 1950 832 1951
rect 820 1948 832 1950
rect 820 1947 821 1948
rect 815 1946 821 1947
rect 831 1947 832 1948
rect 836 1947 837 1951
rect 831 1946 837 1947
rect 1118 1951 1124 1952
rect 1118 1947 1119 1951
rect 1123 1950 1124 1951
rect 1196 1950 1198 1964
rect 1822 1963 1823 1967
rect 1827 1963 1828 1967
rect 1822 1962 1828 1963
rect 1894 1959 1900 1960
rect 1246 1957 1252 1958
rect 1246 1953 1247 1957
rect 1251 1953 1252 1957
rect 1894 1955 1895 1959
rect 1899 1955 1900 1959
rect 1894 1954 1900 1955
rect 2038 1959 2044 1960
rect 2038 1955 2039 1959
rect 2043 1955 2044 1959
rect 2038 1954 2044 1955
rect 2206 1959 2212 1960
rect 2206 1955 2207 1959
rect 2211 1955 2212 1959
rect 2206 1954 2212 1955
rect 2382 1959 2388 1960
rect 2382 1955 2383 1959
rect 2387 1955 2388 1959
rect 2382 1954 2388 1955
rect 2550 1959 2556 1960
rect 2550 1955 2551 1959
rect 2555 1955 2556 1959
rect 2550 1954 2556 1955
rect 2718 1959 2724 1960
rect 2718 1955 2719 1959
rect 2723 1955 2724 1959
rect 2718 1954 2724 1955
rect 2878 1959 2884 1960
rect 2878 1955 2879 1959
rect 2883 1955 2884 1959
rect 2878 1954 2884 1955
rect 3046 1959 3052 1960
rect 3046 1955 3047 1959
rect 3051 1955 3052 1959
rect 3046 1954 3052 1955
rect 3214 1959 3220 1960
rect 3214 1955 3215 1959
rect 3219 1955 3220 1959
rect 3214 1954 3220 1955
rect 1246 1952 1252 1953
rect 1123 1948 1198 1950
rect 1123 1947 1124 1948
rect 1118 1946 1124 1947
rect 1887 1947 1893 1948
rect 1887 1943 1888 1947
rect 1892 1946 1893 1947
rect 1990 1947 1996 1948
rect 1990 1946 1991 1947
rect 1892 1944 1991 1946
rect 1892 1943 1893 1944
rect 1887 1942 1893 1943
rect 1990 1943 1991 1944
rect 1995 1943 1996 1947
rect 1990 1942 1996 1943
rect 2031 1947 2037 1948
rect 2031 1943 2032 1947
rect 2036 1946 2037 1947
rect 2098 1947 2104 1948
rect 2098 1946 2099 1947
rect 2036 1944 2099 1946
rect 2036 1943 2037 1944
rect 2031 1942 2037 1943
rect 2098 1943 2099 1944
rect 2103 1943 2104 1947
rect 2098 1942 2104 1943
rect 2191 1947 2197 1948
rect 2191 1943 2192 1947
rect 2196 1946 2197 1947
rect 2199 1947 2205 1948
rect 2199 1946 2200 1947
rect 2196 1944 2200 1946
rect 2196 1943 2197 1944
rect 2191 1942 2197 1943
rect 2199 1943 2200 1944
rect 2204 1943 2205 1947
rect 2199 1942 2205 1943
rect 2338 1947 2344 1948
rect 2338 1943 2339 1947
rect 2343 1946 2344 1947
rect 2375 1947 2381 1948
rect 2375 1946 2376 1947
rect 2343 1944 2376 1946
rect 2343 1943 2344 1944
rect 2338 1942 2344 1943
rect 2375 1943 2376 1944
rect 2380 1943 2381 1947
rect 2375 1942 2381 1943
rect 2535 1947 2541 1948
rect 2535 1943 2536 1947
rect 2540 1946 2541 1947
rect 2543 1947 2549 1948
rect 2543 1946 2544 1947
rect 2540 1944 2544 1946
rect 2540 1943 2541 1944
rect 2535 1942 2541 1943
rect 2543 1943 2544 1944
rect 2548 1943 2549 1947
rect 2543 1942 2549 1943
rect 2711 1947 2717 1948
rect 2711 1943 2712 1947
rect 2716 1946 2717 1947
rect 2726 1947 2732 1948
rect 2726 1946 2727 1947
rect 2716 1944 2727 1946
rect 2716 1943 2717 1944
rect 2711 1942 2717 1943
rect 2726 1943 2727 1944
rect 2731 1943 2732 1947
rect 2726 1942 2732 1943
rect 2863 1947 2869 1948
rect 2863 1943 2864 1947
rect 2868 1946 2869 1947
rect 2871 1947 2877 1948
rect 2871 1946 2872 1947
rect 2868 1944 2872 1946
rect 2868 1943 2869 1944
rect 2863 1942 2869 1943
rect 2871 1943 2872 1944
rect 2876 1943 2877 1947
rect 2871 1942 2877 1943
rect 3023 1947 3029 1948
rect 3023 1943 3024 1947
rect 3028 1946 3029 1947
rect 3039 1947 3045 1948
rect 3039 1946 3040 1947
rect 3028 1944 3040 1946
rect 3028 1943 3029 1944
rect 3023 1942 3029 1943
rect 3039 1943 3040 1944
rect 3044 1943 3045 1947
rect 3039 1942 3045 1943
rect 3150 1947 3156 1948
rect 3150 1943 3151 1947
rect 3155 1946 3156 1947
rect 3207 1947 3213 1948
rect 3207 1946 3208 1947
rect 3155 1944 3208 1946
rect 3155 1943 3156 1944
rect 3150 1942 3156 1943
rect 3207 1943 3208 1944
rect 3212 1943 3213 1947
rect 3207 1942 3213 1943
rect 2063 1935 2069 1936
rect 2063 1934 2064 1935
rect 1889 1932 2064 1934
rect 134 1931 140 1932
rect 134 1927 135 1931
rect 139 1927 140 1931
rect 134 1926 140 1927
rect 222 1931 228 1932
rect 222 1927 223 1931
rect 227 1927 228 1931
rect 222 1926 228 1927
rect 350 1931 356 1932
rect 350 1927 351 1931
rect 355 1927 356 1931
rect 350 1926 356 1927
rect 494 1931 500 1932
rect 494 1927 495 1931
rect 499 1927 500 1931
rect 494 1926 500 1927
rect 654 1931 660 1932
rect 654 1927 655 1931
rect 659 1927 660 1931
rect 654 1926 660 1927
rect 838 1931 844 1932
rect 838 1927 839 1931
rect 843 1927 844 1931
rect 838 1926 844 1927
rect 1038 1931 1044 1932
rect 1038 1927 1039 1931
rect 1043 1927 1044 1931
rect 1038 1926 1044 1927
rect 1246 1931 1252 1932
rect 1246 1927 1247 1931
rect 1251 1927 1252 1931
rect 1246 1926 1252 1927
rect 1462 1931 1468 1932
rect 1462 1927 1463 1931
rect 1467 1927 1468 1931
rect 1889 1928 1891 1932
rect 2063 1931 2064 1932
rect 2068 1931 2069 1935
rect 2063 1930 2069 1931
rect 1462 1926 1468 1927
rect 1887 1927 1893 1928
rect 562 1923 568 1924
rect 110 1921 116 1922
rect 110 1917 111 1921
rect 115 1917 116 1921
rect 562 1919 563 1923
rect 567 1922 568 1923
rect 1158 1923 1164 1924
rect 567 1920 673 1922
rect 567 1919 568 1920
rect 562 1918 568 1919
rect 1158 1919 1159 1923
rect 1163 1922 1164 1923
rect 1887 1923 1888 1927
rect 1892 1923 1893 1927
rect 1887 1922 1893 1923
rect 1982 1927 1989 1928
rect 1982 1923 1983 1927
rect 1988 1923 1989 1927
rect 1982 1922 1989 1923
rect 2055 1927 2061 1928
rect 2055 1923 2056 1927
rect 2060 1926 2061 1927
rect 2111 1927 2117 1928
rect 2111 1926 2112 1927
rect 2060 1924 2112 1926
rect 2060 1923 2061 1924
rect 2055 1922 2061 1923
rect 2111 1923 2112 1924
rect 2116 1923 2117 1927
rect 2111 1922 2117 1923
rect 2247 1927 2253 1928
rect 2247 1923 2248 1927
rect 2252 1926 2253 1927
rect 2346 1927 2352 1928
rect 2346 1926 2347 1927
rect 2252 1924 2347 1926
rect 2252 1923 2253 1924
rect 2247 1922 2253 1923
rect 2346 1923 2347 1924
rect 2351 1923 2352 1927
rect 2346 1922 2352 1923
rect 2366 1927 2372 1928
rect 2366 1923 2367 1927
rect 2371 1926 2372 1927
rect 2375 1927 2381 1928
rect 2375 1926 2376 1927
rect 2371 1924 2376 1926
rect 2371 1923 2372 1924
rect 2366 1922 2372 1923
rect 2375 1923 2376 1924
rect 2380 1923 2381 1927
rect 2375 1922 2381 1923
rect 2503 1927 2509 1928
rect 2503 1923 2504 1927
rect 2508 1926 2509 1927
rect 2578 1927 2584 1928
rect 2578 1926 2579 1927
rect 2508 1924 2579 1926
rect 2508 1923 2509 1924
rect 2503 1922 2509 1923
rect 2578 1923 2579 1924
rect 2583 1923 2584 1927
rect 2578 1922 2584 1923
rect 2623 1927 2629 1928
rect 2623 1923 2624 1927
rect 2628 1926 2629 1927
rect 2698 1927 2704 1928
rect 2698 1926 2699 1927
rect 2628 1924 2699 1926
rect 2628 1923 2629 1924
rect 2623 1922 2629 1923
rect 2698 1923 2699 1924
rect 2703 1923 2704 1927
rect 2698 1922 2704 1923
rect 2743 1927 2749 1928
rect 2743 1923 2744 1927
rect 2748 1926 2749 1927
rect 2818 1927 2824 1928
rect 2818 1926 2819 1927
rect 2748 1924 2819 1926
rect 2748 1923 2749 1924
rect 2743 1922 2749 1923
rect 2818 1923 2819 1924
rect 2823 1923 2824 1927
rect 2818 1922 2824 1923
rect 2871 1927 2877 1928
rect 2871 1923 2872 1927
rect 2876 1926 2877 1927
rect 2946 1927 2952 1928
rect 2946 1926 2947 1927
rect 2876 1924 2947 1926
rect 2876 1923 2877 1924
rect 2871 1922 2877 1923
rect 2946 1923 2947 1924
rect 2951 1923 2952 1927
rect 2946 1922 2952 1923
rect 2998 1927 3005 1928
rect 2998 1923 2999 1927
rect 3004 1923 3005 1927
rect 2998 1922 3005 1923
rect 1163 1920 1265 1922
rect 1822 1921 1828 1922
rect 1163 1919 1164 1920
rect 1158 1918 1164 1919
rect 110 1916 116 1917
rect 1822 1917 1823 1921
rect 1827 1917 1828 1921
rect 1822 1916 1828 1917
rect 1894 1917 1900 1918
rect 1894 1913 1895 1917
rect 1899 1913 1900 1917
rect 1894 1912 1900 1913
rect 1990 1917 1996 1918
rect 1990 1913 1991 1917
rect 1995 1913 1996 1917
rect 1990 1912 1996 1913
rect 2118 1917 2124 1918
rect 2118 1913 2119 1917
rect 2123 1913 2124 1917
rect 2118 1912 2124 1913
rect 2254 1917 2260 1918
rect 2254 1913 2255 1917
rect 2259 1913 2260 1917
rect 2254 1912 2260 1913
rect 2382 1917 2388 1918
rect 2382 1913 2383 1917
rect 2387 1913 2388 1917
rect 2382 1912 2388 1913
rect 2510 1917 2516 1918
rect 2510 1913 2511 1917
rect 2515 1913 2516 1917
rect 2510 1912 2516 1913
rect 2630 1917 2636 1918
rect 2630 1913 2631 1917
rect 2635 1913 2636 1917
rect 2630 1912 2636 1913
rect 2750 1917 2756 1918
rect 2750 1913 2751 1917
rect 2755 1913 2756 1917
rect 2750 1912 2756 1913
rect 2878 1917 2884 1918
rect 2878 1913 2879 1917
rect 2883 1913 2884 1917
rect 2878 1912 2884 1913
rect 3006 1917 3012 1918
rect 3006 1913 3007 1917
rect 3011 1913 3012 1917
rect 3006 1912 3012 1913
rect 215 1907 221 1908
rect 215 1906 216 1907
rect 110 1904 116 1905
rect 197 1904 216 1906
rect 110 1900 111 1904
rect 115 1900 116 1904
rect 215 1903 216 1904
rect 220 1903 221 1907
rect 343 1907 349 1908
rect 343 1906 344 1907
rect 285 1904 344 1906
rect 215 1902 221 1903
rect 343 1903 344 1904
rect 348 1903 349 1907
rect 487 1907 493 1908
rect 487 1906 488 1907
rect 413 1904 488 1906
rect 343 1902 349 1903
rect 487 1903 488 1904
rect 492 1903 493 1907
rect 647 1907 653 1908
rect 647 1906 648 1907
rect 557 1904 648 1906
rect 487 1902 493 1903
rect 647 1903 648 1904
rect 652 1903 653 1907
rect 1007 1907 1013 1908
rect 1007 1906 1008 1907
rect 901 1904 1008 1906
rect 647 1902 653 1903
rect 1007 1903 1008 1904
rect 1012 1903 1013 1907
rect 1239 1907 1245 1908
rect 1239 1906 1240 1907
rect 1101 1904 1240 1906
rect 1007 1902 1013 1903
rect 1239 1903 1240 1904
rect 1244 1903 1245 1907
rect 1239 1902 1245 1903
rect 1455 1907 1461 1908
rect 1455 1903 1456 1907
rect 1460 1906 1461 1907
rect 1460 1904 1489 1906
rect 1822 1904 1828 1905
rect 1460 1903 1461 1904
rect 1455 1902 1461 1903
rect 110 1899 116 1900
rect 1822 1900 1823 1904
rect 1827 1900 1828 1904
rect 1822 1899 1828 1900
rect 1862 1904 1868 1905
rect 3574 1904 3580 1905
rect 1862 1900 1863 1904
rect 1867 1900 1868 1904
rect 2055 1903 2061 1904
rect 2055 1902 2056 1903
rect 2045 1900 2056 1902
rect 1862 1899 1868 1900
rect 2055 1899 2056 1900
rect 2060 1899 2061 1903
rect 2338 1903 2344 1904
rect 2338 1902 2339 1903
rect 2309 1900 2339 1902
rect 2055 1898 2061 1899
rect 2063 1899 2069 1900
rect 2063 1895 2064 1899
rect 2068 1898 2069 1899
rect 2338 1899 2339 1900
rect 2343 1899 2344 1903
rect 3574 1900 3575 1904
rect 3579 1900 3580 1904
rect 2338 1898 2344 1899
rect 2346 1899 2352 1900
rect 2068 1896 2137 1898
rect 2068 1895 2069 1896
rect 2063 1894 2069 1895
rect 2346 1895 2347 1899
rect 2351 1898 2352 1899
rect 2578 1899 2584 1900
rect 2351 1896 2401 1898
rect 2351 1895 2352 1896
rect 2346 1894 2352 1895
rect 2578 1895 2579 1899
rect 2583 1898 2584 1899
rect 2698 1899 2704 1900
rect 2583 1896 2649 1898
rect 2583 1895 2584 1896
rect 2578 1894 2584 1895
rect 2698 1895 2699 1899
rect 2703 1898 2704 1899
rect 2818 1899 2824 1900
rect 2703 1896 2769 1898
rect 2703 1895 2704 1896
rect 2698 1894 2704 1895
rect 2818 1895 2819 1899
rect 2823 1898 2824 1899
rect 2946 1899 2952 1900
rect 3574 1899 3580 1900
rect 2823 1896 2897 1898
rect 2823 1895 2824 1896
rect 2818 1894 2824 1895
rect 2946 1895 2947 1899
rect 2951 1898 2952 1899
rect 2951 1896 3025 1898
rect 2951 1895 2952 1896
rect 2946 1894 2952 1895
rect 142 1891 148 1892
rect 142 1887 143 1891
rect 147 1887 148 1891
rect 142 1886 148 1887
rect 230 1891 236 1892
rect 230 1887 231 1891
rect 235 1887 236 1891
rect 230 1886 236 1887
rect 358 1891 364 1892
rect 358 1887 359 1891
rect 363 1887 364 1891
rect 358 1886 364 1887
rect 502 1891 508 1892
rect 502 1887 503 1891
rect 507 1887 508 1891
rect 502 1886 508 1887
rect 662 1891 668 1892
rect 662 1887 663 1891
rect 667 1887 668 1891
rect 662 1886 668 1887
rect 846 1891 852 1892
rect 846 1887 847 1891
rect 851 1887 852 1891
rect 846 1886 852 1887
rect 1046 1891 1052 1892
rect 1046 1887 1047 1891
rect 1051 1887 1052 1891
rect 1046 1886 1052 1887
rect 1254 1891 1260 1892
rect 1254 1887 1255 1891
rect 1259 1887 1260 1891
rect 1254 1886 1260 1887
rect 1470 1891 1476 1892
rect 1470 1887 1471 1891
rect 1475 1887 1476 1891
rect 1470 1886 1476 1887
rect 1862 1887 1868 1888
rect 1862 1883 1863 1887
rect 1867 1883 1868 1887
rect 1862 1882 1868 1883
rect 1870 1887 1876 1888
rect 1870 1883 1871 1887
rect 1875 1886 1876 1887
rect 2510 1887 2516 1888
rect 1875 1884 1905 1886
rect 1875 1883 1876 1884
rect 1870 1882 1876 1883
rect 2510 1883 2511 1887
rect 2515 1886 2516 1887
rect 3574 1887 3580 1888
rect 2515 1884 2521 1886
rect 2515 1883 2516 1884
rect 2510 1882 2516 1883
rect 3574 1883 3575 1887
rect 3579 1883 3580 1887
rect 3574 1882 3580 1883
rect 134 1879 141 1880
rect 134 1875 135 1879
rect 140 1875 141 1879
rect 134 1874 141 1875
rect 215 1879 221 1880
rect 215 1875 216 1879
rect 220 1878 221 1879
rect 223 1879 229 1880
rect 223 1878 224 1879
rect 220 1876 224 1878
rect 220 1875 221 1876
rect 215 1874 221 1875
rect 223 1875 224 1876
rect 228 1875 229 1879
rect 223 1874 229 1875
rect 343 1879 349 1880
rect 343 1875 344 1879
rect 348 1878 349 1879
rect 351 1879 357 1880
rect 351 1878 352 1879
rect 348 1876 352 1878
rect 348 1875 349 1876
rect 343 1874 349 1875
rect 351 1875 352 1876
rect 356 1875 357 1879
rect 351 1874 357 1875
rect 487 1879 493 1880
rect 487 1875 488 1879
rect 492 1878 493 1879
rect 495 1879 501 1880
rect 495 1878 496 1879
rect 492 1876 496 1878
rect 492 1875 493 1876
rect 487 1874 493 1875
rect 495 1875 496 1876
rect 500 1875 501 1879
rect 495 1874 501 1875
rect 647 1879 653 1880
rect 647 1875 648 1879
rect 652 1878 653 1879
rect 655 1879 661 1880
rect 655 1878 656 1879
rect 652 1876 656 1878
rect 652 1875 653 1876
rect 647 1874 653 1875
rect 655 1875 656 1876
rect 660 1875 661 1879
rect 655 1874 661 1875
rect 831 1879 837 1880
rect 831 1875 832 1879
rect 836 1878 837 1879
rect 839 1879 845 1880
rect 839 1878 840 1879
rect 836 1876 840 1878
rect 836 1875 837 1876
rect 831 1874 837 1875
rect 839 1875 840 1876
rect 844 1875 845 1879
rect 839 1874 845 1875
rect 1007 1879 1013 1880
rect 1007 1875 1008 1879
rect 1012 1878 1013 1879
rect 1039 1879 1045 1880
rect 1039 1878 1040 1879
rect 1012 1876 1040 1878
rect 1012 1875 1013 1876
rect 1007 1874 1013 1875
rect 1039 1875 1040 1876
rect 1044 1875 1045 1879
rect 1039 1874 1045 1875
rect 1239 1879 1245 1880
rect 1239 1875 1240 1879
rect 1244 1878 1245 1879
rect 1247 1879 1253 1880
rect 1247 1878 1248 1879
rect 1244 1876 1248 1878
rect 1244 1875 1245 1876
rect 1239 1874 1245 1875
rect 1247 1875 1248 1876
rect 1252 1875 1253 1879
rect 1247 1874 1253 1875
rect 1255 1879 1261 1880
rect 1255 1875 1256 1879
rect 1260 1878 1261 1879
rect 1463 1879 1469 1880
rect 1463 1878 1464 1879
rect 1260 1876 1464 1878
rect 1260 1875 1261 1876
rect 1255 1874 1261 1875
rect 1463 1875 1464 1876
rect 1468 1875 1469 1879
rect 1463 1874 1469 1875
rect 1886 1877 1892 1878
rect 1886 1873 1887 1877
rect 1891 1873 1892 1877
rect 1886 1872 1892 1873
rect 1982 1877 1988 1878
rect 1982 1873 1983 1877
rect 1987 1873 1988 1877
rect 1982 1872 1988 1873
rect 2110 1877 2116 1878
rect 2110 1873 2111 1877
rect 2115 1873 2116 1877
rect 2110 1872 2116 1873
rect 2246 1877 2252 1878
rect 2246 1873 2247 1877
rect 2251 1873 2252 1877
rect 2246 1872 2252 1873
rect 2374 1877 2380 1878
rect 2374 1873 2375 1877
rect 2379 1873 2380 1877
rect 2374 1872 2380 1873
rect 2502 1877 2508 1878
rect 2502 1873 2503 1877
rect 2507 1873 2508 1877
rect 2502 1872 2508 1873
rect 2622 1877 2628 1878
rect 2622 1873 2623 1877
rect 2627 1873 2628 1877
rect 2622 1872 2628 1873
rect 2742 1877 2748 1878
rect 2742 1873 2743 1877
rect 2747 1873 2748 1877
rect 2742 1872 2748 1873
rect 2870 1877 2876 1878
rect 2870 1873 2871 1877
rect 2875 1873 2876 1877
rect 2870 1872 2876 1873
rect 2998 1877 3004 1878
rect 2998 1873 2999 1877
rect 3003 1873 3004 1877
rect 2998 1872 3004 1873
rect 1426 1867 1432 1868
rect 1426 1866 1427 1867
rect 1320 1864 1427 1866
rect 135 1859 141 1860
rect 135 1855 136 1859
rect 140 1858 141 1859
rect 210 1859 216 1860
rect 210 1858 211 1859
rect 140 1856 211 1858
rect 140 1855 141 1856
rect 135 1854 141 1855
rect 210 1855 211 1856
rect 215 1855 216 1859
rect 210 1854 216 1855
rect 263 1859 269 1860
rect 263 1855 264 1859
rect 268 1858 269 1859
rect 338 1859 344 1860
rect 338 1858 339 1859
rect 268 1856 339 1858
rect 268 1855 269 1856
rect 263 1854 269 1855
rect 338 1855 339 1856
rect 343 1855 344 1859
rect 338 1854 344 1855
rect 370 1859 376 1860
rect 370 1855 371 1859
rect 375 1858 376 1859
rect 407 1859 413 1860
rect 407 1858 408 1859
rect 375 1856 408 1858
rect 375 1855 376 1856
rect 370 1854 376 1855
rect 407 1855 408 1856
rect 412 1855 413 1859
rect 407 1854 413 1855
rect 551 1859 557 1860
rect 551 1855 552 1859
rect 556 1858 557 1859
rect 647 1859 653 1860
rect 647 1858 648 1859
rect 556 1856 648 1858
rect 556 1855 557 1856
rect 551 1854 557 1855
rect 647 1855 648 1856
rect 652 1855 653 1859
rect 647 1854 653 1855
rect 687 1859 693 1860
rect 687 1855 688 1859
rect 692 1858 693 1859
rect 762 1859 768 1860
rect 762 1858 763 1859
rect 692 1856 763 1858
rect 692 1855 693 1856
rect 687 1854 693 1855
rect 762 1855 763 1856
rect 767 1855 768 1859
rect 762 1854 768 1855
rect 815 1859 821 1860
rect 815 1855 816 1859
rect 820 1858 821 1859
rect 890 1859 896 1860
rect 890 1858 891 1859
rect 820 1856 891 1858
rect 820 1855 821 1856
rect 815 1854 821 1855
rect 890 1855 891 1856
rect 895 1855 896 1859
rect 890 1854 896 1855
rect 935 1859 941 1860
rect 935 1855 936 1859
rect 940 1858 941 1859
rect 950 1859 956 1860
rect 950 1858 951 1859
rect 940 1856 951 1858
rect 940 1855 941 1856
rect 935 1854 941 1855
rect 950 1855 951 1856
rect 955 1855 956 1859
rect 950 1854 956 1855
rect 1047 1859 1053 1860
rect 1047 1855 1048 1859
rect 1052 1858 1053 1859
rect 1110 1859 1116 1860
rect 1110 1858 1111 1859
rect 1052 1856 1111 1858
rect 1052 1855 1053 1856
rect 1047 1854 1053 1855
rect 1110 1855 1111 1856
rect 1115 1855 1116 1859
rect 1110 1854 1116 1855
rect 1119 1859 1125 1860
rect 1119 1855 1120 1859
rect 1124 1858 1125 1859
rect 1151 1859 1157 1860
rect 1151 1858 1152 1859
rect 1124 1856 1152 1858
rect 1124 1855 1125 1856
rect 1119 1854 1125 1855
rect 1151 1855 1152 1856
rect 1156 1855 1157 1859
rect 1151 1854 1157 1855
rect 1255 1859 1261 1860
rect 1255 1855 1256 1859
rect 1260 1858 1261 1859
rect 1320 1858 1322 1864
rect 1426 1863 1427 1864
rect 1431 1863 1432 1867
rect 1426 1862 1432 1863
rect 1260 1856 1322 1858
rect 1327 1859 1333 1860
rect 1260 1855 1261 1856
rect 1255 1854 1261 1855
rect 1327 1855 1328 1859
rect 1332 1858 1333 1859
rect 1351 1859 1357 1860
rect 1351 1858 1352 1859
rect 1332 1856 1352 1858
rect 1332 1855 1333 1856
rect 1327 1854 1333 1855
rect 1351 1855 1352 1856
rect 1356 1855 1357 1859
rect 1351 1854 1357 1855
rect 1447 1859 1453 1860
rect 1447 1855 1448 1859
rect 1452 1858 1453 1859
rect 1455 1859 1461 1860
rect 1455 1858 1456 1859
rect 1452 1856 1456 1858
rect 1452 1855 1453 1856
rect 1447 1854 1453 1855
rect 1455 1855 1456 1856
rect 1460 1855 1461 1859
rect 1455 1854 1461 1855
rect 1543 1859 1549 1860
rect 1543 1855 1544 1859
rect 1548 1858 1549 1859
rect 1618 1859 1624 1860
rect 1618 1858 1619 1859
rect 1548 1856 1619 1858
rect 1548 1855 1549 1856
rect 1543 1854 1549 1855
rect 1618 1855 1619 1856
rect 1623 1855 1624 1859
rect 1618 1854 1624 1855
rect 1639 1859 1645 1860
rect 1639 1855 1640 1859
rect 1644 1858 1645 1859
rect 1714 1859 1720 1860
rect 1714 1858 1715 1859
rect 1644 1856 1715 1858
rect 1644 1855 1645 1856
rect 1639 1854 1645 1855
rect 1714 1855 1715 1856
rect 1719 1855 1720 1859
rect 1714 1854 1720 1855
rect 1727 1859 1733 1860
rect 1727 1855 1728 1859
rect 1732 1858 1733 1859
rect 1870 1859 1876 1860
rect 1870 1858 1871 1859
rect 1732 1856 1871 1858
rect 1732 1855 1733 1856
rect 1727 1854 1733 1855
rect 1870 1855 1871 1856
rect 1875 1855 1876 1859
rect 1870 1854 1876 1855
rect 142 1849 148 1850
rect 142 1845 143 1849
rect 147 1845 148 1849
rect 142 1844 148 1845
rect 270 1849 276 1850
rect 270 1845 271 1849
rect 275 1845 276 1849
rect 270 1844 276 1845
rect 414 1849 420 1850
rect 414 1845 415 1849
rect 419 1845 420 1849
rect 414 1844 420 1845
rect 558 1849 564 1850
rect 558 1845 559 1849
rect 563 1845 564 1849
rect 558 1844 564 1845
rect 694 1849 700 1850
rect 694 1845 695 1849
rect 699 1845 700 1849
rect 694 1844 700 1845
rect 822 1849 828 1850
rect 822 1845 823 1849
rect 827 1845 828 1849
rect 822 1844 828 1845
rect 942 1849 948 1850
rect 942 1845 943 1849
rect 947 1845 948 1849
rect 942 1844 948 1845
rect 1054 1849 1060 1850
rect 1054 1845 1055 1849
rect 1059 1845 1060 1849
rect 1054 1844 1060 1845
rect 1158 1849 1164 1850
rect 1158 1845 1159 1849
rect 1163 1845 1164 1849
rect 1158 1844 1164 1845
rect 1262 1849 1268 1850
rect 1262 1845 1263 1849
rect 1267 1845 1268 1849
rect 1262 1844 1268 1845
rect 1358 1849 1364 1850
rect 1358 1845 1359 1849
rect 1363 1845 1364 1849
rect 1358 1844 1364 1845
rect 1454 1849 1460 1850
rect 1454 1845 1455 1849
rect 1459 1845 1460 1849
rect 1454 1844 1460 1845
rect 1550 1849 1556 1850
rect 1550 1845 1551 1849
rect 1555 1845 1556 1849
rect 1550 1844 1556 1845
rect 1646 1849 1652 1850
rect 1646 1845 1647 1849
rect 1651 1845 1652 1849
rect 1646 1844 1652 1845
rect 1734 1849 1740 1850
rect 1734 1845 1735 1849
rect 1739 1845 1740 1849
rect 1734 1844 1740 1845
rect 2222 1847 2228 1848
rect 2222 1843 2223 1847
rect 2227 1843 2228 1847
rect 2222 1842 2228 1843
rect 2358 1847 2364 1848
rect 2358 1843 2359 1847
rect 2363 1843 2364 1847
rect 2358 1842 2364 1843
rect 2494 1847 2500 1848
rect 2494 1843 2495 1847
rect 2499 1843 2500 1847
rect 2494 1842 2500 1843
rect 2622 1847 2628 1848
rect 2622 1843 2623 1847
rect 2627 1843 2628 1847
rect 2622 1842 2628 1843
rect 2742 1847 2748 1848
rect 2742 1843 2743 1847
rect 2747 1843 2748 1847
rect 2742 1842 2748 1843
rect 2862 1847 2868 1848
rect 2862 1843 2863 1847
rect 2867 1843 2868 1847
rect 2862 1842 2868 1843
rect 2990 1847 2996 1848
rect 2990 1843 2991 1847
rect 2995 1843 2996 1847
rect 2990 1842 2996 1843
rect 2930 1839 2936 1840
rect 1862 1837 1868 1838
rect 110 1836 116 1837
rect 1822 1836 1828 1837
rect 110 1832 111 1836
rect 115 1832 116 1836
rect 1119 1835 1125 1836
rect 1119 1834 1120 1835
rect 1109 1832 1120 1834
rect 110 1831 116 1832
rect 134 1831 140 1832
rect 134 1827 135 1831
rect 139 1830 140 1831
rect 210 1831 216 1832
rect 139 1828 161 1830
rect 139 1827 140 1828
rect 134 1826 140 1827
rect 210 1827 211 1831
rect 215 1830 216 1831
rect 338 1831 344 1832
rect 215 1828 289 1830
rect 215 1827 216 1828
rect 210 1826 216 1827
rect 338 1827 339 1831
rect 343 1830 344 1831
rect 647 1831 653 1832
rect 343 1828 433 1830
rect 343 1827 344 1828
rect 338 1826 344 1827
rect 647 1827 648 1831
rect 652 1830 653 1831
rect 762 1831 768 1832
rect 652 1828 713 1830
rect 652 1827 653 1828
rect 647 1826 653 1827
rect 762 1827 763 1831
rect 767 1830 768 1831
rect 890 1831 896 1832
rect 767 1828 841 1830
rect 767 1827 768 1828
rect 762 1826 768 1827
rect 890 1827 891 1831
rect 895 1830 896 1831
rect 1119 1831 1120 1832
rect 1124 1831 1125 1835
rect 1247 1835 1253 1836
rect 1247 1834 1248 1835
rect 1213 1832 1248 1834
rect 1119 1830 1125 1831
rect 1247 1831 1248 1832
rect 1252 1831 1253 1835
rect 1327 1835 1333 1836
rect 1327 1834 1328 1835
rect 1317 1832 1328 1834
rect 1247 1830 1253 1831
rect 1327 1831 1328 1832
rect 1332 1831 1333 1835
rect 1822 1832 1823 1836
rect 1827 1832 1828 1836
rect 1862 1833 1863 1837
rect 1867 1833 1868 1837
rect 2368 1836 2377 1838
rect 1862 1832 1868 1833
rect 2366 1835 2372 1836
rect 1327 1830 1333 1831
rect 1426 1831 1432 1832
rect 895 1828 961 1830
rect 895 1827 896 1828
rect 890 1826 896 1827
rect 1426 1827 1427 1831
rect 1431 1830 1432 1831
rect 1618 1831 1624 1832
rect 1431 1828 1473 1830
rect 1431 1827 1432 1828
rect 1426 1826 1432 1827
rect 1618 1827 1619 1831
rect 1623 1830 1624 1831
rect 1714 1831 1720 1832
rect 1822 1831 1828 1832
rect 2366 1831 2367 1835
rect 2371 1831 2372 1835
rect 2930 1835 2931 1839
rect 2935 1838 2936 1839
rect 2935 1836 3009 1838
rect 3574 1837 3580 1838
rect 2935 1835 2936 1836
rect 2930 1834 2936 1835
rect 3574 1833 3575 1837
rect 3579 1833 3580 1837
rect 3574 1832 3580 1833
rect 1623 1828 1665 1830
rect 1623 1827 1624 1828
rect 1618 1826 1624 1827
rect 1714 1827 1715 1831
rect 1719 1830 1720 1831
rect 2366 1830 2372 1831
rect 1719 1828 1753 1830
rect 1719 1827 1720 1828
rect 1714 1826 1720 1827
rect 2351 1823 2357 1824
rect 2351 1822 2352 1823
rect 1862 1820 1868 1821
rect 2285 1820 2352 1822
rect 110 1819 116 1820
rect 110 1815 111 1819
rect 115 1815 116 1819
rect 110 1814 116 1815
rect 510 1819 516 1820
rect 510 1815 511 1819
rect 515 1818 516 1819
rect 1550 1819 1556 1820
rect 515 1816 569 1818
rect 515 1815 516 1816
rect 510 1814 516 1815
rect 1550 1815 1551 1819
rect 1555 1818 1556 1819
rect 1822 1819 1828 1820
rect 1555 1816 1561 1818
rect 1555 1815 1556 1816
rect 1550 1814 1556 1815
rect 1822 1815 1823 1819
rect 1827 1815 1828 1819
rect 1862 1816 1863 1820
rect 1867 1816 1868 1820
rect 2351 1819 2352 1820
rect 2356 1819 2357 1823
rect 2615 1823 2621 1824
rect 2615 1822 2616 1823
rect 2557 1820 2616 1822
rect 2351 1818 2357 1819
rect 2615 1819 2616 1820
rect 2620 1819 2621 1823
rect 2735 1823 2741 1824
rect 2735 1822 2736 1823
rect 2685 1820 2736 1822
rect 2615 1818 2621 1819
rect 2735 1819 2736 1820
rect 2740 1819 2741 1823
rect 2855 1823 2861 1824
rect 2855 1822 2856 1823
rect 2805 1820 2856 1822
rect 2735 1818 2741 1819
rect 2855 1819 2856 1820
rect 2860 1819 2861 1823
rect 2983 1823 2989 1824
rect 2983 1822 2984 1823
rect 2925 1820 2984 1822
rect 2855 1818 2861 1819
rect 2983 1819 2984 1820
rect 2988 1819 2989 1823
rect 2983 1818 2989 1819
rect 3574 1820 3580 1821
rect 1862 1815 1868 1816
rect 3574 1816 3575 1820
rect 3579 1816 3580 1820
rect 3574 1815 3580 1816
rect 1822 1814 1828 1815
rect 134 1809 140 1810
rect 134 1805 135 1809
rect 139 1805 140 1809
rect 134 1804 140 1805
rect 262 1809 268 1810
rect 262 1805 263 1809
rect 267 1805 268 1809
rect 262 1804 268 1805
rect 406 1809 412 1810
rect 406 1805 407 1809
rect 411 1805 412 1809
rect 406 1804 412 1805
rect 550 1809 556 1810
rect 550 1805 551 1809
rect 555 1805 556 1809
rect 550 1804 556 1805
rect 686 1809 692 1810
rect 686 1805 687 1809
rect 691 1805 692 1809
rect 686 1804 692 1805
rect 814 1809 820 1810
rect 814 1805 815 1809
rect 819 1805 820 1809
rect 814 1804 820 1805
rect 934 1809 940 1810
rect 934 1805 935 1809
rect 939 1805 940 1809
rect 934 1804 940 1805
rect 1046 1809 1052 1810
rect 1046 1805 1047 1809
rect 1051 1805 1052 1809
rect 1046 1804 1052 1805
rect 1150 1809 1156 1810
rect 1150 1805 1151 1809
rect 1155 1805 1156 1809
rect 1150 1804 1156 1805
rect 1254 1809 1260 1810
rect 1254 1805 1255 1809
rect 1259 1805 1260 1809
rect 1254 1804 1260 1805
rect 1350 1809 1356 1810
rect 1350 1805 1351 1809
rect 1355 1805 1356 1809
rect 1350 1804 1356 1805
rect 1446 1809 1452 1810
rect 1446 1805 1447 1809
rect 1451 1805 1452 1809
rect 1446 1804 1452 1805
rect 1542 1809 1548 1810
rect 1542 1805 1543 1809
rect 1547 1805 1548 1809
rect 1542 1804 1548 1805
rect 1638 1809 1644 1810
rect 1638 1805 1639 1809
rect 1643 1805 1644 1809
rect 1638 1804 1644 1805
rect 1726 1809 1732 1810
rect 1726 1805 1727 1809
rect 1731 1805 1732 1809
rect 1726 1804 1732 1805
rect 2230 1807 2236 1808
rect 1390 1803 1396 1804
rect 1390 1799 1391 1803
rect 1395 1802 1396 1803
rect 1399 1803 1405 1804
rect 1399 1802 1400 1803
rect 1395 1800 1400 1802
rect 1395 1799 1396 1800
rect 1390 1798 1396 1799
rect 1399 1799 1400 1800
rect 1404 1799 1405 1803
rect 2230 1803 2231 1807
rect 2235 1803 2236 1807
rect 2230 1802 2236 1803
rect 2366 1807 2372 1808
rect 2366 1803 2367 1807
rect 2371 1803 2372 1807
rect 2366 1802 2372 1803
rect 2502 1807 2508 1808
rect 2502 1803 2503 1807
rect 2507 1803 2508 1807
rect 2502 1802 2508 1803
rect 2630 1807 2636 1808
rect 2630 1803 2631 1807
rect 2635 1803 2636 1807
rect 2630 1802 2636 1803
rect 2750 1807 2756 1808
rect 2750 1803 2751 1807
rect 2755 1803 2756 1807
rect 2750 1802 2756 1803
rect 2870 1807 2876 1808
rect 2870 1803 2871 1807
rect 2875 1803 2876 1807
rect 2870 1802 2876 1803
rect 2998 1807 3004 1808
rect 2998 1803 2999 1807
rect 3003 1803 3004 1807
rect 2998 1802 3004 1803
rect 1399 1798 1405 1799
rect 2223 1795 2229 1796
rect 2223 1791 2224 1795
rect 2228 1794 2229 1795
rect 2330 1795 2336 1796
rect 2330 1794 2331 1795
rect 2228 1792 2331 1794
rect 2228 1791 2229 1792
rect 2223 1790 2229 1791
rect 2330 1791 2331 1792
rect 2335 1791 2336 1795
rect 2330 1790 2336 1791
rect 2351 1795 2357 1796
rect 2351 1791 2352 1795
rect 2356 1794 2357 1795
rect 2359 1795 2365 1796
rect 2359 1794 2360 1795
rect 2356 1792 2360 1794
rect 2356 1791 2357 1792
rect 2351 1790 2357 1791
rect 2359 1791 2360 1792
rect 2364 1791 2365 1795
rect 2359 1790 2365 1791
rect 2495 1795 2501 1796
rect 2495 1791 2496 1795
rect 2500 1794 2501 1795
rect 2510 1795 2516 1796
rect 2510 1794 2511 1795
rect 2500 1792 2511 1794
rect 2500 1791 2501 1792
rect 2495 1790 2501 1791
rect 2510 1791 2511 1792
rect 2515 1791 2516 1795
rect 2510 1790 2516 1791
rect 2615 1795 2621 1796
rect 2615 1791 2616 1795
rect 2620 1794 2621 1795
rect 2623 1795 2629 1796
rect 2623 1794 2624 1795
rect 2620 1792 2624 1794
rect 2620 1791 2621 1792
rect 2615 1790 2621 1791
rect 2623 1791 2624 1792
rect 2628 1791 2629 1795
rect 2623 1790 2629 1791
rect 2735 1795 2741 1796
rect 2735 1791 2736 1795
rect 2740 1794 2741 1795
rect 2743 1795 2749 1796
rect 2743 1794 2744 1795
rect 2740 1792 2744 1794
rect 2740 1791 2741 1792
rect 2735 1790 2741 1791
rect 2743 1791 2744 1792
rect 2748 1791 2749 1795
rect 2743 1790 2749 1791
rect 2855 1795 2861 1796
rect 2855 1791 2856 1795
rect 2860 1794 2861 1795
rect 2863 1795 2869 1796
rect 2863 1794 2864 1795
rect 2860 1792 2864 1794
rect 2860 1791 2861 1792
rect 2855 1790 2861 1791
rect 2863 1791 2864 1792
rect 2868 1791 2869 1795
rect 2863 1790 2869 1791
rect 2983 1795 2989 1796
rect 2983 1791 2984 1795
rect 2988 1794 2989 1795
rect 2991 1795 2997 1796
rect 2991 1794 2992 1795
rect 2988 1792 2992 1794
rect 2988 1791 2989 1792
rect 2983 1790 2989 1791
rect 2991 1791 2992 1792
rect 2996 1791 2997 1795
rect 2991 1790 2997 1791
rect 2930 1787 2936 1788
rect 2930 1786 2931 1787
rect 2816 1784 2931 1786
rect 2263 1779 2269 1780
rect 134 1775 140 1776
rect 134 1771 135 1775
rect 139 1771 140 1775
rect 134 1770 140 1771
rect 302 1775 308 1776
rect 302 1771 303 1775
rect 307 1771 308 1775
rect 302 1770 308 1771
rect 494 1775 500 1776
rect 494 1771 495 1775
rect 499 1771 500 1775
rect 494 1770 500 1771
rect 686 1775 692 1776
rect 686 1771 687 1775
rect 691 1771 692 1775
rect 686 1770 692 1771
rect 870 1775 876 1776
rect 870 1771 871 1775
rect 875 1771 876 1775
rect 870 1770 876 1771
rect 1046 1775 1052 1776
rect 1046 1771 1047 1775
rect 1051 1771 1052 1775
rect 1046 1770 1052 1771
rect 1214 1775 1220 1776
rect 1214 1771 1215 1775
rect 1219 1771 1220 1775
rect 1214 1770 1220 1771
rect 1374 1775 1380 1776
rect 1374 1771 1375 1775
rect 1379 1771 1380 1775
rect 1374 1770 1380 1771
rect 1534 1775 1540 1776
rect 1534 1771 1535 1775
rect 1539 1771 1540 1775
rect 1534 1770 1540 1771
rect 1702 1775 1708 1776
rect 1702 1771 1703 1775
rect 1707 1771 1708 1775
rect 2263 1775 2264 1779
rect 2268 1778 2269 1779
rect 2338 1779 2344 1780
rect 2338 1778 2339 1779
rect 2268 1776 2339 1778
rect 2268 1775 2269 1776
rect 2263 1774 2269 1775
rect 2338 1775 2339 1776
rect 2343 1775 2344 1779
rect 2338 1774 2344 1775
rect 2351 1779 2357 1780
rect 2351 1775 2352 1779
rect 2356 1778 2357 1779
rect 2426 1779 2432 1780
rect 2426 1778 2427 1779
rect 2356 1776 2427 1778
rect 2356 1775 2357 1776
rect 2351 1774 2357 1775
rect 2426 1775 2427 1776
rect 2431 1775 2432 1779
rect 2426 1774 2432 1775
rect 2447 1779 2453 1780
rect 2447 1775 2448 1779
rect 2452 1778 2453 1779
rect 2522 1779 2528 1780
rect 2522 1778 2523 1779
rect 2452 1776 2523 1778
rect 2452 1775 2453 1776
rect 2447 1774 2453 1775
rect 2522 1775 2523 1776
rect 2527 1775 2528 1779
rect 2522 1774 2528 1775
rect 2551 1779 2557 1780
rect 2551 1775 2552 1779
rect 2556 1778 2557 1779
rect 2631 1779 2637 1780
rect 2631 1778 2632 1779
rect 2556 1776 2632 1778
rect 2556 1775 2557 1776
rect 2551 1774 2557 1775
rect 2631 1775 2632 1776
rect 2636 1775 2637 1779
rect 2631 1774 2637 1775
rect 2655 1779 2661 1780
rect 2655 1775 2656 1779
rect 2660 1778 2661 1779
rect 2722 1779 2728 1780
rect 2722 1778 2723 1779
rect 2660 1776 2723 1778
rect 2660 1775 2661 1776
rect 2655 1774 2661 1775
rect 2722 1775 2723 1776
rect 2727 1775 2728 1779
rect 2722 1774 2728 1775
rect 2751 1779 2757 1780
rect 2751 1775 2752 1779
rect 2756 1778 2757 1779
rect 2816 1778 2818 1784
rect 2930 1783 2931 1784
rect 2935 1783 2936 1787
rect 2930 1782 2936 1783
rect 2756 1776 2818 1778
rect 2823 1779 2829 1780
rect 2756 1775 2757 1776
rect 2751 1774 2757 1775
rect 2823 1775 2824 1779
rect 2828 1778 2829 1779
rect 2855 1779 2861 1780
rect 2855 1778 2856 1779
rect 2828 1776 2856 1778
rect 2828 1775 2829 1776
rect 2823 1774 2829 1775
rect 2855 1775 2856 1776
rect 2860 1775 2861 1779
rect 2855 1774 2861 1775
rect 2927 1779 2933 1780
rect 2927 1775 2928 1779
rect 2932 1778 2933 1779
rect 2959 1779 2965 1780
rect 2959 1778 2960 1779
rect 2932 1776 2960 1778
rect 2932 1775 2933 1776
rect 2927 1774 2933 1775
rect 2959 1775 2960 1776
rect 2964 1775 2965 1779
rect 2959 1774 2965 1775
rect 3031 1779 3037 1780
rect 3031 1775 3032 1779
rect 3036 1778 3037 1779
rect 3063 1779 3069 1780
rect 3063 1778 3064 1779
rect 3036 1776 3064 1778
rect 3036 1775 3037 1776
rect 3031 1774 3037 1775
rect 3063 1775 3064 1776
rect 3068 1775 3069 1779
rect 3063 1774 3069 1775
rect 3151 1779 3157 1780
rect 3151 1775 3152 1779
rect 3156 1778 3157 1779
rect 3167 1779 3173 1780
rect 3167 1778 3168 1779
rect 3156 1776 3168 1778
rect 3156 1775 3157 1776
rect 3151 1774 3157 1775
rect 3167 1775 3168 1776
rect 3172 1775 3173 1779
rect 3167 1774 3173 1775
rect 1702 1770 1708 1771
rect 2270 1769 2276 1770
rect 370 1767 376 1768
rect 370 1766 371 1767
rect 110 1765 116 1766
rect 110 1761 111 1765
rect 115 1761 116 1765
rect 361 1764 371 1766
rect 370 1763 371 1764
rect 375 1763 376 1767
rect 370 1762 376 1763
rect 839 1767 845 1768
rect 839 1763 840 1767
rect 844 1766 845 1767
rect 1114 1767 1120 1768
rect 844 1764 889 1766
rect 844 1763 845 1764
rect 839 1762 845 1763
rect 1114 1763 1115 1767
rect 1119 1766 1120 1767
rect 1119 1764 1233 1766
rect 1822 1765 1828 1766
rect 1119 1763 1120 1764
rect 1114 1762 1120 1763
rect 110 1760 116 1761
rect 1822 1761 1823 1765
rect 1827 1761 1828 1765
rect 2270 1765 2271 1769
rect 2275 1765 2276 1769
rect 2270 1764 2276 1765
rect 2358 1769 2364 1770
rect 2358 1765 2359 1769
rect 2363 1765 2364 1769
rect 2358 1764 2364 1765
rect 2454 1769 2460 1770
rect 2454 1765 2455 1769
rect 2459 1765 2460 1769
rect 2454 1764 2460 1765
rect 2558 1769 2564 1770
rect 2558 1765 2559 1769
rect 2563 1765 2564 1769
rect 2558 1764 2564 1765
rect 2662 1769 2668 1770
rect 2662 1765 2663 1769
rect 2667 1765 2668 1769
rect 2662 1764 2668 1765
rect 2758 1769 2764 1770
rect 2758 1765 2759 1769
rect 2763 1765 2764 1769
rect 2758 1764 2764 1765
rect 2862 1769 2868 1770
rect 2862 1765 2863 1769
rect 2867 1765 2868 1769
rect 2862 1764 2868 1765
rect 2966 1769 2972 1770
rect 2966 1765 2967 1769
rect 2971 1765 2972 1769
rect 2966 1764 2972 1765
rect 3070 1769 3076 1770
rect 3070 1765 3071 1769
rect 3075 1765 3076 1769
rect 3070 1764 3076 1765
rect 3174 1769 3180 1770
rect 3174 1765 3175 1769
rect 3179 1765 3180 1769
rect 3174 1764 3180 1765
rect 1822 1760 1828 1761
rect 1862 1756 1868 1757
rect 3574 1756 3580 1757
rect 1862 1752 1863 1756
rect 1867 1752 1868 1756
rect 2330 1755 2336 1756
rect 2330 1754 2331 1755
rect 2325 1752 2331 1754
rect 295 1751 301 1752
rect 295 1750 296 1751
rect 110 1748 116 1749
rect 197 1748 296 1750
rect 110 1744 111 1748
rect 115 1744 116 1748
rect 295 1747 296 1748
rect 300 1747 301 1751
rect 567 1751 573 1752
rect 567 1750 568 1751
rect 557 1748 568 1750
rect 295 1746 301 1747
rect 567 1747 568 1748
rect 572 1747 573 1751
rect 863 1751 869 1752
rect 863 1750 864 1751
rect 749 1748 864 1750
rect 567 1746 573 1747
rect 863 1747 864 1748
rect 868 1747 869 1751
rect 1207 1751 1213 1752
rect 1207 1750 1208 1751
rect 1109 1748 1208 1750
rect 863 1746 869 1747
rect 1207 1747 1208 1748
rect 1212 1747 1213 1751
rect 1519 1751 1525 1752
rect 1519 1750 1520 1751
rect 1437 1748 1520 1750
rect 1207 1746 1213 1747
rect 1519 1747 1520 1748
rect 1524 1747 1525 1751
rect 1519 1746 1525 1747
rect 1527 1751 1533 1752
rect 1527 1747 1528 1751
rect 1532 1750 1533 1751
rect 1695 1751 1701 1752
rect 1862 1751 1868 1752
rect 2330 1751 2331 1752
rect 2335 1751 2336 1755
rect 2823 1755 2829 1756
rect 2823 1754 2824 1755
rect 2813 1752 2824 1754
rect 1532 1748 1561 1750
rect 1532 1747 1533 1748
rect 1527 1746 1533 1747
rect 1695 1747 1696 1751
rect 1700 1750 1701 1751
rect 2330 1750 2336 1751
rect 2338 1751 2344 1752
rect 1700 1748 1729 1750
rect 1822 1748 1828 1749
rect 1700 1747 1701 1748
rect 1695 1746 1701 1747
rect 110 1743 116 1744
rect 1822 1744 1823 1748
rect 1827 1744 1828 1748
rect 2338 1747 2339 1751
rect 2343 1750 2344 1751
rect 2426 1751 2432 1752
rect 2343 1748 2377 1750
rect 2343 1747 2344 1748
rect 2338 1746 2344 1747
rect 2426 1747 2427 1751
rect 2431 1750 2432 1751
rect 2522 1751 2528 1752
rect 2431 1748 2473 1750
rect 2431 1747 2432 1748
rect 2426 1746 2432 1747
rect 2522 1747 2523 1751
rect 2527 1750 2528 1751
rect 2631 1751 2637 1752
rect 2527 1748 2577 1750
rect 2527 1747 2528 1748
rect 2522 1746 2528 1747
rect 2631 1747 2632 1751
rect 2636 1750 2637 1751
rect 2823 1751 2824 1752
rect 2828 1751 2829 1755
rect 2927 1755 2933 1756
rect 2927 1754 2928 1755
rect 2917 1752 2928 1754
rect 2823 1750 2829 1751
rect 2927 1751 2928 1752
rect 2932 1751 2933 1755
rect 3031 1755 3037 1756
rect 3031 1754 3032 1755
rect 3021 1752 3032 1754
rect 2927 1750 2933 1751
rect 3031 1751 3032 1752
rect 3036 1751 3037 1755
rect 3151 1755 3157 1756
rect 3151 1754 3152 1755
rect 3125 1752 3152 1754
rect 3031 1750 3037 1751
rect 3151 1751 3152 1752
rect 3156 1751 3157 1755
rect 3574 1752 3575 1756
rect 3579 1752 3580 1756
rect 3574 1751 3580 1752
rect 3151 1750 3157 1751
rect 2636 1748 2681 1750
rect 2636 1747 2637 1748
rect 2631 1746 2637 1747
rect 1822 1743 1828 1744
rect 1862 1739 1868 1740
rect 142 1735 148 1736
rect 142 1731 143 1735
rect 147 1731 148 1735
rect 142 1730 148 1731
rect 310 1735 316 1736
rect 310 1731 311 1735
rect 315 1731 316 1735
rect 310 1730 316 1731
rect 502 1735 508 1736
rect 502 1731 503 1735
rect 507 1731 508 1735
rect 502 1730 508 1731
rect 694 1735 700 1736
rect 694 1731 695 1735
rect 699 1731 700 1735
rect 694 1730 700 1731
rect 878 1735 884 1736
rect 878 1731 879 1735
rect 883 1731 884 1735
rect 878 1730 884 1731
rect 1054 1735 1060 1736
rect 1054 1731 1055 1735
rect 1059 1731 1060 1735
rect 1054 1730 1060 1731
rect 1222 1735 1228 1736
rect 1222 1731 1223 1735
rect 1227 1731 1228 1735
rect 1222 1730 1228 1731
rect 1382 1735 1388 1736
rect 1382 1731 1383 1735
rect 1387 1731 1388 1735
rect 1382 1730 1388 1731
rect 1542 1735 1548 1736
rect 1542 1731 1543 1735
rect 1547 1731 1548 1735
rect 1542 1730 1548 1731
rect 1710 1735 1716 1736
rect 1710 1731 1711 1735
rect 1715 1731 1716 1735
rect 1862 1735 1863 1739
rect 1867 1735 1868 1739
rect 3574 1739 3580 1740
rect 1862 1734 1868 1735
rect 3139 1736 3185 1738
rect 1710 1730 1716 1731
rect 2262 1729 2268 1730
rect 2262 1725 2263 1729
rect 2267 1725 2268 1729
rect 2262 1724 2268 1725
rect 2350 1729 2356 1730
rect 2350 1725 2351 1729
rect 2355 1725 2356 1729
rect 2350 1724 2356 1725
rect 2446 1729 2452 1730
rect 2446 1725 2447 1729
rect 2451 1725 2452 1729
rect 2446 1724 2452 1725
rect 2550 1729 2556 1730
rect 2550 1725 2551 1729
rect 2555 1725 2556 1729
rect 2550 1724 2556 1725
rect 2654 1729 2660 1730
rect 2654 1725 2655 1729
rect 2659 1725 2660 1729
rect 2654 1724 2660 1725
rect 2750 1729 2756 1730
rect 2750 1725 2751 1729
rect 2755 1725 2756 1729
rect 2750 1724 2756 1725
rect 2854 1729 2860 1730
rect 2854 1725 2855 1729
rect 2859 1725 2860 1729
rect 2854 1724 2860 1725
rect 2958 1729 2964 1730
rect 2958 1725 2959 1729
rect 2963 1725 2964 1729
rect 2958 1724 2964 1725
rect 3062 1729 3068 1730
rect 3062 1725 3063 1729
rect 3067 1725 3068 1729
rect 3062 1724 3068 1725
rect 134 1723 141 1724
rect 134 1719 135 1723
rect 140 1719 141 1723
rect 134 1718 141 1719
rect 295 1723 301 1724
rect 295 1719 296 1723
rect 300 1722 301 1723
rect 303 1723 309 1724
rect 303 1722 304 1723
rect 300 1720 304 1722
rect 300 1719 301 1720
rect 295 1718 301 1719
rect 303 1719 304 1720
rect 308 1719 309 1723
rect 303 1718 309 1719
rect 495 1723 501 1724
rect 495 1719 496 1723
rect 500 1722 501 1723
rect 510 1723 516 1724
rect 510 1722 511 1723
rect 500 1720 511 1722
rect 500 1719 501 1720
rect 495 1718 501 1719
rect 510 1719 511 1720
rect 515 1719 516 1723
rect 510 1718 516 1719
rect 567 1723 573 1724
rect 567 1719 568 1723
rect 572 1722 573 1723
rect 687 1723 693 1724
rect 687 1722 688 1723
rect 572 1720 688 1722
rect 572 1719 573 1720
rect 567 1718 573 1719
rect 687 1719 688 1720
rect 692 1719 693 1723
rect 687 1718 693 1719
rect 863 1723 869 1724
rect 863 1719 864 1723
rect 868 1722 869 1723
rect 871 1723 877 1724
rect 871 1722 872 1723
rect 868 1720 872 1722
rect 868 1719 869 1720
rect 863 1718 869 1719
rect 871 1719 872 1720
rect 876 1719 877 1723
rect 871 1718 877 1719
rect 1047 1723 1053 1724
rect 1047 1719 1048 1723
rect 1052 1722 1053 1723
rect 1082 1723 1088 1724
rect 1082 1722 1083 1723
rect 1052 1720 1083 1722
rect 1052 1719 1053 1720
rect 1047 1718 1053 1719
rect 1082 1719 1083 1720
rect 1087 1719 1088 1723
rect 1082 1718 1088 1719
rect 1207 1723 1213 1724
rect 1207 1719 1208 1723
rect 1212 1722 1213 1723
rect 1215 1723 1221 1724
rect 1215 1722 1216 1723
rect 1212 1720 1216 1722
rect 1212 1719 1213 1720
rect 1207 1718 1213 1719
rect 1215 1719 1216 1720
rect 1220 1719 1221 1723
rect 1215 1718 1221 1719
rect 1375 1723 1381 1724
rect 1375 1719 1376 1723
rect 1380 1722 1381 1723
rect 1390 1723 1396 1724
rect 1390 1722 1391 1723
rect 1380 1720 1391 1722
rect 1380 1719 1381 1720
rect 1375 1718 1381 1719
rect 1390 1719 1391 1720
rect 1395 1719 1396 1723
rect 1390 1718 1396 1719
rect 1535 1723 1541 1724
rect 1535 1719 1536 1723
rect 1540 1722 1541 1723
rect 1550 1723 1556 1724
rect 1550 1722 1551 1723
rect 1540 1720 1551 1722
rect 1540 1719 1541 1720
rect 1535 1718 1541 1719
rect 1550 1719 1551 1720
rect 1555 1719 1556 1723
rect 1703 1723 1709 1724
rect 1703 1722 1704 1723
rect 1550 1718 1556 1719
rect 1584 1720 1704 1722
rect 1519 1715 1525 1716
rect 1519 1711 1520 1715
rect 1524 1714 1525 1715
rect 1584 1714 1586 1720
rect 1703 1719 1704 1720
rect 1708 1719 1709 1723
rect 1703 1718 1709 1719
rect 2902 1723 2908 1724
rect 2902 1719 2903 1723
rect 2907 1722 2908 1723
rect 3139 1722 3141 1736
rect 3574 1735 3575 1739
rect 3579 1735 3580 1739
rect 3574 1734 3580 1735
rect 3166 1729 3172 1730
rect 3166 1725 3167 1729
rect 3171 1725 3172 1729
rect 3166 1724 3172 1725
rect 2907 1720 3141 1722
rect 2907 1719 2908 1720
rect 2902 1718 2908 1719
rect 1524 1712 1586 1714
rect 1524 1711 1525 1712
rect 1519 1710 1525 1711
rect 127 1707 133 1708
rect 127 1703 128 1707
rect 132 1706 133 1707
rect 135 1707 141 1708
rect 135 1706 136 1707
rect 132 1704 136 1706
rect 132 1703 133 1704
rect 127 1702 133 1703
rect 135 1703 136 1704
rect 140 1703 141 1707
rect 135 1702 141 1703
rect 279 1707 285 1708
rect 279 1703 280 1707
rect 284 1706 285 1707
rect 382 1707 388 1708
rect 382 1706 383 1707
rect 284 1704 383 1706
rect 284 1703 285 1704
rect 279 1702 285 1703
rect 382 1703 383 1704
rect 387 1703 388 1707
rect 382 1702 388 1703
rect 463 1707 469 1708
rect 463 1703 464 1707
rect 468 1706 469 1707
rect 599 1707 605 1708
rect 599 1706 600 1707
rect 468 1704 600 1706
rect 468 1703 469 1704
rect 463 1702 469 1703
rect 599 1703 600 1704
rect 604 1703 605 1707
rect 599 1702 605 1703
rect 647 1707 653 1708
rect 647 1703 648 1707
rect 652 1706 653 1707
rect 750 1707 756 1708
rect 750 1706 751 1707
rect 652 1704 751 1706
rect 652 1703 653 1704
rect 647 1702 653 1703
rect 750 1703 751 1704
rect 755 1703 756 1707
rect 750 1702 756 1703
rect 831 1707 837 1708
rect 831 1703 832 1707
rect 836 1706 837 1707
rect 839 1707 845 1708
rect 839 1706 840 1707
rect 836 1704 840 1706
rect 836 1703 837 1704
rect 831 1702 837 1703
rect 839 1703 840 1704
rect 844 1703 845 1707
rect 839 1702 845 1703
rect 998 1707 1004 1708
rect 998 1703 999 1707
rect 1003 1706 1004 1707
rect 1015 1707 1021 1708
rect 1015 1706 1016 1707
rect 1003 1704 1016 1706
rect 1003 1703 1004 1704
rect 998 1702 1004 1703
rect 1015 1703 1016 1704
rect 1020 1703 1021 1707
rect 1015 1702 1021 1703
rect 1183 1707 1189 1708
rect 1183 1703 1184 1707
rect 1188 1706 1189 1707
rect 1263 1707 1269 1708
rect 1263 1706 1264 1707
rect 1188 1704 1264 1706
rect 1188 1703 1189 1704
rect 1183 1702 1189 1703
rect 1263 1703 1264 1704
rect 1268 1703 1269 1707
rect 1263 1702 1269 1703
rect 1351 1707 1357 1708
rect 1351 1703 1352 1707
rect 1356 1706 1357 1707
rect 1426 1707 1432 1708
rect 1426 1706 1427 1707
rect 1356 1704 1427 1706
rect 1356 1703 1357 1704
rect 1351 1702 1357 1703
rect 1426 1703 1427 1704
rect 1431 1703 1432 1707
rect 1426 1702 1432 1703
rect 1519 1707 1525 1708
rect 1519 1703 1520 1707
rect 1524 1706 1525 1707
rect 1527 1707 1533 1708
rect 1527 1706 1528 1707
rect 1524 1704 1528 1706
rect 1524 1703 1525 1704
rect 1519 1702 1525 1703
rect 1527 1703 1528 1704
rect 1532 1703 1533 1707
rect 1527 1702 1533 1703
rect 1687 1707 1693 1708
rect 1687 1703 1688 1707
rect 1692 1706 1693 1707
rect 1695 1707 1701 1708
rect 1695 1706 1696 1707
rect 1692 1704 1696 1706
rect 1692 1703 1693 1704
rect 1687 1702 1693 1703
rect 1695 1703 1696 1704
rect 1700 1703 1701 1707
rect 1695 1702 1701 1703
rect 2246 1703 2252 1704
rect 2246 1699 2247 1703
rect 2251 1699 2252 1703
rect 2246 1698 2252 1699
rect 2366 1703 2372 1704
rect 2366 1699 2367 1703
rect 2371 1699 2372 1703
rect 2366 1698 2372 1699
rect 2494 1703 2500 1704
rect 2494 1699 2495 1703
rect 2499 1699 2500 1703
rect 2494 1698 2500 1699
rect 2622 1703 2628 1704
rect 2622 1699 2623 1703
rect 2627 1699 2628 1703
rect 2622 1698 2628 1699
rect 2758 1703 2764 1704
rect 2758 1699 2759 1703
rect 2763 1699 2764 1703
rect 2758 1698 2764 1699
rect 2886 1703 2892 1704
rect 2886 1699 2887 1703
rect 2891 1699 2892 1703
rect 2886 1698 2892 1699
rect 3014 1703 3020 1704
rect 3014 1699 3015 1703
rect 3019 1699 3020 1703
rect 3014 1698 3020 1699
rect 3134 1703 3140 1704
rect 3134 1699 3135 1703
rect 3139 1699 3140 1703
rect 3134 1698 3140 1699
rect 3246 1703 3252 1704
rect 3246 1699 3247 1703
rect 3251 1699 3252 1703
rect 3246 1698 3252 1699
rect 3366 1703 3372 1704
rect 3366 1699 3367 1703
rect 3371 1699 3372 1703
rect 3366 1698 3372 1699
rect 3478 1703 3484 1704
rect 3478 1699 3479 1703
rect 3483 1699 3484 1703
rect 3478 1698 3484 1699
rect 142 1697 148 1698
rect 142 1693 143 1697
rect 147 1693 148 1697
rect 142 1692 148 1693
rect 286 1697 292 1698
rect 286 1693 287 1697
rect 291 1693 292 1697
rect 286 1692 292 1693
rect 470 1697 476 1698
rect 470 1693 471 1697
rect 475 1693 476 1697
rect 470 1692 476 1693
rect 654 1697 660 1698
rect 654 1693 655 1697
rect 659 1693 660 1697
rect 654 1692 660 1693
rect 838 1697 844 1698
rect 838 1693 839 1697
rect 843 1693 844 1697
rect 838 1692 844 1693
rect 1022 1697 1028 1698
rect 1022 1693 1023 1697
rect 1027 1693 1028 1697
rect 1022 1692 1028 1693
rect 1190 1697 1196 1698
rect 1190 1693 1191 1697
rect 1195 1693 1196 1697
rect 1190 1692 1196 1693
rect 1358 1697 1364 1698
rect 1358 1693 1359 1697
rect 1363 1693 1364 1697
rect 1358 1692 1364 1693
rect 1526 1697 1532 1698
rect 1526 1693 1527 1697
rect 1531 1693 1532 1697
rect 1526 1692 1532 1693
rect 1694 1697 1700 1698
rect 1694 1693 1695 1697
rect 1699 1693 1700 1697
rect 2722 1695 2728 1696
rect 1694 1692 1700 1693
rect 1862 1693 1868 1694
rect 1862 1689 1863 1693
rect 1867 1689 1868 1693
rect 2722 1691 2723 1695
rect 2727 1694 2728 1695
rect 3351 1695 3357 1696
rect 2727 1692 2777 1694
rect 2727 1691 2728 1692
rect 2722 1690 2728 1691
rect 3351 1691 3352 1695
rect 3356 1694 3357 1695
rect 3356 1692 3385 1694
rect 3574 1693 3580 1694
rect 3356 1691 3357 1692
rect 3351 1690 3357 1691
rect 1862 1688 1868 1689
rect 3574 1689 3575 1693
rect 3579 1689 3580 1693
rect 3574 1688 3580 1689
rect 110 1684 116 1685
rect 1822 1684 1828 1685
rect 110 1680 111 1684
rect 115 1680 116 1684
rect 1082 1683 1088 1684
rect 1082 1682 1083 1683
rect 1077 1680 1083 1682
rect 110 1679 116 1680
rect 134 1679 140 1680
rect 134 1675 135 1679
rect 139 1678 140 1679
rect 382 1679 388 1680
rect 139 1676 161 1678
rect 139 1675 140 1676
rect 134 1674 140 1675
rect 382 1675 383 1679
rect 387 1678 388 1679
rect 599 1679 605 1680
rect 387 1676 489 1678
rect 387 1675 388 1676
rect 382 1674 388 1675
rect 599 1675 600 1679
rect 604 1678 605 1679
rect 750 1679 756 1680
rect 604 1676 673 1678
rect 604 1675 605 1676
rect 599 1674 605 1675
rect 750 1675 751 1679
rect 755 1678 756 1679
rect 1082 1679 1083 1680
rect 1087 1679 1088 1683
rect 1822 1680 1823 1684
rect 1827 1680 1828 1684
rect 1082 1678 1088 1679
rect 1263 1679 1269 1680
rect 755 1676 857 1678
rect 755 1675 756 1676
rect 750 1674 756 1675
rect 1263 1675 1264 1679
rect 1268 1678 1269 1679
rect 1426 1679 1432 1680
rect 1822 1679 1828 1680
rect 2359 1679 2365 1680
rect 1268 1676 1377 1678
rect 1268 1675 1269 1676
rect 1263 1674 1269 1675
rect 1426 1675 1427 1679
rect 1431 1678 1432 1679
rect 2359 1678 2360 1679
rect 1431 1676 1545 1678
rect 1862 1676 1868 1677
rect 2309 1676 2360 1678
rect 1431 1675 1432 1676
rect 1426 1674 1432 1675
rect 1862 1672 1863 1676
rect 1867 1672 1868 1676
rect 2359 1675 2360 1676
rect 2364 1675 2365 1679
rect 2487 1679 2493 1680
rect 2487 1678 2488 1679
rect 2429 1676 2488 1678
rect 2359 1674 2365 1675
rect 2487 1675 2488 1676
rect 2492 1675 2493 1679
rect 2615 1679 2621 1680
rect 2615 1678 2616 1679
rect 2557 1676 2616 1678
rect 2487 1674 2493 1675
rect 2615 1675 2616 1676
rect 2620 1675 2621 1679
rect 2751 1679 2757 1680
rect 2751 1678 2752 1679
rect 2685 1676 2752 1678
rect 2615 1674 2621 1675
rect 2751 1675 2752 1676
rect 2756 1675 2757 1679
rect 3007 1679 3013 1680
rect 3007 1678 3008 1679
rect 2949 1676 3008 1678
rect 2751 1674 2757 1675
rect 3007 1675 3008 1676
rect 3012 1675 3013 1679
rect 3126 1679 3132 1680
rect 3126 1678 3127 1679
rect 3077 1676 3127 1678
rect 3007 1674 3013 1675
rect 3126 1675 3127 1676
rect 3131 1675 3132 1679
rect 3239 1679 3245 1680
rect 3239 1678 3240 1679
rect 3197 1676 3240 1678
rect 3126 1674 3132 1675
rect 3239 1675 3240 1676
rect 3244 1675 3245 1679
rect 3359 1679 3365 1680
rect 3359 1678 3360 1679
rect 3309 1676 3360 1678
rect 3239 1674 3245 1675
rect 3359 1675 3360 1676
rect 3364 1675 3365 1679
rect 3359 1674 3365 1675
rect 3471 1679 3477 1680
rect 3471 1675 3472 1679
rect 3476 1678 3477 1679
rect 3476 1676 3505 1678
rect 3574 1676 3580 1677
rect 3476 1675 3477 1676
rect 3471 1674 3477 1675
rect 1862 1671 1868 1672
rect 3574 1672 3575 1676
rect 3579 1672 3580 1676
rect 3574 1671 3580 1672
rect 110 1667 116 1668
rect 110 1663 111 1667
rect 115 1663 116 1667
rect 110 1662 116 1663
rect 286 1667 292 1668
rect 286 1663 287 1667
rect 291 1666 292 1667
rect 1166 1667 1172 1668
rect 291 1664 297 1666
rect 291 1663 292 1664
rect 286 1662 292 1663
rect 1166 1663 1167 1667
rect 1171 1666 1172 1667
rect 1822 1667 1828 1668
rect 1171 1664 1201 1666
rect 1171 1663 1172 1664
rect 1166 1662 1172 1663
rect 1822 1663 1823 1667
rect 1827 1663 1828 1667
rect 1822 1662 1828 1663
rect 2254 1663 2260 1664
rect 2254 1659 2255 1663
rect 2259 1659 2260 1663
rect 2254 1658 2260 1659
rect 2374 1663 2380 1664
rect 2374 1659 2375 1663
rect 2379 1659 2380 1663
rect 2374 1658 2380 1659
rect 2502 1663 2508 1664
rect 2502 1659 2503 1663
rect 2507 1659 2508 1663
rect 2502 1658 2508 1659
rect 2630 1663 2636 1664
rect 2630 1659 2631 1663
rect 2635 1659 2636 1663
rect 2630 1658 2636 1659
rect 2766 1663 2772 1664
rect 2766 1659 2767 1663
rect 2771 1659 2772 1663
rect 2766 1658 2772 1659
rect 2894 1663 2900 1664
rect 2894 1659 2895 1663
rect 2899 1659 2900 1663
rect 2894 1658 2900 1659
rect 3022 1663 3028 1664
rect 3022 1659 3023 1663
rect 3027 1659 3028 1663
rect 3022 1658 3028 1659
rect 3142 1663 3148 1664
rect 3142 1659 3143 1663
rect 3147 1659 3148 1663
rect 3142 1658 3148 1659
rect 3254 1663 3260 1664
rect 3254 1659 3255 1663
rect 3259 1659 3260 1663
rect 3254 1658 3260 1659
rect 3374 1663 3380 1664
rect 3374 1659 3375 1663
rect 3379 1659 3380 1663
rect 3374 1658 3380 1659
rect 3486 1663 3492 1664
rect 3486 1659 3487 1663
rect 3491 1659 3492 1663
rect 3486 1658 3492 1659
rect 134 1657 140 1658
rect 134 1653 135 1657
rect 139 1653 140 1657
rect 134 1652 140 1653
rect 278 1657 284 1658
rect 278 1653 279 1657
rect 283 1653 284 1657
rect 278 1652 284 1653
rect 462 1657 468 1658
rect 462 1653 463 1657
rect 467 1653 468 1657
rect 462 1652 468 1653
rect 646 1657 652 1658
rect 646 1653 647 1657
rect 651 1653 652 1657
rect 646 1652 652 1653
rect 830 1657 836 1658
rect 830 1653 831 1657
rect 835 1653 836 1657
rect 830 1652 836 1653
rect 1014 1657 1020 1658
rect 1014 1653 1015 1657
rect 1019 1653 1020 1657
rect 1014 1652 1020 1653
rect 1182 1657 1188 1658
rect 1182 1653 1183 1657
rect 1187 1653 1188 1657
rect 1182 1652 1188 1653
rect 1350 1657 1356 1658
rect 1350 1653 1351 1657
rect 1355 1653 1356 1657
rect 1350 1652 1356 1653
rect 1518 1657 1524 1658
rect 1518 1653 1519 1657
rect 1523 1653 1524 1657
rect 1518 1652 1524 1653
rect 1686 1657 1692 1658
rect 1686 1653 1687 1657
rect 1691 1653 1692 1657
rect 1686 1652 1692 1653
rect 1719 1651 1725 1652
rect 1719 1647 1720 1651
rect 1724 1650 1725 1651
rect 1735 1651 1741 1652
rect 1735 1650 1736 1651
rect 1724 1648 1736 1650
rect 1724 1647 1725 1648
rect 1719 1646 1725 1647
rect 1735 1647 1736 1648
rect 1740 1647 1741 1651
rect 1735 1646 1741 1647
rect 2247 1651 2253 1652
rect 2247 1647 2248 1651
rect 2252 1650 2253 1651
rect 2359 1651 2365 1652
rect 2252 1648 2301 1650
rect 2252 1647 2253 1648
rect 2247 1646 2253 1647
rect 2299 1642 2301 1648
rect 2359 1647 2360 1651
rect 2364 1650 2365 1651
rect 2367 1651 2373 1652
rect 2367 1650 2368 1651
rect 2364 1648 2368 1650
rect 2364 1647 2365 1648
rect 2359 1646 2365 1647
rect 2367 1647 2368 1648
rect 2372 1647 2373 1651
rect 2367 1646 2373 1647
rect 2487 1651 2493 1652
rect 2487 1647 2488 1651
rect 2492 1650 2493 1651
rect 2495 1651 2501 1652
rect 2495 1650 2496 1651
rect 2492 1648 2496 1650
rect 2492 1647 2493 1648
rect 2487 1646 2493 1647
rect 2495 1647 2496 1648
rect 2500 1647 2501 1651
rect 2495 1646 2501 1647
rect 2615 1651 2621 1652
rect 2615 1647 2616 1651
rect 2620 1650 2621 1651
rect 2623 1651 2629 1652
rect 2623 1650 2624 1651
rect 2620 1648 2624 1650
rect 2620 1647 2621 1648
rect 2615 1646 2621 1647
rect 2623 1647 2624 1648
rect 2628 1647 2629 1651
rect 2623 1646 2629 1647
rect 2751 1651 2757 1652
rect 2751 1647 2752 1651
rect 2756 1650 2757 1651
rect 2759 1651 2765 1652
rect 2759 1650 2760 1651
rect 2756 1648 2760 1650
rect 2756 1647 2757 1648
rect 2751 1646 2757 1647
rect 2759 1647 2760 1648
rect 2764 1647 2765 1651
rect 2759 1646 2765 1647
rect 2887 1651 2893 1652
rect 2887 1647 2888 1651
rect 2892 1650 2893 1651
rect 2902 1651 2908 1652
rect 2902 1650 2903 1651
rect 2892 1648 2903 1650
rect 2892 1647 2893 1648
rect 2887 1646 2893 1647
rect 2902 1647 2903 1648
rect 2907 1647 2908 1651
rect 2902 1646 2908 1647
rect 3007 1651 3013 1652
rect 3007 1647 3008 1651
rect 3012 1650 3013 1651
rect 3015 1651 3021 1652
rect 3015 1650 3016 1651
rect 3012 1648 3016 1650
rect 3012 1647 3013 1648
rect 3007 1646 3013 1647
rect 3015 1647 3016 1648
rect 3020 1647 3021 1651
rect 3015 1646 3021 1647
rect 3126 1651 3132 1652
rect 3126 1647 3127 1651
rect 3131 1650 3132 1651
rect 3135 1651 3141 1652
rect 3135 1650 3136 1651
rect 3131 1648 3136 1650
rect 3131 1647 3132 1648
rect 3126 1646 3132 1647
rect 3135 1647 3136 1648
rect 3140 1647 3141 1651
rect 3135 1646 3141 1647
rect 3239 1651 3245 1652
rect 3239 1647 3240 1651
rect 3244 1650 3245 1651
rect 3247 1651 3253 1652
rect 3247 1650 3248 1651
rect 3244 1648 3248 1650
rect 3244 1647 3245 1648
rect 3239 1646 3245 1647
rect 3247 1647 3248 1648
rect 3252 1647 3253 1651
rect 3247 1646 3253 1647
rect 3359 1651 3365 1652
rect 3359 1647 3360 1651
rect 3364 1650 3365 1651
rect 3367 1651 3373 1652
rect 3367 1650 3368 1651
rect 3364 1648 3368 1650
rect 3364 1647 3365 1648
rect 3359 1646 3365 1647
rect 3367 1647 3368 1648
rect 3372 1647 3373 1651
rect 3367 1646 3373 1647
rect 3479 1651 3485 1652
rect 3479 1647 3480 1651
rect 3484 1650 3485 1651
rect 3498 1651 3504 1652
rect 3498 1650 3499 1651
rect 3484 1648 3499 1650
rect 3484 1647 3485 1648
rect 3479 1646 3485 1647
rect 3498 1647 3499 1648
rect 3503 1647 3504 1651
rect 3498 1646 3504 1647
rect 2623 1643 2629 1644
rect 2623 1642 2624 1643
rect 2299 1640 2624 1642
rect 2623 1639 2624 1640
rect 2628 1639 2629 1643
rect 3098 1643 3104 1644
rect 3098 1642 3099 1643
rect 2623 1638 2629 1639
rect 2945 1640 3099 1642
rect 2143 1635 2149 1636
rect 2143 1631 2144 1635
rect 2148 1634 2149 1635
rect 2158 1635 2164 1636
rect 2158 1634 2159 1635
rect 2148 1632 2159 1634
rect 2148 1631 2149 1632
rect 2143 1630 2149 1631
rect 2158 1631 2159 1632
rect 2163 1631 2164 1635
rect 2158 1630 2164 1631
rect 2215 1635 2221 1636
rect 2215 1631 2216 1635
rect 2220 1634 2221 1635
rect 2335 1635 2341 1636
rect 2335 1634 2336 1635
rect 2220 1632 2336 1634
rect 2220 1631 2221 1632
rect 2215 1630 2221 1631
rect 2335 1631 2336 1632
rect 2340 1631 2341 1635
rect 2335 1630 2341 1631
rect 2431 1635 2437 1636
rect 2431 1631 2432 1635
rect 2436 1634 2437 1635
rect 2519 1635 2525 1636
rect 2519 1634 2520 1635
rect 2436 1632 2520 1634
rect 2436 1631 2437 1632
rect 2431 1630 2437 1631
rect 2519 1631 2520 1632
rect 2524 1631 2525 1635
rect 2519 1630 2525 1631
rect 2615 1635 2621 1636
rect 2615 1631 2616 1635
rect 2620 1634 2621 1635
rect 2695 1635 2701 1636
rect 2695 1634 2696 1635
rect 2620 1632 2696 1634
rect 2620 1631 2621 1632
rect 2615 1630 2621 1631
rect 2695 1631 2696 1632
rect 2700 1631 2701 1635
rect 2695 1630 2701 1631
rect 2863 1635 2869 1636
rect 2863 1631 2864 1635
rect 2868 1634 2869 1635
rect 2945 1634 2947 1640
rect 3098 1639 3099 1640
rect 3103 1639 3104 1643
rect 3098 1638 3104 1639
rect 2868 1632 2947 1634
rect 2951 1635 2957 1636
rect 2868 1631 2869 1632
rect 2863 1630 2869 1631
rect 2951 1631 2952 1635
rect 2956 1634 2957 1635
rect 3023 1635 3029 1636
rect 3023 1634 3024 1635
rect 2956 1632 3024 1634
rect 2956 1631 2957 1632
rect 2951 1630 2957 1631
rect 3023 1631 3024 1632
rect 3028 1631 3029 1635
rect 3023 1630 3029 1631
rect 3183 1635 3189 1636
rect 3183 1631 3184 1635
rect 3188 1634 3189 1635
rect 3271 1635 3277 1636
rect 3271 1634 3272 1635
rect 3188 1632 3272 1634
rect 3188 1631 3189 1632
rect 3183 1630 3189 1631
rect 3271 1631 3272 1632
rect 3276 1631 3277 1635
rect 3271 1630 3277 1631
rect 3343 1635 3349 1636
rect 3343 1631 3344 1635
rect 3348 1634 3349 1635
rect 3351 1635 3357 1636
rect 3351 1634 3352 1635
rect 3348 1632 3352 1634
rect 3348 1631 3349 1632
rect 3343 1630 3349 1631
rect 3351 1631 3352 1632
rect 3356 1631 3357 1635
rect 3351 1630 3357 1631
rect 3471 1635 3477 1636
rect 3471 1631 3472 1635
rect 3476 1634 3477 1635
rect 3479 1635 3485 1636
rect 3479 1634 3480 1635
rect 3476 1632 3480 1634
rect 3476 1631 3477 1632
rect 3471 1630 3477 1631
rect 3479 1631 3480 1632
rect 3484 1631 3485 1635
rect 3479 1630 3485 1631
rect 134 1627 140 1628
rect 134 1623 135 1627
rect 139 1623 140 1627
rect 134 1622 140 1623
rect 270 1627 276 1628
rect 270 1623 271 1627
rect 275 1623 276 1627
rect 270 1622 276 1623
rect 446 1627 452 1628
rect 446 1623 447 1627
rect 451 1623 452 1627
rect 446 1622 452 1623
rect 630 1627 636 1628
rect 630 1623 631 1627
rect 635 1623 636 1627
rect 630 1622 636 1623
rect 814 1627 820 1628
rect 814 1623 815 1627
rect 819 1623 820 1627
rect 814 1622 820 1623
rect 990 1627 996 1628
rect 990 1623 991 1627
rect 995 1623 996 1627
rect 990 1622 996 1623
rect 1150 1627 1156 1628
rect 1150 1623 1151 1627
rect 1155 1623 1156 1627
rect 1150 1622 1156 1623
rect 1302 1627 1308 1628
rect 1302 1623 1303 1627
rect 1307 1623 1308 1627
rect 1302 1622 1308 1623
rect 1454 1627 1460 1628
rect 1454 1623 1455 1627
rect 1459 1623 1460 1627
rect 1454 1622 1460 1623
rect 1598 1627 1604 1628
rect 1598 1623 1599 1627
rect 1603 1623 1604 1627
rect 1598 1622 1604 1623
rect 1726 1627 1732 1628
rect 1726 1623 1727 1627
rect 1731 1623 1732 1627
rect 1726 1622 1732 1623
rect 2150 1625 2156 1626
rect 2150 1621 2151 1625
rect 2155 1621 2156 1625
rect 2150 1620 2156 1621
rect 2342 1625 2348 1626
rect 2342 1621 2343 1625
rect 2347 1621 2348 1625
rect 2342 1620 2348 1621
rect 2526 1625 2532 1626
rect 2526 1621 2527 1625
rect 2531 1621 2532 1625
rect 2526 1620 2532 1621
rect 2702 1625 2708 1626
rect 2702 1621 2703 1625
rect 2707 1621 2708 1625
rect 2702 1620 2708 1621
rect 2870 1625 2876 1626
rect 2870 1621 2871 1625
rect 2875 1621 2876 1625
rect 2870 1620 2876 1621
rect 3030 1625 3036 1626
rect 3030 1621 3031 1625
rect 3035 1621 3036 1625
rect 3030 1620 3036 1621
rect 3190 1625 3196 1626
rect 3190 1621 3191 1625
rect 3195 1621 3196 1625
rect 3190 1620 3196 1621
rect 3350 1625 3356 1626
rect 3350 1621 3351 1625
rect 3355 1621 3356 1625
rect 3350 1620 3356 1621
rect 3486 1625 3492 1626
rect 3486 1621 3487 1625
rect 3491 1621 3492 1625
rect 3486 1620 3492 1621
rect 127 1619 133 1620
rect 110 1617 116 1618
rect 110 1613 111 1617
rect 115 1613 116 1617
rect 127 1615 128 1619
rect 132 1618 133 1619
rect 767 1619 773 1620
rect 132 1616 153 1618
rect 132 1615 133 1616
rect 127 1614 133 1615
rect 767 1615 768 1619
rect 772 1618 773 1619
rect 1263 1619 1269 1620
rect 772 1616 833 1618
rect 1000 1616 1009 1618
rect 772 1615 773 1616
rect 767 1614 773 1615
rect 998 1615 1004 1616
rect 110 1612 116 1613
rect 998 1611 999 1615
rect 1003 1611 1004 1615
rect 1263 1615 1264 1619
rect 1268 1618 1269 1619
rect 1268 1616 1321 1618
rect 1822 1617 1828 1618
rect 1268 1615 1269 1616
rect 1263 1614 1269 1615
rect 1822 1613 1823 1617
rect 1827 1613 1828 1617
rect 1822 1612 1828 1613
rect 1862 1612 1868 1613
rect 3574 1612 3580 1613
rect 998 1610 1004 1611
rect 1862 1608 1863 1612
rect 1867 1608 1868 1612
rect 2215 1611 2221 1612
rect 2215 1610 2216 1611
rect 2205 1608 2216 1610
rect 1862 1607 1868 1608
rect 2215 1607 2216 1608
rect 2220 1607 2221 1611
rect 2431 1611 2437 1612
rect 2431 1610 2432 1611
rect 2397 1608 2432 1610
rect 2215 1606 2221 1607
rect 2431 1607 2432 1608
rect 2436 1607 2437 1611
rect 2615 1611 2621 1612
rect 2615 1610 2616 1611
rect 2581 1608 2616 1610
rect 2431 1606 2437 1607
rect 2615 1607 2616 1608
rect 2620 1607 2621 1611
rect 2951 1611 2957 1612
rect 2951 1610 2952 1611
rect 2925 1608 2952 1610
rect 2615 1606 2621 1607
rect 2623 1607 2629 1608
rect 439 1603 445 1604
rect 439 1602 440 1603
rect 110 1600 116 1601
rect 333 1600 440 1602
rect 110 1596 111 1600
rect 115 1596 116 1600
rect 439 1599 440 1600
rect 444 1599 445 1603
rect 623 1603 629 1604
rect 623 1602 624 1603
rect 509 1600 624 1602
rect 439 1598 445 1599
rect 623 1599 624 1600
rect 628 1599 629 1603
rect 807 1603 813 1604
rect 807 1602 808 1603
rect 693 1600 808 1602
rect 623 1598 629 1599
rect 807 1599 808 1600
rect 812 1599 813 1603
rect 1295 1603 1301 1604
rect 1295 1602 1296 1603
rect 1213 1600 1296 1602
rect 807 1598 813 1599
rect 1295 1599 1296 1600
rect 1300 1599 1301 1603
rect 1582 1603 1588 1604
rect 1582 1602 1583 1603
rect 1517 1600 1583 1602
rect 1295 1598 1301 1599
rect 1582 1599 1583 1600
rect 1587 1599 1588 1603
rect 1582 1598 1588 1599
rect 1591 1603 1597 1604
rect 1591 1599 1592 1603
rect 1596 1602 1597 1603
rect 1666 1603 1672 1604
rect 1596 1600 1625 1602
rect 1596 1599 1597 1600
rect 1591 1598 1597 1599
rect 1666 1599 1667 1603
rect 1671 1602 1672 1603
rect 2623 1603 2624 1607
rect 2628 1606 2629 1607
rect 2951 1607 2952 1608
rect 2956 1607 2957 1611
rect 3574 1608 3575 1612
rect 3579 1608 3580 1612
rect 2951 1606 2957 1607
rect 3098 1607 3104 1608
rect 2628 1604 2721 1606
rect 2628 1603 2629 1604
rect 2623 1602 2629 1603
rect 3098 1603 3099 1607
rect 3103 1606 3104 1607
rect 3271 1607 3277 1608
rect 3574 1607 3580 1608
rect 3103 1604 3209 1606
rect 3103 1603 3104 1604
rect 3098 1602 3104 1603
rect 3271 1603 3272 1607
rect 3276 1606 3277 1607
rect 3276 1604 3369 1606
rect 3276 1603 3277 1604
rect 3271 1602 3277 1603
rect 1671 1600 1753 1602
rect 1822 1600 1828 1601
rect 1671 1599 1672 1600
rect 1666 1598 1672 1599
rect 110 1595 116 1596
rect 1822 1596 1823 1600
rect 1827 1596 1828 1600
rect 1822 1595 1828 1596
rect 1862 1595 1868 1596
rect 1862 1591 1863 1595
rect 1867 1591 1868 1595
rect 3103 1595 3109 1596
rect 3103 1594 3104 1595
rect 3081 1592 3104 1594
rect 1862 1590 1868 1591
rect 3103 1591 3104 1592
rect 3108 1591 3109 1595
rect 3103 1590 3109 1591
rect 3470 1595 3476 1596
rect 3470 1591 3471 1595
rect 3475 1594 3476 1595
rect 3574 1595 3580 1596
rect 3475 1592 3497 1594
rect 3475 1591 3476 1592
rect 3470 1590 3476 1591
rect 3574 1591 3575 1595
rect 3579 1591 3580 1595
rect 3574 1590 3580 1591
rect 142 1587 148 1588
rect 142 1583 143 1587
rect 147 1583 148 1587
rect 142 1582 148 1583
rect 278 1587 284 1588
rect 278 1583 279 1587
rect 283 1583 284 1587
rect 278 1582 284 1583
rect 454 1587 460 1588
rect 454 1583 455 1587
rect 459 1583 460 1587
rect 454 1582 460 1583
rect 638 1587 644 1588
rect 638 1583 639 1587
rect 643 1583 644 1587
rect 638 1582 644 1583
rect 822 1587 828 1588
rect 822 1583 823 1587
rect 827 1583 828 1587
rect 822 1582 828 1583
rect 998 1587 1004 1588
rect 998 1583 999 1587
rect 1003 1583 1004 1587
rect 998 1582 1004 1583
rect 1158 1587 1164 1588
rect 1158 1583 1159 1587
rect 1163 1583 1164 1587
rect 1158 1582 1164 1583
rect 1310 1587 1316 1588
rect 1310 1583 1311 1587
rect 1315 1583 1316 1587
rect 1310 1582 1316 1583
rect 1462 1587 1468 1588
rect 1462 1583 1463 1587
rect 1467 1583 1468 1587
rect 1462 1582 1468 1583
rect 1606 1587 1612 1588
rect 1606 1583 1607 1587
rect 1611 1583 1612 1587
rect 1606 1582 1612 1583
rect 1734 1587 1740 1588
rect 1734 1583 1735 1587
rect 1739 1583 1740 1587
rect 1734 1582 1740 1583
rect 2142 1585 2148 1586
rect 2142 1581 2143 1585
rect 2147 1581 2148 1585
rect 2142 1580 2148 1581
rect 2334 1585 2340 1586
rect 2334 1581 2335 1585
rect 2339 1581 2340 1585
rect 2334 1580 2340 1581
rect 2518 1585 2524 1586
rect 2518 1581 2519 1585
rect 2523 1581 2524 1585
rect 2518 1580 2524 1581
rect 2694 1585 2700 1586
rect 2694 1581 2695 1585
rect 2699 1581 2700 1585
rect 2694 1580 2700 1581
rect 2862 1585 2868 1586
rect 2862 1581 2863 1585
rect 2867 1581 2868 1585
rect 2862 1580 2868 1581
rect 3022 1585 3028 1586
rect 3022 1581 3023 1585
rect 3027 1581 3028 1585
rect 3022 1580 3028 1581
rect 3182 1585 3188 1586
rect 3182 1581 3183 1585
rect 3187 1581 3188 1585
rect 3182 1580 3188 1581
rect 3342 1585 3348 1586
rect 3342 1581 3343 1585
rect 3347 1581 3348 1585
rect 3342 1580 3348 1581
rect 3478 1585 3484 1586
rect 3478 1581 3479 1585
rect 3483 1581 3484 1585
rect 3478 1580 3484 1581
rect 134 1575 141 1576
rect 134 1571 135 1575
rect 140 1571 141 1575
rect 134 1570 141 1571
rect 271 1575 277 1576
rect 271 1571 272 1575
rect 276 1574 277 1575
rect 286 1575 292 1576
rect 286 1574 287 1575
rect 276 1572 287 1574
rect 276 1571 277 1572
rect 271 1570 277 1571
rect 286 1571 287 1572
rect 291 1571 292 1575
rect 286 1570 292 1571
rect 439 1575 445 1576
rect 439 1571 440 1575
rect 444 1574 445 1575
rect 447 1575 453 1576
rect 447 1574 448 1575
rect 444 1572 448 1574
rect 444 1571 445 1572
rect 439 1570 445 1571
rect 447 1571 448 1572
rect 452 1571 453 1575
rect 447 1570 453 1571
rect 623 1575 629 1576
rect 623 1571 624 1575
rect 628 1574 629 1575
rect 631 1575 637 1576
rect 631 1574 632 1575
rect 628 1572 632 1574
rect 628 1571 629 1572
rect 623 1570 629 1571
rect 631 1571 632 1572
rect 636 1571 637 1575
rect 631 1570 637 1571
rect 807 1575 813 1576
rect 807 1571 808 1575
rect 812 1574 813 1575
rect 815 1575 821 1576
rect 815 1574 816 1575
rect 812 1572 816 1574
rect 812 1571 813 1572
rect 807 1570 813 1571
rect 815 1571 816 1572
rect 820 1571 821 1575
rect 815 1570 821 1571
rect 991 1575 997 1576
rect 991 1571 992 1575
rect 996 1574 997 1575
rect 1026 1575 1032 1576
rect 1026 1574 1027 1575
rect 996 1572 1027 1574
rect 996 1571 997 1572
rect 991 1570 997 1571
rect 1026 1571 1027 1572
rect 1031 1571 1032 1575
rect 1026 1570 1032 1571
rect 1151 1575 1157 1576
rect 1151 1571 1152 1575
rect 1156 1574 1157 1575
rect 1166 1575 1172 1576
rect 1166 1574 1167 1575
rect 1156 1572 1167 1574
rect 1156 1571 1157 1572
rect 1151 1570 1157 1571
rect 1166 1571 1167 1572
rect 1171 1571 1172 1575
rect 1166 1570 1172 1571
rect 1295 1575 1301 1576
rect 1295 1571 1296 1575
rect 1300 1574 1301 1575
rect 1303 1575 1309 1576
rect 1303 1574 1304 1575
rect 1300 1572 1304 1574
rect 1300 1571 1301 1572
rect 1295 1570 1301 1571
rect 1303 1571 1304 1572
rect 1308 1571 1309 1575
rect 1303 1570 1309 1571
rect 1455 1575 1461 1576
rect 1455 1571 1456 1575
rect 1460 1574 1461 1575
rect 1591 1575 1597 1576
rect 1591 1574 1592 1575
rect 1460 1572 1592 1574
rect 1460 1571 1461 1572
rect 1455 1570 1461 1571
rect 1591 1571 1592 1572
rect 1596 1571 1597 1575
rect 1591 1570 1597 1571
rect 1599 1575 1605 1576
rect 1599 1571 1600 1575
rect 1604 1574 1605 1575
rect 1666 1575 1672 1576
rect 1666 1574 1667 1575
rect 1604 1572 1667 1574
rect 1604 1571 1605 1572
rect 1599 1570 1605 1571
rect 1666 1571 1667 1572
rect 1671 1571 1672 1575
rect 1666 1570 1672 1571
rect 1719 1575 1725 1576
rect 1719 1571 1720 1575
rect 1724 1574 1725 1575
rect 1727 1575 1733 1576
rect 1727 1574 1728 1575
rect 1724 1572 1728 1574
rect 1724 1571 1725 1572
rect 1719 1570 1725 1571
rect 1727 1571 1728 1572
rect 1732 1571 1733 1575
rect 1727 1570 1733 1571
rect 2102 1571 2108 1572
rect 2102 1567 2103 1571
rect 2107 1570 2108 1571
rect 2107 1568 2394 1570
rect 2107 1567 2108 1568
rect 2102 1566 2108 1567
rect 135 1563 141 1564
rect 135 1559 136 1563
rect 140 1562 141 1563
rect 210 1563 216 1564
rect 210 1562 211 1563
rect 140 1560 211 1562
rect 140 1559 141 1560
rect 135 1558 141 1559
rect 210 1559 211 1560
rect 215 1559 216 1563
rect 210 1558 216 1559
rect 250 1563 256 1564
rect 250 1559 251 1563
rect 255 1562 256 1563
rect 263 1563 269 1564
rect 263 1562 264 1563
rect 255 1560 264 1562
rect 255 1559 256 1560
rect 250 1558 256 1559
rect 263 1559 264 1560
rect 268 1559 269 1563
rect 263 1558 269 1559
rect 423 1563 429 1564
rect 423 1559 424 1563
rect 428 1562 429 1563
rect 514 1563 520 1564
rect 514 1562 515 1563
rect 428 1560 515 1562
rect 428 1559 429 1560
rect 423 1558 429 1559
rect 514 1559 515 1560
rect 519 1559 520 1563
rect 514 1558 520 1559
rect 591 1563 597 1564
rect 591 1559 592 1563
rect 596 1562 597 1563
rect 666 1563 672 1564
rect 666 1562 667 1563
rect 596 1560 667 1562
rect 596 1559 597 1560
rect 591 1558 597 1559
rect 666 1559 667 1560
rect 671 1559 672 1563
rect 666 1558 672 1559
rect 759 1563 765 1564
rect 759 1559 760 1563
rect 764 1562 765 1563
rect 767 1563 773 1564
rect 767 1562 768 1563
rect 764 1560 768 1562
rect 764 1559 765 1560
rect 759 1558 765 1559
rect 767 1559 768 1560
rect 772 1559 773 1563
rect 767 1558 773 1559
rect 927 1563 933 1564
rect 927 1559 928 1563
rect 932 1562 933 1563
rect 942 1563 948 1564
rect 942 1562 943 1563
rect 932 1560 943 1562
rect 932 1559 933 1560
rect 927 1558 933 1559
rect 942 1559 943 1560
rect 947 1559 948 1563
rect 942 1558 948 1559
rect 1018 1563 1024 1564
rect 1018 1559 1019 1563
rect 1023 1562 1024 1563
rect 1095 1563 1101 1564
rect 1095 1562 1096 1563
rect 1023 1560 1096 1562
rect 1023 1559 1024 1560
rect 1018 1558 1024 1559
rect 1095 1559 1096 1560
rect 1100 1559 1101 1563
rect 1095 1558 1101 1559
rect 1255 1563 1261 1564
rect 1255 1559 1256 1563
rect 1260 1562 1261 1563
rect 1263 1563 1269 1564
rect 1263 1562 1264 1563
rect 1260 1560 1264 1562
rect 1260 1559 1261 1560
rect 1255 1558 1261 1559
rect 1263 1559 1264 1560
rect 1268 1559 1269 1563
rect 1263 1558 1269 1559
rect 1342 1563 1348 1564
rect 1342 1559 1343 1563
rect 1347 1562 1348 1563
rect 1415 1563 1421 1564
rect 1415 1562 1416 1563
rect 1347 1560 1416 1562
rect 1347 1559 1348 1560
rect 1342 1558 1348 1559
rect 1415 1559 1416 1560
rect 1420 1559 1421 1563
rect 1415 1558 1421 1559
rect 1582 1563 1589 1564
rect 1582 1559 1583 1563
rect 1588 1559 1589 1563
rect 1582 1558 1589 1559
rect 1662 1563 1668 1564
rect 1662 1559 1663 1563
rect 1667 1562 1668 1563
rect 1727 1563 1733 1564
rect 1727 1562 1728 1563
rect 1667 1560 1728 1562
rect 1667 1559 1668 1560
rect 1662 1558 1668 1559
rect 1727 1559 1728 1560
rect 1732 1559 1733 1563
rect 1727 1558 1733 1559
rect 2086 1563 2092 1564
rect 2086 1559 2087 1563
rect 2091 1559 2092 1563
rect 2086 1558 2092 1559
rect 2278 1563 2284 1564
rect 2278 1559 2279 1563
rect 2283 1559 2284 1563
rect 2278 1558 2284 1559
rect 2158 1555 2164 1556
rect 2158 1554 2159 1555
rect 142 1553 148 1554
rect 142 1549 143 1553
rect 147 1549 148 1553
rect 142 1548 148 1549
rect 270 1553 276 1554
rect 270 1549 271 1553
rect 275 1549 276 1553
rect 270 1548 276 1549
rect 430 1553 436 1554
rect 430 1549 431 1553
rect 435 1549 436 1553
rect 430 1548 436 1549
rect 598 1553 604 1554
rect 598 1549 599 1553
rect 603 1549 604 1553
rect 598 1548 604 1549
rect 766 1553 772 1554
rect 766 1549 767 1553
rect 771 1549 772 1553
rect 766 1548 772 1549
rect 934 1553 940 1554
rect 934 1549 935 1553
rect 939 1549 940 1553
rect 934 1548 940 1549
rect 1102 1553 1108 1554
rect 1102 1549 1103 1553
rect 1107 1549 1108 1553
rect 1102 1548 1108 1549
rect 1262 1553 1268 1554
rect 1262 1549 1263 1553
rect 1267 1549 1268 1553
rect 1262 1548 1268 1549
rect 1422 1553 1428 1554
rect 1422 1549 1423 1553
rect 1427 1549 1428 1553
rect 1422 1548 1428 1549
rect 1590 1553 1596 1554
rect 1590 1549 1591 1553
rect 1595 1549 1596 1553
rect 1590 1548 1596 1549
rect 1734 1553 1740 1554
rect 1734 1549 1735 1553
rect 1739 1549 1740 1553
rect 1734 1548 1740 1549
rect 1862 1553 1868 1554
rect 1862 1549 1863 1553
rect 1867 1549 1868 1553
rect 2145 1552 2159 1554
rect 2158 1551 2159 1552
rect 2163 1551 2164 1555
rect 2392 1554 2394 1568
rect 2454 1563 2460 1564
rect 2454 1559 2455 1563
rect 2459 1559 2460 1563
rect 2454 1558 2460 1559
rect 2622 1563 2628 1564
rect 2622 1559 2623 1563
rect 2627 1559 2628 1563
rect 2622 1558 2628 1559
rect 2790 1563 2796 1564
rect 2790 1559 2791 1563
rect 2795 1559 2796 1563
rect 2790 1558 2796 1559
rect 2950 1563 2956 1564
rect 2950 1559 2951 1563
rect 2955 1559 2956 1563
rect 2950 1558 2956 1559
rect 3110 1563 3116 1564
rect 3110 1559 3111 1563
rect 3115 1559 3116 1563
rect 3110 1558 3116 1559
rect 3270 1563 3276 1564
rect 3270 1559 3271 1563
rect 3275 1559 3276 1563
rect 3270 1558 3276 1559
rect 3430 1563 3436 1564
rect 3430 1559 3431 1563
rect 3435 1559 3436 1563
rect 3430 1558 3436 1559
rect 3214 1555 3220 1556
rect 2392 1552 2473 1554
rect 2158 1550 2164 1551
rect 3214 1551 3215 1555
rect 3219 1554 3220 1555
rect 3498 1555 3504 1556
rect 3498 1554 3499 1555
rect 3219 1552 3289 1554
rect 3489 1552 3499 1554
rect 3219 1551 3220 1552
rect 3214 1550 3220 1551
rect 3498 1551 3499 1552
rect 3503 1551 3504 1555
rect 3498 1550 3504 1551
rect 3574 1553 3580 1554
rect 1862 1548 1868 1549
rect 3574 1549 3575 1553
rect 3579 1549 3580 1553
rect 3574 1548 3580 1549
rect 110 1540 116 1541
rect 1822 1540 1828 1541
rect 110 1536 111 1540
rect 115 1536 116 1540
rect 1018 1539 1024 1540
rect 1018 1538 1019 1539
rect 989 1536 1019 1538
rect 110 1535 116 1536
rect 134 1535 140 1536
rect 134 1531 135 1535
rect 139 1534 140 1535
rect 210 1535 216 1536
rect 139 1532 161 1534
rect 139 1531 140 1532
rect 134 1530 140 1531
rect 210 1531 211 1535
rect 215 1534 216 1535
rect 514 1535 520 1536
rect 215 1532 289 1534
rect 215 1531 216 1532
rect 210 1530 216 1531
rect 514 1531 515 1535
rect 519 1534 520 1535
rect 666 1535 672 1536
rect 519 1532 617 1534
rect 519 1531 520 1532
rect 514 1530 520 1531
rect 666 1531 667 1535
rect 671 1534 672 1535
rect 1018 1535 1019 1536
rect 1023 1535 1024 1539
rect 1342 1539 1348 1540
rect 1342 1538 1343 1539
rect 1317 1536 1343 1538
rect 1018 1534 1024 1535
rect 1026 1535 1032 1536
rect 671 1532 785 1534
rect 671 1531 672 1532
rect 666 1530 672 1531
rect 1026 1531 1027 1535
rect 1031 1534 1032 1535
rect 1342 1535 1343 1536
rect 1347 1535 1348 1539
rect 1662 1539 1668 1540
rect 1662 1538 1663 1539
rect 1645 1536 1663 1538
rect 1342 1534 1348 1535
rect 1662 1535 1663 1536
rect 1667 1535 1668 1539
rect 1822 1536 1823 1540
rect 1827 1536 1828 1540
rect 2447 1539 2453 1540
rect 2447 1538 2448 1539
rect 1822 1535 1828 1536
rect 1862 1536 1868 1537
rect 2341 1536 2448 1538
rect 1662 1534 1668 1535
rect 1031 1532 1121 1534
rect 1862 1532 1863 1536
rect 1867 1532 1868 1536
rect 2447 1535 2448 1536
rect 2452 1535 2453 1539
rect 2783 1539 2789 1540
rect 2783 1538 2784 1539
rect 2685 1536 2784 1538
rect 2447 1534 2453 1535
rect 2783 1535 2784 1536
rect 2788 1535 2789 1539
rect 2943 1539 2949 1540
rect 2943 1538 2944 1539
rect 2853 1536 2944 1538
rect 2783 1534 2789 1535
rect 2943 1535 2944 1536
rect 2948 1535 2949 1539
rect 3078 1539 3084 1540
rect 3078 1538 3079 1539
rect 3013 1536 3079 1538
rect 2943 1534 2949 1535
rect 3078 1535 3079 1536
rect 3083 1535 3084 1539
rect 3263 1539 3269 1540
rect 3263 1538 3264 1539
rect 3173 1536 3264 1538
rect 3078 1534 3084 1535
rect 3263 1535 3264 1536
rect 3268 1535 3269 1539
rect 3263 1534 3269 1535
rect 3574 1536 3580 1537
rect 1031 1531 1032 1532
rect 1862 1531 1868 1532
rect 3574 1532 3575 1536
rect 3579 1532 3580 1536
rect 3574 1531 3580 1532
rect 1026 1530 1032 1531
rect 110 1523 116 1524
rect 110 1519 111 1523
rect 115 1519 116 1523
rect 110 1518 116 1519
rect 350 1523 356 1524
rect 350 1519 351 1523
rect 355 1522 356 1523
rect 1390 1523 1396 1524
rect 355 1520 441 1522
rect 355 1519 356 1520
rect 350 1518 356 1519
rect 1390 1519 1391 1523
rect 1395 1522 1396 1523
rect 1814 1523 1820 1524
rect 1814 1522 1815 1523
rect 1395 1520 1433 1522
rect 1785 1520 1815 1522
rect 1395 1519 1396 1520
rect 1390 1518 1396 1519
rect 1814 1519 1815 1520
rect 1819 1519 1820 1523
rect 1814 1518 1820 1519
rect 1822 1523 1828 1524
rect 1822 1519 1823 1523
rect 1827 1519 1828 1523
rect 1822 1518 1828 1519
rect 2094 1523 2100 1524
rect 2094 1519 2095 1523
rect 2099 1519 2100 1523
rect 2094 1518 2100 1519
rect 2286 1523 2292 1524
rect 2286 1519 2287 1523
rect 2291 1519 2292 1523
rect 2286 1518 2292 1519
rect 2462 1523 2468 1524
rect 2462 1519 2463 1523
rect 2467 1519 2468 1523
rect 2462 1518 2468 1519
rect 2630 1523 2636 1524
rect 2630 1519 2631 1523
rect 2635 1519 2636 1523
rect 2630 1518 2636 1519
rect 2798 1523 2804 1524
rect 2798 1519 2799 1523
rect 2803 1519 2804 1523
rect 2798 1518 2804 1519
rect 2958 1523 2964 1524
rect 2958 1519 2959 1523
rect 2963 1519 2964 1523
rect 2958 1518 2964 1519
rect 3118 1523 3124 1524
rect 3118 1519 3119 1523
rect 3123 1519 3124 1523
rect 3118 1518 3124 1519
rect 3278 1523 3284 1524
rect 3278 1519 3279 1523
rect 3283 1519 3284 1523
rect 3278 1518 3284 1519
rect 3438 1523 3444 1524
rect 3438 1519 3439 1523
rect 3443 1519 3444 1523
rect 3438 1518 3444 1519
rect 134 1513 140 1514
rect 134 1509 135 1513
rect 139 1509 140 1513
rect 134 1508 140 1509
rect 262 1513 268 1514
rect 262 1509 263 1513
rect 267 1509 268 1513
rect 262 1508 268 1509
rect 422 1513 428 1514
rect 422 1509 423 1513
rect 427 1509 428 1513
rect 422 1508 428 1509
rect 590 1513 596 1514
rect 590 1509 591 1513
rect 595 1509 596 1513
rect 590 1508 596 1509
rect 758 1513 764 1514
rect 758 1509 759 1513
rect 763 1509 764 1513
rect 758 1508 764 1509
rect 926 1513 932 1514
rect 926 1509 927 1513
rect 931 1509 932 1513
rect 926 1508 932 1509
rect 1094 1513 1100 1514
rect 1094 1509 1095 1513
rect 1099 1509 1100 1513
rect 1094 1508 1100 1509
rect 1254 1513 1260 1514
rect 1254 1509 1255 1513
rect 1259 1509 1260 1513
rect 1254 1508 1260 1509
rect 1414 1513 1420 1514
rect 1414 1509 1415 1513
rect 1419 1509 1420 1513
rect 1414 1508 1420 1509
rect 1582 1513 1588 1514
rect 1582 1509 1583 1513
rect 1587 1509 1588 1513
rect 1582 1508 1588 1509
rect 1726 1513 1732 1514
rect 1726 1509 1727 1513
rect 1731 1509 1732 1513
rect 1726 1508 1732 1509
rect 2087 1511 2093 1512
rect 2087 1507 2088 1511
rect 2092 1510 2093 1511
rect 2102 1511 2108 1512
rect 2102 1510 2103 1511
rect 2092 1508 2103 1510
rect 2092 1507 2093 1508
rect 2087 1506 2093 1507
rect 2102 1507 2103 1508
rect 2107 1507 2108 1511
rect 2102 1506 2108 1507
rect 2178 1511 2184 1512
rect 2178 1507 2179 1511
rect 2183 1510 2184 1511
rect 2279 1511 2285 1512
rect 2279 1510 2280 1511
rect 2183 1508 2280 1510
rect 2183 1507 2184 1508
rect 2178 1506 2184 1507
rect 2279 1507 2280 1508
rect 2284 1507 2285 1511
rect 2279 1506 2285 1507
rect 2447 1511 2453 1512
rect 2447 1507 2448 1511
rect 2452 1510 2453 1511
rect 2455 1511 2461 1512
rect 2455 1510 2456 1511
rect 2452 1508 2456 1510
rect 2452 1507 2453 1508
rect 2447 1506 2453 1507
rect 2455 1507 2456 1508
rect 2460 1507 2461 1511
rect 2455 1506 2461 1507
rect 2623 1511 2629 1512
rect 2623 1507 2624 1511
rect 2628 1510 2629 1511
rect 2638 1511 2644 1512
rect 2638 1510 2639 1511
rect 2628 1508 2639 1510
rect 2628 1507 2629 1508
rect 2623 1506 2629 1507
rect 2638 1507 2639 1508
rect 2643 1507 2644 1511
rect 2638 1506 2644 1507
rect 2783 1511 2789 1512
rect 2783 1507 2784 1511
rect 2788 1510 2789 1511
rect 2791 1511 2797 1512
rect 2791 1510 2792 1511
rect 2788 1508 2792 1510
rect 2788 1507 2789 1508
rect 2783 1506 2789 1507
rect 2791 1507 2792 1508
rect 2796 1507 2797 1511
rect 2791 1506 2797 1507
rect 2943 1511 2949 1512
rect 2943 1507 2944 1511
rect 2948 1510 2949 1511
rect 2951 1511 2957 1512
rect 2951 1510 2952 1511
rect 2948 1508 2952 1510
rect 2948 1507 2949 1508
rect 2943 1506 2949 1507
rect 2951 1507 2952 1508
rect 2956 1507 2957 1511
rect 2951 1506 2957 1507
rect 3103 1511 3109 1512
rect 3103 1507 3104 1511
rect 3108 1510 3109 1511
rect 3111 1511 3117 1512
rect 3111 1510 3112 1511
rect 3108 1508 3112 1510
rect 3108 1507 3109 1508
rect 3103 1506 3109 1507
rect 3111 1507 3112 1508
rect 3116 1507 3117 1511
rect 3111 1506 3117 1507
rect 3263 1511 3269 1512
rect 3263 1507 3264 1511
rect 3268 1510 3269 1511
rect 3271 1511 3277 1512
rect 3271 1510 3272 1511
rect 3268 1508 3272 1510
rect 3268 1507 3269 1508
rect 3263 1506 3269 1507
rect 3271 1507 3272 1508
rect 3276 1507 3277 1511
rect 3271 1506 3277 1507
rect 3367 1511 3373 1512
rect 3367 1507 3368 1511
rect 3372 1510 3373 1511
rect 3431 1511 3437 1512
rect 3431 1510 3432 1511
rect 3372 1508 3432 1510
rect 3372 1507 3373 1508
rect 3367 1506 3373 1507
rect 3431 1507 3432 1508
rect 3436 1507 3437 1511
rect 3431 1506 3437 1507
rect 2778 1499 2784 1500
rect 2778 1498 2779 1499
rect 2608 1496 2779 1498
rect 1814 1491 1820 1492
rect 182 1487 188 1488
rect 182 1483 183 1487
rect 187 1483 188 1487
rect 182 1482 188 1483
rect 326 1487 332 1488
rect 326 1483 327 1487
rect 331 1483 332 1487
rect 326 1482 332 1483
rect 470 1487 476 1488
rect 470 1483 471 1487
rect 475 1483 476 1487
rect 470 1482 476 1483
rect 606 1487 612 1488
rect 606 1483 607 1487
rect 611 1483 612 1487
rect 606 1482 612 1483
rect 742 1487 748 1488
rect 742 1483 743 1487
rect 747 1483 748 1487
rect 742 1482 748 1483
rect 870 1487 876 1488
rect 870 1483 871 1487
rect 875 1483 876 1487
rect 870 1482 876 1483
rect 990 1487 996 1488
rect 990 1483 991 1487
rect 995 1483 996 1487
rect 990 1482 996 1483
rect 1118 1487 1124 1488
rect 1118 1483 1119 1487
rect 1123 1483 1124 1487
rect 1118 1482 1124 1483
rect 1246 1487 1252 1488
rect 1246 1483 1247 1487
rect 1251 1483 1252 1487
rect 1246 1482 1252 1483
rect 1374 1487 1380 1488
rect 1374 1483 1375 1487
rect 1379 1483 1380 1487
rect 1814 1487 1815 1491
rect 1819 1490 1820 1491
rect 1887 1491 1893 1492
rect 1887 1490 1888 1491
rect 1819 1488 1888 1490
rect 1819 1487 1820 1488
rect 1814 1486 1820 1487
rect 1887 1487 1888 1488
rect 1892 1487 1893 1491
rect 1887 1486 1893 1487
rect 1959 1491 1965 1492
rect 1959 1487 1960 1491
rect 1964 1490 1965 1491
rect 1983 1491 1989 1492
rect 1983 1490 1984 1491
rect 1964 1488 1984 1490
rect 1964 1487 1965 1488
rect 1959 1486 1965 1487
rect 1983 1487 1984 1488
rect 1988 1487 1989 1491
rect 1983 1486 1989 1487
rect 2111 1491 2117 1492
rect 2111 1487 2112 1491
rect 2116 1490 2117 1491
rect 2186 1491 2192 1492
rect 2186 1490 2187 1491
rect 2116 1488 2187 1490
rect 2116 1487 2117 1488
rect 2111 1486 2117 1487
rect 2186 1487 2187 1488
rect 2191 1487 2192 1491
rect 2186 1486 2192 1487
rect 2239 1491 2245 1492
rect 2239 1487 2240 1491
rect 2244 1490 2245 1491
rect 2335 1491 2341 1492
rect 2335 1490 2336 1491
rect 2244 1488 2336 1490
rect 2244 1487 2245 1488
rect 2239 1486 2245 1487
rect 2335 1487 2336 1488
rect 2340 1487 2341 1491
rect 2335 1486 2341 1487
rect 2375 1491 2381 1492
rect 2375 1487 2376 1491
rect 2380 1490 2381 1491
rect 2390 1491 2396 1492
rect 2390 1490 2391 1491
rect 2380 1488 2391 1490
rect 2380 1487 2381 1488
rect 2375 1486 2381 1487
rect 2390 1487 2391 1488
rect 2395 1487 2396 1491
rect 2390 1486 2396 1487
rect 2527 1491 2533 1492
rect 2527 1487 2528 1491
rect 2532 1490 2533 1491
rect 2608 1490 2610 1496
rect 2778 1495 2779 1496
rect 2783 1495 2784 1499
rect 3218 1499 3224 1500
rect 3218 1498 3219 1499
rect 2778 1494 2784 1495
rect 3008 1496 3219 1498
rect 2532 1488 2610 1490
rect 2615 1491 2621 1492
rect 2532 1487 2533 1488
rect 2527 1486 2533 1487
rect 2615 1487 2616 1491
rect 2620 1490 2621 1491
rect 2695 1491 2701 1492
rect 2695 1490 2696 1491
rect 2620 1488 2696 1490
rect 2620 1487 2621 1488
rect 2615 1486 2621 1487
rect 2695 1487 2696 1488
rect 2700 1487 2701 1491
rect 2695 1486 2701 1487
rect 2879 1491 2885 1492
rect 2879 1487 2880 1491
rect 2884 1490 2885 1491
rect 3008 1490 3010 1496
rect 3218 1495 3219 1496
rect 3223 1495 3224 1499
rect 3218 1494 3224 1495
rect 2884 1488 3010 1490
rect 3078 1491 3085 1492
rect 2884 1487 2885 1488
rect 2879 1486 2885 1487
rect 3078 1487 3079 1491
rect 3084 1487 3085 1491
rect 3078 1486 3085 1487
rect 3191 1491 3197 1492
rect 3191 1487 3192 1491
rect 3196 1490 3197 1491
rect 3287 1491 3293 1492
rect 3287 1490 3288 1491
rect 3196 1488 3288 1490
rect 3196 1487 3197 1488
rect 3191 1486 3197 1487
rect 3287 1487 3288 1488
rect 3292 1487 3293 1491
rect 3287 1486 3293 1487
rect 3470 1491 3476 1492
rect 3470 1487 3471 1491
rect 3475 1490 3476 1491
rect 3479 1491 3485 1492
rect 3479 1490 3480 1491
rect 3475 1488 3480 1490
rect 3475 1487 3476 1488
rect 3470 1486 3476 1487
rect 3479 1487 3480 1488
rect 3484 1487 3485 1491
rect 3479 1486 3485 1487
rect 1374 1482 1380 1483
rect 1894 1481 1900 1482
rect 250 1479 256 1480
rect 250 1478 251 1479
rect 110 1477 116 1478
rect 110 1473 111 1477
rect 115 1473 116 1477
rect 241 1476 251 1478
rect 250 1475 251 1476
rect 255 1475 256 1479
rect 250 1474 256 1475
rect 703 1479 709 1480
rect 703 1475 704 1479
rect 708 1478 709 1479
rect 942 1479 948 1480
rect 942 1478 943 1479
rect 708 1476 761 1478
rect 929 1476 943 1478
rect 708 1475 709 1476
rect 703 1474 709 1475
rect 942 1475 943 1476
rect 947 1475 948 1479
rect 942 1474 948 1475
rect 1822 1477 1828 1478
rect 110 1472 116 1473
rect 1822 1473 1823 1477
rect 1827 1473 1828 1477
rect 1894 1477 1895 1481
rect 1899 1477 1900 1481
rect 1894 1476 1900 1477
rect 1990 1481 1996 1482
rect 1990 1477 1991 1481
rect 1995 1477 1996 1481
rect 1990 1476 1996 1477
rect 2118 1481 2124 1482
rect 2118 1477 2119 1481
rect 2123 1477 2124 1481
rect 2118 1476 2124 1477
rect 2246 1481 2252 1482
rect 2246 1477 2247 1481
rect 2251 1477 2252 1481
rect 2246 1476 2252 1477
rect 2382 1481 2388 1482
rect 2382 1477 2383 1481
rect 2387 1477 2388 1481
rect 2382 1476 2388 1477
rect 2534 1481 2540 1482
rect 2534 1477 2535 1481
rect 2539 1477 2540 1481
rect 2534 1476 2540 1477
rect 2702 1481 2708 1482
rect 2702 1477 2703 1481
rect 2707 1477 2708 1481
rect 2702 1476 2708 1477
rect 2886 1481 2892 1482
rect 2886 1477 2887 1481
rect 2891 1477 2892 1481
rect 2886 1476 2892 1477
rect 3086 1481 3092 1482
rect 3086 1477 3087 1481
rect 3091 1477 3092 1481
rect 3086 1476 3092 1477
rect 3294 1481 3300 1482
rect 3294 1477 3295 1481
rect 3299 1477 3300 1481
rect 3294 1476 3300 1477
rect 3486 1481 3492 1482
rect 3486 1477 3487 1481
rect 3491 1477 3492 1481
rect 3486 1476 3492 1477
rect 1822 1472 1828 1473
rect 1862 1468 1868 1469
rect 3574 1468 3580 1469
rect 1862 1464 1863 1468
rect 1867 1464 1868 1468
rect 1959 1467 1965 1468
rect 1959 1466 1960 1467
rect 1949 1464 1960 1466
rect 463 1463 469 1464
rect 463 1462 464 1463
rect 110 1460 116 1461
rect 389 1460 464 1462
rect 110 1456 111 1460
rect 115 1456 116 1460
rect 463 1459 464 1460
rect 468 1459 469 1463
rect 599 1463 605 1464
rect 599 1462 600 1463
rect 533 1460 600 1462
rect 463 1458 469 1459
rect 599 1459 600 1460
rect 604 1459 605 1463
rect 735 1463 741 1464
rect 735 1462 736 1463
rect 669 1460 736 1462
rect 599 1458 605 1459
rect 735 1459 736 1460
rect 740 1459 741 1463
rect 735 1458 741 1459
rect 938 1463 944 1464
rect 938 1459 939 1463
rect 943 1462 944 1463
rect 1058 1463 1064 1464
rect 943 1460 1017 1462
rect 943 1459 944 1460
rect 938 1458 944 1459
rect 1058 1459 1059 1463
rect 1063 1462 1064 1463
rect 1223 1463 1229 1464
rect 1063 1460 1145 1462
rect 1063 1459 1064 1460
rect 1058 1458 1064 1459
rect 1223 1459 1224 1463
rect 1228 1462 1229 1463
rect 1314 1463 1320 1464
rect 1862 1463 1868 1464
rect 1959 1463 1960 1464
rect 1964 1463 1965 1467
rect 2178 1467 2184 1468
rect 2178 1466 2179 1467
rect 2173 1464 2179 1466
rect 1228 1460 1273 1462
rect 1228 1459 1229 1460
rect 1223 1458 1229 1459
rect 1314 1459 1315 1463
rect 1319 1462 1320 1463
rect 1959 1462 1965 1463
rect 2178 1463 2179 1464
rect 2183 1463 2184 1467
rect 2615 1467 2621 1468
rect 2615 1466 2616 1467
rect 2589 1464 2616 1466
rect 2178 1462 2184 1463
rect 2186 1463 2192 1464
rect 1319 1460 1401 1462
rect 1822 1460 1828 1461
rect 1319 1459 1320 1460
rect 1314 1458 1320 1459
rect 110 1455 116 1456
rect 1822 1456 1823 1460
rect 1827 1456 1828 1460
rect 2186 1459 2187 1463
rect 2191 1462 2192 1463
rect 2335 1463 2341 1464
rect 2191 1460 2265 1462
rect 2191 1459 2192 1460
rect 2186 1458 2192 1459
rect 2335 1459 2336 1463
rect 2340 1462 2341 1463
rect 2615 1463 2616 1464
rect 2620 1463 2621 1467
rect 3191 1467 3197 1468
rect 3191 1466 3192 1467
rect 3141 1464 3192 1466
rect 2615 1462 2621 1463
rect 2778 1463 2784 1464
rect 2340 1460 2401 1462
rect 2340 1459 2341 1460
rect 2335 1458 2341 1459
rect 2778 1459 2779 1463
rect 2783 1462 2784 1463
rect 3191 1463 3192 1464
rect 3196 1463 3197 1467
rect 3574 1464 3575 1468
rect 3579 1464 3580 1468
rect 3191 1462 3197 1463
rect 3218 1463 3224 1464
rect 3574 1463 3580 1464
rect 2783 1460 2905 1462
rect 2783 1459 2784 1460
rect 2778 1458 2784 1459
rect 3218 1459 3219 1463
rect 3223 1462 3224 1463
rect 3223 1460 3313 1462
rect 3223 1459 3224 1460
rect 3218 1458 3224 1459
rect 1822 1455 1828 1456
rect 1862 1451 1868 1452
rect 190 1447 196 1448
rect 190 1443 191 1447
rect 195 1443 196 1447
rect 190 1442 196 1443
rect 334 1447 340 1448
rect 334 1443 335 1447
rect 339 1443 340 1447
rect 334 1442 340 1443
rect 478 1447 484 1448
rect 478 1443 479 1447
rect 483 1443 484 1447
rect 478 1442 484 1443
rect 614 1447 620 1448
rect 614 1443 615 1447
rect 619 1443 620 1447
rect 614 1442 620 1443
rect 750 1447 756 1448
rect 750 1443 751 1447
rect 755 1443 756 1447
rect 750 1442 756 1443
rect 878 1447 884 1448
rect 878 1443 879 1447
rect 883 1443 884 1447
rect 878 1442 884 1443
rect 998 1447 1004 1448
rect 998 1443 999 1447
rect 1003 1443 1004 1447
rect 998 1442 1004 1443
rect 1126 1447 1132 1448
rect 1126 1443 1127 1447
rect 1131 1443 1132 1447
rect 1126 1442 1132 1443
rect 1254 1447 1260 1448
rect 1254 1443 1255 1447
rect 1259 1443 1260 1447
rect 1254 1442 1260 1443
rect 1382 1447 1388 1448
rect 1382 1443 1383 1447
rect 1387 1443 1388 1447
rect 1862 1447 1863 1451
rect 1867 1447 1868 1451
rect 2063 1451 2069 1452
rect 2063 1450 2064 1451
rect 2041 1448 2064 1450
rect 1862 1446 1868 1447
rect 2063 1447 2064 1448
rect 2068 1447 2069 1451
rect 2799 1451 2805 1452
rect 2799 1450 2800 1451
rect 2753 1448 2800 1450
rect 2063 1446 2069 1447
rect 2799 1447 2800 1448
rect 2804 1447 2805 1451
rect 2799 1446 2805 1447
rect 3471 1451 3477 1452
rect 3471 1447 3472 1451
rect 3476 1450 3477 1451
rect 3574 1451 3580 1452
rect 3476 1448 3497 1450
rect 3476 1447 3477 1448
rect 3471 1446 3477 1447
rect 3574 1447 3575 1451
rect 3579 1447 3580 1451
rect 3574 1446 3580 1447
rect 1382 1442 1388 1443
rect 1886 1441 1892 1442
rect 1886 1437 1887 1441
rect 1891 1437 1892 1441
rect 1886 1436 1892 1437
rect 1982 1441 1988 1442
rect 1982 1437 1983 1441
rect 1987 1437 1988 1441
rect 1982 1436 1988 1437
rect 2110 1441 2116 1442
rect 2110 1437 2111 1441
rect 2115 1437 2116 1441
rect 2110 1436 2116 1437
rect 2238 1441 2244 1442
rect 2238 1437 2239 1441
rect 2243 1437 2244 1441
rect 2238 1436 2244 1437
rect 2374 1441 2380 1442
rect 2374 1437 2375 1441
rect 2379 1437 2380 1441
rect 2374 1436 2380 1437
rect 2526 1441 2532 1442
rect 2526 1437 2527 1441
rect 2531 1437 2532 1441
rect 2526 1436 2532 1437
rect 2694 1441 2700 1442
rect 2694 1437 2695 1441
rect 2699 1437 2700 1441
rect 2694 1436 2700 1437
rect 2878 1441 2884 1442
rect 2878 1437 2879 1441
rect 2883 1437 2884 1441
rect 2878 1436 2884 1437
rect 3078 1441 3084 1442
rect 3078 1437 3079 1441
rect 3083 1437 3084 1441
rect 3078 1436 3084 1437
rect 3286 1441 3292 1442
rect 3286 1437 3287 1441
rect 3291 1437 3292 1441
rect 3286 1436 3292 1437
rect 3478 1441 3484 1442
rect 3478 1437 3479 1441
rect 3483 1437 3484 1441
rect 3478 1436 3484 1437
rect 182 1435 189 1436
rect 182 1431 183 1435
rect 188 1431 189 1435
rect 182 1430 189 1431
rect 327 1435 333 1436
rect 327 1431 328 1435
rect 332 1434 333 1435
rect 350 1435 356 1436
rect 350 1434 351 1435
rect 332 1432 351 1434
rect 332 1431 333 1432
rect 327 1430 333 1431
rect 350 1431 351 1432
rect 355 1431 356 1435
rect 350 1430 356 1431
rect 463 1435 469 1436
rect 463 1431 464 1435
rect 468 1434 469 1435
rect 471 1435 477 1436
rect 471 1434 472 1435
rect 468 1432 472 1434
rect 468 1431 469 1432
rect 463 1430 469 1431
rect 471 1431 472 1432
rect 476 1431 477 1435
rect 471 1430 477 1431
rect 599 1435 605 1436
rect 599 1431 600 1435
rect 604 1434 605 1435
rect 607 1435 613 1436
rect 607 1434 608 1435
rect 604 1432 608 1434
rect 604 1431 605 1432
rect 599 1430 605 1431
rect 607 1431 608 1432
rect 612 1431 613 1435
rect 607 1430 613 1431
rect 735 1435 741 1436
rect 735 1431 736 1435
rect 740 1434 741 1435
rect 743 1435 749 1436
rect 743 1434 744 1435
rect 740 1432 744 1434
rect 740 1431 741 1432
rect 735 1430 741 1431
rect 743 1431 744 1432
rect 748 1431 749 1435
rect 743 1430 749 1431
rect 871 1435 877 1436
rect 871 1431 872 1435
rect 876 1434 877 1435
rect 938 1435 944 1436
rect 938 1434 939 1435
rect 876 1432 939 1434
rect 876 1431 877 1432
rect 871 1430 877 1431
rect 938 1431 939 1432
rect 943 1431 944 1435
rect 938 1430 944 1431
rect 991 1435 997 1436
rect 991 1431 992 1435
rect 996 1434 997 1435
rect 1058 1435 1064 1436
rect 1058 1434 1059 1435
rect 996 1432 1059 1434
rect 996 1431 997 1432
rect 991 1430 997 1431
rect 1058 1431 1059 1432
rect 1063 1431 1064 1435
rect 1058 1430 1064 1431
rect 1110 1435 1116 1436
rect 1110 1431 1111 1435
rect 1115 1434 1116 1435
rect 1119 1435 1125 1436
rect 1119 1434 1120 1435
rect 1115 1432 1120 1434
rect 1115 1431 1116 1432
rect 1110 1430 1116 1431
rect 1119 1431 1120 1432
rect 1124 1431 1125 1435
rect 1119 1430 1125 1431
rect 1247 1435 1253 1436
rect 1247 1431 1248 1435
rect 1252 1434 1253 1435
rect 1314 1435 1320 1436
rect 1314 1434 1315 1435
rect 1252 1432 1315 1434
rect 1252 1431 1253 1432
rect 1247 1430 1253 1431
rect 1314 1431 1315 1432
rect 1319 1431 1320 1435
rect 1314 1430 1320 1431
rect 1375 1435 1381 1436
rect 1375 1431 1376 1435
rect 1380 1434 1381 1435
rect 1390 1435 1396 1436
rect 1390 1434 1391 1435
rect 1380 1432 1391 1434
rect 1380 1431 1381 1432
rect 1375 1430 1381 1431
rect 1390 1431 1391 1432
rect 1395 1431 1396 1435
rect 1390 1430 1396 1431
rect 658 1423 664 1424
rect 658 1422 659 1423
rect 520 1420 659 1422
rect 191 1415 197 1416
rect 191 1411 192 1415
rect 196 1414 197 1415
rect 270 1415 276 1416
rect 270 1414 271 1415
rect 196 1412 271 1414
rect 196 1411 197 1412
rect 191 1410 197 1411
rect 270 1411 271 1412
rect 275 1411 276 1415
rect 270 1410 276 1411
rect 298 1415 304 1416
rect 298 1411 299 1415
rect 303 1414 304 1415
rect 327 1415 333 1416
rect 327 1414 328 1415
rect 303 1412 328 1414
rect 303 1411 304 1412
rect 298 1410 304 1411
rect 327 1411 328 1412
rect 332 1411 333 1415
rect 327 1410 333 1411
rect 455 1415 461 1416
rect 455 1411 456 1415
rect 460 1414 461 1415
rect 520 1414 522 1420
rect 658 1419 659 1420
rect 663 1419 664 1423
rect 658 1418 664 1419
rect 460 1412 522 1414
rect 527 1415 533 1416
rect 460 1411 461 1412
rect 455 1410 461 1411
rect 527 1411 528 1415
rect 532 1414 533 1415
rect 575 1415 581 1416
rect 575 1414 576 1415
rect 532 1412 576 1414
rect 532 1411 533 1412
rect 527 1410 533 1411
rect 575 1411 576 1412
rect 580 1411 581 1415
rect 575 1410 581 1411
rect 695 1415 701 1416
rect 695 1411 696 1415
rect 700 1414 701 1415
rect 703 1415 709 1416
rect 703 1414 704 1415
rect 700 1412 704 1414
rect 700 1411 701 1412
rect 695 1410 701 1411
rect 703 1411 704 1412
rect 708 1411 709 1415
rect 703 1410 709 1411
rect 770 1415 776 1416
rect 770 1411 771 1415
rect 775 1414 776 1415
rect 807 1415 813 1416
rect 807 1414 808 1415
rect 775 1412 808 1414
rect 775 1411 776 1412
rect 770 1410 776 1411
rect 807 1411 808 1412
rect 812 1411 813 1415
rect 807 1410 813 1411
rect 879 1415 885 1416
rect 879 1411 880 1415
rect 884 1414 885 1415
rect 911 1415 917 1416
rect 911 1414 912 1415
rect 884 1412 912 1414
rect 884 1411 885 1412
rect 879 1410 885 1411
rect 911 1411 912 1412
rect 916 1411 917 1415
rect 911 1410 917 1411
rect 983 1415 989 1416
rect 983 1411 984 1415
rect 988 1414 989 1415
rect 1007 1415 1013 1416
rect 1007 1414 1008 1415
rect 988 1412 1008 1414
rect 988 1411 989 1412
rect 983 1410 989 1411
rect 1007 1411 1008 1412
rect 1012 1411 1013 1415
rect 1007 1410 1013 1411
rect 1079 1415 1085 1416
rect 1079 1411 1080 1415
rect 1084 1414 1085 1415
rect 1111 1415 1117 1416
rect 1111 1414 1112 1415
rect 1084 1412 1112 1414
rect 1084 1411 1085 1412
rect 1079 1410 1085 1411
rect 1111 1411 1112 1412
rect 1116 1411 1117 1415
rect 1111 1410 1117 1411
rect 1215 1415 1221 1416
rect 1215 1411 1216 1415
rect 1220 1414 1221 1415
rect 1223 1415 1229 1416
rect 1223 1414 1224 1415
rect 1220 1412 1224 1414
rect 1220 1411 1221 1412
rect 1215 1410 1221 1411
rect 1223 1411 1224 1412
rect 1228 1411 1229 1415
rect 1223 1410 1229 1411
rect 1287 1415 1293 1416
rect 1287 1411 1288 1415
rect 1292 1414 1293 1415
rect 1319 1415 1325 1416
rect 1319 1414 1320 1415
rect 1292 1412 1320 1414
rect 1292 1411 1293 1412
rect 1287 1410 1293 1411
rect 1319 1411 1320 1412
rect 1324 1411 1325 1415
rect 1319 1410 1325 1411
rect 1886 1415 1892 1416
rect 1886 1411 1887 1415
rect 1891 1411 1892 1415
rect 1886 1410 1892 1411
rect 1974 1415 1980 1416
rect 1974 1411 1975 1415
rect 1979 1411 1980 1415
rect 1974 1410 1980 1411
rect 2070 1415 2076 1416
rect 2070 1411 2071 1415
rect 2075 1411 2076 1415
rect 2070 1410 2076 1411
rect 2182 1415 2188 1416
rect 2182 1411 2183 1415
rect 2187 1411 2188 1415
rect 2182 1410 2188 1411
rect 2302 1415 2308 1416
rect 2302 1411 2303 1415
rect 2307 1411 2308 1415
rect 2302 1410 2308 1411
rect 2438 1415 2444 1416
rect 2438 1411 2439 1415
rect 2443 1411 2444 1415
rect 2438 1410 2444 1411
rect 2606 1415 2612 1416
rect 2606 1411 2607 1415
rect 2611 1411 2612 1415
rect 2606 1410 2612 1411
rect 2806 1415 2812 1416
rect 2806 1411 2807 1415
rect 2811 1411 2812 1415
rect 2806 1410 2812 1411
rect 3030 1415 3036 1416
rect 3030 1411 3031 1415
rect 3035 1411 3036 1415
rect 3030 1410 3036 1411
rect 3262 1415 3268 1416
rect 3262 1411 3263 1415
rect 3267 1411 3268 1415
rect 3262 1410 3268 1411
rect 3478 1415 3484 1416
rect 3478 1411 3479 1415
rect 3483 1411 3484 1415
rect 3478 1410 3484 1411
rect 2390 1407 2396 1408
rect 2390 1406 2391 1407
rect 198 1405 204 1406
rect 198 1401 199 1405
rect 203 1401 204 1405
rect 198 1400 204 1401
rect 334 1405 340 1406
rect 334 1401 335 1405
rect 339 1401 340 1405
rect 334 1400 340 1401
rect 462 1405 468 1406
rect 462 1401 463 1405
rect 467 1401 468 1405
rect 462 1400 468 1401
rect 582 1405 588 1406
rect 582 1401 583 1405
rect 587 1401 588 1405
rect 582 1400 588 1401
rect 702 1405 708 1406
rect 702 1401 703 1405
rect 707 1401 708 1405
rect 702 1400 708 1401
rect 814 1405 820 1406
rect 814 1401 815 1405
rect 819 1401 820 1405
rect 814 1400 820 1401
rect 918 1405 924 1406
rect 918 1401 919 1405
rect 923 1401 924 1405
rect 918 1400 924 1401
rect 1014 1405 1020 1406
rect 1014 1401 1015 1405
rect 1019 1401 1020 1405
rect 1014 1400 1020 1401
rect 1118 1405 1124 1406
rect 1118 1401 1119 1405
rect 1123 1401 1124 1405
rect 1118 1400 1124 1401
rect 1222 1405 1228 1406
rect 1222 1401 1223 1405
rect 1227 1401 1228 1405
rect 1222 1400 1228 1401
rect 1326 1405 1332 1406
rect 1326 1401 1327 1405
rect 1331 1401 1332 1405
rect 1326 1400 1332 1401
rect 1862 1405 1868 1406
rect 1862 1401 1863 1405
rect 1867 1401 1868 1405
rect 2361 1404 2391 1406
rect 2390 1403 2391 1404
rect 2395 1403 2396 1407
rect 2390 1402 2396 1403
rect 3210 1407 3216 1408
rect 3210 1403 3211 1407
rect 3215 1406 3216 1407
rect 3215 1404 3281 1406
rect 3574 1405 3580 1406
rect 3215 1403 3216 1404
rect 3210 1402 3216 1403
rect 1862 1400 1868 1401
rect 3574 1401 3575 1405
rect 3579 1401 3580 1405
rect 3574 1400 3580 1401
rect 110 1392 116 1393
rect 1822 1392 1828 1393
rect 110 1388 111 1392
rect 115 1388 116 1392
rect 527 1391 533 1392
rect 527 1390 528 1391
rect 517 1388 528 1390
rect 110 1387 116 1388
rect 182 1387 188 1388
rect 182 1383 183 1387
rect 187 1386 188 1387
rect 270 1387 276 1388
rect 187 1384 217 1386
rect 187 1383 188 1384
rect 182 1382 188 1383
rect 270 1383 271 1387
rect 275 1386 276 1387
rect 527 1387 528 1388
rect 532 1387 533 1391
rect 879 1391 885 1392
rect 879 1390 880 1391
rect 869 1388 880 1390
rect 527 1386 533 1387
rect 658 1387 664 1388
rect 275 1384 353 1386
rect 275 1383 276 1384
rect 270 1382 276 1383
rect 658 1383 659 1387
rect 663 1386 664 1387
rect 879 1387 880 1388
rect 884 1387 885 1391
rect 983 1391 989 1392
rect 983 1390 984 1391
rect 973 1388 984 1390
rect 879 1386 885 1387
rect 983 1387 984 1388
rect 988 1387 989 1391
rect 1079 1391 1085 1392
rect 1079 1390 1080 1391
rect 1069 1388 1080 1390
rect 983 1386 989 1387
rect 1079 1387 1080 1388
rect 1084 1387 1085 1391
rect 1287 1391 1293 1392
rect 1287 1390 1288 1391
rect 1277 1388 1288 1390
rect 1079 1386 1085 1387
rect 1110 1387 1116 1388
rect 663 1384 721 1386
rect 663 1383 664 1384
rect 658 1382 664 1383
rect 1110 1383 1111 1387
rect 1115 1386 1116 1387
rect 1287 1387 1288 1388
rect 1292 1387 1293 1391
rect 1822 1388 1823 1392
rect 1827 1388 1828 1392
rect 1879 1391 1885 1392
rect 1822 1387 1828 1388
rect 1862 1388 1868 1389
rect 1287 1386 1293 1387
rect 1115 1384 1137 1386
rect 1862 1384 1863 1388
rect 1867 1384 1868 1388
rect 1879 1387 1880 1391
rect 1884 1390 1885 1391
rect 1954 1391 1960 1392
rect 1884 1388 1913 1390
rect 1884 1387 1885 1388
rect 1879 1386 1885 1387
rect 1954 1387 1955 1391
rect 1959 1390 1960 1391
rect 2042 1391 2048 1392
rect 1959 1388 2001 1390
rect 1959 1387 1960 1388
rect 1954 1386 1960 1387
rect 2042 1387 2043 1391
rect 2047 1390 2048 1391
rect 2250 1391 2256 1392
rect 2250 1390 2251 1391
rect 2047 1388 2097 1390
rect 2245 1388 2251 1390
rect 2047 1387 2048 1388
rect 2042 1386 2048 1387
rect 2250 1387 2251 1388
rect 2255 1387 2256 1391
rect 2250 1386 2256 1387
rect 2370 1391 2376 1392
rect 2370 1387 2371 1391
rect 2375 1390 2376 1391
rect 2506 1391 2512 1392
rect 2375 1388 2465 1390
rect 2375 1387 2376 1388
rect 2370 1386 2376 1387
rect 2506 1387 2507 1391
rect 2511 1390 2512 1391
rect 3023 1391 3029 1392
rect 3023 1390 3024 1391
rect 2511 1388 2633 1390
rect 2869 1388 3024 1390
rect 2511 1387 2512 1388
rect 2506 1386 2512 1387
rect 3023 1387 3024 1388
rect 3028 1387 3029 1391
rect 3254 1391 3260 1392
rect 3254 1390 3255 1391
rect 3093 1388 3255 1390
rect 3023 1386 3029 1387
rect 3254 1387 3255 1388
rect 3259 1387 3260 1391
rect 3254 1386 3260 1387
rect 3470 1391 3476 1392
rect 3470 1387 3471 1391
rect 3475 1390 3476 1391
rect 3475 1388 3505 1390
rect 3574 1388 3580 1389
rect 3475 1387 3476 1388
rect 3470 1386 3476 1387
rect 1115 1383 1116 1384
rect 1862 1383 1868 1384
rect 3574 1384 3575 1388
rect 3579 1384 3580 1388
rect 3574 1383 3580 1384
rect 1110 1382 1116 1383
rect 110 1375 116 1376
rect 110 1371 111 1375
rect 115 1371 116 1375
rect 687 1375 693 1376
rect 687 1374 688 1375
rect 633 1372 688 1374
rect 110 1370 116 1371
rect 687 1371 688 1372
rect 692 1371 693 1375
rect 687 1370 693 1371
rect 1822 1375 1828 1376
rect 1822 1371 1823 1375
rect 1827 1371 1828 1375
rect 1822 1370 1828 1371
rect 1894 1375 1900 1376
rect 1894 1371 1895 1375
rect 1899 1371 1900 1375
rect 1894 1370 1900 1371
rect 1982 1375 1988 1376
rect 1982 1371 1983 1375
rect 1987 1371 1988 1375
rect 1982 1370 1988 1371
rect 2078 1375 2084 1376
rect 2078 1371 2079 1375
rect 2083 1371 2084 1375
rect 2078 1370 2084 1371
rect 2190 1375 2196 1376
rect 2190 1371 2191 1375
rect 2195 1371 2196 1375
rect 2190 1370 2196 1371
rect 2310 1375 2316 1376
rect 2310 1371 2311 1375
rect 2315 1371 2316 1375
rect 2310 1370 2316 1371
rect 2446 1375 2452 1376
rect 2446 1371 2447 1375
rect 2451 1371 2452 1375
rect 2446 1370 2452 1371
rect 2614 1375 2620 1376
rect 2614 1371 2615 1375
rect 2619 1371 2620 1375
rect 2614 1370 2620 1371
rect 2814 1375 2820 1376
rect 2814 1371 2815 1375
rect 2819 1371 2820 1375
rect 2814 1370 2820 1371
rect 3038 1375 3044 1376
rect 3038 1371 3039 1375
rect 3043 1371 3044 1375
rect 3038 1370 3044 1371
rect 3270 1375 3276 1376
rect 3270 1371 3271 1375
rect 3275 1371 3276 1375
rect 3270 1370 3276 1371
rect 3486 1375 3492 1376
rect 3486 1371 3487 1375
rect 3491 1371 3492 1375
rect 3486 1370 3492 1371
rect 190 1365 196 1366
rect 190 1361 191 1365
rect 195 1361 196 1365
rect 190 1360 196 1361
rect 326 1365 332 1366
rect 326 1361 327 1365
rect 331 1361 332 1365
rect 326 1360 332 1361
rect 454 1365 460 1366
rect 454 1361 455 1365
rect 459 1361 460 1365
rect 454 1360 460 1361
rect 574 1365 580 1366
rect 574 1361 575 1365
rect 579 1361 580 1365
rect 574 1360 580 1361
rect 694 1365 700 1366
rect 694 1361 695 1365
rect 699 1361 700 1365
rect 694 1360 700 1361
rect 806 1365 812 1366
rect 806 1361 807 1365
rect 811 1361 812 1365
rect 806 1360 812 1361
rect 910 1365 916 1366
rect 910 1361 911 1365
rect 915 1361 916 1365
rect 910 1360 916 1361
rect 1006 1365 1012 1366
rect 1006 1361 1007 1365
rect 1011 1361 1012 1365
rect 1006 1360 1012 1361
rect 1110 1365 1116 1366
rect 1110 1361 1111 1365
rect 1115 1361 1116 1365
rect 1110 1360 1116 1361
rect 1214 1365 1220 1366
rect 1214 1361 1215 1365
rect 1219 1361 1220 1365
rect 1214 1360 1220 1361
rect 1318 1365 1324 1366
rect 1318 1361 1319 1365
rect 1323 1361 1324 1365
rect 1318 1360 1324 1361
rect 1887 1363 1893 1364
rect 1366 1359 1373 1360
rect 1366 1355 1367 1359
rect 1372 1355 1373 1359
rect 1887 1359 1888 1363
rect 1892 1362 1893 1363
rect 1954 1363 1960 1364
rect 1954 1362 1955 1363
rect 1892 1360 1955 1362
rect 1892 1359 1893 1360
rect 1887 1358 1893 1359
rect 1954 1359 1955 1360
rect 1959 1359 1960 1363
rect 1954 1358 1960 1359
rect 1975 1363 1981 1364
rect 1975 1359 1976 1363
rect 1980 1362 1981 1363
rect 2042 1363 2048 1364
rect 2042 1362 2043 1363
rect 1980 1360 2043 1362
rect 1980 1359 1981 1360
rect 1975 1358 1981 1359
rect 2042 1359 2043 1360
rect 2047 1359 2048 1363
rect 2042 1358 2048 1359
rect 2063 1363 2069 1364
rect 2063 1359 2064 1363
rect 2068 1362 2069 1363
rect 2071 1363 2077 1364
rect 2071 1362 2072 1363
rect 2068 1360 2072 1362
rect 2068 1359 2069 1360
rect 2063 1358 2069 1359
rect 2071 1359 2072 1360
rect 2076 1359 2077 1363
rect 2071 1358 2077 1359
rect 2183 1363 2189 1364
rect 2183 1359 2184 1363
rect 2188 1362 2189 1363
rect 2191 1363 2197 1364
rect 2191 1362 2192 1363
rect 2188 1360 2192 1362
rect 2188 1359 2189 1360
rect 2183 1358 2189 1359
rect 2191 1359 2192 1360
rect 2196 1359 2197 1363
rect 2191 1358 2197 1359
rect 2250 1363 2256 1364
rect 2250 1359 2251 1363
rect 2255 1362 2256 1363
rect 2303 1363 2309 1364
rect 2303 1362 2304 1363
rect 2255 1360 2304 1362
rect 2255 1359 2256 1360
rect 2250 1358 2256 1359
rect 2303 1359 2304 1360
rect 2308 1359 2309 1363
rect 2303 1358 2309 1359
rect 2439 1363 2445 1364
rect 2439 1359 2440 1363
rect 2444 1362 2445 1363
rect 2506 1363 2512 1364
rect 2506 1362 2507 1363
rect 2444 1360 2507 1362
rect 2444 1359 2445 1360
rect 2439 1358 2445 1359
rect 2506 1359 2507 1360
rect 2511 1359 2512 1363
rect 2506 1358 2512 1359
rect 2607 1363 2613 1364
rect 2607 1359 2608 1363
rect 2612 1362 2613 1363
rect 2774 1363 2780 1364
rect 2774 1362 2775 1363
rect 2612 1360 2775 1362
rect 2612 1359 2613 1360
rect 2607 1358 2613 1359
rect 2774 1359 2775 1360
rect 2779 1359 2780 1363
rect 2774 1358 2780 1359
rect 2799 1363 2805 1364
rect 2799 1359 2800 1363
rect 2804 1362 2805 1363
rect 2807 1363 2813 1364
rect 2807 1362 2808 1363
rect 2804 1360 2808 1362
rect 2804 1359 2805 1360
rect 2799 1358 2805 1359
rect 2807 1359 2808 1360
rect 2812 1359 2813 1363
rect 2807 1358 2813 1359
rect 3023 1363 3029 1364
rect 3023 1359 3024 1363
rect 3028 1362 3029 1363
rect 3031 1363 3037 1364
rect 3031 1362 3032 1363
rect 3028 1360 3032 1362
rect 3028 1359 3029 1360
rect 3023 1358 3029 1359
rect 3031 1359 3032 1360
rect 3036 1359 3037 1363
rect 3031 1358 3037 1359
rect 3254 1363 3260 1364
rect 3254 1359 3255 1363
rect 3259 1362 3260 1363
rect 3263 1363 3269 1364
rect 3263 1362 3264 1363
rect 3259 1360 3264 1362
rect 3259 1359 3260 1360
rect 3254 1358 3260 1359
rect 3263 1359 3264 1360
rect 3268 1359 3269 1363
rect 3263 1358 3269 1359
rect 3471 1363 3477 1364
rect 3471 1359 3472 1363
rect 3476 1362 3477 1363
rect 3479 1363 3485 1364
rect 3479 1362 3480 1363
rect 3476 1360 3480 1362
rect 3476 1359 3477 1360
rect 3471 1358 3477 1359
rect 3479 1359 3480 1360
rect 3484 1359 3485 1363
rect 3479 1358 3485 1359
rect 1366 1354 1373 1355
rect 1879 1347 1885 1348
rect 1879 1343 1880 1347
rect 1884 1346 1885 1347
rect 1887 1347 1893 1348
rect 1887 1346 1888 1347
rect 1884 1344 1888 1346
rect 1884 1343 1885 1344
rect 1879 1342 1885 1343
rect 1887 1343 1888 1344
rect 1892 1343 1893 1347
rect 1887 1342 1893 1343
rect 1959 1347 1965 1348
rect 1959 1343 1960 1347
rect 1964 1346 1965 1347
rect 1975 1347 1981 1348
rect 1975 1346 1976 1347
rect 1964 1344 1976 1346
rect 1964 1343 1965 1344
rect 1959 1342 1965 1343
rect 1975 1343 1976 1344
rect 1980 1343 1981 1347
rect 1975 1342 1981 1343
rect 2047 1347 2053 1348
rect 2047 1343 2048 1347
rect 2052 1346 2053 1347
rect 2095 1347 2101 1348
rect 2095 1346 2096 1347
rect 2052 1344 2096 1346
rect 2052 1343 2053 1344
rect 2047 1342 2053 1343
rect 2095 1343 2096 1344
rect 2100 1343 2101 1347
rect 2095 1342 2101 1343
rect 2167 1347 2173 1348
rect 2167 1343 2168 1347
rect 2172 1346 2173 1347
rect 2215 1347 2221 1348
rect 2215 1346 2216 1347
rect 2172 1344 2216 1346
rect 2172 1343 2173 1344
rect 2167 1342 2173 1343
rect 2215 1343 2216 1344
rect 2220 1343 2221 1347
rect 2215 1342 2221 1343
rect 2351 1347 2357 1348
rect 2351 1343 2352 1347
rect 2356 1346 2357 1347
rect 2370 1347 2376 1348
rect 2370 1346 2371 1347
rect 2356 1344 2371 1346
rect 2356 1343 2357 1344
rect 2351 1342 2357 1343
rect 2370 1343 2371 1344
rect 2375 1343 2376 1347
rect 2370 1342 2376 1343
rect 2431 1347 2437 1348
rect 2431 1343 2432 1347
rect 2436 1346 2437 1347
rect 2503 1347 2509 1348
rect 2503 1346 2504 1347
rect 2436 1344 2504 1346
rect 2436 1343 2437 1344
rect 2431 1342 2437 1343
rect 2503 1343 2504 1344
rect 2508 1343 2509 1347
rect 2503 1342 2509 1343
rect 2599 1347 2605 1348
rect 2599 1343 2600 1347
rect 2604 1346 2605 1347
rect 2679 1347 2685 1348
rect 2679 1346 2680 1347
rect 2604 1344 2680 1346
rect 2604 1343 2605 1344
rect 2599 1342 2605 1343
rect 2679 1343 2680 1344
rect 2684 1343 2685 1347
rect 2679 1342 2685 1343
rect 2775 1347 2781 1348
rect 2775 1343 2776 1347
rect 2780 1346 2781 1347
rect 2863 1347 2869 1348
rect 2863 1346 2864 1347
rect 2780 1344 2864 1346
rect 2780 1343 2781 1344
rect 2775 1342 2781 1343
rect 2863 1343 2864 1344
rect 2868 1343 2869 1347
rect 2863 1342 2869 1343
rect 2967 1347 2973 1348
rect 2967 1343 2968 1347
rect 2972 1346 2973 1347
rect 3063 1347 3069 1348
rect 3063 1346 3064 1347
rect 2972 1344 3064 1346
rect 2972 1343 2973 1344
rect 2967 1342 2973 1343
rect 3063 1343 3064 1344
rect 3068 1343 3069 1347
rect 3063 1342 3069 1343
rect 3254 1347 3260 1348
rect 3254 1343 3255 1347
rect 3259 1346 3260 1347
rect 3271 1347 3277 1348
rect 3271 1346 3272 1347
rect 3259 1344 3272 1346
rect 3259 1343 3260 1344
rect 3254 1342 3260 1343
rect 3271 1343 3272 1344
rect 3276 1343 3277 1347
rect 3271 1342 3277 1343
rect 3470 1347 3476 1348
rect 3470 1343 3471 1347
rect 3475 1346 3476 1347
rect 3479 1347 3485 1348
rect 3479 1346 3480 1347
rect 3475 1344 3480 1346
rect 3475 1343 3476 1344
rect 3470 1342 3476 1343
rect 3479 1343 3480 1344
rect 3484 1343 3485 1347
rect 3479 1342 3485 1343
rect 230 1339 236 1340
rect 230 1335 231 1339
rect 235 1335 236 1339
rect 230 1334 236 1335
rect 382 1339 388 1340
rect 382 1335 383 1339
rect 387 1335 388 1339
rect 382 1334 388 1335
rect 542 1339 548 1340
rect 542 1335 543 1339
rect 547 1335 548 1339
rect 542 1334 548 1335
rect 702 1339 708 1340
rect 702 1335 703 1339
rect 707 1335 708 1339
rect 702 1334 708 1335
rect 870 1339 876 1340
rect 870 1335 871 1339
rect 875 1335 876 1339
rect 870 1334 876 1335
rect 1038 1339 1044 1340
rect 1038 1335 1039 1339
rect 1043 1335 1044 1339
rect 1038 1334 1044 1335
rect 1206 1339 1212 1340
rect 1206 1335 1207 1339
rect 1211 1335 1212 1339
rect 1206 1334 1212 1335
rect 1374 1339 1380 1340
rect 1374 1335 1375 1339
rect 1379 1335 1380 1339
rect 1374 1334 1380 1335
rect 1894 1337 1900 1338
rect 1894 1333 1895 1337
rect 1899 1333 1900 1337
rect 1894 1332 1900 1333
rect 1982 1337 1988 1338
rect 1982 1333 1983 1337
rect 1987 1333 1988 1337
rect 1982 1332 1988 1333
rect 2102 1337 2108 1338
rect 2102 1333 2103 1337
rect 2107 1333 2108 1337
rect 2102 1332 2108 1333
rect 2222 1337 2228 1338
rect 2222 1333 2223 1337
rect 2227 1333 2228 1337
rect 2222 1332 2228 1333
rect 2358 1337 2364 1338
rect 2358 1333 2359 1337
rect 2363 1333 2364 1337
rect 2358 1332 2364 1333
rect 2510 1337 2516 1338
rect 2510 1333 2511 1337
rect 2515 1333 2516 1337
rect 2510 1332 2516 1333
rect 2686 1337 2692 1338
rect 2686 1333 2687 1337
rect 2691 1333 2692 1337
rect 2686 1332 2692 1333
rect 2870 1337 2876 1338
rect 2870 1333 2871 1337
rect 2875 1333 2876 1337
rect 2870 1332 2876 1333
rect 3070 1337 3076 1338
rect 3070 1333 3071 1337
rect 3075 1333 3076 1337
rect 3070 1332 3076 1333
rect 3278 1337 3284 1338
rect 3278 1333 3279 1337
rect 3283 1333 3284 1337
rect 3278 1332 3284 1333
rect 3486 1337 3492 1338
rect 3486 1333 3487 1337
rect 3491 1333 3492 1337
rect 3486 1332 3492 1333
rect 298 1331 304 1332
rect 298 1330 299 1331
rect 110 1329 116 1330
rect 110 1325 111 1329
rect 115 1325 116 1329
rect 289 1328 299 1330
rect 298 1327 299 1328
rect 303 1327 304 1331
rect 770 1331 776 1332
rect 770 1330 771 1331
rect 761 1328 771 1330
rect 298 1326 304 1327
rect 770 1327 771 1328
rect 775 1327 776 1331
rect 770 1326 776 1327
rect 1822 1329 1828 1330
rect 110 1324 116 1325
rect 1822 1325 1823 1329
rect 1827 1325 1828 1329
rect 1822 1324 1828 1325
rect 1862 1324 1868 1325
rect 3574 1324 3580 1325
rect 1862 1320 1863 1324
rect 1867 1320 1868 1324
rect 1959 1323 1965 1324
rect 1959 1322 1960 1323
rect 1949 1320 1960 1322
rect 1862 1319 1868 1320
rect 1959 1319 1960 1320
rect 1964 1319 1965 1323
rect 2047 1323 2053 1324
rect 2047 1322 2048 1323
rect 2037 1320 2048 1322
rect 1959 1318 1965 1319
rect 2047 1319 2048 1320
rect 2052 1319 2053 1323
rect 2167 1323 2173 1324
rect 2167 1322 2168 1323
rect 2157 1320 2168 1322
rect 2047 1318 2053 1319
rect 2167 1319 2168 1320
rect 2172 1319 2173 1323
rect 2431 1323 2437 1324
rect 2431 1322 2432 1323
rect 2413 1320 2432 1322
rect 2167 1318 2173 1319
rect 2191 1319 2197 1320
rect 319 1315 325 1316
rect 110 1312 116 1313
rect 110 1308 111 1312
rect 115 1308 116 1312
rect 319 1311 320 1315
rect 324 1314 325 1315
rect 450 1315 456 1316
rect 324 1312 409 1314
rect 324 1311 325 1312
rect 319 1310 325 1311
rect 450 1311 451 1315
rect 455 1314 456 1315
rect 798 1315 804 1316
rect 455 1312 569 1314
rect 455 1311 456 1312
rect 450 1310 456 1311
rect 798 1311 799 1315
rect 803 1314 804 1315
rect 999 1315 1005 1316
rect 803 1312 897 1314
rect 803 1311 804 1312
rect 798 1310 804 1311
rect 999 1311 1000 1315
rect 1004 1314 1005 1315
rect 1106 1315 1112 1316
rect 1004 1312 1065 1314
rect 1004 1311 1005 1312
rect 999 1310 1005 1311
rect 1106 1311 1107 1315
rect 1111 1314 1112 1315
rect 1274 1315 1280 1316
rect 1111 1312 1233 1314
rect 1111 1311 1112 1312
rect 1106 1310 1112 1311
rect 1274 1311 1275 1315
rect 1279 1314 1280 1315
rect 2191 1315 2192 1319
rect 2196 1318 2197 1319
rect 2431 1319 2432 1320
rect 2436 1319 2437 1323
rect 2599 1323 2605 1324
rect 2599 1322 2600 1323
rect 2565 1320 2600 1322
rect 2431 1318 2437 1319
rect 2599 1319 2600 1320
rect 2604 1319 2605 1323
rect 2775 1323 2781 1324
rect 2775 1322 2776 1323
rect 2741 1320 2776 1322
rect 2599 1318 2605 1319
rect 2775 1319 2776 1320
rect 2780 1319 2781 1323
rect 2967 1323 2973 1324
rect 2967 1322 2968 1323
rect 2925 1320 2968 1322
rect 2775 1318 2781 1319
rect 2967 1319 2968 1320
rect 2972 1319 2973 1323
rect 3367 1323 3373 1324
rect 3367 1322 3368 1323
rect 3333 1320 3368 1322
rect 2967 1318 2973 1319
rect 3367 1319 3368 1320
rect 3372 1319 3373 1323
rect 3574 1320 3575 1324
rect 3579 1320 3580 1324
rect 3574 1319 3580 1320
rect 3367 1318 3373 1319
rect 2196 1316 2241 1318
rect 2196 1315 2197 1316
rect 2191 1314 2197 1315
rect 1279 1312 1401 1314
rect 1822 1312 1828 1313
rect 1279 1311 1280 1312
rect 1274 1310 1280 1311
rect 110 1307 116 1308
rect 1822 1308 1823 1312
rect 1827 1308 1828 1312
rect 1822 1307 1828 1308
rect 1862 1307 1868 1308
rect 1862 1303 1863 1307
rect 1867 1303 1868 1307
rect 1862 1302 1868 1303
rect 2958 1307 2964 1308
rect 2958 1303 2959 1307
rect 2963 1306 2964 1307
rect 3454 1307 3460 1308
rect 2963 1304 3081 1306
rect 2963 1303 2964 1304
rect 2958 1302 2964 1303
rect 3454 1303 3455 1307
rect 3459 1306 3460 1307
rect 3574 1307 3580 1308
rect 3459 1304 3497 1306
rect 3459 1303 3460 1304
rect 3454 1302 3460 1303
rect 3574 1303 3575 1307
rect 3579 1303 3580 1307
rect 3574 1302 3580 1303
rect 238 1299 244 1300
rect 238 1295 239 1299
rect 243 1295 244 1299
rect 238 1294 244 1295
rect 390 1299 396 1300
rect 390 1295 391 1299
rect 395 1295 396 1299
rect 390 1294 396 1295
rect 550 1299 556 1300
rect 550 1295 551 1299
rect 555 1295 556 1299
rect 550 1294 556 1295
rect 710 1299 716 1300
rect 710 1295 711 1299
rect 715 1295 716 1299
rect 710 1294 716 1295
rect 878 1299 884 1300
rect 878 1295 879 1299
rect 883 1295 884 1299
rect 878 1294 884 1295
rect 1046 1299 1052 1300
rect 1046 1295 1047 1299
rect 1051 1295 1052 1299
rect 1046 1294 1052 1295
rect 1214 1299 1220 1300
rect 1214 1295 1215 1299
rect 1219 1295 1220 1299
rect 1214 1294 1220 1295
rect 1382 1299 1388 1300
rect 1382 1295 1383 1299
rect 1387 1295 1388 1299
rect 1382 1294 1388 1295
rect 1886 1297 1892 1298
rect 1886 1293 1887 1297
rect 1891 1293 1892 1297
rect 1886 1292 1892 1293
rect 1974 1297 1980 1298
rect 1974 1293 1975 1297
rect 1979 1293 1980 1297
rect 1974 1292 1980 1293
rect 2094 1297 2100 1298
rect 2094 1293 2095 1297
rect 2099 1293 2100 1297
rect 2094 1292 2100 1293
rect 2214 1297 2220 1298
rect 2214 1293 2215 1297
rect 2219 1293 2220 1297
rect 2214 1292 2220 1293
rect 2350 1297 2356 1298
rect 2350 1293 2351 1297
rect 2355 1293 2356 1297
rect 2350 1292 2356 1293
rect 2502 1297 2508 1298
rect 2502 1293 2503 1297
rect 2507 1293 2508 1297
rect 2502 1292 2508 1293
rect 2678 1297 2684 1298
rect 2678 1293 2679 1297
rect 2683 1293 2684 1297
rect 2678 1292 2684 1293
rect 2862 1297 2868 1298
rect 2862 1293 2863 1297
rect 2867 1293 2868 1297
rect 2862 1292 2868 1293
rect 3062 1297 3068 1298
rect 3062 1293 3063 1297
rect 3067 1293 3068 1297
rect 3062 1292 3068 1293
rect 3270 1297 3276 1298
rect 3270 1293 3271 1297
rect 3275 1293 3276 1297
rect 3270 1292 3276 1293
rect 3478 1297 3484 1298
rect 3478 1293 3479 1297
rect 3483 1293 3484 1297
rect 3478 1292 3484 1293
rect 231 1287 237 1288
rect 231 1283 232 1287
rect 236 1286 237 1287
rect 319 1287 325 1288
rect 319 1286 320 1287
rect 236 1284 320 1286
rect 236 1283 237 1284
rect 231 1282 237 1283
rect 319 1283 320 1284
rect 324 1283 325 1287
rect 319 1282 325 1283
rect 383 1287 389 1288
rect 383 1283 384 1287
rect 388 1286 389 1287
rect 450 1287 456 1288
rect 450 1286 451 1287
rect 388 1284 451 1286
rect 388 1283 389 1284
rect 383 1282 389 1283
rect 450 1283 451 1284
rect 455 1283 456 1287
rect 450 1282 456 1283
rect 543 1287 549 1288
rect 543 1283 544 1287
rect 548 1286 549 1287
rect 558 1287 564 1288
rect 558 1286 559 1287
rect 548 1284 559 1286
rect 548 1283 549 1284
rect 543 1282 549 1283
rect 558 1283 559 1284
rect 563 1283 564 1287
rect 558 1282 564 1283
rect 687 1287 693 1288
rect 687 1283 688 1287
rect 692 1286 693 1287
rect 703 1287 709 1288
rect 703 1286 704 1287
rect 692 1284 704 1286
rect 692 1283 693 1284
rect 687 1282 693 1283
rect 703 1283 704 1284
rect 708 1283 709 1287
rect 703 1282 709 1283
rect 871 1287 877 1288
rect 871 1283 872 1287
rect 876 1286 877 1287
rect 898 1287 904 1288
rect 898 1286 899 1287
rect 876 1284 899 1286
rect 876 1283 877 1284
rect 871 1282 877 1283
rect 898 1283 899 1284
rect 903 1283 904 1287
rect 898 1282 904 1283
rect 1039 1287 1045 1288
rect 1039 1283 1040 1287
rect 1044 1286 1045 1287
rect 1106 1287 1112 1288
rect 1106 1286 1107 1287
rect 1044 1284 1107 1286
rect 1044 1283 1045 1284
rect 1039 1282 1045 1283
rect 1106 1283 1107 1284
rect 1111 1283 1112 1287
rect 1106 1282 1112 1283
rect 1207 1287 1213 1288
rect 1207 1283 1208 1287
rect 1212 1286 1213 1287
rect 1274 1287 1280 1288
rect 1274 1286 1275 1287
rect 1212 1284 1275 1286
rect 1212 1283 1213 1284
rect 1207 1282 1213 1283
rect 1274 1283 1275 1284
rect 1279 1283 1280 1287
rect 1274 1282 1280 1283
rect 1366 1287 1372 1288
rect 1366 1283 1367 1287
rect 1371 1286 1372 1287
rect 1375 1287 1381 1288
rect 1375 1286 1376 1287
rect 1371 1284 1376 1286
rect 1371 1283 1372 1284
rect 1366 1282 1372 1283
rect 1375 1283 1376 1284
rect 1380 1283 1381 1287
rect 1375 1282 1381 1283
rect 198 1275 204 1276
rect 198 1271 199 1275
rect 203 1274 204 1275
rect 207 1275 213 1276
rect 207 1274 208 1275
rect 203 1272 208 1274
rect 203 1271 204 1272
rect 198 1270 204 1271
rect 207 1271 208 1272
rect 212 1271 213 1275
rect 207 1270 213 1271
rect 287 1275 293 1276
rect 287 1271 288 1275
rect 292 1274 293 1275
rect 351 1275 357 1276
rect 351 1274 352 1275
rect 292 1272 352 1274
rect 292 1271 293 1272
rect 287 1270 293 1271
rect 351 1271 352 1272
rect 356 1271 357 1275
rect 351 1270 357 1271
rect 439 1275 445 1276
rect 439 1271 440 1275
rect 444 1274 445 1275
rect 511 1275 517 1276
rect 511 1274 512 1275
rect 444 1272 512 1274
rect 444 1271 445 1272
rect 439 1270 445 1271
rect 511 1271 512 1272
rect 516 1271 517 1275
rect 511 1270 517 1271
rect 583 1275 589 1276
rect 583 1271 584 1275
rect 588 1274 589 1275
rect 671 1275 677 1276
rect 671 1274 672 1275
rect 588 1272 672 1274
rect 588 1271 589 1272
rect 583 1270 589 1271
rect 671 1271 672 1272
rect 676 1271 677 1275
rect 671 1270 677 1271
rect 759 1275 765 1276
rect 759 1271 760 1275
rect 764 1274 765 1275
rect 831 1275 837 1276
rect 831 1274 832 1275
rect 764 1272 832 1274
rect 764 1271 765 1272
rect 759 1270 765 1271
rect 831 1271 832 1272
rect 836 1271 837 1275
rect 831 1270 837 1271
rect 991 1275 997 1276
rect 991 1271 992 1275
rect 996 1274 997 1275
rect 999 1275 1005 1276
rect 999 1274 1000 1275
rect 996 1272 1000 1274
rect 996 1271 997 1272
rect 991 1270 997 1271
rect 999 1271 1000 1272
rect 1004 1271 1005 1275
rect 999 1270 1005 1271
rect 1071 1275 1077 1276
rect 1071 1271 1072 1275
rect 1076 1274 1077 1275
rect 1143 1275 1149 1276
rect 1143 1274 1144 1275
rect 1076 1272 1144 1274
rect 1076 1271 1077 1272
rect 1071 1270 1077 1271
rect 1143 1271 1144 1272
rect 1148 1271 1149 1275
rect 1143 1270 1149 1271
rect 1223 1275 1229 1276
rect 1223 1271 1224 1275
rect 1228 1274 1229 1275
rect 1287 1275 1293 1276
rect 1287 1274 1288 1275
rect 1228 1272 1288 1274
rect 1228 1271 1229 1272
rect 1223 1270 1229 1271
rect 1287 1271 1288 1272
rect 1292 1271 1293 1275
rect 1287 1270 1293 1271
rect 1367 1275 1373 1276
rect 1367 1271 1368 1275
rect 1372 1274 1373 1275
rect 1431 1275 1437 1276
rect 1431 1274 1432 1275
rect 1372 1272 1432 1274
rect 1372 1271 1373 1272
rect 1367 1270 1373 1271
rect 1431 1271 1432 1272
rect 1436 1271 1437 1275
rect 1431 1270 1437 1271
rect 1575 1275 1581 1276
rect 1575 1271 1576 1275
rect 1580 1274 1581 1275
rect 1583 1275 1589 1276
rect 1583 1274 1584 1275
rect 1580 1272 1584 1274
rect 1580 1271 1581 1272
rect 1575 1270 1581 1271
rect 1583 1271 1584 1272
rect 1588 1271 1589 1275
rect 1583 1270 1589 1271
rect 214 1265 220 1266
rect 214 1261 215 1265
rect 219 1261 220 1265
rect 214 1260 220 1261
rect 358 1265 364 1266
rect 358 1261 359 1265
rect 363 1261 364 1265
rect 358 1260 364 1261
rect 518 1265 524 1266
rect 518 1261 519 1265
rect 523 1261 524 1265
rect 518 1260 524 1261
rect 678 1265 684 1266
rect 678 1261 679 1265
rect 683 1261 684 1265
rect 678 1260 684 1261
rect 838 1265 844 1266
rect 838 1261 839 1265
rect 843 1261 844 1265
rect 838 1260 844 1261
rect 998 1265 1004 1266
rect 998 1261 999 1265
rect 1003 1261 1004 1265
rect 998 1260 1004 1261
rect 1150 1265 1156 1266
rect 1150 1261 1151 1265
rect 1155 1261 1156 1265
rect 1150 1260 1156 1261
rect 1294 1265 1300 1266
rect 1294 1261 1295 1265
rect 1299 1261 1300 1265
rect 1294 1260 1300 1261
rect 1438 1265 1444 1266
rect 1438 1261 1439 1265
rect 1443 1261 1444 1265
rect 1438 1260 1444 1261
rect 1590 1265 1596 1266
rect 1590 1261 1591 1265
rect 1595 1261 1596 1265
rect 1590 1260 1596 1261
rect 2054 1263 2060 1264
rect 2054 1259 2055 1263
rect 2059 1259 2060 1263
rect 2054 1258 2060 1259
rect 2142 1263 2148 1264
rect 2142 1259 2143 1263
rect 2147 1259 2148 1263
rect 2142 1258 2148 1259
rect 2238 1263 2244 1264
rect 2238 1259 2239 1263
rect 2243 1259 2244 1263
rect 2238 1258 2244 1259
rect 2334 1263 2340 1264
rect 2334 1259 2335 1263
rect 2339 1259 2340 1263
rect 2334 1258 2340 1259
rect 2430 1263 2436 1264
rect 2430 1259 2431 1263
rect 2435 1259 2436 1263
rect 2430 1258 2436 1259
rect 2550 1263 2556 1264
rect 2550 1259 2551 1263
rect 2555 1259 2556 1263
rect 2550 1258 2556 1259
rect 2686 1263 2692 1264
rect 2686 1259 2687 1263
rect 2691 1259 2692 1263
rect 2686 1258 2692 1259
rect 2854 1263 2860 1264
rect 2854 1259 2855 1263
rect 2859 1259 2860 1263
rect 2854 1258 2860 1259
rect 3038 1263 3044 1264
rect 3038 1259 3039 1263
rect 3043 1259 3044 1263
rect 3038 1258 3044 1259
rect 3230 1263 3236 1264
rect 3230 1259 3231 1263
rect 3235 1259 3236 1263
rect 3230 1258 3236 1259
rect 3430 1263 3436 1264
rect 3430 1259 3431 1263
rect 3435 1259 3436 1263
rect 3430 1258 3436 1259
rect 2122 1255 2128 1256
rect 1862 1253 1868 1254
rect 110 1252 116 1253
rect 1822 1252 1828 1253
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 287 1251 293 1252
rect 287 1250 288 1251
rect 269 1248 288 1250
rect 110 1247 116 1248
rect 287 1247 288 1248
rect 292 1247 293 1251
rect 439 1251 445 1252
rect 439 1250 440 1251
rect 413 1248 440 1250
rect 287 1246 293 1247
rect 439 1247 440 1248
rect 444 1247 445 1251
rect 583 1251 589 1252
rect 583 1250 584 1251
rect 573 1248 584 1250
rect 439 1246 445 1247
rect 583 1247 584 1248
rect 588 1247 589 1251
rect 759 1251 765 1252
rect 759 1250 760 1251
rect 733 1248 760 1250
rect 583 1246 589 1247
rect 759 1247 760 1248
rect 764 1247 765 1251
rect 898 1251 904 1252
rect 898 1250 899 1251
rect 893 1248 899 1250
rect 759 1246 765 1247
rect 898 1247 899 1248
rect 903 1247 904 1251
rect 1071 1251 1077 1252
rect 1071 1250 1072 1251
rect 1053 1248 1072 1250
rect 898 1246 904 1247
rect 1071 1247 1072 1248
rect 1076 1247 1077 1251
rect 1223 1251 1229 1252
rect 1223 1250 1224 1251
rect 1205 1248 1224 1250
rect 1071 1246 1077 1247
rect 1223 1247 1224 1248
rect 1228 1247 1229 1251
rect 1367 1251 1373 1252
rect 1367 1250 1368 1251
rect 1349 1248 1368 1250
rect 1223 1246 1229 1247
rect 1367 1247 1368 1248
rect 1372 1247 1373 1251
rect 1575 1251 1581 1252
rect 1575 1250 1576 1251
rect 1493 1248 1576 1250
rect 1367 1246 1373 1247
rect 1575 1247 1576 1248
rect 1580 1247 1581 1251
rect 1822 1248 1823 1252
rect 1827 1248 1828 1252
rect 1862 1249 1863 1253
rect 1867 1249 1868 1253
rect 2122 1251 2123 1255
rect 2127 1254 2128 1255
rect 3106 1255 3112 1256
rect 2127 1252 2161 1254
rect 2127 1251 2128 1252
rect 2122 1250 2128 1251
rect 3106 1251 3107 1255
rect 3111 1254 3112 1255
rect 3111 1252 3249 1254
rect 3574 1253 3580 1254
rect 3111 1251 3112 1252
rect 3106 1250 3112 1251
rect 1862 1248 1868 1249
rect 3574 1249 3575 1253
rect 3579 1249 3580 1253
rect 3574 1248 3580 1249
rect 1822 1247 1828 1248
rect 1575 1246 1581 1247
rect 2135 1239 2141 1240
rect 2135 1238 2136 1239
rect 1862 1236 1868 1237
rect 2117 1236 2136 1238
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 110 1230 116 1231
rect 1590 1235 1596 1236
rect 1590 1231 1591 1235
rect 1595 1234 1596 1235
rect 1822 1235 1828 1236
rect 1595 1232 1601 1234
rect 1595 1231 1596 1232
rect 1590 1230 1596 1231
rect 1822 1231 1823 1235
rect 1827 1231 1828 1235
rect 1862 1232 1863 1236
rect 1867 1232 1868 1236
rect 2135 1235 2136 1236
rect 2140 1235 2141 1239
rect 2135 1234 2141 1235
rect 2210 1239 2216 1240
rect 2210 1235 2211 1239
rect 2215 1238 2216 1239
rect 2327 1239 2333 1240
rect 2215 1236 2265 1238
rect 2215 1235 2216 1236
rect 2210 1234 2216 1235
rect 2327 1235 2328 1239
rect 2332 1238 2333 1239
rect 2402 1239 2408 1240
rect 2332 1236 2361 1238
rect 2332 1235 2333 1236
rect 2327 1234 2333 1235
rect 2402 1235 2403 1239
rect 2407 1238 2408 1239
rect 2679 1239 2685 1240
rect 2679 1238 2680 1239
rect 2407 1236 2457 1238
rect 2613 1236 2680 1238
rect 2407 1235 2408 1236
rect 2402 1234 2408 1235
rect 2679 1235 2680 1236
rect 2684 1235 2685 1239
rect 2847 1239 2853 1240
rect 2847 1238 2848 1239
rect 2749 1236 2848 1238
rect 2679 1234 2685 1235
rect 2847 1235 2848 1236
rect 2852 1235 2853 1239
rect 3031 1239 3037 1240
rect 3031 1238 3032 1239
rect 2917 1236 3032 1238
rect 2847 1234 2853 1235
rect 3031 1235 3032 1236
rect 3036 1235 3037 1239
rect 3223 1239 3229 1240
rect 3223 1238 3224 1239
rect 3101 1236 3224 1238
rect 3031 1234 3037 1235
rect 3223 1235 3224 1236
rect 3228 1235 3229 1239
rect 3498 1239 3504 1240
rect 3498 1238 3499 1239
rect 3493 1236 3499 1238
rect 3223 1234 3229 1235
rect 3498 1235 3499 1236
rect 3503 1235 3504 1239
rect 3498 1234 3504 1235
rect 3574 1236 3580 1237
rect 1862 1231 1868 1232
rect 3574 1232 3575 1236
rect 3579 1232 3580 1236
rect 3574 1231 3580 1232
rect 1822 1230 1828 1231
rect 206 1225 212 1226
rect 206 1221 207 1225
rect 211 1221 212 1225
rect 206 1220 212 1221
rect 350 1225 356 1226
rect 350 1221 351 1225
rect 355 1221 356 1225
rect 350 1220 356 1221
rect 510 1225 516 1226
rect 510 1221 511 1225
rect 515 1221 516 1225
rect 510 1220 516 1221
rect 670 1225 676 1226
rect 670 1221 671 1225
rect 675 1221 676 1225
rect 670 1220 676 1221
rect 830 1225 836 1226
rect 830 1221 831 1225
rect 835 1221 836 1225
rect 830 1220 836 1221
rect 990 1225 996 1226
rect 990 1221 991 1225
rect 995 1221 996 1225
rect 990 1220 996 1221
rect 1142 1225 1148 1226
rect 1142 1221 1143 1225
rect 1147 1221 1148 1225
rect 1142 1220 1148 1221
rect 1286 1225 1292 1226
rect 1286 1221 1287 1225
rect 1291 1221 1292 1225
rect 1286 1220 1292 1221
rect 1430 1225 1436 1226
rect 1430 1221 1431 1225
rect 1435 1221 1436 1225
rect 1430 1220 1436 1221
rect 1582 1225 1588 1226
rect 1582 1221 1583 1225
rect 1587 1221 1588 1225
rect 1582 1220 1588 1221
rect 2062 1223 2068 1224
rect 2062 1219 2063 1223
rect 2067 1219 2068 1223
rect 2062 1218 2068 1219
rect 2150 1223 2156 1224
rect 2150 1219 2151 1223
rect 2155 1219 2156 1223
rect 2150 1218 2156 1219
rect 2246 1223 2252 1224
rect 2246 1219 2247 1223
rect 2251 1219 2252 1223
rect 2246 1218 2252 1219
rect 2342 1223 2348 1224
rect 2342 1219 2343 1223
rect 2347 1219 2348 1223
rect 2342 1218 2348 1219
rect 2438 1223 2444 1224
rect 2438 1219 2439 1223
rect 2443 1219 2444 1223
rect 2438 1218 2444 1219
rect 2558 1223 2564 1224
rect 2558 1219 2559 1223
rect 2563 1219 2564 1223
rect 2558 1218 2564 1219
rect 2694 1223 2700 1224
rect 2694 1219 2695 1223
rect 2699 1219 2700 1223
rect 2694 1218 2700 1219
rect 2862 1223 2868 1224
rect 2862 1219 2863 1223
rect 2867 1219 2868 1223
rect 2862 1218 2868 1219
rect 3046 1223 3052 1224
rect 3046 1219 3047 1223
rect 3051 1219 3052 1223
rect 3046 1218 3052 1219
rect 3238 1223 3244 1224
rect 3238 1219 3239 1223
rect 3243 1219 3244 1223
rect 3238 1218 3244 1219
rect 3438 1223 3444 1224
rect 3438 1219 3439 1223
rect 3443 1219 3444 1223
rect 3438 1218 3444 1219
rect 2055 1211 2061 1212
rect 2055 1207 2056 1211
rect 2060 1210 2061 1211
rect 2122 1211 2128 1212
rect 2122 1210 2123 1211
rect 2060 1208 2123 1210
rect 2060 1207 2061 1208
rect 2055 1206 2061 1207
rect 2122 1207 2123 1208
rect 2127 1207 2128 1211
rect 2122 1206 2128 1207
rect 2143 1211 2149 1212
rect 2143 1207 2144 1211
rect 2148 1210 2149 1211
rect 2210 1211 2216 1212
rect 2210 1210 2211 1211
rect 2148 1208 2211 1210
rect 2148 1207 2149 1208
rect 2143 1206 2149 1207
rect 2210 1207 2211 1208
rect 2215 1207 2216 1211
rect 2210 1206 2216 1207
rect 2239 1211 2245 1212
rect 2239 1207 2240 1211
rect 2244 1210 2245 1211
rect 2327 1211 2333 1212
rect 2327 1210 2328 1211
rect 2244 1208 2328 1210
rect 2244 1207 2245 1208
rect 2239 1206 2245 1207
rect 2327 1207 2328 1208
rect 2332 1207 2333 1211
rect 2327 1206 2333 1207
rect 2335 1211 2341 1212
rect 2335 1207 2336 1211
rect 2340 1210 2341 1211
rect 2402 1211 2408 1212
rect 2402 1210 2403 1211
rect 2340 1208 2403 1210
rect 2340 1207 2341 1208
rect 2335 1206 2341 1207
rect 2402 1207 2403 1208
rect 2407 1207 2408 1211
rect 2402 1206 2408 1207
rect 2431 1211 2437 1212
rect 2431 1207 2432 1211
rect 2436 1210 2437 1211
rect 2474 1211 2480 1212
rect 2474 1210 2475 1211
rect 2436 1208 2475 1210
rect 2436 1207 2437 1208
rect 2431 1206 2437 1207
rect 2474 1207 2475 1208
rect 2479 1207 2480 1211
rect 2474 1206 2480 1207
rect 2551 1211 2557 1212
rect 2551 1207 2552 1211
rect 2556 1210 2557 1211
rect 2566 1211 2572 1212
rect 2566 1210 2567 1211
rect 2556 1208 2567 1210
rect 2556 1207 2557 1208
rect 2551 1206 2557 1207
rect 2566 1207 2567 1208
rect 2571 1207 2572 1211
rect 2566 1206 2572 1207
rect 2679 1211 2685 1212
rect 2679 1207 2680 1211
rect 2684 1210 2685 1211
rect 2687 1211 2693 1212
rect 2687 1210 2688 1211
rect 2684 1208 2688 1210
rect 2684 1207 2685 1208
rect 2679 1206 2685 1207
rect 2687 1207 2688 1208
rect 2692 1207 2693 1211
rect 2687 1206 2693 1207
rect 2847 1211 2853 1212
rect 2847 1207 2848 1211
rect 2852 1210 2853 1211
rect 2855 1211 2861 1212
rect 2855 1210 2856 1211
rect 2852 1208 2856 1210
rect 2852 1207 2853 1208
rect 2847 1206 2853 1207
rect 2855 1207 2856 1208
rect 2860 1207 2861 1211
rect 2855 1206 2861 1207
rect 3031 1211 3037 1212
rect 3031 1207 3032 1211
rect 3036 1210 3037 1211
rect 3039 1211 3045 1212
rect 3039 1210 3040 1211
rect 3036 1208 3040 1210
rect 3036 1207 3037 1208
rect 3031 1206 3037 1207
rect 3039 1207 3040 1208
rect 3044 1207 3045 1211
rect 3039 1206 3045 1207
rect 3223 1211 3229 1212
rect 3223 1207 3224 1211
rect 3228 1210 3229 1211
rect 3231 1211 3237 1212
rect 3231 1210 3232 1211
rect 3228 1208 3232 1210
rect 3228 1207 3229 1208
rect 3223 1206 3229 1207
rect 3231 1207 3232 1208
rect 3236 1207 3237 1211
rect 3231 1206 3237 1207
rect 3431 1211 3437 1212
rect 3431 1207 3432 1211
rect 3436 1210 3437 1211
rect 3454 1211 3460 1212
rect 3454 1210 3455 1211
rect 3436 1208 3455 1210
rect 3436 1207 3437 1208
rect 3431 1206 3437 1207
rect 3454 1207 3455 1208
rect 3459 1207 3460 1211
rect 3454 1206 3460 1207
rect 2223 1203 2229 1204
rect 2223 1202 2224 1203
rect 2128 1200 2224 1202
rect 134 1195 140 1196
rect 134 1191 135 1195
rect 139 1191 140 1195
rect 134 1190 140 1191
rect 270 1195 276 1196
rect 270 1191 271 1195
rect 275 1191 276 1195
rect 270 1190 276 1191
rect 422 1195 428 1196
rect 422 1191 423 1195
rect 427 1191 428 1195
rect 422 1190 428 1191
rect 574 1195 580 1196
rect 574 1191 575 1195
rect 579 1191 580 1195
rect 574 1190 580 1191
rect 726 1195 732 1196
rect 726 1191 727 1195
rect 731 1191 732 1195
rect 726 1190 732 1191
rect 886 1195 892 1196
rect 886 1191 887 1195
rect 891 1191 892 1195
rect 886 1190 892 1191
rect 1054 1195 1060 1196
rect 1054 1191 1055 1195
rect 1059 1191 1060 1195
rect 1054 1190 1060 1191
rect 1230 1195 1236 1196
rect 1230 1191 1231 1195
rect 1235 1191 1236 1195
rect 1230 1190 1236 1191
rect 1414 1195 1420 1196
rect 1414 1191 1415 1195
rect 1419 1191 1420 1195
rect 1414 1190 1420 1191
rect 1598 1195 1604 1196
rect 1598 1191 1599 1195
rect 1603 1191 1604 1195
rect 1598 1190 1604 1191
rect 2031 1195 2037 1196
rect 2031 1191 2032 1195
rect 2036 1194 2037 1195
rect 2128 1194 2130 1200
rect 2223 1199 2224 1200
rect 2228 1199 2229 1203
rect 2223 1198 2229 1199
rect 2036 1192 2130 1194
rect 2135 1195 2141 1196
rect 2036 1191 2037 1192
rect 2031 1190 2037 1191
rect 2135 1191 2136 1195
rect 2140 1194 2141 1195
rect 2143 1195 2149 1196
rect 2143 1194 2144 1195
rect 2140 1192 2144 1194
rect 2140 1191 2141 1192
rect 2135 1190 2141 1191
rect 2143 1191 2144 1192
rect 2148 1191 2149 1195
rect 2143 1190 2149 1191
rect 2215 1195 2221 1196
rect 2215 1191 2216 1195
rect 2220 1194 2221 1195
rect 2271 1195 2277 1196
rect 2271 1194 2272 1195
rect 2220 1192 2272 1194
rect 2220 1191 2221 1192
rect 2215 1190 2221 1191
rect 2271 1191 2272 1192
rect 2276 1191 2277 1195
rect 2271 1190 2277 1191
rect 2407 1195 2413 1196
rect 2407 1191 2408 1195
rect 2412 1194 2413 1195
rect 2482 1195 2488 1196
rect 2482 1194 2483 1195
rect 2412 1192 2483 1194
rect 2412 1191 2413 1192
rect 2407 1190 2413 1191
rect 2482 1191 2483 1192
rect 2487 1191 2488 1195
rect 2482 1190 2488 1191
rect 2542 1195 2548 1196
rect 2542 1191 2543 1195
rect 2547 1194 2548 1195
rect 2551 1195 2557 1196
rect 2551 1194 2552 1195
rect 2547 1192 2552 1194
rect 2547 1191 2548 1192
rect 2542 1190 2548 1191
rect 2551 1191 2552 1192
rect 2556 1191 2557 1195
rect 2551 1190 2557 1191
rect 2703 1195 2709 1196
rect 2703 1191 2704 1195
rect 2708 1194 2709 1195
rect 2778 1195 2784 1196
rect 2778 1194 2779 1195
rect 2708 1192 2779 1194
rect 2708 1191 2709 1192
rect 2703 1190 2709 1191
rect 2778 1191 2779 1192
rect 2783 1191 2784 1195
rect 2778 1190 2784 1191
rect 2855 1195 2861 1196
rect 2855 1191 2856 1195
rect 2860 1194 2861 1195
rect 2934 1195 2940 1196
rect 2934 1194 2935 1195
rect 2860 1192 2935 1194
rect 2860 1191 2861 1192
rect 2855 1190 2861 1191
rect 2934 1191 2935 1192
rect 2939 1191 2940 1195
rect 2934 1190 2940 1191
rect 3007 1195 3013 1196
rect 3007 1191 3008 1195
rect 3012 1194 3013 1195
rect 3106 1195 3112 1196
rect 3106 1194 3107 1195
rect 3012 1192 3107 1194
rect 3012 1191 3013 1192
rect 3007 1190 3013 1191
rect 3106 1191 3107 1192
rect 3111 1191 3112 1195
rect 3106 1190 3112 1191
rect 3159 1195 3165 1196
rect 3159 1191 3160 1195
rect 3164 1194 3165 1195
rect 3246 1195 3252 1196
rect 3246 1194 3247 1195
rect 3164 1192 3247 1194
rect 3164 1191 3165 1192
rect 3159 1190 3165 1191
rect 3246 1191 3247 1192
rect 3251 1191 3252 1195
rect 3246 1190 3252 1191
rect 3311 1195 3317 1196
rect 3311 1191 3312 1195
rect 3316 1194 3317 1195
rect 3319 1195 3325 1196
rect 3319 1194 3320 1195
rect 3316 1192 3320 1194
rect 3316 1191 3317 1192
rect 3311 1190 3317 1191
rect 3319 1191 3320 1192
rect 3324 1191 3325 1195
rect 3319 1190 3325 1191
rect 3479 1195 3485 1196
rect 3479 1191 3480 1195
rect 3484 1194 3485 1195
rect 3498 1195 3504 1196
rect 3498 1194 3499 1195
rect 3484 1192 3499 1194
rect 3484 1191 3485 1192
rect 3479 1190 3485 1191
rect 3498 1191 3499 1192
rect 3503 1191 3504 1195
rect 3498 1190 3504 1191
rect 202 1187 208 1188
rect 202 1186 203 1187
rect 110 1185 116 1186
rect 110 1181 111 1185
rect 115 1181 116 1185
rect 193 1184 203 1186
rect 202 1183 203 1184
rect 207 1183 208 1187
rect 202 1182 208 1183
rect 1822 1185 1828 1186
rect 110 1180 116 1181
rect 1822 1181 1823 1185
rect 1827 1181 1828 1185
rect 1822 1180 1828 1181
rect 2038 1185 2044 1186
rect 2038 1181 2039 1185
rect 2043 1181 2044 1185
rect 2038 1180 2044 1181
rect 2150 1185 2156 1186
rect 2150 1181 2151 1185
rect 2155 1181 2156 1185
rect 2150 1180 2156 1181
rect 2278 1185 2284 1186
rect 2278 1181 2279 1185
rect 2283 1181 2284 1185
rect 2278 1180 2284 1181
rect 2414 1185 2420 1186
rect 2414 1181 2415 1185
rect 2419 1181 2420 1185
rect 2414 1180 2420 1181
rect 2558 1185 2564 1186
rect 2558 1181 2559 1185
rect 2563 1181 2564 1185
rect 2558 1180 2564 1181
rect 2710 1185 2716 1186
rect 2710 1181 2711 1185
rect 2715 1181 2716 1185
rect 2710 1180 2716 1181
rect 2862 1185 2868 1186
rect 2862 1181 2863 1185
rect 2867 1181 2868 1185
rect 2862 1180 2868 1181
rect 3014 1185 3020 1186
rect 3014 1181 3015 1185
rect 3019 1181 3020 1185
rect 3014 1180 3020 1181
rect 3166 1185 3172 1186
rect 3166 1181 3167 1185
rect 3171 1181 3172 1185
rect 3166 1180 3172 1181
rect 3326 1185 3332 1186
rect 3326 1181 3327 1185
rect 3331 1181 3332 1185
rect 3326 1180 3332 1181
rect 3486 1185 3492 1186
rect 3486 1181 3487 1185
rect 3491 1181 3492 1185
rect 3486 1180 3492 1181
rect 3254 1175 3260 1176
rect 3254 1174 3255 1175
rect 1862 1172 1868 1173
rect 3220 1172 3255 1174
rect 202 1171 208 1172
rect 110 1168 116 1169
rect 110 1164 111 1168
rect 115 1164 116 1168
rect 202 1167 203 1171
rect 207 1170 208 1171
rect 338 1171 344 1172
rect 207 1168 297 1170
rect 207 1167 208 1168
rect 202 1166 208 1167
rect 338 1167 339 1171
rect 343 1170 344 1171
rect 654 1171 660 1172
rect 654 1170 655 1171
rect 343 1168 449 1170
rect 637 1168 655 1170
rect 343 1167 344 1168
rect 338 1166 344 1167
rect 654 1167 655 1168
rect 659 1167 660 1171
rect 654 1166 660 1167
rect 679 1171 685 1172
rect 679 1167 680 1171
rect 684 1170 685 1171
rect 794 1171 800 1172
rect 684 1168 753 1170
rect 684 1167 685 1168
rect 679 1166 685 1167
rect 794 1167 795 1171
rect 799 1170 800 1171
rect 954 1171 960 1172
rect 799 1168 913 1170
rect 799 1167 800 1168
rect 794 1166 800 1167
rect 954 1167 955 1171
rect 959 1170 960 1171
rect 1122 1171 1128 1172
rect 959 1168 1081 1170
rect 959 1167 960 1168
rect 954 1166 960 1167
rect 1122 1167 1123 1171
rect 1127 1170 1128 1171
rect 1391 1171 1397 1172
rect 1127 1168 1257 1170
rect 1127 1167 1128 1168
rect 1122 1166 1128 1167
rect 1391 1167 1392 1171
rect 1396 1170 1397 1171
rect 1538 1171 1544 1172
rect 1396 1168 1441 1170
rect 1396 1167 1397 1168
rect 1391 1166 1397 1167
rect 1538 1167 1539 1171
rect 1543 1170 1544 1171
rect 1543 1168 1625 1170
rect 1822 1168 1828 1169
rect 1543 1167 1544 1168
rect 1538 1166 1544 1167
rect 110 1163 116 1164
rect 1822 1164 1823 1168
rect 1827 1164 1828 1168
rect 1862 1168 1863 1172
rect 1867 1168 1868 1172
rect 2215 1171 2221 1172
rect 2215 1170 2216 1171
rect 2205 1168 2216 1170
rect 1862 1167 1868 1168
rect 2215 1167 2216 1168
rect 2220 1167 2221 1171
rect 2474 1171 2480 1172
rect 2474 1170 2475 1171
rect 2469 1168 2475 1170
rect 2215 1166 2221 1167
rect 2223 1167 2229 1168
rect 1822 1163 1828 1164
rect 2223 1163 2224 1167
rect 2228 1166 2229 1167
rect 2474 1167 2475 1168
rect 2479 1167 2480 1171
rect 3220 1169 3222 1172
rect 3254 1171 3255 1172
rect 3259 1171 3260 1175
rect 3254 1170 3260 1171
rect 3574 1172 3580 1173
rect 3574 1168 3575 1172
rect 3579 1168 3580 1172
rect 2474 1166 2480 1167
rect 2482 1167 2488 1168
rect 2228 1164 2297 1166
rect 2228 1163 2229 1164
rect 2223 1162 2229 1163
rect 2482 1163 2483 1167
rect 2487 1166 2488 1167
rect 2778 1167 2784 1168
rect 2487 1164 2577 1166
rect 2487 1163 2488 1164
rect 2482 1162 2488 1163
rect 2778 1163 2779 1167
rect 2783 1166 2784 1167
rect 2934 1167 2940 1168
rect 2783 1164 2881 1166
rect 2783 1163 2784 1164
rect 2778 1162 2784 1163
rect 2934 1163 2935 1167
rect 2939 1166 2940 1167
rect 3246 1167 3252 1168
rect 3574 1167 3580 1168
rect 2939 1164 3033 1166
rect 2939 1163 2940 1164
rect 2934 1162 2940 1163
rect 3246 1163 3247 1167
rect 3251 1166 3252 1167
rect 3251 1164 3345 1166
rect 3251 1163 3252 1164
rect 3246 1162 3252 1163
rect 142 1155 148 1156
rect 142 1151 143 1155
rect 147 1151 148 1155
rect 142 1150 148 1151
rect 278 1155 284 1156
rect 278 1151 279 1155
rect 283 1151 284 1155
rect 278 1150 284 1151
rect 430 1155 436 1156
rect 430 1151 431 1155
rect 435 1151 436 1155
rect 430 1150 436 1151
rect 582 1155 588 1156
rect 582 1151 583 1155
rect 587 1151 588 1155
rect 582 1150 588 1151
rect 734 1155 740 1156
rect 734 1151 735 1155
rect 739 1151 740 1155
rect 734 1150 740 1151
rect 894 1155 900 1156
rect 894 1151 895 1155
rect 899 1151 900 1155
rect 894 1150 900 1151
rect 1062 1155 1068 1156
rect 1062 1151 1063 1155
rect 1067 1151 1068 1155
rect 1062 1150 1068 1151
rect 1238 1155 1244 1156
rect 1238 1151 1239 1155
rect 1243 1151 1244 1155
rect 1238 1150 1244 1151
rect 1422 1155 1428 1156
rect 1422 1151 1423 1155
rect 1427 1151 1428 1155
rect 1422 1150 1428 1151
rect 1606 1155 1612 1156
rect 1606 1151 1607 1155
rect 1611 1151 1612 1155
rect 1606 1150 1612 1151
rect 1862 1155 1868 1156
rect 1862 1151 1863 1155
rect 1867 1151 1868 1155
rect 1862 1150 1868 1151
rect 1958 1155 1964 1156
rect 1958 1151 1959 1155
rect 1963 1154 1964 1155
rect 2710 1155 2716 1156
rect 1963 1152 2049 1154
rect 1963 1151 1964 1152
rect 1958 1150 1964 1151
rect 2710 1151 2711 1155
rect 2715 1154 2716 1155
rect 3471 1155 3477 1156
rect 2715 1152 2721 1154
rect 2715 1151 2716 1152
rect 2710 1150 2716 1151
rect 3471 1151 3472 1155
rect 3476 1154 3477 1155
rect 3574 1155 3580 1156
rect 3476 1152 3497 1154
rect 3476 1151 3477 1152
rect 3471 1150 3477 1151
rect 3574 1151 3575 1155
rect 3579 1151 3580 1155
rect 3574 1150 3580 1151
rect 2030 1145 2036 1146
rect 135 1143 141 1144
rect 135 1139 136 1143
rect 140 1142 141 1143
rect 202 1143 208 1144
rect 202 1142 203 1143
rect 140 1140 203 1142
rect 140 1139 141 1140
rect 135 1138 141 1139
rect 202 1139 203 1140
rect 207 1139 208 1143
rect 202 1138 208 1139
rect 271 1143 277 1144
rect 271 1139 272 1143
rect 276 1142 277 1143
rect 338 1143 344 1144
rect 338 1142 339 1143
rect 276 1140 339 1142
rect 276 1139 277 1140
rect 271 1138 277 1139
rect 338 1139 339 1140
rect 343 1139 344 1143
rect 338 1138 344 1139
rect 359 1143 365 1144
rect 359 1139 360 1143
rect 364 1142 365 1143
rect 423 1143 429 1144
rect 423 1142 424 1143
rect 364 1140 424 1142
rect 364 1139 365 1140
rect 359 1138 365 1139
rect 423 1139 424 1140
rect 428 1139 429 1143
rect 423 1138 429 1139
rect 575 1143 581 1144
rect 575 1139 576 1143
rect 580 1142 581 1143
rect 679 1143 685 1144
rect 679 1142 680 1143
rect 580 1140 680 1142
rect 580 1139 581 1140
rect 575 1138 581 1139
rect 679 1139 680 1140
rect 684 1139 685 1143
rect 679 1138 685 1139
rect 727 1143 733 1144
rect 727 1139 728 1143
rect 732 1142 733 1143
rect 794 1143 800 1144
rect 794 1142 795 1143
rect 732 1140 795 1142
rect 732 1139 733 1140
rect 727 1138 733 1139
rect 794 1139 795 1140
rect 799 1139 800 1143
rect 794 1138 800 1139
rect 887 1143 893 1144
rect 887 1139 888 1143
rect 892 1142 893 1143
rect 954 1143 960 1144
rect 954 1142 955 1143
rect 892 1140 955 1142
rect 892 1139 893 1140
rect 887 1138 893 1139
rect 954 1139 955 1140
rect 959 1139 960 1143
rect 954 1138 960 1139
rect 1055 1143 1061 1144
rect 1055 1139 1056 1143
rect 1060 1142 1061 1143
rect 1122 1143 1128 1144
rect 1122 1142 1123 1143
rect 1060 1140 1123 1142
rect 1060 1139 1061 1140
rect 1055 1138 1061 1139
rect 1122 1139 1123 1140
rect 1127 1139 1128 1143
rect 1122 1138 1128 1139
rect 1231 1143 1237 1144
rect 1231 1139 1232 1143
rect 1236 1142 1237 1143
rect 1266 1143 1272 1144
rect 1266 1142 1267 1143
rect 1236 1140 1267 1142
rect 1236 1139 1237 1140
rect 1231 1138 1237 1139
rect 1266 1139 1267 1140
rect 1271 1139 1272 1143
rect 1266 1138 1272 1139
rect 1415 1143 1421 1144
rect 1415 1139 1416 1143
rect 1420 1142 1421 1143
rect 1538 1143 1544 1144
rect 1538 1142 1539 1143
rect 1420 1140 1539 1142
rect 1420 1139 1421 1140
rect 1415 1138 1421 1139
rect 1538 1139 1539 1140
rect 1543 1139 1544 1143
rect 1538 1138 1544 1139
rect 1590 1143 1596 1144
rect 1590 1139 1591 1143
rect 1595 1142 1596 1143
rect 1599 1143 1605 1144
rect 1599 1142 1600 1143
rect 1595 1140 1600 1142
rect 1595 1139 1596 1140
rect 1590 1138 1596 1139
rect 1599 1139 1600 1140
rect 1604 1139 1605 1143
rect 2030 1141 2031 1145
rect 2035 1141 2036 1145
rect 2030 1140 2036 1141
rect 2142 1145 2148 1146
rect 2142 1141 2143 1145
rect 2147 1141 2148 1145
rect 2142 1140 2148 1141
rect 2270 1145 2276 1146
rect 2270 1141 2271 1145
rect 2275 1141 2276 1145
rect 2270 1140 2276 1141
rect 2406 1145 2412 1146
rect 2406 1141 2407 1145
rect 2411 1141 2412 1145
rect 2406 1140 2412 1141
rect 2550 1145 2556 1146
rect 2550 1141 2551 1145
rect 2555 1141 2556 1145
rect 2550 1140 2556 1141
rect 2702 1145 2708 1146
rect 2702 1141 2703 1145
rect 2707 1141 2708 1145
rect 2702 1140 2708 1141
rect 2854 1145 2860 1146
rect 2854 1141 2855 1145
rect 2859 1141 2860 1145
rect 2854 1140 2860 1141
rect 3006 1145 3012 1146
rect 3006 1141 3007 1145
rect 3011 1141 3012 1145
rect 3006 1140 3012 1141
rect 3158 1145 3164 1146
rect 3158 1141 3159 1145
rect 3163 1141 3164 1145
rect 3158 1140 3164 1141
rect 3318 1145 3324 1146
rect 3318 1141 3319 1145
rect 3323 1141 3324 1145
rect 3318 1140 3324 1141
rect 3478 1145 3484 1146
rect 3478 1141 3479 1145
rect 3483 1141 3484 1145
rect 3478 1140 3484 1141
rect 1599 1138 1605 1139
rect 127 1131 133 1132
rect 127 1127 128 1131
rect 132 1130 133 1131
rect 135 1131 141 1132
rect 135 1130 136 1131
rect 132 1128 136 1130
rect 132 1127 133 1128
rect 127 1126 133 1127
rect 135 1127 136 1128
rect 140 1127 141 1131
rect 135 1126 141 1127
rect 215 1131 221 1132
rect 215 1127 216 1131
rect 220 1130 221 1131
rect 287 1131 293 1132
rect 287 1130 288 1131
rect 220 1128 288 1130
rect 220 1127 221 1128
rect 215 1126 221 1127
rect 287 1127 288 1128
rect 292 1127 293 1131
rect 287 1126 293 1127
rect 471 1131 477 1132
rect 471 1127 472 1131
rect 476 1130 477 1131
rect 594 1131 600 1132
rect 594 1130 595 1131
rect 476 1128 595 1130
rect 476 1127 477 1128
rect 471 1126 477 1127
rect 594 1127 595 1128
rect 599 1127 600 1131
rect 594 1126 600 1127
rect 654 1131 661 1132
rect 654 1127 655 1131
rect 660 1127 661 1131
rect 654 1126 661 1127
rect 751 1131 757 1132
rect 751 1127 752 1131
rect 756 1130 757 1131
rect 839 1131 845 1132
rect 839 1130 840 1131
rect 756 1128 840 1130
rect 756 1127 757 1128
rect 751 1126 757 1127
rect 839 1127 840 1128
rect 844 1127 845 1131
rect 839 1126 845 1127
rect 966 1131 972 1132
rect 966 1127 967 1131
rect 971 1130 972 1131
rect 1023 1131 1029 1132
rect 1023 1130 1024 1131
rect 971 1128 1024 1130
rect 971 1127 972 1128
rect 966 1126 972 1127
rect 1023 1127 1024 1128
rect 1028 1127 1029 1131
rect 1023 1126 1029 1127
rect 1119 1131 1125 1132
rect 1119 1127 1120 1131
rect 1124 1130 1125 1131
rect 1199 1131 1205 1132
rect 1199 1130 1200 1131
rect 1124 1128 1200 1130
rect 1124 1127 1125 1128
rect 1119 1126 1125 1127
rect 1199 1127 1200 1128
rect 1204 1127 1205 1131
rect 1199 1126 1205 1127
rect 1383 1131 1389 1132
rect 1383 1127 1384 1131
rect 1388 1130 1389 1131
rect 1391 1131 1397 1132
rect 1391 1130 1392 1131
rect 1388 1128 1392 1130
rect 1388 1127 1389 1128
rect 1383 1126 1389 1127
rect 1391 1127 1392 1128
rect 1396 1127 1397 1131
rect 1391 1126 1397 1127
rect 1495 1131 1501 1132
rect 1495 1127 1496 1131
rect 1500 1130 1501 1131
rect 1567 1131 1573 1132
rect 1567 1130 1568 1131
rect 1500 1128 1568 1130
rect 1500 1127 1501 1128
rect 1495 1126 1501 1127
rect 1567 1127 1568 1128
rect 1572 1127 1573 1131
rect 1567 1126 1573 1127
rect 1655 1131 1661 1132
rect 1655 1127 1656 1131
rect 1660 1130 1661 1131
rect 1727 1131 1733 1132
rect 1727 1130 1728 1131
rect 1660 1128 1728 1130
rect 1660 1127 1661 1128
rect 1655 1126 1661 1127
rect 1727 1127 1728 1128
rect 1732 1127 1733 1131
rect 1727 1126 1733 1127
rect 142 1121 148 1122
rect 142 1117 143 1121
rect 147 1117 148 1121
rect 142 1116 148 1117
rect 294 1121 300 1122
rect 294 1117 295 1121
rect 299 1117 300 1121
rect 294 1116 300 1117
rect 478 1121 484 1122
rect 478 1117 479 1121
rect 483 1117 484 1121
rect 478 1116 484 1117
rect 662 1121 668 1122
rect 662 1117 663 1121
rect 667 1117 668 1121
rect 662 1116 668 1117
rect 846 1121 852 1122
rect 846 1117 847 1121
rect 851 1117 852 1121
rect 846 1116 852 1117
rect 1030 1121 1036 1122
rect 1030 1117 1031 1121
rect 1035 1117 1036 1121
rect 1030 1116 1036 1117
rect 1206 1121 1212 1122
rect 1206 1117 1207 1121
rect 1211 1117 1212 1121
rect 1206 1116 1212 1117
rect 1390 1121 1396 1122
rect 1390 1117 1391 1121
rect 1395 1117 1396 1121
rect 1390 1116 1396 1117
rect 1574 1121 1580 1122
rect 1574 1117 1575 1121
rect 1579 1117 1580 1121
rect 1574 1116 1580 1117
rect 1734 1121 1740 1122
rect 1734 1117 1735 1121
rect 1739 1117 1740 1121
rect 1734 1116 1740 1117
rect 1942 1111 1948 1112
rect 110 1108 116 1109
rect 1822 1108 1828 1109
rect 110 1104 111 1108
rect 115 1104 116 1108
rect 215 1107 221 1108
rect 215 1106 216 1107
rect 197 1104 216 1106
rect 110 1103 116 1104
rect 215 1103 216 1104
rect 220 1103 221 1107
rect 359 1107 365 1108
rect 359 1106 360 1107
rect 349 1104 360 1106
rect 215 1102 221 1103
rect 359 1103 360 1104
rect 364 1103 365 1107
rect 751 1107 757 1108
rect 751 1106 752 1107
rect 717 1104 752 1106
rect 359 1102 365 1103
rect 751 1103 752 1104
rect 756 1103 757 1107
rect 1119 1107 1125 1108
rect 1119 1106 1120 1107
rect 1085 1104 1120 1106
rect 751 1102 757 1103
rect 1119 1103 1120 1104
rect 1124 1103 1125 1107
rect 1266 1107 1272 1108
rect 1266 1106 1267 1107
rect 1261 1104 1267 1106
rect 1119 1102 1125 1103
rect 1266 1103 1267 1104
rect 1271 1103 1272 1107
rect 1495 1107 1501 1108
rect 1495 1106 1496 1107
rect 1445 1104 1496 1106
rect 1266 1102 1272 1103
rect 1495 1103 1496 1104
rect 1500 1103 1501 1107
rect 1655 1107 1661 1108
rect 1655 1106 1656 1107
rect 1629 1104 1656 1106
rect 1495 1102 1501 1103
rect 1655 1103 1656 1104
rect 1660 1103 1661 1107
rect 1822 1104 1823 1108
rect 1827 1104 1828 1108
rect 1942 1107 1943 1111
rect 1947 1107 1948 1111
rect 1942 1106 1948 1107
rect 2086 1111 2092 1112
rect 2086 1107 2087 1111
rect 2091 1107 2092 1111
rect 2086 1106 2092 1107
rect 2230 1111 2236 1112
rect 2230 1107 2231 1111
rect 2235 1107 2236 1111
rect 2230 1106 2236 1107
rect 2382 1111 2388 1112
rect 2382 1107 2383 1111
rect 2387 1107 2388 1111
rect 2382 1106 2388 1107
rect 2534 1111 2540 1112
rect 2534 1107 2535 1111
rect 2539 1107 2540 1111
rect 2534 1106 2540 1107
rect 2686 1111 2692 1112
rect 2686 1107 2687 1111
rect 2691 1107 2692 1111
rect 2686 1106 2692 1107
rect 2838 1111 2844 1112
rect 2838 1107 2839 1111
rect 2843 1107 2844 1111
rect 2838 1106 2844 1107
rect 2990 1111 2996 1112
rect 2990 1107 2991 1111
rect 2995 1107 2996 1111
rect 2990 1106 2996 1107
rect 3150 1111 3156 1112
rect 3150 1107 3151 1111
rect 3155 1107 3156 1111
rect 3150 1106 3156 1107
rect 3318 1111 3324 1112
rect 3318 1107 3319 1111
rect 3323 1107 3324 1111
rect 3318 1106 3324 1107
rect 3478 1111 3484 1112
rect 3478 1107 3479 1111
rect 3483 1107 3484 1111
rect 3478 1106 3484 1107
rect 1822 1103 1828 1104
rect 2154 1103 2160 1104
rect 1655 1102 1661 1103
rect 1862 1101 1868 1102
rect 1862 1097 1863 1101
rect 1867 1097 1868 1101
rect 2154 1099 2155 1103
rect 2159 1102 2160 1103
rect 3078 1103 3084 1104
rect 2159 1100 2249 1102
rect 2544 1100 2553 1102
rect 2159 1099 2160 1100
rect 2154 1098 2160 1099
rect 2542 1099 2548 1100
rect 1862 1096 1868 1097
rect 2542 1095 2543 1099
rect 2547 1095 2548 1099
rect 3078 1099 3079 1103
rect 3083 1102 3084 1103
rect 3311 1103 3317 1104
rect 3083 1100 3169 1102
rect 3083 1099 3084 1100
rect 3078 1098 3084 1099
rect 3311 1099 3312 1103
rect 3316 1102 3317 1103
rect 3316 1100 3337 1102
rect 3574 1101 3580 1102
rect 3316 1099 3317 1100
rect 3311 1098 3317 1099
rect 3574 1097 3575 1101
rect 3579 1097 3580 1101
rect 3574 1096 3580 1097
rect 2542 1094 2548 1095
rect 110 1091 116 1092
rect 110 1087 111 1091
rect 115 1087 116 1091
rect 110 1086 116 1087
rect 362 1091 368 1092
rect 362 1087 363 1091
rect 367 1090 368 1091
rect 1719 1091 1725 1092
rect 367 1088 489 1090
rect 740 1088 857 1090
rect 367 1087 368 1088
rect 362 1086 368 1087
rect 134 1081 140 1082
rect 134 1077 135 1081
rect 139 1077 140 1081
rect 134 1076 140 1077
rect 286 1081 292 1082
rect 286 1077 287 1081
rect 291 1077 292 1081
rect 286 1076 292 1077
rect 470 1081 476 1082
rect 470 1077 471 1081
rect 475 1077 476 1081
rect 470 1076 476 1077
rect 654 1081 660 1082
rect 654 1077 655 1081
rect 659 1077 660 1081
rect 654 1076 660 1077
rect 594 1075 600 1076
rect 594 1071 595 1075
rect 599 1074 600 1075
rect 740 1074 742 1088
rect 1719 1087 1720 1091
rect 1724 1090 1725 1091
rect 1822 1091 1828 1092
rect 1724 1088 1745 1090
rect 1724 1087 1725 1088
rect 1719 1086 1725 1087
rect 1822 1087 1823 1091
rect 1827 1087 1828 1091
rect 1822 1086 1828 1087
rect 2079 1087 2085 1088
rect 2079 1086 2080 1087
rect 1862 1084 1868 1085
rect 2005 1084 2080 1086
rect 838 1081 844 1082
rect 838 1077 839 1081
rect 843 1077 844 1081
rect 838 1076 844 1077
rect 1022 1081 1028 1082
rect 1022 1077 1023 1081
rect 1027 1077 1028 1081
rect 1022 1076 1028 1077
rect 1198 1081 1204 1082
rect 1198 1077 1199 1081
rect 1203 1077 1204 1081
rect 1198 1076 1204 1077
rect 1382 1081 1388 1082
rect 1382 1077 1383 1081
rect 1387 1077 1388 1081
rect 1382 1076 1388 1077
rect 1566 1081 1572 1082
rect 1566 1077 1567 1081
rect 1571 1077 1572 1081
rect 1566 1076 1572 1077
rect 1726 1081 1732 1082
rect 1726 1077 1727 1081
rect 1731 1077 1732 1081
rect 1862 1080 1863 1084
rect 1867 1080 1868 1084
rect 2079 1083 2080 1084
rect 2084 1083 2085 1087
rect 2223 1087 2229 1088
rect 2223 1086 2224 1087
rect 2149 1084 2224 1086
rect 2079 1082 2085 1083
rect 2223 1083 2224 1084
rect 2228 1083 2229 1087
rect 2527 1087 2533 1088
rect 2527 1086 2528 1087
rect 2445 1084 2528 1086
rect 2223 1082 2229 1083
rect 2527 1083 2528 1084
rect 2532 1083 2533 1087
rect 2831 1087 2837 1088
rect 2831 1086 2832 1087
rect 2749 1084 2832 1086
rect 2527 1082 2533 1083
rect 2831 1083 2832 1084
rect 2836 1083 2837 1087
rect 2983 1087 2989 1088
rect 2983 1086 2984 1087
rect 2901 1084 2984 1086
rect 2831 1082 2837 1083
rect 2983 1083 2984 1084
rect 2988 1083 2989 1087
rect 3143 1087 3149 1088
rect 3143 1086 3144 1087
rect 3053 1084 3144 1086
rect 2983 1082 2989 1083
rect 3143 1083 3144 1084
rect 3148 1083 3149 1087
rect 3143 1082 3149 1083
rect 3470 1087 3476 1088
rect 3470 1083 3471 1087
rect 3475 1086 3476 1087
rect 3475 1084 3505 1086
rect 3574 1084 3580 1085
rect 3475 1083 3476 1084
rect 3470 1082 3476 1083
rect 1862 1079 1868 1080
rect 3574 1080 3575 1084
rect 3579 1080 3580 1084
rect 3574 1079 3580 1080
rect 1726 1076 1732 1077
rect 599 1072 742 1074
rect 599 1071 600 1072
rect 594 1070 600 1071
rect 1950 1071 1956 1072
rect 1950 1067 1951 1071
rect 1955 1067 1956 1071
rect 1950 1066 1956 1067
rect 2094 1071 2100 1072
rect 2094 1067 2095 1071
rect 2099 1067 2100 1071
rect 2094 1066 2100 1067
rect 2238 1071 2244 1072
rect 2238 1067 2239 1071
rect 2243 1067 2244 1071
rect 2238 1066 2244 1067
rect 2390 1071 2396 1072
rect 2390 1067 2391 1071
rect 2395 1067 2396 1071
rect 2390 1066 2396 1067
rect 2542 1071 2548 1072
rect 2542 1067 2543 1071
rect 2547 1067 2548 1071
rect 2542 1066 2548 1067
rect 2694 1071 2700 1072
rect 2694 1067 2695 1071
rect 2699 1067 2700 1071
rect 2694 1066 2700 1067
rect 2846 1071 2852 1072
rect 2846 1067 2847 1071
rect 2851 1067 2852 1071
rect 2846 1066 2852 1067
rect 2998 1071 3004 1072
rect 2998 1067 2999 1071
rect 3003 1067 3004 1071
rect 2998 1066 3004 1067
rect 3158 1071 3164 1072
rect 3158 1067 3159 1071
rect 3163 1067 3164 1071
rect 3158 1066 3164 1067
rect 3326 1071 3332 1072
rect 3326 1067 3327 1071
rect 3331 1067 3332 1071
rect 3326 1066 3332 1067
rect 3486 1071 3492 1072
rect 3486 1067 3487 1071
rect 3491 1067 3492 1071
rect 3486 1066 3492 1067
rect 134 1059 140 1060
rect 134 1055 135 1059
rect 139 1055 140 1059
rect 134 1054 140 1055
rect 270 1059 276 1060
rect 270 1055 271 1059
rect 275 1055 276 1059
rect 270 1054 276 1055
rect 430 1059 436 1060
rect 430 1055 431 1059
rect 435 1055 436 1059
rect 430 1054 436 1055
rect 582 1059 588 1060
rect 582 1055 583 1059
rect 587 1055 588 1059
rect 582 1054 588 1055
rect 734 1059 740 1060
rect 734 1055 735 1059
rect 739 1055 740 1059
rect 734 1054 740 1055
rect 886 1059 892 1060
rect 886 1055 887 1059
rect 891 1055 892 1059
rect 886 1054 892 1055
rect 1046 1059 1052 1060
rect 1046 1055 1047 1059
rect 1051 1055 1052 1059
rect 1046 1054 1052 1055
rect 1214 1059 1220 1060
rect 1214 1055 1215 1059
rect 1219 1055 1220 1059
rect 1214 1054 1220 1055
rect 1382 1059 1388 1060
rect 1382 1055 1383 1059
rect 1387 1055 1388 1059
rect 1382 1054 1388 1055
rect 1558 1059 1564 1060
rect 1558 1055 1559 1059
rect 1563 1055 1564 1059
rect 1558 1054 1564 1055
rect 1726 1059 1732 1060
rect 1726 1055 1727 1059
rect 1731 1055 1732 1059
rect 1726 1054 1732 1055
rect 1943 1059 1949 1060
rect 1943 1055 1944 1059
rect 1948 1058 1949 1059
rect 1958 1059 1964 1060
rect 1958 1058 1959 1059
rect 1948 1056 1959 1058
rect 1948 1055 1949 1056
rect 1943 1054 1949 1055
rect 1958 1055 1959 1056
rect 1963 1055 1964 1059
rect 1958 1054 1964 1055
rect 2079 1059 2085 1060
rect 2079 1055 2080 1059
rect 2084 1058 2085 1059
rect 2087 1059 2093 1060
rect 2087 1058 2088 1059
rect 2084 1056 2088 1058
rect 2084 1055 2085 1056
rect 2079 1054 2085 1055
rect 2087 1055 2088 1056
rect 2092 1055 2093 1059
rect 2087 1054 2093 1055
rect 2223 1059 2229 1060
rect 2223 1055 2224 1059
rect 2228 1058 2229 1059
rect 2231 1059 2237 1060
rect 2231 1058 2232 1059
rect 2228 1056 2232 1058
rect 2228 1055 2229 1056
rect 2223 1054 2229 1055
rect 2231 1055 2232 1056
rect 2236 1055 2237 1059
rect 2231 1054 2237 1055
rect 2383 1059 2389 1060
rect 2383 1055 2384 1059
rect 2388 1058 2389 1059
rect 2391 1059 2397 1060
rect 2391 1058 2392 1059
rect 2388 1056 2392 1058
rect 2388 1055 2389 1056
rect 2383 1054 2389 1055
rect 2391 1055 2392 1056
rect 2396 1055 2397 1059
rect 2391 1054 2397 1055
rect 2527 1059 2533 1060
rect 2527 1055 2528 1059
rect 2532 1058 2533 1059
rect 2535 1059 2541 1060
rect 2535 1058 2536 1059
rect 2532 1056 2536 1058
rect 2532 1055 2533 1056
rect 2527 1054 2533 1055
rect 2535 1055 2536 1056
rect 2540 1055 2541 1059
rect 2535 1054 2541 1055
rect 2687 1059 2693 1060
rect 2687 1055 2688 1059
rect 2692 1058 2693 1059
rect 2710 1059 2716 1060
rect 2710 1058 2711 1059
rect 2692 1056 2711 1058
rect 2692 1055 2693 1056
rect 2687 1054 2693 1055
rect 2710 1055 2711 1056
rect 2715 1055 2716 1059
rect 2710 1054 2716 1055
rect 2831 1059 2837 1060
rect 2831 1055 2832 1059
rect 2836 1058 2837 1059
rect 2839 1059 2845 1060
rect 2839 1058 2840 1059
rect 2836 1056 2840 1058
rect 2836 1055 2837 1056
rect 2831 1054 2837 1055
rect 2839 1055 2840 1056
rect 2844 1055 2845 1059
rect 2839 1054 2845 1055
rect 2983 1059 2989 1060
rect 2983 1055 2984 1059
rect 2988 1058 2989 1059
rect 2991 1059 2997 1060
rect 2991 1058 2992 1059
rect 2988 1056 2992 1058
rect 2988 1055 2989 1056
rect 2983 1054 2989 1055
rect 2991 1055 2992 1056
rect 2996 1055 2997 1059
rect 2991 1054 2997 1055
rect 3143 1059 3149 1060
rect 3143 1055 3144 1059
rect 3148 1058 3149 1059
rect 3151 1059 3157 1060
rect 3151 1058 3152 1059
rect 3148 1056 3152 1058
rect 3148 1055 3149 1056
rect 3143 1054 3149 1055
rect 3151 1055 3152 1056
rect 3156 1055 3157 1059
rect 3151 1054 3157 1055
rect 3319 1059 3325 1060
rect 3319 1055 3320 1059
rect 3324 1058 3325 1059
rect 3327 1059 3333 1060
rect 3327 1058 3328 1059
rect 3324 1056 3328 1058
rect 3324 1055 3325 1056
rect 3319 1054 3325 1055
rect 3327 1055 3328 1056
rect 3332 1055 3333 1059
rect 3327 1054 3333 1055
rect 3471 1059 3477 1060
rect 3471 1055 3472 1059
rect 3476 1058 3477 1059
rect 3479 1059 3485 1060
rect 3479 1058 3480 1059
rect 3476 1056 3480 1058
rect 3476 1055 3477 1056
rect 3471 1054 3477 1055
rect 3479 1055 3480 1056
rect 3484 1055 3485 1059
rect 3479 1054 3485 1055
rect 127 1051 133 1052
rect 110 1049 116 1050
rect 110 1045 111 1049
rect 115 1045 116 1049
rect 127 1047 128 1051
rect 132 1050 133 1051
rect 966 1051 972 1052
rect 966 1050 967 1051
rect 132 1048 153 1050
rect 945 1048 967 1050
rect 132 1047 133 1048
rect 127 1046 133 1047
rect 966 1047 967 1048
rect 971 1047 972 1051
rect 966 1046 972 1047
rect 1282 1051 1288 1052
rect 1282 1047 1283 1051
rect 1287 1050 1288 1051
rect 1287 1048 1401 1050
rect 1822 1049 1828 1050
rect 1287 1047 1288 1048
rect 1282 1046 1288 1047
rect 110 1044 116 1045
rect 1822 1045 1823 1049
rect 1827 1045 1828 1049
rect 1822 1044 1828 1045
rect 423 1035 429 1036
rect 423 1034 424 1035
rect 110 1032 116 1033
rect 333 1032 424 1034
rect 110 1028 111 1032
rect 115 1028 116 1032
rect 423 1031 424 1032
rect 428 1031 429 1035
rect 575 1035 581 1036
rect 575 1034 576 1035
rect 493 1032 576 1034
rect 423 1030 429 1031
rect 575 1031 576 1032
rect 580 1031 581 1035
rect 727 1035 733 1036
rect 727 1034 728 1035
rect 645 1032 728 1034
rect 575 1030 581 1031
rect 727 1031 728 1032
rect 732 1031 733 1035
rect 814 1035 820 1036
rect 814 1034 815 1035
rect 797 1032 815 1034
rect 727 1030 733 1031
rect 814 1031 815 1032
rect 819 1031 820 1035
rect 814 1030 820 1031
rect 954 1035 960 1036
rect 954 1031 955 1035
rect 959 1034 960 1035
rect 1375 1035 1381 1036
rect 1375 1034 1376 1035
rect 959 1032 1073 1034
rect 1277 1032 1376 1034
rect 959 1031 960 1032
rect 954 1030 960 1031
rect 1375 1031 1376 1032
rect 1380 1031 1381 1035
rect 1646 1035 1652 1036
rect 1646 1034 1647 1035
rect 1621 1032 1647 1034
rect 1375 1030 1381 1031
rect 1646 1031 1647 1032
rect 1651 1031 1652 1035
rect 1646 1030 1652 1031
rect 1655 1035 1661 1036
rect 1655 1031 1656 1035
rect 1660 1034 1661 1035
rect 1911 1035 1917 1036
rect 1660 1032 1753 1034
rect 1822 1032 1828 1033
rect 1660 1031 1661 1032
rect 1655 1030 1661 1031
rect 110 1027 116 1028
rect 1822 1028 1823 1032
rect 1827 1028 1828 1032
rect 1911 1031 1912 1035
rect 1916 1034 1917 1035
rect 1986 1035 1992 1036
rect 1986 1034 1987 1035
rect 1916 1032 1987 1034
rect 1916 1031 1917 1032
rect 1911 1030 1917 1031
rect 1986 1031 1987 1032
rect 1991 1031 1992 1035
rect 1986 1030 1992 1031
rect 2119 1035 2125 1036
rect 2119 1031 2120 1035
rect 2124 1034 2125 1035
rect 2154 1035 2160 1036
rect 2154 1034 2155 1035
rect 2124 1032 2155 1034
rect 2124 1031 2125 1032
rect 2119 1030 2125 1031
rect 2154 1031 2155 1032
rect 2159 1031 2160 1035
rect 2154 1030 2160 1031
rect 2319 1035 2325 1036
rect 2319 1031 2320 1035
rect 2324 1034 2325 1035
rect 2423 1035 2429 1036
rect 2423 1034 2424 1035
rect 2324 1032 2424 1034
rect 2324 1031 2325 1032
rect 2319 1030 2325 1031
rect 2423 1031 2424 1032
rect 2428 1031 2429 1035
rect 2423 1030 2429 1031
rect 2511 1035 2517 1036
rect 2511 1031 2512 1035
rect 2516 1034 2517 1035
rect 2526 1035 2532 1036
rect 2526 1034 2527 1035
rect 2516 1032 2527 1034
rect 2516 1031 2517 1032
rect 2511 1030 2517 1031
rect 2526 1031 2527 1032
rect 2531 1031 2532 1035
rect 2526 1030 2532 1031
rect 2687 1035 2693 1036
rect 2687 1031 2688 1035
rect 2692 1034 2693 1035
rect 2702 1035 2708 1036
rect 2702 1034 2703 1035
rect 2692 1032 2703 1034
rect 2692 1031 2693 1032
rect 2687 1030 2693 1031
rect 2702 1031 2703 1032
rect 2707 1031 2708 1035
rect 2702 1030 2708 1031
rect 2775 1035 2781 1036
rect 2775 1031 2776 1035
rect 2780 1034 2781 1035
rect 2855 1035 2861 1036
rect 2855 1034 2856 1035
rect 2780 1032 2856 1034
rect 2780 1031 2781 1032
rect 2775 1030 2781 1031
rect 2855 1031 2856 1032
rect 2860 1031 2861 1035
rect 2855 1030 2861 1031
rect 2943 1035 2949 1036
rect 2943 1031 2944 1035
rect 2948 1034 2949 1035
rect 3015 1035 3021 1036
rect 3015 1034 3016 1035
rect 2948 1032 3016 1034
rect 2948 1031 2949 1032
rect 2943 1030 2949 1031
rect 3015 1031 3016 1032
rect 3020 1031 3021 1035
rect 3015 1030 3021 1031
rect 3087 1035 3093 1036
rect 3087 1031 3088 1035
rect 3092 1034 3093 1035
rect 3175 1035 3181 1036
rect 3175 1034 3176 1035
rect 3092 1032 3176 1034
rect 3092 1031 3093 1032
rect 3087 1030 3093 1031
rect 3175 1031 3176 1032
rect 3180 1031 3181 1035
rect 3175 1030 3181 1031
rect 3335 1035 3341 1036
rect 3335 1031 3336 1035
rect 3340 1034 3341 1035
rect 3350 1035 3356 1036
rect 3350 1034 3351 1035
rect 3340 1032 3351 1034
rect 3340 1031 3341 1032
rect 3335 1030 3341 1031
rect 3350 1031 3351 1032
rect 3355 1031 3356 1035
rect 3350 1030 3356 1031
rect 3470 1035 3476 1036
rect 3470 1031 3471 1035
rect 3475 1034 3476 1035
rect 3479 1035 3485 1036
rect 3479 1034 3480 1035
rect 3475 1032 3480 1034
rect 3475 1031 3476 1032
rect 3470 1030 3476 1031
rect 3479 1031 3480 1032
rect 3484 1031 3485 1035
rect 3479 1030 3485 1031
rect 1822 1027 1828 1028
rect 1918 1025 1924 1026
rect 1918 1021 1919 1025
rect 1923 1021 1924 1025
rect 1918 1020 1924 1021
rect 2126 1025 2132 1026
rect 2126 1021 2127 1025
rect 2131 1021 2132 1025
rect 2126 1020 2132 1021
rect 2326 1025 2332 1026
rect 2326 1021 2327 1025
rect 2331 1021 2332 1025
rect 2326 1020 2332 1021
rect 2518 1025 2524 1026
rect 2518 1021 2519 1025
rect 2523 1021 2524 1025
rect 2518 1020 2524 1021
rect 2694 1025 2700 1026
rect 2694 1021 2695 1025
rect 2699 1021 2700 1025
rect 2694 1020 2700 1021
rect 2862 1025 2868 1026
rect 2862 1021 2863 1025
rect 2867 1021 2868 1025
rect 2862 1020 2868 1021
rect 3022 1025 3028 1026
rect 3022 1021 3023 1025
rect 3027 1021 3028 1025
rect 3022 1020 3028 1021
rect 3182 1025 3188 1026
rect 3182 1021 3183 1025
rect 3187 1021 3188 1025
rect 3182 1020 3188 1021
rect 3342 1025 3348 1026
rect 3342 1021 3343 1025
rect 3347 1021 3348 1025
rect 3342 1020 3348 1021
rect 3486 1025 3492 1026
rect 3486 1021 3487 1025
rect 3491 1021 3492 1025
rect 3486 1020 3492 1021
rect 142 1019 148 1020
rect 142 1015 143 1019
rect 147 1015 148 1019
rect 142 1014 148 1015
rect 278 1019 284 1020
rect 278 1015 279 1019
rect 283 1015 284 1019
rect 278 1014 284 1015
rect 438 1019 444 1020
rect 438 1015 439 1019
rect 443 1015 444 1019
rect 438 1014 444 1015
rect 590 1019 596 1020
rect 590 1015 591 1019
rect 595 1015 596 1019
rect 590 1014 596 1015
rect 742 1019 748 1020
rect 742 1015 743 1019
rect 747 1015 748 1019
rect 742 1014 748 1015
rect 894 1019 900 1020
rect 894 1015 895 1019
rect 899 1015 900 1019
rect 894 1014 900 1015
rect 1054 1019 1060 1020
rect 1054 1015 1055 1019
rect 1059 1015 1060 1019
rect 1054 1014 1060 1015
rect 1222 1019 1228 1020
rect 1222 1015 1223 1019
rect 1227 1015 1228 1019
rect 1222 1014 1228 1015
rect 1390 1019 1396 1020
rect 1390 1015 1391 1019
rect 1395 1015 1396 1019
rect 1390 1014 1396 1015
rect 1566 1019 1572 1020
rect 1566 1015 1567 1019
rect 1571 1015 1572 1019
rect 1566 1014 1572 1015
rect 1734 1019 1740 1020
rect 1734 1015 1735 1019
rect 1739 1015 1740 1019
rect 1734 1014 1740 1015
rect 1862 1012 1868 1013
rect 3574 1012 3580 1013
rect 1862 1008 1863 1012
rect 1867 1008 1868 1012
rect 2391 1011 2397 1012
rect 2391 1010 2392 1011
rect 2381 1008 2392 1010
rect 135 1007 141 1008
rect 135 1003 136 1007
rect 140 1006 141 1007
rect 223 1007 229 1008
rect 223 1006 224 1007
rect 140 1004 224 1006
rect 140 1003 141 1004
rect 135 1002 141 1003
rect 223 1003 224 1004
rect 228 1003 229 1007
rect 223 1002 229 1003
rect 271 1007 277 1008
rect 271 1003 272 1007
rect 276 1006 277 1007
rect 362 1007 368 1008
rect 362 1006 363 1007
rect 276 1004 363 1006
rect 276 1003 277 1004
rect 271 1002 277 1003
rect 362 1003 363 1004
rect 367 1003 368 1007
rect 362 1002 368 1003
rect 423 1007 429 1008
rect 423 1003 424 1007
rect 428 1006 429 1007
rect 431 1007 437 1008
rect 431 1006 432 1007
rect 428 1004 432 1006
rect 428 1003 429 1004
rect 423 1002 429 1003
rect 431 1003 432 1004
rect 436 1003 437 1007
rect 431 1002 437 1003
rect 575 1007 581 1008
rect 575 1003 576 1007
rect 580 1006 581 1007
rect 583 1007 589 1008
rect 583 1006 584 1007
rect 580 1004 584 1006
rect 580 1003 581 1004
rect 575 1002 581 1003
rect 583 1003 584 1004
rect 588 1003 589 1007
rect 583 1002 589 1003
rect 727 1007 733 1008
rect 727 1003 728 1007
rect 732 1006 733 1007
rect 735 1007 741 1008
rect 735 1006 736 1007
rect 732 1004 736 1006
rect 732 1003 733 1004
rect 727 1002 733 1003
rect 735 1003 736 1004
rect 740 1003 741 1007
rect 735 1002 741 1003
rect 887 1007 893 1008
rect 887 1003 888 1007
rect 892 1006 893 1007
rect 954 1007 960 1008
rect 954 1006 955 1007
rect 892 1004 955 1006
rect 892 1003 893 1004
rect 887 1002 893 1003
rect 954 1003 955 1004
rect 959 1003 960 1007
rect 954 1002 960 1003
rect 1047 1007 1053 1008
rect 1047 1003 1048 1007
rect 1052 1006 1053 1007
rect 1062 1007 1068 1008
rect 1062 1006 1063 1007
rect 1052 1004 1063 1006
rect 1052 1003 1053 1004
rect 1047 1002 1053 1003
rect 1062 1003 1063 1004
rect 1067 1003 1068 1007
rect 1062 1002 1068 1003
rect 1215 1007 1221 1008
rect 1215 1003 1216 1007
rect 1220 1006 1221 1007
rect 1230 1007 1236 1008
rect 1230 1006 1231 1007
rect 1220 1004 1231 1006
rect 1220 1003 1221 1004
rect 1215 1002 1221 1003
rect 1230 1003 1231 1004
rect 1235 1003 1236 1007
rect 1230 1002 1236 1003
rect 1375 1007 1381 1008
rect 1375 1003 1376 1007
rect 1380 1006 1381 1007
rect 1383 1007 1389 1008
rect 1383 1006 1384 1007
rect 1380 1004 1384 1006
rect 1380 1003 1381 1004
rect 1375 1002 1381 1003
rect 1383 1003 1384 1004
rect 1388 1003 1389 1007
rect 1383 1002 1389 1003
rect 1559 1007 1565 1008
rect 1559 1003 1560 1007
rect 1564 1006 1565 1007
rect 1655 1007 1661 1008
rect 1655 1006 1656 1007
rect 1564 1004 1656 1006
rect 1564 1003 1565 1004
rect 1559 1002 1565 1003
rect 1655 1003 1656 1004
rect 1660 1003 1661 1007
rect 1655 1002 1661 1003
rect 1719 1007 1725 1008
rect 1719 1003 1720 1007
rect 1724 1006 1725 1007
rect 1727 1007 1733 1008
rect 1862 1007 1868 1008
rect 1986 1007 1992 1008
rect 1727 1006 1728 1007
rect 1724 1004 1728 1006
rect 1724 1003 1725 1004
rect 1719 1002 1725 1003
rect 1727 1003 1728 1004
rect 1732 1003 1733 1007
rect 1727 1002 1733 1003
rect 1986 1003 1987 1007
rect 1991 1006 1992 1007
rect 2391 1007 2392 1008
rect 2396 1007 2397 1011
rect 2775 1011 2781 1012
rect 2775 1010 2776 1011
rect 2749 1008 2776 1010
rect 2391 1006 2397 1007
rect 2423 1007 2429 1008
rect 1991 1004 2145 1006
rect 1991 1003 1992 1004
rect 1986 1002 1992 1003
rect 2423 1003 2424 1007
rect 2428 1006 2429 1007
rect 2775 1007 2776 1008
rect 2780 1007 2781 1011
rect 2943 1011 2949 1012
rect 2943 1010 2944 1011
rect 2917 1008 2944 1010
rect 2775 1006 2781 1007
rect 2943 1007 2944 1008
rect 2948 1007 2949 1011
rect 3087 1011 3093 1012
rect 3087 1010 3088 1011
rect 3077 1008 3088 1010
rect 2943 1006 2949 1007
rect 3087 1007 3088 1008
rect 3092 1007 3093 1011
rect 3574 1008 3575 1012
rect 3579 1008 3580 1012
rect 3087 1006 3093 1007
rect 3327 1007 3333 1008
rect 3574 1007 3580 1008
rect 2428 1004 2537 1006
rect 2428 1003 2429 1004
rect 2423 1002 2429 1003
rect 3327 1003 3328 1007
rect 3332 1006 3333 1007
rect 3332 1004 3361 1006
rect 3332 1003 3333 1004
rect 3327 1002 3333 1003
rect 1578 999 1584 1000
rect 1578 998 1579 999
rect 1388 996 1579 998
rect 127 991 133 992
rect 127 987 128 991
rect 132 990 133 991
rect 135 991 141 992
rect 135 990 136 991
rect 132 988 136 990
rect 132 987 133 988
rect 127 986 133 987
rect 135 987 136 988
rect 140 987 141 991
rect 135 986 141 987
rect 215 991 221 992
rect 215 987 216 991
rect 220 990 221 991
rect 279 991 285 992
rect 279 990 280 991
rect 220 988 280 990
rect 220 987 221 988
rect 215 986 221 987
rect 279 987 280 988
rect 284 987 285 991
rect 279 986 285 987
rect 455 991 461 992
rect 455 987 456 991
rect 460 990 461 991
rect 535 991 541 992
rect 535 990 536 991
rect 460 988 536 990
rect 460 987 461 988
rect 455 986 461 987
rect 535 987 536 988
rect 540 987 541 991
rect 535 986 541 987
rect 639 991 645 992
rect 639 987 640 991
rect 644 990 645 991
rect 727 991 733 992
rect 727 990 728 991
rect 644 988 728 990
rect 644 987 645 988
rect 639 986 645 987
rect 727 987 728 988
rect 732 987 733 991
rect 727 986 733 987
rect 814 991 821 992
rect 814 987 815 991
rect 820 987 821 991
rect 814 986 821 987
rect 991 991 997 992
rect 991 987 992 991
rect 996 990 997 991
rect 1006 991 1012 992
rect 1006 990 1007 991
rect 996 988 1007 990
rect 996 987 997 988
rect 991 986 997 987
rect 1006 987 1007 988
rect 1011 987 1012 991
rect 1006 986 1012 987
rect 1079 991 1085 992
rect 1079 987 1080 991
rect 1084 990 1085 991
rect 1159 991 1165 992
rect 1159 990 1160 991
rect 1084 988 1160 990
rect 1084 987 1085 988
rect 1079 986 1085 987
rect 1159 987 1160 988
rect 1164 987 1165 991
rect 1159 986 1165 987
rect 1319 991 1325 992
rect 1319 987 1320 991
rect 1324 990 1325 991
rect 1388 990 1390 996
rect 1578 995 1579 996
rect 1583 995 1584 999
rect 1578 994 1584 995
rect 1862 995 1868 996
rect 1324 988 1390 990
rect 1399 991 1405 992
rect 1324 987 1325 988
rect 1319 986 1325 987
rect 1399 987 1400 991
rect 1404 990 1405 991
rect 1479 991 1485 992
rect 1479 990 1480 991
rect 1404 988 1480 990
rect 1404 987 1405 988
rect 1399 986 1405 987
rect 1479 987 1480 988
rect 1484 987 1485 991
rect 1479 986 1485 987
rect 1646 991 1653 992
rect 1646 987 1647 991
rect 1652 987 1653 991
rect 1862 991 1863 995
rect 1867 991 1868 995
rect 1862 990 1868 991
rect 1902 995 1908 996
rect 1902 991 1903 995
rect 1907 994 1908 995
rect 3110 995 3116 996
rect 1907 992 1929 994
rect 1907 991 1908 992
rect 1902 990 1908 991
rect 3110 991 3111 995
rect 3115 994 3116 995
rect 3471 995 3477 996
rect 3115 992 3193 994
rect 3115 991 3116 992
rect 3110 990 3116 991
rect 3471 991 3472 995
rect 3476 994 3477 995
rect 3574 995 3580 996
rect 3476 992 3497 994
rect 3476 991 3477 992
rect 3471 990 3477 991
rect 3574 991 3575 995
rect 3579 991 3580 995
rect 3574 990 3580 991
rect 1646 986 1653 987
rect 1910 985 1916 986
rect 142 981 148 982
rect 142 977 143 981
rect 147 977 148 981
rect 142 976 148 977
rect 286 981 292 982
rect 286 977 287 981
rect 291 977 292 981
rect 286 976 292 977
rect 462 981 468 982
rect 462 977 463 981
rect 467 977 468 981
rect 462 976 468 977
rect 646 981 652 982
rect 646 977 647 981
rect 651 977 652 981
rect 646 976 652 977
rect 822 981 828 982
rect 822 977 823 981
rect 827 977 828 981
rect 822 976 828 977
rect 998 981 1004 982
rect 998 977 999 981
rect 1003 977 1004 981
rect 998 976 1004 977
rect 1166 981 1172 982
rect 1166 977 1167 981
rect 1171 977 1172 981
rect 1166 976 1172 977
rect 1326 981 1332 982
rect 1326 977 1327 981
rect 1331 977 1332 981
rect 1326 976 1332 977
rect 1486 981 1492 982
rect 1486 977 1487 981
rect 1491 977 1492 981
rect 1486 976 1492 977
rect 1654 981 1660 982
rect 1654 977 1655 981
rect 1659 977 1660 981
rect 1910 981 1911 985
rect 1915 981 1916 985
rect 1910 980 1916 981
rect 2118 985 2124 986
rect 2118 981 2119 985
rect 2123 981 2124 985
rect 2118 980 2124 981
rect 2318 985 2324 986
rect 2318 981 2319 985
rect 2323 981 2324 985
rect 2318 980 2324 981
rect 2510 985 2516 986
rect 2510 981 2511 985
rect 2515 981 2516 985
rect 2510 980 2516 981
rect 2686 985 2692 986
rect 2686 981 2687 985
rect 2691 981 2692 985
rect 2686 980 2692 981
rect 2854 985 2860 986
rect 2854 981 2855 985
rect 2859 981 2860 985
rect 2854 980 2860 981
rect 3014 985 3020 986
rect 3014 981 3015 985
rect 3019 981 3020 985
rect 3014 980 3020 981
rect 3174 985 3180 986
rect 3174 981 3175 985
rect 3179 981 3180 985
rect 3174 980 3180 981
rect 3334 985 3340 986
rect 3334 981 3335 985
rect 3339 981 3340 985
rect 3334 980 3340 981
rect 3478 985 3484 986
rect 3478 981 3479 985
rect 3483 981 3484 985
rect 3478 980 3484 981
rect 1654 976 1660 977
rect 110 968 116 969
rect 1822 968 1828 969
rect 110 964 111 968
rect 115 964 116 968
rect 215 967 221 968
rect 215 966 216 967
rect 197 964 216 966
rect 110 963 116 964
rect 215 963 216 964
rect 220 963 221 967
rect 1079 967 1085 968
rect 1079 966 1080 967
rect 1053 964 1080 966
rect 215 962 221 963
rect 223 963 229 964
rect 223 959 224 963
rect 228 962 229 963
rect 535 963 541 964
rect 228 960 305 962
rect 228 959 229 960
rect 223 958 229 959
rect 535 959 536 963
rect 540 962 541 963
rect 727 963 733 964
rect 540 960 665 962
rect 540 959 541 960
rect 535 958 541 959
rect 727 959 728 963
rect 732 962 733 963
rect 1079 963 1080 964
rect 1084 963 1085 967
rect 1230 967 1236 968
rect 1230 966 1231 967
rect 1221 964 1231 966
rect 1079 962 1085 963
rect 1230 963 1231 964
rect 1235 963 1236 967
rect 1399 967 1405 968
rect 1399 966 1400 967
rect 1381 964 1400 966
rect 1230 962 1236 963
rect 1399 963 1400 964
rect 1404 963 1405 967
rect 1822 964 1823 968
rect 1827 964 1828 968
rect 1399 962 1405 963
rect 1578 963 1584 964
rect 1822 963 1828 964
rect 732 960 841 962
rect 732 959 733 960
rect 727 958 733 959
rect 1578 959 1579 963
rect 1583 962 1584 963
rect 1583 960 1673 962
rect 1583 959 1584 960
rect 1578 958 1584 959
rect 1886 959 1892 960
rect 1886 955 1887 959
rect 1891 955 1892 959
rect 1886 954 1892 955
rect 2070 959 2076 960
rect 2070 955 2071 959
rect 2075 955 2076 959
rect 2070 954 2076 955
rect 2262 959 2268 960
rect 2262 955 2263 959
rect 2267 955 2268 959
rect 2262 954 2268 955
rect 2454 959 2460 960
rect 2454 955 2455 959
rect 2459 955 2460 959
rect 2454 954 2460 955
rect 2630 959 2636 960
rect 2630 955 2631 959
rect 2635 955 2636 959
rect 2630 954 2636 955
rect 2798 959 2804 960
rect 2798 955 2799 959
rect 2803 955 2804 959
rect 2798 954 2804 955
rect 2950 959 2956 960
rect 2950 955 2951 959
rect 2955 955 2956 959
rect 2950 954 2956 955
rect 3094 959 3100 960
rect 3094 955 3095 959
rect 3099 955 3100 959
rect 3094 954 3100 955
rect 3230 959 3236 960
rect 3230 955 3231 959
rect 3235 955 3236 959
rect 3230 954 3236 955
rect 3366 959 3372 960
rect 3366 955 3367 959
rect 3371 955 3372 959
rect 3366 954 3372 955
rect 3478 959 3484 960
rect 3478 955 3479 959
rect 3483 955 3484 959
rect 3478 954 3484 955
rect 110 951 116 952
rect 110 947 111 951
rect 115 947 116 951
rect 599 951 605 952
rect 599 950 600 951
rect 513 948 600 950
rect 110 946 116 947
rect 599 947 600 948
rect 604 947 605 951
rect 599 946 605 947
rect 1822 951 1828 952
rect 1822 947 1823 951
rect 1827 947 1828 951
rect 2526 951 2532 952
rect 1822 946 1828 947
rect 1862 949 1868 950
rect 1862 945 1863 949
rect 1867 945 1868 949
rect 2526 947 2527 951
rect 2531 950 2532 951
rect 3350 951 3356 952
rect 2531 948 2649 950
rect 2531 947 2532 948
rect 2526 946 2532 947
rect 3350 947 3351 951
rect 3355 950 3356 951
rect 3355 948 3385 950
rect 3574 949 3580 950
rect 3355 947 3356 948
rect 3350 946 3356 947
rect 1862 944 1868 945
rect 3574 945 3575 949
rect 3579 945 3580 949
rect 3574 944 3580 945
rect 134 941 140 942
rect 134 937 135 941
rect 139 937 140 941
rect 134 936 140 937
rect 278 941 284 942
rect 278 937 279 941
rect 283 937 284 941
rect 278 936 284 937
rect 454 941 460 942
rect 454 937 455 941
rect 459 937 460 941
rect 454 936 460 937
rect 638 941 644 942
rect 638 937 639 941
rect 643 937 644 941
rect 638 936 644 937
rect 814 941 820 942
rect 814 937 815 941
rect 819 937 820 941
rect 814 936 820 937
rect 990 941 996 942
rect 990 937 991 941
rect 995 937 996 941
rect 990 936 996 937
rect 1158 941 1164 942
rect 1158 937 1159 941
rect 1163 937 1164 941
rect 1158 936 1164 937
rect 1318 941 1324 942
rect 1318 937 1319 941
rect 1323 937 1324 941
rect 1318 936 1324 937
rect 1478 941 1484 942
rect 1478 937 1479 941
rect 1483 937 1484 941
rect 1478 936 1484 937
rect 1646 941 1652 942
rect 1646 937 1647 941
rect 1651 937 1652 941
rect 1646 936 1652 937
rect 1527 935 1533 936
rect 1527 931 1528 935
rect 1532 934 1533 935
rect 1543 935 1549 936
rect 1543 934 1544 935
rect 1532 932 1544 934
rect 1532 931 1533 932
rect 1527 930 1533 931
rect 1543 931 1544 932
rect 1548 931 1549 935
rect 2063 935 2069 936
rect 2063 934 2064 935
rect 1543 930 1549 931
rect 1862 932 1868 933
rect 1949 932 2064 934
rect 1862 928 1863 932
rect 1867 928 1868 932
rect 2063 931 2064 932
rect 2068 931 2069 935
rect 2174 935 2180 936
rect 2174 934 2175 935
rect 2133 932 2175 934
rect 2063 930 2069 931
rect 2174 931 2175 932
rect 2179 931 2180 935
rect 2447 935 2453 936
rect 2447 934 2448 935
rect 2325 932 2448 934
rect 2174 930 2180 931
rect 2447 931 2448 932
rect 2452 931 2453 935
rect 2623 935 2629 936
rect 2623 934 2624 935
rect 2517 932 2624 934
rect 2447 930 2453 931
rect 2623 931 2624 932
rect 2628 931 2629 935
rect 2943 935 2949 936
rect 2943 934 2944 935
rect 2861 932 2944 934
rect 2623 930 2629 931
rect 2943 931 2944 932
rect 2948 931 2949 935
rect 3087 935 3093 936
rect 3087 934 3088 935
rect 3013 932 3088 934
rect 2943 930 2949 931
rect 3087 931 3088 932
rect 3092 931 3093 935
rect 3223 935 3229 936
rect 3223 934 3224 935
rect 3157 932 3224 934
rect 3087 930 3093 931
rect 3223 931 3224 932
rect 3228 931 3229 935
rect 3359 935 3365 936
rect 3359 934 3360 935
rect 3293 932 3360 934
rect 3223 930 3229 931
rect 3359 931 3360 932
rect 3364 931 3365 935
rect 3359 930 3365 931
rect 3470 935 3476 936
rect 3470 931 3471 935
rect 3475 934 3476 935
rect 3475 932 3505 934
rect 3574 932 3580 933
rect 3475 931 3476 932
rect 3470 930 3476 931
rect 1862 927 1868 928
rect 3574 928 3575 932
rect 3579 928 3580 932
rect 3574 927 3580 928
rect 1894 919 1900 920
rect 1894 915 1895 919
rect 1899 915 1900 919
rect 1894 914 1900 915
rect 2078 919 2084 920
rect 2078 915 2079 919
rect 2083 915 2084 919
rect 2078 914 2084 915
rect 2270 919 2276 920
rect 2270 915 2271 919
rect 2275 915 2276 919
rect 2270 914 2276 915
rect 2462 919 2468 920
rect 2462 915 2463 919
rect 2467 915 2468 919
rect 2462 914 2468 915
rect 2638 919 2644 920
rect 2638 915 2639 919
rect 2643 915 2644 919
rect 2638 914 2644 915
rect 2806 919 2812 920
rect 2806 915 2807 919
rect 2811 915 2812 919
rect 2806 914 2812 915
rect 2958 919 2964 920
rect 2958 915 2959 919
rect 2963 915 2964 919
rect 2958 914 2964 915
rect 3102 919 3108 920
rect 3102 915 3103 919
rect 3107 915 3108 919
rect 3102 914 3108 915
rect 3238 919 3244 920
rect 3238 915 3239 919
rect 3243 915 3244 919
rect 3238 914 3244 915
rect 3374 919 3380 920
rect 3374 915 3375 919
rect 3379 915 3380 919
rect 3374 914 3380 915
rect 3486 919 3492 920
rect 3486 915 3487 919
rect 3491 915 3492 919
rect 3486 914 3492 915
rect 134 911 140 912
rect 134 907 135 911
rect 139 907 140 911
rect 134 906 140 907
rect 270 911 276 912
rect 270 907 271 911
rect 275 907 276 911
rect 270 906 276 907
rect 438 911 444 912
rect 438 907 439 911
rect 443 907 444 911
rect 438 906 444 907
rect 606 911 612 912
rect 606 907 607 911
rect 611 907 612 911
rect 606 906 612 907
rect 774 911 780 912
rect 774 907 775 911
rect 779 907 780 911
rect 774 906 780 907
rect 934 911 940 912
rect 934 907 935 911
rect 939 907 940 911
rect 934 906 940 907
rect 1094 911 1100 912
rect 1094 907 1095 911
rect 1099 907 1100 911
rect 1094 906 1100 907
rect 1246 911 1252 912
rect 1246 907 1247 911
rect 1251 907 1252 911
rect 1246 906 1252 907
rect 1398 911 1404 912
rect 1398 907 1399 911
rect 1403 907 1404 911
rect 1398 906 1404 907
rect 1550 911 1556 912
rect 1550 907 1551 911
rect 1555 907 1556 911
rect 1550 906 1556 907
rect 1887 907 1893 908
rect 127 903 133 904
rect 110 901 116 902
rect 110 897 111 901
rect 115 897 116 901
rect 127 899 128 903
rect 132 902 133 903
rect 706 903 712 904
rect 132 900 153 902
rect 132 899 133 900
rect 127 898 133 899
rect 706 899 707 903
rect 711 902 712 903
rect 1006 903 1012 904
rect 1006 902 1007 903
rect 711 900 793 902
rect 993 900 1007 902
rect 711 899 712 900
rect 706 898 712 899
rect 1006 899 1007 900
rect 1011 899 1012 903
rect 1887 903 1888 907
rect 1892 906 1893 907
rect 1902 907 1908 908
rect 1902 906 1903 907
rect 1892 904 1903 906
rect 1892 903 1893 904
rect 1887 902 1893 903
rect 1902 903 1903 904
rect 1907 903 1908 907
rect 1902 902 1908 903
rect 2063 907 2069 908
rect 2063 903 2064 907
rect 2068 906 2069 907
rect 2071 907 2077 908
rect 2071 906 2072 907
rect 2068 904 2072 906
rect 2068 903 2069 904
rect 2063 902 2069 903
rect 2071 903 2072 904
rect 2076 903 2077 907
rect 2071 902 2077 903
rect 2263 907 2269 908
rect 2263 903 2264 907
rect 2268 906 2269 907
rect 2287 907 2293 908
rect 2287 906 2288 907
rect 2268 904 2288 906
rect 2268 903 2269 904
rect 2263 902 2269 903
rect 2287 903 2288 904
rect 2292 903 2293 907
rect 2287 902 2293 903
rect 2447 907 2453 908
rect 2447 903 2448 907
rect 2452 906 2453 907
rect 2455 907 2461 908
rect 2455 906 2456 907
rect 2452 904 2456 906
rect 2452 903 2453 904
rect 2447 902 2453 903
rect 2455 903 2456 904
rect 2460 903 2461 907
rect 2455 902 2461 903
rect 2623 907 2629 908
rect 2623 903 2624 907
rect 2628 906 2629 907
rect 2631 907 2637 908
rect 2631 906 2632 907
rect 2628 904 2632 906
rect 2628 903 2629 904
rect 2623 902 2629 903
rect 2631 903 2632 904
rect 2636 903 2637 907
rect 2631 902 2637 903
rect 2799 907 2805 908
rect 2799 903 2800 907
rect 2804 906 2805 907
rect 2814 907 2820 908
rect 2814 906 2815 907
rect 2804 904 2815 906
rect 2804 903 2805 904
rect 2799 902 2805 903
rect 2814 903 2815 904
rect 2819 903 2820 907
rect 2814 902 2820 903
rect 2943 907 2949 908
rect 2943 903 2944 907
rect 2948 906 2949 907
rect 2951 907 2957 908
rect 2951 906 2952 907
rect 2948 904 2952 906
rect 2948 903 2949 904
rect 2943 902 2949 903
rect 2951 903 2952 904
rect 2956 903 2957 907
rect 2951 902 2957 903
rect 3087 907 3093 908
rect 3087 903 3088 907
rect 3092 906 3093 907
rect 3095 907 3101 908
rect 3095 906 3096 907
rect 3092 904 3096 906
rect 3092 903 3093 904
rect 3087 902 3093 903
rect 3095 903 3096 904
rect 3100 903 3101 907
rect 3095 902 3101 903
rect 3223 907 3229 908
rect 3223 903 3224 907
rect 3228 906 3229 907
rect 3231 907 3237 908
rect 3231 906 3232 907
rect 3228 904 3232 906
rect 3228 903 3229 904
rect 3223 902 3229 903
rect 3231 903 3232 904
rect 3236 903 3237 907
rect 3231 902 3237 903
rect 3359 907 3365 908
rect 3359 903 3360 907
rect 3364 906 3365 907
rect 3367 907 3373 908
rect 3367 906 3368 907
rect 3364 904 3368 906
rect 3364 903 3365 904
rect 3359 902 3365 903
rect 3367 903 3368 904
rect 3372 903 3373 907
rect 3367 902 3373 903
rect 3471 907 3477 908
rect 3471 903 3472 907
rect 3476 906 3477 907
rect 3479 907 3485 908
rect 3479 906 3480 907
rect 3476 904 3480 906
rect 3476 903 3477 904
rect 3471 902 3477 903
rect 3479 903 3480 904
rect 3484 903 3485 907
rect 3479 902 3485 903
rect 1006 898 1012 899
rect 1822 901 1828 902
rect 110 896 116 897
rect 1822 897 1823 901
rect 1827 897 1828 901
rect 1822 896 1828 897
rect 202 887 208 888
rect 110 884 116 885
rect 110 880 111 884
rect 115 880 116 884
rect 202 883 203 887
rect 207 886 208 887
rect 338 887 344 888
rect 207 884 297 886
rect 207 883 208 884
rect 202 882 208 883
rect 338 883 339 887
rect 343 886 344 887
rect 767 887 773 888
rect 767 886 768 887
rect 343 884 465 886
rect 669 884 768 886
rect 343 883 344 884
rect 338 882 344 883
rect 767 883 768 884
rect 772 883 773 887
rect 767 882 773 883
rect 1002 887 1008 888
rect 1002 883 1003 887
rect 1007 886 1008 887
rect 1391 887 1397 888
rect 1391 886 1392 887
rect 1007 884 1121 886
rect 1309 884 1392 886
rect 1007 883 1008 884
rect 1002 882 1008 883
rect 1391 883 1392 884
rect 1396 883 1397 887
rect 1479 887 1485 888
rect 1479 886 1480 887
rect 1461 884 1480 886
rect 1391 882 1397 883
rect 1479 883 1480 884
rect 1484 883 1485 887
rect 1479 882 1485 883
rect 1494 887 1500 888
rect 1494 883 1495 887
rect 1499 886 1500 887
rect 1887 887 1893 888
rect 1499 884 1577 886
rect 1822 884 1828 885
rect 1499 883 1500 884
rect 1494 882 1500 883
rect 110 879 116 880
rect 1822 880 1823 884
rect 1827 880 1828 884
rect 1887 883 1888 887
rect 1892 886 1893 887
rect 1962 887 1968 888
rect 1962 886 1963 887
rect 1892 884 1963 886
rect 1892 883 1893 884
rect 1887 882 1893 883
rect 1962 883 1963 884
rect 1967 883 1968 887
rect 1962 882 1968 883
rect 2015 887 2021 888
rect 2015 883 2016 887
rect 2020 886 2021 887
rect 2103 887 2109 888
rect 2103 886 2104 887
rect 2020 884 2104 886
rect 2020 883 2021 884
rect 2015 882 2021 883
rect 2103 883 2104 884
rect 2108 883 2109 887
rect 2103 882 2109 883
rect 2174 887 2181 888
rect 2174 883 2175 887
rect 2180 883 2181 887
rect 2174 882 2181 883
rect 2343 887 2349 888
rect 2343 883 2344 887
rect 2348 886 2349 887
rect 2438 887 2444 888
rect 2438 886 2439 887
rect 2348 884 2439 886
rect 2348 883 2349 884
rect 2343 882 2349 883
rect 2438 883 2439 884
rect 2443 883 2444 887
rect 2438 882 2444 883
rect 2511 887 2517 888
rect 2511 883 2512 887
rect 2516 886 2517 887
rect 2606 887 2612 888
rect 2606 886 2607 887
rect 2516 884 2607 886
rect 2516 883 2517 884
rect 2511 882 2517 883
rect 2606 883 2607 884
rect 2611 883 2612 887
rect 2606 882 2612 883
rect 2679 887 2685 888
rect 2679 883 2680 887
rect 2684 886 2685 887
rect 2694 887 2700 888
rect 2694 886 2695 887
rect 2684 884 2695 886
rect 2684 883 2685 884
rect 2679 882 2685 883
rect 2694 883 2695 884
rect 2699 883 2700 887
rect 2694 882 2700 883
rect 2831 887 2837 888
rect 2831 883 2832 887
rect 2836 886 2837 887
rect 2906 887 2912 888
rect 2906 886 2907 887
rect 2836 884 2907 886
rect 2836 883 2837 884
rect 2831 882 2837 883
rect 2906 883 2907 884
rect 2911 883 2912 887
rect 2906 882 2912 883
rect 2975 887 2981 888
rect 2975 883 2976 887
rect 2980 886 2981 887
rect 3050 887 3056 888
rect 3050 886 3051 887
rect 2980 884 3051 886
rect 2980 883 2981 884
rect 2975 882 2981 883
rect 3050 883 3051 884
rect 3055 883 3056 887
rect 3050 882 3056 883
rect 3111 887 3117 888
rect 3111 883 3112 887
rect 3116 886 3117 887
rect 3198 887 3204 888
rect 3198 886 3199 887
rect 3116 884 3199 886
rect 3116 883 3117 884
rect 3111 882 3117 883
rect 3198 883 3199 884
rect 3203 883 3204 887
rect 3198 882 3204 883
rect 3239 887 3245 888
rect 3239 883 3240 887
rect 3244 886 3245 887
rect 3314 887 3320 888
rect 3314 886 3315 887
rect 3244 884 3315 886
rect 3244 883 3245 884
rect 3239 882 3245 883
rect 3314 883 3315 884
rect 3319 883 3320 887
rect 3314 882 3320 883
rect 3351 887 3357 888
rect 3351 883 3352 887
rect 3356 886 3357 887
rect 3367 887 3373 888
rect 3367 886 3368 887
rect 3356 884 3368 886
rect 3356 883 3357 884
rect 3351 882 3357 883
rect 3367 883 3368 884
rect 3372 883 3373 887
rect 3367 882 3373 883
rect 3470 887 3476 888
rect 3470 883 3471 887
rect 3475 886 3476 887
rect 3479 887 3485 888
rect 3479 886 3480 887
rect 3475 884 3480 886
rect 3475 883 3476 884
rect 3470 882 3476 883
rect 3479 883 3480 884
rect 3484 883 3485 887
rect 3479 882 3485 883
rect 1822 879 1828 880
rect 1894 877 1900 878
rect 1894 873 1895 877
rect 1899 873 1900 877
rect 1894 872 1900 873
rect 2022 877 2028 878
rect 2022 873 2023 877
rect 2027 873 2028 877
rect 2022 872 2028 873
rect 2182 877 2188 878
rect 2182 873 2183 877
rect 2187 873 2188 877
rect 2182 872 2188 873
rect 2350 877 2356 878
rect 2350 873 2351 877
rect 2355 873 2356 877
rect 2350 872 2356 873
rect 2518 877 2524 878
rect 2518 873 2519 877
rect 2523 873 2524 877
rect 2518 872 2524 873
rect 2686 877 2692 878
rect 2686 873 2687 877
rect 2691 873 2692 877
rect 2686 872 2692 873
rect 2838 877 2844 878
rect 2838 873 2839 877
rect 2843 873 2844 877
rect 2838 872 2844 873
rect 2982 877 2988 878
rect 2982 873 2983 877
rect 2987 873 2988 877
rect 2982 872 2988 873
rect 3118 877 3124 878
rect 3118 873 3119 877
rect 3123 873 3124 877
rect 3118 872 3124 873
rect 3246 877 3252 878
rect 3246 873 3247 877
rect 3251 873 3252 877
rect 3246 872 3252 873
rect 3374 877 3380 878
rect 3374 873 3375 877
rect 3379 873 3380 877
rect 3374 872 3380 873
rect 3486 877 3492 878
rect 3486 873 3487 877
rect 3491 873 3492 877
rect 3486 872 3492 873
rect 142 871 148 872
rect 142 867 143 871
rect 147 867 148 871
rect 142 866 148 867
rect 278 871 284 872
rect 278 867 279 871
rect 283 867 284 871
rect 278 866 284 867
rect 446 871 452 872
rect 446 867 447 871
rect 451 867 452 871
rect 446 866 452 867
rect 614 871 620 872
rect 614 867 615 871
rect 619 867 620 871
rect 614 866 620 867
rect 782 871 788 872
rect 782 867 783 871
rect 787 867 788 871
rect 782 866 788 867
rect 942 871 948 872
rect 942 867 943 871
rect 947 867 948 871
rect 942 866 948 867
rect 1102 871 1108 872
rect 1102 867 1103 871
rect 1107 867 1108 871
rect 1102 866 1108 867
rect 1254 871 1260 872
rect 1254 867 1255 871
rect 1259 867 1260 871
rect 1254 866 1260 867
rect 1406 871 1412 872
rect 1406 867 1407 871
rect 1411 867 1412 871
rect 1406 866 1412 867
rect 1558 871 1564 872
rect 1558 867 1559 871
rect 1563 867 1564 871
rect 1558 866 1564 867
rect 1862 864 1868 865
rect 1862 860 1863 864
rect 1867 860 1868 864
rect 3574 864 3580 865
rect 3574 860 3575 864
rect 3579 860 3580 864
rect 135 859 141 860
rect 135 855 136 859
rect 140 858 141 859
rect 198 859 204 860
rect 198 858 199 859
rect 140 856 199 858
rect 140 855 141 856
rect 135 854 141 855
rect 198 855 199 856
rect 203 855 204 859
rect 198 854 204 855
rect 207 859 213 860
rect 207 855 208 859
rect 212 858 213 859
rect 271 859 277 860
rect 271 858 272 859
rect 212 856 272 858
rect 212 855 213 856
rect 207 854 213 855
rect 271 855 272 856
rect 276 855 277 859
rect 271 854 277 855
rect 439 859 445 860
rect 439 855 440 859
rect 444 858 445 859
rect 454 859 460 860
rect 454 858 455 859
rect 444 856 455 858
rect 444 855 445 856
rect 439 854 445 855
rect 454 855 455 856
rect 459 855 460 859
rect 454 854 460 855
rect 599 859 605 860
rect 599 855 600 859
rect 604 858 605 859
rect 607 859 613 860
rect 607 858 608 859
rect 604 856 608 858
rect 604 855 605 856
rect 599 854 605 855
rect 607 855 608 856
rect 612 855 613 859
rect 607 854 613 855
rect 767 859 773 860
rect 767 855 768 859
rect 772 858 773 859
rect 775 859 781 860
rect 775 858 776 859
rect 772 856 776 858
rect 772 855 773 856
rect 767 854 773 855
rect 775 855 776 856
rect 780 855 781 859
rect 775 854 781 855
rect 935 859 941 860
rect 935 855 936 859
rect 940 858 941 859
rect 1002 859 1008 860
rect 1002 858 1003 859
rect 940 856 1003 858
rect 940 855 941 856
rect 935 854 941 855
rect 1002 855 1003 856
rect 1007 855 1008 859
rect 1002 854 1008 855
rect 1047 859 1053 860
rect 1047 855 1048 859
rect 1052 858 1053 859
rect 1095 859 1101 860
rect 1095 858 1096 859
rect 1052 856 1096 858
rect 1052 855 1053 856
rect 1047 854 1053 855
rect 1095 855 1096 856
rect 1100 855 1101 859
rect 1095 854 1101 855
rect 1247 859 1253 860
rect 1247 855 1248 859
rect 1252 858 1253 859
rect 1262 859 1268 860
rect 1262 858 1263 859
rect 1252 856 1263 858
rect 1252 855 1253 856
rect 1247 854 1253 855
rect 1262 855 1263 856
rect 1267 855 1268 859
rect 1262 854 1268 855
rect 1391 859 1397 860
rect 1391 855 1392 859
rect 1396 858 1397 859
rect 1399 859 1405 860
rect 1399 858 1400 859
rect 1396 856 1400 858
rect 1396 855 1397 856
rect 1391 854 1397 855
rect 1399 855 1400 856
rect 1404 855 1405 859
rect 1399 854 1405 855
rect 1543 859 1549 860
rect 1543 855 1544 859
rect 1548 858 1549 859
rect 1551 859 1557 860
rect 1862 859 1868 860
rect 1962 859 1968 860
rect 1551 858 1552 859
rect 1548 856 1552 858
rect 1548 855 1549 856
rect 1543 854 1549 855
rect 1551 855 1552 856
rect 1556 855 1557 859
rect 1551 854 1557 855
rect 1962 855 1963 859
rect 1967 858 1968 859
rect 2103 859 2109 860
rect 1967 856 2041 858
rect 1967 855 1968 856
rect 1962 854 1968 855
rect 2103 855 2104 859
rect 2108 858 2109 859
rect 2287 859 2293 860
rect 2108 856 2201 858
rect 2108 855 2109 856
rect 2103 854 2109 855
rect 2287 855 2288 859
rect 2292 858 2293 859
rect 2438 859 2444 860
rect 2292 856 2369 858
rect 2292 855 2293 856
rect 2287 854 2293 855
rect 2438 855 2439 859
rect 2443 858 2444 859
rect 2606 859 2612 860
rect 2443 856 2537 858
rect 2443 855 2444 856
rect 2438 854 2444 855
rect 2606 855 2607 859
rect 2611 858 2612 859
rect 2906 859 2912 860
rect 2611 856 2705 858
rect 2611 855 2612 856
rect 2606 854 2612 855
rect 2906 855 2907 859
rect 2911 858 2912 859
rect 3050 859 3056 860
rect 2911 856 3001 858
rect 2911 855 2912 856
rect 2906 854 2912 855
rect 3050 855 3051 859
rect 3055 858 3056 859
rect 3198 859 3204 860
rect 3055 856 3137 858
rect 3055 855 3056 856
rect 3050 854 3056 855
rect 3198 855 3199 859
rect 3203 858 3204 859
rect 3314 859 3320 860
rect 3574 859 3580 860
rect 3203 856 3265 858
rect 3203 855 3204 856
rect 3198 854 3204 855
rect 3314 855 3315 859
rect 3319 858 3320 859
rect 3319 856 3393 858
rect 3319 855 3320 856
rect 3314 854 3320 855
rect 127 847 133 848
rect 127 843 128 847
rect 132 846 133 847
rect 135 847 141 848
rect 135 846 136 847
rect 132 844 136 846
rect 132 843 133 844
rect 127 842 133 843
rect 135 843 136 844
rect 140 843 141 847
rect 135 842 141 843
rect 279 847 285 848
rect 279 843 280 847
rect 284 846 285 847
rect 338 847 344 848
rect 338 846 339 847
rect 284 844 339 846
rect 284 843 285 844
rect 279 842 285 843
rect 338 843 339 844
rect 343 843 344 847
rect 338 842 344 843
rect 375 847 381 848
rect 375 843 376 847
rect 380 846 381 847
rect 455 847 461 848
rect 455 846 456 847
rect 380 844 456 846
rect 380 843 381 844
rect 375 842 381 843
rect 455 843 456 844
rect 460 843 461 847
rect 455 842 461 843
rect 543 847 549 848
rect 543 843 544 847
rect 548 846 549 847
rect 631 847 637 848
rect 631 846 632 847
rect 548 844 632 846
rect 548 843 549 844
rect 543 842 549 843
rect 631 843 632 844
rect 636 843 637 847
rect 631 842 637 843
rect 719 847 725 848
rect 719 843 720 847
rect 724 846 725 847
rect 799 847 805 848
rect 799 846 800 847
rect 724 844 800 846
rect 724 843 725 844
rect 719 842 725 843
rect 799 843 800 844
rect 804 843 805 847
rect 799 842 805 843
rect 975 847 981 848
rect 975 843 976 847
rect 980 846 981 847
rect 1058 847 1064 848
rect 1058 846 1059 847
rect 980 844 1059 846
rect 980 843 981 844
rect 975 842 981 843
rect 1058 843 1059 844
rect 1063 843 1064 847
rect 1058 842 1064 843
rect 1151 847 1157 848
rect 1151 843 1152 847
rect 1156 846 1157 847
rect 1166 847 1172 848
rect 1166 846 1167 847
rect 1156 844 1167 846
rect 1156 843 1157 844
rect 1151 842 1157 843
rect 1166 843 1167 844
rect 1171 843 1172 847
rect 1166 842 1172 843
rect 1327 847 1333 848
rect 1327 843 1328 847
rect 1332 846 1333 847
rect 1407 847 1413 848
rect 1407 846 1408 847
rect 1332 844 1408 846
rect 1332 843 1333 844
rect 1327 842 1333 843
rect 1407 843 1408 844
rect 1412 843 1413 847
rect 1407 842 1413 843
rect 1479 847 1485 848
rect 1479 843 1480 847
rect 1484 846 1485 847
rect 1503 847 1509 848
rect 1503 846 1504 847
rect 1484 844 1504 846
rect 1484 843 1485 844
rect 1479 842 1485 843
rect 1503 843 1504 844
rect 1508 843 1509 847
rect 1503 842 1509 843
rect 1862 847 1868 848
rect 1862 843 1863 847
rect 1867 843 1868 847
rect 1862 842 1868 843
rect 1879 847 1885 848
rect 1879 843 1880 847
rect 1884 846 1885 847
rect 2806 847 2812 848
rect 1884 844 1905 846
rect 1884 843 1885 844
rect 1879 842 1885 843
rect 2806 843 2807 847
rect 2811 846 2812 847
rect 3471 847 3477 848
rect 2811 844 2849 846
rect 2811 843 2812 844
rect 2806 842 2812 843
rect 3471 843 3472 847
rect 3476 846 3477 847
rect 3574 847 3580 848
rect 3476 844 3497 846
rect 3476 843 3477 844
rect 3471 842 3477 843
rect 3574 843 3575 847
rect 3579 843 3580 847
rect 3574 842 3580 843
rect 142 837 148 838
rect 142 833 143 837
rect 147 833 148 837
rect 142 832 148 833
rect 286 837 292 838
rect 286 833 287 837
rect 291 833 292 837
rect 286 832 292 833
rect 462 837 468 838
rect 462 833 463 837
rect 467 833 468 837
rect 462 832 468 833
rect 638 837 644 838
rect 638 833 639 837
rect 643 833 644 837
rect 638 832 644 833
rect 806 837 812 838
rect 806 833 807 837
rect 811 833 812 837
rect 806 832 812 833
rect 982 837 988 838
rect 982 833 983 837
rect 987 833 988 837
rect 982 832 988 833
rect 1158 837 1164 838
rect 1158 833 1159 837
rect 1163 833 1164 837
rect 1158 832 1164 833
rect 1334 837 1340 838
rect 1334 833 1335 837
rect 1339 833 1340 837
rect 1334 832 1340 833
rect 1510 837 1516 838
rect 1510 833 1511 837
rect 1515 833 1516 837
rect 1510 832 1516 833
rect 1886 837 1892 838
rect 1886 833 1887 837
rect 1891 833 1892 837
rect 1886 832 1892 833
rect 2014 837 2020 838
rect 2014 833 2015 837
rect 2019 833 2020 837
rect 2014 832 2020 833
rect 2174 837 2180 838
rect 2174 833 2175 837
rect 2179 833 2180 837
rect 2174 832 2180 833
rect 2342 837 2348 838
rect 2342 833 2343 837
rect 2347 833 2348 837
rect 2342 832 2348 833
rect 2510 837 2516 838
rect 2510 833 2511 837
rect 2515 833 2516 837
rect 2510 832 2516 833
rect 2678 837 2684 838
rect 2678 833 2679 837
rect 2683 833 2684 837
rect 2678 832 2684 833
rect 2830 837 2836 838
rect 2830 833 2831 837
rect 2835 833 2836 837
rect 2830 832 2836 833
rect 2974 837 2980 838
rect 2974 833 2975 837
rect 2979 833 2980 837
rect 2974 832 2980 833
rect 3110 837 3116 838
rect 3110 833 3111 837
rect 3115 833 3116 837
rect 3110 832 3116 833
rect 3238 837 3244 838
rect 3238 833 3239 837
rect 3243 833 3244 837
rect 3238 832 3244 833
rect 3366 837 3372 838
rect 3366 833 3367 837
rect 3371 833 3372 837
rect 3366 832 3372 833
rect 3478 837 3484 838
rect 3478 833 3479 837
rect 3483 833 3484 837
rect 3478 832 3484 833
rect 110 824 116 825
rect 1822 824 1828 825
rect 110 820 111 824
rect 115 820 116 824
rect 207 823 213 824
rect 207 822 208 823
rect 197 820 208 822
rect 110 819 116 820
rect 207 819 208 820
rect 212 819 213 823
rect 375 823 381 824
rect 375 822 376 823
rect 341 820 376 822
rect 207 818 213 819
rect 375 819 376 820
rect 380 819 381 823
rect 543 823 549 824
rect 543 822 544 823
rect 517 820 544 822
rect 375 818 381 819
rect 543 819 544 820
rect 548 819 549 823
rect 719 823 725 824
rect 719 822 720 823
rect 693 820 720 822
rect 543 818 549 819
rect 719 819 720 820
rect 724 819 725 823
rect 1047 823 1053 824
rect 1047 822 1048 823
rect 1037 820 1048 822
rect 719 818 725 819
rect 1047 819 1048 820
rect 1052 819 1053 823
rect 1822 820 1823 824
rect 1827 820 1828 824
rect 1047 818 1053 819
rect 1058 819 1064 820
rect 1058 815 1059 819
rect 1063 818 1064 819
rect 1407 819 1413 820
rect 1822 819 1828 820
rect 1063 816 1177 818
rect 1063 815 1064 816
rect 1058 814 1064 815
rect 1407 815 1408 819
rect 1412 818 1413 819
rect 1412 816 1529 818
rect 1412 815 1413 816
rect 1407 814 1413 815
rect 110 807 116 808
rect 110 803 111 807
rect 115 803 116 807
rect 110 802 116 803
rect 790 807 796 808
rect 790 803 791 807
rect 795 806 796 807
rect 1294 807 1300 808
rect 795 804 817 806
rect 795 803 796 804
rect 790 802 796 803
rect 1294 803 1295 807
rect 1299 806 1300 807
rect 1822 807 1828 808
rect 1299 804 1345 806
rect 1299 803 1300 804
rect 1294 802 1300 803
rect 1822 803 1823 807
rect 1827 803 1828 807
rect 1822 802 1828 803
rect 1886 807 1892 808
rect 1886 803 1887 807
rect 1891 803 1892 807
rect 1886 802 1892 803
rect 2070 807 2076 808
rect 2070 803 2071 807
rect 2075 803 2076 807
rect 2070 802 2076 803
rect 2262 807 2268 808
rect 2262 803 2263 807
rect 2267 803 2268 807
rect 2262 802 2268 803
rect 2446 807 2452 808
rect 2446 803 2447 807
rect 2451 803 2452 807
rect 2446 802 2452 803
rect 2622 807 2628 808
rect 2622 803 2623 807
rect 2627 803 2628 807
rect 2622 802 2628 803
rect 2790 807 2796 808
rect 2790 803 2791 807
rect 2795 803 2796 807
rect 2790 802 2796 803
rect 2942 807 2948 808
rect 2942 803 2943 807
rect 2947 803 2948 807
rect 2942 802 2948 803
rect 3086 807 3092 808
rect 3086 803 3087 807
rect 3091 803 3092 807
rect 3086 802 3092 803
rect 3222 807 3228 808
rect 3222 803 3223 807
rect 3227 803 3228 807
rect 3222 802 3228 803
rect 3358 807 3364 808
rect 3358 803 3359 807
rect 3363 803 3364 807
rect 3358 802 3364 803
rect 3478 807 3484 808
rect 3478 803 3479 807
rect 3483 803 3484 807
rect 3478 802 3484 803
rect 1954 799 1960 800
rect 134 797 140 798
rect 134 793 135 797
rect 139 793 140 797
rect 134 792 140 793
rect 278 797 284 798
rect 278 793 279 797
rect 283 793 284 797
rect 278 792 284 793
rect 454 797 460 798
rect 454 793 455 797
rect 459 793 460 797
rect 454 792 460 793
rect 630 797 636 798
rect 630 793 631 797
rect 635 793 636 797
rect 630 792 636 793
rect 798 797 804 798
rect 798 793 799 797
rect 803 793 804 797
rect 798 792 804 793
rect 974 797 980 798
rect 974 793 975 797
rect 979 793 980 797
rect 974 792 980 793
rect 1150 797 1156 798
rect 1150 793 1151 797
rect 1155 793 1156 797
rect 1150 792 1156 793
rect 1326 797 1332 798
rect 1326 793 1327 797
rect 1331 793 1332 797
rect 1326 792 1332 793
rect 1502 797 1508 798
rect 1502 793 1503 797
rect 1507 793 1508 797
rect 1502 792 1508 793
rect 1862 797 1868 798
rect 1862 793 1863 797
rect 1867 793 1868 797
rect 1954 795 1955 799
rect 1959 798 1960 799
rect 2694 799 2700 800
rect 2694 798 2695 799
rect 1959 796 2089 798
rect 2681 796 2695 798
rect 1959 795 1960 796
rect 1954 794 1960 795
rect 2694 795 2695 796
rect 2699 795 2700 799
rect 2694 794 2700 795
rect 3351 799 3357 800
rect 3351 795 3352 799
rect 3356 798 3357 799
rect 3356 796 3377 798
rect 3574 797 3580 798
rect 3356 795 3357 796
rect 3351 794 3357 795
rect 1862 792 1868 793
rect 3574 793 3575 797
rect 3579 793 3580 797
rect 3574 792 3580 793
rect 2063 783 2069 784
rect 2063 782 2064 783
rect 1862 780 1868 781
rect 1949 780 2064 782
rect 1862 776 1863 780
rect 1867 776 1868 780
rect 2063 779 2064 780
rect 2068 779 2069 783
rect 2439 783 2445 784
rect 2439 782 2440 783
rect 2325 780 2440 782
rect 2063 778 2069 779
rect 2439 779 2440 780
rect 2444 779 2445 783
rect 2615 783 2621 784
rect 2615 782 2616 783
rect 2509 780 2616 782
rect 2439 778 2445 779
rect 2615 779 2616 780
rect 2620 779 2621 783
rect 2935 783 2941 784
rect 2935 782 2936 783
rect 2853 780 2936 782
rect 2615 778 2621 779
rect 2935 779 2936 780
rect 2940 779 2941 783
rect 3079 783 3085 784
rect 3079 782 3080 783
rect 3005 780 3080 782
rect 2935 778 2941 779
rect 3079 779 3080 780
rect 3084 779 3085 783
rect 3158 783 3164 784
rect 3158 782 3159 783
rect 3149 780 3159 782
rect 3079 778 3085 779
rect 3158 779 3159 780
rect 3163 779 3164 783
rect 3351 783 3357 784
rect 3351 782 3352 783
rect 3285 780 3352 782
rect 3158 778 3164 779
rect 3351 779 3352 780
rect 3356 779 3357 783
rect 3351 778 3357 779
rect 3426 783 3432 784
rect 3426 779 3427 783
rect 3431 782 3432 783
rect 3431 780 3505 782
rect 3574 780 3580 781
rect 3431 779 3432 780
rect 3426 778 3432 779
rect 1862 775 1868 776
rect 3574 776 3575 780
rect 3579 776 3580 780
rect 3574 775 3580 776
rect 134 771 140 772
rect 134 767 135 771
rect 139 767 140 771
rect 134 766 140 767
rect 270 771 276 772
rect 270 767 271 771
rect 275 767 276 771
rect 270 766 276 767
rect 438 771 444 772
rect 438 767 439 771
rect 443 767 444 771
rect 438 766 444 767
rect 606 771 612 772
rect 606 767 607 771
rect 611 767 612 771
rect 606 766 612 767
rect 774 771 780 772
rect 774 767 775 771
rect 779 767 780 771
rect 774 766 780 767
rect 934 771 940 772
rect 934 767 935 771
rect 939 767 940 771
rect 934 766 940 767
rect 1086 771 1092 772
rect 1086 767 1087 771
rect 1091 767 1092 771
rect 1086 766 1092 767
rect 1238 771 1244 772
rect 1238 767 1239 771
rect 1243 767 1244 771
rect 1238 766 1244 767
rect 1390 771 1396 772
rect 1390 767 1391 771
rect 1395 767 1396 771
rect 1390 766 1396 767
rect 1550 771 1556 772
rect 1550 767 1551 771
rect 1555 767 1556 771
rect 1550 766 1556 767
rect 1894 767 1900 768
rect 127 763 133 764
rect 110 761 116 762
rect 110 757 111 761
rect 115 757 116 761
rect 127 759 128 763
rect 132 762 133 763
rect 1166 763 1172 764
rect 1166 762 1167 763
rect 132 760 153 762
rect 1145 760 1167 762
rect 132 759 133 760
rect 127 758 133 759
rect 1166 759 1167 760
rect 1171 759 1172 763
rect 1894 763 1895 767
rect 1899 763 1900 767
rect 1894 762 1900 763
rect 2078 767 2084 768
rect 2078 763 2079 767
rect 2083 763 2084 767
rect 2078 762 2084 763
rect 2270 767 2276 768
rect 2270 763 2271 767
rect 2275 763 2276 767
rect 2270 762 2276 763
rect 2454 767 2460 768
rect 2454 763 2455 767
rect 2459 763 2460 767
rect 2454 762 2460 763
rect 2630 767 2636 768
rect 2630 763 2631 767
rect 2635 763 2636 767
rect 2630 762 2636 763
rect 2798 767 2804 768
rect 2798 763 2799 767
rect 2803 763 2804 767
rect 2798 762 2804 763
rect 2950 767 2956 768
rect 2950 763 2951 767
rect 2955 763 2956 767
rect 2950 762 2956 763
rect 3094 767 3100 768
rect 3094 763 3095 767
rect 3099 763 3100 767
rect 3094 762 3100 763
rect 3230 767 3236 768
rect 3230 763 3231 767
rect 3235 763 3236 767
rect 3230 762 3236 763
rect 3366 767 3372 768
rect 3366 763 3367 767
rect 3371 763 3372 767
rect 3366 762 3372 763
rect 3486 767 3492 768
rect 3486 763 3487 767
rect 3491 763 3492 767
rect 3486 762 3492 763
rect 1166 758 1172 759
rect 1822 761 1828 762
rect 110 756 116 757
rect 1822 757 1823 761
rect 1827 757 1828 761
rect 1822 756 1828 757
rect 1879 755 1885 756
rect 1879 751 1880 755
rect 1884 754 1885 755
rect 1887 755 1893 756
rect 1887 754 1888 755
rect 1884 752 1888 754
rect 1884 751 1885 752
rect 1879 750 1885 751
rect 1887 751 1888 752
rect 1892 751 1893 755
rect 1887 750 1893 751
rect 2063 755 2069 756
rect 2063 751 2064 755
rect 2068 754 2069 755
rect 2071 755 2077 756
rect 2071 754 2072 755
rect 2068 752 2072 754
rect 2068 751 2069 752
rect 2063 750 2069 751
rect 2071 751 2072 752
rect 2076 751 2077 755
rect 2071 750 2077 751
rect 2254 755 2260 756
rect 2254 751 2255 755
rect 2259 754 2260 755
rect 2263 755 2269 756
rect 2263 754 2264 755
rect 2259 752 2264 754
rect 2259 751 2260 752
rect 2254 750 2260 751
rect 2263 751 2264 752
rect 2268 751 2269 755
rect 2263 750 2269 751
rect 2439 755 2445 756
rect 2439 751 2440 755
rect 2444 754 2445 755
rect 2447 755 2453 756
rect 2447 754 2448 755
rect 2444 752 2448 754
rect 2444 751 2445 752
rect 2439 750 2445 751
rect 2447 751 2448 752
rect 2452 751 2453 755
rect 2447 750 2453 751
rect 2615 755 2621 756
rect 2615 751 2616 755
rect 2620 754 2621 755
rect 2623 755 2629 756
rect 2623 754 2624 755
rect 2620 752 2624 754
rect 2620 751 2621 752
rect 2615 750 2621 751
rect 2623 751 2624 752
rect 2628 751 2629 755
rect 2623 750 2629 751
rect 2791 755 2797 756
rect 2791 751 2792 755
rect 2796 754 2797 755
rect 2806 755 2812 756
rect 2806 754 2807 755
rect 2796 752 2807 754
rect 2796 751 2797 752
rect 2791 750 2797 751
rect 2806 751 2807 752
rect 2811 751 2812 755
rect 2806 750 2812 751
rect 2935 755 2941 756
rect 2935 751 2936 755
rect 2940 754 2941 755
rect 2943 755 2949 756
rect 2943 754 2944 755
rect 2940 752 2944 754
rect 2940 751 2941 752
rect 2935 750 2941 751
rect 2943 751 2944 752
rect 2948 751 2949 755
rect 2943 750 2949 751
rect 3079 755 3085 756
rect 3079 751 3080 755
rect 3084 754 3085 755
rect 3087 755 3093 756
rect 3087 754 3088 755
rect 3084 752 3088 754
rect 3084 751 3085 752
rect 3079 750 3085 751
rect 3087 751 3088 752
rect 3092 751 3093 755
rect 3087 750 3093 751
rect 3223 755 3229 756
rect 3223 751 3224 755
rect 3228 754 3229 755
rect 3351 755 3357 756
rect 3228 752 3346 754
rect 3228 751 3229 752
rect 3223 750 3229 751
rect 202 747 208 748
rect 110 744 116 745
rect 110 740 111 744
rect 115 740 116 744
rect 202 743 203 747
rect 207 746 208 747
rect 431 747 437 748
rect 207 744 297 746
rect 207 743 208 744
rect 202 742 208 743
rect 431 743 432 747
rect 436 746 437 747
rect 506 747 512 748
rect 436 744 465 746
rect 436 743 437 744
rect 431 742 437 743
rect 506 743 507 747
rect 511 746 512 747
rect 674 747 680 748
rect 511 744 633 746
rect 511 743 512 744
rect 506 742 512 743
rect 674 743 675 747
rect 679 746 680 747
rect 1079 747 1085 748
rect 1079 746 1080 747
rect 679 744 801 746
rect 997 744 1080 746
rect 679 743 680 744
rect 674 742 680 743
rect 1079 743 1080 744
rect 1084 743 1085 747
rect 1383 747 1389 748
rect 1383 746 1384 747
rect 1301 744 1384 746
rect 1079 742 1085 743
rect 1383 743 1384 744
rect 1388 743 1389 747
rect 1543 747 1549 748
rect 1543 746 1544 747
rect 1453 744 1544 746
rect 1383 742 1389 743
rect 1543 743 1544 744
rect 1548 743 1549 747
rect 1618 747 1624 748
rect 1618 746 1619 747
rect 1613 744 1619 746
rect 1543 742 1549 743
rect 1618 743 1619 744
rect 1623 743 1624 747
rect 3344 746 3346 752
rect 3351 751 3352 755
rect 3356 754 3357 755
rect 3359 755 3365 756
rect 3359 754 3360 755
rect 3356 752 3360 754
rect 3356 751 3357 752
rect 3351 750 3357 751
rect 3359 751 3360 752
rect 3364 751 3365 755
rect 3359 750 3365 751
rect 3463 755 3469 756
rect 3463 751 3464 755
rect 3468 754 3469 755
rect 3479 755 3485 756
rect 3479 754 3480 755
rect 3468 752 3480 754
rect 3468 751 3469 752
rect 3463 750 3469 751
rect 3479 751 3480 752
rect 3484 751 3485 755
rect 3479 750 3485 751
rect 3426 747 3432 748
rect 3426 746 3427 747
rect 1618 742 1624 743
rect 1822 744 1828 745
rect 3344 744 3427 746
rect 110 739 116 740
rect 1822 740 1823 744
rect 1827 740 1828 744
rect 1822 739 1828 740
rect 1887 743 1893 744
rect 1887 739 1888 743
rect 1892 742 1893 743
rect 1954 743 1960 744
rect 1954 742 1955 743
rect 1892 740 1955 742
rect 1892 739 1893 740
rect 1887 738 1893 739
rect 1954 739 1955 740
rect 1959 739 1960 743
rect 1954 738 1960 739
rect 1983 743 1989 744
rect 1983 739 1984 743
rect 1988 742 1989 743
rect 2063 743 2069 744
rect 2063 742 2064 743
rect 1988 740 2064 742
rect 1988 739 1989 740
rect 1983 738 1989 739
rect 2063 739 2064 740
rect 2068 739 2069 743
rect 2063 738 2069 739
rect 2255 743 2261 744
rect 2255 739 2256 743
rect 2260 742 2261 743
rect 2374 743 2380 744
rect 2374 742 2375 743
rect 2260 740 2375 742
rect 2260 739 2261 740
rect 2255 738 2261 739
rect 2374 739 2375 740
rect 2379 739 2380 743
rect 2374 738 2380 739
rect 2439 743 2445 744
rect 2439 739 2440 743
rect 2444 742 2445 743
rect 2462 743 2468 744
rect 2462 742 2463 743
rect 2444 740 2463 742
rect 2444 739 2445 740
rect 2439 738 2445 739
rect 2462 739 2463 740
rect 2467 739 2468 743
rect 2462 738 2468 739
rect 2615 743 2621 744
rect 2615 739 2616 743
rect 2620 742 2621 743
rect 2646 743 2652 744
rect 2646 742 2647 743
rect 2620 740 2647 742
rect 2620 739 2621 740
rect 2615 738 2621 739
rect 2646 739 2647 740
rect 2651 739 2652 743
rect 2646 738 2652 739
rect 2711 743 2717 744
rect 2711 739 2712 743
rect 2716 742 2717 743
rect 2791 743 2797 744
rect 2791 742 2792 743
rect 2716 740 2792 742
rect 2716 739 2717 740
rect 2711 738 2717 739
rect 2791 739 2792 740
rect 2796 739 2797 743
rect 2791 738 2797 739
rect 2967 743 2973 744
rect 2967 739 2968 743
rect 2972 742 2973 743
rect 3054 743 3060 744
rect 3054 742 3055 743
rect 2972 740 3055 742
rect 2972 739 2973 740
rect 2967 738 2973 739
rect 3054 739 3055 740
rect 3059 739 3060 743
rect 3054 738 3060 739
rect 3143 743 3149 744
rect 3143 739 3144 743
rect 3148 742 3149 743
rect 3158 743 3164 744
rect 3158 742 3159 743
rect 3148 740 3159 742
rect 3148 739 3149 740
rect 3143 738 3149 739
rect 3158 739 3159 740
rect 3163 739 3164 743
rect 3158 738 3164 739
rect 3239 743 3245 744
rect 3239 739 3240 743
rect 3244 742 3245 743
rect 3319 743 3325 744
rect 3319 742 3320 743
rect 3244 740 3320 742
rect 3244 739 3245 740
rect 3239 738 3245 739
rect 3319 739 3320 740
rect 3324 739 3325 743
rect 3426 743 3427 744
rect 3431 743 3432 747
rect 3426 742 3432 743
rect 3471 743 3477 744
rect 3319 738 3325 739
rect 3471 739 3472 743
rect 3476 742 3477 743
rect 3479 743 3485 744
rect 3479 742 3480 743
rect 3476 740 3480 742
rect 3476 739 3477 740
rect 3471 738 3477 739
rect 3479 739 3480 740
rect 3484 739 3485 743
rect 3479 738 3485 739
rect 1894 733 1900 734
rect 142 731 148 732
rect 142 727 143 731
rect 147 727 148 731
rect 142 726 148 727
rect 278 731 284 732
rect 278 727 279 731
rect 283 727 284 731
rect 278 726 284 727
rect 446 731 452 732
rect 446 727 447 731
rect 451 727 452 731
rect 446 726 452 727
rect 614 731 620 732
rect 614 727 615 731
rect 619 727 620 731
rect 614 726 620 727
rect 782 731 788 732
rect 782 727 783 731
rect 787 727 788 731
rect 782 726 788 727
rect 942 731 948 732
rect 942 727 943 731
rect 947 727 948 731
rect 942 726 948 727
rect 1094 731 1100 732
rect 1094 727 1095 731
rect 1099 727 1100 731
rect 1094 726 1100 727
rect 1246 731 1252 732
rect 1246 727 1247 731
rect 1251 727 1252 731
rect 1246 726 1252 727
rect 1398 731 1404 732
rect 1398 727 1399 731
rect 1403 727 1404 731
rect 1398 726 1404 727
rect 1558 731 1564 732
rect 1558 727 1559 731
rect 1563 727 1564 731
rect 1894 729 1895 733
rect 1899 729 1900 733
rect 1894 728 1900 729
rect 2070 733 2076 734
rect 2070 729 2071 733
rect 2075 729 2076 733
rect 2070 728 2076 729
rect 2262 733 2268 734
rect 2262 729 2263 733
rect 2267 729 2268 733
rect 2262 728 2268 729
rect 2446 733 2452 734
rect 2446 729 2447 733
rect 2451 729 2452 733
rect 2446 728 2452 729
rect 2622 733 2628 734
rect 2622 729 2623 733
rect 2627 729 2628 733
rect 2622 728 2628 729
rect 2798 733 2804 734
rect 2798 729 2799 733
rect 2803 729 2804 733
rect 2798 728 2804 729
rect 2974 733 2980 734
rect 2974 729 2975 733
rect 2979 729 2980 733
rect 2974 728 2980 729
rect 3150 733 3156 734
rect 3150 729 3151 733
rect 3155 729 3156 733
rect 3150 728 3156 729
rect 3326 733 3332 734
rect 3326 729 3327 733
rect 3331 729 3332 733
rect 3326 728 3332 729
rect 3486 733 3492 734
rect 3486 729 3487 733
rect 3491 729 3492 733
rect 3486 728 3492 729
rect 1558 726 1564 727
rect 1862 720 1868 721
rect 3574 720 3580 721
rect 135 719 141 720
rect 135 715 136 719
rect 140 718 141 719
rect 202 719 208 720
rect 202 718 203 719
rect 140 716 203 718
rect 140 715 141 716
rect 135 714 141 715
rect 202 715 203 716
rect 207 715 208 719
rect 202 714 208 715
rect 270 719 277 720
rect 270 715 271 719
rect 276 715 277 719
rect 270 714 277 715
rect 439 719 445 720
rect 439 715 440 719
rect 444 718 445 719
rect 506 719 512 720
rect 506 718 507 719
rect 444 716 507 718
rect 444 715 445 716
rect 439 714 445 715
rect 506 715 507 716
rect 511 715 512 719
rect 506 714 512 715
rect 607 719 613 720
rect 607 715 608 719
rect 612 718 613 719
rect 674 719 680 720
rect 674 718 675 719
rect 612 716 675 718
rect 612 715 613 716
rect 607 714 613 715
rect 674 715 675 716
rect 679 715 680 719
rect 674 714 680 715
rect 775 719 781 720
rect 775 715 776 719
rect 780 718 781 719
rect 790 719 796 720
rect 790 718 791 719
rect 780 716 791 718
rect 780 715 781 716
rect 775 714 781 715
rect 790 715 791 716
rect 795 715 796 719
rect 790 714 796 715
rect 935 719 941 720
rect 935 715 936 719
rect 940 718 941 719
rect 943 719 949 720
rect 943 718 944 719
rect 940 716 944 718
rect 940 715 941 716
rect 935 714 941 715
rect 943 715 944 716
rect 948 715 949 719
rect 943 714 949 715
rect 1079 719 1085 720
rect 1079 715 1080 719
rect 1084 718 1085 719
rect 1087 719 1093 720
rect 1087 718 1088 719
rect 1084 716 1088 718
rect 1084 715 1085 716
rect 1079 714 1085 715
rect 1087 715 1088 716
rect 1092 715 1093 719
rect 1087 714 1093 715
rect 1239 719 1245 720
rect 1239 715 1240 719
rect 1244 718 1245 719
rect 1294 719 1300 720
rect 1294 718 1295 719
rect 1244 716 1295 718
rect 1244 715 1245 716
rect 1239 714 1245 715
rect 1294 715 1295 716
rect 1299 715 1300 719
rect 1294 714 1300 715
rect 1383 719 1389 720
rect 1383 715 1384 719
rect 1388 718 1389 719
rect 1391 719 1397 720
rect 1391 718 1392 719
rect 1388 716 1392 718
rect 1388 715 1389 716
rect 1383 714 1389 715
rect 1391 715 1392 716
rect 1396 715 1397 719
rect 1391 714 1397 715
rect 1543 719 1549 720
rect 1543 715 1544 719
rect 1548 718 1549 719
rect 1551 719 1557 720
rect 1551 718 1552 719
rect 1548 716 1552 718
rect 1548 715 1549 716
rect 1543 714 1549 715
rect 1551 715 1552 716
rect 1556 715 1557 719
rect 1862 716 1863 720
rect 1867 716 1868 720
rect 1983 719 1989 720
rect 1983 718 1984 719
rect 1949 716 1984 718
rect 1862 715 1868 716
rect 1983 715 1984 716
rect 1988 715 1989 719
rect 2711 719 2717 720
rect 2711 718 2712 719
rect 2677 716 2712 718
rect 1551 714 1557 715
rect 1983 714 1989 715
rect 2254 715 2260 716
rect 2254 711 2255 715
rect 2259 714 2260 715
rect 2374 715 2380 716
rect 2259 712 2281 714
rect 2259 711 2260 712
rect 2254 710 2260 711
rect 2374 711 2375 715
rect 2379 714 2380 715
rect 2711 715 2712 716
rect 2716 715 2717 719
rect 3239 719 3245 720
rect 3239 718 3240 719
rect 3205 716 3240 718
rect 2711 714 2717 715
rect 3239 715 3240 716
rect 3244 715 3245 719
rect 3574 716 3575 720
rect 3579 716 3580 720
rect 3239 714 3245 715
rect 3258 715 3264 716
rect 3574 715 3580 716
rect 2379 712 2465 714
rect 2379 711 2380 712
rect 2374 710 2380 711
rect 3258 711 3259 715
rect 3263 714 3264 715
rect 3263 712 3345 714
rect 3263 711 3264 712
rect 3258 710 3264 711
rect 127 703 133 704
rect 127 699 128 703
rect 132 702 133 703
rect 135 703 141 704
rect 135 702 136 703
rect 132 700 136 702
rect 132 699 133 700
rect 127 698 133 699
rect 135 699 136 700
rect 140 699 141 703
rect 135 698 141 699
rect 214 703 220 704
rect 214 699 215 703
rect 219 702 220 703
rect 279 703 285 704
rect 279 702 280 703
rect 219 700 280 702
rect 219 699 220 700
rect 214 698 220 699
rect 279 699 280 700
rect 284 699 285 703
rect 279 698 285 699
rect 431 703 437 704
rect 431 699 432 703
rect 436 702 437 703
rect 447 703 453 704
rect 447 702 448 703
rect 436 700 448 702
rect 436 699 437 700
rect 431 698 437 699
rect 447 699 448 700
rect 452 699 453 703
rect 447 698 453 699
rect 526 703 532 704
rect 526 699 527 703
rect 531 702 532 703
rect 615 703 621 704
rect 615 702 616 703
rect 531 700 616 702
rect 531 699 532 700
rect 526 698 532 699
rect 615 699 616 700
rect 620 699 621 703
rect 615 698 621 699
rect 710 703 716 704
rect 710 699 711 703
rect 715 702 716 703
rect 783 703 789 704
rect 783 702 784 703
rect 715 700 784 702
rect 715 699 716 700
rect 710 698 716 699
rect 783 699 784 700
rect 788 699 789 703
rect 783 698 789 699
rect 951 703 957 704
rect 951 699 952 703
rect 956 702 957 703
rect 1026 703 1032 704
rect 1026 702 1027 703
rect 956 700 1027 702
rect 956 699 957 700
rect 951 698 957 699
rect 1026 699 1027 700
rect 1031 699 1032 703
rect 1026 698 1032 699
rect 1103 703 1109 704
rect 1103 699 1104 703
rect 1108 702 1109 703
rect 1111 703 1117 704
rect 1111 702 1112 703
rect 1108 700 1112 702
rect 1108 699 1109 700
rect 1103 698 1109 699
rect 1111 699 1112 700
rect 1116 699 1117 703
rect 1111 698 1117 699
rect 1271 703 1277 704
rect 1271 699 1272 703
rect 1276 702 1277 703
rect 1362 703 1368 704
rect 1362 702 1363 703
rect 1276 700 1363 702
rect 1276 699 1277 700
rect 1271 698 1277 699
rect 1362 699 1363 700
rect 1367 699 1368 703
rect 1362 698 1368 699
rect 1431 703 1437 704
rect 1431 699 1432 703
rect 1436 702 1437 703
rect 1514 703 1520 704
rect 1514 702 1515 703
rect 1436 700 1515 702
rect 1436 699 1437 700
rect 1431 698 1437 699
rect 1514 699 1515 700
rect 1519 699 1520 703
rect 1514 698 1520 699
rect 1591 703 1597 704
rect 1591 699 1592 703
rect 1596 702 1597 703
rect 1618 703 1624 704
rect 1618 702 1619 703
rect 1596 700 1619 702
rect 1596 699 1597 700
rect 1591 698 1597 699
rect 1618 699 1619 700
rect 1623 699 1624 703
rect 1618 698 1624 699
rect 1862 703 1868 704
rect 1862 699 1863 703
rect 1867 699 1868 703
rect 2927 703 2933 704
rect 2927 702 2928 703
rect 2849 700 2928 702
rect 1862 698 1868 699
rect 2927 699 2928 700
rect 2932 699 2933 703
rect 3471 703 3477 704
rect 2927 698 2933 699
rect 2936 700 2985 702
rect 142 693 148 694
rect 142 689 143 693
rect 147 689 148 693
rect 142 688 148 689
rect 286 693 292 694
rect 286 689 287 693
rect 291 689 292 693
rect 286 688 292 689
rect 454 693 460 694
rect 454 689 455 693
rect 459 689 460 693
rect 454 688 460 689
rect 622 693 628 694
rect 622 689 623 693
rect 627 689 628 693
rect 622 688 628 689
rect 790 693 796 694
rect 790 689 791 693
rect 795 689 796 693
rect 790 688 796 689
rect 958 693 964 694
rect 958 689 959 693
rect 963 689 964 693
rect 958 688 964 689
rect 1118 693 1124 694
rect 1118 689 1119 693
rect 1123 689 1124 693
rect 1118 688 1124 689
rect 1278 693 1284 694
rect 1278 689 1279 693
rect 1283 689 1284 693
rect 1278 688 1284 689
rect 1438 693 1444 694
rect 1438 689 1439 693
rect 1443 689 1444 693
rect 1438 688 1444 689
rect 1598 693 1604 694
rect 1598 689 1599 693
rect 1603 689 1604 693
rect 1598 688 1604 689
rect 1886 693 1892 694
rect 1886 689 1887 693
rect 1891 689 1892 693
rect 1886 688 1892 689
rect 2062 693 2068 694
rect 2062 689 2063 693
rect 2067 689 2068 693
rect 2062 688 2068 689
rect 2254 693 2260 694
rect 2254 689 2255 693
rect 2259 689 2260 693
rect 2254 688 2260 689
rect 2438 693 2444 694
rect 2438 689 2439 693
rect 2443 689 2444 693
rect 2438 688 2444 689
rect 2614 693 2620 694
rect 2614 689 2615 693
rect 2619 689 2620 693
rect 2614 688 2620 689
rect 2790 693 2796 694
rect 2790 689 2791 693
rect 2795 689 2796 693
rect 2790 688 2796 689
rect 2110 687 2117 688
rect 2110 683 2111 687
rect 2116 683 2117 687
rect 2110 682 2117 683
rect 2646 687 2652 688
rect 2646 683 2647 687
rect 2651 686 2652 687
rect 2936 686 2938 700
rect 3471 699 3472 703
rect 3476 702 3477 703
rect 3574 703 3580 704
rect 3476 700 3497 702
rect 3476 699 3477 700
rect 3471 698 3477 699
rect 3574 699 3575 703
rect 3579 699 3580 703
rect 3574 698 3580 699
rect 2966 693 2972 694
rect 2966 689 2967 693
rect 2971 689 2972 693
rect 2966 688 2972 689
rect 3142 693 3148 694
rect 3142 689 3143 693
rect 3147 689 3148 693
rect 3142 688 3148 689
rect 3318 693 3324 694
rect 3318 689 3319 693
rect 3323 689 3324 693
rect 3318 688 3324 689
rect 3478 693 3484 694
rect 3478 689 3479 693
rect 3483 689 3484 693
rect 3478 688 3484 689
rect 2651 684 2938 686
rect 2651 683 2652 684
rect 2646 682 2652 683
rect 110 680 116 681
rect 1822 680 1828 681
rect 110 676 111 680
rect 115 676 116 680
rect 214 679 220 680
rect 214 678 215 679
rect 197 676 215 678
rect 110 675 116 676
rect 214 675 215 676
rect 219 675 220 679
rect 526 679 532 680
rect 526 678 527 679
rect 509 676 527 678
rect 214 674 220 675
rect 270 675 276 676
rect 270 671 271 675
rect 275 674 276 675
rect 526 675 527 676
rect 531 675 532 679
rect 710 679 716 680
rect 710 678 711 679
rect 677 676 711 678
rect 526 674 532 675
rect 710 675 711 676
rect 715 675 716 679
rect 1822 676 1823 680
rect 1827 676 1828 680
rect 710 674 716 675
rect 943 675 949 676
rect 275 672 305 674
rect 275 671 276 672
rect 270 670 276 671
rect 943 671 944 675
rect 948 674 949 675
rect 1026 675 1032 676
rect 948 672 977 674
rect 948 671 949 672
rect 943 670 949 671
rect 1026 671 1027 675
rect 1031 674 1032 675
rect 1362 675 1368 676
rect 1031 672 1137 674
rect 1031 671 1032 672
rect 1026 670 1032 671
rect 1362 671 1363 675
rect 1367 674 1368 675
rect 1514 675 1520 676
rect 1822 675 1828 676
rect 1367 672 1457 674
rect 1367 671 1368 672
rect 1362 670 1368 671
rect 1514 671 1515 675
rect 1519 674 1520 675
rect 1519 672 1617 674
rect 1519 671 1520 672
rect 1514 670 1520 671
rect 1886 667 1892 668
rect 110 663 116 664
rect 110 659 111 663
rect 115 659 116 663
rect 110 658 116 659
rect 790 663 796 664
rect 790 659 791 663
rect 795 662 796 663
rect 1263 663 1269 664
rect 795 660 801 662
rect 795 659 796 660
rect 790 658 796 659
rect 1263 659 1264 663
rect 1268 662 1269 663
rect 1822 663 1828 664
rect 1268 660 1289 662
rect 1268 659 1269 660
rect 1263 658 1269 659
rect 1822 659 1823 663
rect 1827 659 1828 663
rect 1886 663 1887 667
rect 1891 663 1892 667
rect 1886 662 1892 663
rect 1974 667 1980 668
rect 1974 663 1975 667
rect 1979 663 1980 667
rect 1974 662 1980 663
rect 2094 667 2100 668
rect 2094 663 2095 667
rect 2099 663 2100 667
rect 2094 662 2100 663
rect 2222 667 2228 668
rect 2222 663 2223 667
rect 2227 663 2228 667
rect 2222 662 2228 663
rect 2350 667 2356 668
rect 2350 663 2351 667
rect 2355 663 2356 667
rect 2350 662 2356 663
rect 2478 667 2484 668
rect 2478 663 2479 667
rect 2483 663 2484 667
rect 2478 662 2484 663
rect 2614 667 2620 668
rect 2614 663 2615 667
rect 2619 663 2620 667
rect 2614 662 2620 663
rect 2766 667 2772 668
rect 2766 663 2767 667
rect 2771 663 2772 667
rect 2766 662 2772 663
rect 2934 667 2940 668
rect 2934 663 2935 667
rect 2939 663 2940 667
rect 2934 662 2940 663
rect 3118 667 3124 668
rect 3118 663 3119 667
rect 3123 663 3124 667
rect 3118 662 3124 663
rect 3310 667 3316 668
rect 3310 663 3311 667
rect 3315 663 3316 667
rect 3310 662 3316 663
rect 3478 667 3484 668
rect 3478 663 3479 667
rect 3483 663 3484 667
rect 3478 662 3484 663
rect 1822 658 1828 659
rect 2462 659 2468 660
rect 1862 657 1868 658
rect 134 653 140 654
rect 134 649 135 653
rect 139 649 140 653
rect 134 648 140 649
rect 278 653 284 654
rect 278 649 279 653
rect 283 649 284 653
rect 278 648 284 649
rect 446 653 452 654
rect 446 649 447 653
rect 451 649 452 653
rect 446 648 452 649
rect 614 653 620 654
rect 614 649 615 653
rect 619 649 620 653
rect 614 648 620 649
rect 782 653 788 654
rect 782 649 783 653
rect 787 649 788 653
rect 782 648 788 649
rect 950 653 956 654
rect 950 649 951 653
rect 955 649 956 653
rect 950 648 956 649
rect 1110 653 1116 654
rect 1110 649 1111 653
rect 1115 649 1116 653
rect 1110 648 1116 649
rect 1270 653 1276 654
rect 1270 649 1271 653
rect 1275 649 1276 653
rect 1270 648 1276 649
rect 1430 653 1436 654
rect 1430 649 1431 653
rect 1435 649 1436 653
rect 1430 648 1436 649
rect 1590 653 1596 654
rect 1590 649 1591 653
rect 1595 649 1596 653
rect 1862 653 1863 657
rect 1867 653 1868 657
rect 2462 655 2463 659
rect 2467 658 2468 659
rect 2467 656 2497 658
rect 3574 657 3580 658
rect 2467 655 2468 656
rect 2462 654 2468 655
rect 1862 652 1868 653
rect 3574 653 3575 657
rect 3579 653 3580 657
rect 3574 652 3580 653
rect 1590 648 1596 649
rect 1879 643 1885 644
rect 1862 640 1868 641
rect 1862 636 1863 640
rect 1867 636 1868 640
rect 1879 639 1880 643
rect 1884 642 1885 643
rect 1954 643 1960 644
rect 1884 640 1913 642
rect 1884 639 1885 640
rect 1879 638 1885 639
rect 1954 639 1955 643
rect 1959 642 1960 643
rect 2042 643 2048 644
rect 1959 640 2001 642
rect 1959 639 1960 640
rect 1954 638 1960 639
rect 2042 639 2043 643
rect 2047 642 2048 643
rect 2343 643 2349 644
rect 2343 642 2344 643
rect 2047 640 2121 642
rect 2285 640 2344 642
rect 2047 639 2048 640
rect 2042 638 2048 639
rect 2343 639 2344 640
rect 2348 639 2349 643
rect 2471 643 2477 644
rect 2471 642 2472 643
rect 2413 640 2472 642
rect 2343 638 2349 639
rect 2471 639 2472 640
rect 2476 639 2477 643
rect 2759 643 2765 644
rect 2759 642 2760 643
rect 2677 640 2760 642
rect 2471 638 2477 639
rect 2759 639 2760 640
rect 2764 639 2765 643
rect 2834 643 2840 644
rect 2834 642 2835 643
rect 2829 640 2835 642
rect 2759 638 2765 639
rect 2834 639 2835 640
rect 2839 639 2840 643
rect 3111 643 3117 644
rect 3111 642 3112 643
rect 2997 640 3112 642
rect 2834 638 2840 639
rect 3111 639 3112 640
rect 3116 639 3117 643
rect 3226 643 3232 644
rect 3226 642 3227 643
rect 3181 640 3227 642
rect 3111 638 3117 639
rect 3226 639 3227 640
rect 3231 639 3232 643
rect 3226 638 3232 639
rect 3234 643 3240 644
rect 3234 639 3235 643
rect 3239 642 3240 643
rect 3470 643 3476 644
rect 3239 640 3337 642
rect 3239 639 3240 640
rect 3234 638 3240 639
rect 3470 639 3471 643
rect 3475 642 3476 643
rect 3475 640 3505 642
rect 3574 640 3580 641
rect 3475 639 3476 640
rect 3470 638 3476 639
rect 1862 635 1868 636
rect 3574 636 3575 640
rect 3579 636 3580 640
rect 3574 635 3580 636
rect 1894 627 1900 628
rect 134 623 140 624
rect 134 619 135 623
rect 139 619 140 623
rect 134 618 140 619
rect 286 623 292 624
rect 286 619 287 623
rect 291 619 292 623
rect 286 618 292 619
rect 454 623 460 624
rect 454 619 455 623
rect 459 619 460 623
rect 454 618 460 619
rect 630 623 636 624
rect 630 619 631 623
rect 635 619 636 623
rect 630 618 636 619
rect 798 623 804 624
rect 798 619 799 623
rect 803 619 804 623
rect 798 618 804 619
rect 966 623 972 624
rect 966 619 967 623
rect 971 619 972 623
rect 966 618 972 619
rect 1118 623 1124 624
rect 1118 619 1119 623
rect 1123 619 1124 623
rect 1118 618 1124 619
rect 1270 623 1276 624
rect 1270 619 1271 623
rect 1275 619 1276 623
rect 1270 618 1276 619
rect 1414 623 1420 624
rect 1414 619 1415 623
rect 1419 619 1420 623
rect 1414 618 1420 619
rect 1558 623 1564 624
rect 1558 619 1559 623
rect 1563 619 1564 623
rect 1558 618 1564 619
rect 1710 623 1716 624
rect 1710 619 1711 623
rect 1715 619 1716 623
rect 1894 623 1895 627
rect 1899 623 1900 627
rect 1894 622 1900 623
rect 1982 627 1988 628
rect 1982 623 1983 627
rect 1987 623 1988 627
rect 1982 622 1988 623
rect 2102 627 2108 628
rect 2102 623 2103 627
rect 2107 623 2108 627
rect 2102 622 2108 623
rect 2230 627 2236 628
rect 2230 623 2231 627
rect 2235 623 2236 627
rect 2230 622 2236 623
rect 2358 627 2364 628
rect 2358 623 2359 627
rect 2363 623 2364 627
rect 2358 622 2364 623
rect 2486 627 2492 628
rect 2486 623 2487 627
rect 2491 623 2492 627
rect 2486 622 2492 623
rect 2622 627 2628 628
rect 2622 623 2623 627
rect 2627 623 2628 627
rect 2622 622 2628 623
rect 2774 627 2780 628
rect 2774 623 2775 627
rect 2779 623 2780 627
rect 2774 622 2780 623
rect 2942 627 2948 628
rect 2942 623 2943 627
rect 2947 623 2948 627
rect 2942 622 2948 623
rect 3126 627 3132 628
rect 3126 623 3127 627
rect 3131 623 3132 627
rect 3126 622 3132 623
rect 3318 627 3324 628
rect 3318 623 3319 627
rect 3323 623 3324 627
rect 3318 622 3324 623
rect 3486 627 3492 628
rect 3486 623 3487 627
rect 3491 623 3492 627
rect 3486 622 3492 623
rect 1710 618 1716 619
rect 127 615 133 616
rect 110 613 116 614
rect 110 609 111 613
rect 115 609 116 613
rect 127 611 128 615
rect 132 614 133 615
rect 1103 615 1109 616
rect 132 612 153 614
rect 132 611 133 612
rect 127 610 133 611
rect 1103 611 1104 615
rect 1108 614 1109 615
rect 1638 615 1644 616
rect 1108 612 1137 614
rect 1108 611 1109 612
rect 1103 610 1109 611
rect 1638 611 1639 615
rect 1643 614 1644 615
rect 1887 615 1893 616
rect 1643 612 1729 614
rect 1822 613 1828 614
rect 1643 611 1644 612
rect 1638 610 1644 611
rect 110 608 116 609
rect 1822 609 1823 613
rect 1827 609 1828 613
rect 1887 611 1888 615
rect 1892 614 1893 615
rect 1954 615 1960 616
rect 1954 614 1955 615
rect 1892 612 1955 614
rect 1892 611 1893 612
rect 1887 610 1893 611
rect 1954 611 1955 612
rect 1959 611 1960 615
rect 1954 610 1960 611
rect 1975 615 1981 616
rect 1975 611 1976 615
rect 1980 614 1981 615
rect 2042 615 2048 616
rect 2042 614 2043 615
rect 1980 612 2043 614
rect 1980 611 1981 612
rect 1975 610 1981 611
rect 2042 611 2043 612
rect 2047 611 2048 615
rect 2042 610 2048 611
rect 2095 615 2101 616
rect 2095 611 2096 615
rect 2100 614 2101 615
rect 2110 615 2116 616
rect 2110 614 2111 615
rect 2100 612 2111 614
rect 2100 611 2101 612
rect 2095 610 2101 611
rect 2110 611 2111 612
rect 2115 611 2116 615
rect 2110 610 2116 611
rect 2206 615 2212 616
rect 2206 611 2207 615
rect 2211 614 2212 615
rect 2223 615 2229 616
rect 2223 614 2224 615
rect 2211 612 2224 614
rect 2211 611 2212 612
rect 2206 610 2212 611
rect 2223 611 2224 612
rect 2228 611 2229 615
rect 2223 610 2229 611
rect 2343 615 2349 616
rect 2343 611 2344 615
rect 2348 614 2349 615
rect 2351 615 2357 616
rect 2351 614 2352 615
rect 2348 612 2352 614
rect 2348 611 2349 612
rect 2343 610 2349 611
rect 2351 611 2352 612
rect 2356 611 2357 615
rect 2351 610 2357 611
rect 2471 615 2477 616
rect 2471 611 2472 615
rect 2476 614 2477 615
rect 2479 615 2485 616
rect 2479 614 2480 615
rect 2476 612 2480 614
rect 2476 611 2477 612
rect 2471 610 2477 611
rect 2479 611 2480 612
rect 2484 611 2485 615
rect 2479 610 2485 611
rect 2615 615 2621 616
rect 2615 611 2616 615
rect 2620 614 2621 615
rect 2630 615 2636 616
rect 2630 614 2631 615
rect 2620 612 2631 614
rect 2620 611 2621 612
rect 2615 610 2621 611
rect 2630 611 2631 612
rect 2635 611 2636 615
rect 2630 610 2636 611
rect 2759 615 2765 616
rect 2759 611 2760 615
rect 2764 614 2765 615
rect 2767 615 2773 616
rect 2767 614 2768 615
rect 2764 612 2768 614
rect 2764 611 2765 612
rect 2759 610 2765 611
rect 2767 611 2768 612
rect 2772 611 2773 615
rect 2767 610 2773 611
rect 2927 615 2933 616
rect 2927 611 2928 615
rect 2932 614 2933 615
rect 2935 615 2941 616
rect 2935 614 2936 615
rect 2932 612 2936 614
rect 2932 611 2933 612
rect 2927 610 2933 611
rect 2935 611 2936 612
rect 2940 611 2941 615
rect 2935 610 2941 611
rect 3111 615 3117 616
rect 3111 611 3112 615
rect 3116 614 3117 615
rect 3119 615 3125 616
rect 3119 614 3120 615
rect 3116 612 3120 614
rect 3116 611 3117 612
rect 3111 610 3117 611
rect 3119 611 3120 612
rect 3124 611 3125 615
rect 3119 610 3125 611
rect 3226 615 3232 616
rect 3226 611 3227 615
rect 3231 614 3232 615
rect 3311 615 3317 616
rect 3311 614 3312 615
rect 3231 612 3312 614
rect 3231 611 3232 612
rect 3226 610 3232 611
rect 3311 611 3312 612
rect 3316 611 3317 615
rect 3311 610 3317 611
rect 3471 615 3477 616
rect 3471 611 3472 615
rect 3476 614 3477 615
rect 3479 615 3485 616
rect 3479 614 3480 615
rect 3476 612 3480 614
rect 3476 611 3477 612
rect 3471 610 3477 611
rect 3479 611 3480 612
rect 3484 611 3485 615
rect 3479 610 3485 611
rect 1822 608 1828 609
rect 3175 607 3181 608
rect 3175 606 3176 607
rect 2784 604 3176 606
rect 202 599 208 600
rect 110 596 116 597
rect 110 592 111 596
rect 115 592 116 596
rect 202 595 203 599
rect 207 598 208 599
rect 447 599 453 600
rect 207 596 313 598
rect 207 595 208 596
rect 202 594 208 595
rect 447 595 448 599
rect 452 598 453 599
rect 522 599 528 600
rect 452 596 481 598
rect 452 595 453 596
rect 447 594 453 595
rect 522 595 523 599
rect 527 598 528 599
rect 698 599 704 600
rect 527 596 657 598
rect 527 595 528 596
rect 522 594 528 595
rect 698 595 699 599
rect 703 598 704 599
rect 1111 599 1117 600
rect 1111 598 1112 599
rect 703 596 825 598
rect 1029 596 1112 598
rect 703 595 704 596
rect 698 594 704 595
rect 1111 595 1112 596
rect 1116 595 1117 599
rect 1407 599 1413 600
rect 1407 598 1408 599
rect 1333 596 1408 598
rect 1111 594 1117 595
rect 1407 595 1408 596
rect 1412 595 1413 599
rect 1551 599 1557 600
rect 1551 598 1552 599
rect 1477 596 1552 598
rect 1407 594 1413 595
rect 1551 595 1552 596
rect 1556 595 1557 599
rect 1703 599 1709 600
rect 1703 598 1704 599
rect 1621 596 1704 598
rect 1551 594 1557 595
rect 1703 595 1704 596
rect 1708 595 1709 599
rect 1879 599 1885 600
rect 1703 594 1709 595
rect 1822 596 1828 597
rect 110 591 116 592
rect 1822 592 1823 596
rect 1827 592 1828 596
rect 1879 595 1880 599
rect 1884 598 1885 599
rect 1887 599 1893 600
rect 1887 598 1888 599
rect 1884 596 1888 598
rect 1884 595 1885 596
rect 1879 594 1885 595
rect 1887 595 1888 596
rect 1892 595 1893 599
rect 1887 594 1893 595
rect 2039 599 2045 600
rect 2039 595 2040 599
rect 2044 598 2045 599
rect 2054 599 2060 600
rect 2054 598 2055 599
rect 2044 596 2055 598
rect 2044 595 2045 596
rect 2039 594 2045 595
rect 2054 595 2055 596
rect 2059 595 2060 599
rect 2054 594 2060 595
rect 2127 599 2133 600
rect 2127 595 2128 599
rect 2132 598 2133 599
rect 2207 599 2213 600
rect 2207 598 2208 599
rect 2132 596 2208 598
rect 2132 595 2133 596
rect 2127 594 2133 595
rect 2207 595 2208 596
rect 2212 595 2213 599
rect 2207 594 2213 595
rect 2383 599 2389 600
rect 2383 595 2384 599
rect 2388 598 2389 599
rect 2487 599 2493 600
rect 2487 598 2488 599
rect 2388 596 2488 598
rect 2388 595 2389 596
rect 2383 594 2389 595
rect 2487 595 2488 596
rect 2492 595 2493 599
rect 2487 594 2493 595
rect 2575 599 2581 600
rect 2575 595 2576 599
rect 2580 598 2581 599
rect 2784 598 2786 604
rect 3175 603 3176 604
rect 3180 603 3181 607
rect 3175 602 3181 603
rect 2580 596 2786 598
rect 2791 599 2797 600
rect 2580 595 2581 596
rect 2575 594 2581 595
rect 2791 595 2792 599
rect 2796 598 2797 599
rect 2834 599 2840 600
rect 2834 598 2835 599
rect 2796 596 2835 598
rect 2796 595 2797 596
rect 2791 594 2797 595
rect 2834 595 2835 596
rect 2839 595 2840 599
rect 2834 594 2840 595
rect 2911 599 2917 600
rect 2911 595 2912 599
rect 2916 598 2917 599
rect 3015 599 3021 600
rect 3015 598 3016 599
rect 2916 596 3016 598
rect 2916 595 2917 596
rect 2911 594 2917 595
rect 3015 595 3016 596
rect 3020 595 3021 599
rect 3015 594 3021 595
rect 3087 599 3093 600
rect 3087 595 3088 599
rect 3092 598 3093 599
rect 3247 599 3253 600
rect 3247 598 3248 599
rect 3092 596 3248 598
rect 3092 595 3093 596
rect 3087 594 3093 595
rect 3247 595 3248 596
rect 3252 595 3253 599
rect 3247 594 3253 595
rect 3470 599 3476 600
rect 3470 595 3471 599
rect 3475 598 3476 599
rect 3479 599 3485 600
rect 3479 598 3480 599
rect 3475 596 3480 598
rect 3475 595 3476 596
rect 3470 594 3476 595
rect 3479 595 3480 596
rect 3484 595 3485 599
rect 3479 594 3485 595
rect 1822 591 1828 592
rect 1894 589 1900 590
rect 1894 585 1895 589
rect 1899 585 1900 589
rect 1894 584 1900 585
rect 2046 589 2052 590
rect 2046 585 2047 589
rect 2051 585 2052 589
rect 2046 584 2052 585
rect 2214 589 2220 590
rect 2214 585 2215 589
rect 2219 585 2220 589
rect 2214 584 2220 585
rect 2390 589 2396 590
rect 2390 585 2391 589
rect 2395 585 2396 589
rect 2390 584 2396 585
rect 2582 589 2588 590
rect 2582 585 2583 589
rect 2587 585 2588 589
rect 2582 584 2588 585
rect 2798 589 2804 590
rect 2798 585 2799 589
rect 2803 585 2804 589
rect 2798 584 2804 585
rect 3022 589 3028 590
rect 3022 585 3023 589
rect 3027 585 3028 589
rect 3022 584 3028 585
rect 3254 589 3260 590
rect 3254 585 3255 589
rect 3259 585 3260 589
rect 3254 584 3260 585
rect 3486 589 3492 590
rect 3486 585 3487 589
rect 3491 585 3492 589
rect 3486 584 3492 585
rect 142 583 148 584
rect 142 579 143 583
rect 147 579 148 583
rect 142 578 148 579
rect 294 583 300 584
rect 294 579 295 583
rect 299 579 300 583
rect 294 578 300 579
rect 462 583 468 584
rect 462 579 463 583
rect 467 579 468 583
rect 462 578 468 579
rect 638 583 644 584
rect 638 579 639 583
rect 643 579 644 583
rect 638 578 644 579
rect 806 583 812 584
rect 806 579 807 583
rect 811 579 812 583
rect 806 578 812 579
rect 974 583 980 584
rect 974 579 975 583
rect 979 579 980 583
rect 974 578 980 579
rect 1126 583 1132 584
rect 1126 579 1127 583
rect 1131 579 1132 583
rect 1126 578 1132 579
rect 1278 583 1284 584
rect 1278 579 1279 583
rect 1283 579 1284 583
rect 1278 578 1284 579
rect 1422 583 1428 584
rect 1422 579 1423 583
rect 1427 579 1428 583
rect 1422 578 1428 579
rect 1566 583 1572 584
rect 1566 579 1567 583
rect 1571 579 1572 583
rect 1566 578 1572 579
rect 1718 583 1724 584
rect 1718 579 1719 583
rect 1723 579 1724 583
rect 1718 578 1724 579
rect 1862 576 1868 577
rect 3574 576 3580 577
rect 1862 572 1863 576
rect 1867 572 1868 576
rect 2127 575 2133 576
rect 2127 574 2128 575
rect 2101 572 2128 574
rect 135 571 141 572
rect 135 567 136 571
rect 140 570 141 571
rect 202 571 208 572
rect 202 570 203 571
rect 140 568 203 570
rect 140 567 141 568
rect 135 566 141 567
rect 202 567 203 568
rect 207 567 208 571
rect 202 566 208 567
rect 287 571 293 572
rect 287 567 288 571
rect 292 570 293 571
rect 295 571 301 572
rect 295 570 296 571
rect 292 568 296 570
rect 292 567 293 568
rect 287 566 293 567
rect 295 567 296 568
rect 300 567 301 571
rect 295 566 301 567
rect 455 571 461 572
rect 455 567 456 571
rect 460 570 461 571
rect 522 571 528 572
rect 522 570 523 571
rect 460 568 523 570
rect 460 567 461 568
rect 455 566 461 567
rect 522 567 523 568
rect 527 567 528 571
rect 522 566 528 567
rect 631 571 637 572
rect 631 567 632 571
rect 636 570 637 571
rect 698 571 704 572
rect 698 570 699 571
rect 636 568 699 570
rect 636 567 637 568
rect 631 566 637 567
rect 698 567 699 568
rect 703 567 704 571
rect 698 566 704 567
rect 790 571 796 572
rect 790 567 791 571
rect 795 570 796 571
rect 799 571 805 572
rect 799 570 800 571
rect 795 568 800 570
rect 795 567 796 568
rect 790 566 796 567
rect 799 567 800 568
rect 804 567 805 571
rect 799 566 805 567
rect 967 571 973 572
rect 967 567 968 571
rect 972 570 973 571
rect 986 571 992 572
rect 986 570 987 571
rect 972 568 987 570
rect 972 567 973 568
rect 967 566 973 567
rect 986 567 987 568
rect 991 567 992 571
rect 986 566 992 567
rect 1111 571 1117 572
rect 1111 567 1112 571
rect 1116 570 1117 571
rect 1119 571 1125 572
rect 1119 570 1120 571
rect 1116 568 1120 570
rect 1116 567 1117 568
rect 1111 566 1117 567
rect 1119 567 1120 568
rect 1124 567 1125 571
rect 1119 566 1125 567
rect 1263 571 1269 572
rect 1263 567 1264 571
rect 1268 570 1269 571
rect 1271 571 1277 572
rect 1271 570 1272 571
rect 1268 568 1272 570
rect 1268 567 1269 568
rect 1263 566 1269 567
rect 1271 567 1272 568
rect 1276 567 1277 571
rect 1271 566 1277 567
rect 1407 571 1413 572
rect 1407 567 1408 571
rect 1412 570 1413 571
rect 1415 571 1421 572
rect 1415 570 1416 571
rect 1412 568 1416 570
rect 1412 567 1413 568
rect 1407 566 1413 567
rect 1415 567 1416 568
rect 1420 567 1421 571
rect 1415 566 1421 567
rect 1551 571 1557 572
rect 1551 567 1552 571
rect 1556 570 1557 571
rect 1559 571 1565 572
rect 1559 570 1560 571
rect 1556 568 1560 570
rect 1556 567 1557 568
rect 1551 566 1557 567
rect 1559 567 1560 568
rect 1564 567 1565 571
rect 1559 566 1565 567
rect 1703 571 1709 572
rect 1703 567 1704 571
rect 1708 570 1709 571
rect 1711 571 1717 572
rect 1862 571 1868 572
rect 2127 571 2128 572
rect 2132 571 2133 575
rect 2911 575 2917 576
rect 2911 574 2912 575
rect 2853 572 2912 574
rect 1711 570 1712 571
rect 1708 568 1712 570
rect 1708 567 1709 568
rect 1703 566 1709 567
rect 1711 567 1712 568
rect 1716 567 1717 571
rect 2127 570 2133 571
rect 2206 571 2212 572
rect 1711 566 1717 567
rect 2206 567 2207 571
rect 2211 570 2212 571
rect 2487 571 2493 572
rect 2211 568 2233 570
rect 2211 567 2212 568
rect 2206 566 2212 567
rect 2487 567 2488 571
rect 2492 570 2493 571
rect 2911 571 2912 572
rect 2916 571 2917 575
rect 3087 575 3093 576
rect 3087 574 3088 575
rect 3077 572 3088 574
rect 2911 570 2917 571
rect 3087 571 3088 572
rect 3092 571 3093 575
rect 3574 572 3575 576
rect 3579 572 3580 576
rect 3087 570 3093 571
rect 3175 571 3181 572
rect 2492 568 2601 570
rect 2492 567 2493 568
rect 2487 566 2493 567
rect 3175 567 3176 571
rect 3180 570 3181 571
rect 3463 571 3469 572
rect 3574 571 3580 572
rect 3180 568 3273 570
rect 3180 567 3181 568
rect 3175 566 3181 567
rect 3463 567 3464 571
rect 3468 570 3469 571
rect 3468 568 3505 570
rect 3468 567 3469 568
rect 3463 566 3469 567
rect 1862 559 1868 560
rect 135 555 141 556
rect 135 551 136 555
rect 140 554 141 555
rect 143 555 149 556
rect 143 554 144 555
rect 140 552 144 554
rect 140 551 141 552
rect 135 550 141 551
rect 143 551 144 552
rect 148 551 149 555
rect 143 550 149 551
rect 231 555 237 556
rect 231 551 232 555
rect 236 554 237 555
rect 303 555 309 556
rect 303 554 304 555
rect 236 552 304 554
rect 236 551 237 552
rect 231 550 237 551
rect 303 551 304 552
rect 308 551 309 555
rect 303 550 309 551
rect 447 555 453 556
rect 447 551 448 555
rect 452 554 453 555
rect 463 555 469 556
rect 463 554 464 555
rect 452 552 464 554
rect 452 551 453 552
rect 447 550 453 551
rect 463 551 464 552
rect 468 551 469 555
rect 463 550 469 551
rect 551 555 557 556
rect 551 551 552 555
rect 556 554 557 555
rect 623 555 629 556
rect 623 554 624 555
rect 556 552 624 554
rect 556 551 557 552
rect 551 550 557 551
rect 623 551 624 552
rect 628 551 629 555
rect 623 550 629 551
rect 703 555 709 556
rect 703 551 704 555
rect 708 554 709 555
rect 775 555 781 556
rect 775 554 776 555
rect 708 552 776 554
rect 708 551 709 552
rect 703 550 709 551
rect 775 551 776 552
rect 780 551 781 555
rect 775 550 781 551
rect 919 555 925 556
rect 919 551 920 555
rect 924 554 925 555
rect 994 555 1000 556
rect 994 554 995 555
rect 924 552 995 554
rect 924 551 925 552
rect 919 550 925 551
rect 994 551 995 552
rect 999 551 1000 555
rect 994 550 1000 551
rect 1055 555 1061 556
rect 1055 551 1056 555
rect 1060 554 1061 555
rect 1074 555 1080 556
rect 1074 554 1075 555
rect 1060 552 1075 554
rect 1060 551 1061 552
rect 1055 550 1061 551
rect 1074 551 1075 552
rect 1079 551 1080 555
rect 1074 550 1080 551
rect 1183 555 1189 556
rect 1183 551 1184 555
rect 1188 554 1189 555
rect 1198 555 1204 556
rect 1198 554 1199 555
rect 1188 552 1199 554
rect 1188 551 1189 552
rect 1183 550 1189 551
rect 1198 551 1199 552
rect 1203 551 1204 555
rect 1198 550 1204 551
rect 1255 555 1261 556
rect 1255 551 1256 555
rect 1260 554 1261 555
rect 1303 555 1309 556
rect 1303 554 1304 555
rect 1260 552 1304 554
rect 1260 551 1261 552
rect 1255 550 1261 551
rect 1303 551 1304 552
rect 1308 551 1309 555
rect 1303 550 1309 551
rect 1375 555 1381 556
rect 1375 551 1376 555
rect 1380 554 1381 555
rect 1415 555 1421 556
rect 1415 554 1416 555
rect 1380 552 1416 554
rect 1380 551 1381 552
rect 1375 550 1381 551
rect 1415 551 1416 552
rect 1420 551 1421 555
rect 1415 550 1421 551
rect 1527 555 1533 556
rect 1527 551 1528 555
rect 1532 554 1533 555
rect 1602 555 1608 556
rect 1602 554 1603 555
rect 1532 552 1603 554
rect 1532 551 1533 552
rect 1527 550 1533 551
rect 1602 551 1603 552
rect 1607 551 1608 555
rect 1602 550 1608 551
rect 1639 555 1645 556
rect 1639 551 1640 555
rect 1644 554 1645 555
rect 1670 555 1676 556
rect 1670 554 1671 555
rect 1644 552 1671 554
rect 1644 551 1645 552
rect 1639 550 1645 551
rect 1670 551 1671 552
rect 1675 551 1676 555
rect 1670 550 1676 551
rect 1727 555 1733 556
rect 1727 551 1728 555
rect 1732 554 1733 555
rect 1862 555 1863 559
rect 1867 555 1868 559
rect 2479 559 2485 560
rect 2479 558 2480 559
rect 1862 554 1868 555
rect 1872 556 1905 558
rect 2441 556 2480 558
rect 1732 552 1818 554
rect 1732 551 1733 552
rect 1727 550 1733 551
rect 1816 550 1818 552
rect 1872 550 1874 556
rect 2479 555 2480 556
rect 2484 555 2485 559
rect 2479 554 2485 555
rect 3574 559 3580 560
rect 3574 555 3575 559
rect 3579 555 3580 559
rect 3574 554 3580 555
rect 1816 548 1874 550
rect 1886 549 1892 550
rect 150 545 156 546
rect 150 541 151 545
rect 155 541 156 545
rect 150 540 156 541
rect 310 545 316 546
rect 310 541 311 545
rect 315 541 316 545
rect 310 540 316 541
rect 470 545 476 546
rect 470 541 471 545
rect 475 541 476 545
rect 470 540 476 541
rect 630 545 636 546
rect 630 541 631 545
rect 635 541 636 545
rect 630 540 636 541
rect 782 545 788 546
rect 782 541 783 545
rect 787 541 788 545
rect 782 540 788 541
rect 926 545 932 546
rect 926 541 927 545
rect 931 541 932 545
rect 926 540 932 541
rect 1062 545 1068 546
rect 1062 541 1063 545
rect 1067 541 1068 545
rect 1062 540 1068 541
rect 1190 545 1196 546
rect 1190 541 1191 545
rect 1195 541 1196 545
rect 1190 540 1196 541
rect 1310 545 1316 546
rect 1310 541 1311 545
rect 1315 541 1316 545
rect 1310 540 1316 541
rect 1422 545 1428 546
rect 1422 541 1423 545
rect 1427 541 1428 545
rect 1422 540 1428 541
rect 1534 545 1540 546
rect 1534 541 1535 545
rect 1539 541 1540 545
rect 1534 540 1540 541
rect 1646 545 1652 546
rect 1646 541 1647 545
rect 1651 541 1652 545
rect 1646 540 1652 541
rect 1734 545 1740 546
rect 1734 541 1735 545
rect 1739 541 1740 545
rect 1886 545 1887 549
rect 1891 545 1892 549
rect 1886 544 1892 545
rect 2038 549 2044 550
rect 2038 545 2039 549
rect 2043 545 2044 549
rect 2038 544 2044 545
rect 2206 549 2212 550
rect 2206 545 2207 549
rect 2211 545 2212 549
rect 2206 544 2212 545
rect 2382 549 2388 550
rect 2382 545 2383 549
rect 2387 545 2388 549
rect 2382 544 2388 545
rect 2574 549 2580 550
rect 2574 545 2575 549
rect 2579 545 2580 549
rect 2574 544 2580 545
rect 2790 549 2796 550
rect 2790 545 2791 549
rect 2795 545 2796 549
rect 2790 544 2796 545
rect 3014 549 3020 550
rect 3014 545 3015 549
rect 3019 545 3020 549
rect 3014 544 3020 545
rect 3246 549 3252 550
rect 3246 545 3247 549
rect 3251 545 3252 549
rect 3246 544 3252 545
rect 3478 549 3484 550
rect 3478 545 3479 549
rect 3483 545 3484 549
rect 3478 544 3484 545
rect 1734 540 1740 541
rect 110 532 116 533
rect 1822 532 1828 533
rect 110 528 111 532
rect 115 528 116 532
rect 231 531 237 532
rect 231 530 232 531
rect 205 528 232 530
rect 110 527 116 528
rect 231 527 232 528
rect 236 527 237 531
rect 551 531 557 532
rect 551 530 552 531
rect 525 528 552 530
rect 231 526 237 527
rect 295 527 301 528
rect 295 523 296 527
rect 300 526 301 527
rect 551 527 552 528
rect 556 527 557 531
rect 703 531 709 532
rect 703 530 704 531
rect 685 528 704 530
rect 551 526 557 527
rect 703 527 704 528
rect 708 527 709 531
rect 986 531 992 532
rect 986 530 987 531
rect 981 528 987 530
rect 703 526 709 527
rect 986 527 987 528
rect 991 527 992 531
rect 1255 531 1261 532
rect 1255 530 1256 531
rect 1245 528 1256 530
rect 986 526 992 527
rect 994 527 1000 528
rect 300 524 329 526
rect 300 523 301 524
rect 295 522 301 523
rect 994 523 995 527
rect 999 526 1000 527
rect 1255 527 1256 528
rect 1260 527 1261 531
rect 1375 531 1381 532
rect 1375 530 1376 531
rect 1365 528 1376 530
rect 1255 526 1261 527
rect 1375 527 1376 528
rect 1380 527 1381 531
rect 1822 528 1823 532
rect 1827 528 1828 532
rect 1375 526 1381 527
rect 1602 527 1608 528
rect 1822 527 1828 528
rect 2054 527 2060 528
rect 999 524 1081 526
rect 999 523 1000 524
rect 994 522 1000 523
rect 1602 523 1603 527
rect 1607 526 1608 527
rect 1607 524 1665 526
rect 1607 523 1608 524
rect 1602 522 1608 523
rect 2054 523 2055 527
rect 2059 526 2060 527
rect 2059 524 2350 526
rect 2059 523 2060 524
rect 2054 522 2060 523
rect 2190 519 2196 520
rect 110 515 116 516
rect 110 511 111 515
rect 115 511 116 515
rect 110 510 116 511
rect 782 515 788 516
rect 782 511 783 515
rect 787 514 788 515
rect 1490 515 1496 516
rect 787 512 793 514
rect 787 511 788 512
rect 782 510 788 511
rect 1490 511 1491 515
rect 1495 514 1496 515
rect 1822 515 1828 516
rect 1495 512 1545 514
rect 1720 512 1745 514
rect 1495 511 1496 512
rect 1490 510 1496 511
rect 142 505 148 506
rect 142 501 143 505
rect 147 501 148 505
rect 142 500 148 501
rect 302 505 308 506
rect 302 501 303 505
rect 307 501 308 505
rect 302 500 308 501
rect 462 505 468 506
rect 462 501 463 505
rect 467 501 468 505
rect 462 500 468 501
rect 622 505 628 506
rect 622 501 623 505
rect 627 501 628 505
rect 622 500 628 501
rect 774 505 780 506
rect 774 501 775 505
rect 779 501 780 505
rect 774 500 780 501
rect 918 505 924 506
rect 918 501 919 505
rect 923 501 924 505
rect 918 500 924 501
rect 1054 505 1060 506
rect 1054 501 1055 505
rect 1059 501 1060 505
rect 1054 500 1060 501
rect 1182 505 1188 506
rect 1182 501 1183 505
rect 1187 501 1188 505
rect 1182 500 1188 501
rect 1302 505 1308 506
rect 1302 501 1303 505
rect 1307 501 1308 505
rect 1302 500 1308 501
rect 1414 505 1420 506
rect 1414 501 1415 505
rect 1419 501 1420 505
rect 1414 500 1420 501
rect 1526 505 1532 506
rect 1526 501 1527 505
rect 1531 501 1532 505
rect 1526 500 1532 501
rect 1638 505 1644 506
rect 1638 501 1639 505
rect 1643 501 1644 505
rect 1638 500 1644 501
rect 1454 499 1460 500
rect 1454 495 1455 499
rect 1459 498 1460 499
rect 1463 499 1469 500
rect 1463 498 1464 499
rect 1459 496 1464 498
rect 1459 495 1460 496
rect 1454 494 1460 495
rect 1463 495 1464 496
rect 1468 495 1469 499
rect 1720 498 1722 512
rect 1822 511 1823 515
rect 1827 511 1828 515
rect 2190 515 2191 519
rect 2195 515 2196 519
rect 2190 514 2196 515
rect 2278 519 2284 520
rect 2278 515 2279 519
rect 2283 515 2284 519
rect 2278 514 2284 515
rect 1822 510 1828 511
rect 2348 510 2350 524
rect 2374 519 2380 520
rect 2374 515 2375 519
rect 2379 515 2380 519
rect 2374 514 2380 515
rect 2486 519 2492 520
rect 2486 515 2487 519
rect 2491 515 2492 519
rect 2486 514 2492 515
rect 2630 519 2636 520
rect 2630 515 2631 519
rect 2635 515 2636 519
rect 2630 514 2636 515
rect 2806 519 2812 520
rect 2806 515 2807 519
rect 2811 515 2812 519
rect 2806 514 2812 515
rect 3006 519 3012 520
rect 3006 515 3007 519
rect 3011 515 3012 519
rect 3006 514 3012 515
rect 3214 519 3220 520
rect 3214 515 3215 519
rect 3219 515 3220 519
rect 3214 514 3220 515
rect 3430 519 3436 520
rect 3430 515 3431 519
rect 3435 515 3436 519
rect 3430 514 3436 515
rect 1862 509 1868 510
rect 1726 505 1732 506
rect 1726 501 1727 505
rect 1731 501 1732 505
rect 1862 505 1863 509
rect 1867 505 1868 509
rect 2348 508 2393 510
rect 3574 509 3580 510
rect 1862 504 1868 505
rect 3574 505 3575 509
rect 3579 505 3580 509
rect 3574 504 3580 505
rect 1726 500 1732 501
rect 1463 494 1469 495
rect 1696 496 1722 498
rect 1670 491 1676 492
rect 1670 487 1671 491
rect 1675 490 1676 491
rect 1696 490 1698 496
rect 2271 495 2277 496
rect 2271 494 2272 495
rect 1675 488 1698 490
rect 1862 492 1868 493
rect 2253 492 2272 494
rect 1862 488 1863 492
rect 1867 488 1868 492
rect 2271 491 2272 492
rect 2276 491 2277 495
rect 2346 495 2352 496
rect 2346 494 2347 495
rect 2341 492 2347 494
rect 2271 490 2277 491
rect 2346 491 2347 492
rect 2351 491 2352 495
rect 2623 495 2629 496
rect 2623 494 2624 495
rect 2549 492 2624 494
rect 2346 490 2352 491
rect 2623 491 2624 492
rect 2628 491 2629 495
rect 2799 495 2805 496
rect 2799 494 2800 495
rect 2693 492 2800 494
rect 2623 490 2629 491
rect 2799 491 2800 492
rect 2804 491 2805 495
rect 2983 495 2989 496
rect 2983 494 2984 495
rect 2869 492 2984 494
rect 2799 490 2805 491
rect 2983 491 2984 492
rect 2988 491 2989 495
rect 3175 495 3181 496
rect 3175 494 3176 495
rect 3069 492 3176 494
rect 2983 490 2989 491
rect 3175 491 3176 492
rect 3180 491 3181 495
rect 3175 490 3181 491
rect 3186 495 3192 496
rect 3186 491 3187 495
rect 3191 494 3192 495
rect 3498 495 3504 496
rect 3498 494 3499 495
rect 3191 492 3241 494
rect 3493 492 3499 494
rect 3191 491 3192 492
rect 3186 490 3192 491
rect 3498 491 3499 492
rect 3503 491 3504 495
rect 3498 490 3504 491
rect 3574 492 3580 493
rect 1675 487 1676 488
rect 1862 487 1868 488
rect 3574 488 3575 492
rect 3579 488 3580 492
rect 3574 487 3580 488
rect 1670 486 1676 487
rect 2198 479 2204 480
rect 158 475 164 476
rect 158 471 159 475
rect 163 471 164 475
rect 158 470 164 471
rect 310 475 316 476
rect 310 471 311 475
rect 315 471 316 475
rect 310 470 316 471
rect 462 475 468 476
rect 462 471 463 475
rect 467 471 468 475
rect 462 470 468 471
rect 614 475 620 476
rect 614 471 615 475
rect 619 471 620 475
rect 614 470 620 471
rect 758 475 764 476
rect 758 471 759 475
rect 763 471 764 475
rect 758 470 764 471
rect 886 475 892 476
rect 886 471 887 475
rect 891 471 892 475
rect 886 470 892 471
rect 1006 475 1012 476
rect 1006 471 1007 475
rect 1011 471 1012 475
rect 1006 470 1012 471
rect 1126 475 1132 476
rect 1126 471 1127 475
rect 1131 471 1132 475
rect 1126 470 1132 471
rect 1238 475 1244 476
rect 1238 471 1239 475
rect 1243 471 1244 475
rect 1238 470 1244 471
rect 1342 475 1348 476
rect 1342 471 1343 475
rect 1347 471 1348 475
rect 1342 470 1348 471
rect 1438 475 1444 476
rect 1438 471 1439 475
rect 1443 471 1444 475
rect 1438 470 1444 471
rect 1542 475 1548 476
rect 1542 471 1543 475
rect 1547 471 1548 475
rect 1542 470 1548 471
rect 1638 475 1644 476
rect 1638 471 1639 475
rect 1643 471 1644 475
rect 1638 470 1644 471
rect 1726 475 1732 476
rect 1726 471 1727 475
rect 1731 471 1732 475
rect 2198 475 2199 479
rect 2203 475 2204 479
rect 2198 474 2204 475
rect 2286 479 2292 480
rect 2286 475 2287 479
rect 2291 475 2292 479
rect 2286 474 2292 475
rect 2382 479 2388 480
rect 2382 475 2383 479
rect 2387 475 2388 479
rect 2382 474 2388 475
rect 2494 479 2500 480
rect 2494 475 2495 479
rect 2499 475 2500 479
rect 2494 474 2500 475
rect 2638 479 2644 480
rect 2638 475 2639 479
rect 2643 475 2644 479
rect 2638 474 2644 475
rect 2814 479 2820 480
rect 2814 475 2815 479
rect 2819 475 2820 479
rect 2814 474 2820 475
rect 3014 479 3020 480
rect 3014 475 3015 479
rect 3019 475 3020 479
rect 3014 474 3020 475
rect 3222 479 3228 480
rect 3222 475 3223 479
rect 3227 475 3228 479
rect 3222 474 3228 475
rect 3438 479 3444 480
rect 3438 475 3439 479
rect 3443 475 3444 479
rect 3438 474 3444 475
rect 1726 470 1732 471
rect 135 467 141 468
rect 110 465 116 466
rect 110 461 111 465
rect 115 461 116 465
rect 135 463 136 467
rect 140 466 141 467
rect 1074 467 1080 468
rect 1074 466 1075 467
rect 140 464 177 466
rect 1065 464 1075 466
rect 140 463 141 464
rect 135 462 141 463
rect 1074 463 1075 464
rect 1079 463 1080 467
rect 2119 467 2125 468
rect 1074 462 1080 463
rect 1822 465 1828 466
rect 110 460 116 461
rect 1822 461 1823 465
rect 1827 461 1828 465
rect 2119 463 2120 467
rect 2124 466 2125 467
rect 2191 467 2197 468
rect 2191 466 2192 467
rect 2124 464 2192 466
rect 2124 463 2125 464
rect 2119 462 2125 463
rect 2191 463 2192 464
rect 2196 463 2197 467
rect 2191 462 2197 463
rect 2271 467 2277 468
rect 2271 463 2272 467
rect 2276 466 2277 467
rect 2279 467 2285 468
rect 2279 466 2280 467
rect 2276 464 2280 466
rect 2276 463 2277 464
rect 2271 462 2277 463
rect 2279 463 2280 464
rect 2284 463 2285 467
rect 2279 462 2285 463
rect 2346 467 2352 468
rect 2346 463 2347 467
rect 2351 466 2352 467
rect 2375 467 2381 468
rect 2375 466 2376 467
rect 2351 464 2376 466
rect 2351 463 2352 464
rect 2346 462 2352 463
rect 2375 463 2376 464
rect 2380 463 2381 467
rect 2375 462 2381 463
rect 2479 467 2485 468
rect 2479 463 2480 467
rect 2484 466 2485 467
rect 2487 467 2493 468
rect 2487 466 2488 467
rect 2484 464 2488 466
rect 2484 463 2485 464
rect 2479 462 2485 463
rect 2487 463 2488 464
rect 2492 463 2493 467
rect 2487 462 2493 463
rect 2623 467 2629 468
rect 2623 463 2624 467
rect 2628 466 2629 467
rect 2631 467 2637 468
rect 2631 466 2632 467
rect 2628 464 2632 466
rect 2628 463 2629 464
rect 2623 462 2629 463
rect 2631 463 2632 464
rect 2636 463 2637 467
rect 2631 462 2637 463
rect 2799 467 2805 468
rect 2799 463 2800 467
rect 2804 466 2805 467
rect 2807 467 2813 468
rect 2807 466 2808 467
rect 2804 464 2808 466
rect 2804 463 2805 464
rect 2799 462 2805 463
rect 2807 463 2808 464
rect 2812 463 2813 467
rect 2807 462 2813 463
rect 2983 467 2989 468
rect 2983 463 2984 467
rect 2988 466 2989 467
rect 3007 467 3013 468
rect 3007 466 3008 467
rect 2988 464 3008 466
rect 2988 463 2989 464
rect 2983 462 2989 463
rect 3007 463 3008 464
rect 3012 463 3013 467
rect 3007 462 3013 463
rect 3175 467 3181 468
rect 3175 463 3176 467
rect 3180 466 3181 467
rect 3215 467 3221 468
rect 3215 466 3216 467
rect 3180 464 3216 466
rect 3180 463 3181 464
rect 3175 462 3181 463
rect 3215 463 3216 464
rect 3220 463 3221 467
rect 3215 462 3221 463
rect 3423 467 3429 468
rect 3423 463 3424 467
rect 3428 466 3429 467
rect 3431 467 3437 468
rect 3431 466 3432 467
rect 3428 464 3432 466
rect 3428 463 3429 464
rect 3423 462 3429 463
rect 3431 463 3432 464
rect 3436 463 3437 467
rect 3431 462 3437 463
rect 1822 460 1828 461
rect 1816 452 1834 454
rect 247 451 253 452
rect 110 448 116 449
rect 110 444 111 448
rect 115 444 116 448
rect 247 447 248 451
rect 252 450 253 451
rect 542 451 548 452
rect 542 450 543 451
rect 252 448 337 450
rect 525 448 543 450
rect 252 447 253 448
rect 247 446 253 447
rect 542 447 543 448
rect 547 447 548 451
rect 542 446 548 447
rect 551 451 557 452
rect 551 447 552 451
rect 556 450 557 451
rect 698 451 704 452
rect 556 448 641 450
rect 556 447 557 448
rect 551 446 557 447
rect 698 447 699 451
rect 703 450 704 451
rect 999 451 1005 452
rect 999 450 1000 451
rect 703 448 785 450
rect 949 448 1000 450
rect 703 447 704 448
rect 698 446 704 447
rect 999 447 1000 448
rect 1004 447 1005 451
rect 1231 451 1237 452
rect 1231 450 1232 451
rect 1189 448 1232 450
rect 999 446 1005 447
rect 1231 447 1232 448
rect 1236 447 1237 451
rect 1335 451 1341 452
rect 1335 450 1336 451
rect 1301 448 1336 450
rect 1231 446 1237 447
rect 1335 447 1336 448
rect 1340 447 1341 451
rect 1430 451 1436 452
rect 1430 450 1431 451
rect 1405 448 1431 450
rect 1335 446 1341 447
rect 1430 447 1431 448
rect 1435 447 1436 451
rect 1535 451 1541 452
rect 1535 450 1536 451
rect 1501 448 1536 450
rect 1430 446 1436 447
rect 1535 447 1536 448
rect 1540 447 1541 451
rect 1631 451 1637 452
rect 1631 450 1632 451
rect 1605 448 1632 450
rect 1535 446 1541 447
rect 1631 447 1632 448
rect 1636 447 1637 451
rect 1711 451 1717 452
rect 1711 450 1712 451
rect 1701 448 1712 450
rect 1631 446 1637 447
rect 1711 447 1712 448
rect 1716 447 1717 451
rect 1816 450 1818 452
rect 1789 448 1818 450
rect 1822 448 1828 449
rect 1711 446 1717 447
rect 110 443 116 444
rect 1822 444 1823 448
rect 1827 444 1828 448
rect 1832 446 1834 452
rect 1887 447 1893 448
rect 1887 446 1888 447
rect 1832 444 1888 446
rect 1822 443 1828 444
rect 1887 443 1888 444
rect 1892 443 1893 447
rect 1887 442 1893 443
rect 2031 447 2037 448
rect 2031 443 2032 447
rect 2036 446 2037 447
rect 2127 447 2133 448
rect 2127 446 2128 447
rect 2036 444 2128 446
rect 2036 443 2037 444
rect 2031 442 2037 443
rect 2127 443 2128 444
rect 2132 443 2133 447
rect 2127 442 2133 443
rect 2199 447 2205 448
rect 2199 443 2200 447
rect 2204 446 2205 447
rect 2218 447 2224 448
rect 2218 446 2219 447
rect 2204 444 2219 446
rect 2204 443 2205 444
rect 2199 442 2205 443
rect 2218 443 2219 444
rect 2223 443 2224 447
rect 2218 442 2224 443
rect 2375 447 2381 448
rect 2375 443 2376 447
rect 2380 446 2381 447
rect 2390 447 2396 448
rect 2390 446 2391 447
rect 2380 444 2391 446
rect 2380 443 2381 444
rect 2375 442 2381 443
rect 2390 443 2391 444
rect 2395 443 2396 447
rect 2390 442 2396 443
rect 2479 447 2485 448
rect 2479 443 2480 447
rect 2484 446 2485 447
rect 2567 447 2573 448
rect 2567 446 2568 447
rect 2484 444 2568 446
rect 2484 443 2485 444
rect 2479 442 2485 443
rect 2567 443 2568 444
rect 2572 443 2573 447
rect 2567 442 2573 443
rect 2679 447 2685 448
rect 2679 443 2680 447
rect 2684 446 2685 447
rect 2775 447 2781 448
rect 2775 446 2776 447
rect 2684 444 2776 446
rect 2684 443 2685 444
rect 2679 442 2685 443
rect 2775 443 2776 444
rect 2780 443 2781 447
rect 2775 442 2781 443
rect 2895 447 2901 448
rect 2895 443 2896 447
rect 2900 446 2901 447
rect 2999 447 3005 448
rect 2999 446 3000 447
rect 2900 444 3000 446
rect 2900 443 2901 444
rect 2895 442 2901 443
rect 2999 443 3000 444
rect 3004 443 3005 447
rect 2999 442 3005 443
rect 3079 447 3085 448
rect 3079 443 3080 447
rect 3084 446 3085 447
rect 3231 447 3237 448
rect 3231 446 3232 447
rect 3084 444 3232 446
rect 3084 443 3085 444
rect 3079 442 3085 443
rect 3231 443 3232 444
rect 3236 443 3237 447
rect 3231 442 3237 443
rect 3463 447 3469 448
rect 3463 443 3464 447
rect 3468 446 3469 447
rect 3498 447 3504 448
rect 3498 446 3499 447
rect 3468 444 3499 446
rect 3468 443 3469 444
rect 3463 442 3469 443
rect 3498 443 3499 444
rect 3503 443 3504 447
rect 3498 442 3504 443
rect 1894 437 1900 438
rect 166 435 172 436
rect 166 431 167 435
rect 171 431 172 435
rect 166 430 172 431
rect 318 435 324 436
rect 318 431 319 435
rect 323 431 324 435
rect 318 430 324 431
rect 470 435 476 436
rect 470 431 471 435
rect 475 431 476 435
rect 470 430 476 431
rect 622 435 628 436
rect 622 431 623 435
rect 627 431 628 435
rect 622 430 628 431
rect 766 435 772 436
rect 766 431 767 435
rect 771 431 772 435
rect 766 430 772 431
rect 894 435 900 436
rect 894 431 895 435
rect 899 431 900 435
rect 894 430 900 431
rect 1014 435 1020 436
rect 1014 431 1015 435
rect 1019 431 1020 435
rect 1014 430 1020 431
rect 1134 435 1140 436
rect 1134 431 1135 435
rect 1139 431 1140 435
rect 1134 430 1140 431
rect 1246 435 1252 436
rect 1246 431 1247 435
rect 1251 431 1252 435
rect 1246 430 1252 431
rect 1350 435 1356 436
rect 1350 431 1351 435
rect 1355 431 1356 435
rect 1350 430 1356 431
rect 1446 435 1452 436
rect 1446 431 1447 435
rect 1451 431 1452 435
rect 1446 430 1452 431
rect 1550 435 1556 436
rect 1550 431 1551 435
rect 1555 431 1556 435
rect 1550 430 1556 431
rect 1646 435 1652 436
rect 1646 431 1647 435
rect 1651 431 1652 435
rect 1646 430 1652 431
rect 1734 435 1740 436
rect 1734 431 1735 435
rect 1739 431 1740 435
rect 1894 433 1895 437
rect 1899 433 1900 437
rect 1894 432 1900 433
rect 2038 437 2044 438
rect 2038 433 2039 437
rect 2043 433 2044 437
rect 2038 432 2044 433
rect 2206 437 2212 438
rect 2206 433 2207 437
rect 2211 433 2212 437
rect 2206 432 2212 433
rect 2382 437 2388 438
rect 2382 433 2383 437
rect 2387 433 2388 437
rect 2382 432 2388 433
rect 2574 437 2580 438
rect 2574 433 2575 437
rect 2579 433 2580 437
rect 2574 432 2580 433
rect 2782 437 2788 438
rect 2782 433 2783 437
rect 2787 433 2788 437
rect 2782 432 2788 433
rect 3006 437 3012 438
rect 3006 433 3007 437
rect 3011 433 3012 437
rect 3006 432 3012 433
rect 3238 437 3244 438
rect 3238 433 3239 437
rect 3243 433 3244 437
rect 3238 432 3244 433
rect 3470 437 3476 438
rect 3470 433 3471 437
rect 3475 433 3476 437
rect 3470 432 3476 433
rect 1734 430 1740 431
rect 1862 424 1868 425
rect 3574 424 3580 425
rect 159 423 165 424
rect 159 419 160 423
rect 164 422 165 423
rect 247 423 253 424
rect 247 422 248 423
rect 164 420 248 422
rect 164 419 165 420
rect 159 418 165 419
rect 247 419 248 420
rect 252 419 253 423
rect 247 418 253 419
rect 311 423 317 424
rect 311 419 312 423
rect 316 422 317 423
rect 330 423 336 424
rect 330 422 331 423
rect 316 420 331 422
rect 316 419 317 420
rect 311 418 317 419
rect 330 419 331 420
rect 335 419 336 423
rect 330 418 336 419
rect 463 423 469 424
rect 463 419 464 423
rect 468 422 469 423
rect 551 423 557 424
rect 551 422 552 423
rect 468 420 552 422
rect 468 419 469 420
rect 463 418 469 419
rect 551 419 552 420
rect 556 419 557 423
rect 551 418 557 419
rect 615 423 621 424
rect 615 419 616 423
rect 620 422 621 423
rect 698 423 704 424
rect 698 422 699 423
rect 620 420 699 422
rect 620 419 621 420
rect 615 418 621 419
rect 698 419 699 420
rect 703 419 704 423
rect 698 418 704 419
rect 759 423 765 424
rect 759 419 760 423
rect 764 422 765 423
rect 782 423 788 424
rect 782 422 783 423
rect 764 420 783 422
rect 764 419 765 420
rect 759 418 765 419
rect 782 419 783 420
rect 787 419 788 423
rect 782 418 788 419
rect 887 423 893 424
rect 887 419 888 423
rect 892 422 893 423
rect 902 423 908 424
rect 902 422 903 423
rect 892 420 903 422
rect 892 419 893 420
rect 887 418 893 419
rect 902 419 903 420
rect 907 419 908 423
rect 902 418 908 419
rect 999 423 1005 424
rect 999 419 1000 423
rect 1004 422 1005 423
rect 1007 423 1013 424
rect 1007 422 1008 423
rect 1004 420 1008 422
rect 1004 419 1005 420
rect 999 418 1005 419
rect 1007 419 1008 420
rect 1012 419 1013 423
rect 1007 418 1013 419
rect 1127 423 1133 424
rect 1127 419 1128 423
rect 1132 422 1133 423
rect 1142 423 1148 424
rect 1142 422 1143 423
rect 1132 420 1143 422
rect 1132 419 1133 420
rect 1127 418 1133 419
rect 1142 419 1143 420
rect 1147 419 1148 423
rect 1142 418 1148 419
rect 1231 423 1237 424
rect 1231 419 1232 423
rect 1236 422 1237 423
rect 1239 423 1245 424
rect 1239 422 1240 423
rect 1236 420 1240 422
rect 1236 419 1237 420
rect 1231 418 1237 419
rect 1239 419 1240 420
rect 1244 419 1245 423
rect 1239 418 1245 419
rect 1335 423 1341 424
rect 1335 419 1336 423
rect 1340 422 1341 423
rect 1343 423 1349 424
rect 1343 422 1344 423
rect 1340 420 1344 422
rect 1340 419 1341 420
rect 1335 418 1341 419
rect 1343 419 1344 420
rect 1348 419 1349 423
rect 1343 418 1349 419
rect 1439 423 1445 424
rect 1439 419 1440 423
rect 1444 422 1445 423
rect 1454 423 1460 424
rect 1454 422 1455 423
rect 1444 420 1455 422
rect 1444 419 1445 420
rect 1439 418 1445 419
rect 1454 419 1455 420
rect 1459 419 1460 423
rect 1454 418 1460 419
rect 1535 423 1541 424
rect 1535 419 1536 423
rect 1540 422 1541 423
rect 1543 423 1549 424
rect 1543 422 1544 423
rect 1540 420 1544 422
rect 1540 419 1541 420
rect 1535 418 1541 419
rect 1543 419 1544 420
rect 1548 419 1549 423
rect 1543 418 1549 419
rect 1631 423 1637 424
rect 1631 419 1632 423
rect 1636 422 1637 423
rect 1639 423 1645 424
rect 1639 422 1640 423
rect 1636 420 1640 422
rect 1636 419 1637 420
rect 1631 418 1637 419
rect 1639 419 1640 420
rect 1644 419 1645 423
rect 1639 418 1645 419
rect 1711 423 1717 424
rect 1711 419 1712 423
rect 1716 422 1717 423
rect 1727 423 1733 424
rect 1727 422 1728 423
rect 1716 420 1728 422
rect 1716 419 1717 420
rect 1711 418 1717 419
rect 1727 419 1728 420
rect 1732 419 1733 423
rect 1862 420 1863 424
rect 1867 420 1868 424
rect 2119 423 2125 424
rect 2119 422 2120 423
rect 2093 420 2120 422
rect 1862 419 1868 420
rect 2119 419 2120 420
rect 2124 419 2125 423
rect 2479 423 2485 424
rect 2479 422 2480 423
rect 2437 420 2480 422
rect 1727 418 1733 419
rect 2119 418 2125 419
rect 2127 419 2133 420
rect 2127 415 2128 419
rect 2132 418 2133 419
rect 2479 419 2480 420
rect 2484 419 2485 423
rect 2679 423 2685 424
rect 2679 422 2680 423
rect 2629 420 2680 422
rect 2479 418 2485 419
rect 2679 419 2680 420
rect 2684 419 2685 423
rect 2895 423 2901 424
rect 2895 422 2896 423
rect 2837 420 2896 422
rect 2679 418 2685 419
rect 2895 419 2896 420
rect 2900 419 2901 423
rect 3079 423 3085 424
rect 3079 422 3080 423
rect 3061 420 3080 422
rect 2895 418 2901 419
rect 3079 419 3080 420
rect 3084 419 3085 423
rect 3574 420 3575 424
rect 3579 420 3580 424
rect 3574 419 3580 420
rect 3079 418 3085 419
rect 2132 416 2225 418
rect 2132 415 2133 416
rect 2127 414 2133 415
rect 143 411 149 412
rect 143 407 144 411
rect 148 410 149 411
rect 158 411 164 412
rect 158 410 159 411
rect 148 408 159 410
rect 148 407 149 408
rect 143 406 149 407
rect 158 407 159 408
rect 163 407 164 411
rect 158 406 164 407
rect 215 411 221 412
rect 215 407 216 411
rect 220 410 221 411
rect 263 411 269 412
rect 263 410 264 411
rect 220 408 264 410
rect 220 407 221 408
rect 215 406 221 407
rect 263 407 264 408
rect 268 407 269 411
rect 263 406 269 407
rect 391 411 397 412
rect 391 407 392 411
rect 396 410 397 411
rect 399 411 405 412
rect 399 410 400 411
rect 396 408 400 410
rect 396 407 397 408
rect 391 406 397 407
rect 399 407 400 408
rect 404 407 405 411
rect 399 406 405 407
rect 542 411 549 412
rect 542 407 543 411
rect 548 407 549 411
rect 542 406 549 407
rect 646 411 652 412
rect 646 407 647 411
rect 651 410 652 411
rect 703 411 709 412
rect 703 410 704 411
rect 651 408 704 410
rect 651 407 652 408
rect 646 406 652 407
rect 703 407 704 408
rect 708 407 709 411
rect 703 406 709 407
rect 799 411 805 412
rect 799 407 800 411
rect 804 410 805 411
rect 879 411 885 412
rect 879 410 880 411
rect 804 408 880 410
rect 804 407 805 408
rect 799 406 805 407
rect 879 407 880 408
rect 884 407 885 411
rect 879 406 885 407
rect 1055 411 1061 412
rect 1055 407 1056 411
rect 1060 410 1061 411
rect 1082 411 1088 412
rect 1082 410 1083 411
rect 1060 408 1083 410
rect 1060 407 1061 408
rect 1055 406 1061 407
rect 1082 407 1083 408
rect 1087 407 1088 411
rect 1082 406 1088 407
rect 1151 411 1157 412
rect 1151 407 1152 411
rect 1156 410 1157 411
rect 1239 411 1245 412
rect 1239 410 1240 411
rect 1156 408 1240 410
rect 1156 407 1157 408
rect 1151 406 1157 407
rect 1239 407 1240 408
rect 1244 407 1245 411
rect 1239 406 1245 407
rect 1430 411 1437 412
rect 1430 407 1431 411
rect 1436 407 1437 411
rect 1430 406 1437 407
rect 1535 411 1541 412
rect 1535 407 1536 411
rect 1540 410 1541 411
rect 1631 411 1637 412
rect 1631 410 1632 411
rect 1540 408 1632 410
rect 1540 407 1541 408
rect 1535 406 1541 407
rect 1631 407 1632 408
rect 1636 407 1637 411
rect 1631 406 1637 407
rect 1862 407 1868 408
rect 1862 403 1863 407
rect 1867 403 1868 407
rect 1862 402 1868 403
rect 1879 407 1885 408
rect 1879 403 1880 407
rect 1884 406 1885 407
rect 3178 407 3184 408
rect 1884 404 1905 406
rect 1884 403 1885 404
rect 1879 402 1885 403
rect 3178 403 3179 407
rect 3183 406 3184 407
rect 3470 407 3476 408
rect 3183 404 3249 406
rect 3183 403 3184 404
rect 3178 402 3184 403
rect 3470 403 3471 407
rect 3475 406 3476 407
rect 3574 407 3580 408
rect 3475 404 3481 406
rect 3475 403 3476 404
rect 3470 402 3476 403
rect 3574 403 3575 407
rect 3579 403 3580 407
rect 3574 402 3580 403
rect 150 401 156 402
rect 150 397 151 401
rect 155 397 156 401
rect 150 396 156 397
rect 270 401 276 402
rect 270 397 271 401
rect 275 397 276 401
rect 270 396 276 397
rect 406 401 412 402
rect 406 397 407 401
rect 411 397 412 401
rect 406 396 412 397
rect 550 401 556 402
rect 550 397 551 401
rect 555 397 556 401
rect 550 396 556 397
rect 710 401 716 402
rect 710 397 711 401
rect 715 397 716 401
rect 710 396 716 397
rect 886 401 892 402
rect 886 397 887 401
rect 891 397 892 401
rect 886 396 892 397
rect 1062 401 1068 402
rect 1062 397 1063 401
rect 1067 397 1068 401
rect 1062 396 1068 397
rect 1246 401 1252 402
rect 1246 397 1247 401
rect 1251 397 1252 401
rect 1246 396 1252 397
rect 1438 401 1444 402
rect 1438 397 1439 401
rect 1443 397 1444 401
rect 1438 396 1444 397
rect 1638 401 1644 402
rect 1638 397 1639 401
rect 1643 397 1644 401
rect 1638 396 1644 397
rect 1886 397 1892 398
rect 1886 393 1887 397
rect 1891 393 1892 397
rect 1886 392 1892 393
rect 2030 397 2036 398
rect 2030 393 2031 397
rect 2035 393 2036 397
rect 2030 392 2036 393
rect 2198 397 2204 398
rect 2198 393 2199 397
rect 2203 393 2204 397
rect 2198 392 2204 393
rect 2374 397 2380 398
rect 2374 393 2375 397
rect 2379 393 2380 397
rect 2374 392 2380 393
rect 2566 397 2572 398
rect 2566 393 2567 397
rect 2571 393 2572 397
rect 2566 392 2572 393
rect 2774 397 2780 398
rect 2774 393 2775 397
rect 2779 393 2780 397
rect 2774 392 2780 393
rect 2998 397 3004 398
rect 2998 393 2999 397
rect 3003 393 3004 397
rect 2998 392 3004 393
rect 3230 397 3236 398
rect 3230 393 3231 397
rect 3235 393 3236 397
rect 3230 392 3236 393
rect 3462 397 3468 398
rect 3462 393 3463 397
rect 3467 393 3468 397
rect 3462 392 3468 393
rect 110 388 116 389
rect 1822 388 1828 389
rect 110 384 111 388
rect 115 384 116 388
rect 215 387 221 388
rect 215 386 216 387
rect 205 384 216 386
rect 110 383 116 384
rect 215 383 216 384
rect 220 383 221 387
rect 330 387 336 388
rect 330 386 331 387
rect 325 384 331 386
rect 215 382 221 383
rect 330 383 331 384
rect 335 383 336 387
rect 646 387 652 388
rect 646 386 647 387
rect 605 384 647 386
rect 330 382 336 383
rect 338 383 344 384
rect 338 379 339 383
rect 343 382 344 383
rect 646 383 647 384
rect 651 383 652 387
rect 799 387 805 388
rect 799 386 800 387
rect 765 384 800 386
rect 646 382 652 383
rect 799 383 800 384
rect 804 383 805 387
rect 1151 387 1157 388
rect 1151 386 1152 387
rect 1117 384 1152 386
rect 799 382 805 383
rect 1151 383 1152 384
rect 1156 383 1157 387
rect 1535 387 1541 388
rect 1535 386 1536 387
rect 1493 384 1536 386
rect 1151 382 1157 383
rect 1162 383 1168 384
rect 343 380 425 382
rect 343 379 344 380
rect 338 378 344 379
rect 1162 379 1163 383
rect 1167 382 1168 383
rect 1535 383 1536 384
rect 1540 383 1541 387
rect 1822 384 1823 388
rect 1827 384 1828 388
rect 1822 383 1828 384
rect 1902 383 1908 384
rect 1535 382 1541 383
rect 1167 380 1265 382
rect 1167 379 1168 380
rect 1162 378 1168 379
rect 1902 379 1903 383
rect 1907 382 1908 383
rect 1907 380 2134 382
rect 1907 379 1908 380
rect 1902 378 1908 379
rect 1886 375 1892 376
rect 110 371 116 372
rect 110 367 111 371
rect 115 367 116 371
rect 110 366 116 367
rect 854 371 860 372
rect 854 367 855 371
rect 859 370 860 371
rect 1822 371 1828 372
rect 859 368 897 370
rect 859 367 860 368
rect 854 366 860 367
rect 1822 367 1823 371
rect 1827 367 1828 371
rect 1886 371 1887 375
rect 1891 371 1892 375
rect 1886 370 1892 371
rect 1974 375 1980 376
rect 1974 371 1975 375
rect 1979 371 1980 375
rect 1974 370 1980 371
rect 2062 375 2068 376
rect 2062 371 2063 375
rect 2067 371 2068 375
rect 2062 370 2068 371
rect 1822 366 1828 367
rect 2132 366 2134 380
rect 2150 375 2156 376
rect 2150 371 2151 375
rect 2155 371 2156 375
rect 2150 370 2156 371
rect 2262 375 2268 376
rect 2262 371 2263 375
rect 2267 371 2268 375
rect 2262 370 2268 371
rect 2382 375 2388 376
rect 2382 371 2383 375
rect 2387 371 2388 375
rect 2382 370 2388 371
rect 2518 375 2524 376
rect 2518 371 2519 375
rect 2523 371 2524 375
rect 2518 370 2524 371
rect 2670 375 2676 376
rect 2670 371 2671 375
rect 2675 371 2676 375
rect 2670 370 2676 371
rect 2846 375 2852 376
rect 2846 371 2847 375
rect 2851 371 2852 375
rect 2846 370 2852 371
rect 3030 375 3036 376
rect 3030 371 3031 375
rect 3035 371 3036 375
rect 3030 370 3036 371
rect 3230 375 3236 376
rect 3230 371 3231 375
rect 3235 371 3236 375
rect 3230 370 3236 371
rect 3430 375 3436 376
rect 3430 371 3431 375
rect 3435 371 3436 375
rect 3430 370 3436 371
rect 2218 367 2224 368
rect 1862 365 1868 366
rect 142 361 148 362
rect 142 357 143 361
rect 147 357 148 361
rect 142 356 148 357
rect 262 361 268 362
rect 262 357 263 361
rect 267 357 268 361
rect 262 356 268 357
rect 398 361 404 362
rect 398 357 399 361
rect 403 357 404 361
rect 398 356 404 357
rect 542 361 548 362
rect 542 357 543 361
rect 547 357 548 361
rect 542 356 548 357
rect 702 361 708 362
rect 702 357 703 361
rect 707 357 708 361
rect 702 356 708 357
rect 878 361 884 362
rect 878 357 879 361
rect 883 357 884 361
rect 878 356 884 357
rect 1054 361 1060 362
rect 1054 357 1055 361
rect 1059 357 1060 361
rect 1054 356 1060 357
rect 1238 361 1244 362
rect 1238 357 1239 361
rect 1243 357 1244 361
rect 1238 356 1244 357
rect 1430 361 1436 362
rect 1430 357 1431 361
rect 1435 357 1436 361
rect 1430 356 1436 357
rect 1630 361 1636 362
rect 1630 357 1631 361
rect 1635 357 1636 361
rect 1862 361 1863 365
rect 1867 361 1868 365
rect 2132 364 2169 366
rect 2218 363 2219 367
rect 2223 366 2224 367
rect 3423 367 3429 368
rect 2223 364 2281 366
rect 2223 363 2224 364
rect 2218 362 2224 363
rect 3423 363 3424 367
rect 3428 366 3429 367
rect 3428 364 3449 366
rect 3574 365 3580 366
rect 3428 363 3429 364
rect 3423 362 3429 363
rect 1862 360 1868 361
rect 3574 361 3575 365
rect 3579 361 3580 365
rect 3574 360 3580 361
rect 1630 356 1636 357
rect 1663 355 1669 356
rect 1663 351 1664 355
rect 1668 354 1669 355
rect 1679 355 1685 356
rect 1679 354 1680 355
rect 1668 352 1680 354
rect 1668 351 1669 352
rect 1663 350 1669 351
rect 1679 351 1680 352
rect 1684 351 1685 355
rect 1679 350 1685 351
rect 1967 351 1973 352
rect 1967 350 1968 351
rect 1862 348 1868 349
rect 1949 348 1968 350
rect 1862 344 1863 348
rect 1867 344 1868 348
rect 1967 347 1968 348
rect 1972 347 1973 351
rect 2055 351 2061 352
rect 2055 350 2056 351
rect 2037 348 2056 350
rect 1967 346 1973 347
rect 2055 347 2056 348
rect 2060 347 2061 351
rect 2143 351 2149 352
rect 2143 350 2144 351
rect 2125 348 2144 350
rect 2055 346 2061 347
rect 2143 347 2144 348
rect 2148 347 2149 351
rect 2143 346 2149 347
rect 2351 351 2357 352
rect 2351 347 2352 351
rect 2356 350 2357 351
rect 2450 351 2456 352
rect 2356 348 2409 350
rect 2356 347 2357 348
rect 2351 346 2357 347
rect 2450 347 2451 351
rect 2455 350 2456 351
rect 2839 351 2845 352
rect 2839 350 2840 351
rect 2455 348 2545 350
rect 2733 348 2840 350
rect 2455 347 2456 348
rect 2450 346 2456 347
rect 2839 347 2840 348
rect 2844 347 2845 351
rect 3023 351 3029 352
rect 3023 350 3024 351
rect 2909 348 3024 350
rect 2839 346 2845 347
rect 3023 347 3024 348
rect 3028 347 3029 351
rect 3150 351 3156 352
rect 3150 350 3151 351
rect 3093 348 3151 350
rect 3023 346 3029 347
rect 3150 347 3151 348
rect 3155 347 3156 351
rect 3150 346 3156 347
rect 3158 351 3164 352
rect 3158 347 3159 351
rect 3163 350 3164 351
rect 3163 348 3257 350
rect 3574 348 3580 349
rect 3163 347 3164 348
rect 3158 346 3164 347
rect 1862 343 1868 344
rect 3574 344 3575 348
rect 3579 344 3580 348
rect 3574 343 3580 344
rect 1894 335 1900 336
rect 1894 331 1895 335
rect 1899 331 1900 335
rect 1894 330 1900 331
rect 1982 335 1988 336
rect 1982 331 1983 335
rect 1987 331 1988 335
rect 1982 330 1988 331
rect 2070 335 2076 336
rect 2070 331 2071 335
rect 2075 331 2076 335
rect 2070 330 2076 331
rect 2158 335 2164 336
rect 2158 331 2159 335
rect 2163 331 2164 335
rect 2158 330 2164 331
rect 2270 335 2276 336
rect 2270 331 2271 335
rect 2275 331 2276 335
rect 2270 330 2276 331
rect 2390 335 2396 336
rect 2390 331 2391 335
rect 2395 331 2396 335
rect 2390 330 2396 331
rect 2526 335 2532 336
rect 2526 331 2527 335
rect 2531 331 2532 335
rect 2526 330 2532 331
rect 2678 335 2684 336
rect 2678 331 2679 335
rect 2683 331 2684 335
rect 2678 330 2684 331
rect 2854 335 2860 336
rect 2854 331 2855 335
rect 2859 331 2860 335
rect 2854 330 2860 331
rect 3038 335 3044 336
rect 3038 331 3039 335
rect 3043 331 3044 335
rect 3038 330 3044 331
rect 3238 335 3244 336
rect 3238 331 3239 335
rect 3243 331 3244 335
rect 3238 330 3244 331
rect 3438 335 3444 336
rect 3438 331 3439 335
rect 3443 331 3444 335
rect 3438 330 3444 331
rect 134 323 140 324
rect 134 319 135 323
rect 139 319 140 323
rect 134 318 140 319
rect 222 323 228 324
rect 222 319 223 323
rect 227 319 228 323
rect 222 318 228 319
rect 310 323 316 324
rect 310 319 311 323
rect 315 319 316 323
rect 310 318 316 319
rect 398 323 404 324
rect 398 319 399 323
rect 403 319 404 323
rect 398 318 404 319
rect 486 323 492 324
rect 486 319 487 323
rect 491 319 492 323
rect 486 318 492 319
rect 574 323 580 324
rect 574 319 575 323
rect 579 319 580 323
rect 574 318 580 319
rect 662 323 668 324
rect 662 319 663 323
rect 667 319 668 323
rect 662 318 668 319
rect 750 323 756 324
rect 750 319 751 323
rect 755 319 756 323
rect 750 318 756 319
rect 838 323 844 324
rect 838 319 839 323
rect 843 319 844 323
rect 838 318 844 319
rect 926 323 932 324
rect 926 319 927 323
rect 931 319 932 323
rect 926 318 932 319
rect 1014 323 1020 324
rect 1014 319 1015 323
rect 1019 319 1020 323
rect 1014 318 1020 319
rect 1102 323 1108 324
rect 1102 319 1103 323
rect 1107 319 1108 323
rect 1102 318 1108 319
rect 1190 323 1196 324
rect 1190 319 1191 323
rect 1195 319 1196 323
rect 1190 318 1196 319
rect 1286 323 1292 324
rect 1286 319 1287 323
rect 1291 319 1292 323
rect 1286 318 1292 319
rect 1382 323 1388 324
rect 1382 319 1383 323
rect 1387 319 1388 323
rect 1382 318 1388 319
rect 1478 323 1484 324
rect 1478 319 1479 323
rect 1483 319 1484 323
rect 1478 318 1484 319
rect 1574 323 1580 324
rect 1574 319 1575 323
rect 1579 319 1580 323
rect 1574 318 1580 319
rect 1670 323 1676 324
rect 1670 319 1671 323
rect 1675 319 1676 323
rect 1670 318 1676 319
rect 1879 323 1885 324
rect 1879 319 1880 323
rect 1884 322 1885 323
rect 1887 323 1893 324
rect 1887 322 1888 323
rect 1884 320 1888 322
rect 1884 319 1885 320
rect 1879 318 1885 319
rect 1887 319 1888 320
rect 1892 319 1893 323
rect 1887 318 1893 319
rect 1967 323 1973 324
rect 1967 319 1968 323
rect 1972 322 1973 323
rect 1975 323 1981 324
rect 1975 322 1976 323
rect 1972 320 1976 322
rect 1972 319 1973 320
rect 1967 318 1973 319
rect 1975 319 1976 320
rect 1980 319 1981 323
rect 1975 318 1981 319
rect 2055 323 2061 324
rect 2055 319 2056 323
rect 2060 322 2061 323
rect 2063 323 2069 324
rect 2063 322 2064 323
rect 2060 320 2064 322
rect 2060 319 2061 320
rect 2055 318 2061 319
rect 2063 319 2064 320
rect 2068 319 2069 323
rect 2063 318 2069 319
rect 2143 323 2149 324
rect 2143 319 2144 323
rect 2148 322 2149 323
rect 2151 323 2157 324
rect 2151 322 2152 323
rect 2148 320 2152 322
rect 2148 319 2149 320
rect 2143 318 2149 319
rect 2151 319 2152 320
rect 2156 319 2157 323
rect 2151 318 2157 319
rect 2263 323 2269 324
rect 2263 319 2264 323
rect 2268 322 2269 323
rect 2351 323 2357 324
rect 2351 322 2352 323
rect 2268 320 2352 322
rect 2268 319 2269 320
rect 2263 318 2269 319
rect 2351 319 2352 320
rect 2356 319 2357 323
rect 2351 318 2357 319
rect 2383 323 2389 324
rect 2383 319 2384 323
rect 2388 322 2389 323
rect 2450 323 2456 324
rect 2450 322 2451 323
rect 2388 320 2451 322
rect 2388 319 2389 320
rect 2383 318 2389 319
rect 2450 319 2451 320
rect 2455 319 2456 323
rect 2450 318 2456 319
rect 2519 323 2525 324
rect 2519 319 2520 323
rect 2524 322 2525 323
rect 2534 323 2540 324
rect 2534 322 2535 323
rect 2524 320 2535 322
rect 2524 319 2525 320
rect 2519 318 2525 319
rect 2534 319 2535 320
rect 2539 319 2540 323
rect 2534 318 2540 319
rect 2671 323 2677 324
rect 2671 319 2672 323
rect 2676 322 2677 323
rect 2686 323 2692 324
rect 2686 322 2687 323
rect 2676 320 2687 322
rect 2676 319 2677 320
rect 2671 318 2677 319
rect 2686 319 2687 320
rect 2691 319 2692 323
rect 2686 318 2692 319
rect 2839 323 2845 324
rect 2839 319 2840 323
rect 2844 322 2845 323
rect 2847 323 2853 324
rect 2847 322 2848 323
rect 2844 320 2848 322
rect 2844 319 2845 320
rect 2839 318 2845 319
rect 2847 319 2848 320
rect 2852 319 2853 323
rect 2847 318 2853 319
rect 3023 323 3029 324
rect 3023 319 3024 323
rect 3028 322 3029 323
rect 3031 323 3037 324
rect 3031 322 3032 323
rect 3028 320 3032 322
rect 3028 319 3029 320
rect 3023 318 3029 319
rect 3031 319 3032 320
rect 3036 319 3037 323
rect 3031 318 3037 319
rect 3150 323 3156 324
rect 3150 319 3151 323
rect 3155 322 3156 323
rect 3231 323 3237 324
rect 3231 322 3232 323
rect 3155 320 3232 322
rect 3155 319 3156 320
rect 3150 318 3156 319
rect 3231 319 3232 320
rect 3236 319 3237 323
rect 3231 318 3237 319
rect 3426 323 3437 324
rect 3426 319 3427 323
rect 3431 319 3432 323
rect 3436 319 3437 323
rect 3426 318 3437 319
rect 391 315 397 316
rect 110 313 116 314
rect 110 309 111 313
rect 115 309 116 313
rect 391 311 392 315
rect 396 314 397 315
rect 730 315 736 316
rect 396 312 417 314
rect 396 311 397 312
rect 391 310 397 311
rect 730 311 731 315
rect 735 314 736 315
rect 1082 315 1088 316
rect 1082 314 1083 315
rect 735 312 769 314
rect 1073 312 1083 314
rect 735 311 736 312
rect 730 310 736 311
rect 1082 311 1083 312
rect 1087 311 1088 315
rect 1082 310 1088 311
rect 1822 313 1828 314
rect 110 308 116 309
rect 1822 309 1823 313
rect 1827 309 1828 313
rect 1822 308 1828 309
rect 1887 311 1893 312
rect 1887 307 1888 311
rect 1892 310 1893 311
rect 1902 311 1908 312
rect 1902 310 1903 311
rect 1892 308 1903 310
rect 1892 307 1893 308
rect 1887 306 1893 307
rect 1902 307 1903 308
rect 1907 307 1908 311
rect 1902 306 1908 307
rect 1959 311 1965 312
rect 1959 307 1960 311
rect 1964 310 1965 311
rect 1975 311 1981 312
rect 1975 310 1976 311
rect 1964 308 1976 310
rect 1964 307 1965 308
rect 1959 306 1965 307
rect 1975 307 1976 308
rect 1980 307 1981 311
rect 1975 306 1981 307
rect 2047 311 2053 312
rect 2047 307 2048 311
rect 2052 310 2053 311
rect 2063 311 2069 312
rect 2063 310 2064 311
rect 2052 308 2064 310
rect 2052 307 2053 308
rect 2047 306 2053 307
rect 2063 307 2064 308
rect 2068 307 2069 311
rect 2063 306 2069 307
rect 2135 311 2141 312
rect 2135 307 2136 311
rect 2140 310 2141 311
rect 2151 311 2157 312
rect 2151 310 2152 311
rect 2140 308 2152 310
rect 2140 307 2141 308
rect 2135 306 2141 307
rect 2151 307 2152 308
rect 2156 307 2157 311
rect 2151 306 2157 307
rect 2223 311 2229 312
rect 2223 307 2224 311
rect 2228 310 2229 311
rect 2239 311 2245 312
rect 2239 310 2240 311
rect 2228 308 2240 310
rect 2228 307 2229 308
rect 2223 306 2229 307
rect 2239 307 2240 308
rect 2244 307 2245 311
rect 2239 306 2245 307
rect 2351 311 2357 312
rect 2351 307 2352 311
rect 2356 310 2357 311
rect 2366 311 2372 312
rect 2366 310 2367 311
rect 2356 308 2367 310
rect 2356 307 2357 308
rect 2351 306 2357 307
rect 2366 307 2367 308
rect 2371 307 2372 311
rect 2366 306 2372 307
rect 2423 311 2429 312
rect 2423 307 2424 311
rect 2428 310 2429 311
rect 2463 311 2469 312
rect 2463 310 2464 311
rect 2428 308 2464 310
rect 2428 307 2429 308
rect 2423 306 2429 307
rect 2463 307 2464 308
rect 2468 307 2469 311
rect 2463 306 2469 307
rect 2575 311 2581 312
rect 2575 307 2576 311
rect 2580 310 2581 311
rect 2602 311 2608 312
rect 2602 310 2603 311
rect 2580 308 2603 310
rect 2580 307 2581 308
rect 2575 306 2581 307
rect 2602 307 2603 308
rect 2607 307 2608 311
rect 2602 306 2608 307
rect 2687 311 2693 312
rect 2687 307 2688 311
rect 2692 310 2693 311
rect 2702 311 2708 312
rect 2702 310 2703 311
rect 2692 308 2703 310
rect 2692 307 2693 308
rect 2687 306 2693 307
rect 2702 307 2703 308
rect 2707 307 2708 311
rect 2702 306 2708 307
rect 2759 311 2765 312
rect 2759 307 2760 311
rect 2764 310 2765 311
rect 2799 311 2805 312
rect 2799 310 2800 311
rect 2764 308 2800 310
rect 2764 307 2765 308
rect 2759 306 2765 307
rect 2799 307 2800 308
rect 2804 307 2805 311
rect 2799 306 2805 307
rect 2871 311 2877 312
rect 2871 307 2872 311
rect 2876 310 2877 311
rect 2911 311 2917 312
rect 2911 310 2912 311
rect 2876 308 2912 310
rect 2876 307 2877 308
rect 2871 306 2877 307
rect 2911 307 2912 308
rect 2916 307 2917 311
rect 2911 306 2917 307
rect 2983 311 2989 312
rect 2983 307 2984 311
rect 2988 310 2989 311
rect 3031 311 3037 312
rect 3031 310 3032 311
rect 2988 308 3032 310
rect 2988 307 2989 308
rect 2983 306 2989 307
rect 3031 307 3032 308
rect 3036 307 3037 311
rect 3031 306 3037 307
rect 3103 311 3109 312
rect 3103 307 3104 311
rect 3108 310 3109 311
rect 3151 311 3157 312
rect 3151 310 3152 311
rect 3108 308 3152 310
rect 3108 307 3109 308
rect 3103 306 3109 307
rect 3151 307 3152 308
rect 3156 307 3157 311
rect 3151 306 3157 307
rect 1894 301 1900 302
rect 215 299 221 300
rect 215 298 216 299
rect 110 296 116 297
rect 197 296 216 298
rect 110 292 111 296
rect 115 292 116 296
rect 215 295 216 296
rect 220 295 221 299
rect 303 299 309 300
rect 303 298 304 299
rect 285 296 304 298
rect 215 294 221 295
rect 303 295 304 296
rect 308 295 309 299
rect 391 299 397 300
rect 391 298 392 299
rect 373 296 392 298
rect 303 294 309 295
rect 391 295 392 296
rect 396 295 397 299
rect 567 299 573 300
rect 567 298 568 299
rect 549 296 568 298
rect 391 294 397 295
rect 567 295 568 296
rect 572 295 573 299
rect 655 299 661 300
rect 655 298 656 299
rect 637 296 656 298
rect 567 294 573 295
rect 655 295 656 296
rect 660 295 661 299
rect 743 299 749 300
rect 743 298 744 299
rect 725 296 744 298
rect 655 294 661 295
rect 743 295 744 296
rect 748 295 749 299
rect 743 294 749 295
rect 818 299 824 300
rect 818 295 819 299
rect 823 298 824 299
rect 1007 299 1013 300
rect 1007 298 1008 299
rect 823 296 865 298
rect 989 296 1008 298
rect 823 295 824 296
rect 818 294 824 295
rect 1007 295 1008 296
rect 1012 295 1013 299
rect 1007 294 1013 295
rect 1082 299 1088 300
rect 1082 295 1083 299
rect 1087 298 1088 299
rect 1170 299 1176 300
rect 1087 296 1129 298
rect 1087 295 1088 296
rect 1082 294 1088 295
rect 1170 295 1171 299
rect 1175 298 1176 299
rect 1375 299 1381 300
rect 1375 298 1376 299
rect 1175 296 1217 298
rect 1349 296 1376 298
rect 1175 295 1176 296
rect 1170 294 1176 295
rect 1375 295 1376 296
rect 1380 295 1381 299
rect 1471 299 1477 300
rect 1471 298 1472 299
rect 1445 296 1472 298
rect 1375 294 1381 295
rect 1471 295 1472 296
rect 1476 295 1477 299
rect 1551 299 1557 300
rect 1551 298 1552 299
rect 1541 296 1552 298
rect 1471 294 1477 295
rect 1551 295 1552 296
rect 1556 295 1557 299
rect 1551 294 1557 295
rect 1562 299 1568 300
rect 1562 295 1563 299
rect 1567 298 1568 299
rect 1642 299 1648 300
rect 1567 296 1601 298
rect 1567 295 1568 296
rect 1562 294 1568 295
rect 1642 295 1643 299
rect 1647 298 1648 299
rect 1647 296 1697 298
rect 1894 297 1895 301
rect 1899 297 1900 301
rect 1822 296 1828 297
rect 1894 296 1900 297
rect 1982 301 1988 302
rect 1982 297 1983 301
rect 1987 297 1988 301
rect 1982 296 1988 297
rect 2070 301 2076 302
rect 2070 297 2071 301
rect 2075 297 2076 301
rect 2070 296 2076 297
rect 2158 301 2164 302
rect 2158 297 2159 301
rect 2163 297 2164 301
rect 2158 296 2164 297
rect 2246 301 2252 302
rect 2246 297 2247 301
rect 2251 297 2252 301
rect 2246 296 2252 297
rect 2358 301 2364 302
rect 2358 297 2359 301
rect 2363 297 2364 301
rect 2358 296 2364 297
rect 2470 301 2476 302
rect 2470 297 2471 301
rect 2475 297 2476 301
rect 2470 296 2476 297
rect 2582 301 2588 302
rect 2582 297 2583 301
rect 2587 297 2588 301
rect 2582 296 2588 297
rect 2694 301 2700 302
rect 2694 297 2695 301
rect 2699 297 2700 301
rect 2694 296 2700 297
rect 2806 301 2812 302
rect 2806 297 2807 301
rect 2811 297 2812 301
rect 2806 296 2812 297
rect 2918 301 2924 302
rect 2918 297 2919 301
rect 2923 297 2924 301
rect 2918 296 2924 297
rect 3038 301 3044 302
rect 3038 297 3039 301
rect 3043 297 3044 301
rect 3038 296 3044 297
rect 3158 301 3164 302
rect 3158 297 3159 301
rect 3163 297 3164 301
rect 3158 296 3164 297
rect 1647 295 1648 296
rect 1642 294 1648 295
rect 110 291 116 292
rect 1822 292 1823 296
rect 1827 292 1828 296
rect 1822 291 1828 292
rect 1862 288 1868 289
rect 3574 288 3580 289
rect 1862 284 1863 288
rect 1867 284 1868 288
rect 1959 287 1965 288
rect 1959 286 1960 287
rect 1949 284 1960 286
rect 142 283 148 284
rect 142 279 143 283
rect 147 279 148 283
rect 142 278 148 279
rect 230 283 236 284
rect 230 279 231 283
rect 235 279 236 283
rect 230 278 236 279
rect 318 283 324 284
rect 318 279 319 283
rect 323 279 324 283
rect 318 278 324 279
rect 406 283 412 284
rect 406 279 407 283
rect 411 279 412 283
rect 406 278 412 279
rect 494 283 500 284
rect 494 279 495 283
rect 499 279 500 283
rect 494 278 500 279
rect 582 283 588 284
rect 582 279 583 283
rect 587 279 588 283
rect 582 278 588 279
rect 670 283 676 284
rect 670 279 671 283
rect 675 279 676 283
rect 670 278 676 279
rect 758 283 764 284
rect 758 279 759 283
rect 763 279 764 283
rect 758 278 764 279
rect 846 283 852 284
rect 846 279 847 283
rect 851 279 852 283
rect 846 278 852 279
rect 934 283 940 284
rect 934 279 935 283
rect 939 279 940 283
rect 934 278 940 279
rect 1022 283 1028 284
rect 1022 279 1023 283
rect 1027 279 1028 283
rect 1022 278 1028 279
rect 1110 283 1116 284
rect 1110 279 1111 283
rect 1115 279 1116 283
rect 1110 278 1116 279
rect 1198 283 1204 284
rect 1198 279 1199 283
rect 1203 279 1204 283
rect 1198 278 1204 279
rect 1294 283 1300 284
rect 1294 279 1295 283
rect 1299 279 1300 283
rect 1294 278 1300 279
rect 1390 283 1396 284
rect 1390 279 1391 283
rect 1395 279 1396 283
rect 1390 278 1396 279
rect 1486 283 1492 284
rect 1486 279 1487 283
rect 1491 279 1492 283
rect 1486 278 1492 279
rect 1582 283 1588 284
rect 1582 279 1583 283
rect 1587 279 1588 283
rect 1582 278 1588 279
rect 1678 283 1684 284
rect 1862 283 1868 284
rect 1959 283 1960 284
rect 1964 283 1965 287
rect 2047 287 2053 288
rect 2047 286 2048 287
rect 2037 284 2048 286
rect 1678 279 1679 283
rect 1683 279 1684 283
rect 1959 282 1965 283
rect 2047 283 2048 284
rect 2052 283 2053 287
rect 2135 287 2141 288
rect 2135 286 2136 287
rect 2125 284 2136 286
rect 2047 282 2053 283
rect 2135 283 2136 284
rect 2140 283 2141 287
rect 2223 287 2229 288
rect 2223 286 2224 287
rect 2213 284 2224 286
rect 2135 282 2141 283
rect 2223 283 2224 284
rect 2228 283 2229 287
rect 2423 287 2429 288
rect 2423 286 2424 287
rect 2413 284 2424 286
rect 2223 282 2229 283
rect 2423 283 2424 284
rect 2428 283 2429 287
rect 2534 287 2540 288
rect 2534 286 2535 287
rect 2525 284 2535 286
rect 2423 282 2429 283
rect 2534 283 2535 284
rect 2539 283 2540 287
rect 2759 287 2765 288
rect 2759 286 2760 287
rect 2749 284 2760 286
rect 2534 282 2540 283
rect 2542 283 2548 284
rect 1678 278 1684 279
rect 2542 279 2543 283
rect 2547 282 2548 283
rect 2759 283 2760 284
rect 2764 283 2765 287
rect 2871 287 2877 288
rect 2871 286 2872 287
rect 2861 284 2872 286
rect 2759 282 2765 283
rect 2871 283 2872 284
rect 2876 283 2877 287
rect 2983 287 2989 288
rect 2983 286 2984 287
rect 2973 284 2984 286
rect 2871 282 2877 283
rect 2983 283 2984 284
rect 2988 283 2989 287
rect 3103 287 3109 288
rect 3103 286 3104 287
rect 3093 284 3104 286
rect 2983 282 2989 283
rect 3103 283 3104 284
rect 3108 283 3109 287
rect 3574 284 3575 288
rect 3579 284 3580 288
rect 3574 283 3580 284
rect 3103 282 3109 283
rect 2547 280 2601 282
rect 2547 279 2548 280
rect 2542 278 2548 279
rect 134 271 141 272
rect 134 267 135 271
rect 140 267 141 271
rect 134 266 141 267
rect 215 271 221 272
rect 215 267 216 271
rect 220 270 221 271
rect 223 271 229 272
rect 223 270 224 271
rect 220 268 224 270
rect 220 267 221 268
rect 215 266 221 267
rect 223 267 224 268
rect 228 267 229 271
rect 223 266 229 267
rect 303 271 309 272
rect 303 267 304 271
rect 308 270 309 271
rect 311 271 317 272
rect 311 270 312 271
rect 308 268 312 270
rect 308 267 309 268
rect 303 266 309 267
rect 311 267 312 268
rect 316 267 317 271
rect 311 266 317 267
rect 391 271 397 272
rect 391 267 392 271
rect 396 270 397 271
rect 399 271 405 272
rect 399 270 400 271
rect 396 268 400 270
rect 396 267 397 268
rect 391 266 397 267
rect 399 267 400 268
rect 404 267 405 271
rect 399 266 405 267
rect 487 271 493 272
rect 487 267 488 271
rect 492 270 493 271
rect 567 271 573 272
rect 492 268 558 270
rect 492 267 493 268
rect 487 266 493 267
rect 556 262 558 268
rect 567 267 568 271
rect 572 270 573 271
rect 575 271 581 272
rect 575 270 576 271
rect 572 268 576 270
rect 572 267 573 268
rect 567 266 573 267
rect 575 267 576 268
rect 580 267 581 271
rect 575 266 581 267
rect 655 271 661 272
rect 655 267 656 271
rect 660 270 661 271
rect 663 271 669 272
rect 663 270 664 271
rect 660 268 664 270
rect 660 267 661 268
rect 655 266 661 267
rect 663 267 664 268
rect 668 267 669 271
rect 663 266 669 267
rect 751 271 757 272
rect 751 267 752 271
rect 756 270 757 271
rect 818 271 824 272
rect 818 270 819 271
rect 756 268 819 270
rect 756 267 757 268
rect 751 266 757 267
rect 818 267 819 268
rect 823 267 824 271
rect 818 266 824 267
rect 839 271 845 272
rect 839 267 840 271
rect 844 270 845 271
rect 854 271 860 272
rect 854 270 855 271
rect 844 268 855 270
rect 844 267 845 268
rect 839 266 845 267
rect 854 267 855 268
rect 859 267 860 271
rect 854 266 860 267
rect 927 271 933 272
rect 927 267 928 271
rect 932 270 933 271
rect 1007 271 1013 272
rect 932 268 1002 270
rect 932 267 933 268
rect 927 266 933 267
rect 730 263 736 264
rect 730 262 731 263
rect 556 260 731 262
rect 730 259 731 260
rect 735 259 736 263
rect 730 258 736 259
rect 738 263 744 264
rect 738 259 739 263
rect 743 262 744 263
rect 919 263 925 264
rect 919 262 920 263
rect 743 260 920 262
rect 743 259 744 260
rect 738 258 744 259
rect 919 259 920 260
rect 924 259 925 263
rect 1000 262 1002 268
rect 1007 267 1008 271
rect 1012 270 1013 271
rect 1015 271 1021 272
rect 1015 270 1016 271
rect 1012 268 1016 270
rect 1012 267 1013 268
rect 1007 266 1013 267
rect 1015 267 1016 268
rect 1020 267 1021 271
rect 1015 266 1021 267
rect 1103 271 1109 272
rect 1103 267 1104 271
rect 1108 270 1109 271
rect 1170 271 1176 272
rect 1170 270 1171 271
rect 1108 268 1171 270
rect 1108 267 1109 268
rect 1103 266 1109 267
rect 1170 267 1171 268
rect 1175 267 1176 271
rect 1170 266 1176 267
rect 1190 271 1197 272
rect 1190 267 1191 271
rect 1196 267 1197 271
rect 1190 266 1197 267
rect 1287 271 1293 272
rect 1287 267 1288 271
rect 1292 270 1293 271
rect 1302 271 1308 272
rect 1302 270 1303 271
rect 1292 268 1303 270
rect 1292 267 1293 268
rect 1287 266 1293 267
rect 1302 267 1303 268
rect 1307 267 1308 271
rect 1302 266 1308 267
rect 1375 271 1381 272
rect 1375 267 1376 271
rect 1380 270 1381 271
rect 1383 271 1389 272
rect 1383 270 1384 271
rect 1380 268 1384 270
rect 1380 267 1381 268
rect 1375 266 1381 267
rect 1383 267 1384 268
rect 1388 267 1389 271
rect 1383 266 1389 267
rect 1471 271 1477 272
rect 1471 267 1472 271
rect 1476 270 1477 271
rect 1479 271 1485 272
rect 1479 270 1480 271
rect 1476 268 1480 270
rect 1476 267 1477 268
rect 1471 266 1477 267
rect 1479 267 1480 268
rect 1484 267 1485 271
rect 1479 266 1485 267
rect 1575 271 1581 272
rect 1575 267 1576 271
rect 1580 270 1581 271
rect 1642 271 1648 272
rect 1642 270 1643 271
rect 1580 268 1643 270
rect 1580 267 1581 268
rect 1575 266 1581 267
rect 1642 267 1643 268
rect 1647 267 1648 271
rect 1642 266 1648 267
rect 1663 271 1669 272
rect 1663 267 1664 271
rect 1668 270 1669 271
rect 1671 271 1677 272
rect 1671 270 1672 271
rect 1668 268 1672 270
rect 1668 267 1669 268
rect 1663 266 1669 267
rect 1671 267 1672 268
rect 1676 267 1677 271
rect 1671 266 1677 267
rect 1862 271 1868 272
rect 1862 267 1863 271
rect 1867 267 1868 271
rect 1862 266 1868 267
rect 2226 271 2232 272
rect 2226 267 2227 271
rect 2231 270 2232 271
rect 3106 271 3112 272
rect 2231 268 2257 270
rect 2231 267 2232 268
rect 2226 266 2232 267
rect 3106 267 3107 271
rect 3111 270 3112 271
rect 3574 271 3580 272
rect 3111 268 3169 270
rect 3111 267 3112 268
rect 3106 266 3112 267
rect 3574 267 3575 271
rect 3579 267 3580 271
rect 3574 266 3580 267
rect 1082 263 1088 264
rect 1082 262 1083 263
rect 1000 260 1083 262
rect 919 258 925 259
rect 1082 259 1083 260
rect 1087 259 1088 263
rect 1082 258 1088 259
rect 1886 261 1892 262
rect 1886 257 1887 261
rect 1891 257 1892 261
rect 1886 256 1892 257
rect 1974 261 1980 262
rect 1974 257 1975 261
rect 1979 257 1980 261
rect 1974 256 1980 257
rect 2062 261 2068 262
rect 2062 257 2063 261
rect 2067 257 2068 261
rect 2062 256 2068 257
rect 2150 261 2156 262
rect 2150 257 2151 261
rect 2155 257 2156 261
rect 2150 256 2156 257
rect 2238 261 2244 262
rect 2238 257 2239 261
rect 2243 257 2244 261
rect 2238 256 2244 257
rect 2350 261 2356 262
rect 2350 257 2351 261
rect 2355 257 2356 261
rect 2350 256 2356 257
rect 2462 261 2468 262
rect 2462 257 2463 261
rect 2467 257 2468 261
rect 2462 256 2468 257
rect 2574 261 2580 262
rect 2574 257 2575 261
rect 2579 257 2580 261
rect 2574 256 2580 257
rect 2686 261 2692 262
rect 2686 257 2687 261
rect 2691 257 2692 261
rect 2686 256 2692 257
rect 2798 261 2804 262
rect 2798 257 2799 261
rect 2803 257 2804 261
rect 2798 256 2804 257
rect 2910 261 2916 262
rect 2910 257 2911 261
rect 2915 257 2916 261
rect 2910 256 2916 257
rect 3030 261 3036 262
rect 3030 257 3031 261
rect 3035 257 3036 261
rect 3030 256 3036 257
rect 3150 261 3156 262
rect 3150 257 3151 261
rect 3155 257 3156 261
rect 3150 256 3156 257
rect 135 255 141 256
rect 135 251 136 255
rect 140 254 141 255
rect 210 255 216 256
rect 210 254 211 255
rect 140 252 211 254
rect 140 251 141 252
rect 135 250 141 251
rect 210 251 211 252
rect 215 251 216 255
rect 210 250 216 251
rect 223 255 229 256
rect 223 251 224 255
rect 228 254 229 255
rect 298 255 304 256
rect 298 254 299 255
rect 228 252 299 254
rect 228 251 229 252
rect 223 250 229 251
rect 298 251 299 252
rect 303 251 304 255
rect 298 250 304 251
rect 311 255 317 256
rect 311 251 312 255
rect 316 254 317 255
rect 386 255 392 256
rect 386 254 387 255
rect 316 252 387 254
rect 316 251 317 252
rect 311 250 317 251
rect 386 251 387 252
rect 391 251 392 255
rect 386 250 392 251
rect 399 255 405 256
rect 399 251 400 255
rect 404 254 405 255
rect 474 255 480 256
rect 474 254 475 255
rect 404 252 475 254
rect 404 251 405 252
rect 399 250 405 251
rect 474 251 475 252
rect 479 251 480 255
rect 474 250 480 251
rect 487 255 493 256
rect 487 251 488 255
rect 492 254 493 255
rect 562 255 568 256
rect 562 254 563 255
rect 492 252 563 254
rect 492 251 493 252
rect 487 250 493 251
rect 562 251 563 252
rect 567 251 568 255
rect 562 250 568 251
rect 575 255 581 256
rect 575 251 576 255
rect 580 254 581 255
rect 650 255 656 256
rect 650 254 651 255
rect 580 252 651 254
rect 580 251 581 252
rect 575 250 581 251
rect 650 251 651 252
rect 655 251 656 255
rect 650 250 656 251
rect 663 255 669 256
rect 663 251 664 255
rect 668 254 669 255
rect 734 255 740 256
rect 734 254 735 255
rect 668 252 735 254
rect 668 251 669 252
rect 663 250 669 251
rect 734 251 735 252
rect 739 251 740 255
rect 734 250 740 251
rect 743 255 749 256
rect 743 251 744 255
rect 748 254 749 255
rect 751 255 757 256
rect 751 254 752 255
rect 748 252 752 254
rect 748 251 749 252
rect 743 250 749 251
rect 751 251 752 252
rect 756 251 757 255
rect 751 250 757 251
rect 823 255 829 256
rect 823 251 824 255
rect 828 254 829 255
rect 839 255 845 256
rect 839 254 840 255
rect 828 252 840 254
rect 828 251 829 252
rect 823 250 829 251
rect 839 251 840 252
rect 844 251 845 255
rect 839 250 845 251
rect 911 255 917 256
rect 911 251 912 255
rect 916 254 917 255
rect 927 255 933 256
rect 927 254 928 255
rect 916 252 928 254
rect 916 251 917 252
rect 911 250 917 251
rect 927 251 928 252
rect 932 251 933 255
rect 927 250 933 251
rect 1015 255 1021 256
rect 1015 251 1016 255
rect 1020 254 1021 255
rect 1030 255 1036 256
rect 1030 254 1031 255
rect 1020 252 1031 254
rect 1020 251 1021 252
rect 1015 250 1021 251
rect 1030 251 1031 252
rect 1035 251 1036 255
rect 1030 250 1036 251
rect 1087 255 1093 256
rect 1087 251 1088 255
rect 1092 254 1093 255
rect 1103 255 1109 256
rect 1103 254 1104 255
rect 1092 252 1104 254
rect 1092 251 1093 252
rect 1087 250 1093 251
rect 1103 251 1104 252
rect 1108 251 1109 255
rect 1103 250 1109 251
rect 1175 255 1181 256
rect 1175 251 1176 255
rect 1180 254 1181 255
rect 1191 255 1197 256
rect 1191 254 1192 255
rect 1180 252 1192 254
rect 1180 251 1181 252
rect 1175 250 1181 251
rect 1191 251 1192 252
rect 1196 251 1197 255
rect 1191 250 1197 251
rect 1279 255 1285 256
rect 1279 251 1280 255
rect 1284 254 1285 255
rect 1354 255 1360 256
rect 1354 254 1355 255
rect 1284 252 1355 254
rect 1284 251 1285 252
rect 1279 250 1285 251
rect 1354 251 1355 252
rect 1359 251 1360 255
rect 1354 250 1360 251
rect 1367 255 1373 256
rect 1367 251 1368 255
rect 1372 254 1373 255
rect 1442 255 1448 256
rect 1442 254 1443 255
rect 1372 252 1443 254
rect 1372 251 1373 252
rect 1367 250 1373 251
rect 1442 251 1443 252
rect 1447 251 1448 255
rect 1442 250 1448 251
rect 1455 255 1461 256
rect 1455 251 1456 255
rect 1460 254 1461 255
rect 1534 255 1540 256
rect 1534 254 1535 255
rect 1460 252 1535 254
rect 1460 251 1461 252
rect 1455 250 1461 251
rect 1534 251 1535 252
rect 1539 251 1540 255
rect 1534 250 1540 251
rect 1543 255 1549 256
rect 1543 251 1544 255
rect 1548 254 1549 255
rect 1551 255 1557 256
rect 1551 254 1552 255
rect 1548 252 1552 254
rect 1548 251 1549 252
rect 1543 250 1549 251
rect 1551 251 1552 252
rect 1556 251 1557 255
rect 1551 250 1557 251
rect 1615 255 1621 256
rect 1615 251 1616 255
rect 1620 254 1621 255
rect 1631 255 1637 256
rect 1631 254 1632 255
rect 1620 252 1632 254
rect 1620 251 1621 252
rect 1615 250 1621 251
rect 1631 251 1632 252
rect 1636 251 1637 255
rect 1631 250 1637 251
rect 1706 255 1712 256
rect 1706 251 1707 255
rect 1711 254 1712 255
rect 1719 255 1725 256
rect 1719 254 1720 255
rect 1711 252 1720 254
rect 1711 251 1712 252
rect 1706 250 1712 251
rect 1719 251 1720 252
rect 1724 251 1725 255
rect 1719 250 1725 251
rect 142 245 148 246
rect 142 241 143 245
rect 147 241 148 245
rect 142 240 148 241
rect 230 245 236 246
rect 230 241 231 245
rect 235 241 236 245
rect 230 240 236 241
rect 318 245 324 246
rect 318 241 319 245
rect 323 241 324 245
rect 318 240 324 241
rect 406 245 412 246
rect 406 241 407 245
rect 411 241 412 245
rect 406 240 412 241
rect 494 245 500 246
rect 494 241 495 245
rect 499 241 500 245
rect 494 240 500 241
rect 582 245 588 246
rect 582 241 583 245
rect 587 241 588 245
rect 582 240 588 241
rect 670 245 676 246
rect 670 241 671 245
rect 675 241 676 245
rect 670 240 676 241
rect 758 245 764 246
rect 758 241 759 245
rect 763 241 764 245
rect 758 240 764 241
rect 846 245 852 246
rect 846 241 847 245
rect 851 241 852 245
rect 846 240 852 241
rect 934 245 940 246
rect 934 241 935 245
rect 939 241 940 245
rect 934 240 940 241
rect 1022 245 1028 246
rect 1022 241 1023 245
rect 1027 241 1028 245
rect 1022 240 1028 241
rect 1110 245 1116 246
rect 1110 241 1111 245
rect 1115 241 1116 245
rect 1110 240 1116 241
rect 1198 245 1204 246
rect 1198 241 1199 245
rect 1203 241 1204 245
rect 1198 240 1204 241
rect 1286 245 1292 246
rect 1286 241 1287 245
rect 1291 241 1292 245
rect 1286 240 1292 241
rect 1374 245 1380 246
rect 1374 241 1375 245
rect 1379 241 1380 245
rect 1374 240 1380 241
rect 1462 245 1468 246
rect 1462 241 1463 245
rect 1467 241 1468 245
rect 1462 240 1468 241
rect 1550 245 1556 246
rect 1550 241 1551 245
rect 1555 241 1556 245
rect 1550 240 1556 241
rect 1638 245 1644 246
rect 1638 241 1639 245
rect 1643 241 1644 245
rect 1638 240 1644 241
rect 1726 245 1732 246
rect 1726 241 1727 245
rect 1731 241 1732 245
rect 1726 240 1732 241
rect 1886 239 1892 240
rect 1886 235 1887 239
rect 1891 235 1892 239
rect 1886 234 1892 235
rect 1974 239 1980 240
rect 1974 235 1975 239
rect 1979 235 1980 239
rect 1974 234 1980 235
rect 2062 239 2068 240
rect 2062 235 2063 239
rect 2067 235 2068 239
rect 2062 234 2068 235
rect 2150 239 2156 240
rect 2150 235 2151 239
rect 2155 235 2156 239
rect 2150 234 2156 235
rect 2262 239 2268 240
rect 2262 235 2263 239
rect 2267 235 2268 239
rect 2262 234 2268 235
rect 2398 239 2404 240
rect 2398 235 2399 239
rect 2403 235 2404 239
rect 2398 234 2404 235
rect 2534 239 2540 240
rect 2534 235 2535 239
rect 2539 235 2540 239
rect 2534 234 2540 235
rect 2678 239 2684 240
rect 2678 235 2679 239
rect 2683 235 2684 239
rect 2678 234 2684 235
rect 2814 239 2820 240
rect 2814 235 2815 239
rect 2819 235 2820 239
rect 2814 234 2820 235
rect 2950 239 2956 240
rect 2950 235 2951 239
rect 2955 235 2956 239
rect 2950 234 2956 235
rect 3086 239 3092 240
rect 3086 235 3087 239
rect 3091 235 3092 239
rect 3086 234 3092 235
rect 3222 239 3228 240
rect 3222 235 3223 239
rect 3227 235 3228 239
rect 3222 234 3228 235
rect 3358 239 3364 240
rect 3358 235 3359 239
rect 3363 235 3364 239
rect 3358 234 3364 235
rect 3478 239 3484 240
rect 3478 235 3479 239
rect 3483 235 3484 239
rect 3478 234 3484 235
rect 110 232 116 233
rect 1822 232 1828 233
rect 110 228 111 232
rect 115 228 116 232
rect 823 231 829 232
rect 823 230 824 231
rect 813 228 824 230
rect 110 227 116 228
rect 134 227 140 228
rect 134 223 135 227
rect 139 226 140 227
rect 210 227 216 228
rect 139 224 161 226
rect 139 223 140 224
rect 134 222 140 223
rect 210 223 211 227
rect 215 226 216 227
rect 298 227 304 228
rect 215 224 249 226
rect 215 223 216 224
rect 210 222 216 223
rect 298 223 299 227
rect 303 226 304 227
rect 386 227 392 228
rect 303 224 337 226
rect 303 223 304 224
rect 298 222 304 223
rect 386 223 387 227
rect 391 226 392 227
rect 474 227 480 228
rect 391 224 425 226
rect 391 223 392 224
rect 386 222 392 223
rect 474 223 475 227
rect 479 226 480 227
rect 562 227 568 228
rect 479 224 513 226
rect 479 223 480 224
rect 474 222 480 223
rect 562 223 563 227
rect 567 226 568 227
rect 650 227 656 228
rect 567 224 601 226
rect 567 223 568 224
rect 562 222 568 223
rect 650 223 651 227
rect 655 226 656 227
rect 823 227 824 228
rect 828 227 829 231
rect 911 231 917 232
rect 911 230 912 231
rect 901 228 912 230
rect 823 226 829 227
rect 911 227 912 228
rect 916 227 917 231
rect 1087 231 1093 232
rect 1087 230 1088 231
rect 1077 228 1088 230
rect 911 226 917 227
rect 919 227 925 228
rect 655 224 689 226
rect 655 223 656 224
rect 650 222 656 223
rect 919 223 920 227
rect 924 226 925 227
rect 1087 227 1088 228
rect 1092 227 1093 231
rect 1175 231 1181 232
rect 1175 230 1176 231
rect 1165 228 1176 230
rect 1087 226 1093 227
rect 1175 227 1176 228
rect 1180 227 1181 231
rect 1615 231 1621 232
rect 1615 230 1616 231
rect 1605 228 1616 230
rect 1175 226 1181 227
rect 1190 227 1196 228
rect 924 224 953 226
rect 924 223 925 224
rect 919 222 925 223
rect 1190 223 1191 227
rect 1195 226 1196 227
rect 1266 227 1272 228
rect 1195 224 1217 226
rect 1195 223 1196 224
rect 1190 222 1196 223
rect 1266 223 1267 227
rect 1271 226 1272 227
rect 1354 227 1360 228
rect 1271 224 1305 226
rect 1271 223 1272 224
rect 1266 222 1272 223
rect 1354 223 1355 227
rect 1359 226 1360 227
rect 1442 227 1448 228
rect 1359 224 1393 226
rect 1359 223 1360 224
rect 1354 222 1360 223
rect 1442 223 1443 227
rect 1447 226 1448 227
rect 1615 227 1616 228
rect 1620 227 1621 231
rect 1822 228 1823 232
rect 1827 228 1828 232
rect 2602 231 2608 232
rect 1822 227 1828 228
rect 1862 229 1868 230
rect 1615 226 1621 227
rect 1447 224 1481 226
rect 1862 225 1863 229
rect 1867 225 1868 229
rect 2602 227 2603 231
rect 2607 230 2608 231
rect 3190 231 3196 232
rect 2607 228 2697 230
rect 2607 227 2608 228
rect 2602 226 2608 227
rect 3190 227 3191 231
rect 3195 230 3196 231
rect 3426 231 3432 232
rect 3426 230 3427 231
rect 3195 228 3241 230
rect 3417 228 3427 230
rect 3195 227 3196 228
rect 3190 226 3196 227
rect 3426 227 3427 228
rect 3431 227 3432 231
rect 3426 226 3432 227
rect 3574 229 3580 230
rect 1862 224 1868 225
rect 3574 225 3575 229
rect 3579 225 3580 229
rect 3574 224 3580 225
rect 1447 223 1448 224
rect 1442 222 1448 223
rect 110 215 116 216
rect 110 211 111 215
rect 115 211 116 215
rect 1706 215 1712 216
rect 1706 214 1707 215
rect 1689 212 1707 214
rect 110 210 116 211
rect 1706 211 1707 212
rect 1711 211 1712 215
rect 1706 210 1712 211
rect 1726 215 1732 216
rect 1726 211 1727 215
rect 1731 214 1732 215
rect 1822 215 1828 216
rect 1731 212 1737 214
rect 1731 211 1732 212
rect 1726 210 1732 211
rect 1822 211 1823 215
rect 1827 211 1828 215
rect 1967 215 1973 216
rect 1967 214 1968 215
rect 1822 210 1828 211
rect 1862 212 1868 213
rect 1949 212 1968 214
rect 1862 208 1863 212
rect 1867 208 1868 212
rect 1967 211 1968 212
rect 1972 211 1973 215
rect 2055 215 2061 216
rect 2055 214 2056 215
rect 2037 212 2056 214
rect 1967 210 1973 211
rect 2055 211 2056 212
rect 2060 211 2061 215
rect 2143 215 2149 216
rect 2143 214 2144 215
rect 2125 212 2144 214
rect 2055 210 2061 211
rect 2143 211 2144 212
rect 2148 211 2149 215
rect 2255 215 2261 216
rect 2255 214 2256 215
rect 2213 212 2256 214
rect 2143 210 2149 211
rect 2255 211 2256 212
rect 2260 211 2261 215
rect 2391 215 2397 216
rect 2391 214 2392 215
rect 2325 212 2392 214
rect 2255 210 2261 211
rect 2391 211 2392 212
rect 2396 211 2397 215
rect 2527 215 2533 216
rect 2527 214 2528 215
rect 2461 212 2528 214
rect 2391 210 2397 211
rect 2527 211 2528 212
rect 2532 211 2533 215
rect 2671 215 2677 216
rect 2671 214 2672 215
rect 2597 212 2672 214
rect 2527 210 2533 211
rect 2671 211 2672 212
rect 2676 211 2677 215
rect 2943 215 2949 216
rect 2943 214 2944 215
rect 2877 212 2944 214
rect 2671 210 2677 211
rect 2943 211 2944 212
rect 2948 211 2949 215
rect 3079 215 3085 216
rect 3079 214 3080 215
rect 3013 212 3080 214
rect 2943 210 2949 211
rect 3079 211 3080 212
rect 3084 211 3085 215
rect 3215 215 3221 216
rect 3215 214 3216 215
rect 3149 212 3216 214
rect 3079 210 3085 211
rect 3215 211 3216 212
rect 3220 211 3221 215
rect 3215 210 3221 211
rect 3471 215 3477 216
rect 3471 211 3472 215
rect 3476 214 3477 215
rect 3476 212 3505 214
rect 3574 212 3580 213
rect 3476 211 3477 212
rect 3471 210 3477 211
rect 1862 207 1868 208
rect 3574 208 3575 212
rect 3579 208 3580 212
rect 3574 207 3580 208
rect 134 205 140 206
rect 134 201 135 205
rect 139 201 140 205
rect 134 200 140 201
rect 222 205 228 206
rect 222 201 223 205
rect 227 201 228 205
rect 222 200 228 201
rect 310 205 316 206
rect 310 201 311 205
rect 315 201 316 205
rect 310 200 316 201
rect 398 205 404 206
rect 398 201 399 205
rect 403 201 404 205
rect 398 200 404 201
rect 486 205 492 206
rect 486 201 487 205
rect 491 201 492 205
rect 486 200 492 201
rect 574 205 580 206
rect 574 201 575 205
rect 579 201 580 205
rect 574 200 580 201
rect 662 205 668 206
rect 662 201 663 205
rect 667 201 668 205
rect 662 200 668 201
rect 750 205 756 206
rect 750 201 751 205
rect 755 201 756 205
rect 750 200 756 201
rect 838 205 844 206
rect 838 201 839 205
rect 843 201 844 205
rect 838 200 844 201
rect 926 205 932 206
rect 926 201 927 205
rect 931 201 932 205
rect 926 200 932 201
rect 1014 205 1020 206
rect 1014 201 1015 205
rect 1019 201 1020 205
rect 1014 200 1020 201
rect 1102 205 1108 206
rect 1102 201 1103 205
rect 1107 201 1108 205
rect 1102 200 1108 201
rect 1190 205 1196 206
rect 1190 201 1191 205
rect 1195 201 1196 205
rect 1190 200 1196 201
rect 1278 205 1284 206
rect 1278 201 1279 205
rect 1283 201 1284 205
rect 1278 200 1284 201
rect 1366 205 1372 206
rect 1366 201 1367 205
rect 1371 201 1372 205
rect 1366 200 1372 201
rect 1454 205 1460 206
rect 1454 201 1455 205
rect 1459 201 1460 205
rect 1454 200 1460 201
rect 1542 205 1548 206
rect 1542 201 1543 205
rect 1547 201 1548 205
rect 1542 200 1548 201
rect 1630 205 1636 206
rect 1630 201 1631 205
rect 1635 201 1636 205
rect 1630 200 1636 201
rect 1718 205 1724 206
rect 1718 201 1719 205
rect 1723 201 1724 205
rect 1718 200 1724 201
rect 1534 199 1540 200
rect 1534 195 1535 199
rect 1539 198 1540 199
rect 1726 199 1732 200
rect 1726 198 1727 199
rect 1539 196 1727 198
rect 1539 195 1540 196
rect 1534 194 1540 195
rect 1726 195 1727 196
rect 1731 195 1732 199
rect 1726 194 1732 195
rect 1894 199 1900 200
rect 1894 195 1895 199
rect 1899 195 1900 199
rect 1894 194 1900 195
rect 1982 199 1988 200
rect 1982 195 1983 199
rect 1987 195 1988 199
rect 1982 194 1988 195
rect 2070 199 2076 200
rect 2070 195 2071 199
rect 2075 195 2076 199
rect 2070 194 2076 195
rect 2158 199 2164 200
rect 2158 195 2159 199
rect 2163 195 2164 199
rect 2158 194 2164 195
rect 2270 199 2276 200
rect 2270 195 2271 199
rect 2275 195 2276 199
rect 2270 194 2276 195
rect 2406 199 2412 200
rect 2406 195 2407 199
rect 2411 195 2412 199
rect 2406 194 2412 195
rect 2542 199 2548 200
rect 2542 195 2543 199
rect 2547 195 2548 199
rect 2542 194 2548 195
rect 2686 199 2692 200
rect 2686 195 2687 199
rect 2691 195 2692 199
rect 2686 194 2692 195
rect 2822 199 2828 200
rect 2822 195 2823 199
rect 2827 195 2828 199
rect 2822 194 2828 195
rect 2958 199 2964 200
rect 2958 195 2959 199
rect 2963 195 2964 199
rect 2958 194 2964 195
rect 3094 199 3100 200
rect 3094 195 3095 199
rect 3099 195 3100 199
rect 3094 194 3100 195
rect 3230 199 3236 200
rect 3230 195 3231 199
rect 3235 195 3236 199
rect 3230 194 3236 195
rect 3366 199 3372 200
rect 3366 195 3367 199
rect 3371 195 3372 199
rect 3366 194 3372 195
rect 3486 199 3492 200
rect 3486 195 3487 199
rect 3491 195 3492 199
rect 3486 194 3492 195
rect 1887 187 1893 188
rect 1887 183 1888 187
rect 1892 186 1893 187
rect 1902 187 1908 188
rect 1902 186 1903 187
rect 1892 184 1903 186
rect 1892 183 1893 184
rect 1887 182 1893 183
rect 1902 183 1903 184
rect 1907 183 1908 187
rect 1902 182 1908 183
rect 1967 187 1973 188
rect 1967 183 1968 187
rect 1972 186 1973 187
rect 1975 187 1981 188
rect 1975 186 1976 187
rect 1972 184 1976 186
rect 1972 183 1973 184
rect 1967 182 1973 183
rect 1975 183 1976 184
rect 1980 183 1981 187
rect 1975 182 1981 183
rect 2055 187 2061 188
rect 2055 183 2056 187
rect 2060 186 2061 187
rect 2063 187 2069 188
rect 2063 186 2064 187
rect 2060 184 2064 186
rect 2060 183 2061 184
rect 2055 182 2061 183
rect 2063 183 2064 184
rect 2068 183 2069 187
rect 2063 182 2069 183
rect 2143 187 2149 188
rect 2143 183 2144 187
rect 2148 186 2149 187
rect 2151 187 2157 188
rect 2151 186 2152 187
rect 2148 184 2152 186
rect 2148 183 2149 184
rect 2143 182 2149 183
rect 2151 183 2152 184
rect 2156 183 2157 187
rect 2151 182 2157 183
rect 2255 187 2261 188
rect 2255 183 2256 187
rect 2260 186 2261 187
rect 2263 187 2269 188
rect 2263 186 2264 187
rect 2260 184 2264 186
rect 2260 183 2261 184
rect 2255 182 2261 183
rect 2263 183 2264 184
rect 2268 183 2269 187
rect 2263 182 2269 183
rect 2391 187 2397 188
rect 2391 183 2392 187
rect 2396 186 2397 187
rect 2399 187 2405 188
rect 2399 186 2400 187
rect 2396 184 2400 186
rect 2396 183 2397 184
rect 2391 182 2397 183
rect 2399 183 2400 184
rect 2404 183 2405 187
rect 2399 182 2405 183
rect 2527 187 2533 188
rect 2527 183 2528 187
rect 2532 186 2533 187
rect 2535 187 2541 188
rect 2535 186 2536 187
rect 2532 184 2536 186
rect 2532 183 2533 184
rect 2527 182 2533 183
rect 2535 183 2536 184
rect 2540 183 2541 187
rect 2535 182 2541 183
rect 2671 187 2677 188
rect 2671 183 2672 187
rect 2676 186 2677 187
rect 2679 187 2685 188
rect 2679 186 2680 187
rect 2676 184 2680 186
rect 2676 183 2677 184
rect 2671 182 2677 183
rect 2679 183 2680 184
rect 2684 183 2685 187
rect 2679 182 2685 183
rect 2815 187 2821 188
rect 2815 183 2816 187
rect 2820 186 2821 187
rect 2830 187 2836 188
rect 2830 186 2831 187
rect 2820 184 2831 186
rect 2820 183 2821 184
rect 2815 182 2821 183
rect 2830 183 2831 184
rect 2835 183 2836 187
rect 2830 182 2836 183
rect 2943 187 2949 188
rect 2943 183 2944 187
rect 2948 186 2949 187
rect 2951 187 2957 188
rect 2951 186 2952 187
rect 2948 184 2952 186
rect 2948 183 2949 184
rect 2943 182 2949 183
rect 2951 183 2952 184
rect 2956 183 2957 187
rect 2951 182 2957 183
rect 3079 187 3085 188
rect 3079 183 3080 187
rect 3084 186 3085 187
rect 3087 187 3093 188
rect 3087 186 3088 187
rect 3084 184 3088 186
rect 3084 183 3085 184
rect 3079 182 3085 183
rect 3087 183 3088 184
rect 3092 183 3093 187
rect 3087 182 3093 183
rect 3215 187 3221 188
rect 3215 183 3216 187
rect 3220 186 3221 187
rect 3223 187 3229 188
rect 3223 186 3224 187
rect 3220 184 3224 186
rect 3220 183 3221 184
rect 3215 182 3221 183
rect 3223 183 3224 184
rect 3228 183 3229 187
rect 3223 182 3229 183
rect 3359 187 3365 188
rect 3359 183 3360 187
rect 3364 186 3365 187
rect 3374 187 3380 188
rect 3374 186 3375 187
rect 3364 184 3375 186
rect 3364 183 3365 184
rect 3359 182 3365 183
rect 3374 183 3375 184
rect 3379 183 3380 187
rect 3374 182 3380 183
rect 3470 187 3476 188
rect 3470 183 3471 187
rect 3475 186 3476 187
rect 3479 187 3485 188
rect 3479 186 3480 187
rect 3475 184 3480 186
rect 3475 183 3476 184
rect 3470 182 3476 183
rect 3479 183 3480 184
rect 3484 183 3485 187
rect 3479 182 3485 183
rect 2775 143 2781 144
rect 2775 139 2776 143
rect 2780 142 2781 143
rect 2790 143 2796 144
rect 2790 142 2791 143
rect 2780 140 2791 142
rect 2780 139 2781 140
rect 2775 138 2781 139
rect 2790 139 2791 140
rect 2795 139 2796 143
rect 2790 138 2796 139
rect 2847 143 2853 144
rect 2847 139 2848 143
rect 2852 142 2853 143
rect 2863 143 2869 144
rect 2863 142 2864 143
rect 2852 140 2864 142
rect 2852 139 2853 140
rect 2847 138 2853 139
rect 2863 139 2864 140
rect 2868 139 2869 143
rect 2863 138 2869 139
rect 2935 143 2941 144
rect 2935 139 2936 143
rect 2940 142 2941 143
rect 2951 143 2957 144
rect 2951 142 2952 143
rect 2940 140 2952 142
rect 2940 139 2941 140
rect 2935 138 2941 139
rect 2951 139 2952 140
rect 2956 139 2957 143
rect 2951 138 2957 139
rect 3023 143 3029 144
rect 3023 139 3024 143
rect 3028 142 3029 143
rect 3039 143 3045 144
rect 3039 142 3040 143
rect 3028 140 3040 142
rect 3028 139 3029 140
rect 3023 138 3029 139
rect 3039 139 3040 140
rect 3044 139 3045 143
rect 3039 138 3045 139
rect 3111 143 3117 144
rect 3111 139 3112 143
rect 3116 142 3117 143
rect 3127 143 3133 144
rect 3127 142 3128 143
rect 3116 140 3128 142
rect 3116 139 3117 140
rect 3111 138 3117 139
rect 3127 139 3128 140
rect 3132 139 3133 143
rect 3127 138 3133 139
rect 3199 143 3205 144
rect 3199 139 3200 143
rect 3204 142 3205 143
rect 3215 143 3221 144
rect 3215 142 3216 143
rect 3204 140 3216 142
rect 3204 139 3205 140
rect 3199 138 3205 139
rect 3215 139 3216 140
rect 3220 139 3221 143
rect 3215 138 3221 139
rect 3287 143 3293 144
rect 3287 139 3288 143
rect 3292 142 3293 143
rect 3303 143 3309 144
rect 3303 142 3304 143
rect 3292 140 3304 142
rect 3292 139 3293 140
rect 3287 138 3293 139
rect 3303 139 3304 140
rect 3308 139 3309 143
rect 3303 138 3309 139
rect 3391 143 3397 144
rect 3391 139 3392 143
rect 3396 142 3397 143
rect 3458 143 3464 144
rect 3458 142 3459 143
rect 3396 140 3459 142
rect 3396 139 3397 140
rect 3391 138 3397 139
rect 3458 139 3459 140
rect 3463 139 3464 143
rect 3458 138 3464 139
rect 3471 143 3477 144
rect 3471 139 3472 143
rect 3476 142 3477 143
rect 3479 143 3485 144
rect 3479 142 3480 143
rect 3476 140 3480 142
rect 3476 139 3477 140
rect 3471 138 3477 139
rect 3479 139 3480 140
rect 3484 139 3485 143
rect 3479 138 3485 139
rect 2782 133 2788 134
rect 2782 129 2783 133
rect 2787 129 2788 133
rect 2782 128 2788 129
rect 2870 133 2876 134
rect 2870 129 2871 133
rect 2875 129 2876 133
rect 2870 128 2876 129
rect 2958 133 2964 134
rect 2958 129 2959 133
rect 2963 129 2964 133
rect 2958 128 2964 129
rect 3046 133 3052 134
rect 3046 129 3047 133
rect 3051 129 3052 133
rect 3046 128 3052 129
rect 3134 133 3140 134
rect 3134 129 3135 133
rect 3139 129 3140 133
rect 3134 128 3140 129
rect 3222 133 3228 134
rect 3222 129 3223 133
rect 3227 129 3228 133
rect 3222 128 3228 129
rect 3310 133 3316 134
rect 3310 129 3311 133
rect 3315 129 3316 133
rect 3310 128 3316 129
rect 3398 133 3404 134
rect 3398 129 3399 133
rect 3403 129 3404 133
rect 3398 128 3404 129
rect 3486 133 3492 134
rect 3486 129 3487 133
rect 3491 129 3492 133
rect 3486 128 3492 129
rect 1862 120 1868 121
rect 3574 120 3580 121
rect 1862 116 1863 120
rect 1867 116 1868 120
rect 2847 119 2853 120
rect 2847 118 2848 119
rect 2837 116 2848 118
rect 1862 115 1868 116
rect 2847 115 2848 116
rect 2852 115 2853 119
rect 2935 119 2941 120
rect 2935 118 2936 119
rect 2925 116 2936 118
rect 2847 114 2853 115
rect 2935 115 2936 116
rect 2940 115 2941 119
rect 3023 119 3029 120
rect 3023 118 3024 119
rect 3013 116 3024 118
rect 2935 114 2941 115
rect 3023 115 3024 116
rect 3028 115 3029 119
rect 3111 119 3117 120
rect 3111 118 3112 119
rect 3101 116 3112 118
rect 3023 114 3029 115
rect 3111 115 3112 116
rect 3116 115 3117 119
rect 3199 119 3205 120
rect 3199 118 3200 119
rect 3189 116 3200 118
rect 3111 114 3117 115
rect 3199 115 3200 116
rect 3204 115 3205 119
rect 3287 119 3293 120
rect 3287 118 3288 119
rect 3277 116 3288 118
rect 3199 114 3205 115
rect 3287 115 3288 116
rect 3292 115 3293 119
rect 3374 119 3380 120
rect 3374 118 3375 119
rect 3365 116 3375 118
rect 3287 114 3293 115
rect 3374 115 3375 116
rect 3379 115 3380 119
rect 3374 114 3380 115
rect 3458 119 3464 120
rect 3458 115 3459 119
rect 3463 115 3464 119
rect 3574 116 3575 120
rect 3579 116 3580 120
rect 3574 115 3580 116
rect 3458 114 3464 115
rect 3460 112 3505 114
rect 1862 103 1868 104
rect 1862 99 1863 103
rect 1867 99 1868 103
rect 1862 98 1868 99
rect 3574 103 3580 104
rect 3574 99 3575 103
rect 3579 99 3580 103
rect 3574 98 3580 99
rect 2774 93 2780 94
rect 2774 89 2775 93
rect 2779 89 2780 93
rect 2774 88 2780 89
rect 2862 93 2868 94
rect 2862 89 2863 93
rect 2867 89 2868 93
rect 2862 88 2868 89
rect 2950 93 2956 94
rect 2950 89 2951 93
rect 2955 89 2956 93
rect 2950 88 2956 89
rect 3038 93 3044 94
rect 3038 89 3039 93
rect 3043 89 3044 93
rect 3038 88 3044 89
rect 3126 93 3132 94
rect 3126 89 3127 93
rect 3131 89 3132 93
rect 3126 88 3132 89
rect 3214 93 3220 94
rect 3214 89 3215 93
rect 3219 89 3220 93
rect 3214 88 3220 89
rect 3302 93 3308 94
rect 3302 89 3303 93
rect 3307 89 3308 93
rect 3302 88 3308 89
rect 3390 93 3396 94
rect 3390 89 3391 93
rect 3395 89 3396 93
rect 3390 88 3396 89
rect 3478 93 3484 94
rect 3478 89 3479 93
rect 3483 89 3484 93
rect 3478 88 3484 89
<< m3c >>
rect 135 3655 139 3659
rect 223 3655 227 3659
rect 111 3645 115 3649
rect 203 3647 207 3651
rect 1823 3645 1827 3649
rect 111 3628 115 3632
rect 1823 3628 1827 3632
rect 143 3615 147 3619
rect 231 3615 235 3619
rect 199 3591 203 3595
rect 143 3581 147 3585
rect 231 3581 235 3585
rect 319 3581 323 3585
rect 407 3581 411 3585
rect 495 3581 499 3585
rect 1887 3579 1891 3583
rect 1975 3579 1979 3583
rect 2063 3579 2067 3583
rect 2151 3579 2155 3583
rect 2239 3579 2243 3583
rect 2327 3579 2331 3583
rect 2431 3579 2435 3583
rect 2535 3579 2539 3583
rect 2631 3579 2635 3583
rect 2727 3579 2731 3583
rect 2823 3579 2827 3583
rect 2919 3579 2923 3583
rect 3015 3579 3019 3583
rect 3119 3579 3123 3583
rect 3223 3579 3227 3583
rect 111 3568 115 3572
rect 1823 3568 1827 3572
rect 1863 3569 1867 3573
rect 2499 3571 2503 3575
rect 3575 3569 3579 3573
rect 111 3551 115 3555
rect 135 3541 139 3545
rect 223 3541 227 3545
rect 311 3541 315 3545
rect 399 3541 403 3545
rect 267 3535 271 3539
rect 1823 3551 1827 3555
rect 1863 3552 1867 3556
rect 3187 3555 3191 3559
rect 3215 3555 3219 3559
rect 3575 3552 3579 3556
rect 487 3541 491 3545
rect 1895 3539 1899 3543
rect 1983 3539 1987 3543
rect 2071 3539 2075 3543
rect 2159 3539 2163 3543
rect 2247 3539 2251 3543
rect 2335 3539 2339 3543
rect 2439 3539 2443 3543
rect 2543 3539 2547 3543
rect 2639 3539 2643 3543
rect 2735 3539 2739 3543
rect 2831 3539 2835 3543
rect 2927 3539 2931 3543
rect 3023 3539 3027 3543
rect 3127 3539 3131 3543
rect 3231 3539 3235 3543
rect 1887 3527 1888 3531
rect 1888 3527 1891 3531
rect 3187 3527 3191 3531
rect 247 3519 251 3523
rect 375 3519 379 3523
rect 503 3519 507 3523
rect 623 3519 627 3523
rect 743 3519 747 3523
rect 863 3519 867 3523
rect 975 3519 979 3523
rect 1079 3519 1083 3523
rect 1175 3519 1179 3523
rect 1271 3519 1275 3523
rect 1367 3519 1371 3523
rect 1471 3519 1475 3523
rect 1575 3519 1579 3523
rect 111 3509 115 3513
rect 1539 3511 1543 3515
rect 1963 3515 1967 3519
rect 1991 3515 1995 3519
rect 2111 3515 2115 3519
rect 2291 3515 2295 3519
rect 2723 3515 2727 3519
rect 2799 3515 2803 3519
rect 3003 3515 3007 3519
rect 3183 3515 3187 3519
rect 3215 3515 3216 3519
rect 3216 3515 3219 3519
rect 1823 3509 1827 3513
rect 1895 3505 1899 3509
rect 1983 3505 1987 3509
rect 2103 3505 2107 3509
rect 2231 3505 2235 3509
rect 2367 3505 2371 3509
rect 2511 3505 2515 3509
rect 2655 3505 2659 3509
rect 2791 3505 2795 3509
rect 2935 3505 2939 3509
rect 3079 3505 3083 3509
rect 3223 3505 3227 3509
rect 111 3492 115 3496
rect 571 3495 575 3499
rect 735 3495 739 3499
rect 967 3495 971 3499
rect 1823 3492 1827 3496
rect 1863 3492 1867 3496
rect 1887 3487 1891 3491
rect 1963 3487 1967 3491
rect 2291 3491 2295 3495
rect 3575 3492 3579 3496
rect 2723 3487 2727 3491
rect 3003 3487 3007 3491
rect 3183 3487 3187 3491
rect 255 3479 259 3483
rect 383 3479 387 3483
rect 511 3479 515 3483
rect 631 3479 635 3483
rect 751 3479 755 3483
rect 871 3479 875 3483
rect 983 3479 987 3483
rect 1087 3479 1091 3483
rect 1183 3479 1187 3483
rect 1279 3479 1283 3483
rect 1375 3479 1379 3483
rect 1479 3479 1483 3483
rect 1583 3479 1587 3483
rect 267 3467 271 3471
rect 571 3471 575 3475
rect 1863 3475 1867 3479
rect 2887 3475 2891 3479
rect 3575 3475 3579 3479
rect 967 3467 971 3471
rect 1887 3465 1891 3469
rect 1975 3465 1979 3469
rect 2095 3465 2099 3469
rect 2223 3465 2227 3469
rect 2359 3465 2363 3469
rect 2503 3465 2507 3469
rect 2647 3465 2651 3469
rect 2783 3465 2787 3469
rect 2927 3465 2931 3469
rect 3071 3465 3075 3469
rect 3215 3465 3219 3469
rect 243 3455 247 3459
rect 371 3455 375 3459
rect 651 3459 655 3463
rect 683 3451 687 3455
rect 735 3455 736 3459
rect 736 3455 739 3459
rect 963 3455 967 3459
rect 1251 3455 1255 3459
rect 1439 3455 1443 3459
rect 1539 3455 1543 3459
rect 175 3445 179 3449
rect 303 3445 307 3449
rect 447 3445 451 3449
rect 591 3445 595 3449
rect 743 3445 747 3449
rect 895 3445 899 3449
rect 1039 3445 1043 3449
rect 1183 3445 1187 3449
rect 1327 3445 1331 3449
rect 1479 3445 1483 3449
rect 111 3432 115 3436
rect 243 3427 247 3431
rect 371 3427 375 3431
rect 651 3431 655 3435
rect 1823 3432 1827 3436
rect 1887 3435 1891 3439
rect 2023 3435 2027 3439
rect 2191 3435 2195 3439
rect 2367 3435 2371 3439
rect 2543 3435 2547 3439
rect 2711 3435 2715 3439
rect 2871 3435 2875 3439
rect 3031 3435 3035 3439
rect 3191 3435 3195 3439
rect 3359 3435 3363 3439
rect 683 3427 687 3431
rect 963 3427 967 3431
rect 1251 3427 1255 3431
rect 1471 3427 1475 3431
rect 1863 3425 1867 3429
rect 1991 3427 1995 3431
rect 2799 3427 2803 3431
rect 3259 3427 3263 3431
rect 3575 3425 3579 3429
rect 111 3415 115 3419
rect 151 3415 155 3419
rect 1823 3415 1827 3419
rect 167 3405 171 3409
rect 295 3405 299 3409
rect 439 3405 443 3409
rect 583 3405 587 3409
rect 735 3405 739 3409
rect 887 3405 891 3409
rect 1031 3405 1035 3409
rect 1175 3405 1179 3409
rect 1319 3405 1323 3409
rect 1471 3405 1475 3409
rect 1863 3408 1867 3412
rect 2091 3411 2095 3415
rect 2259 3411 2263 3415
rect 2435 3411 2439 3415
rect 3575 3408 3579 3412
rect 1223 3399 1224 3403
rect 1224 3399 1227 3403
rect 1895 3395 1899 3399
rect 2031 3395 2035 3399
rect 2199 3395 2203 3399
rect 2375 3395 2379 3399
rect 2551 3395 2555 3399
rect 2719 3395 2723 3399
rect 2879 3395 2883 3399
rect 3039 3395 3043 3399
rect 3199 3395 3203 3399
rect 3367 3395 3371 3399
rect 135 3383 139 3387
rect 263 3383 267 3387
rect 407 3383 411 3387
rect 567 3383 571 3387
rect 727 3383 731 3387
rect 887 3383 891 3387
rect 1047 3383 1051 3387
rect 1207 3383 1211 3387
rect 1367 3383 1371 3387
rect 1527 3383 1531 3387
rect 1887 3383 1888 3387
rect 1888 3383 1891 3387
rect 2259 3383 2263 3387
rect 2435 3383 2439 3387
rect 2711 3383 2712 3387
rect 2712 3383 2715 3387
rect 2887 3383 2891 3387
rect 111 3373 115 3377
rect 683 3375 687 3379
rect 1823 3373 1827 3377
rect 111 3356 115 3360
rect 2091 3363 2095 3367
rect 2887 3363 2891 3367
rect 3047 3363 3051 3367
rect 1823 3356 1827 3360
rect 1895 3353 1899 3357
rect 2031 3353 2035 3357
rect 2199 3353 2203 3357
rect 2375 3353 2379 3357
rect 2551 3353 2555 3357
rect 2719 3353 2723 3357
rect 2879 3353 2883 3357
rect 3039 3353 3043 3357
rect 3191 3353 3195 3357
rect 3343 3353 3347 3357
rect 3487 3353 3491 3357
rect 143 3343 147 3347
rect 271 3343 275 3347
rect 415 3343 419 3347
rect 575 3343 579 3347
rect 735 3343 739 3347
rect 895 3343 899 3347
rect 1055 3343 1059 3347
rect 1215 3343 1219 3347
rect 1375 3343 1379 3347
rect 1535 3343 1539 3347
rect 1863 3340 1867 3344
rect 151 3331 155 3335
rect 1223 3331 1227 3335
rect 1887 3335 1891 3339
rect 2711 3335 2715 3339
rect 3575 3340 3579 3344
rect 1863 3323 1867 3327
rect 2479 3323 2483 3327
rect 3411 3323 3415 3327
rect 3575 3323 3579 3327
rect 215 3315 219 3319
rect 1079 3315 1083 3319
rect 1175 3315 1179 3319
rect 1427 3315 1431 3319
rect 1887 3313 1891 3317
rect 2023 3313 2027 3317
rect 2191 3313 2195 3317
rect 2367 3313 2371 3317
rect 2543 3313 2547 3317
rect 2711 3313 2715 3317
rect 2871 3313 2875 3317
rect 3031 3313 3035 3317
rect 3183 3313 3187 3317
rect 3335 3313 3339 3317
rect 3479 3313 3483 3317
rect 207 3305 211 3309
rect 335 3305 339 3309
rect 479 3305 483 3309
rect 639 3305 643 3309
rect 807 3305 811 3309
rect 983 3305 987 3309
rect 1167 3305 1171 3309
rect 1351 3305 1355 3309
rect 1543 3305 1547 3309
rect 111 3292 115 3296
rect 1823 3292 1827 3296
rect 1079 3287 1083 3291
rect 1887 3291 1891 3295
rect 1427 3287 1431 3291
rect 2007 3291 2011 3295
rect 2151 3291 2155 3295
rect 2303 3291 2307 3295
rect 2463 3291 2467 3295
rect 2631 3291 2635 3295
rect 2799 3291 2803 3295
rect 2967 3291 2971 3295
rect 3135 3291 3139 3295
rect 3311 3291 3315 3295
rect 3479 3291 3483 3295
rect 1863 3281 1867 3285
rect 2539 3283 2543 3287
rect 2887 3283 2891 3287
rect 111 3275 115 3279
rect 199 3265 203 3269
rect 327 3265 331 3269
rect 471 3265 475 3269
rect 631 3265 635 3269
rect 1823 3275 1827 3279
rect 3479 3279 3483 3283
rect 3575 3281 3579 3285
rect 799 3265 803 3269
rect 975 3265 979 3269
rect 1159 3265 1163 3269
rect 1343 3265 1347 3269
rect 1535 3265 1539 3269
rect 1863 3264 1867 3268
rect 1955 3267 1959 3271
rect 2235 3267 2239 3271
rect 2867 3267 2871 3271
rect 3055 3267 3059 3271
rect 3575 3264 3579 3268
rect 1895 3251 1899 3255
rect 2015 3251 2019 3255
rect 2159 3251 2163 3255
rect 2311 3251 2315 3255
rect 2471 3251 2475 3255
rect 2639 3251 2643 3255
rect 2807 3251 2811 3255
rect 2975 3251 2979 3255
rect 3143 3251 3147 3255
rect 3319 3251 3323 3255
rect 3487 3251 3491 3255
rect 367 3239 371 3243
rect 503 3239 507 3243
rect 639 3239 643 3243
rect 783 3239 787 3243
rect 935 3239 939 3243
rect 1095 3239 1099 3243
rect 1255 3239 1259 3243
rect 1415 3239 1419 3243
rect 1575 3239 1579 3243
rect 1951 3239 1955 3243
rect 1959 3239 1963 3243
rect 2167 3239 2171 3243
rect 2235 3239 2239 3243
rect 2867 3239 2871 3243
rect 3055 3239 3059 3243
rect 3259 3239 3263 3243
rect 3411 3239 3415 3243
rect 111 3229 115 3233
rect 711 3231 715 3235
rect 1175 3231 1179 3235
rect 1823 3229 1827 3233
rect 111 3212 115 3216
rect 1163 3215 1167 3219
rect 1647 3215 1651 3219
rect 1967 3219 1971 3223
rect 2031 3219 2035 3223
rect 2183 3219 2187 3223
rect 2243 3219 2247 3223
rect 2399 3219 2403 3223
rect 2527 3219 2531 3223
rect 2791 3219 2795 3223
rect 2943 3219 2947 3223
rect 3083 3219 3087 3223
rect 3251 3219 3255 3223
rect 3479 3219 3480 3223
rect 3480 3219 3483 3223
rect 1823 3212 1827 3216
rect 1895 3209 1899 3213
rect 2023 3209 2027 3213
rect 2175 3209 2179 3213
rect 2327 3209 2331 3213
rect 2463 3209 2467 3213
rect 2599 3209 2603 3213
rect 2735 3209 2739 3213
rect 2871 3209 2875 3213
rect 3015 3209 3019 3213
rect 3167 3209 3171 3213
rect 3327 3209 3331 3213
rect 3487 3209 3491 3213
rect 375 3199 379 3203
rect 511 3199 515 3203
rect 647 3199 651 3203
rect 791 3199 795 3203
rect 943 3199 947 3203
rect 1103 3199 1107 3203
rect 1263 3199 1267 3203
rect 1423 3199 1427 3203
rect 1583 3199 1587 3203
rect 1863 3196 1867 3200
rect 1959 3195 1963 3199
rect 951 3187 955 3191
rect 1967 3191 1971 3195
rect 2243 3195 2247 3199
rect 2399 3195 2403 3199
rect 2527 3195 2531 3199
rect 2943 3195 2947 3199
rect 3083 3195 3087 3199
rect 3251 3195 3255 3199
rect 3575 3196 3579 3200
rect 3259 3191 3263 3195
rect 1863 3179 1867 3183
rect 2531 3179 2535 3183
rect 3575 3179 3579 3183
rect 487 3167 491 3171
rect 1367 3167 1371 3171
rect 1539 3167 1543 3171
rect 1647 3167 1651 3171
rect 1887 3169 1891 3173
rect 2015 3169 2019 3173
rect 2167 3169 2171 3173
rect 2319 3169 2323 3173
rect 2455 3169 2459 3173
rect 2591 3169 2595 3173
rect 2727 3169 2731 3173
rect 2863 3169 2867 3173
rect 3007 3169 3011 3173
rect 3159 3169 3163 3173
rect 3319 3169 3323 3173
rect 3479 3169 3483 3173
rect 447 3157 451 3161
rect 559 3157 563 3161
rect 687 3157 691 3161
rect 823 3157 827 3161
rect 975 3157 979 3161
rect 1135 3157 1139 3161
rect 1295 3157 1299 3161
rect 1463 3157 1467 3161
rect 1639 3157 1643 3161
rect 111 3144 115 3148
rect 1823 3144 1827 3148
rect 1887 3143 1891 3147
rect 1539 3139 1543 3143
rect 2047 3143 2051 3147
rect 2199 3143 2203 3147
rect 2351 3143 2355 3147
rect 2511 3143 2515 3147
rect 2679 3143 2683 3147
rect 2871 3143 2875 3147
rect 3071 3143 3075 3147
rect 3287 3143 3291 3147
rect 3479 3143 3483 3147
rect 1863 3133 1867 3137
rect 2031 3135 2035 3139
rect 2791 3135 2795 3139
rect 3575 3133 3579 3137
rect 111 3127 115 3131
rect 891 3127 895 3131
rect 1823 3127 1827 3131
rect 439 3117 443 3121
rect 551 3117 555 3121
rect 679 3117 683 3121
rect 815 3117 819 3121
rect 967 3117 971 3121
rect 1127 3117 1131 3121
rect 1287 3117 1291 3121
rect 1455 3117 1459 3121
rect 1631 3117 1635 3121
rect 1863 3116 1867 3120
rect 2747 3119 2751 3123
rect 2939 3119 2943 3123
rect 3471 3119 3475 3123
rect 3575 3116 3579 3120
rect 1895 3103 1899 3107
rect 2055 3103 2059 3107
rect 2207 3103 2211 3107
rect 2359 3103 2363 3107
rect 2519 3103 2523 3107
rect 2687 3103 2691 3107
rect 2879 3103 2883 3107
rect 3079 3103 3083 3107
rect 3295 3103 3299 3107
rect 3487 3103 3491 3107
rect 551 3087 555 3091
rect 663 3087 667 3091
rect 783 3087 787 3091
rect 903 3087 907 3091
rect 1031 3087 1035 3091
rect 1159 3087 1163 3091
rect 1287 3087 1291 3091
rect 1423 3087 1427 3091
rect 1559 3087 1563 3091
rect 1695 3087 1699 3091
rect 2215 3091 2219 3095
rect 2939 3091 2943 3095
rect 3303 3091 3307 3095
rect 111 3077 115 3081
rect 1367 3079 1371 3083
rect 1823 3077 1827 3081
rect 2007 3071 2011 3075
rect 2183 3071 2187 3075
rect 2503 3071 2507 3075
rect 2747 3071 2751 3075
rect 3247 3071 3251 3075
rect 3471 3071 3475 3075
rect 111 3060 115 3064
rect 1763 3063 1767 3067
rect 1823 3060 1827 3064
rect 1919 3061 1923 3065
rect 2087 3061 2091 3065
rect 2279 3061 2283 3065
rect 2487 3061 2491 3065
rect 2719 3061 2723 3065
rect 2975 3061 2979 3065
rect 3239 3061 3243 3065
rect 3487 3061 3491 3065
rect 559 3047 563 3051
rect 671 3047 675 3051
rect 791 3047 795 3051
rect 911 3047 915 3051
rect 1039 3047 1043 3051
rect 1167 3047 1171 3051
rect 1295 3047 1299 3051
rect 1431 3047 1435 3051
rect 1567 3047 1571 3051
rect 1703 3047 1707 3051
rect 1863 3048 1867 3052
rect 2007 3043 2011 3047
rect 2183 3043 2187 3047
rect 2899 3043 2903 3047
rect 3303 3047 3307 3051
rect 3575 3048 3579 3052
rect 567 3035 571 3039
rect 1175 3035 1179 3039
rect 1863 3031 1867 3035
rect 2431 3031 2435 3035
rect 3575 3031 3579 3035
rect 771 3019 775 3023
rect 899 3019 903 3023
rect 1307 3019 1311 3023
rect 1439 3019 1443 3023
rect 1595 3019 1599 3023
rect 1763 3019 1767 3023
rect 1911 3021 1915 3025
rect 2079 3021 2083 3025
rect 2271 3021 2275 3025
rect 2479 3021 2483 3025
rect 2711 3021 2715 3025
rect 2967 3021 2971 3025
rect 3231 3021 3235 3025
rect 3479 3021 3483 3025
rect 575 3009 579 3013
rect 703 3009 707 3013
rect 831 3009 835 3013
rect 967 3009 971 3013
rect 1103 3009 1107 3013
rect 1239 3009 1243 3013
rect 1367 3009 1371 3013
rect 1495 3009 1499 3013
rect 1623 3009 1627 3013
rect 1735 3009 1739 3013
rect 111 2996 115 3000
rect 1823 2996 1827 3000
rect 771 2991 775 2995
rect 899 2991 903 2995
rect 1175 2991 1179 2995
rect 1307 2991 1311 2995
rect 1439 2991 1443 2995
rect 2023 2995 2027 2999
rect 2159 2995 2163 2999
rect 2287 2995 2291 2999
rect 2415 2995 2419 2999
rect 2535 2995 2539 2999
rect 2663 2995 2667 2999
rect 2807 2995 2811 2999
rect 2967 2995 2971 2999
rect 3143 2995 3147 2999
rect 3319 2995 3323 2999
rect 3479 2995 3483 2999
rect 1863 2985 1867 2989
rect 3247 2987 3251 2991
rect 3575 2985 3579 2989
rect 111 2979 115 2983
rect 511 2979 515 2983
rect 1691 2979 1695 2983
rect 1823 2979 1827 2983
rect 567 2969 571 2973
rect 695 2969 699 2973
rect 823 2969 827 2973
rect 959 2969 963 2973
rect 1095 2969 1099 2973
rect 1231 2969 1235 2973
rect 1359 2969 1363 2973
rect 1487 2969 1491 2973
rect 1615 2969 1619 2973
rect 1727 2969 1731 2973
rect 1863 2968 1867 2972
rect 3471 2971 3475 2975
rect 3575 2968 3579 2972
rect 2031 2955 2035 2959
rect 2167 2955 2171 2959
rect 2295 2955 2299 2959
rect 2423 2955 2427 2959
rect 2543 2955 2547 2959
rect 2671 2955 2675 2959
rect 2815 2955 2819 2959
rect 2975 2955 2979 2959
rect 3151 2955 3155 2959
rect 3327 2955 3331 2959
rect 3487 2955 3491 2959
rect 495 2947 499 2951
rect 639 2947 643 2951
rect 783 2947 787 2951
rect 919 2947 923 2951
rect 1055 2947 1059 2951
rect 1183 2947 1187 2951
rect 1303 2947 1307 2951
rect 1415 2947 1419 2951
rect 1527 2947 1531 2951
rect 1639 2947 1643 2951
rect 1727 2947 1731 2951
rect 111 2937 115 2941
rect 1595 2939 1599 2943
rect 2431 2943 2435 2947
rect 1823 2937 1827 2941
rect 111 2920 115 2924
rect 631 2923 635 2927
rect 1823 2920 1827 2924
rect 2319 2923 2323 2927
rect 2563 2923 2567 2927
rect 3471 2923 3475 2927
rect 1895 2913 1899 2917
rect 2175 2913 2179 2917
rect 2495 2913 2499 2917
rect 2823 2913 2827 2917
rect 3167 2913 3171 2917
rect 3487 2913 3491 2917
rect 503 2907 507 2911
rect 647 2907 651 2911
rect 791 2907 795 2911
rect 927 2907 931 2911
rect 1063 2907 1067 2911
rect 1191 2907 1195 2911
rect 1311 2907 1315 2911
rect 1423 2907 1427 2911
rect 1535 2907 1539 2911
rect 1647 2907 1651 2911
rect 1735 2907 1739 2911
rect 1863 2900 1867 2904
rect 3575 2900 3579 2904
rect 511 2895 515 2899
rect 631 2895 635 2899
rect 1167 2895 1171 2899
rect 1691 2895 1695 2899
rect 2319 2895 2323 2899
rect 2563 2895 2567 2899
rect 395 2879 399 2883
rect 523 2879 527 2883
rect 671 2879 675 2883
rect 799 2879 803 2883
rect 1015 2879 1019 2883
rect 1503 2879 1507 2883
rect 1863 2883 1867 2887
rect 3071 2883 3075 2887
rect 3575 2883 3579 2887
rect 327 2869 331 2873
rect 455 2869 459 2873
rect 591 2869 595 2873
rect 727 2869 731 2873
rect 871 2869 875 2873
rect 1007 2869 1011 2873
rect 1143 2869 1147 2873
rect 1279 2869 1283 2873
rect 1415 2869 1419 2873
rect 1551 2869 1555 2873
rect 1887 2873 1891 2877
rect 2167 2873 2171 2877
rect 2487 2873 2491 2877
rect 2815 2873 2819 2877
rect 3159 2873 3163 2877
rect 3479 2873 3483 2877
rect 111 2856 115 2860
rect 395 2851 399 2855
rect 523 2851 527 2855
rect 671 2851 675 2855
rect 799 2851 803 2855
rect 1503 2855 1507 2859
rect 1823 2856 1827 2860
rect 2687 2859 2691 2863
rect 1511 2851 1515 2855
rect 1887 2851 1891 2855
rect 2023 2851 2027 2855
rect 2191 2851 2195 2855
rect 2359 2851 2363 2855
rect 2519 2851 2523 2855
rect 2671 2851 2675 2855
rect 2807 2851 2811 2855
rect 2935 2851 2939 2855
rect 111 2839 115 2843
rect 1823 2839 1827 2843
rect 1863 2841 1867 2845
rect 3055 2851 3059 2855
rect 3167 2851 3171 2855
rect 3279 2851 3283 2855
rect 3391 2851 3395 2855
rect 3479 2851 3483 2855
rect 3575 2841 3579 2845
rect 319 2829 323 2833
rect 447 2829 451 2833
rect 583 2829 587 2833
rect 719 2829 723 2833
rect 863 2829 867 2833
rect 999 2829 1003 2833
rect 1135 2829 1139 2833
rect 1271 2829 1275 2833
rect 1407 2829 1411 2833
rect 1543 2829 1547 2833
rect 1863 2824 1867 2828
rect 2091 2827 2095 2831
rect 3235 2827 3239 2831
rect 3347 2827 3351 2831
rect 3471 2827 3475 2831
rect 3575 2824 3579 2828
rect 1015 2807 1019 2811
rect 1895 2811 1899 2815
rect 2031 2811 2035 2815
rect 2199 2811 2203 2815
rect 2367 2811 2371 2815
rect 2527 2811 2531 2815
rect 2679 2811 2683 2815
rect 2815 2811 2819 2815
rect 2943 2811 2947 2815
rect 3063 2811 3067 2815
rect 3175 2811 3179 2815
rect 3287 2811 3291 2815
rect 3399 2811 3403 2815
rect 3487 2811 3491 2815
rect 167 2799 171 2803
rect 295 2799 299 2803
rect 423 2799 427 2803
rect 559 2799 563 2803
rect 695 2799 699 2803
rect 823 2799 827 2803
rect 951 2799 955 2803
rect 1079 2799 1083 2803
rect 1207 2799 1211 2803
rect 1343 2799 1347 2803
rect 2687 2799 2691 2803
rect 3071 2799 3075 2803
rect 3235 2799 3239 2803
rect 3347 2799 3351 2803
rect 3427 2799 3431 2803
rect 111 2789 115 2793
rect 1823 2789 1827 2793
rect 2091 2787 2095 2791
rect 2339 2787 2343 2791
rect 2507 2787 2511 2791
rect 2563 2787 2567 2791
rect 2847 2787 2851 2791
rect 3435 2787 3439 2791
rect 3471 2787 3475 2791
rect 111 2772 115 2776
rect 363 2775 367 2779
rect 627 2775 631 2779
rect 647 2775 651 2779
rect 1895 2777 1899 2781
rect 2063 2777 2067 2781
rect 2255 2777 2259 2781
rect 2439 2777 2443 2781
rect 2615 2777 2619 2781
rect 2783 2777 2787 2781
rect 2935 2777 2939 2781
rect 3079 2777 3083 2781
rect 3223 2777 3227 2781
rect 3367 2777 3371 2781
rect 3487 2777 3491 2781
rect 1823 2772 1827 2776
rect 1863 2764 1867 2768
rect 175 2759 179 2763
rect 303 2759 307 2763
rect 431 2759 435 2763
rect 567 2759 571 2763
rect 703 2759 707 2763
rect 831 2759 835 2763
rect 959 2759 963 2763
rect 1087 2759 1091 2763
rect 1215 2759 1219 2763
rect 1351 2759 1355 2763
rect 2339 2759 2343 2763
rect 2507 2759 2511 2763
rect 3427 2763 3431 2767
rect 3575 2764 3579 2768
rect 3435 2759 3439 2763
rect 183 2747 187 2751
rect 627 2747 631 2751
rect 1863 2747 1867 2751
rect 3575 2747 3579 2751
rect 211 2727 215 2731
rect 1887 2737 1891 2741
rect 2055 2737 2059 2741
rect 2247 2737 2251 2741
rect 2431 2737 2435 2741
rect 2607 2737 2611 2741
rect 2775 2737 2779 2741
rect 2927 2737 2931 2741
rect 3071 2737 3075 2741
rect 3215 2737 3219 2741
rect 3359 2737 3363 2741
rect 3479 2737 3483 2741
rect 363 2727 367 2731
rect 2975 2731 2976 2735
rect 2976 2731 2979 2735
rect 2847 2723 2851 2727
rect 143 2717 147 2721
rect 231 2717 235 2721
rect 351 2717 355 2721
rect 479 2717 483 2721
rect 615 2717 619 2721
rect 759 2717 763 2721
rect 903 2717 907 2721
rect 1047 2717 1051 2721
rect 1887 2711 1891 2715
rect 2047 2711 2051 2715
rect 2207 2711 2211 2715
rect 2359 2711 2363 2715
rect 2495 2711 2499 2715
rect 2623 2711 2627 2715
rect 2743 2711 2747 2715
rect 2863 2711 2867 2715
rect 2983 2711 2987 2715
rect 3103 2711 3107 2715
rect 111 2704 115 2708
rect 211 2699 215 2703
rect 1823 2704 1827 2708
rect 1863 2701 1867 2705
rect 2563 2703 2567 2707
rect 3051 2703 3055 2707
rect 3575 2701 3579 2705
rect 111 2687 115 2691
rect 1823 2687 1827 2691
rect 1863 2684 1867 2688
rect 1955 2687 1959 2691
rect 2691 2687 2695 2691
rect 2699 2687 2703 2691
rect 2811 2687 2815 2691
rect 3575 2684 3579 2688
rect 135 2677 139 2681
rect 223 2677 227 2681
rect 343 2677 347 2681
rect 471 2677 475 2681
rect 607 2677 611 2681
rect 751 2677 755 2681
rect 895 2677 899 2681
rect 1039 2677 1043 2681
rect 1895 2671 1899 2675
rect 2055 2671 2059 2675
rect 2215 2671 2219 2675
rect 2367 2671 2371 2675
rect 2503 2671 2507 2675
rect 2631 2671 2635 2675
rect 2751 2671 2755 2675
rect 2871 2671 2875 2675
rect 2991 2671 2995 2675
rect 3111 2671 3115 2675
rect 1955 2659 1959 2663
rect 2327 2659 2331 2663
rect 2699 2659 2703 2663
rect 2811 2659 2815 2663
rect 135 2651 139 2655
rect 231 2651 235 2655
rect 351 2651 355 2655
rect 471 2651 475 2655
rect 583 2651 587 2655
rect 695 2651 699 2655
rect 799 2651 803 2655
rect 903 2651 907 2655
rect 999 2651 1003 2655
rect 1103 2651 1107 2655
rect 1207 2651 1211 2655
rect 1311 2651 1315 2655
rect 2975 2659 2979 2663
rect 111 2641 115 2645
rect 423 2643 427 2647
rect 1275 2643 1279 2647
rect 1823 2641 1827 2645
rect 2315 2639 2319 2643
rect 2523 2639 2527 2643
rect 3051 2651 3055 2655
rect 2691 2639 2695 2643
rect 111 2624 115 2628
rect 1895 2629 1899 2633
rect 1999 2629 2003 2633
rect 2119 2629 2123 2633
rect 2239 2629 2243 2633
rect 2351 2629 2355 2633
rect 2455 2629 2459 2633
rect 2551 2629 2555 2633
rect 2655 2629 2659 2633
rect 2759 2629 2763 2633
rect 2863 2629 2867 2633
rect 1823 2624 1827 2628
rect 1863 2616 1867 2620
rect 143 2611 147 2615
rect 239 2611 243 2615
rect 359 2611 363 2615
rect 479 2611 483 2615
rect 591 2611 595 2615
rect 703 2611 707 2615
rect 807 2611 811 2615
rect 911 2611 915 2615
rect 1007 2611 1011 2615
rect 1111 2611 1115 2615
rect 1215 2611 1219 2615
rect 1319 2611 1323 2615
rect 2315 2615 2319 2619
rect 2327 2611 2331 2615
rect 2523 2611 2527 2615
rect 3575 2616 3579 2620
rect 619 2599 623 2603
rect 747 2599 751 2603
rect 1863 2599 1867 2603
rect 3575 2599 3579 2603
rect 1887 2589 1891 2593
rect 1991 2589 1995 2593
rect 2111 2589 2115 2593
rect 2231 2589 2235 2593
rect 2343 2589 2347 2593
rect 2447 2589 2451 2593
rect 2543 2589 2547 2593
rect 2647 2589 2651 2593
rect 2751 2589 2755 2593
rect 2855 2589 2859 2593
rect 211 2583 215 2587
rect 339 2583 343 2587
rect 423 2583 427 2587
rect 651 2583 655 2587
rect 663 2583 667 2587
rect 815 2583 819 2587
rect 995 2583 999 2587
rect 1119 2583 1123 2587
rect 1275 2583 1279 2587
rect 2487 2583 2491 2587
rect 143 2573 147 2577
rect 271 2573 275 2577
rect 415 2573 419 2577
rect 551 2573 555 2577
rect 679 2573 683 2577
rect 807 2573 811 2577
rect 927 2573 931 2577
rect 1047 2573 1051 2577
rect 1175 2573 1179 2577
rect 111 2560 115 2564
rect 211 2555 215 2559
rect 339 2555 343 2559
rect 619 2559 623 2563
rect 1823 2560 1827 2564
rect 1887 2563 1891 2567
rect 1991 2563 1995 2567
rect 2111 2563 2115 2567
rect 2231 2563 2235 2567
rect 2351 2563 2355 2567
rect 2471 2563 2475 2567
rect 2591 2563 2595 2567
rect 2711 2563 2715 2567
rect 2831 2563 2835 2567
rect 651 2555 655 2559
rect 747 2555 751 2559
rect 995 2555 999 2559
rect 1119 2555 1123 2559
rect 1863 2553 1867 2557
rect 2779 2555 2783 2559
rect 3575 2553 3579 2557
rect 111 2543 115 2547
rect 887 2543 891 2547
rect 1823 2543 1827 2547
rect 135 2533 139 2537
rect 263 2533 267 2537
rect 407 2533 411 2537
rect 543 2533 547 2537
rect 671 2533 675 2537
rect 799 2533 803 2537
rect 919 2533 923 2537
rect 1039 2533 1043 2537
rect 1167 2533 1171 2537
rect 1863 2536 1867 2540
rect 1955 2539 1959 2543
rect 2179 2539 2183 2543
rect 2327 2539 2331 2543
rect 3575 2536 3579 2540
rect 1895 2523 1899 2527
rect 1999 2523 2003 2527
rect 2119 2523 2123 2527
rect 2239 2523 2243 2527
rect 2359 2523 2363 2527
rect 2479 2523 2483 2527
rect 2599 2523 2603 2527
rect 2719 2523 2723 2527
rect 2839 2523 2843 2527
rect 135 2511 139 2515
rect 279 2511 283 2515
rect 439 2511 443 2515
rect 591 2511 595 2515
rect 735 2511 739 2515
rect 871 2511 875 2515
rect 1007 2511 1011 2515
rect 1143 2511 1147 2515
rect 1279 2511 1283 2515
rect 1955 2511 1959 2515
rect 2179 2511 2183 2515
rect 2327 2511 2331 2515
rect 2335 2511 2339 2515
rect 2487 2511 2491 2515
rect 111 2501 115 2505
rect 663 2503 667 2507
rect 815 2503 819 2507
rect 1219 2503 1223 2507
rect 1823 2501 1827 2505
rect 2495 2495 2499 2499
rect 111 2484 115 2488
rect 1823 2484 1827 2488
rect 1895 2485 1899 2489
rect 2031 2485 2035 2489
rect 2191 2485 2195 2489
rect 2343 2485 2347 2489
rect 2487 2485 2491 2489
rect 2623 2485 2627 2489
rect 2751 2485 2755 2489
rect 2879 2485 2883 2489
rect 3015 2485 3019 2489
rect 143 2471 147 2475
rect 287 2471 291 2475
rect 447 2471 451 2475
rect 599 2471 603 2475
rect 743 2471 747 2475
rect 879 2471 883 2475
rect 1015 2471 1019 2475
rect 1151 2471 1155 2475
rect 1287 2471 1291 2475
rect 1863 2472 1867 2476
rect 2335 2467 2339 2471
rect 3575 2472 3579 2476
rect 583 2459 587 2463
rect 795 2459 799 2463
rect 887 2459 891 2463
rect 1863 2455 1867 2459
rect 2031 2455 2035 2459
rect 2967 2455 2971 2459
rect 3575 2455 3579 2459
rect 259 2447 263 2451
rect 391 2447 395 2451
rect 679 2447 683 2451
rect 767 2447 771 2451
rect 887 2447 891 2451
rect 1007 2447 1011 2451
rect 1887 2445 1891 2449
rect 2023 2445 2027 2449
rect 2183 2445 2187 2449
rect 2335 2445 2339 2449
rect 2479 2445 2483 2449
rect 2615 2445 2619 2449
rect 2743 2445 2747 2449
rect 2871 2445 2875 2449
rect 3007 2445 3011 2449
rect 191 2437 195 2441
rect 319 2437 323 2441
rect 455 2437 459 2441
rect 591 2437 595 2441
rect 727 2437 731 2441
rect 863 2437 867 2441
rect 999 2437 1003 2441
rect 1135 2437 1139 2441
rect 1271 2437 1275 2441
rect 1407 2437 1411 2441
rect 111 2424 115 2428
rect 259 2419 263 2423
rect 391 2419 395 2423
rect 583 2419 587 2423
rect 679 2419 683 2423
rect 795 2419 799 2423
rect 1823 2424 1827 2428
rect 1887 2423 1891 2427
rect 2015 2423 2019 2427
rect 2175 2423 2179 2427
rect 2335 2423 2339 2427
rect 2495 2423 2499 2427
rect 2647 2423 2651 2427
rect 2799 2423 2803 2427
rect 2951 2423 2955 2427
rect 3111 2423 3115 2427
rect 1863 2413 1867 2417
rect 3019 2415 3023 2419
rect 3575 2413 3579 2417
rect 111 2407 115 2411
rect 175 2407 179 2411
rect 1339 2407 1343 2411
rect 1823 2407 1827 2411
rect 183 2397 187 2401
rect 311 2397 315 2401
rect 447 2397 451 2401
rect 583 2397 587 2401
rect 719 2397 723 2401
rect 855 2397 859 2401
rect 991 2397 995 2401
rect 1127 2397 1131 2401
rect 1263 2397 1267 2401
rect 1399 2397 1403 2401
rect 1863 2396 1867 2400
rect 1955 2399 1959 2403
rect 1963 2399 1967 2403
rect 2243 2399 2247 2403
rect 2403 2399 2407 2403
rect 3575 2396 3579 2400
rect 1895 2383 1899 2387
rect 2023 2383 2027 2387
rect 2183 2383 2187 2387
rect 2343 2383 2347 2387
rect 2503 2383 2507 2387
rect 2655 2383 2659 2387
rect 2807 2383 2811 2387
rect 2959 2383 2963 2387
rect 3119 2383 3123 2387
rect 1963 2371 1967 2375
rect 2031 2371 2035 2375
rect 2243 2371 2247 2375
rect 2403 2371 2407 2375
rect 2663 2371 2667 2375
rect 159 2363 163 2367
rect 247 2363 251 2367
rect 335 2363 339 2367
rect 439 2363 443 2367
rect 559 2363 563 2367
rect 687 2363 691 2367
rect 815 2363 819 2367
rect 951 2363 955 2367
rect 1079 2363 1083 2367
rect 1207 2363 1211 2367
rect 1327 2363 1331 2367
rect 1455 2363 1459 2367
rect 1583 2363 1587 2367
rect 111 2353 115 2357
rect 767 2355 771 2359
rect 887 2355 891 2359
rect 1523 2355 1527 2359
rect 1823 2353 1827 2357
rect 1955 2355 1959 2359
rect 2479 2363 2483 2367
rect 2567 2355 2571 2359
rect 2711 2355 2715 2359
rect 1927 2345 1931 2349
rect 2087 2345 2091 2349
rect 2247 2345 2251 2349
rect 2407 2345 2411 2349
rect 2559 2345 2563 2349
rect 2703 2345 2707 2349
rect 2831 2345 2835 2349
rect 2951 2345 2955 2349
rect 3071 2345 3075 2349
rect 3183 2345 3187 2349
rect 3287 2345 3291 2349
rect 3399 2345 3403 2349
rect 3487 2345 3491 2349
rect 111 2336 115 2340
rect 227 2339 231 2343
rect 315 2339 319 2343
rect 403 2339 407 2343
rect 655 2339 659 2343
rect 763 2339 767 2343
rect 1155 2339 1159 2343
rect 1403 2339 1407 2343
rect 1531 2339 1535 2343
rect 1823 2336 1827 2340
rect 1863 2332 1867 2336
rect 3575 2332 3579 2336
rect 167 2323 171 2327
rect 255 2323 259 2327
rect 343 2323 347 2327
rect 447 2323 451 2327
rect 567 2323 571 2327
rect 695 2323 699 2327
rect 823 2323 827 2327
rect 959 2323 963 2327
rect 1087 2323 1091 2327
rect 1215 2323 1219 2327
rect 1335 2323 1339 2327
rect 1463 2323 1467 2327
rect 1591 2323 1595 2327
rect 175 2311 179 2315
rect 227 2311 231 2315
rect 315 2311 319 2315
rect 403 2311 407 2315
rect 655 2311 659 2315
rect 763 2311 767 2315
rect 1135 2311 1139 2315
rect 1155 2311 1159 2315
rect 1403 2311 1407 2315
rect 1531 2311 1535 2315
rect 1863 2315 1867 2319
rect 2479 2315 2483 2319
rect 3183 2315 3187 2319
rect 3575 2315 3579 2319
rect 1919 2305 1923 2309
rect 2079 2305 2083 2309
rect 2239 2305 2243 2309
rect 2399 2305 2403 2309
rect 2551 2305 2555 2309
rect 2695 2305 2699 2309
rect 2823 2305 2827 2309
rect 2943 2305 2947 2309
rect 3063 2305 3067 2309
rect 3175 2305 3179 2309
rect 3279 2305 3283 2309
rect 3391 2305 3395 2309
rect 3479 2305 3483 2309
rect 703 2291 707 2295
rect 1031 2291 1035 2295
rect 1183 2291 1187 2295
rect 695 2281 699 2285
rect 863 2281 867 2285
rect 1023 2281 1027 2285
rect 1175 2281 1179 2285
rect 1319 2281 1323 2285
rect 1463 2281 1467 2285
rect 1599 2281 1603 2285
rect 1735 2281 1739 2285
rect 1975 2279 1979 2283
rect 2143 2279 2147 2283
rect 2311 2279 2315 2283
rect 2479 2279 2483 2283
rect 2639 2279 2643 2283
rect 2783 2279 2787 2283
rect 2919 2279 2923 2283
rect 3039 2279 3043 2283
rect 3159 2279 3163 2283
rect 3271 2279 3275 2283
rect 3383 2279 3387 2283
rect 3479 2279 3483 2283
rect 111 2268 115 2272
rect 939 2263 943 2267
rect 1823 2268 1827 2272
rect 1863 2269 1867 2273
rect 2567 2271 2571 2275
rect 3111 2271 3115 2275
rect 3575 2269 3579 2273
rect 111 2251 115 2255
rect 1667 2251 1671 2255
rect 1823 2251 1827 2255
rect 1863 2252 1867 2256
rect 2043 2255 2047 2259
rect 2051 2255 2055 2259
rect 3151 2255 3155 2259
rect 3339 2255 3343 2259
rect 3471 2255 3475 2259
rect 3575 2252 3579 2256
rect 687 2241 691 2245
rect 855 2241 859 2245
rect 1015 2241 1019 2245
rect 1167 2241 1171 2245
rect 1311 2241 1315 2245
rect 1455 2241 1459 2245
rect 1591 2241 1595 2245
rect 1727 2241 1731 2245
rect 1983 2239 1987 2243
rect 2151 2239 2155 2243
rect 2319 2239 2323 2243
rect 2487 2239 2491 2243
rect 2647 2239 2651 2243
rect 2791 2239 2795 2243
rect 2927 2239 2931 2243
rect 3047 2239 3051 2243
rect 3167 2239 3171 2243
rect 3279 2239 3283 2243
rect 3391 2239 3395 2243
rect 3487 2239 3491 2243
rect 2051 2227 2055 2231
rect 2403 2227 2407 2231
rect 2799 2227 2803 2231
rect 3151 2227 3155 2231
rect 3339 2227 3343 2231
rect 535 2211 539 2215
rect 719 2211 723 2215
rect 895 2211 899 2215
rect 1071 2211 1075 2215
rect 1239 2211 1243 2215
rect 1407 2211 1411 2215
rect 1575 2211 1579 2215
rect 1727 2211 1731 2215
rect 2043 2215 2047 2219
rect 2587 2215 2591 2219
rect 2839 2215 2843 2219
rect 3111 2215 3115 2219
rect 3471 2215 3475 2219
rect 111 2201 115 2205
rect 1031 2203 1035 2207
rect 1643 2203 1647 2207
rect 1823 2201 1827 2205
rect 2007 2205 2011 2209
rect 2167 2205 2171 2209
rect 2335 2205 2339 2209
rect 2519 2205 2523 2209
rect 2711 2205 2715 2209
rect 2903 2205 2907 2209
rect 3103 2205 3107 2209
rect 3303 2205 3307 2209
rect 3487 2205 3491 2209
rect 1863 2192 1867 2196
rect 111 2184 115 2188
rect 1823 2184 1827 2188
rect 2403 2187 2407 2191
rect 2587 2187 2591 2191
rect 3575 2192 3579 2196
rect 543 2171 547 2175
rect 727 2171 731 2175
rect 903 2171 907 2175
rect 1079 2171 1083 2175
rect 1247 2171 1251 2175
rect 1415 2171 1419 2175
rect 1583 2171 1587 2175
rect 1735 2171 1739 2175
rect 1863 2175 1867 2179
rect 2235 2175 2239 2179
rect 3575 2175 3579 2179
rect 1999 2165 2003 2169
rect 2159 2165 2163 2169
rect 2327 2165 2331 2169
rect 2511 2165 2515 2169
rect 2703 2165 2707 2169
rect 2895 2165 2899 2169
rect 3095 2165 3099 2169
rect 3295 2165 3299 2169
rect 3479 2165 3483 2169
rect 575 2159 579 2163
rect 1255 2159 1259 2163
rect 551 2147 555 2151
rect 1239 2147 1243 2151
rect 1539 2147 1543 2151
rect 1643 2147 1647 2151
rect 495 2137 499 2141
rect 623 2137 627 2141
rect 759 2137 763 2141
rect 895 2137 899 2141
rect 1039 2137 1043 2141
rect 1183 2137 1187 2141
rect 1327 2137 1331 2141
rect 1471 2137 1475 2141
rect 1623 2137 1627 2141
rect 2023 2135 2027 2139
rect 2167 2135 2171 2139
rect 2319 2135 2323 2139
rect 2471 2135 2475 2139
rect 2615 2135 2619 2139
rect 2759 2135 2763 2139
rect 2895 2135 2899 2139
rect 3023 2135 3027 2139
rect 3143 2135 3147 2139
rect 3263 2135 3267 2139
rect 3383 2135 3387 2139
rect 3479 2135 3483 2139
rect 111 2124 115 2128
rect 1823 2124 1827 2128
rect 1863 2125 1867 2129
rect 2839 2127 2843 2131
rect 3451 2127 3455 2131
rect 3575 2125 3579 2129
rect 1539 2119 1543 2123
rect 111 2107 115 2111
rect 1039 2107 1043 2111
rect 1399 2107 1403 2111
rect 1823 2107 1827 2111
rect 1863 2108 1867 2112
rect 2107 2111 2111 2115
rect 2827 2111 2831 2115
rect 2963 2111 2967 2115
rect 3091 2111 3095 2115
rect 3211 2111 3215 2115
rect 3471 2111 3475 2115
rect 3575 2108 3579 2112
rect 487 2097 491 2101
rect 615 2097 619 2101
rect 751 2097 755 2101
rect 887 2097 891 2101
rect 1031 2097 1035 2101
rect 1175 2097 1179 2101
rect 1319 2097 1323 2101
rect 1463 2097 1467 2101
rect 1615 2097 1619 2101
rect 1239 2091 1243 2095
rect 2031 2095 2035 2099
rect 2175 2095 2179 2099
rect 2327 2095 2331 2099
rect 2479 2095 2483 2099
rect 2623 2095 2627 2099
rect 2767 2095 2771 2099
rect 2903 2095 2907 2099
rect 3031 2095 3035 2099
rect 3151 2095 3155 2099
rect 3271 2095 3275 2099
rect 3391 2095 3395 2099
rect 3487 2095 3491 2099
rect 2107 2083 2111 2087
rect 2235 2083 2239 2087
rect 2303 2083 2307 2087
rect 2963 2083 2967 2087
rect 3091 2083 3095 2087
rect 3211 2083 3215 2087
rect 3451 2083 3455 2087
rect 319 2071 323 2075
rect 431 2071 435 2075
rect 551 2071 555 2075
rect 679 2071 683 2075
rect 799 2071 803 2075
rect 919 2071 923 2075
rect 1039 2071 1043 2075
rect 1159 2071 1163 2075
rect 1279 2071 1283 2075
rect 1407 2071 1411 2075
rect 111 2061 115 2065
rect 767 2063 771 2067
rect 2611 2067 2615 2071
rect 2827 2067 2831 2071
rect 3347 2067 3351 2071
rect 3459 2067 3463 2071
rect 3471 2067 3475 2071
rect 1823 2061 1827 2065
rect 1983 2057 1987 2061
rect 2143 2057 2147 2061
rect 2311 2057 2315 2061
rect 2471 2057 2475 2061
rect 2631 2057 2635 2061
rect 2775 2057 2779 2061
rect 2911 2057 2915 2061
rect 3039 2057 3043 2061
rect 3159 2057 3163 2061
rect 3279 2057 3283 2061
rect 3391 2057 3395 2061
rect 3487 2057 3491 2061
rect 111 2044 115 2048
rect 1127 2047 1131 2051
rect 1227 2047 1231 2051
rect 1347 2047 1351 2051
rect 1823 2044 1827 2048
rect 1863 2044 1867 2048
rect 2303 2039 2307 2043
rect 3575 2044 3579 2048
rect 3347 2039 3351 2043
rect 3459 2039 3463 2043
rect 327 2031 331 2035
rect 439 2031 443 2035
rect 559 2031 563 2035
rect 687 2031 691 2035
rect 807 2031 811 2035
rect 927 2031 931 2035
rect 1047 2031 1051 2035
rect 1167 2031 1171 2035
rect 1287 2031 1291 2035
rect 1415 2031 1419 2035
rect 1863 2027 1867 2031
rect 3575 2027 3579 2031
rect 1227 2019 1231 2023
rect 1347 2019 1351 2023
rect 1399 2019 1403 2023
rect 1975 2017 1979 2021
rect 2135 2017 2139 2021
rect 2303 2017 2307 2021
rect 2463 2017 2467 2021
rect 2623 2017 2627 2021
rect 2767 2017 2771 2021
rect 2903 2017 2907 2021
rect 3031 2017 3035 2021
rect 3151 2017 3155 2021
rect 3271 2017 3275 2021
rect 3383 2017 3387 2021
rect 3479 2017 3483 2021
rect 239 2003 243 2007
rect 843 2003 847 2007
rect 963 2003 967 2007
rect 1119 2003 1123 2007
rect 1127 2003 1128 2007
rect 1128 2003 1131 2007
rect 183 1993 187 1997
rect 295 1993 299 1997
rect 415 1993 419 1997
rect 535 1993 539 1997
rect 655 1993 659 1997
rect 775 1993 779 1997
rect 895 1993 899 1997
rect 1015 1993 1019 1997
rect 1135 1993 1139 1997
rect 1255 1993 1259 1997
rect 1887 1995 1891 1999
rect 2031 1995 2035 1999
rect 2199 1995 2203 1999
rect 2375 1995 2379 1999
rect 2543 1995 2547 1999
rect 2711 1995 2715 1999
rect 2871 1995 2875 1999
rect 3039 1995 3043 1999
rect 3207 1995 3211 1999
rect 1863 1985 1867 1989
rect 2611 1987 2615 1991
rect 3575 1985 3579 1989
rect 111 1980 115 1984
rect 843 1975 847 1979
rect 963 1975 967 1979
rect 1823 1980 1827 1984
rect 1863 1968 1867 1972
rect 1983 1971 1987 1975
rect 1991 1971 1995 1975
rect 2099 1971 2103 1975
rect 2999 1971 3003 1975
rect 3151 1971 3155 1975
rect 3159 1971 3163 1975
rect 111 1963 115 1967
rect 3575 1968 3579 1972
rect 175 1953 179 1957
rect 287 1953 291 1957
rect 407 1953 411 1957
rect 527 1953 531 1957
rect 647 1953 651 1957
rect 767 1953 771 1957
rect 887 1953 891 1957
rect 1007 1953 1011 1957
rect 1127 1953 1131 1957
rect 1119 1947 1123 1951
rect 1823 1963 1827 1967
rect 1247 1953 1251 1957
rect 1895 1955 1899 1959
rect 2039 1955 2043 1959
rect 2207 1955 2211 1959
rect 2383 1955 2387 1959
rect 2551 1955 2555 1959
rect 2719 1955 2723 1959
rect 2879 1955 2883 1959
rect 3047 1955 3051 1959
rect 3215 1955 3219 1959
rect 1991 1943 1995 1947
rect 2099 1943 2103 1947
rect 2339 1943 2343 1947
rect 2727 1943 2731 1947
rect 3151 1943 3155 1947
rect 135 1927 139 1931
rect 223 1927 227 1931
rect 351 1927 355 1931
rect 495 1927 499 1931
rect 655 1927 659 1931
rect 839 1927 843 1931
rect 1039 1927 1043 1931
rect 1247 1927 1251 1931
rect 1463 1927 1467 1931
rect 111 1917 115 1921
rect 563 1919 567 1923
rect 1159 1919 1163 1923
rect 1983 1923 1984 1927
rect 1984 1923 1987 1927
rect 2347 1923 2351 1927
rect 2367 1923 2371 1927
rect 2579 1923 2583 1927
rect 2699 1923 2703 1927
rect 2819 1923 2823 1927
rect 2947 1923 2951 1927
rect 2999 1923 3000 1927
rect 3000 1923 3003 1927
rect 1823 1917 1827 1921
rect 1895 1913 1899 1917
rect 1991 1913 1995 1917
rect 2119 1913 2123 1917
rect 2255 1913 2259 1917
rect 2383 1913 2387 1917
rect 2511 1913 2515 1917
rect 2631 1913 2635 1917
rect 2751 1913 2755 1917
rect 2879 1913 2883 1917
rect 3007 1913 3011 1917
rect 111 1900 115 1904
rect 1823 1900 1827 1904
rect 1863 1900 1867 1904
rect 2339 1899 2343 1903
rect 3575 1900 3579 1904
rect 2347 1895 2351 1899
rect 2579 1895 2583 1899
rect 2699 1895 2703 1899
rect 2819 1895 2823 1899
rect 2947 1895 2951 1899
rect 143 1887 147 1891
rect 231 1887 235 1891
rect 359 1887 363 1891
rect 503 1887 507 1891
rect 663 1887 667 1891
rect 847 1887 851 1891
rect 1047 1887 1051 1891
rect 1255 1887 1259 1891
rect 1471 1887 1475 1891
rect 1863 1883 1867 1887
rect 1871 1883 1875 1887
rect 2511 1883 2515 1887
rect 3575 1883 3579 1887
rect 135 1875 136 1879
rect 136 1875 139 1879
rect 1887 1873 1891 1877
rect 1983 1873 1987 1877
rect 2111 1873 2115 1877
rect 2247 1873 2251 1877
rect 2375 1873 2379 1877
rect 2503 1873 2507 1877
rect 2623 1873 2627 1877
rect 2743 1873 2747 1877
rect 2871 1873 2875 1877
rect 2999 1873 3003 1877
rect 211 1855 215 1859
rect 339 1855 343 1859
rect 371 1855 375 1859
rect 763 1855 767 1859
rect 891 1855 895 1859
rect 951 1855 955 1859
rect 1111 1855 1115 1859
rect 1427 1863 1431 1867
rect 1619 1855 1623 1859
rect 1715 1855 1719 1859
rect 1871 1855 1875 1859
rect 143 1845 147 1849
rect 271 1845 275 1849
rect 415 1845 419 1849
rect 559 1845 563 1849
rect 695 1845 699 1849
rect 823 1845 827 1849
rect 943 1845 947 1849
rect 1055 1845 1059 1849
rect 1159 1845 1163 1849
rect 1263 1845 1267 1849
rect 1359 1845 1363 1849
rect 1455 1845 1459 1849
rect 1551 1845 1555 1849
rect 1647 1845 1651 1849
rect 1735 1845 1739 1849
rect 2223 1843 2227 1847
rect 2359 1843 2363 1847
rect 2495 1843 2499 1847
rect 2623 1843 2627 1847
rect 2743 1843 2747 1847
rect 2863 1843 2867 1847
rect 2991 1843 2995 1847
rect 111 1832 115 1836
rect 135 1827 139 1831
rect 211 1827 215 1831
rect 339 1827 343 1831
rect 763 1827 767 1831
rect 891 1827 895 1831
rect 1823 1832 1827 1836
rect 1863 1833 1867 1837
rect 1427 1827 1431 1831
rect 1619 1827 1623 1831
rect 2367 1831 2371 1835
rect 2931 1835 2935 1839
rect 3575 1833 3579 1837
rect 1715 1827 1719 1831
rect 111 1815 115 1819
rect 511 1815 515 1819
rect 1551 1815 1555 1819
rect 1823 1815 1827 1819
rect 1863 1816 1867 1820
rect 3575 1816 3579 1820
rect 135 1805 139 1809
rect 263 1805 267 1809
rect 407 1805 411 1809
rect 551 1805 555 1809
rect 687 1805 691 1809
rect 815 1805 819 1809
rect 935 1805 939 1809
rect 1047 1805 1051 1809
rect 1151 1805 1155 1809
rect 1255 1805 1259 1809
rect 1351 1805 1355 1809
rect 1447 1805 1451 1809
rect 1543 1805 1547 1809
rect 1639 1805 1643 1809
rect 1727 1805 1731 1809
rect 1391 1799 1395 1803
rect 2231 1803 2235 1807
rect 2367 1803 2371 1807
rect 2503 1803 2507 1807
rect 2631 1803 2635 1807
rect 2751 1803 2755 1807
rect 2871 1803 2875 1807
rect 2999 1803 3003 1807
rect 2331 1791 2335 1795
rect 2511 1791 2515 1795
rect 135 1771 139 1775
rect 303 1771 307 1775
rect 495 1771 499 1775
rect 687 1771 691 1775
rect 871 1771 875 1775
rect 1047 1771 1051 1775
rect 1215 1771 1219 1775
rect 1375 1771 1379 1775
rect 1535 1771 1539 1775
rect 1703 1771 1707 1775
rect 2339 1775 2343 1779
rect 2427 1775 2431 1779
rect 2523 1775 2527 1779
rect 2723 1775 2727 1779
rect 2931 1783 2935 1787
rect 111 1761 115 1765
rect 371 1763 375 1767
rect 1115 1763 1119 1767
rect 1823 1761 1827 1765
rect 2271 1765 2275 1769
rect 2359 1765 2363 1769
rect 2455 1765 2459 1769
rect 2559 1765 2563 1769
rect 2663 1765 2667 1769
rect 2759 1765 2763 1769
rect 2863 1765 2867 1769
rect 2967 1765 2971 1769
rect 3071 1765 3075 1769
rect 3175 1765 3179 1769
rect 1863 1752 1867 1756
rect 111 1744 115 1748
rect 2331 1751 2335 1755
rect 1823 1744 1827 1748
rect 2339 1747 2343 1751
rect 2427 1747 2431 1751
rect 2523 1747 2527 1751
rect 3575 1752 3579 1756
rect 143 1731 147 1735
rect 311 1731 315 1735
rect 503 1731 507 1735
rect 695 1731 699 1735
rect 879 1731 883 1735
rect 1055 1731 1059 1735
rect 1223 1731 1227 1735
rect 1383 1731 1387 1735
rect 1543 1731 1547 1735
rect 1711 1731 1715 1735
rect 1863 1735 1867 1739
rect 2263 1725 2267 1729
rect 2351 1725 2355 1729
rect 2447 1725 2451 1729
rect 2551 1725 2555 1729
rect 2655 1725 2659 1729
rect 2751 1725 2755 1729
rect 2855 1725 2859 1729
rect 2959 1725 2963 1729
rect 3063 1725 3067 1729
rect 135 1719 136 1723
rect 136 1719 139 1723
rect 511 1719 515 1723
rect 1083 1719 1087 1723
rect 1391 1719 1395 1723
rect 1551 1719 1555 1723
rect 2903 1719 2907 1723
rect 3575 1735 3579 1739
rect 3167 1725 3171 1729
rect 383 1703 387 1707
rect 751 1703 755 1707
rect 999 1703 1003 1707
rect 1427 1703 1431 1707
rect 2247 1699 2251 1703
rect 2367 1699 2371 1703
rect 2495 1699 2499 1703
rect 2623 1699 2627 1703
rect 2759 1699 2763 1703
rect 2887 1699 2891 1703
rect 3015 1699 3019 1703
rect 3135 1699 3139 1703
rect 3247 1699 3251 1703
rect 3367 1699 3371 1703
rect 3479 1699 3483 1703
rect 143 1693 147 1697
rect 287 1693 291 1697
rect 471 1693 475 1697
rect 655 1693 659 1697
rect 839 1693 843 1697
rect 1023 1693 1027 1697
rect 1191 1693 1195 1697
rect 1359 1693 1363 1697
rect 1527 1693 1531 1697
rect 1695 1693 1699 1697
rect 1863 1689 1867 1693
rect 2723 1691 2727 1695
rect 3575 1689 3579 1693
rect 111 1680 115 1684
rect 135 1675 139 1679
rect 383 1675 387 1679
rect 751 1675 755 1679
rect 1083 1679 1087 1683
rect 1823 1680 1827 1684
rect 1427 1675 1431 1679
rect 1863 1672 1867 1676
rect 3127 1675 3131 1679
rect 3575 1672 3579 1676
rect 111 1663 115 1667
rect 287 1663 291 1667
rect 1167 1663 1171 1667
rect 1823 1663 1827 1667
rect 2255 1659 2259 1663
rect 2375 1659 2379 1663
rect 2503 1659 2507 1663
rect 2631 1659 2635 1663
rect 2767 1659 2771 1663
rect 2895 1659 2899 1663
rect 3023 1659 3027 1663
rect 3143 1659 3147 1663
rect 3255 1659 3259 1663
rect 3375 1659 3379 1663
rect 3487 1659 3491 1663
rect 135 1653 139 1657
rect 279 1653 283 1657
rect 463 1653 467 1657
rect 647 1653 651 1657
rect 831 1653 835 1657
rect 1015 1653 1019 1657
rect 1183 1653 1187 1657
rect 1351 1653 1355 1657
rect 1519 1653 1523 1657
rect 1687 1653 1691 1657
rect 2903 1647 2907 1651
rect 3127 1647 3131 1651
rect 3499 1647 3503 1651
rect 2159 1631 2163 1635
rect 3099 1639 3103 1643
rect 135 1623 139 1627
rect 271 1623 275 1627
rect 447 1623 451 1627
rect 631 1623 635 1627
rect 815 1623 819 1627
rect 991 1623 995 1627
rect 1151 1623 1155 1627
rect 1303 1623 1307 1627
rect 1455 1623 1459 1627
rect 1599 1623 1603 1627
rect 1727 1623 1731 1627
rect 2151 1621 2155 1625
rect 2343 1621 2347 1625
rect 2527 1621 2531 1625
rect 2703 1621 2707 1625
rect 2871 1621 2875 1625
rect 3031 1621 3035 1625
rect 3191 1621 3195 1625
rect 3351 1621 3355 1625
rect 3487 1621 3491 1625
rect 111 1613 115 1617
rect 999 1611 1003 1615
rect 1823 1613 1827 1617
rect 1863 1608 1867 1612
rect 111 1596 115 1600
rect 1583 1599 1587 1603
rect 1667 1599 1671 1603
rect 3575 1608 3579 1612
rect 3099 1603 3103 1607
rect 1823 1596 1827 1600
rect 1863 1591 1867 1595
rect 3471 1591 3475 1595
rect 3575 1591 3579 1595
rect 143 1583 147 1587
rect 279 1583 283 1587
rect 455 1583 459 1587
rect 639 1583 643 1587
rect 823 1583 827 1587
rect 999 1583 1003 1587
rect 1159 1583 1163 1587
rect 1311 1583 1315 1587
rect 1463 1583 1467 1587
rect 1607 1583 1611 1587
rect 1735 1583 1739 1587
rect 2143 1581 2147 1585
rect 2335 1581 2339 1585
rect 2519 1581 2523 1585
rect 2695 1581 2699 1585
rect 2863 1581 2867 1585
rect 3023 1581 3027 1585
rect 3183 1581 3187 1585
rect 3343 1581 3347 1585
rect 3479 1581 3483 1585
rect 135 1571 136 1575
rect 136 1571 139 1575
rect 287 1571 291 1575
rect 1027 1571 1031 1575
rect 1167 1571 1171 1575
rect 1667 1571 1671 1575
rect 2103 1567 2107 1571
rect 211 1559 215 1563
rect 251 1559 255 1563
rect 515 1559 519 1563
rect 667 1559 671 1563
rect 943 1559 947 1563
rect 1019 1559 1023 1563
rect 1343 1559 1347 1563
rect 1583 1559 1584 1563
rect 1584 1559 1587 1563
rect 1663 1559 1667 1563
rect 2087 1559 2091 1563
rect 2279 1559 2283 1563
rect 143 1549 147 1553
rect 271 1549 275 1553
rect 431 1549 435 1553
rect 599 1549 603 1553
rect 767 1549 771 1553
rect 935 1549 939 1553
rect 1103 1549 1107 1553
rect 1263 1549 1267 1553
rect 1423 1549 1427 1553
rect 1591 1549 1595 1553
rect 1735 1549 1739 1553
rect 1863 1549 1867 1553
rect 2159 1551 2163 1555
rect 2455 1559 2459 1563
rect 2623 1559 2627 1563
rect 2791 1559 2795 1563
rect 2951 1559 2955 1563
rect 3111 1559 3115 1563
rect 3271 1559 3275 1563
rect 3431 1559 3435 1563
rect 3215 1551 3219 1555
rect 3499 1551 3503 1555
rect 3575 1549 3579 1553
rect 111 1536 115 1540
rect 135 1531 139 1535
rect 211 1531 215 1535
rect 515 1531 519 1535
rect 667 1531 671 1535
rect 1019 1535 1023 1539
rect 1027 1531 1031 1535
rect 1343 1535 1347 1539
rect 1663 1535 1667 1539
rect 1823 1536 1827 1540
rect 1863 1532 1867 1536
rect 3079 1535 3083 1539
rect 3575 1532 3579 1536
rect 111 1519 115 1523
rect 351 1519 355 1523
rect 1391 1519 1395 1523
rect 1815 1519 1819 1523
rect 1823 1519 1827 1523
rect 2095 1519 2099 1523
rect 2287 1519 2291 1523
rect 2463 1519 2467 1523
rect 2631 1519 2635 1523
rect 2799 1519 2803 1523
rect 2959 1519 2963 1523
rect 3119 1519 3123 1523
rect 3279 1519 3283 1523
rect 3439 1519 3443 1523
rect 135 1509 139 1513
rect 263 1509 267 1513
rect 423 1509 427 1513
rect 591 1509 595 1513
rect 759 1509 763 1513
rect 927 1509 931 1513
rect 1095 1509 1099 1513
rect 1255 1509 1259 1513
rect 1415 1509 1419 1513
rect 1583 1509 1587 1513
rect 1727 1509 1731 1513
rect 2103 1507 2107 1511
rect 2179 1507 2183 1511
rect 2639 1507 2643 1511
rect 183 1483 187 1487
rect 327 1483 331 1487
rect 471 1483 475 1487
rect 607 1483 611 1487
rect 743 1483 747 1487
rect 871 1483 875 1487
rect 991 1483 995 1487
rect 1119 1483 1123 1487
rect 1247 1483 1251 1487
rect 1375 1483 1379 1487
rect 1815 1487 1819 1491
rect 2187 1487 2191 1491
rect 2391 1487 2395 1491
rect 2779 1495 2783 1499
rect 3219 1495 3223 1499
rect 3079 1487 3080 1491
rect 3080 1487 3083 1491
rect 3471 1487 3475 1491
rect 111 1473 115 1477
rect 251 1475 255 1479
rect 943 1475 947 1479
rect 1823 1473 1827 1477
rect 1895 1477 1899 1481
rect 1991 1477 1995 1481
rect 2119 1477 2123 1481
rect 2247 1477 2251 1481
rect 2383 1477 2387 1481
rect 2535 1477 2539 1481
rect 2703 1477 2707 1481
rect 2887 1477 2891 1481
rect 3087 1477 3091 1481
rect 3295 1477 3299 1481
rect 3487 1477 3491 1481
rect 1863 1464 1867 1468
rect 111 1456 115 1460
rect 939 1459 943 1463
rect 1059 1459 1063 1463
rect 1315 1459 1319 1463
rect 2179 1463 2183 1467
rect 1823 1456 1827 1460
rect 2187 1459 2191 1463
rect 2779 1459 2783 1463
rect 3575 1464 3579 1468
rect 3219 1459 3223 1463
rect 191 1443 195 1447
rect 335 1443 339 1447
rect 479 1443 483 1447
rect 615 1443 619 1447
rect 751 1443 755 1447
rect 879 1443 883 1447
rect 999 1443 1003 1447
rect 1127 1443 1131 1447
rect 1255 1443 1259 1447
rect 1383 1443 1387 1447
rect 1863 1447 1867 1451
rect 3575 1447 3579 1451
rect 1887 1437 1891 1441
rect 1983 1437 1987 1441
rect 2111 1437 2115 1441
rect 2239 1437 2243 1441
rect 2375 1437 2379 1441
rect 2527 1437 2531 1441
rect 2695 1437 2699 1441
rect 2879 1437 2883 1441
rect 3079 1437 3083 1441
rect 3287 1437 3291 1441
rect 3479 1437 3483 1441
rect 183 1431 184 1435
rect 184 1431 187 1435
rect 351 1431 355 1435
rect 939 1431 943 1435
rect 1059 1431 1063 1435
rect 1111 1431 1115 1435
rect 1315 1431 1319 1435
rect 1391 1431 1395 1435
rect 271 1411 275 1415
rect 299 1411 303 1415
rect 659 1419 663 1423
rect 771 1411 775 1415
rect 1887 1411 1891 1415
rect 1975 1411 1979 1415
rect 2071 1411 2075 1415
rect 2183 1411 2187 1415
rect 2303 1411 2307 1415
rect 2439 1411 2443 1415
rect 2607 1411 2611 1415
rect 2807 1411 2811 1415
rect 3031 1411 3035 1415
rect 3263 1411 3267 1415
rect 3479 1411 3483 1415
rect 199 1401 203 1405
rect 335 1401 339 1405
rect 463 1401 467 1405
rect 583 1401 587 1405
rect 703 1401 707 1405
rect 815 1401 819 1405
rect 919 1401 923 1405
rect 1015 1401 1019 1405
rect 1119 1401 1123 1405
rect 1223 1401 1227 1405
rect 1327 1401 1331 1405
rect 1863 1401 1867 1405
rect 2391 1403 2395 1407
rect 3211 1403 3215 1407
rect 3575 1401 3579 1405
rect 111 1388 115 1392
rect 183 1383 187 1387
rect 271 1383 275 1387
rect 659 1383 663 1387
rect 1111 1383 1115 1387
rect 1823 1388 1827 1392
rect 1863 1384 1867 1388
rect 1955 1387 1959 1391
rect 2043 1387 2047 1391
rect 2251 1387 2255 1391
rect 2371 1387 2375 1391
rect 2507 1387 2511 1391
rect 3255 1387 3259 1391
rect 3471 1387 3475 1391
rect 3575 1384 3579 1388
rect 111 1371 115 1375
rect 1823 1371 1827 1375
rect 1895 1371 1899 1375
rect 1983 1371 1987 1375
rect 2079 1371 2083 1375
rect 2191 1371 2195 1375
rect 2311 1371 2315 1375
rect 2447 1371 2451 1375
rect 2615 1371 2619 1375
rect 2815 1371 2819 1375
rect 3039 1371 3043 1375
rect 3271 1371 3275 1375
rect 3487 1371 3491 1375
rect 191 1361 195 1365
rect 327 1361 331 1365
rect 455 1361 459 1365
rect 575 1361 579 1365
rect 695 1361 699 1365
rect 807 1361 811 1365
rect 911 1361 915 1365
rect 1007 1361 1011 1365
rect 1111 1361 1115 1365
rect 1215 1361 1219 1365
rect 1319 1361 1323 1365
rect 1367 1355 1368 1359
rect 1368 1355 1371 1359
rect 1955 1359 1959 1363
rect 2043 1359 2047 1363
rect 2251 1359 2255 1363
rect 2507 1359 2511 1363
rect 2775 1359 2779 1363
rect 3255 1359 3259 1363
rect 2371 1343 2375 1347
rect 3255 1343 3259 1347
rect 3471 1343 3475 1347
rect 231 1335 235 1339
rect 383 1335 387 1339
rect 543 1335 547 1339
rect 703 1335 707 1339
rect 871 1335 875 1339
rect 1039 1335 1043 1339
rect 1207 1335 1211 1339
rect 1375 1335 1379 1339
rect 1895 1333 1899 1337
rect 1983 1333 1987 1337
rect 2103 1333 2107 1337
rect 2223 1333 2227 1337
rect 2359 1333 2363 1337
rect 2511 1333 2515 1337
rect 2687 1333 2691 1337
rect 2871 1333 2875 1337
rect 3071 1333 3075 1337
rect 3279 1333 3283 1337
rect 3487 1333 3491 1337
rect 111 1325 115 1329
rect 299 1327 303 1331
rect 771 1327 775 1331
rect 1823 1325 1827 1329
rect 1863 1320 1867 1324
rect 111 1308 115 1312
rect 451 1311 455 1315
rect 799 1311 803 1315
rect 1107 1311 1111 1315
rect 1275 1311 1279 1315
rect 3575 1320 3579 1324
rect 1823 1308 1827 1312
rect 1863 1303 1867 1307
rect 2959 1303 2963 1307
rect 3455 1303 3459 1307
rect 3575 1303 3579 1307
rect 239 1295 243 1299
rect 391 1295 395 1299
rect 551 1295 555 1299
rect 711 1295 715 1299
rect 879 1295 883 1299
rect 1047 1295 1051 1299
rect 1215 1295 1219 1299
rect 1383 1295 1387 1299
rect 1887 1293 1891 1297
rect 1975 1293 1979 1297
rect 2095 1293 2099 1297
rect 2215 1293 2219 1297
rect 2351 1293 2355 1297
rect 2503 1293 2507 1297
rect 2679 1293 2683 1297
rect 2863 1293 2867 1297
rect 3063 1293 3067 1297
rect 3271 1293 3275 1297
rect 3479 1293 3483 1297
rect 451 1283 455 1287
rect 559 1283 563 1287
rect 899 1283 903 1287
rect 1107 1283 1111 1287
rect 1275 1283 1279 1287
rect 1367 1283 1371 1287
rect 199 1271 203 1275
rect 215 1261 219 1265
rect 359 1261 363 1265
rect 519 1261 523 1265
rect 679 1261 683 1265
rect 839 1261 843 1265
rect 999 1261 1003 1265
rect 1151 1261 1155 1265
rect 1295 1261 1299 1265
rect 1439 1261 1443 1265
rect 1591 1261 1595 1265
rect 2055 1259 2059 1263
rect 2143 1259 2147 1263
rect 2239 1259 2243 1263
rect 2335 1259 2339 1263
rect 2431 1259 2435 1263
rect 2551 1259 2555 1263
rect 2687 1259 2691 1263
rect 2855 1259 2859 1263
rect 3039 1259 3043 1263
rect 3231 1259 3235 1263
rect 3431 1259 3435 1263
rect 111 1248 115 1252
rect 899 1247 903 1251
rect 1823 1248 1827 1252
rect 1863 1249 1867 1253
rect 2123 1251 2127 1255
rect 3107 1251 3111 1255
rect 3575 1249 3579 1253
rect 111 1231 115 1235
rect 1591 1231 1595 1235
rect 1823 1231 1827 1235
rect 1863 1232 1867 1236
rect 2211 1235 2215 1239
rect 2403 1235 2407 1239
rect 3499 1235 3503 1239
rect 3575 1232 3579 1236
rect 207 1221 211 1225
rect 351 1221 355 1225
rect 511 1221 515 1225
rect 671 1221 675 1225
rect 831 1221 835 1225
rect 991 1221 995 1225
rect 1143 1221 1147 1225
rect 1287 1221 1291 1225
rect 1431 1221 1435 1225
rect 1583 1221 1587 1225
rect 2063 1219 2067 1223
rect 2151 1219 2155 1223
rect 2247 1219 2251 1223
rect 2343 1219 2347 1223
rect 2439 1219 2443 1223
rect 2559 1219 2563 1223
rect 2695 1219 2699 1223
rect 2863 1219 2867 1223
rect 3047 1219 3051 1223
rect 3239 1219 3243 1223
rect 3439 1219 3443 1223
rect 2123 1207 2127 1211
rect 2211 1207 2215 1211
rect 2403 1207 2407 1211
rect 2475 1207 2479 1211
rect 2567 1207 2571 1211
rect 3455 1207 3459 1211
rect 135 1191 139 1195
rect 271 1191 275 1195
rect 423 1191 427 1195
rect 575 1191 579 1195
rect 727 1191 731 1195
rect 887 1191 891 1195
rect 1055 1191 1059 1195
rect 1231 1191 1235 1195
rect 1415 1191 1419 1195
rect 1599 1191 1603 1195
rect 2483 1191 2487 1195
rect 2543 1191 2547 1195
rect 2779 1191 2783 1195
rect 2935 1191 2939 1195
rect 3107 1191 3111 1195
rect 3247 1191 3251 1195
rect 3499 1191 3503 1195
rect 111 1181 115 1185
rect 203 1183 207 1187
rect 1823 1181 1827 1185
rect 2039 1181 2043 1185
rect 2151 1181 2155 1185
rect 2279 1181 2283 1185
rect 2415 1181 2419 1185
rect 2559 1181 2563 1185
rect 2711 1181 2715 1185
rect 2863 1181 2867 1185
rect 3015 1181 3019 1185
rect 3167 1181 3171 1185
rect 3327 1181 3331 1185
rect 3487 1181 3491 1185
rect 111 1164 115 1168
rect 203 1167 207 1171
rect 339 1167 343 1171
rect 655 1167 659 1171
rect 795 1167 799 1171
rect 955 1167 959 1171
rect 1123 1167 1127 1171
rect 1539 1167 1543 1171
rect 1823 1164 1827 1168
rect 1863 1168 1867 1172
rect 2475 1167 2479 1171
rect 3255 1171 3259 1175
rect 3575 1168 3579 1172
rect 2483 1163 2487 1167
rect 2779 1163 2783 1167
rect 2935 1163 2939 1167
rect 3247 1163 3251 1167
rect 143 1151 147 1155
rect 279 1151 283 1155
rect 431 1151 435 1155
rect 583 1151 587 1155
rect 735 1151 739 1155
rect 895 1151 899 1155
rect 1063 1151 1067 1155
rect 1239 1151 1243 1155
rect 1423 1151 1427 1155
rect 1607 1151 1611 1155
rect 1863 1151 1867 1155
rect 1959 1151 1963 1155
rect 2711 1151 2715 1155
rect 3575 1151 3579 1155
rect 203 1139 207 1143
rect 339 1139 343 1143
rect 795 1139 799 1143
rect 955 1139 959 1143
rect 1123 1139 1127 1143
rect 1267 1139 1271 1143
rect 1539 1139 1543 1143
rect 1591 1139 1595 1143
rect 2031 1141 2035 1145
rect 2143 1141 2147 1145
rect 2271 1141 2275 1145
rect 2407 1141 2411 1145
rect 2551 1141 2555 1145
rect 2703 1141 2707 1145
rect 2855 1141 2859 1145
rect 3007 1141 3011 1145
rect 3159 1141 3163 1145
rect 3319 1141 3323 1145
rect 3479 1141 3483 1145
rect 595 1127 599 1131
rect 655 1127 656 1131
rect 656 1127 659 1131
rect 967 1127 971 1131
rect 143 1117 147 1121
rect 295 1117 299 1121
rect 479 1117 483 1121
rect 663 1117 667 1121
rect 847 1117 851 1121
rect 1031 1117 1035 1121
rect 1207 1117 1211 1121
rect 1391 1117 1395 1121
rect 1575 1117 1579 1121
rect 1735 1117 1739 1121
rect 111 1104 115 1108
rect 1267 1103 1271 1107
rect 1823 1104 1827 1108
rect 1943 1107 1947 1111
rect 2087 1107 2091 1111
rect 2231 1107 2235 1111
rect 2383 1107 2387 1111
rect 2535 1107 2539 1111
rect 2687 1107 2691 1111
rect 2839 1107 2843 1111
rect 2991 1107 2995 1111
rect 3151 1107 3155 1111
rect 3319 1107 3323 1111
rect 3479 1107 3483 1111
rect 1863 1097 1867 1101
rect 2155 1099 2159 1103
rect 2543 1095 2547 1099
rect 3079 1099 3083 1103
rect 3575 1097 3579 1101
rect 111 1087 115 1091
rect 363 1087 367 1091
rect 135 1077 139 1081
rect 287 1077 291 1081
rect 471 1077 475 1081
rect 655 1077 659 1081
rect 595 1071 599 1075
rect 1823 1087 1827 1091
rect 839 1077 843 1081
rect 1023 1077 1027 1081
rect 1199 1077 1203 1081
rect 1383 1077 1387 1081
rect 1567 1077 1571 1081
rect 1727 1077 1731 1081
rect 1863 1080 1867 1084
rect 3471 1083 3475 1087
rect 3575 1080 3579 1084
rect 1951 1067 1955 1071
rect 2095 1067 2099 1071
rect 2239 1067 2243 1071
rect 2391 1067 2395 1071
rect 2543 1067 2547 1071
rect 2695 1067 2699 1071
rect 2847 1067 2851 1071
rect 2999 1067 3003 1071
rect 3159 1067 3163 1071
rect 3327 1067 3331 1071
rect 3487 1067 3491 1071
rect 135 1055 139 1059
rect 271 1055 275 1059
rect 431 1055 435 1059
rect 583 1055 587 1059
rect 735 1055 739 1059
rect 887 1055 891 1059
rect 1047 1055 1051 1059
rect 1215 1055 1219 1059
rect 1383 1055 1387 1059
rect 1559 1055 1563 1059
rect 1727 1055 1731 1059
rect 1959 1055 1963 1059
rect 2711 1055 2715 1059
rect 111 1045 115 1049
rect 967 1047 971 1051
rect 1283 1047 1287 1051
rect 1823 1045 1827 1049
rect 111 1028 115 1032
rect 815 1031 819 1035
rect 955 1031 959 1035
rect 1647 1031 1651 1035
rect 1823 1028 1827 1032
rect 1987 1031 1991 1035
rect 2155 1031 2159 1035
rect 2527 1031 2531 1035
rect 2703 1031 2707 1035
rect 3351 1031 3355 1035
rect 3471 1031 3475 1035
rect 1919 1021 1923 1025
rect 2127 1021 2131 1025
rect 2327 1021 2331 1025
rect 2519 1021 2523 1025
rect 2695 1021 2699 1025
rect 2863 1021 2867 1025
rect 3023 1021 3027 1025
rect 3183 1021 3187 1025
rect 3343 1021 3347 1025
rect 3487 1021 3491 1025
rect 143 1015 147 1019
rect 279 1015 283 1019
rect 439 1015 443 1019
rect 591 1015 595 1019
rect 743 1015 747 1019
rect 895 1015 899 1019
rect 1055 1015 1059 1019
rect 1223 1015 1227 1019
rect 1391 1015 1395 1019
rect 1567 1015 1571 1019
rect 1735 1015 1739 1019
rect 1863 1008 1867 1012
rect 363 1003 367 1007
rect 955 1003 959 1007
rect 1063 1003 1067 1007
rect 1231 1003 1235 1007
rect 1987 1003 1991 1007
rect 3575 1008 3579 1012
rect 815 987 816 991
rect 816 987 819 991
rect 1007 987 1011 991
rect 1579 995 1583 999
rect 1647 987 1648 991
rect 1648 987 1651 991
rect 1863 991 1867 995
rect 1903 991 1907 995
rect 3111 991 3115 995
rect 3575 991 3579 995
rect 143 977 147 981
rect 287 977 291 981
rect 463 977 467 981
rect 647 977 651 981
rect 823 977 827 981
rect 999 977 1003 981
rect 1167 977 1171 981
rect 1327 977 1331 981
rect 1487 977 1491 981
rect 1655 977 1659 981
rect 1911 981 1915 985
rect 2119 981 2123 985
rect 2319 981 2323 985
rect 2511 981 2515 985
rect 2687 981 2691 985
rect 2855 981 2859 985
rect 3015 981 3019 985
rect 3175 981 3179 985
rect 3335 981 3339 985
rect 3479 981 3483 985
rect 111 964 115 968
rect 1231 963 1235 967
rect 1823 964 1827 968
rect 1579 959 1583 963
rect 1887 955 1891 959
rect 2071 955 2075 959
rect 2263 955 2267 959
rect 2455 955 2459 959
rect 2631 955 2635 959
rect 2799 955 2803 959
rect 2951 955 2955 959
rect 3095 955 3099 959
rect 3231 955 3235 959
rect 3367 955 3371 959
rect 3479 955 3483 959
rect 111 947 115 951
rect 1823 947 1827 951
rect 1863 945 1867 949
rect 2527 947 2531 951
rect 3351 947 3355 951
rect 3575 945 3579 949
rect 135 937 139 941
rect 279 937 283 941
rect 455 937 459 941
rect 639 937 643 941
rect 815 937 819 941
rect 991 937 995 941
rect 1159 937 1163 941
rect 1319 937 1323 941
rect 1479 937 1483 941
rect 1647 937 1651 941
rect 1863 928 1867 932
rect 2175 931 2179 935
rect 3471 931 3475 935
rect 3575 928 3579 932
rect 1895 915 1899 919
rect 2079 915 2083 919
rect 2271 915 2275 919
rect 2463 915 2467 919
rect 2639 915 2643 919
rect 2807 915 2811 919
rect 2959 915 2963 919
rect 3103 915 3107 919
rect 3239 915 3243 919
rect 3375 915 3379 919
rect 3487 915 3491 919
rect 135 907 139 911
rect 271 907 275 911
rect 439 907 443 911
rect 607 907 611 911
rect 775 907 779 911
rect 935 907 939 911
rect 1095 907 1099 911
rect 1247 907 1251 911
rect 1399 907 1403 911
rect 1551 907 1555 911
rect 111 897 115 901
rect 707 899 711 903
rect 1007 899 1011 903
rect 1903 903 1907 907
rect 2815 903 2819 907
rect 1823 897 1827 901
rect 111 880 115 884
rect 203 883 207 887
rect 339 883 343 887
rect 1003 883 1007 887
rect 1495 883 1499 887
rect 1823 880 1827 884
rect 1963 883 1967 887
rect 2175 883 2176 887
rect 2176 883 2179 887
rect 2439 883 2443 887
rect 2607 883 2611 887
rect 2695 883 2699 887
rect 2907 883 2911 887
rect 3051 883 3055 887
rect 3199 883 3203 887
rect 3315 883 3319 887
rect 3471 883 3475 887
rect 1895 873 1899 877
rect 2023 873 2027 877
rect 2183 873 2187 877
rect 2351 873 2355 877
rect 2519 873 2523 877
rect 2687 873 2691 877
rect 2839 873 2843 877
rect 2983 873 2987 877
rect 3119 873 3123 877
rect 3247 873 3251 877
rect 3375 873 3379 877
rect 3487 873 3491 877
rect 143 867 147 871
rect 279 867 283 871
rect 447 867 451 871
rect 615 867 619 871
rect 783 867 787 871
rect 943 867 947 871
rect 1103 867 1107 871
rect 1255 867 1259 871
rect 1407 867 1411 871
rect 1559 867 1563 871
rect 1863 860 1867 864
rect 3575 860 3579 864
rect 199 855 203 859
rect 455 855 459 859
rect 1003 855 1007 859
rect 1263 855 1267 859
rect 1963 855 1967 859
rect 2439 855 2443 859
rect 2607 855 2611 859
rect 2907 855 2911 859
rect 3051 855 3055 859
rect 3199 855 3203 859
rect 3315 855 3319 859
rect 339 843 343 847
rect 1059 843 1063 847
rect 1167 843 1171 847
rect 1863 843 1867 847
rect 2807 843 2811 847
rect 3575 843 3579 847
rect 143 833 147 837
rect 287 833 291 837
rect 463 833 467 837
rect 639 833 643 837
rect 807 833 811 837
rect 983 833 987 837
rect 1159 833 1163 837
rect 1335 833 1339 837
rect 1511 833 1515 837
rect 1887 833 1891 837
rect 2015 833 2019 837
rect 2175 833 2179 837
rect 2343 833 2347 837
rect 2511 833 2515 837
rect 2679 833 2683 837
rect 2831 833 2835 837
rect 2975 833 2979 837
rect 3111 833 3115 837
rect 3239 833 3243 837
rect 3367 833 3371 837
rect 3479 833 3483 837
rect 111 820 115 824
rect 1823 820 1827 824
rect 1059 815 1063 819
rect 111 803 115 807
rect 791 803 795 807
rect 1295 803 1299 807
rect 1823 803 1827 807
rect 1887 803 1891 807
rect 2071 803 2075 807
rect 2263 803 2267 807
rect 2447 803 2451 807
rect 2623 803 2627 807
rect 2791 803 2795 807
rect 2943 803 2947 807
rect 3087 803 3091 807
rect 3223 803 3227 807
rect 3359 803 3363 807
rect 3479 803 3483 807
rect 135 793 139 797
rect 279 793 283 797
rect 455 793 459 797
rect 631 793 635 797
rect 799 793 803 797
rect 975 793 979 797
rect 1151 793 1155 797
rect 1327 793 1331 797
rect 1503 793 1507 797
rect 1863 793 1867 797
rect 1955 795 1959 799
rect 2695 795 2699 799
rect 3575 793 3579 797
rect 1863 776 1867 780
rect 3159 779 3163 783
rect 3427 779 3431 783
rect 3575 776 3579 780
rect 135 767 139 771
rect 271 767 275 771
rect 439 767 443 771
rect 607 767 611 771
rect 775 767 779 771
rect 935 767 939 771
rect 1087 767 1091 771
rect 1239 767 1243 771
rect 1391 767 1395 771
rect 1551 767 1555 771
rect 111 757 115 761
rect 1167 759 1171 763
rect 1895 763 1899 767
rect 2079 763 2083 767
rect 2271 763 2275 767
rect 2455 763 2459 767
rect 2631 763 2635 767
rect 2799 763 2803 767
rect 2951 763 2955 767
rect 3095 763 3099 767
rect 3231 763 3235 767
rect 3367 763 3371 767
rect 3487 763 3491 767
rect 1823 757 1827 761
rect 2255 751 2259 755
rect 2807 751 2811 755
rect 111 740 115 744
rect 203 743 207 747
rect 507 743 511 747
rect 675 743 679 747
rect 1619 743 1623 747
rect 1823 740 1827 744
rect 1955 739 1959 743
rect 2375 739 2379 743
rect 2463 739 2467 743
rect 2647 739 2651 743
rect 3055 739 3059 743
rect 3159 739 3163 743
rect 3427 743 3431 747
rect 143 727 147 731
rect 279 727 283 731
rect 447 727 451 731
rect 615 727 619 731
rect 783 727 787 731
rect 943 727 947 731
rect 1095 727 1099 731
rect 1247 727 1251 731
rect 1399 727 1403 731
rect 1559 727 1563 731
rect 1895 729 1899 733
rect 2071 729 2075 733
rect 2263 729 2267 733
rect 2447 729 2451 733
rect 2623 729 2627 733
rect 2799 729 2803 733
rect 2975 729 2979 733
rect 3151 729 3155 733
rect 3327 729 3331 733
rect 3487 729 3491 733
rect 203 715 207 719
rect 271 715 272 719
rect 272 715 275 719
rect 507 715 511 719
rect 675 715 679 719
rect 791 715 795 719
rect 1295 715 1299 719
rect 1863 716 1867 720
rect 2255 711 2259 715
rect 2375 711 2379 715
rect 3575 716 3579 720
rect 3259 711 3263 715
rect 215 699 219 703
rect 527 699 531 703
rect 711 699 715 703
rect 1027 699 1031 703
rect 1363 699 1367 703
rect 1515 699 1519 703
rect 1619 699 1623 703
rect 1863 699 1867 703
rect 143 689 147 693
rect 287 689 291 693
rect 455 689 459 693
rect 623 689 627 693
rect 791 689 795 693
rect 959 689 963 693
rect 1119 689 1123 693
rect 1279 689 1283 693
rect 1439 689 1443 693
rect 1599 689 1603 693
rect 1887 689 1891 693
rect 2063 689 2067 693
rect 2255 689 2259 693
rect 2439 689 2443 693
rect 2615 689 2619 693
rect 2791 689 2795 693
rect 2111 683 2112 687
rect 2112 683 2115 687
rect 2647 683 2651 687
rect 3575 699 3579 703
rect 2967 689 2971 693
rect 3143 689 3147 693
rect 3319 689 3323 693
rect 3479 689 3483 693
rect 111 676 115 680
rect 215 675 219 679
rect 271 671 275 675
rect 527 675 531 679
rect 711 675 715 679
rect 1823 676 1827 680
rect 1027 671 1031 675
rect 1363 671 1367 675
rect 1515 671 1519 675
rect 111 659 115 663
rect 791 659 795 663
rect 1823 659 1827 663
rect 1887 663 1891 667
rect 1975 663 1979 667
rect 2095 663 2099 667
rect 2223 663 2227 667
rect 2351 663 2355 667
rect 2479 663 2483 667
rect 2615 663 2619 667
rect 2767 663 2771 667
rect 2935 663 2939 667
rect 3119 663 3123 667
rect 3311 663 3315 667
rect 3479 663 3483 667
rect 135 649 139 653
rect 279 649 283 653
rect 447 649 451 653
rect 615 649 619 653
rect 783 649 787 653
rect 951 649 955 653
rect 1111 649 1115 653
rect 1271 649 1275 653
rect 1431 649 1435 653
rect 1591 649 1595 653
rect 1863 653 1867 657
rect 2463 655 2467 659
rect 3575 653 3579 657
rect 1863 636 1867 640
rect 1955 639 1959 643
rect 2043 639 2047 643
rect 2835 639 2839 643
rect 3227 639 3231 643
rect 3235 639 3239 643
rect 3471 639 3475 643
rect 3575 636 3579 640
rect 135 619 139 623
rect 287 619 291 623
rect 455 619 459 623
rect 631 619 635 623
rect 799 619 803 623
rect 967 619 971 623
rect 1119 619 1123 623
rect 1271 619 1275 623
rect 1415 619 1419 623
rect 1559 619 1563 623
rect 1711 619 1715 623
rect 1895 623 1899 627
rect 1983 623 1987 627
rect 2103 623 2107 627
rect 2231 623 2235 627
rect 2359 623 2363 627
rect 2487 623 2491 627
rect 2623 623 2627 627
rect 2775 623 2779 627
rect 2943 623 2947 627
rect 3127 623 3131 627
rect 3319 623 3323 627
rect 3487 623 3491 627
rect 111 609 115 613
rect 1639 611 1643 615
rect 1823 609 1827 613
rect 1955 611 1959 615
rect 2043 611 2047 615
rect 2111 611 2115 615
rect 2207 611 2211 615
rect 2631 611 2635 615
rect 3227 611 3231 615
rect 111 592 115 596
rect 203 595 207 599
rect 523 595 527 599
rect 699 595 703 599
rect 1823 592 1827 596
rect 2055 595 2059 599
rect 2835 595 2839 599
rect 3471 595 3475 599
rect 1895 585 1899 589
rect 2047 585 2051 589
rect 2215 585 2219 589
rect 2391 585 2395 589
rect 2583 585 2587 589
rect 2799 585 2803 589
rect 3023 585 3027 589
rect 3255 585 3259 589
rect 3487 585 3491 589
rect 143 579 147 583
rect 295 579 299 583
rect 463 579 467 583
rect 639 579 643 583
rect 807 579 811 583
rect 975 579 979 583
rect 1127 579 1131 583
rect 1279 579 1283 583
rect 1423 579 1427 583
rect 1567 579 1571 583
rect 1719 579 1723 583
rect 1863 572 1867 576
rect 203 567 207 571
rect 523 567 527 571
rect 699 567 703 571
rect 791 567 795 571
rect 987 567 991 571
rect 2207 567 2211 571
rect 3575 572 3579 576
rect 995 551 999 555
rect 1075 551 1079 555
rect 1199 551 1203 555
rect 1603 551 1607 555
rect 1671 551 1675 555
rect 1863 555 1867 559
rect 3575 555 3579 559
rect 151 541 155 545
rect 311 541 315 545
rect 471 541 475 545
rect 631 541 635 545
rect 783 541 787 545
rect 927 541 931 545
rect 1063 541 1067 545
rect 1191 541 1195 545
rect 1311 541 1315 545
rect 1423 541 1427 545
rect 1535 541 1539 545
rect 1647 541 1651 545
rect 1735 541 1739 545
rect 1887 545 1891 549
rect 2039 545 2043 549
rect 2207 545 2211 549
rect 2383 545 2387 549
rect 2575 545 2579 549
rect 2791 545 2795 549
rect 3015 545 3019 549
rect 3247 545 3251 549
rect 3479 545 3483 549
rect 111 528 115 532
rect 987 527 991 531
rect 995 523 999 527
rect 1823 528 1827 532
rect 1603 523 1607 527
rect 2055 523 2059 527
rect 111 511 115 515
rect 783 511 787 515
rect 1491 511 1495 515
rect 143 501 147 505
rect 303 501 307 505
rect 463 501 467 505
rect 623 501 627 505
rect 775 501 779 505
rect 919 501 923 505
rect 1055 501 1059 505
rect 1183 501 1187 505
rect 1303 501 1307 505
rect 1415 501 1419 505
rect 1527 501 1531 505
rect 1639 501 1643 505
rect 1455 495 1459 499
rect 1823 511 1827 515
rect 2191 515 2195 519
rect 2279 515 2283 519
rect 2375 515 2379 519
rect 2487 515 2491 519
rect 2631 515 2635 519
rect 2807 515 2811 519
rect 3007 515 3011 519
rect 3215 515 3219 519
rect 3431 515 3435 519
rect 1727 501 1731 505
rect 1863 505 1867 509
rect 3575 505 3579 509
rect 1671 487 1675 491
rect 1863 488 1867 492
rect 2347 491 2351 495
rect 3187 491 3191 495
rect 3499 491 3503 495
rect 3575 488 3579 492
rect 159 471 163 475
rect 311 471 315 475
rect 463 471 467 475
rect 615 471 619 475
rect 759 471 763 475
rect 887 471 891 475
rect 1007 471 1011 475
rect 1127 471 1131 475
rect 1239 471 1243 475
rect 1343 471 1347 475
rect 1439 471 1443 475
rect 1543 471 1547 475
rect 1639 471 1643 475
rect 1727 471 1731 475
rect 2199 475 2203 479
rect 2287 475 2291 479
rect 2383 475 2387 479
rect 2495 475 2499 479
rect 2639 475 2643 479
rect 2815 475 2819 479
rect 3015 475 3019 479
rect 3223 475 3227 479
rect 3439 475 3443 479
rect 111 461 115 465
rect 1075 463 1079 467
rect 1823 461 1827 465
rect 2347 463 2351 467
rect 111 444 115 448
rect 543 447 547 451
rect 699 447 703 451
rect 1431 447 1435 451
rect 1823 444 1827 448
rect 2219 443 2223 447
rect 2391 443 2395 447
rect 3499 443 3503 447
rect 167 431 171 435
rect 319 431 323 435
rect 471 431 475 435
rect 623 431 627 435
rect 767 431 771 435
rect 895 431 899 435
rect 1015 431 1019 435
rect 1135 431 1139 435
rect 1247 431 1251 435
rect 1351 431 1355 435
rect 1447 431 1451 435
rect 1551 431 1555 435
rect 1647 431 1651 435
rect 1735 431 1739 435
rect 1895 433 1899 437
rect 2039 433 2043 437
rect 2207 433 2211 437
rect 2383 433 2387 437
rect 2575 433 2579 437
rect 2783 433 2787 437
rect 3007 433 3011 437
rect 3239 433 3243 437
rect 3471 433 3475 437
rect 331 419 335 423
rect 699 419 703 423
rect 783 419 787 423
rect 903 419 907 423
rect 1143 419 1147 423
rect 1455 419 1459 423
rect 1863 420 1867 424
rect 3575 420 3579 424
rect 159 407 163 411
rect 543 407 544 411
rect 544 407 547 411
rect 647 407 651 411
rect 1083 407 1087 411
rect 1431 407 1432 411
rect 1432 407 1435 411
rect 1863 403 1867 407
rect 3179 403 3183 407
rect 3471 403 3475 407
rect 3575 403 3579 407
rect 151 397 155 401
rect 271 397 275 401
rect 407 397 411 401
rect 551 397 555 401
rect 711 397 715 401
rect 887 397 891 401
rect 1063 397 1067 401
rect 1247 397 1251 401
rect 1439 397 1443 401
rect 1639 397 1643 401
rect 1887 393 1891 397
rect 2031 393 2035 397
rect 2199 393 2203 397
rect 2375 393 2379 397
rect 2567 393 2571 397
rect 2775 393 2779 397
rect 2999 393 3003 397
rect 3231 393 3235 397
rect 3463 393 3467 397
rect 111 384 115 388
rect 331 383 335 387
rect 339 379 343 383
rect 647 383 651 387
rect 1163 379 1167 383
rect 1823 384 1827 388
rect 1903 379 1907 383
rect 111 367 115 371
rect 855 367 859 371
rect 1823 367 1827 371
rect 1887 371 1891 375
rect 1975 371 1979 375
rect 2063 371 2067 375
rect 2151 371 2155 375
rect 2263 371 2267 375
rect 2383 371 2387 375
rect 2519 371 2523 375
rect 2671 371 2675 375
rect 2847 371 2851 375
rect 3031 371 3035 375
rect 3231 371 3235 375
rect 3431 371 3435 375
rect 143 357 147 361
rect 263 357 267 361
rect 399 357 403 361
rect 543 357 547 361
rect 703 357 707 361
rect 879 357 883 361
rect 1055 357 1059 361
rect 1239 357 1243 361
rect 1431 357 1435 361
rect 1631 357 1635 361
rect 1863 361 1867 365
rect 2219 363 2223 367
rect 3575 361 3579 365
rect 1863 344 1867 348
rect 2451 347 2455 351
rect 3151 347 3155 351
rect 3159 347 3163 351
rect 3575 344 3579 348
rect 1895 331 1899 335
rect 1983 331 1987 335
rect 2071 331 2075 335
rect 2159 331 2163 335
rect 2271 331 2275 335
rect 2391 331 2395 335
rect 2527 331 2531 335
rect 2679 331 2683 335
rect 2855 331 2859 335
rect 3039 331 3043 335
rect 3239 331 3243 335
rect 3439 331 3443 335
rect 135 319 139 323
rect 223 319 227 323
rect 311 319 315 323
rect 399 319 403 323
rect 487 319 491 323
rect 575 319 579 323
rect 663 319 667 323
rect 751 319 755 323
rect 839 319 843 323
rect 927 319 931 323
rect 1015 319 1019 323
rect 1103 319 1107 323
rect 1191 319 1195 323
rect 1287 319 1291 323
rect 1383 319 1387 323
rect 1479 319 1483 323
rect 1575 319 1579 323
rect 1671 319 1675 323
rect 2451 319 2455 323
rect 2535 319 2539 323
rect 2687 319 2691 323
rect 3151 319 3155 323
rect 3427 319 3431 323
rect 111 309 115 313
rect 731 311 735 315
rect 1083 311 1087 315
rect 1823 309 1827 313
rect 1903 307 1907 311
rect 2367 307 2371 311
rect 2603 307 2607 311
rect 2703 307 2707 311
rect 111 292 115 296
rect 819 295 823 299
rect 1083 295 1087 299
rect 1171 295 1175 299
rect 1563 295 1567 299
rect 1643 295 1647 299
rect 1895 297 1899 301
rect 1983 297 1987 301
rect 2071 297 2075 301
rect 2159 297 2163 301
rect 2247 297 2251 301
rect 2359 297 2363 301
rect 2471 297 2475 301
rect 2583 297 2587 301
rect 2695 297 2699 301
rect 2807 297 2811 301
rect 2919 297 2923 301
rect 3039 297 3043 301
rect 3159 297 3163 301
rect 1823 292 1827 296
rect 1863 284 1867 288
rect 143 279 147 283
rect 231 279 235 283
rect 319 279 323 283
rect 407 279 411 283
rect 495 279 499 283
rect 583 279 587 283
rect 671 279 675 283
rect 759 279 763 283
rect 847 279 851 283
rect 935 279 939 283
rect 1023 279 1027 283
rect 1111 279 1115 283
rect 1199 279 1203 283
rect 1295 279 1299 283
rect 1391 279 1395 283
rect 1487 279 1491 283
rect 1583 279 1587 283
rect 1679 279 1683 283
rect 2535 283 2539 287
rect 2543 279 2547 283
rect 3575 284 3579 288
rect 135 267 136 271
rect 136 267 139 271
rect 819 267 823 271
rect 855 267 859 271
rect 731 259 735 263
rect 739 259 743 263
rect 1171 267 1175 271
rect 1191 267 1192 271
rect 1192 267 1195 271
rect 1303 267 1307 271
rect 1643 267 1647 271
rect 1863 267 1867 271
rect 2227 267 2231 271
rect 3107 267 3111 271
rect 3575 267 3579 271
rect 1083 259 1087 263
rect 1887 257 1891 261
rect 1975 257 1979 261
rect 2063 257 2067 261
rect 2151 257 2155 261
rect 2239 257 2243 261
rect 2351 257 2355 261
rect 2463 257 2467 261
rect 2575 257 2579 261
rect 2687 257 2691 261
rect 2799 257 2803 261
rect 2911 257 2915 261
rect 3031 257 3035 261
rect 3151 257 3155 261
rect 211 251 215 255
rect 299 251 303 255
rect 387 251 391 255
rect 475 251 479 255
rect 563 251 567 255
rect 651 251 655 255
rect 735 251 739 255
rect 1031 251 1035 255
rect 1355 251 1359 255
rect 1443 251 1447 255
rect 1535 251 1539 255
rect 1707 251 1711 255
rect 143 241 147 245
rect 231 241 235 245
rect 319 241 323 245
rect 407 241 411 245
rect 495 241 499 245
rect 583 241 587 245
rect 671 241 675 245
rect 759 241 763 245
rect 847 241 851 245
rect 935 241 939 245
rect 1023 241 1027 245
rect 1111 241 1115 245
rect 1199 241 1203 245
rect 1287 241 1291 245
rect 1375 241 1379 245
rect 1463 241 1467 245
rect 1551 241 1555 245
rect 1639 241 1643 245
rect 1727 241 1731 245
rect 1887 235 1891 239
rect 1975 235 1979 239
rect 2063 235 2067 239
rect 2151 235 2155 239
rect 2263 235 2267 239
rect 2399 235 2403 239
rect 2535 235 2539 239
rect 2679 235 2683 239
rect 2815 235 2819 239
rect 2951 235 2955 239
rect 3087 235 3091 239
rect 3223 235 3227 239
rect 3359 235 3363 239
rect 3479 235 3483 239
rect 111 228 115 232
rect 135 223 139 227
rect 211 223 215 227
rect 299 223 303 227
rect 387 223 391 227
rect 475 223 479 227
rect 563 223 567 227
rect 651 223 655 227
rect 1191 223 1195 227
rect 1267 223 1271 227
rect 1355 223 1359 227
rect 1443 223 1447 227
rect 1823 228 1827 232
rect 1863 225 1867 229
rect 2603 227 2607 231
rect 3191 227 3195 231
rect 3427 227 3431 231
rect 3575 225 3579 229
rect 111 211 115 215
rect 1707 211 1711 215
rect 1727 211 1731 215
rect 1823 211 1827 215
rect 1863 208 1867 212
rect 3575 208 3579 212
rect 135 201 139 205
rect 223 201 227 205
rect 311 201 315 205
rect 399 201 403 205
rect 487 201 491 205
rect 575 201 579 205
rect 663 201 667 205
rect 751 201 755 205
rect 839 201 843 205
rect 927 201 931 205
rect 1015 201 1019 205
rect 1103 201 1107 205
rect 1191 201 1195 205
rect 1279 201 1283 205
rect 1367 201 1371 205
rect 1455 201 1459 205
rect 1543 201 1547 205
rect 1631 201 1635 205
rect 1719 201 1723 205
rect 1535 195 1539 199
rect 1727 195 1731 199
rect 1895 195 1899 199
rect 1983 195 1987 199
rect 2071 195 2075 199
rect 2159 195 2163 199
rect 2271 195 2275 199
rect 2407 195 2411 199
rect 2543 195 2547 199
rect 2687 195 2691 199
rect 2823 195 2827 199
rect 2959 195 2963 199
rect 3095 195 3099 199
rect 3231 195 3235 199
rect 3367 195 3371 199
rect 3487 195 3491 199
rect 1903 183 1907 187
rect 2831 183 2835 187
rect 3375 183 3379 187
rect 3471 183 3475 187
rect 2791 139 2795 143
rect 3459 139 3463 143
rect 2783 129 2787 133
rect 2871 129 2875 133
rect 2959 129 2963 133
rect 3047 129 3051 133
rect 3135 129 3139 133
rect 3223 129 3227 133
rect 3311 129 3315 133
rect 3399 129 3403 133
rect 3487 129 3491 133
rect 1863 116 1867 120
rect 3375 115 3379 119
rect 3459 115 3463 119
rect 3575 116 3579 120
rect 1863 99 1867 103
rect 3575 99 3579 103
rect 2775 89 2779 93
rect 2863 89 2867 93
rect 2951 89 2955 93
rect 3039 89 3043 93
rect 3127 89 3131 93
rect 3215 89 3219 93
rect 3303 89 3307 93
rect 3391 89 3395 93
rect 3479 89 3483 93
<< m3 >>
rect 111 3670 115 3671
rect 111 3665 115 3666
rect 135 3670 139 3671
rect 135 3665 139 3666
rect 223 3670 227 3671
rect 223 3665 227 3666
rect 1823 3670 1827 3671
rect 1823 3665 1827 3666
rect 112 3650 114 3665
rect 136 3660 138 3665
rect 224 3660 226 3665
rect 134 3659 140 3660
rect 134 3655 135 3659
rect 139 3655 140 3659
rect 134 3654 140 3655
rect 222 3659 228 3660
rect 222 3655 223 3659
rect 227 3655 228 3659
rect 222 3654 228 3655
rect 202 3651 208 3652
rect 110 3649 116 3650
rect 110 3645 111 3649
rect 115 3645 116 3649
rect 202 3647 203 3651
rect 207 3647 208 3651
rect 1824 3650 1826 3665
rect 202 3646 208 3647
rect 1822 3649 1828 3650
rect 110 3644 116 3645
rect 110 3632 116 3633
rect 110 3628 111 3632
rect 115 3628 116 3632
rect 110 3627 116 3628
rect 112 3603 114 3627
rect 142 3619 148 3620
rect 142 3615 143 3619
rect 147 3615 148 3619
rect 142 3614 148 3615
rect 144 3603 146 3614
rect 111 3602 115 3603
rect 111 3597 115 3598
rect 143 3602 147 3603
rect 143 3597 147 3598
rect 112 3573 114 3597
rect 144 3586 146 3597
rect 204 3596 206 3646
rect 1822 3645 1823 3649
rect 1827 3645 1828 3649
rect 1822 3644 1828 3645
rect 1822 3632 1828 3633
rect 1822 3628 1823 3632
rect 1827 3628 1828 3632
rect 1822 3627 1828 3628
rect 230 3619 236 3620
rect 230 3615 231 3619
rect 235 3615 236 3619
rect 230 3614 236 3615
rect 232 3603 234 3614
rect 1824 3603 1826 3627
rect 231 3602 235 3603
rect 231 3597 235 3598
rect 319 3602 323 3603
rect 319 3597 323 3598
rect 407 3602 411 3603
rect 407 3597 411 3598
rect 495 3602 499 3603
rect 495 3597 499 3598
rect 1823 3602 1827 3603
rect 1823 3597 1827 3598
rect 198 3595 206 3596
rect 198 3591 199 3595
rect 203 3593 206 3595
rect 203 3591 204 3593
rect 198 3590 204 3591
rect 232 3586 234 3597
rect 320 3586 322 3597
rect 408 3586 410 3597
rect 496 3586 498 3597
rect 142 3585 148 3586
rect 142 3581 143 3585
rect 147 3581 148 3585
rect 142 3580 148 3581
rect 230 3585 236 3586
rect 230 3581 231 3585
rect 235 3581 236 3585
rect 230 3580 236 3581
rect 318 3585 324 3586
rect 318 3581 319 3585
rect 323 3581 324 3585
rect 318 3580 324 3581
rect 406 3585 412 3586
rect 406 3581 407 3585
rect 411 3581 412 3585
rect 406 3580 412 3581
rect 494 3585 500 3586
rect 494 3581 495 3585
rect 499 3581 500 3585
rect 494 3580 500 3581
rect 1824 3573 1826 3597
rect 1863 3594 1867 3595
rect 1863 3589 1867 3590
rect 1887 3594 1891 3595
rect 1887 3589 1891 3590
rect 1975 3594 1979 3595
rect 1975 3589 1979 3590
rect 2063 3594 2067 3595
rect 2063 3589 2067 3590
rect 2151 3594 2155 3595
rect 2151 3589 2155 3590
rect 2239 3594 2243 3595
rect 2239 3589 2243 3590
rect 2327 3594 2331 3595
rect 2327 3589 2331 3590
rect 2431 3594 2435 3595
rect 2431 3589 2435 3590
rect 2535 3594 2539 3595
rect 2535 3589 2539 3590
rect 2631 3594 2635 3595
rect 2631 3589 2635 3590
rect 2727 3594 2731 3595
rect 2727 3589 2731 3590
rect 2823 3594 2827 3595
rect 2823 3589 2827 3590
rect 2919 3594 2923 3595
rect 2919 3589 2923 3590
rect 3015 3594 3019 3595
rect 3015 3589 3019 3590
rect 3119 3594 3123 3595
rect 3119 3589 3123 3590
rect 3223 3594 3227 3595
rect 3223 3589 3227 3590
rect 3575 3594 3579 3595
rect 3575 3589 3579 3590
rect 1864 3574 1866 3589
rect 1888 3584 1890 3589
rect 1976 3584 1978 3589
rect 2064 3584 2066 3589
rect 2152 3584 2154 3589
rect 2240 3584 2242 3589
rect 2328 3584 2330 3589
rect 2432 3584 2434 3589
rect 2536 3584 2538 3589
rect 2632 3584 2634 3589
rect 2728 3584 2730 3589
rect 2824 3584 2826 3589
rect 2920 3584 2922 3589
rect 3016 3584 3018 3589
rect 3120 3584 3122 3589
rect 3224 3584 3226 3589
rect 1886 3583 1892 3584
rect 1886 3579 1887 3583
rect 1891 3579 1892 3583
rect 1886 3578 1892 3579
rect 1974 3583 1980 3584
rect 1974 3579 1975 3583
rect 1979 3579 1980 3583
rect 1974 3578 1980 3579
rect 2062 3583 2068 3584
rect 2062 3579 2063 3583
rect 2067 3579 2068 3583
rect 2062 3578 2068 3579
rect 2150 3583 2156 3584
rect 2150 3579 2151 3583
rect 2155 3579 2156 3583
rect 2150 3578 2156 3579
rect 2238 3583 2244 3584
rect 2238 3579 2239 3583
rect 2243 3579 2244 3583
rect 2238 3578 2244 3579
rect 2326 3583 2332 3584
rect 2326 3579 2327 3583
rect 2331 3579 2332 3583
rect 2326 3578 2332 3579
rect 2430 3583 2436 3584
rect 2430 3579 2431 3583
rect 2435 3579 2436 3583
rect 2430 3578 2436 3579
rect 2534 3583 2540 3584
rect 2534 3579 2535 3583
rect 2539 3579 2540 3583
rect 2534 3578 2540 3579
rect 2630 3583 2636 3584
rect 2630 3579 2631 3583
rect 2635 3579 2636 3583
rect 2630 3578 2636 3579
rect 2726 3583 2732 3584
rect 2726 3579 2727 3583
rect 2731 3579 2732 3583
rect 2726 3578 2732 3579
rect 2822 3583 2828 3584
rect 2822 3579 2823 3583
rect 2827 3579 2828 3583
rect 2822 3578 2828 3579
rect 2918 3583 2924 3584
rect 2918 3579 2919 3583
rect 2923 3579 2924 3583
rect 2918 3578 2924 3579
rect 3014 3583 3020 3584
rect 3014 3579 3015 3583
rect 3019 3579 3020 3583
rect 3014 3578 3020 3579
rect 3118 3583 3124 3584
rect 3118 3579 3119 3583
rect 3123 3579 3124 3583
rect 3118 3578 3124 3579
rect 3222 3583 3228 3584
rect 3222 3579 3223 3583
rect 3227 3579 3228 3583
rect 3222 3578 3228 3579
rect 2498 3575 2504 3576
rect 1862 3573 1868 3574
rect 110 3572 116 3573
rect 110 3568 111 3572
rect 115 3568 116 3572
rect 110 3567 116 3568
rect 1822 3572 1828 3573
rect 1822 3568 1823 3572
rect 1827 3568 1828 3572
rect 1862 3569 1863 3573
rect 1867 3569 1868 3573
rect 2498 3571 2499 3575
rect 2503 3571 2504 3575
rect 3576 3574 3578 3589
rect 2498 3570 2504 3571
rect 3574 3573 3580 3574
rect 1862 3568 1868 3569
rect 1822 3567 1828 3568
rect 2500 3557 2502 3570
rect 3574 3569 3575 3573
rect 3579 3569 3580 3573
rect 3574 3568 3580 3569
rect 3186 3559 3192 3560
rect 1862 3556 1868 3557
rect 110 3555 116 3556
rect 110 3551 111 3555
rect 115 3551 116 3555
rect 110 3550 116 3551
rect 1822 3555 1828 3556
rect 1822 3551 1823 3555
rect 1827 3551 1828 3555
rect 1862 3552 1863 3556
rect 1867 3552 1868 3556
rect 1862 3551 1868 3552
rect 2111 3556 2115 3557
rect 2111 3551 2115 3552
rect 2499 3556 2503 3557
rect 3186 3555 3187 3559
rect 3191 3555 3192 3559
rect 3186 3554 3192 3555
rect 3214 3559 3220 3560
rect 3214 3555 3215 3559
rect 3219 3555 3220 3559
rect 3214 3554 3220 3555
rect 3574 3556 3580 3557
rect 2499 3551 2503 3552
rect 1822 3550 1828 3551
rect 112 3535 114 3550
rect 134 3545 140 3546
rect 134 3541 135 3545
rect 139 3541 140 3545
rect 134 3540 140 3541
rect 222 3545 228 3546
rect 222 3541 223 3545
rect 227 3541 228 3545
rect 222 3540 228 3541
rect 310 3545 316 3546
rect 310 3541 311 3545
rect 315 3541 316 3545
rect 310 3540 316 3541
rect 398 3545 404 3546
rect 398 3541 399 3545
rect 403 3541 404 3545
rect 398 3540 404 3541
rect 486 3545 492 3546
rect 486 3541 487 3545
rect 491 3541 492 3545
rect 486 3540 492 3541
rect 136 3535 138 3540
rect 224 3535 226 3540
rect 266 3539 272 3540
rect 266 3535 267 3539
rect 271 3535 272 3539
rect 312 3535 314 3540
rect 400 3535 402 3540
rect 488 3535 490 3540
rect 1824 3535 1826 3550
rect 111 3534 115 3535
rect 111 3529 115 3530
rect 135 3534 139 3535
rect 135 3529 139 3530
rect 223 3534 227 3535
rect 223 3529 227 3530
rect 247 3534 251 3535
rect 266 3534 272 3535
rect 311 3534 315 3535
rect 247 3529 251 3530
rect 112 3514 114 3529
rect 248 3524 250 3529
rect 246 3523 252 3524
rect 246 3519 247 3523
rect 251 3519 252 3523
rect 246 3518 252 3519
rect 110 3513 116 3514
rect 110 3509 111 3513
rect 115 3509 116 3513
rect 110 3508 116 3509
rect 110 3496 116 3497
rect 110 3492 111 3496
rect 115 3492 116 3496
rect 110 3491 116 3492
rect 112 3467 114 3491
rect 254 3483 260 3484
rect 254 3479 255 3483
rect 259 3479 260 3483
rect 254 3478 260 3479
rect 256 3467 258 3478
rect 268 3472 270 3534
rect 311 3529 315 3530
rect 375 3534 379 3535
rect 375 3529 379 3530
rect 399 3534 403 3535
rect 399 3529 403 3530
rect 487 3534 491 3535
rect 487 3529 491 3530
rect 503 3534 507 3535
rect 503 3529 507 3530
rect 623 3534 627 3535
rect 623 3529 627 3530
rect 743 3534 747 3535
rect 743 3529 747 3530
rect 863 3534 867 3535
rect 863 3529 867 3530
rect 975 3534 979 3535
rect 975 3529 979 3530
rect 1079 3534 1083 3535
rect 1079 3529 1083 3530
rect 1175 3534 1179 3535
rect 1175 3529 1179 3530
rect 1271 3534 1275 3535
rect 1271 3529 1275 3530
rect 1367 3534 1371 3535
rect 1367 3529 1371 3530
rect 1471 3534 1475 3535
rect 1471 3529 1475 3530
rect 1575 3534 1579 3535
rect 1575 3529 1579 3530
rect 1823 3534 1827 3535
rect 1823 3529 1827 3530
rect 376 3524 378 3529
rect 504 3524 506 3529
rect 624 3524 626 3529
rect 744 3524 746 3529
rect 864 3524 866 3529
rect 976 3524 978 3529
rect 1080 3524 1082 3529
rect 1176 3524 1178 3529
rect 1272 3524 1274 3529
rect 1368 3524 1370 3529
rect 1472 3524 1474 3529
rect 1576 3524 1578 3529
rect 374 3523 380 3524
rect 374 3519 375 3523
rect 379 3519 380 3523
rect 374 3518 380 3519
rect 502 3523 508 3524
rect 502 3519 503 3523
rect 507 3519 508 3523
rect 502 3518 508 3519
rect 622 3523 628 3524
rect 622 3519 623 3523
rect 627 3519 628 3523
rect 622 3518 628 3519
rect 742 3523 748 3524
rect 742 3519 743 3523
rect 747 3519 748 3523
rect 742 3518 748 3519
rect 862 3523 868 3524
rect 862 3519 863 3523
rect 867 3519 868 3523
rect 862 3518 868 3519
rect 974 3523 980 3524
rect 974 3519 975 3523
rect 979 3519 980 3523
rect 974 3518 980 3519
rect 1078 3523 1084 3524
rect 1078 3519 1079 3523
rect 1083 3519 1084 3523
rect 1078 3518 1084 3519
rect 1174 3523 1180 3524
rect 1174 3519 1175 3523
rect 1179 3519 1180 3523
rect 1174 3518 1180 3519
rect 1270 3523 1276 3524
rect 1270 3519 1271 3523
rect 1275 3519 1276 3523
rect 1270 3518 1276 3519
rect 1366 3523 1372 3524
rect 1366 3519 1367 3523
rect 1371 3519 1372 3523
rect 1366 3518 1372 3519
rect 1470 3523 1476 3524
rect 1470 3519 1471 3523
rect 1475 3519 1476 3523
rect 1470 3518 1476 3519
rect 1574 3523 1580 3524
rect 1574 3519 1575 3523
rect 1579 3519 1580 3523
rect 1574 3518 1580 3519
rect 1538 3515 1544 3516
rect 1538 3511 1539 3515
rect 1543 3511 1544 3515
rect 1824 3514 1826 3529
rect 1864 3527 1866 3551
rect 1894 3543 1900 3544
rect 1894 3539 1895 3543
rect 1899 3539 1900 3543
rect 1894 3538 1900 3539
rect 1982 3543 1988 3544
rect 1982 3539 1983 3543
rect 1987 3539 1988 3543
rect 1982 3538 1988 3539
rect 2070 3543 2076 3544
rect 2070 3539 2071 3543
rect 2075 3539 2076 3543
rect 2070 3538 2076 3539
rect 1886 3531 1892 3532
rect 1886 3527 1887 3531
rect 1891 3527 1892 3531
rect 1896 3527 1898 3538
rect 1984 3527 1986 3538
rect 2072 3527 2074 3538
rect 1863 3526 1867 3527
rect 1886 3526 1892 3527
rect 1895 3526 1899 3527
rect 1863 3521 1867 3522
rect 1538 3510 1544 3511
rect 1822 3513 1828 3514
rect 570 3499 576 3500
rect 570 3495 571 3499
rect 575 3495 576 3499
rect 570 3494 576 3495
rect 734 3499 740 3500
rect 734 3495 735 3499
rect 739 3495 740 3499
rect 734 3494 740 3495
rect 966 3499 972 3500
rect 966 3495 967 3499
rect 971 3495 972 3499
rect 966 3494 972 3495
rect 382 3483 388 3484
rect 382 3479 383 3483
rect 387 3479 388 3483
rect 382 3478 388 3479
rect 510 3483 516 3484
rect 510 3479 511 3483
rect 515 3479 516 3483
rect 510 3478 516 3479
rect 266 3471 272 3472
rect 266 3467 267 3471
rect 271 3467 272 3471
rect 384 3467 386 3478
rect 512 3467 514 3478
rect 572 3476 574 3494
rect 630 3483 636 3484
rect 630 3479 631 3483
rect 635 3479 636 3483
rect 630 3478 636 3479
rect 570 3475 576 3476
rect 570 3471 571 3475
rect 575 3471 576 3475
rect 570 3470 576 3471
rect 632 3467 634 3478
rect 111 3466 115 3467
rect 111 3461 115 3462
rect 175 3466 179 3467
rect 175 3461 179 3462
rect 255 3466 259 3467
rect 266 3466 272 3467
rect 303 3466 307 3467
rect 255 3461 259 3462
rect 303 3461 307 3462
rect 383 3466 387 3467
rect 383 3461 387 3462
rect 447 3466 451 3467
rect 447 3461 451 3462
rect 511 3466 515 3467
rect 511 3461 515 3462
rect 591 3466 595 3467
rect 591 3461 595 3462
rect 631 3466 635 3467
rect 631 3461 635 3462
rect 650 3463 656 3464
rect 112 3437 114 3461
rect 176 3450 178 3461
rect 242 3459 248 3460
rect 242 3455 243 3459
rect 247 3455 248 3459
rect 242 3454 248 3455
rect 174 3449 180 3450
rect 174 3445 175 3449
rect 179 3445 180 3449
rect 174 3444 180 3445
rect 110 3436 116 3437
rect 110 3432 111 3436
rect 115 3432 116 3436
rect 244 3432 246 3454
rect 304 3450 306 3461
rect 370 3459 376 3460
rect 370 3455 371 3459
rect 375 3455 376 3459
rect 370 3454 376 3455
rect 302 3449 308 3450
rect 302 3445 303 3449
rect 307 3445 308 3449
rect 302 3444 308 3445
rect 372 3432 374 3454
rect 448 3450 450 3461
rect 592 3450 594 3461
rect 650 3459 651 3463
rect 655 3459 656 3463
rect 736 3460 738 3494
rect 750 3483 756 3484
rect 750 3479 751 3483
rect 755 3479 756 3483
rect 750 3478 756 3479
rect 870 3483 876 3484
rect 870 3479 871 3483
rect 875 3479 876 3483
rect 870 3478 876 3479
rect 752 3467 754 3478
rect 872 3467 874 3478
rect 968 3472 970 3494
rect 982 3483 988 3484
rect 982 3479 983 3483
rect 987 3479 988 3483
rect 982 3478 988 3479
rect 1086 3483 1092 3484
rect 1086 3479 1087 3483
rect 1091 3479 1092 3483
rect 1086 3478 1092 3479
rect 1182 3483 1188 3484
rect 1182 3479 1183 3483
rect 1187 3479 1188 3483
rect 1182 3478 1188 3479
rect 1278 3483 1284 3484
rect 1278 3479 1279 3483
rect 1283 3479 1284 3483
rect 1278 3478 1284 3479
rect 1374 3483 1380 3484
rect 1374 3479 1375 3483
rect 1379 3479 1380 3483
rect 1374 3478 1380 3479
rect 1478 3483 1484 3484
rect 1478 3479 1479 3483
rect 1483 3479 1484 3483
rect 1478 3478 1484 3479
rect 966 3471 972 3472
rect 966 3467 967 3471
rect 971 3467 972 3471
rect 984 3467 986 3478
rect 1088 3467 1090 3478
rect 1184 3467 1186 3478
rect 1280 3467 1282 3478
rect 1376 3467 1378 3478
rect 1480 3467 1482 3478
rect 743 3466 747 3467
rect 743 3461 747 3462
rect 751 3466 755 3467
rect 751 3461 755 3462
rect 871 3466 875 3467
rect 871 3461 875 3462
rect 895 3466 899 3467
rect 966 3466 972 3467
rect 983 3466 987 3467
rect 895 3461 899 3462
rect 983 3461 987 3462
rect 1039 3466 1043 3467
rect 1039 3461 1043 3462
rect 1087 3466 1091 3467
rect 1087 3461 1091 3462
rect 1183 3466 1187 3467
rect 1183 3461 1187 3462
rect 1279 3466 1283 3467
rect 1279 3461 1283 3462
rect 1327 3466 1331 3467
rect 1327 3461 1331 3462
rect 1375 3466 1379 3467
rect 1375 3461 1379 3462
rect 1479 3466 1483 3467
rect 1479 3461 1483 3462
rect 650 3458 656 3459
rect 734 3459 740 3460
rect 446 3449 452 3450
rect 446 3445 447 3449
rect 451 3445 452 3449
rect 446 3444 452 3445
rect 590 3449 596 3450
rect 590 3445 591 3449
rect 595 3445 596 3449
rect 590 3444 596 3445
rect 652 3436 654 3458
rect 682 3455 688 3456
rect 682 3451 683 3455
rect 687 3451 688 3455
rect 734 3455 735 3459
rect 739 3455 740 3459
rect 734 3454 740 3455
rect 682 3450 688 3451
rect 744 3450 746 3461
rect 896 3450 898 3461
rect 962 3459 968 3460
rect 962 3455 963 3459
rect 967 3455 968 3459
rect 962 3454 968 3455
rect 650 3435 656 3436
rect 110 3431 116 3432
rect 242 3431 248 3432
rect 242 3427 243 3431
rect 247 3427 248 3431
rect 242 3426 248 3427
rect 370 3431 376 3432
rect 370 3427 371 3431
rect 375 3427 376 3431
rect 650 3431 651 3435
rect 655 3431 656 3435
rect 684 3432 686 3450
rect 742 3449 748 3450
rect 742 3445 743 3449
rect 747 3445 748 3449
rect 742 3444 748 3445
rect 894 3449 900 3450
rect 894 3445 895 3449
rect 899 3445 900 3449
rect 894 3444 900 3445
rect 964 3432 966 3454
rect 1040 3450 1042 3461
rect 1184 3450 1186 3461
rect 1250 3459 1256 3460
rect 1250 3455 1251 3459
rect 1255 3455 1256 3459
rect 1250 3454 1256 3455
rect 1038 3449 1044 3450
rect 1038 3445 1039 3449
rect 1043 3445 1044 3449
rect 1038 3444 1044 3445
rect 1182 3449 1188 3450
rect 1182 3445 1183 3449
rect 1187 3445 1188 3449
rect 1182 3444 1188 3445
rect 1252 3432 1254 3454
rect 1328 3450 1330 3461
rect 1438 3459 1444 3460
rect 1438 3455 1439 3459
rect 1443 3455 1444 3459
rect 1438 3454 1444 3455
rect 1326 3449 1332 3450
rect 1326 3445 1327 3449
rect 1331 3445 1332 3449
rect 1326 3444 1332 3445
rect 1440 3437 1442 3454
rect 1480 3450 1482 3461
rect 1540 3460 1542 3510
rect 1822 3509 1823 3513
rect 1827 3509 1828 3513
rect 1822 3508 1828 3509
rect 1864 3497 1866 3521
rect 1822 3496 1828 3497
rect 1822 3492 1823 3496
rect 1827 3492 1828 3496
rect 1822 3491 1828 3492
rect 1862 3496 1868 3497
rect 1862 3492 1863 3496
rect 1867 3492 1868 3496
rect 1888 3492 1890 3526
rect 1895 3521 1899 3522
rect 1983 3526 1987 3527
rect 1983 3521 1987 3522
rect 2071 3526 2075 3527
rect 2071 3521 2075 3522
rect 2103 3526 2107 3527
rect 2103 3521 2107 3522
rect 1896 3510 1898 3521
rect 1962 3519 1968 3520
rect 1962 3515 1963 3519
rect 1967 3515 1968 3519
rect 1962 3514 1968 3515
rect 1894 3509 1900 3510
rect 1894 3505 1895 3509
rect 1899 3505 1900 3509
rect 1894 3504 1900 3505
rect 1964 3492 1966 3514
rect 1984 3510 1986 3521
rect 1990 3519 1996 3520
rect 1990 3515 1991 3519
rect 1995 3515 1996 3519
rect 1990 3514 1996 3515
rect 1982 3509 1988 3510
rect 1982 3505 1983 3509
rect 1987 3505 1988 3509
rect 1982 3504 1988 3505
rect 1862 3491 1868 3492
rect 1886 3491 1892 3492
rect 1582 3483 1588 3484
rect 1582 3479 1583 3483
rect 1587 3479 1588 3483
rect 1582 3478 1588 3479
rect 1584 3467 1586 3478
rect 1824 3467 1826 3491
rect 1886 3487 1887 3491
rect 1891 3487 1892 3491
rect 1886 3486 1892 3487
rect 1962 3491 1968 3492
rect 1962 3487 1963 3491
rect 1967 3487 1968 3491
rect 1962 3486 1968 3487
rect 1862 3479 1868 3480
rect 1862 3475 1863 3479
rect 1867 3475 1868 3479
rect 1862 3474 1868 3475
rect 1583 3466 1587 3467
rect 1583 3461 1587 3462
rect 1823 3466 1827 3467
rect 1823 3461 1827 3462
rect 1538 3459 1544 3460
rect 1538 3455 1539 3459
rect 1543 3455 1544 3459
rect 1538 3454 1544 3455
rect 1478 3449 1484 3450
rect 1478 3445 1479 3449
rect 1483 3445 1484 3449
rect 1478 3444 1484 3445
rect 1824 3437 1826 3461
rect 1864 3451 1866 3474
rect 1886 3469 1892 3470
rect 1886 3465 1887 3469
rect 1891 3465 1892 3469
rect 1886 3464 1892 3465
rect 1974 3469 1980 3470
rect 1974 3465 1975 3469
rect 1979 3465 1980 3469
rect 1974 3464 1980 3465
rect 1888 3451 1890 3464
rect 1976 3451 1978 3464
rect 1863 3450 1867 3451
rect 1863 3445 1867 3446
rect 1887 3450 1891 3451
rect 1887 3445 1891 3446
rect 1975 3450 1979 3451
rect 1975 3445 1979 3446
rect 1439 3436 1443 3437
rect 1471 3436 1475 3437
rect 1822 3436 1828 3437
rect 1822 3432 1823 3436
rect 1827 3432 1828 3436
rect 650 3430 656 3431
rect 682 3431 688 3432
rect 370 3426 376 3427
rect 682 3427 683 3431
rect 687 3427 688 3431
rect 682 3426 688 3427
rect 962 3431 968 3432
rect 962 3427 963 3431
rect 967 3427 968 3431
rect 962 3426 968 3427
rect 1250 3431 1256 3432
rect 1439 3431 1443 3432
rect 1470 3431 1476 3432
rect 1822 3431 1828 3432
rect 1250 3427 1251 3431
rect 1255 3427 1256 3431
rect 1250 3426 1256 3427
rect 1470 3427 1471 3431
rect 1475 3427 1476 3431
rect 1864 3430 1866 3445
rect 1888 3440 1890 3445
rect 1886 3439 1892 3440
rect 1886 3435 1887 3439
rect 1891 3435 1892 3439
rect 1886 3434 1892 3435
rect 1992 3432 1994 3514
rect 2104 3510 2106 3521
rect 2112 3520 2114 3551
rect 2158 3543 2164 3544
rect 2158 3539 2159 3543
rect 2163 3539 2164 3543
rect 2158 3538 2164 3539
rect 2246 3543 2252 3544
rect 2246 3539 2247 3543
rect 2251 3539 2252 3543
rect 2246 3538 2252 3539
rect 2334 3543 2340 3544
rect 2334 3539 2335 3543
rect 2339 3539 2340 3543
rect 2334 3538 2340 3539
rect 2438 3543 2444 3544
rect 2438 3539 2439 3543
rect 2443 3539 2444 3543
rect 2438 3538 2444 3539
rect 2542 3543 2548 3544
rect 2542 3539 2543 3543
rect 2547 3539 2548 3543
rect 2542 3538 2548 3539
rect 2638 3543 2644 3544
rect 2638 3539 2639 3543
rect 2643 3539 2644 3543
rect 2638 3538 2644 3539
rect 2734 3543 2740 3544
rect 2734 3539 2735 3543
rect 2739 3539 2740 3543
rect 2734 3538 2740 3539
rect 2830 3543 2836 3544
rect 2830 3539 2831 3543
rect 2835 3539 2836 3543
rect 2830 3538 2836 3539
rect 2926 3543 2932 3544
rect 2926 3539 2927 3543
rect 2931 3539 2932 3543
rect 2926 3538 2932 3539
rect 3022 3543 3028 3544
rect 3022 3539 3023 3543
rect 3027 3539 3028 3543
rect 3022 3538 3028 3539
rect 3126 3543 3132 3544
rect 3126 3539 3127 3543
rect 3131 3539 3132 3543
rect 3126 3538 3132 3539
rect 2160 3527 2162 3538
rect 2248 3527 2250 3538
rect 2336 3527 2338 3538
rect 2440 3527 2442 3538
rect 2544 3527 2546 3538
rect 2640 3527 2642 3538
rect 2736 3527 2738 3538
rect 2832 3527 2834 3538
rect 2928 3527 2930 3538
rect 3024 3527 3026 3538
rect 3128 3527 3130 3538
rect 3188 3532 3190 3554
rect 3186 3531 3192 3532
rect 3186 3527 3187 3531
rect 3191 3527 3192 3531
rect 2159 3526 2163 3527
rect 2159 3521 2163 3522
rect 2231 3526 2235 3527
rect 2231 3521 2235 3522
rect 2247 3526 2251 3527
rect 2247 3521 2251 3522
rect 2335 3526 2339 3527
rect 2335 3521 2339 3522
rect 2367 3526 2371 3527
rect 2367 3521 2371 3522
rect 2439 3526 2443 3527
rect 2439 3521 2443 3522
rect 2511 3526 2515 3527
rect 2511 3521 2515 3522
rect 2543 3526 2547 3527
rect 2543 3521 2547 3522
rect 2639 3526 2643 3527
rect 2639 3521 2643 3522
rect 2655 3526 2659 3527
rect 2655 3521 2659 3522
rect 2735 3526 2739 3527
rect 2735 3521 2739 3522
rect 2791 3526 2795 3527
rect 2791 3521 2795 3522
rect 2831 3526 2835 3527
rect 2831 3521 2835 3522
rect 2927 3526 2931 3527
rect 2927 3521 2931 3522
rect 2935 3526 2939 3527
rect 2935 3521 2939 3522
rect 3023 3526 3027 3527
rect 3023 3521 3027 3522
rect 3079 3526 3083 3527
rect 3079 3521 3083 3522
rect 3127 3526 3131 3527
rect 3186 3526 3192 3527
rect 3127 3521 3131 3522
rect 2110 3519 2116 3520
rect 2110 3515 2111 3519
rect 2115 3515 2116 3519
rect 2110 3514 2116 3515
rect 2232 3510 2234 3521
rect 2290 3519 2296 3520
rect 2290 3515 2291 3519
rect 2295 3515 2296 3519
rect 2290 3514 2296 3515
rect 2102 3509 2108 3510
rect 2102 3505 2103 3509
rect 2107 3505 2108 3509
rect 2102 3504 2108 3505
rect 2230 3509 2236 3510
rect 2230 3505 2231 3509
rect 2235 3505 2236 3509
rect 2230 3504 2236 3505
rect 2292 3496 2294 3514
rect 2368 3510 2370 3521
rect 2512 3510 2514 3521
rect 2656 3510 2658 3521
rect 2722 3519 2728 3520
rect 2722 3515 2723 3519
rect 2727 3515 2728 3519
rect 2722 3514 2728 3515
rect 2366 3509 2372 3510
rect 2366 3505 2367 3509
rect 2371 3505 2372 3509
rect 2366 3504 2372 3505
rect 2510 3509 2516 3510
rect 2510 3505 2511 3509
rect 2515 3505 2516 3509
rect 2510 3504 2516 3505
rect 2654 3509 2660 3510
rect 2654 3505 2655 3509
rect 2659 3505 2660 3509
rect 2654 3504 2660 3505
rect 2290 3495 2296 3496
rect 2290 3491 2291 3495
rect 2295 3491 2296 3495
rect 2724 3492 2726 3514
rect 2792 3510 2794 3521
rect 2798 3519 2804 3520
rect 2798 3515 2799 3519
rect 2803 3515 2804 3519
rect 2798 3514 2804 3515
rect 2790 3509 2796 3510
rect 2790 3505 2791 3509
rect 2795 3505 2796 3509
rect 2790 3504 2796 3505
rect 2290 3490 2296 3491
rect 2722 3491 2728 3492
rect 2722 3487 2723 3491
rect 2727 3487 2728 3491
rect 2722 3486 2728 3487
rect 2094 3469 2100 3470
rect 2094 3465 2095 3469
rect 2099 3465 2100 3469
rect 2094 3464 2100 3465
rect 2222 3469 2228 3470
rect 2222 3465 2223 3469
rect 2227 3465 2228 3469
rect 2222 3464 2228 3465
rect 2358 3469 2364 3470
rect 2358 3465 2359 3469
rect 2363 3465 2364 3469
rect 2358 3464 2364 3465
rect 2502 3469 2508 3470
rect 2502 3465 2503 3469
rect 2507 3465 2508 3469
rect 2502 3464 2508 3465
rect 2646 3469 2652 3470
rect 2646 3465 2647 3469
rect 2651 3465 2652 3469
rect 2646 3464 2652 3465
rect 2782 3469 2788 3470
rect 2782 3465 2783 3469
rect 2787 3465 2788 3469
rect 2782 3464 2788 3465
rect 2096 3451 2098 3464
rect 2224 3451 2226 3464
rect 2360 3451 2362 3464
rect 2504 3451 2506 3464
rect 2648 3451 2650 3464
rect 2784 3451 2786 3464
rect 2023 3450 2027 3451
rect 2023 3445 2027 3446
rect 2095 3450 2099 3451
rect 2095 3445 2099 3446
rect 2191 3450 2195 3451
rect 2191 3445 2195 3446
rect 2223 3450 2227 3451
rect 2223 3445 2227 3446
rect 2359 3450 2363 3451
rect 2359 3445 2363 3446
rect 2367 3450 2371 3451
rect 2367 3445 2371 3446
rect 2503 3450 2507 3451
rect 2503 3445 2507 3446
rect 2543 3450 2547 3451
rect 2543 3445 2547 3446
rect 2647 3450 2651 3451
rect 2647 3445 2651 3446
rect 2711 3450 2715 3451
rect 2711 3445 2715 3446
rect 2783 3450 2787 3451
rect 2783 3445 2787 3446
rect 2024 3440 2026 3445
rect 2192 3440 2194 3445
rect 2368 3440 2370 3445
rect 2544 3440 2546 3445
rect 2712 3440 2714 3445
rect 2022 3439 2028 3440
rect 2022 3435 2023 3439
rect 2027 3435 2028 3439
rect 2022 3434 2028 3435
rect 2190 3439 2196 3440
rect 2190 3435 2191 3439
rect 2195 3435 2196 3439
rect 2190 3434 2196 3435
rect 2366 3439 2372 3440
rect 2366 3435 2367 3439
rect 2371 3435 2372 3439
rect 2366 3434 2372 3435
rect 2542 3439 2548 3440
rect 2542 3435 2543 3439
rect 2547 3435 2548 3439
rect 2542 3434 2548 3435
rect 2710 3439 2716 3440
rect 2710 3435 2711 3439
rect 2715 3435 2716 3439
rect 2710 3434 2716 3435
rect 2800 3432 2802 3514
rect 2936 3510 2938 3521
rect 3002 3519 3008 3520
rect 3002 3515 3003 3519
rect 3007 3515 3008 3519
rect 3002 3514 3008 3515
rect 2934 3509 2940 3510
rect 2934 3505 2935 3509
rect 2939 3505 2940 3509
rect 2934 3504 2940 3505
rect 3004 3492 3006 3514
rect 3080 3510 3082 3521
rect 3216 3520 3218 3554
rect 3574 3552 3575 3556
rect 3579 3552 3580 3556
rect 3574 3551 3580 3552
rect 3230 3543 3236 3544
rect 3230 3539 3231 3543
rect 3235 3539 3236 3543
rect 3230 3538 3236 3539
rect 3232 3527 3234 3538
rect 3576 3527 3578 3551
rect 3223 3526 3227 3527
rect 3223 3521 3227 3522
rect 3231 3526 3235 3527
rect 3231 3521 3235 3522
rect 3575 3526 3579 3527
rect 3575 3521 3579 3522
rect 3182 3519 3188 3520
rect 3182 3515 3183 3519
rect 3187 3515 3188 3519
rect 3182 3514 3188 3515
rect 3214 3519 3220 3520
rect 3214 3515 3215 3519
rect 3219 3515 3220 3519
rect 3214 3514 3220 3515
rect 3078 3509 3084 3510
rect 3078 3505 3079 3509
rect 3083 3505 3084 3509
rect 3078 3504 3084 3505
rect 3184 3492 3186 3514
rect 3224 3510 3226 3521
rect 3222 3509 3228 3510
rect 3222 3505 3223 3509
rect 3227 3505 3228 3509
rect 3222 3504 3228 3505
rect 3576 3497 3578 3521
rect 3574 3496 3580 3497
rect 3574 3492 3575 3496
rect 3579 3492 3580 3496
rect 3002 3491 3008 3492
rect 3002 3487 3003 3491
rect 3007 3487 3008 3491
rect 3002 3486 3008 3487
rect 3182 3491 3188 3492
rect 3574 3491 3580 3492
rect 3182 3487 3183 3491
rect 3187 3487 3188 3491
rect 3182 3486 3188 3487
rect 2886 3479 2892 3480
rect 2886 3475 2887 3479
rect 2891 3475 2892 3479
rect 2886 3474 2892 3475
rect 3574 3479 3580 3480
rect 3574 3475 3575 3479
rect 3579 3475 3580 3479
rect 3574 3474 3580 3475
rect 2871 3450 2875 3451
rect 2871 3445 2875 3446
rect 2872 3440 2874 3445
rect 2870 3439 2876 3440
rect 2870 3435 2871 3439
rect 2875 3435 2876 3439
rect 2870 3434 2876 3435
rect 1990 3431 1996 3432
rect 1470 3426 1476 3427
rect 1862 3429 1868 3430
rect 1862 3425 1863 3429
rect 1867 3425 1868 3429
rect 1990 3427 1991 3431
rect 1995 3427 1996 3431
rect 1990 3426 1996 3427
rect 2798 3431 2804 3432
rect 2798 3427 2799 3431
rect 2803 3427 2804 3431
rect 2798 3426 2804 3427
rect 1862 3424 1868 3425
rect 110 3419 116 3420
rect 110 3415 111 3419
rect 115 3415 116 3419
rect 110 3414 116 3415
rect 150 3419 156 3420
rect 150 3415 151 3419
rect 155 3415 156 3419
rect 150 3414 156 3415
rect 1822 3419 1828 3420
rect 1822 3415 1823 3419
rect 1827 3415 1828 3419
rect 1822 3414 1828 3415
rect 2090 3415 2096 3416
rect 112 3399 114 3414
rect 111 3398 115 3399
rect 111 3393 115 3394
rect 135 3398 139 3399
rect 135 3393 139 3394
rect 112 3378 114 3393
rect 136 3388 138 3393
rect 134 3387 140 3388
rect 134 3383 135 3387
rect 139 3383 140 3387
rect 134 3382 140 3383
rect 110 3377 116 3378
rect 110 3373 111 3377
rect 115 3373 116 3377
rect 110 3372 116 3373
rect 110 3360 116 3361
rect 110 3356 111 3360
rect 115 3356 116 3360
rect 110 3355 116 3356
rect 112 3327 114 3355
rect 142 3347 148 3348
rect 142 3343 143 3347
rect 147 3343 148 3347
rect 142 3342 148 3343
rect 144 3327 146 3342
rect 152 3336 154 3414
rect 166 3409 172 3410
rect 166 3405 167 3409
rect 171 3405 172 3409
rect 166 3404 172 3405
rect 294 3409 300 3410
rect 294 3405 295 3409
rect 299 3405 300 3409
rect 294 3404 300 3405
rect 438 3409 444 3410
rect 438 3405 439 3409
rect 443 3405 444 3409
rect 438 3404 444 3405
rect 582 3409 588 3410
rect 582 3405 583 3409
rect 587 3405 588 3409
rect 582 3404 588 3405
rect 734 3409 740 3410
rect 734 3405 735 3409
rect 739 3405 740 3409
rect 734 3404 740 3405
rect 886 3409 892 3410
rect 886 3405 887 3409
rect 891 3405 892 3409
rect 886 3404 892 3405
rect 1030 3409 1036 3410
rect 1030 3405 1031 3409
rect 1035 3405 1036 3409
rect 1030 3404 1036 3405
rect 1174 3409 1180 3410
rect 1174 3405 1175 3409
rect 1179 3405 1180 3409
rect 1174 3404 1180 3405
rect 1318 3409 1324 3410
rect 1318 3405 1319 3409
rect 1323 3405 1324 3409
rect 1318 3404 1324 3405
rect 1470 3409 1476 3410
rect 1470 3405 1471 3409
rect 1475 3405 1476 3409
rect 1470 3404 1476 3405
rect 168 3399 170 3404
rect 296 3399 298 3404
rect 440 3399 442 3404
rect 584 3399 586 3404
rect 736 3399 738 3404
rect 888 3399 890 3404
rect 1032 3399 1034 3404
rect 1176 3399 1178 3404
rect 1222 3403 1228 3404
rect 1222 3399 1223 3403
rect 1227 3399 1228 3403
rect 1320 3399 1322 3404
rect 1472 3399 1474 3404
rect 1824 3399 1826 3414
rect 1862 3412 1868 3413
rect 1862 3408 1863 3412
rect 1867 3408 1868 3412
rect 2090 3411 2091 3415
rect 2095 3411 2096 3415
rect 2090 3410 2096 3411
rect 2258 3415 2264 3416
rect 2258 3411 2259 3415
rect 2263 3411 2264 3415
rect 2258 3410 2264 3411
rect 2434 3415 2440 3416
rect 2434 3411 2435 3415
rect 2439 3411 2440 3415
rect 2434 3410 2440 3411
rect 1862 3407 1868 3408
rect 167 3398 171 3399
rect 167 3393 171 3394
rect 263 3398 267 3399
rect 263 3393 267 3394
rect 295 3398 299 3399
rect 295 3393 299 3394
rect 407 3398 411 3399
rect 407 3393 411 3394
rect 439 3398 443 3399
rect 439 3393 443 3394
rect 567 3398 571 3399
rect 567 3393 571 3394
rect 583 3398 587 3399
rect 583 3393 587 3394
rect 727 3398 731 3399
rect 727 3393 731 3394
rect 735 3398 739 3399
rect 735 3393 739 3394
rect 887 3398 891 3399
rect 887 3393 891 3394
rect 1031 3398 1035 3399
rect 1031 3393 1035 3394
rect 1047 3398 1051 3399
rect 1047 3393 1051 3394
rect 1175 3398 1179 3399
rect 1175 3393 1179 3394
rect 1207 3398 1211 3399
rect 1222 3398 1228 3399
rect 1319 3398 1323 3399
rect 1207 3393 1211 3394
rect 264 3388 266 3393
rect 408 3388 410 3393
rect 568 3388 570 3393
rect 728 3388 730 3393
rect 888 3388 890 3393
rect 1048 3388 1050 3393
rect 1208 3388 1210 3393
rect 262 3387 268 3388
rect 262 3383 263 3387
rect 267 3383 268 3387
rect 262 3382 268 3383
rect 406 3387 412 3388
rect 406 3383 407 3387
rect 411 3383 412 3387
rect 406 3382 412 3383
rect 566 3387 572 3388
rect 566 3383 567 3387
rect 571 3383 572 3387
rect 566 3382 572 3383
rect 726 3387 732 3388
rect 726 3383 727 3387
rect 731 3383 732 3387
rect 726 3382 732 3383
rect 886 3387 892 3388
rect 886 3383 887 3387
rect 891 3383 892 3387
rect 886 3382 892 3383
rect 1046 3387 1052 3388
rect 1046 3383 1047 3387
rect 1051 3383 1052 3387
rect 1046 3382 1052 3383
rect 1206 3387 1212 3388
rect 1206 3383 1207 3387
rect 1211 3383 1212 3387
rect 1206 3382 1212 3383
rect 682 3379 688 3380
rect 682 3375 683 3379
rect 687 3375 688 3379
rect 682 3374 688 3375
rect 270 3347 276 3348
rect 270 3343 271 3347
rect 275 3343 276 3347
rect 270 3342 276 3343
rect 414 3347 420 3348
rect 414 3343 415 3347
rect 419 3343 420 3347
rect 414 3342 420 3343
rect 574 3347 580 3348
rect 574 3343 575 3347
rect 579 3343 580 3347
rect 574 3342 580 3343
rect 215 3340 219 3341
rect 150 3335 156 3336
rect 215 3335 219 3336
rect 150 3331 151 3335
rect 155 3331 156 3335
rect 150 3330 156 3331
rect 111 3326 115 3327
rect 111 3321 115 3322
rect 143 3326 147 3327
rect 143 3321 147 3322
rect 207 3326 211 3327
rect 207 3321 211 3322
rect 112 3297 114 3321
rect 208 3310 210 3321
rect 216 3320 218 3335
rect 272 3327 274 3342
rect 416 3327 418 3342
rect 576 3327 578 3342
rect 684 3341 686 3374
rect 734 3347 740 3348
rect 734 3343 735 3347
rect 739 3343 740 3347
rect 734 3342 740 3343
rect 894 3347 900 3348
rect 894 3343 895 3347
rect 899 3343 900 3347
rect 894 3342 900 3343
rect 1054 3347 1060 3348
rect 1054 3343 1055 3347
rect 1059 3343 1060 3347
rect 1054 3342 1060 3343
rect 1214 3347 1220 3348
rect 1214 3343 1215 3347
rect 1219 3343 1220 3347
rect 1214 3342 1220 3343
rect 683 3340 687 3341
rect 683 3335 687 3336
rect 736 3327 738 3342
rect 896 3327 898 3342
rect 1056 3327 1058 3342
rect 1216 3327 1218 3342
rect 1224 3336 1226 3398
rect 1319 3393 1323 3394
rect 1367 3398 1371 3399
rect 1367 3393 1371 3394
rect 1471 3398 1475 3399
rect 1471 3393 1475 3394
rect 1527 3398 1531 3399
rect 1527 3393 1531 3394
rect 1823 3398 1827 3399
rect 1823 3393 1827 3394
rect 1368 3388 1370 3393
rect 1528 3388 1530 3393
rect 1366 3387 1372 3388
rect 1366 3383 1367 3387
rect 1371 3383 1372 3387
rect 1366 3382 1372 3383
rect 1526 3387 1532 3388
rect 1526 3383 1527 3387
rect 1531 3383 1532 3387
rect 1526 3382 1532 3383
rect 1824 3378 1826 3393
rect 1822 3377 1828 3378
rect 1822 3373 1823 3377
rect 1827 3373 1828 3377
rect 1864 3375 1866 3407
rect 1894 3399 1900 3400
rect 1894 3395 1895 3399
rect 1899 3395 1900 3399
rect 1894 3394 1900 3395
rect 2030 3399 2036 3400
rect 2030 3395 2031 3399
rect 2035 3395 2036 3399
rect 2030 3394 2036 3395
rect 1886 3387 1892 3388
rect 1886 3383 1887 3387
rect 1891 3383 1892 3387
rect 1886 3382 1892 3383
rect 1822 3372 1828 3373
rect 1863 3374 1867 3375
rect 1863 3369 1867 3370
rect 1822 3360 1828 3361
rect 1822 3356 1823 3360
rect 1827 3356 1828 3360
rect 1822 3355 1828 3356
rect 1374 3347 1380 3348
rect 1374 3343 1375 3347
rect 1379 3343 1380 3347
rect 1374 3342 1380 3343
rect 1534 3347 1540 3348
rect 1534 3343 1535 3347
rect 1539 3343 1540 3347
rect 1534 3342 1540 3343
rect 1222 3335 1228 3336
rect 1222 3331 1223 3335
rect 1227 3331 1228 3335
rect 1222 3330 1228 3331
rect 1376 3327 1378 3342
rect 1536 3327 1538 3342
rect 1824 3327 1826 3355
rect 1864 3345 1866 3369
rect 1862 3344 1868 3345
rect 1862 3340 1863 3344
rect 1867 3340 1868 3344
rect 1888 3340 1890 3382
rect 1896 3375 1898 3394
rect 2032 3375 2034 3394
rect 1895 3374 1899 3375
rect 1895 3369 1899 3370
rect 2031 3374 2035 3375
rect 2031 3369 2035 3370
rect 1896 3358 1898 3369
rect 2032 3358 2034 3369
rect 2092 3368 2094 3410
rect 2198 3399 2204 3400
rect 2198 3395 2199 3399
rect 2203 3395 2204 3399
rect 2198 3394 2204 3395
rect 2200 3375 2202 3394
rect 2260 3388 2262 3410
rect 2374 3399 2380 3400
rect 2374 3395 2375 3399
rect 2379 3395 2380 3399
rect 2374 3394 2380 3395
rect 2258 3387 2264 3388
rect 2258 3383 2259 3387
rect 2263 3383 2264 3387
rect 2258 3382 2264 3383
rect 2376 3375 2378 3394
rect 2436 3388 2438 3410
rect 2550 3399 2556 3400
rect 2550 3395 2551 3399
rect 2555 3395 2556 3399
rect 2550 3394 2556 3395
rect 2718 3399 2724 3400
rect 2718 3395 2719 3399
rect 2723 3395 2724 3399
rect 2718 3394 2724 3395
rect 2878 3399 2884 3400
rect 2878 3395 2879 3399
rect 2883 3395 2884 3399
rect 2878 3394 2884 3395
rect 2434 3387 2440 3388
rect 2434 3383 2435 3387
rect 2439 3383 2440 3387
rect 2434 3382 2440 3383
rect 2552 3375 2554 3394
rect 2710 3387 2716 3388
rect 2710 3383 2711 3387
rect 2715 3383 2716 3387
rect 2710 3382 2716 3383
rect 2199 3374 2203 3375
rect 2199 3369 2203 3370
rect 2375 3374 2379 3375
rect 2375 3369 2379 3370
rect 2551 3374 2555 3375
rect 2551 3369 2555 3370
rect 2090 3367 2096 3368
rect 2090 3363 2091 3367
rect 2095 3363 2096 3367
rect 2090 3362 2096 3363
rect 2200 3358 2202 3369
rect 2376 3358 2378 3369
rect 2552 3358 2554 3369
rect 1894 3357 1900 3358
rect 1894 3353 1895 3357
rect 1899 3353 1900 3357
rect 1894 3352 1900 3353
rect 2030 3357 2036 3358
rect 2030 3353 2031 3357
rect 2035 3353 2036 3357
rect 2030 3352 2036 3353
rect 2198 3357 2204 3358
rect 2198 3353 2199 3357
rect 2203 3353 2204 3357
rect 2198 3352 2204 3353
rect 2374 3357 2380 3358
rect 2374 3353 2375 3357
rect 2379 3353 2380 3357
rect 2374 3352 2380 3353
rect 2550 3357 2556 3358
rect 2550 3353 2551 3357
rect 2555 3353 2556 3357
rect 2550 3352 2556 3353
rect 2712 3340 2714 3382
rect 2720 3375 2722 3394
rect 2880 3375 2882 3394
rect 2888 3388 2890 3474
rect 2926 3469 2932 3470
rect 2926 3465 2927 3469
rect 2931 3465 2932 3469
rect 2926 3464 2932 3465
rect 3070 3469 3076 3470
rect 3070 3465 3071 3469
rect 3075 3465 3076 3469
rect 3070 3464 3076 3465
rect 3214 3469 3220 3470
rect 3214 3465 3215 3469
rect 3219 3465 3220 3469
rect 3214 3464 3220 3465
rect 2928 3451 2930 3464
rect 3072 3451 3074 3464
rect 3216 3451 3218 3464
rect 3576 3451 3578 3474
rect 2927 3450 2931 3451
rect 2927 3445 2931 3446
rect 3031 3450 3035 3451
rect 3031 3445 3035 3446
rect 3071 3450 3075 3451
rect 3071 3445 3075 3446
rect 3191 3450 3195 3451
rect 3191 3445 3195 3446
rect 3215 3450 3219 3451
rect 3215 3445 3219 3446
rect 3359 3450 3363 3451
rect 3359 3445 3363 3446
rect 3575 3450 3579 3451
rect 3575 3445 3579 3446
rect 3032 3440 3034 3445
rect 3192 3440 3194 3445
rect 3360 3440 3362 3445
rect 3030 3439 3036 3440
rect 3030 3435 3031 3439
rect 3035 3435 3036 3439
rect 3030 3434 3036 3435
rect 3190 3439 3196 3440
rect 3190 3435 3191 3439
rect 3195 3435 3196 3439
rect 3190 3434 3196 3435
rect 3358 3439 3364 3440
rect 3358 3435 3359 3439
rect 3363 3435 3364 3439
rect 3358 3434 3364 3435
rect 3258 3431 3264 3432
rect 3258 3427 3259 3431
rect 3263 3427 3264 3431
rect 3576 3430 3578 3445
rect 3258 3426 3264 3427
rect 3574 3429 3580 3430
rect 3038 3399 3044 3400
rect 3038 3395 3039 3399
rect 3043 3395 3044 3399
rect 3198 3399 3204 3400
rect 3038 3394 3044 3395
rect 3047 3396 3051 3397
rect 2886 3387 2892 3388
rect 2886 3383 2887 3387
rect 2891 3383 2892 3387
rect 2886 3382 2892 3383
rect 3040 3375 3042 3394
rect 3198 3395 3199 3399
rect 3203 3395 3204 3399
rect 3260 3397 3262 3426
rect 3574 3425 3575 3429
rect 3579 3425 3580 3429
rect 3574 3424 3580 3425
rect 3574 3412 3580 3413
rect 3574 3408 3575 3412
rect 3579 3408 3580 3412
rect 3574 3407 3580 3408
rect 3366 3399 3372 3400
rect 3198 3394 3204 3395
rect 3259 3396 3263 3397
rect 3047 3391 3051 3392
rect 2719 3374 2723 3375
rect 2719 3369 2723 3370
rect 2879 3374 2883 3375
rect 2879 3369 2883 3370
rect 3039 3374 3043 3375
rect 3039 3369 3043 3370
rect 2720 3358 2722 3369
rect 2880 3358 2882 3369
rect 2886 3367 2892 3368
rect 2886 3363 2887 3367
rect 2891 3363 2892 3367
rect 2886 3362 2892 3363
rect 2718 3357 2724 3358
rect 2718 3353 2719 3357
rect 2723 3353 2724 3357
rect 2718 3352 2724 3353
rect 2878 3357 2884 3358
rect 2878 3353 2879 3357
rect 2883 3353 2884 3357
rect 2878 3352 2884 3353
rect 1862 3339 1868 3340
rect 1886 3339 1892 3340
rect 1886 3335 1887 3339
rect 1891 3335 1892 3339
rect 1886 3334 1892 3335
rect 2710 3339 2716 3340
rect 2710 3335 2711 3339
rect 2715 3335 2716 3339
rect 2710 3334 2716 3335
rect 1862 3327 1868 3328
rect 271 3326 275 3327
rect 271 3321 275 3322
rect 335 3326 339 3327
rect 335 3321 339 3322
rect 415 3326 419 3327
rect 415 3321 419 3322
rect 479 3326 483 3327
rect 479 3321 483 3322
rect 575 3326 579 3327
rect 575 3321 579 3322
rect 639 3326 643 3327
rect 639 3321 643 3322
rect 735 3326 739 3327
rect 735 3321 739 3322
rect 807 3326 811 3327
rect 807 3321 811 3322
rect 895 3326 899 3327
rect 895 3321 899 3322
rect 983 3326 987 3327
rect 983 3321 987 3322
rect 1055 3326 1059 3327
rect 1055 3321 1059 3322
rect 1167 3326 1171 3327
rect 1167 3321 1171 3322
rect 1215 3326 1219 3327
rect 1215 3321 1219 3322
rect 1351 3326 1355 3327
rect 1351 3321 1355 3322
rect 1375 3326 1379 3327
rect 1375 3321 1379 3322
rect 1535 3326 1539 3327
rect 1535 3321 1539 3322
rect 1543 3326 1547 3327
rect 1543 3321 1547 3322
rect 1823 3326 1827 3327
rect 1862 3323 1863 3327
rect 1867 3323 1868 3327
rect 1862 3322 1868 3323
rect 2478 3327 2484 3328
rect 2478 3323 2479 3327
rect 2483 3323 2484 3327
rect 2478 3322 2484 3323
rect 1823 3321 1827 3322
rect 214 3319 220 3320
rect 214 3315 215 3319
rect 219 3315 220 3319
rect 214 3314 220 3315
rect 336 3310 338 3321
rect 480 3310 482 3321
rect 640 3310 642 3321
rect 808 3310 810 3321
rect 984 3310 986 3321
rect 1078 3319 1084 3320
rect 1078 3315 1079 3319
rect 1083 3315 1084 3319
rect 1078 3314 1084 3315
rect 206 3309 212 3310
rect 206 3305 207 3309
rect 211 3305 212 3309
rect 206 3304 212 3305
rect 334 3309 340 3310
rect 334 3305 335 3309
rect 339 3305 340 3309
rect 334 3304 340 3305
rect 478 3309 484 3310
rect 478 3305 479 3309
rect 483 3305 484 3309
rect 478 3304 484 3305
rect 638 3309 644 3310
rect 638 3305 639 3309
rect 643 3305 644 3309
rect 638 3304 644 3305
rect 806 3309 812 3310
rect 806 3305 807 3309
rect 811 3305 812 3309
rect 806 3304 812 3305
rect 982 3309 988 3310
rect 982 3305 983 3309
rect 987 3305 988 3309
rect 982 3304 988 3305
rect 110 3296 116 3297
rect 110 3292 111 3296
rect 115 3292 116 3296
rect 1080 3292 1082 3314
rect 1168 3310 1170 3321
rect 1174 3319 1180 3320
rect 1174 3315 1175 3319
rect 1179 3315 1180 3319
rect 1174 3314 1180 3315
rect 1166 3309 1172 3310
rect 1166 3305 1167 3309
rect 1171 3305 1172 3309
rect 1166 3304 1172 3305
rect 110 3291 116 3292
rect 1078 3291 1084 3292
rect 1078 3287 1079 3291
rect 1083 3287 1084 3291
rect 1078 3286 1084 3287
rect 110 3279 116 3280
rect 110 3275 111 3279
rect 115 3275 116 3279
rect 110 3274 116 3275
rect 112 3255 114 3274
rect 198 3269 204 3270
rect 198 3265 199 3269
rect 203 3265 204 3269
rect 198 3264 204 3265
rect 326 3269 332 3270
rect 326 3265 327 3269
rect 331 3265 332 3269
rect 326 3264 332 3265
rect 470 3269 476 3270
rect 470 3265 471 3269
rect 475 3265 476 3269
rect 470 3264 476 3265
rect 630 3269 636 3270
rect 630 3265 631 3269
rect 635 3265 636 3269
rect 630 3264 636 3265
rect 798 3269 804 3270
rect 798 3265 799 3269
rect 803 3265 804 3269
rect 798 3264 804 3265
rect 974 3269 980 3270
rect 974 3265 975 3269
rect 979 3265 980 3269
rect 974 3264 980 3265
rect 1158 3269 1164 3270
rect 1158 3265 1159 3269
rect 1163 3265 1164 3269
rect 1158 3264 1164 3265
rect 200 3255 202 3264
rect 328 3255 330 3264
rect 472 3255 474 3264
rect 632 3255 634 3264
rect 800 3255 802 3264
rect 976 3255 978 3264
rect 1160 3255 1162 3264
rect 111 3254 115 3255
rect 111 3249 115 3250
rect 199 3254 203 3255
rect 199 3249 203 3250
rect 327 3254 331 3255
rect 327 3249 331 3250
rect 367 3254 371 3255
rect 367 3249 371 3250
rect 471 3254 475 3255
rect 471 3249 475 3250
rect 503 3254 507 3255
rect 503 3249 507 3250
rect 631 3254 635 3255
rect 631 3249 635 3250
rect 639 3254 643 3255
rect 639 3249 643 3250
rect 783 3254 787 3255
rect 783 3249 787 3250
rect 799 3254 803 3255
rect 799 3249 803 3250
rect 935 3254 939 3255
rect 935 3249 939 3250
rect 975 3254 979 3255
rect 975 3249 979 3250
rect 1095 3254 1099 3255
rect 1095 3249 1099 3250
rect 1159 3254 1163 3255
rect 1159 3249 1163 3250
rect 112 3234 114 3249
rect 368 3244 370 3249
rect 504 3244 506 3249
rect 640 3244 642 3249
rect 784 3244 786 3249
rect 936 3244 938 3249
rect 1096 3244 1098 3249
rect 366 3243 372 3244
rect 366 3239 367 3243
rect 371 3239 372 3243
rect 366 3238 372 3239
rect 502 3243 508 3244
rect 502 3239 503 3243
rect 507 3239 508 3243
rect 502 3238 508 3239
rect 638 3243 644 3244
rect 638 3239 639 3243
rect 643 3239 644 3243
rect 638 3238 644 3239
rect 782 3243 788 3244
rect 782 3239 783 3243
rect 787 3239 788 3243
rect 782 3238 788 3239
rect 934 3243 940 3244
rect 934 3239 935 3243
rect 939 3239 940 3243
rect 934 3238 940 3239
rect 1094 3243 1100 3244
rect 1094 3239 1095 3243
rect 1099 3239 1100 3243
rect 1094 3238 1100 3239
rect 1176 3236 1178 3314
rect 1352 3310 1354 3321
rect 1426 3319 1432 3320
rect 1426 3315 1427 3319
rect 1431 3315 1432 3319
rect 1426 3314 1432 3315
rect 1350 3309 1356 3310
rect 1350 3305 1351 3309
rect 1355 3305 1356 3309
rect 1350 3304 1356 3305
rect 1428 3292 1430 3314
rect 1544 3310 1546 3321
rect 1542 3309 1548 3310
rect 1542 3305 1543 3309
rect 1547 3305 1548 3309
rect 1542 3304 1548 3305
rect 1824 3297 1826 3321
rect 1864 3307 1866 3322
rect 1886 3317 1892 3318
rect 1886 3313 1887 3317
rect 1891 3313 1892 3317
rect 1886 3312 1892 3313
rect 2022 3317 2028 3318
rect 2022 3313 2023 3317
rect 2027 3313 2028 3317
rect 2022 3312 2028 3313
rect 2190 3317 2196 3318
rect 2190 3313 2191 3317
rect 2195 3313 2196 3317
rect 2190 3312 2196 3313
rect 2366 3317 2372 3318
rect 2366 3313 2367 3317
rect 2371 3313 2372 3317
rect 2366 3312 2372 3313
rect 1888 3307 1890 3312
rect 2024 3307 2026 3312
rect 2192 3307 2194 3312
rect 2368 3307 2370 3312
rect 1863 3306 1867 3307
rect 1863 3301 1867 3302
rect 1887 3306 1891 3307
rect 1887 3301 1891 3302
rect 2007 3306 2011 3307
rect 2007 3301 2011 3302
rect 2023 3306 2027 3307
rect 2023 3301 2027 3302
rect 2151 3306 2155 3307
rect 2151 3301 2155 3302
rect 2191 3306 2195 3307
rect 2191 3301 2195 3302
rect 2303 3306 2307 3307
rect 2303 3301 2307 3302
rect 2367 3306 2371 3307
rect 2367 3301 2371 3302
rect 2463 3306 2467 3307
rect 2463 3301 2467 3302
rect 1822 3296 1828 3297
rect 1822 3292 1823 3296
rect 1827 3292 1828 3296
rect 1426 3291 1432 3292
rect 1822 3291 1828 3292
rect 1426 3287 1427 3291
rect 1431 3287 1432 3291
rect 1426 3286 1432 3287
rect 1864 3286 1866 3301
rect 1888 3296 1890 3301
rect 2008 3296 2010 3301
rect 2152 3296 2154 3301
rect 2304 3296 2306 3301
rect 2464 3296 2466 3301
rect 1886 3295 1892 3296
rect 1886 3291 1887 3295
rect 1891 3291 1892 3295
rect 1886 3290 1892 3291
rect 2006 3295 2012 3296
rect 2006 3291 2007 3295
rect 2011 3291 2012 3295
rect 2006 3290 2012 3291
rect 2150 3295 2156 3296
rect 2150 3291 2151 3295
rect 2155 3291 2156 3295
rect 2150 3290 2156 3291
rect 2302 3295 2308 3296
rect 2302 3291 2303 3295
rect 2307 3291 2308 3295
rect 2302 3290 2308 3291
rect 2462 3295 2468 3296
rect 2462 3291 2463 3295
rect 2467 3291 2468 3295
rect 2462 3290 2468 3291
rect 1862 3285 1868 3286
rect 1862 3281 1863 3285
rect 1867 3281 1868 3285
rect 1862 3280 1868 3281
rect 1822 3279 1828 3280
rect 1822 3275 1823 3279
rect 1827 3275 1828 3279
rect 1822 3274 1828 3275
rect 2183 3276 2187 3277
rect 1342 3269 1348 3270
rect 1342 3265 1343 3269
rect 1347 3265 1348 3269
rect 1342 3264 1348 3265
rect 1534 3269 1540 3270
rect 1534 3265 1535 3269
rect 1539 3265 1540 3269
rect 1534 3264 1540 3265
rect 1344 3255 1346 3264
rect 1536 3255 1538 3264
rect 1824 3255 1826 3274
rect 1954 3271 1960 3272
rect 2183 3271 2187 3272
rect 2234 3271 2240 3272
rect 1862 3268 1868 3269
rect 1862 3264 1863 3268
rect 1867 3264 1868 3268
rect 1954 3267 1955 3271
rect 1959 3267 1960 3271
rect 1954 3266 1960 3267
rect 1862 3263 1868 3264
rect 1255 3254 1259 3255
rect 1255 3249 1259 3250
rect 1343 3254 1347 3255
rect 1343 3249 1347 3250
rect 1415 3254 1419 3255
rect 1415 3249 1419 3250
rect 1535 3254 1539 3255
rect 1535 3249 1539 3250
rect 1575 3254 1579 3255
rect 1575 3249 1579 3250
rect 1823 3254 1827 3255
rect 1823 3249 1827 3250
rect 1256 3244 1258 3249
rect 1416 3244 1418 3249
rect 1576 3244 1578 3249
rect 1254 3243 1260 3244
rect 1254 3239 1255 3243
rect 1259 3239 1260 3243
rect 1254 3238 1260 3239
rect 1414 3243 1420 3244
rect 1414 3239 1415 3243
rect 1419 3239 1420 3243
rect 1414 3238 1420 3239
rect 1574 3243 1580 3244
rect 1574 3239 1575 3243
rect 1579 3239 1580 3243
rect 1574 3238 1580 3239
rect 710 3235 716 3236
rect 110 3233 116 3234
rect 110 3229 111 3233
rect 115 3229 116 3233
rect 710 3231 711 3235
rect 715 3231 716 3235
rect 710 3230 716 3231
rect 1174 3235 1180 3236
rect 1174 3231 1175 3235
rect 1179 3231 1180 3235
rect 1824 3234 1826 3249
rect 1174 3230 1180 3231
rect 1822 3233 1828 3234
rect 110 3228 116 3229
rect 110 3216 116 3217
rect 110 3212 111 3216
rect 115 3212 116 3216
rect 110 3211 116 3212
rect 112 3179 114 3211
rect 374 3203 380 3204
rect 374 3199 375 3203
rect 379 3199 380 3203
rect 374 3198 380 3199
rect 510 3203 516 3204
rect 510 3199 511 3203
rect 515 3199 516 3203
rect 510 3198 516 3199
rect 646 3203 652 3204
rect 646 3199 647 3203
rect 651 3199 652 3203
rect 646 3198 652 3199
rect 376 3179 378 3198
rect 487 3196 491 3197
rect 487 3191 491 3192
rect 111 3178 115 3179
rect 111 3173 115 3174
rect 375 3178 379 3179
rect 375 3173 379 3174
rect 447 3178 451 3179
rect 447 3173 451 3174
rect 112 3149 114 3173
rect 448 3162 450 3173
rect 488 3172 490 3191
rect 512 3179 514 3198
rect 648 3179 650 3198
rect 712 3197 714 3230
rect 1822 3229 1823 3233
rect 1827 3229 1828 3233
rect 1864 3231 1866 3263
rect 1894 3255 1900 3256
rect 1894 3251 1895 3255
rect 1899 3251 1900 3255
rect 1956 3251 1958 3266
rect 1894 3250 1900 3251
rect 1896 3231 1898 3250
rect 1952 3249 1958 3251
rect 2014 3255 2020 3256
rect 2014 3251 2015 3255
rect 2019 3251 2020 3255
rect 2014 3250 2020 3251
rect 2158 3255 2164 3256
rect 2158 3251 2159 3255
rect 2163 3251 2164 3255
rect 2158 3250 2164 3251
rect 2167 3252 2171 3253
rect 1952 3244 1954 3249
rect 1950 3243 1956 3244
rect 1950 3239 1951 3243
rect 1955 3239 1956 3243
rect 1950 3238 1956 3239
rect 1958 3243 1964 3244
rect 1958 3239 1959 3243
rect 1963 3239 1964 3243
rect 1958 3238 1964 3239
rect 1822 3228 1828 3229
rect 1863 3230 1867 3231
rect 1863 3225 1867 3226
rect 1895 3230 1899 3231
rect 1895 3225 1899 3226
rect 1162 3219 1168 3220
rect 1162 3215 1163 3219
rect 1167 3215 1168 3219
rect 1162 3214 1168 3215
rect 1646 3219 1652 3220
rect 1646 3215 1647 3219
rect 1651 3215 1652 3219
rect 1646 3214 1652 3215
rect 1822 3216 1828 3217
rect 1164 3205 1166 3214
rect 951 3204 955 3205
rect 1163 3204 1167 3205
rect 790 3203 796 3204
rect 790 3199 791 3203
rect 795 3199 796 3203
rect 790 3198 796 3199
rect 942 3203 948 3204
rect 942 3199 943 3203
rect 947 3199 948 3203
rect 951 3199 955 3200
rect 1102 3203 1108 3204
rect 1102 3199 1103 3203
rect 1107 3199 1108 3203
rect 1163 3199 1167 3200
rect 1262 3203 1268 3204
rect 1262 3199 1263 3203
rect 1267 3199 1268 3203
rect 942 3198 948 3199
rect 711 3196 715 3197
rect 711 3191 715 3192
rect 792 3179 794 3198
rect 944 3179 946 3198
rect 952 3192 954 3199
rect 1102 3198 1108 3199
rect 1262 3198 1268 3199
rect 1422 3203 1428 3204
rect 1422 3199 1423 3203
rect 1427 3199 1428 3203
rect 1422 3198 1428 3199
rect 1582 3203 1588 3204
rect 1582 3199 1583 3203
rect 1587 3199 1588 3203
rect 1582 3198 1588 3199
rect 950 3191 956 3192
rect 950 3187 951 3191
rect 955 3187 956 3191
rect 950 3186 956 3187
rect 1104 3179 1106 3198
rect 1264 3179 1266 3198
rect 1424 3179 1426 3198
rect 1584 3179 1586 3198
rect 511 3178 515 3179
rect 511 3173 515 3174
rect 559 3178 563 3179
rect 559 3173 563 3174
rect 647 3178 651 3179
rect 647 3173 651 3174
rect 687 3178 691 3179
rect 687 3173 691 3174
rect 791 3178 795 3179
rect 791 3173 795 3174
rect 823 3178 827 3179
rect 823 3173 827 3174
rect 943 3178 947 3179
rect 943 3173 947 3174
rect 975 3178 979 3179
rect 975 3173 979 3174
rect 1103 3178 1107 3179
rect 1103 3173 1107 3174
rect 1135 3178 1139 3179
rect 1135 3173 1139 3174
rect 1263 3178 1267 3179
rect 1263 3173 1267 3174
rect 1295 3178 1299 3179
rect 1295 3173 1299 3174
rect 1423 3178 1427 3179
rect 1423 3173 1427 3174
rect 1463 3178 1467 3179
rect 1463 3173 1467 3174
rect 1583 3178 1587 3179
rect 1583 3173 1587 3174
rect 1639 3178 1643 3179
rect 1639 3173 1643 3174
rect 486 3171 492 3172
rect 486 3167 487 3171
rect 491 3167 492 3171
rect 486 3166 492 3167
rect 560 3162 562 3173
rect 688 3162 690 3173
rect 824 3162 826 3173
rect 976 3162 978 3173
rect 1136 3162 1138 3173
rect 1296 3162 1298 3173
rect 1366 3171 1372 3172
rect 1366 3167 1367 3171
rect 1371 3167 1372 3171
rect 1366 3166 1372 3167
rect 446 3161 452 3162
rect 446 3157 447 3161
rect 451 3157 452 3161
rect 446 3156 452 3157
rect 558 3161 564 3162
rect 558 3157 559 3161
rect 563 3157 564 3161
rect 558 3156 564 3157
rect 686 3161 692 3162
rect 686 3157 687 3161
rect 691 3157 692 3161
rect 686 3156 692 3157
rect 822 3161 828 3162
rect 822 3157 823 3161
rect 827 3157 828 3161
rect 822 3156 828 3157
rect 974 3161 980 3162
rect 974 3157 975 3161
rect 979 3157 980 3161
rect 974 3156 980 3157
rect 1134 3161 1140 3162
rect 1134 3157 1135 3161
rect 1139 3157 1140 3161
rect 1134 3156 1140 3157
rect 1294 3161 1300 3162
rect 1294 3157 1295 3161
rect 1299 3157 1300 3161
rect 1294 3156 1300 3157
rect 110 3148 116 3149
rect 110 3144 111 3148
rect 115 3144 116 3148
rect 110 3143 116 3144
rect 110 3131 116 3132
rect 110 3127 111 3131
rect 115 3127 116 3131
rect 110 3126 116 3127
rect 890 3131 896 3132
rect 890 3127 891 3131
rect 895 3127 896 3131
rect 890 3126 896 3127
rect 112 3103 114 3126
rect 438 3121 444 3122
rect 438 3117 439 3121
rect 443 3117 444 3121
rect 438 3116 444 3117
rect 550 3121 556 3122
rect 550 3117 551 3121
rect 555 3117 556 3121
rect 550 3116 556 3117
rect 678 3121 684 3122
rect 678 3117 679 3121
rect 683 3117 684 3121
rect 678 3116 684 3117
rect 814 3121 820 3122
rect 814 3117 815 3121
rect 819 3117 820 3121
rect 814 3116 820 3117
rect 440 3103 442 3116
rect 552 3103 554 3116
rect 680 3103 682 3116
rect 816 3103 818 3116
rect 111 3102 115 3103
rect 111 3097 115 3098
rect 439 3102 443 3103
rect 439 3097 443 3098
rect 551 3102 555 3103
rect 551 3097 555 3098
rect 663 3102 667 3103
rect 663 3097 667 3098
rect 679 3102 683 3103
rect 679 3097 683 3098
rect 783 3102 787 3103
rect 783 3097 787 3098
rect 815 3102 819 3103
rect 815 3097 819 3098
rect 112 3082 114 3097
rect 552 3092 554 3097
rect 664 3092 666 3097
rect 784 3092 786 3097
rect 550 3091 556 3092
rect 550 3087 551 3091
rect 555 3087 556 3091
rect 550 3086 556 3087
rect 662 3091 668 3092
rect 662 3087 663 3091
rect 667 3087 668 3091
rect 662 3086 668 3087
rect 782 3091 788 3092
rect 782 3087 783 3091
rect 787 3087 788 3091
rect 782 3086 788 3087
rect 110 3081 116 3082
rect 110 3077 111 3081
rect 115 3077 116 3081
rect 892 3077 894 3126
rect 966 3121 972 3122
rect 966 3117 967 3121
rect 971 3117 972 3121
rect 966 3116 972 3117
rect 1126 3121 1132 3122
rect 1126 3117 1127 3121
rect 1131 3117 1132 3121
rect 1126 3116 1132 3117
rect 1286 3121 1292 3122
rect 1286 3117 1287 3121
rect 1291 3117 1292 3121
rect 1286 3116 1292 3117
rect 968 3103 970 3116
rect 1128 3103 1130 3116
rect 1288 3103 1290 3116
rect 903 3102 907 3103
rect 903 3097 907 3098
rect 967 3102 971 3103
rect 967 3097 971 3098
rect 1031 3102 1035 3103
rect 1031 3097 1035 3098
rect 1127 3102 1131 3103
rect 1127 3097 1131 3098
rect 1159 3102 1163 3103
rect 1159 3097 1163 3098
rect 1287 3102 1291 3103
rect 1287 3097 1291 3098
rect 904 3092 906 3097
rect 1032 3092 1034 3097
rect 1160 3092 1162 3097
rect 1288 3092 1290 3097
rect 902 3091 908 3092
rect 902 3087 903 3091
rect 907 3087 908 3091
rect 902 3086 908 3087
rect 1030 3091 1036 3092
rect 1030 3087 1031 3091
rect 1035 3087 1036 3091
rect 1030 3086 1036 3087
rect 1158 3091 1164 3092
rect 1158 3087 1159 3091
rect 1163 3087 1164 3091
rect 1158 3086 1164 3087
rect 1286 3091 1292 3092
rect 1286 3087 1287 3091
rect 1291 3087 1292 3091
rect 1286 3086 1292 3087
rect 1368 3084 1370 3166
rect 1464 3162 1466 3173
rect 1538 3171 1544 3172
rect 1538 3167 1539 3171
rect 1543 3167 1544 3171
rect 1538 3166 1544 3167
rect 1462 3161 1468 3162
rect 1462 3157 1463 3161
rect 1467 3157 1468 3161
rect 1462 3156 1468 3157
rect 1540 3144 1542 3166
rect 1640 3162 1642 3173
rect 1648 3172 1650 3214
rect 1822 3212 1823 3216
rect 1827 3212 1828 3216
rect 1822 3211 1828 3212
rect 1824 3179 1826 3211
rect 1864 3201 1866 3225
rect 1896 3214 1898 3225
rect 1894 3213 1900 3214
rect 1894 3209 1895 3213
rect 1899 3209 1900 3213
rect 1894 3208 1900 3209
rect 1862 3200 1868 3201
rect 1960 3200 1962 3238
rect 2016 3231 2018 3250
rect 2160 3231 2162 3250
rect 2167 3247 2171 3248
rect 2168 3244 2170 3247
rect 2166 3243 2172 3244
rect 2166 3239 2167 3243
rect 2171 3239 2172 3243
rect 2166 3238 2172 3239
rect 2015 3230 2019 3231
rect 2015 3225 2019 3226
rect 2023 3230 2027 3231
rect 2023 3225 2027 3226
rect 2159 3230 2163 3231
rect 2159 3225 2163 3226
rect 2175 3230 2179 3231
rect 2175 3225 2179 3226
rect 1966 3223 1972 3224
rect 1966 3219 1967 3223
rect 1971 3219 1972 3223
rect 1966 3218 1972 3219
rect 1862 3196 1863 3200
rect 1867 3196 1868 3200
rect 1862 3195 1868 3196
rect 1958 3199 1964 3200
rect 1958 3195 1959 3199
rect 1963 3195 1964 3199
rect 1968 3196 1970 3218
rect 2024 3214 2026 3225
rect 2030 3223 2036 3224
rect 2030 3219 2031 3223
rect 2035 3219 2036 3223
rect 2030 3218 2036 3219
rect 2022 3213 2028 3214
rect 2022 3209 2023 3213
rect 2027 3209 2028 3213
rect 2022 3208 2028 3209
rect 1958 3194 1964 3195
rect 1966 3195 1972 3196
rect 1966 3191 1967 3195
rect 1971 3191 1972 3195
rect 1966 3190 1972 3191
rect 1862 3183 1868 3184
rect 1862 3179 1863 3183
rect 1867 3179 1868 3183
rect 1823 3178 1827 3179
rect 1862 3178 1868 3179
rect 1823 3173 1827 3174
rect 1646 3171 1652 3172
rect 1646 3167 1647 3171
rect 1651 3167 1652 3171
rect 1646 3166 1652 3167
rect 1638 3161 1644 3162
rect 1638 3157 1639 3161
rect 1643 3157 1644 3161
rect 1638 3156 1644 3157
rect 1824 3149 1826 3173
rect 1864 3159 1866 3178
rect 1886 3173 1892 3174
rect 1886 3169 1887 3173
rect 1891 3169 1892 3173
rect 1886 3168 1892 3169
rect 2014 3173 2020 3174
rect 2014 3169 2015 3173
rect 2019 3169 2020 3173
rect 2014 3168 2020 3169
rect 1888 3159 1890 3168
rect 2016 3159 2018 3168
rect 1863 3158 1867 3159
rect 1863 3153 1867 3154
rect 1887 3158 1891 3159
rect 1887 3153 1891 3154
rect 2015 3158 2019 3159
rect 2015 3153 2019 3154
rect 1822 3148 1828 3149
rect 1822 3144 1823 3148
rect 1827 3144 1828 3148
rect 1538 3143 1544 3144
rect 1822 3143 1828 3144
rect 1538 3139 1539 3143
rect 1543 3139 1544 3143
rect 1538 3138 1544 3139
rect 1864 3138 1866 3153
rect 1888 3148 1890 3153
rect 1886 3147 1892 3148
rect 1886 3143 1887 3147
rect 1891 3143 1892 3147
rect 1886 3142 1892 3143
rect 2032 3140 2034 3218
rect 2176 3214 2178 3225
rect 2184 3224 2186 3271
rect 2234 3267 2235 3271
rect 2239 3267 2240 3271
rect 2234 3266 2240 3267
rect 2236 3244 2238 3266
rect 2310 3255 2316 3256
rect 2310 3251 2311 3255
rect 2315 3251 2316 3255
rect 2310 3250 2316 3251
rect 2470 3255 2476 3256
rect 2470 3251 2471 3255
rect 2475 3251 2476 3255
rect 2480 3253 2482 3322
rect 2542 3317 2548 3318
rect 2542 3313 2543 3317
rect 2547 3313 2548 3317
rect 2542 3312 2548 3313
rect 2710 3317 2716 3318
rect 2710 3313 2711 3317
rect 2715 3313 2716 3317
rect 2710 3312 2716 3313
rect 2870 3317 2876 3318
rect 2870 3313 2871 3317
rect 2875 3313 2876 3317
rect 2870 3312 2876 3313
rect 2544 3307 2546 3312
rect 2712 3307 2714 3312
rect 2872 3307 2874 3312
rect 2543 3306 2547 3307
rect 2543 3301 2547 3302
rect 2631 3306 2635 3307
rect 2631 3301 2635 3302
rect 2711 3306 2715 3307
rect 2711 3301 2715 3302
rect 2799 3306 2803 3307
rect 2799 3301 2803 3302
rect 2871 3306 2875 3307
rect 2871 3301 2875 3302
rect 2632 3296 2634 3301
rect 2800 3296 2802 3301
rect 2630 3295 2636 3296
rect 2630 3291 2631 3295
rect 2635 3291 2636 3295
rect 2630 3290 2636 3291
rect 2798 3295 2804 3296
rect 2798 3291 2799 3295
rect 2803 3291 2804 3295
rect 2798 3290 2804 3291
rect 2888 3288 2890 3362
rect 3040 3358 3042 3369
rect 3048 3368 3050 3391
rect 3200 3375 3202 3394
rect 3366 3395 3367 3399
rect 3371 3395 3372 3399
rect 3366 3394 3372 3395
rect 3259 3391 3263 3392
rect 3368 3375 3370 3394
rect 3576 3375 3578 3407
rect 3191 3374 3195 3375
rect 3191 3369 3195 3370
rect 3199 3374 3203 3375
rect 3199 3369 3203 3370
rect 3343 3374 3347 3375
rect 3343 3369 3347 3370
rect 3367 3374 3371 3375
rect 3367 3369 3371 3370
rect 3487 3374 3491 3375
rect 3487 3369 3491 3370
rect 3575 3374 3579 3375
rect 3575 3369 3579 3370
rect 3046 3367 3052 3368
rect 3046 3363 3047 3367
rect 3051 3363 3052 3367
rect 3046 3362 3052 3363
rect 3192 3358 3194 3369
rect 3344 3358 3346 3369
rect 3488 3358 3490 3369
rect 3038 3357 3044 3358
rect 3038 3353 3039 3357
rect 3043 3353 3044 3357
rect 3038 3352 3044 3353
rect 3190 3357 3196 3358
rect 3190 3353 3191 3357
rect 3195 3353 3196 3357
rect 3190 3352 3196 3353
rect 3342 3357 3348 3358
rect 3342 3353 3343 3357
rect 3347 3353 3348 3357
rect 3342 3352 3348 3353
rect 3486 3357 3492 3358
rect 3486 3353 3487 3357
rect 3491 3353 3492 3357
rect 3486 3352 3492 3353
rect 3576 3345 3578 3369
rect 3574 3344 3580 3345
rect 3574 3340 3575 3344
rect 3579 3340 3580 3344
rect 3574 3339 3580 3340
rect 3410 3327 3416 3328
rect 3410 3323 3411 3327
rect 3415 3323 3416 3327
rect 3410 3322 3416 3323
rect 3574 3327 3580 3328
rect 3574 3323 3575 3327
rect 3579 3323 3580 3327
rect 3574 3322 3580 3323
rect 3030 3317 3036 3318
rect 3030 3313 3031 3317
rect 3035 3313 3036 3317
rect 3030 3312 3036 3313
rect 3182 3317 3188 3318
rect 3182 3313 3183 3317
rect 3187 3313 3188 3317
rect 3182 3312 3188 3313
rect 3334 3317 3340 3318
rect 3334 3313 3335 3317
rect 3339 3313 3340 3317
rect 3334 3312 3340 3313
rect 3032 3307 3034 3312
rect 3184 3307 3186 3312
rect 3336 3307 3338 3312
rect 2967 3306 2971 3307
rect 2967 3301 2971 3302
rect 3031 3306 3035 3307
rect 3031 3301 3035 3302
rect 3135 3306 3139 3307
rect 3135 3301 3139 3302
rect 3183 3306 3187 3307
rect 3183 3301 3187 3302
rect 3311 3306 3315 3307
rect 3311 3301 3315 3302
rect 3335 3306 3339 3307
rect 3335 3301 3339 3302
rect 2968 3296 2970 3301
rect 3136 3296 3138 3301
rect 3312 3296 3314 3301
rect 2966 3295 2972 3296
rect 2966 3291 2967 3295
rect 2971 3291 2972 3295
rect 2966 3290 2972 3291
rect 3134 3295 3140 3296
rect 3134 3291 3135 3295
rect 3139 3291 3140 3295
rect 3134 3290 3140 3291
rect 3310 3295 3316 3296
rect 3310 3291 3311 3295
rect 3315 3291 3316 3295
rect 3310 3290 3316 3291
rect 2538 3287 2544 3288
rect 2538 3283 2539 3287
rect 2543 3283 2544 3287
rect 2538 3282 2544 3283
rect 2886 3287 2892 3288
rect 2886 3283 2887 3287
rect 2891 3283 2892 3287
rect 2886 3282 2892 3283
rect 2540 3277 2542 3282
rect 2539 3276 2543 3277
rect 2539 3271 2543 3272
rect 2866 3271 2872 3272
rect 2866 3267 2867 3271
rect 2871 3267 2872 3271
rect 2866 3266 2872 3267
rect 3054 3271 3060 3272
rect 3054 3267 3055 3271
rect 3059 3267 3060 3271
rect 3054 3266 3060 3267
rect 2638 3255 2644 3256
rect 2470 3250 2476 3251
rect 2479 3252 2483 3253
rect 2234 3243 2240 3244
rect 2234 3239 2235 3243
rect 2239 3239 2240 3243
rect 2234 3238 2240 3239
rect 2312 3231 2314 3250
rect 2472 3231 2474 3250
rect 2638 3251 2639 3255
rect 2643 3251 2644 3255
rect 2638 3250 2644 3251
rect 2806 3255 2812 3256
rect 2806 3251 2807 3255
rect 2811 3251 2812 3255
rect 2806 3250 2812 3251
rect 2479 3247 2483 3248
rect 2640 3231 2642 3250
rect 2808 3231 2810 3250
rect 2868 3244 2870 3266
rect 2974 3255 2980 3256
rect 2974 3251 2975 3255
rect 2979 3251 2980 3255
rect 2974 3250 2980 3251
rect 2866 3243 2872 3244
rect 2866 3239 2867 3243
rect 2871 3239 2872 3243
rect 2866 3238 2872 3239
rect 2976 3231 2978 3250
rect 3056 3244 3058 3266
rect 3142 3255 3148 3256
rect 3142 3251 3143 3255
rect 3147 3251 3148 3255
rect 3142 3250 3148 3251
rect 3318 3255 3324 3256
rect 3318 3251 3319 3255
rect 3323 3251 3324 3255
rect 3318 3250 3324 3251
rect 3054 3243 3060 3244
rect 3054 3239 3055 3243
rect 3059 3239 3060 3243
rect 3054 3238 3060 3239
rect 3144 3231 3146 3250
rect 3258 3243 3264 3244
rect 3258 3239 3259 3243
rect 3263 3239 3264 3243
rect 3258 3238 3264 3239
rect 2311 3230 2315 3231
rect 2311 3225 2315 3226
rect 2327 3230 2331 3231
rect 2327 3225 2331 3226
rect 2463 3230 2467 3231
rect 2463 3225 2467 3226
rect 2471 3230 2475 3231
rect 2471 3225 2475 3226
rect 2599 3230 2603 3231
rect 2599 3225 2603 3226
rect 2639 3230 2643 3231
rect 2639 3225 2643 3226
rect 2735 3230 2739 3231
rect 2735 3225 2739 3226
rect 2807 3230 2811 3231
rect 2807 3225 2811 3226
rect 2871 3230 2875 3231
rect 2871 3225 2875 3226
rect 2975 3230 2979 3231
rect 2975 3225 2979 3226
rect 3015 3230 3019 3231
rect 3015 3225 3019 3226
rect 3143 3230 3147 3231
rect 3143 3225 3147 3226
rect 3167 3230 3171 3231
rect 3167 3225 3171 3226
rect 2182 3223 2188 3224
rect 2182 3219 2183 3223
rect 2187 3219 2188 3223
rect 2182 3218 2188 3219
rect 2242 3223 2248 3224
rect 2242 3219 2243 3223
rect 2247 3219 2248 3223
rect 2242 3218 2248 3219
rect 2174 3213 2180 3214
rect 2174 3209 2175 3213
rect 2179 3209 2180 3213
rect 2174 3208 2180 3209
rect 2244 3200 2246 3218
rect 2328 3214 2330 3225
rect 2398 3223 2404 3224
rect 2398 3219 2399 3223
rect 2403 3219 2404 3223
rect 2398 3218 2404 3219
rect 2326 3213 2332 3214
rect 2326 3209 2327 3213
rect 2331 3209 2332 3213
rect 2326 3208 2332 3209
rect 2400 3200 2402 3218
rect 2464 3214 2466 3225
rect 2526 3223 2532 3224
rect 2526 3219 2527 3223
rect 2531 3219 2532 3223
rect 2526 3218 2532 3219
rect 2462 3213 2468 3214
rect 2462 3209 2463 3213
rect 2467 3209 2468 3213
rect 2462 3208 2468 3209
rect 2528 3200 2530 3218
rect 2600 3214 2602 3225
rect 2736 3214 2738 3225
rect 2790 3223 2796 3224
rect 2790 3219 2791 3223
rect 2795 3219 2796 3223
rect 2790 3218 2796 3219
rect 2598 3213 2604 3214
rect 2598 3209 2599 3213
rect 2603 3209 2604 3213
rect 2598 3208 2604 3209
rect 2734 3213 2740 3214
rect 2734 3209 2735 3213
rect 2739 3209 2740 3213
rect 2734 3208 2740 3209
rect 2242 3199 2248 3200
rect 2242 3195 2243 3199
rect 2247 3195 2248 3199
rect 2242 3194 2248 3195
rect 2398 3199 2404 3200
rect 2398 3195 2399 3199
rect 2403 3195 2404 3199
rect 2398 3194 2404 3195
rect 2526 3199 2532 3200
rect 2526 3195 2527 3199
rect 2531 3195 2532 3199
rect 2526 3194 2532 3195
rect 2530 3183 2536 3184
rect 2530 3179 2531 3183
rect 2535 3179 2536 3183
rect 2530 3178 2536 3179
rect 2166 3173 2172 3174
rect 2166 3169 2167 3173
rect 2171 3169 2172 3173
rect 2166 3168 2172 3169
rect 2318 3173 2324 3174
rect 2318 3169 2319 3173
rect 2323 3169 2324 3173
rect 2318 3168 2324 3169
rect 2454 3173 2460 3174
rect 2454 3169 2455 3173
rect 2459 3169 2460 3173
rect 2454 3168 2460 3169
rect 2168 3159 2170 3168
rect 2320 3159 2322 3168
rect 2456 3159 2458 3168
rect 2047 3158 2051 3159
rect 2047 3153 2051 3154
rect 2167 3158 2171 3159
rect 2167 3153 2171 3154
rect 2199 3158 2203 3159
rect 2199 3153 2203 3154
rect 2319 3158 2323 3159
rect 2319 3153 2323 3154
rect 2351 3158 2355 3159
rect 2351 3153 2355 3154
rect 2455 3158 2459 3159
rect 2455 3153 2459 3154
rect 2511 3158 2515 3159
rect 2511 3153 2515 3154
rect 2048 3148 2050 3153
rect 2200 3148 2202 3153
rect 2352 3148 2354 3153
rect 2512 3148 2514 3153
rect 2046 3147 2052 3148
rect 2046 3143 2047 3147
rect 2051 3143 2052 3147
rect 2046 3142 2052 3143
rect 2198 3147 2204 3148
rect 2198 3143 2199 3147
rect 2203 3143 2204 3147
rect 2198 3142 2204 3143
rect 2350 3147 2356 3148
rect 2350 3143 2351 3147
rect 2355 3143 2356 3147
rect 2350 3142 2356 3143
rect 2510 3147 2516 3148
rect 2510 3143 2511 3147
rect 2515 3143 2516 3147
rect 2510 3142 2516 3143
rect 2030 3139 2036 3140
rect 1862 3137 1868 3138
rect 1862 3133 1863 3137
rect 1867 3133 1868 3137
rect 2030 3135 2031 3139
rect 2035 3135 2036 3139
rect 2030 3134 2036 3135
rect 1862 3132 1868 3133
rect 1822 3131 1828 3132
rect 1822 3127 1823 3131
rect 1827 3127 1828 3131
rect 1822 3126 1828 3127
rect 1454 3121 1460 3122
rect 1454 3117 1455 3121
rect 1459 3117 1460 3121
rect 1454 3116 1460 3117
rect 1630 3121 1636 3122
rect 1630 3117 1631 3121
rect 1635 3117 1636 3121
rect 1630 3116 1636 3117
rect 1456 3103 1458 3116
rect 1632 3103 1634 3116
rect 1824 3103 1826 3126
rect 1862 3120 1868 3121
rect 1862 3116 1863 3120
rect 1867 3116 1868 3120
rect 1862 3115 1868 3116
rect 1423 3102 1427 3103
rect 1423 3097 1427 3098
rect 1455 3102 1459 3103
rect 1455 3097 1459 3098
rect 1559 3102 1563 3103
rect 1559 3097 1563 3098
rect 1631 3102 1635 3103
rect 1631 3097 1635 3098
rect 1695 3102 1699 3103
rect 1695 3097 1699 3098
rect 1823 3102 1827 3103
rect 1823 3097 1827 3098
rect 1424 3092 1426 3097
rect 1560 3092 1562 3097
rect 1696 3092 1698 3097
rect 1422 3091 1428 3092
rect 1422 3087 1423 3091
rect 1427 3087 1428 3091
rect 1422 3086 1428 3087
rect 1558 3091 1564 3092
rect 1558 3087 1559 3091
rect 1563 3087 1564 3091
rect 1558 3086 1564 3087
rect 1694 3091 1700 3092
rect 1694 3087 1695 3091
rect 1699 3087 1700 3091
rect 1694 3086 1700 3087
rect 1366 3083 1372 3084
rect 1366 3079 1367 3083
rect 1371 3079 1372 3083
rect 1824 3082 1826 3097
rect 1864 3083 1866 3115
rect 1894 3107 1900 3108
rect 1894 3103 1895 3107
rect 1899 3103 1900 3107
rect 1894 3102 1900 3103
rect 2054 3107 2060 3108
rect 2054 3103 2055 3107
rect 2059 3103 2060 3107
rect 2054 3102 2060 3103
rect 2206 3107 2212 3108
rect 2206 3103 2207 3107
rect 2211 3103 2212 3107
rect 2206 3102 2212 3103
rect 2358 3107 2364 3108
rect 2358 3103 2359 3107
rect 2363 3103 2364 3107
rect 2358 3102 2364 3103
rect 2518 3107 2524 3108
rect 2518 3103 2519 3107
rect 2523 3103 2524 3107
rect 2518 3102 2524 3103
rect 1896 3083 1898 3102
rect 2056 3083 2058 3102
rect 2208 3083 2210 3102
rect 2215 3100 2219 3101
rect 2214 3095 2220 3096
rect 2214 3091 2215 3095
rect 2219 3091 2220 3095
rect 2214 3090 2220 3091
rect 2360 3083 2362 3102
rect 2520 3083 2522 3102
rect 2532 3101 2534 3178
rect 2590 3173 2596 3174
rect 2590 3169 2591 3173
rect 2595 3169 2596 3173
rect 2590 3168 2596 3169
rect 2726 3173 2732 3174
rect 2726 3169 2727 3173
rect 2731 3169 2732 3173
rect 2726 3168 2732 3169
rect 2592 3159 2594 3168
rect 2728 3159 2730 3168
rect 2591 3158 2595 3159
rect 2591 3153 2595 3154
rect 2679 3158 2683 3159
rect 2679 3153 2683 3154
rect 2727 3158 2731 3159
rect 2727 3153 2731 3154
rect 2680 3148 2682 3153
rect 2678 3147 2684 3148
rect 2678 3143 2679 3147
rect 2683 3143 2684 3147
rect 2678 3142 2684 3143
rect 2792 3140 2794 3218
rect 2872 3214 2874 3225
rect 2942 3223 2948 3224
rect 2942 3219 2943 3223
rect 2947 3219 2948 3223
rect 2942 3218 2948 3219
rect 2870 3213 2876 3214
rect 2870 3209 2871 3213
rect 2875 3209 2876 3213
rect 2870 3208 2876 3209
rect 2944 3200 2946 3218
rect 3016 3214 3018 3225
rect 3082 3223 3088 3224
rect 3082 3219 3083 3223
rect 3087 3219 3088 3223
rect 3082 3218 3088 3219
rect 3014 3213 3020 3214
rect 3014 3209 3015 3213
rect 3019 3209 3020 3213
rect 3014 3208 3020 3209
rect 3084 3200 3086 3218
rect 3168 3214 3170 3225
rect 3250 3223 3256 3224
rect 3250 3219 3251 3223
rect 3255 3219 3256 3223
rect 3250 3218 3256 3219
rect 3166 3213 3172 3214
rect 3166 3209 3167 3213
rect 3171 3209 3172 3213
rect 3166 3208 3172 3209
rect 3252 3200 3254 3218
rect 2942 3199 2948 3200
rect 2942 3195 2943 3199
rect 2947 3195 2948 3199
rect 2942 3194 2948 3195
rect 3082 3199 3088 3200
rect 3082 3195 3083 3199
rect 3087 3195 3088 3199
rect 3082 3194 3088 3195
rect 3250 3199 3256 3200
rect 3250 3195 3251 3199
rect 3255 3195 3256 3199
rect 3260 3196 3262 3238
rect 3320 3231 3322 3250
rect 3412 3244 3414 3322
rect 3478 3317 3484 3318
rect 3478 3313 3479 3317
rect 3483 3313 3484 3317
rect 3478 3312 3484 3313
rect 3480 3307 3482 3312
rect 3576 3307 3578 3322
rect 3479 3306 3483 3307
rect 3479 3301 3483 3302
rect 3575 3306 3579 3307
rect 3575 3301 3579 3302
rect 3480 3296 3482 3301
rect 3478 3295 3484 3296
rect 3478 3291 3479 3295
rect 3483 3291 3484 3295
rect 3478 3290 3484 3291
rect 3576 3286 3578 3301
rect 3574 3285 3580 3286
rect 3478 3283 3484 3284
rect 3478 3279 3479 3283
rect 3483 3279 3484 3283
rect 3574 3281 3575 3285
rect 3579 3281 3580 3285
rect 3574 3280 3580 3281
rect 3478 3278 3484 3279
rect 3410 3243 3416 3244
rect 3410 3239 3411 3243
rect 3415 3239 3416 3243
rect 3410 3238 3416 3239
rect 3319 3230 3323 3231
rect 3319 3225 3323 3226
rect 3327 3230 3331 3231
rect 3327 3225 3331 3226
rect 3328 3214 3330 3225
rect 3480 3224 3482 3278
rect 3574 3268 3580 3269
rect 3574 3264 3575 3268
rect 3579 3264 3580 3268
rect 3574 3263 3580 3264
rect 3486 3255 3492 3256
rect 3486 3251 3487 3255
rect 3491 3251 3492 3255
rect 3486 3250 3492 3251
rect 3488 3231 3490 3250
rect 3576 3231 3578 3263
rect 3487 3230 3491 3231
rect 3487 3225 3491 3226
rect 3575 3230 3579 3231
rect 3575 3225 3579 3226
rect 3478 3223 3484 3224
rect 3478 3219 3479 3223
rect 3483 3219 3484 3223
rect 3478 3218 3484 3219
rect 3488 3214 3490 3225
rect 3326 3213 3332 3214
rect 3326 3209 3327 3213
rect 3331 3209 3332 3213
rect 3326 3208 3332 3209
rect 3486 3213 3492 3214
rect 3486 3209 3487 3213
rect 3491 3209 3492 3213
rect 3486 3208 3492 3209
rect 3576 3201 3578 3225
rect 3574 3200 3580 3201
rect 3574 3196 3575 3200
rect 3579 3196 3580 3200
rect 3250 3194 3256 3195
rect 3258 3195 3264 3196
rect 3574 3195 3580 3196
rect 3258 3191 3259 3195
rect 3263 3191 3264 3195
rect 3258 3190 3264 3191
rect 3574 3183 3580 3184
rect 3574 3179 3575 3183
rect 3579 3179 3580 3183
rect 3574 3178 3580 3179
rect 2862 3173 2868 3174
rect 2862 3169 2863 3173
rect 2867 3169 2868 3173
rect 2862 3168 2868 3169
rect 3006 3173 3012 3174
rect 3006 3169 3007 3173
rect 3011 3169 3012 3173
rect 3006 3168 3012 3169
rect 3158 3173 3164 3174
rect 3158 3169 3159 3173
rect 3163 3169 3164 3173
rect 3158 3168 3164 3169
rect 3318 3173 3324 3174
rect 3318 3169 3319 3173
rect 3323 3169 3324 3173
rect 3318 3168 3324 3169
rect 3478 3173 3484 3174
rect 3478 3169 3479 3173
rect 3483 3169 3484 3173
rect 3478 3168 3484 3169
rect 2864 3159 2866 3168
rect 3008 3159 3010 3168
rect 3160 3159 3162 3168
rect 3320 3159 3322 3168
rect 3480 3159 3482 3168
rect 3576 3159 3578 3178
rect 2863 3158 2867 3159
rect 2863 3153 2867 3154
rect 2871 3158 2875 3159
rect 2871 3153 2875 3154
rect 3007 3158 3011 3159
rect 3007 3153 3011 3154
rect 3071 3158 3075 3159
rect 3071 3153 3075 3154
rect 3159 3158 3163 3159
rect 3159 3153 3163 3154
rect 3287 3158 3291 3159
rect 3287 3153 3291 3154
rect 3319 3158 3323 3159
rect 3319 3153 3323 3154
rect 3479 3158 3483 3159
rect 3479 3153 3483 3154
rect 3575 3158 3579 3159
rect 3575 3153 3579 3154
rect 2872 3148 2874 3153
rect 3072 3148 3074 3153
rect 3288 3148 3290 3153
rect 3480 3148 3482 3153
rect 2870 3147 2876 3148
rect 2870 3143 2871 3147
rect 2875 3143 2876 3147
rect 2870 3142 2876 3143
rect 3070 3147 3076 3148
rect 3070 3143 3071 3147
rect 3075 3143 3076 3147
rect 3070 3142 3076 3143
rect 3286 3147 3292 3148
rect 3286 3143 3287 3147
rect 3291 3143 3292 3147
rect 3286 3142 3292 3143
rect 3478 3147 3484 3148
rect 3478 3143 3479 3147
rect 3483 3143 3484 3147
rect 3478 3142 3484 3143
rect 2790 3139 2796 3140
rect 2790 3135 2791 3139
rect 2795 3135 2796 3139
rect 3576 3138 3578 3153
rect 2790 3134 2796 3135
rect 3574 3137 3580 3138
rect 3574 3133 3575 3137
rect 3579 3133 3580 3137
rect 3574 3132 3580 3133
rect 2746 3123 2752 3124
rect 2746 3119 2747 3123
rect 2751 3119 2752 3123
rect 2746 3118 2752 3119
rect 2938 3123 2944 3124
rect 2938 3119 2939 3123
rect 2943 3119 2944 3123
rect 2938 3118 2944 3119
rect 3470 3123 3476 3124
rect 3470 3119 3471 3123
rect 3475 3119 3476 3123
rect 3470 3118 3476 3119
rect 3574 3120 3580 3121
rect 2686 3107 2692 3108
rect 2686 3103 2687 3107
rect 2691 3103 2692 3107
rect 2686 3102 2692 3103
rect 2531 3100 2535 3101
rect 2531 3095 2535 3096
rect 2688 3083 2690 3102
rect 1863 3082 1867 3083
rect 1366 3078 1372 3079
rect 1822 3081 1828 3082
rect 1822 3077 1823 3081
rect 1827 3077 1828 3081
rect 1863 3077 1867 3078
rect 1895 3082 1899 3083
rect 1895 3077 1899 3078
rect 1919 3082 1923 3083
rect 1919 3077 1923 3078
rect 2055 3082 2059 3083
rect 2055 3077 2059 3078
rect 2087 3082 2091 3083
rect 2087 3077 2091 3078
rect 2207 3082 2211 3083
rect 2207 3077 2211 3078
rect 2279 3082 2283 3083
rect 2279 3077 2283 3078
rect 2359 3082 2363 3083
rect 2359 3077 2363 3078
rect 2487 3082 2491 3083
rect 2487 3077 2491 3078
rect 2519 3082 2523 3083
rect 2519 3077 2523 3078
rect 2687 3082 2691 3083
rect 2687 3077 2691 3078
rect 2719 3082 2723 3083
rect 2719 3077 2723 3078
rect 110 3076 116 3077
rect 567 3076 571 3077
rect 567 3071 571 3072
rect 891 3076 895 3077
rect 1822 3076 1828 3077
rect 891 3071 895 3072
rect 110 3064 116 3065
rect 110 3060 111 3064
rect 115 3060 116 3064
rect 110 3059 116 3060
rect 112 3031 114 3059
rect 558 3051 564 3052
rect 558 3047 559 3051
rect 563 3047 564 3051
rect 558 3046 564 3047
rect 560 3031 562 3046
rect 568 3040 570 3071
rect 1762 3067 1768 3068
rect 1762 3063 1763 3067
rect 1767 3063 1768 3067
rect 1762 3062 1768 3063
rect 1822 3064 1828 3065
rect 670 3051 676 3052
rect 670 3047 671 3051
rect 675 3047 676 3051
rect 670 3046 676 3047
rect 790 3051 796 3052
rect 790 3047 791 3051
rect 795 3047 796 3051
rect 790 3046 796 3047
rect 910 3051 916 3052
rect 910 3047 911 3051
rect 915 3047 916 3051
rect 910 3046 916 3047
rect 1038 3051 1044 3052
rect 1038 3047 1039 3051
rect 1043 3047 1044 3051
rect 1038 3046 1044 3047
rect 1166 3051 1172 3052
rect 1166 3047 1167 3051
rect 1171 3047 1172 3051
rect 1166 3046 1172 3047
rect 1294 3051 1300 3052
rect 1294 3047 1295 3051
rect 1299 3047 1300 3051
rect 1294 3046 1300 3047
rect 1430 3051 1436 3052
rect 1430 3047 1431 3051
rect 1435 3047 1436 3051
rect 1430 3046 1436 3047
rect 1566 3051 1572 3052
rect 1566 3047 1567 3051
rect 1571 3047 1572 3051
rect 1566 3046 1572 3047
rect 1702 3051 1708 3052
rect 1702 3047 1703 3051
rect 1707 3047 1708 3051
rect 1702 3046 1708 3047
rect 566 3039 572 3040
rect 566 3035 567 3039
rect 571 3035 572 3039
rect 566 3034 572 3035
rect 672 3031 674 3046
rect 792 3031 794 3046
rect 912 3031 914 3046
rect 1040 3031 1042 3046
rect 1168 3031 1170 3046
rect 1174 3039 1180 3040
rect 1174 3035 1175 3039
rect 1179 3035 1180 3039
rect 1174 3034 1180 3035
rect 111 3030 115 3031
rect 111 3025 115 3026
rect 559 3030 563 3031
rect 559 3025 563 3026
rect 575 3030 579 3031
rect 575 3025 579 3026
rect 671 3030 675 3031
rect 671 3025 675 3026
rect 703 3030 707 3031
rect 703 3025 707 3026
rect 791 3030 795 3031
rect 791 3025 795 3026
rect 831 3030 835 3031
rect 831 3025 835 3026
rect 911 3030 915 3031
rect 911 3025 915 3026
rect 967 3030 971 3031
rect 967 3025 971 3026
rect 1039 3030 1043 3031
rect 1039 3025 1043 3026
rect 1103 3030 1107 3031
rect 1103 3025 1107 3026
rect 1167 3030 1171 3031
rect 1167 3025 1171 3026
rect 112 3001 114 3025
rect 576 3014 578 3025
rect 704 3014 706 3025
rect 770 3023 776 3024
rect 770 3019 771 3023
rect 775 3019 776 3023
rect 770 3018 776 3019
rect 574 3013 580 3014
rect 574 3009 575 3013
rect 579 3009 580 3013
rect 574 3008 580 3009
rect 702 3013 708 3014
rect 702 3009 703 3013
rect 707 3009 708 3013
rect 702 3008 708 3009
rect 110 3000 116 3001
rect 110 2996 111 3000
rect 115 2996 116 3000
rect 772 2996 774 3018
rect 832 3014 834 3025
rect 898 3023 904 3024
rect 898 3019 899 3023
rect 903 3019 904 3023
rect 898 3018 904 3019
rect 830 3013 836 3014
rect 830 3009 831 3013
rect 835 3009 836 3013
rect 830 3008 836 3009
rect 900 2996 902 3018
rect 968 3014 970 3025
rect 1104 3014 1106 3025
rect 966 3013 972 3014
rect 966 3009 967 3013
rect 971 3009 972 3013
rect 966 3008 972 3009
rect 1102 3013 1108 3014
rect 1102 3009 1103 3013
rect 1107 3009 1108 3013
rect 1102 3008 1108 3009
rect 1176 2996 1178 3034
rect 1296 3031 1298 3046
rect 1432 3031 1434 3046
rect 1568 3031 1570 3046
rect 1704 3031 1706 3046
rect 1239 3030 1243 3031
rect 1239 3025 1243 3026
rect 1295 3030 1299 3031
rect 1295 3025 1299 3026
rect 1367 3030 1371 3031
rect 1367 3025 1371 3026
rect 1431 3030 1435 3031
rect 1431 3025 1435 3026
rect 1495 3030 1499 3031
rect 1495 3025 1499 3026
rect 1567 3030 1571 3031
rect 1567 3025 1571 3026
rect 1623 3030 1627 3031
rect 1623 3025 1627 3026
rect 1703 3030 1707 3031
rect 1703 3025 1707 3026
rect 1735 3030 1739 3031
rect 1735 3025 1739 3026
rect 1240 3014 1242 3025
rect 1306 3023 1312 3024
rect 1306 3019 1307 3023
rect 1311 3019 1312 3023
rect 1306 3018 1312 3019
rect 1238 3013 1244 3014
rect 1238 3009 1239 3013
rect 1243 3009 1244 3013
rect 1238 3008 1244 3009
rect 1308 2996 1310 3018
rect 1368 3014 1370 3025
rect 1438 3023 1444 3024
rect 1438 3019 1439 3023
rect 1443 3019 1444 3023
rect 1438 3018 1444 3019
rect 1366 3013 1372 3014
rect 1366 3009 1367 3013
rect 1371 3009 1372 3013
rect 1366 3008 1372 3009
rect 1440 2996 1442 3018
rect 1496 3014 1498 3025
rect 1594 3023 1600 3024
rect 1594 3019 1595 3023
rect 1599 3019 1600 3023
rect 1594 3018 1600 3019
rect 1494 3013 1500 3014
rect 1494 3009 1495 3013
rect 1499 3009 1500 3013
rect 1494 3008 1500 3009
rect 110 2995 116 2996
rect 770 2995 776 2996
rect 770 2991 771 2995
rect 775 2991 776 2995
rect 770 2990 776 2991
rect 898 2995 904 2996
rect 898 2991 899 2995
rect 903 2991 904 2995
rect 898 2990 904 2991
rect 1174 2995 1180 2996
rect 1174 2991 1175 2995
rect 1179 2991 1180 2995
rect 1174 2990 1180 2991
rect 1306 2995 1312 2996
rect 1306 2991 1307 2995
rect 1311 2991 1312 2995
rect 1306 2990 1312 2991
rect 1438 2995 1444 2996
rect 1438 2991 1439 2995
rect 1443 2991 1444 2995
rect 1438 2990 1444 2991
rect 110 2983 116 2984
rect 110 2979 111 2983
rect 115 2979 116 2983
rect 110 2978 116 2979
rect 510 2983 516 2984
rect 510 2979 511 2983
rect 515 2979 516 2983
rect 510 2978 516 2979
rect 112 2963 114 2978
rect 111 2962 115 2963
rect 111 2957 115 2958
rect 495 2962 499 2963
rect 495 2957 499 2958
rect 112 2942 114 2957
rect 496 2952 498 2957
rect 494 2951 500 2952
rect 494 2947 495 2951
rect 499 2947 500 2951
rect 494 2946 500 2947
rect 110 2941 116 2942
rect 110 2937 111 2941
rect 115 2937 116 2941
rect 110 2936 116 2937
rect 110 2924 116 2925
rect 110 2920 111 2924
rect 115 2920 116 2924
rect 110 2919 116 2920
rect 112 2891 114 2919
rect 502 2911 508 2912
rect 502 2907 503 2911
rect 507 2907 508 2911
rect 502 2906 508 2907
rect 504 2891 506 2906
rect 512 2900 514 2978
rect 566 2973 572 2974
rect 566 2969 567 2973
rect 571 2969 572 2973
rect 566 2968 572 2969
rect 694 2973 700 2974
rect 694 2969 695 2973
rect 699 2969 700 2973
rect 694 2968 700 2969
rect 822 2973 828 2974
rect 822 2969 823 2973
rect 827 2969 828 2973
rect 822 2968 828 2969
rect 958 2973 964 2974
rect 958 2969 959 2973
rect 963 2969 964 2973
rect 958 2968 964 2969
rect 1094 2973 1100 2974
rect 1094 2969 1095 2973
rect 1099 2969 1100 2973
rect 1094 2968 1100 2969
rect 1230 2973 1236 2974
rect 1230 2969 1231 2973
rect 1235 2969 1236 2973
rect 1230 2968 1236 2969
rect 1358 2973 1364 2974
rect 1358 2969 1359 2973
rect 1363 2969 1364 2973
rect 1358 2968 1364 2969
rect 1486 2973 1492 2974
rect 1486 2969 1487 2973
rect 1491 2969 1492 2973
rect 1486 2968 1492 2969
rect 568 2963 570 2968
rect 696 2963 698 2968
rect 824 2963 826 2968
rect 960 2963 962 2968
rect 1096 2963 1098 2968
rect 1232 2963 1234 2968
rect 1360 2963 1362 2968
rect 1488 2963 1490 2968
rect 567 2962 571 2963
rect 567 2957 571 2958
rect 639 2962 643 2963
rect 639 2957 643 2958
rect 695 2962 699 2963
rect 695 2957 699 2958
rect 783 2962 787 2963
rect 783 2957 787 2958
rect 823 2962 827 2963
rect 823 2957 827 2958
rect 919 2962 923 2963
rect 919 2957 923 2958
rect 959 2962 963 2963
rect 959 2957 963 2958
rect 1055 2962 1059 2963
rect 1055 2957 1059 2958
rect 1095 2962 1099 2963
rect 1095 2957 1099 2958
rect 1183 2962 1187 2963
rect 1183 2957 1187 2958
rect 1231 2962 1235 2963
rect 1231 2957 1235 2958
rect 1303 2962 1307 2963
rect 1303 2957 1307 2958
rect 1359 2962 1363 2963
rect 1359 2957 1363 2958
rect 1415 2962 1419 2963
rect 1415 2957 1419 2958
rect 1487 2962 1491 2963
rect 1487 2957 1491 2958
rect 1527 2962 1531 2963
rect 1527 2957 1531 2958
rect 640 2952 642 2957
rect 784 2952 786 2957
rect 920 2952 922 2957
rect 1056 2952 1058 2957
rect 1184 2952 1186 2957
rect 1304 2952 1306 2957
rect 1416 2952 1418 2957
rect 1528 2952 1530 2957
rect 638 2951 644 2952
rect 638 2947 639 2951
rect 643 2947 644 2951
rect 638 2946 644 2947
rect 782 2951 788 2952
rect 782 2947 783 2951
rect 787 2947 788 2951
rect 782 2946 788 2947
rect 918 2951 924 2952
rect 918 2947 919 2951
rect 923 2947 924 2951
rect 918 2946 924 2947
rect 1054 2951 1060 2952
rect 1054 2947 1055 2951
rect 1059 2947 1060 2951
rect 1054 2946 1060 2947
rect 1182 2951 1188 2952
rect 1182 2947 1183 2951
rect 1187 2947 1188 2951
rect 1182 2946 1188 2947
rect 1302 2951 1308 2952
rect 1302 2947 1303 2951
rect 1307 2947 1308 2951
rect 1302 2946 1308 2947
rect 1414 2951 1420 2952
rect 1414 2947 1415 2951
rect 1419 2947 1420 2951
rect 1414 2946 1420 2947
rect 1526 2951 1532 2952
rect 1526 2947 1527 2951
rect 1531 2947 1532 2951
rect 1526 2946 1532 2947
rect 1596 2944 1598 3018
rect 1624 3014 1626 3025
rect 1736 3014 1738 3025
rect 1764 3024 1766 3062
rect 1822 3060 1823 3064
rect 1827 3060 1828 3064
rect 1822 3059 1828 3060
rect 1824 3031 1826 3059
rect 1864 3053 1866 3077
rect 1920 3066 1922 3077
rect 2006 3075 2012 3076
rect 2006 3071 2007 3075
rect 2011 3071 2012 3075
rect 2006 3070 2012 3071
rect 1918 3065 1924 3066
rect 1918 3061 1919 3065
rect 1923 3061 1924 3065
rect 1918 3060 1924 3061
rect 1862 3052 1868 3053
rect 1862 3048 1863 3052
rect 1867 3048 1868 3052
rect 2008 3048 2010 3070
rect 2088 3066 2090 3077
rect 2182 3075 2188 3076
rect 2182 3071 2183 3075
rect 2187 3071 2188 3075
rect 2182 3070 2188 3071
rect 2086 3065 2092 3066
rect 2086 3061 2087 3065
rect 2091 3061 2092 3065
rect 2086 3060 2092 3061
rect 2184 3048 2186 3070
rect 2280 3066 2282 3077
rect 2488 3066 2490 3077
rect 2502 3075 2508 3076
rect 2502 3071 2503 3075
rect 2507 3071 2508 3075
rect 2502 3070 2508 3071
rect 2278 3065 2284 3066
rect 2278 3061 2279 3065
rect 2283 3061 2284 3065
rect 2278 3060 2284 3061
rect 2486 3065 2492 3066
rect 2486 3061 2487 3065
rect 2491 3061 2492 3065
rect 2486 3060 2492 3061
rect 2504 3053 2506 3070
rect 2720 3066 2722 3077
rect 2748 3076 2750 3118
rect 2878 3107 2884 3108
rect 2878 3103 2879 3107
rect 2883 3103 2884 3107
rect 2878 3102 2884 3103
rect 2880 3083 2882 3102
rect 2940 3096 2942 3118
rect 3078 3107 3084 3108
rect 3078 3103 3079 3107
rect 3083 3103 3084 3107
rect 3078 3102 3084 3103
rect 3294 3107 3300 3108
rect 3294 3103 3295 3107
rect 3299 3103 3300 3107
rect 3294 3102 3300 3103
rect 2938 3095 2944 3096
rect 2938 3091 2939 3095
rect 2943 3091 2944 3095
rect 2938 3090 2944 3091
rect 3080 3083 3082 3102
rect 3296 3083 3298 3102
rect 3302 3095 3308 3096
rect 3302 3091 3303 3095
rect 3307 3091 3308 3095
rect 3302 3090 3308 3091
rect 2879 3082 2883 3083
rect 2879 3077 2883 3078
rect 2975 3082 2979 3083
rect 2975 3077 2979 3078
rect 3079 3082 3083 3083
rect 3079 3077 3083 3078
rect 3239 3082 3243 3083
rect 3239 3077 3243 3078
rect 3295 3082 3299 3083
rect 3295 3077 3299 3078
rect 2746 3075 2752 3076
rect 2746 3071 2747 3075
rect 2751 3071 2752 3075
rect 2746 3070 2752 3071
rect 2976 3066 2978 3077
rect 3240 3066 3242 3077
rect 3246 3075 3252 3076
rect 3246 3071 3247 3075
rect 3251 3071 3252 3075
rect 3246 3070 3252 3071
rect 2718 3065 2724 3066
rect 2718 3061 2719 3065
rect 2723 3061 2724 3065
rect 2718 3060 2724 3061
rect 2974 3065 2980 3066
rect 2974 3061 2975 3065
rect 2979 3061 2980 3065
rect 2974 3060 2980 3061
rect 3238 3065 3244 3066
rect 3238 3061 3239 3065
rect 3243 3061 3244 3065
rect 3238 3060 3244 3061
rect 2503 3052 2507 3053
rect 2899 3052 2903 3053
rect 1862 3047 1868 3048
rect 2006 3047 2012 3048
rect 2006 3043 2007 3047
rect 2011 3043 2012 3047
rect 2006 3042 2012 3043
rect 2182 3047 2188 3048
rect 2503 3047 2507 3048
rect 2898 3047 2904 3048
rect 2182 3043 2183 3047
rect 2187 3043 2188 3047
rect 2182 3042 2188 3043
rect 2898 3043 2899 3047
rect 2903 3043 2904 3047
rect 2898 3042 2904 3043
rect 1862 3035 1868 3036
rect 1862 3031 1863 3035
rect 1867 3031 1868 3035
rect 1823 3030 1827 3031
rect 1862 3030 1868 3031
rect 2430 3035 2436 3036
rect 2430 3031 2431 3035
rect 2435 3031 2436 3035
rect 2430 3030 2436 3031
rect 1823 3025 1827 3026
rect 1762 3023 1768 3024
rect 1762 3019 1763 3023
rect 1767 3019 1768 3023
rect 1762 3018 1768 3019
rect 1622 3013 1628 3014
rect 1622 3009 1623 3013
rect 1627 3009 1628 3013
rect 1622 3008 1628 3009
rect 1734 3013 1740 3014
rect 1734 3009 1735 3013
rect 1739 3009 1740 3013
rect 1734 3008 1740 3009
rect 1824 3001 1826 3025
rect 1864 3011 1866 3030
rect 1910 3025 1916 3026
rect 1910 3021 1911 3025
rect 1915 3021 1916 3025
rect 1910 3020 1916 3021
rect 2078 3025 2084 3026
rect 2078 3021 2079 3025
rect 2083 3021 2084 3025
rect 2078 3020 2084 3021
rect 2270 3025 2276 3026
rect 2270 3021 2271 3025
rect 2275 3021 2276 3025
rect 2270 3020 2276 3021
rect 1912 3011 1914 3020
rect 2080 3011 2082 3020
rect 2272 3011 2274 3020
rect 1863 3010 1867 3011
rect 1863 3005 1867 3006
rect 1911 3010 1915 3011
rect 1911 3005 1915 3006
rect 2023 3010 2027 3011
rect 2023 3005 2027 3006
rect 2079 3010 2083 3011
rect 2079 3005 2083 3006
rect 2159 3010 2163 3011
rect 2159 3005 2163 3006
rect 2271 3010 2275 3011
rect 2271 3005 2275 3006
rect 2287 3010 2291 3011
rect 2287 3005 2291 3006
rect 2415 3010 2419 3011
rect 2415 3005 2419 3006
rect 1822 3000 1828 3001
rect 1822 2996 1823 3000
rect 1827 2996 1828 3000
rect 1822 2995 1828 2996
rect 1864 2990 1866 3005
rect 2024 3000 2026 3005
rect 2160 3000 2162 3005
rect 2288 3000 2290 3005
rect 2416 3000 2418 3005
rect 2022 2999 2028 3000
rect 2022 2995 2023 2999
rect 2027 2995 2028 2999
rect 2022 2994 2028 2995
rect 2158 2999 2164 3000
rect 2158 2995 2159 2999
rect 2163 2995 2164 2999
rect 2158 2994 2164 2995
rect 2286 2999 2292 3000
rect 2286 2995 2287 2999
rect 2291 2995 2292 2999
rect 2286 2994 2292 2995
rect 2414 2999 2420 3000
rect 2414 2995 2415 2999
rect 2419 2995 2420 2999
rect 2414 2994 2420 2995
rect 1862 2989 1868 2990
rect 1862 2985 1863 2989
rect 1867 2985 1868 2989
rect 1862 2984 1868 2985
rect 1690 2983 1696 2984
rect 1690 2979 1691 2983
rect 1695 2979 1696 2983
rect 1690 2978 1696 2979
rect 1822 2983 1828 2984
rect 1822 2979 1823 2983
rect 1827 2979 1828 2983
rect 1822 2978 1828 2979
rect 1614 2973 1620 2974
rect 1614 2969 1615 2973
rect 1619 2969 1620 2973
rect 1614 2968 1620 2969
rect 1616 2963 1618 2968
rect 1615 2962 1619 2963
rect 1615 2957 1619 2958
rect 1639 2962 1643 2963
rect 1639 2957 1643 2958
rect 1640 2952 1642 2957
rect 1638 2951 1644 2952
rect 1638 2947 1639 2951
rect 1643 2947 1644 2951
rect 1638 2946 1644 2947
rect 1594 2943 1600 2944
rect 1594 2939 1595 2943
rect 1599 2939 1600 2943
rect 1594 2938 1600 2939
rect 630 2927 636 2928
rect 630 2923 631 2927
rect 635 2923 636 2927
rect 630 2922 636 2923
rect 632 2900 634 2922
rect 646 2911 652 2912
rect 646 2907 647 2911
rect 651 2907 652 2911
rect 646 2906 652 2907
rect 790 2911 796 2912
rect 790 2907 791 2911
rect 795 2907 796 2911
rect 790 2906 796 2907
rect 926 2911 932 2912
rect 926 2907 927 2911
rect 931 2907 932 2911
rect 926 2906 932 2907
rect 1062 2911 1068 2912
rect 1062 2907 1063 2911
rect 1067 2907 1068 2911
rect 1062 2906 1068 2907
rect 1190 2911 1196 2912
rect 1190 2907 1191 2911
rect 1195 2907 1196 2911
rect 1190 2906 1196 2907
rect 1310 2911 1316 2912
rect 1310 2907 1311 2911
rect 1315 2907 1316 2911
rect 1310 2906 1316 2907
rect 1422 2911 1428 2912
rect 1422 2907 1423 2911
rect 1427 2907 1428 2911
rect 1422 2906 1428 2907
rect 1534 2911 1540 2912
rect 1534 2907 1535 2911
rect 1539 2907 1540 2911
rect 1534 2906 1540 2907
rect 1646 2911 1652 2912
rect 1646 2907 1647 2911
rect 1651 2907 1652 2911
rect 1646 2906 1652 2907
rect 510 2899 516 2900
rect 510 2895 511 2899
rect 515 2895 516 2899
rect 510 2894 516 2895
rect 630 2899 636 2900
rect 630 2895 631 2899
rect 635 2895 636 2899
rect 630 2894 636 2895
rect 648 2891 650 2906
rect 792 2891 794 2906
rect 928 2891 930 2906
rect 1064 2891 1066 2906
rect 1166 2899 1172 2900
rect 1166 2895 1167 2899
rect 1171 2895 1172 2899
rect 1166 2894 1172 2895
rect 111 2890 115 2891
rect 111 2885 115 2886
rect 327 2890 331 2891
rect 327 2885 331 2886
rect 455 2890 459 2891
rect 455 2885 459 2886
rect 503 2890 507 2891
rect 503 2885 507 2886
rect 591 2890 595 2891
rect 591 2885 595 2886
rect 647 2890 651 2891
rect 647 2885 651 2886
rect 727 2890 731 2891
rect 727 2885 731 2886
rect 791 2890 795 2891
rect 791 2885 795 2886
rect 871 2890 875 2891
rect 871 2885 875 2886
rect 927 2890 931 2891
rect 927 2885 931 2886
rect 1007 2890 1011 2891
rect 1007 2885 1011 2886
rect 1063 2890 1067 2891
rect 1063 2885 1067 2886
rect 1143 2890 1147 2891
rect 1143 2885 1147 2886
rect 112 2861 114 2885
rect 328 2874 330 2885
rect 394 2883 400 2884
rect 394 2879 395 2883
rect 399 2879 400 2883
rect 394 2878 400 2879
rect 326 2873 332 2874
rect 326 2869 327 2873
rect 331 2869 332 2873
rect 326 2868 332 2869
rect 110 2860 116 2861
rect 110 2856 111 2860
rect 115 2856 116 2860
rect 396 2856 398 2878
rect 456 2874 458 2885
rect 522 2883 528 2884
rect 522 2879 523 2883
rect 527 2879 528 2883
rect 522 2878 528 2879
rect 454 2873 460 2874
rect 454 2869 455 2873
rect 459 2869 460 2873
rect 454 2868 460 2869
rect 524 2856 526 2878
rect 592 2874 594 2885
rect 670 2883 676 2884
rect 670 2879 671 2883
rect 675 2879 676 2883
rect 670 2878 676 2879
rect 590 2873 596 2874
rect 590 2869 591 2873
rect 595 2869 596 2873
rect 590 2868 596 2869
rect 672 2856 674 2878
rect 728 2874 730 2885
rect 798 2883 804 2884
rect 798 2879 799 2883
rect 803 2879 804 2883
rect 798 2878 804 2879
rect 726 2873 732 2874
rect 726 2869 727 2873
rect 731 2869 732 2873
rect 726 2868 732 2869
rect 800 2856 802 2878
rect 872 2874 874 2885
rect 1008 2874 1010 2885
rect 1014 2883 1020 2884
rect 1014 2879 1015 2883
rect 1019 2879 1020 2883
rect 1014 2878 1020 2879
rect 870 2873 876 2874
rect 870 2869 871 2873
rect 875 2869 876 2873
rect 870 2868 876 2869
rect 1006 2873 1012 2874
rect 1006 2869 1007 2873
rect 1011 2869 1012 2873
rect 1006 2868 1012 2869
rect 110 2855 116 2856
rect 394 2855 400 2856
rect 394 2851 395 2855
rect 399 2851 400 2855
rect 394 2850 400 2851
rect 522 2855 528 2856
rect 522 2851 523 2855
rect 527 2851 528 2855
rect 522 2850 528 2851
rect 670 2855 676 2856
rect 670 2851 671 2855
rect 675 2851 676 2855
rect 670 2850 676 2851
rect 798 2855 804 2856
rect 798 2851 799 2855
rect 803 2851 804 2855
rect 798 2850 804 2851
rect 110 2843 116 2844
rect 110 2839 111 2843
rect 115 2839 116 2843
rect 110 2838 116 2839
rect 112 2815 114 2838
rect 318 2833 324 2834
rect 318 2829 319 2833
rect 323 2829 324 2833
rect 318 2828 324 2829
rect 446 2833 452 2834
rect 446 2829 447 2833
rect 451 2829 452 2833
rect 446 2828 452 2829
rect 582 2833 588 2834
rect 582 2829 583 2833
rect 587 2829 588 2833
rect 582 2828 588 2829
rect 718 2833 724 2834
rect 718 2829 719 2833
rect 723 2829 724 2833
rect 718 2828 724 2829
rect 862 2833 868 2834
rect 862 2829 863 2833
rect 867 2829 868 2833
rect 862 2828 868 2829
rect 998 2833 1004 2834
rect 998 2829 999 2833
rect 1003 2829 1004 2833
rect 998 2828 1004 2829
rect 320 2815 322 2828
rect 448 2815 450 2828
rect 584 2815 586 2828
rect 720 2815 722 2828
rect 864 2815 866 2828
rect 1000 2815 1002 2828
rect 111 2814 115 2815
rect 111 2809 115 2810
rect 167 2814 171 2815
rect 167 2809 171 2810
rect 295 2814 299 2815
rect 295 2809 299 2810
rect 319 2814 323 2815
rect 319 2809 323 2810
rect 423 2814 427 2815
rect 423 2809 427 2810
rect 447 2814 451 2815
rect 447 2809 451 2810
rect 559 2814 563 2815
rect 559 2809 563 2810
rect 583 2814 587 2815
rect 583 2809 587 2810
rect 695 2814 699 2815
rect 695 2809 699 2810
rect 719 2814 723 2815
rect 719 2809 723 2810
rect 823 2814 827 2815
rect 823 2809 827 2810
rect 863 2814 867 2815
rect 863 2809 867 2810
rect 951 2814 955 2815
rect 951 2809 955 2810
rect 999 2814 1003 2815
rect 1016 2812 1018 2878
rect 1144 2874 1146 2885
rect 1142 2873 1148 2874
rect 1142 2869 1143 2873
rect 1147 2869 1148 2873
rect 1168 2869 1170 2894
rect 1192 2891 1194 2906
rect 1312 2891 1314 2906
rect 1424 2891 1426 2906
rect 1536 2891 1538 2906
rect 1648 2891 1650 2906
rect 1692 2900 1694 2978
rect 1726 2973 1732 2974
rect 1726 2969 1727 2973
rect 1731 2969 1732 2973
rect 1726 2968 1732 2969
rect 1728 2963 1730 2968
rect 1824 2963 1826 2978
rect 1862 2972 1868 2973
rect 1862 2968 1863 2972
rect 1867 2968 1868 2972
rect 1862 2967 1868 2968
rect 1727 2962 1731 2963
rect 1727 2957 1731 2958
rect 1823 2962 1827 2963
rect 1823 2957 1827 2958
rect 1728 2952 1730 2957
rect 1726 2951 1732 2952
rect 1726 2947 1727 2951
rect 1731 2947 1732 2951
rect 1726 2946 1732 2947
rect 1824 2942 1826 2957
rect 1822 2941 1828 2942
rect 1822 2937 1823 2941
rect 1827 2937 1828 2941
rect 1822 2936 1828 2937
rect 1864 2935 1866 2967
rect 2030 2959 2036 2960
rect 2030 2955 2031 2959
rect 2035 2955 2036 2959
rect 2030 2954 2036 2955
rect 2166 2959 2172 2960
rect 2166 2955 2167 2959
rect 2171 2955 2172 2959
rect 2166 2954 2172 2955
rect 2294 2959 2300 2960
rect 2294 2955 2295 2959
rect 2299 2955 2300 2959
rect 2294 2954 2300 2955
rect 2422 2959 2428 2960
rect 2422 2955 2423 2959
rect 2427 2955 2428 2959
rect 2422 2954 2428 2955
rect 2032 2935 2034 2954
rect 2168 2935 2170 2954
rect 2296 2935 2298 2954
rect 2424 2935 2426 2954
rect 2432 2948 2434 3030
rect 2478 3025 2484 3026
rect 2478 3021 2479 3025
rect 2483 3021 2484 3025
rect 2478 3020 2484 3021
rect 2710 3025 2716 3026
rect 2710 3021 2711 3025
rect 2715 3021 2716 3025
rect 2710 3020 2716 3021
rect 2966 3025 2972 3026
rect 2966 3021 2967 3025
rect 2971 3021 2972 3025
rect 2966 3020 2972 3021
rect 3230 3025 3236 3026
rect 3230 3021 3231 3025
rect 3235 3021 3236 3025
rect 3230 3020 3236 3021
rect 2480 3011 2482 3020
rect 2712 3011 2714 3020
rect 2968 3011 2970 3020
rect 3232 3011 3234 3020
rect 2479 3010 2483 3011
rect 2479 3005 2483 3006
rect 2535 3010 2539 3011
rect 2535 3005 2539 3006
rect 2663 3010 2667 3011
rect 2663 3005 2667 3006
rect 2711 3010 2715 3011
rect 2711 3005 2715 3006
rect 2807 3010 2811 3011
rect 2807 3005 2811 3006
rect 2967 3010 2971 3011
rect 2967 3005 2971 3006
rect 3143 3010 3147 3011
rect 3143 3005 3147 3006
rect 3231 3010 3235 3011
rect 3231 3005 3235 3006
rect 2536 3000 2538 3005
rect 2664 3000 2666 3005
rect 2808 3000 2810 3005
rect 2968 3000 2970 3005
rect 3144 3000 3146 3005
rect 2534 2999 2540 3000
rect 2534 2995 2535 2999
rect 2539 2995 2540 2999
rect 2534 2994 2540 2995
rect 2662 2999 2668 3000
rect 2662 2995 2663 2999
rect 2667 2995 2668 2999
rect 2662 2994 2668 2995
rect 2806 2999 2812 3000
rect 2806 2995 2807 2999
rect 2811 2995 2812 2999
rect 2806 2994 2812 2995
rect 2966 2999 2972 3000
rect 2966 2995 2967 2999
rect 2971 2995 2972 2999
rect 2966 2994 2972 2995
rect 3142 2999 3148 3000
rect 3142 2995 3143 2999
rect 3147 2995 3148 2999
rect 3142 2994 3148 2995
rect 3248 2992 3250 3070
rect 3304 3052 3306 3090
rect 3472 3076 3474 3118
rect 3574 3116 3575 3120
rect 3579 3116 3580 3120
rect 3574 3115 3580 3116
rect 3486 3107 3492 3108
rect 3486 3103 3487 3107
rect 3491 3103 3492 3107
rect 3486 3102 3492 3103
rect 3488 3083 3490 3102
rect 3576 3083 3578 3115
rect 3487 3082 3491 3083
rect 3487 3077 3491 3078
rect 3575 3082 3579 3083
rect 3575 3077 3579 3078
rect 3470 3075 3476 3076
rect 3470 3071 3471 3075
rect 3475 3071 3476 3075
rect 3470 3070 3476 3071
rect 3488 3066 3490 3077
rect 3486 3065 3492 3066
rect 3486 3061 3487 3065
rect 3491 3061 3492 3065
rect 3486 3060 3492 3061
rect 3576 3053 3578 3077
rect 3574 3052 3580 3053
rect 3302 3051 3308 3052
rect 3302 3047 3303 3051
rect 3307 3047 3308 3051
rect 3574 3048 3575 3052
rect 3579 3048 3580 3052
rect 3574 3047 3580 3048
rect 3302 3046 3308 3047
rect 3574 3035 3580 3036
rect 3574 3031 3575 3035
rect 3579 3031 3580 3035
rect 3574 3030 3580 3031
rect 3478 3025 3484 3026
rect 3478 3021 3479 3025
rect 3483 3021 3484 3025
rect 3478 3020 3484 3021
rect 3480 3011 3482 3020
rect 3576 3011 3578 3030
rect 3319 3010 3323 3011
rect 3319 3005 3323 3006
rect 3479 3010 3483 3011
rect 3479 3005 3483 3006
rect 3575 3010 3579 3011
rect 3575 3005 3579 3006
rect 3320 3000 3322 3005
rect 3480 3000 3482 3005
rect 3318 2999 3324 3000
rect 3318 2995 3319 2999
rect 3323 2995 3324 2999
rect 3318 2994 3324 2995
rect 3478 2999 3484 3000
rect 3478 2995 3479 2999
rect 3483 2995 3484 2999
rect 3478 2994 3484 2995
rect 3246 2991 3252 2992
rect 3246 2987 3247 2991
rect 3251 2987 3252 2991
rect 3576 2990 3578 3005
rect 3246 2986 3252 2987
rect 3574 2989 3580 2990
rect 3574 2985 3575 2989
rect 3579 2985 3580 2989
rect 3574 2984 3580 2985
rect 3470 2975 3476 2976
rect 3470 2971 3471 2975
rect 3475 2971 3476 2975
rect 3470 2970 3476 2971
rect 3574 2972 3580 2973
rect 2542 2959 2548 2960
rect 2542 2955 2543 2959
rect 2547 2955 2548 2959
rect 2542 2954 2548 2955
rect 2670 2959 2676 2960
rect 2670 2955 2671 2959
rect 2675 2955 2676 2959
rect 2670 2954 2676 2955
rect 2814 2959 2820 2960
rect 2814 2955 2815 2959
rect 2819 2955 2820 2959
rect 2814 2954 2820 2955
rect 2974 2959 2980 2960
rect 2974 2955 2975 2959
rect 2979 2955 2980 2959
rect 2974 2954 2980 2955
rect 3150 2959 3156 2960
rect 3150 2955 3151 2959
rect 3155 2955 3156 2959
rect 3150 2954 3156 2955
rect 3326 2959 3332 2960
rect 3326 2955 3327 2959
rect 3331 2955 3332 2959
rect 3326 2954 3332 2955
rect 2430 2947 2436 2948
rect 2430 2943 2431 2947
rect 2435 2943 2436 2947
rect 2430 2942 2436 2943
rect 2544 2935 2546 2954
rect 2672 2935 2674 2954
rect 2816 2935 2818 2954
rect 2976 2935 2978 2954
rect 3152 2935 3154 2954
rect 3328 2935 3330 2954
rect 1863 2934 1867 2935
rect 1863 2929 1867 2930
rect 1895 2934 1899 2935
rect 1895 2929 1899 2930
rect 2031 2934 2035 2935
rect 2031 2929 2035 2930
rect 2167 2934 2171 2935
rect 2167 2929 2171 2930
rect 2175 2934 2179 2935
rect 2175 2929 2179 2930
rect 2295 2934 2299 2935
rect 2295 2929 2299 2930
rect 2423 2934 2427 2935
rect 2423 2929 2427 2930
rect 2495 2934 2499 2935
rect 2495 2929 2499 2930
rect 2543 2934 2547 2935
rect 2543 2929 2547 2930
rect 2671 2934 2675 2935
rect 2671 2929 2675 2930
rect 2815 2934 2819 2935
rect 2815 2929 2819 2930
rect 2823 2934 2827 2935
rect 2823 2929 2827 2930
rect 2975 2934 2979 2935
rect 2975 2929 2979 2930
rect 3151 2934 3155 2935
rect 3151 2929 3155 2930
rect 3167 2934 3171 2935
rect 3167 2929 3171 2930
rect 3327 2934 3331 2935
rect 3327 2929 3331 2930
rect 1822 2924 1828 2925
rect 1822 2920 1823 2924
rect 1827 2920 1828 2924
rect 1822 2919 1828 2920
rect 1734 2911 1740 2912
rect 1734 2907 1735 2911
rect 1739 2907 1740 2911
rect 1734 2906 1740 2907
rect 1690 2899 1696 2900
rect 1690 2895 1691 2899
rect 1695 2895 1696 2899
rect 1690 2894 1696 2895
rect 1736 2891 1738 2906
rect 1824 2891 1826 2919
rect 1864 2905 1866 2929
rect 1896 2918 1898 2929
rect 2176 2918 2178 2929
rect 2318 2927 2324 2928
rect 2318 2923 2319 2927
rect 2323 2923 2324 2927
rect 2318 2922 2324 2923
rect 1894 2917 1900 2918
rect 1894 2913 1895 2917
rect 1899 2913 1900 2917
rect 1894 2912 1900 2913
rect 2174 2917 2180 2918
rect 2174 2913 2175 2917
rect 2179 2913 2180 2917
rect 2174 2912 2180 2913
rect 1862 2904 1868 2905
rect 1862 2900 1863 2904
rect 1867 2900 1868 2904
rect 2320 2900 2322 2922
rect 2496 2918 2498 2929
rect 2562 2927 2568 2928
rect 2562 2923 2563 2927
rect 2567 2923 2568 2927
rect 2562 2922 2568 2923
rect 2494 2917 2500 2918
rect 2494 2913 2495 2917
rect 2499 2913 2500 2917
rect 2494 2912 2500 2913
rect 2564 2900 2566 2922
rect 2824 2918 2826 2929
rect 3168 2918 3170 2929
rect 3472 2928 3474 2970
rect 3574 2968 3575 2972
rect 3579 2968 3580 2972
rect 3574 2967 3580 2968
rect 3486 2959 3492 2960
rect 3486 2955 3487 2959
rect 3491 2955 3492 2959
rect 3486 2954 3492 2955
rect 3488 2935 3490 2954
rect 3576 2935 3578 2967
rect 3487 2934 3491 2935
rect 3487 2929 3491 2930
rect 3575 2934 3579 2935
rect 3575 2929 3579 2930
rect 3470 2927 3476 2928
rect 3470 2923 3471 2927
rect 3475 2923 3476 2927
rect 3470 2922 3476 2923
rect 3488 2918 3490 2929
rect 2822 2917 2828 2918
rect 2822 2913 2823 2917
rect 2827 2913 2828 2917
rect 2822 2912 2828 2913
rect 3166 2917 3172 2918
rect 3166 2913 3167 2917
rect 3171 2913 3172 2917
rect 3166 2912 3172 2913
rect 3486 2917 3492 2918
rect 3486 2913 3487 2917
rect 3491 2913 3492 2917
rect 3486 2912 3492 2913
rect 3576 2905 3578 2929
rect 3574 2904 3580 2905
rect 3574 2900 3575 2904
rect 3579 2900 3580 2904
rect 1862 2899 1868 2900
rect 2318 2899 2324 2900
rect 2318 2895 2319 2899
rect 2323 2895 2324 2899
rect 2318 2894 2324 2895
rect 2562 2899 2568 2900
rect 3574 2899 3580 2900
rect 2562 2895 2563 2899
rect 2567 2895 2568 2899
rect 2562 2894 2568 2895
rect 1191 2890 1195 2891
rect 1191 2885 1195 2886
rect 1279 2890 1283 2891
rect 1279 2885 1283 2886
rect 1311 2890 1315 2891
rect 1311 2885 1315 2886
rect 1415 2890 1419 2891
rect 1415 2885 1419 2886
rect 1423 2890 1427 2891
rect 1423 2885 1427 2886
rect 1535 2890 1539 2891
rect 1535 2885 1539 2886
rect 1551 2890 1555 2891
rect 1551 2885 1555 2886
rect 1647 2890 1651 2891
rect 1647 2885 1651 2886
rect 1735 2890 1739 2891
rect 1735 2885 1739 2886
rect 1823 2890 1827 2891
rect 1823 2885 1827 2886
rect 1862 2887 1868 2888
rect 1280 2874 1282 2885
rect 1416 2874 1418 2885
rect 1502 2883 1508 2884
rect 1502 2879 1503 2883
rect 1507 2879 1508 2883
rect 1502 2878 1508 2879
rect 1278 2873 1284 2874
rect 1278 2869 1279 2873
rect 1283 2869 1284 2873
rect 1142 2868 1148 2869
rect 1167 2868 1171 2869
rect 1278 2868 1284 2869
rect 1414 2873 1420 2874
rect 1414 2869 1415 2873
rect 1419 2869 1420 2873
rect 1414 2868 1420 2869
rect 1167 2863 1171 2864
rect 1504 2860 1506 2878
rect 1552 2874 1554 2885
rect 1550 2873 1556 2874
rect 1550 2869 1551 2873
rect 1555 2869 1556 2873
rect 1511 2868 1515 2869
rect 1550 2868 1556 2869
rect 1511 2863 1515 2864
rect 1502 2859 1508 2860
rect 1502 2855 1503 2859
rect 1507 2855 1508 2859
rect 1512 2856 1514 2863
rect 1824 2861 1826 2885
rect 1862 2883 1863 2887
rect 1867 2883 1868 2887
rect 1862 2882 1868 2883
rect 3070 2887 3076 2888
rect 3070 2883 3071 2887
rect 3075 2883 3076 2887
rect 3070 2882 3076 2883
rect 3574 2887 3580 2888
rect 3574 2883 3575 2887
rect 3579 2883 3580 2887
rect 3574 2882 3580 2883
rect 1864 2867 1866 2882
rect 1886 2877 1892 2878
rect 1886 2873 1887 2877
rect 1891 2873 1892 2877
rect 1886 2872 1892 2873
rect 2166 2877 2172 2878
rect 2166 2873 2167 2877
rect 2171 2873 2172 2877
rect 2166 2872 2172 2873
rect 2486 2877 2492 2878
rect 2486 2873 2487 2877
rect 2491 2873 2492 2877
rect 2486 2872 2492 2873
rect 2814 2877 2820 2878
rect 2814 2873 2815 2877
rect 2819 2873 2820 2877
rect 2814 2872 2820 2873
rect 1888 2867 1890 2872
rect 2168 2867 2170 2872
rect 2488 2867 2490 2872
rect 2816 2867 2818 2872
rect 1863 2866 1867 2867
rect 1863 2861 1867 2862
rect 1887 2866 1891 2867
rect 1887 2861 1891 2862
rect 2023 2866 2027 2867
rect 2023 2861 2027 2862
rect 2167 2866 2171 2867
rect 2167 2861 2171 2862
rect 2191 2866 2195 2867
rect 2191 2861 2195 2862
rect 2359 2866 2363 2867
rect 2359 2861 2363 2862
rect 2487 2866 2491 2867
rect 2487 2861 2491 2862
rect 2519 2866 2523 2867
rect 2519 2861 2523 2862
rect 2671 2866 2675 2867
rect 2807 2866 2811 2867
rect 2671 2861 2675 2862
rect 2686 2863 2692 2864
rect 1822 2860 1828 2861
rect 1822 2856 1823 2860
rect 1827 2856 1828 2860
rect 1502 2854 1508 2855
rect 1510 2855 1516 2856
rect 1822 2855 1828 2856
rect 1510 2851 1511 2855
rect 1515 2851 1516 2855
rect 1510 2850 1516 2851
rect 1864 2846 1866 2861
rect 1888 2856 1890 2861
rect 2024 2856 2026 2861
rect 2192 2856 2194 2861
rect 2360 2856 2362 2861
rect 2520 2856 2522 2861
rect 2672 2856 2674 2861
rect 2686 2859 2687 2863
rect 2691 2859 2692 2863
rect 2807 2861 2811 2862
rect 2815 2866 2819 2867
rect 2815 2861 2819 2862
rect 2935 2866 2939 2867
rect 2935 2861 2939 2862
rect 3055 2866 3059 2867
rect 3055 2861 3059 2862
rect 2686 2858 2692 2859
rect 1886 2855 1892 2856
rect 1886 2851 1887 2855
rect 1891 2851 1892 2855
rect 1886 2850 1892 2851
rect 2022 2855 2028 2856
rect 2022 2851 2023 2855
rect 2027 2851 2028 2855
rect 2022 2850 2028 2851
rect 2190 2855 2196 2856
rect 2190 2851 2191 2855
rect 2195 2851 2196 2855
rect 2190 2850 2196 2851
rect 2358 2855 2364 2856
rect 2358 2851 2359 2855
rect 2363 2851 2364 2855
rect 2358 2850 2364 2851
rect 2518 2855 2524 2856
rect 2518 2851 2519 2855
rect 2523 2851 2524 2855
rect 2518 2850 2524 2851
rect 2670 2855 2676 2856
rect 2670 2851 2671 2855
rect 2675 2851 2676 2855
rect 2670 2850 2676 2851
rect 1862 2845 1868 2846
rect 1822 2843 1828 2844
rect 1822 2839 1823 2843
rect 1827 2839 1828 2843
rect 1862 2841 1863 2845
rect 1867 2841 1868 2845
rect 1862 2840 1868 2841
rect 1822 2838 1828 2839
rect 1134 2833 1140 2834
rect 1134 2829 1135 2833
rect 1139 2829 1140 2833
rect 1134 2828 1140 2829
rect 1270 2833 1276 2834
rect 1270 2829 1271 2833
rect 1275 2829 1276 2833
rect 1270 2828 1276 2829
rect 1406 2833 1412 2834
rect 1406 2829 1407 2833
rect 1411 2829 1412 2833
rect 1406 2828 1412 2829
rect 1542 2833 1548 2834
rect 1542 2829 1543 2833
rect 1547 2829 1548 2833
rect 1542 2828 1548 2829
rect 1136 2815 1138 2828
rect 1272 2815 1274 2828
rect 1408 2815 1410 2828
rect 1544 2815 1546 2828
rect 1824 2815 1826 2838
rect 2090 2831 2096 2832
rect 1862 2828 1868 2829
rect 1862 2824 1863 2828
rect 1867 2824 1868 2828
rect 2090 2827 2091 2831
rect 2095 2827 2096 2831
rect 2090 2826 2096 2827
rect 1862 2823 1868 2824
rect 1079 2814 1083 2815
rect 999 2809 1003 2810
rect 1014 2811 1020 2812
rect 112 2794 114 2809
rect 168 2804 170 2809
rect 296 2804 298 2809
rect 424 2804 426 2809
rect 560 2804 562 2809
rect 696 2804 698 2809
rect 824 2804 826 2809
rect 952 2804 954 2809
rect 1014 2807 1015 2811
rect 1019 2807 1020 2811
rect 1079 2809 1083 2810
rect 1135 2814 1139 2815
rect 1135 2809 1139 2810
rect 1207 2814 1211 2815
rect 1207 2809 1211 2810
rect 1271 2814 1275 2815
rect 1271 2809 1275 2810
rect 1343 2814 1347 2815
rect 1343 2809 1347 2810
rect 1407 2814 1411 2815
rect 1407 2809 1411 2810
rect 1543 2814 1547 2815
rect 1543 2809 1547 2810
rect 1823 2814 1827 2815
rect 1823 2809 1827 2810
rect 1014 2806 1020 2807
rect 1080 2804 1082 2809
rect 1208 2804 1210 2809
rect 1344 2804 1346 2809
rect 166 2803 172 2804
rect 166 2799 167 2803
rect 171 2799 172 2803
rect 166 2798 172 2799
rect 294 2803 300 2804
rect 294 2799 295 2803
rect 299 2799 300 2803
rect 294 2798 300 2799
rect 422 2803 428 2804
rect 422 2799 423 2803
rect 427 2799 428 2803
rect 422 2798 428 2799
rect 558 2803 564 2804
rect 558 2799 559 2803
rect 563 2799 564 2803
rect 558 2798 564 2799
rect 694 2803 700 2804
rect 694 2799 695 2803
rect 699 2799 700 2803
rect 694 2798 700 2799
rect 822 2803 828 2804
rect 822 2799 823 2803
rect 827 2799 828 2803
rect 822 2798 828 2799
rect 950 2803 956 2804
rect 950 2799 951 2803
rect 955 2799 956 2803
rect 950 2798 956 2799
rect 1078 2803 1084 2804
rect 1078 2799 1079 2803
rect 1083 2799 1084 2803
rect 1078 2798 1084 2799
rect 1206 2803 1212 2804
rect 1206 2799 1207 2803
rect 1211 2799 1212 2803
rect 1206 2798 1212 2799
rect 1342 2803 1348 2804
rect 1342 2799 1343 2803
rect 1347 2799 1348 2803
rect 1342 2798 1348 2799
rect 1824 2794 1826 2809
rect 1864 2799 1866 2823
rect 1894 2815 1900 2816
rect 1894 2811 1895 2815
rect 1899 2811 1900 2815
rect 1894 2810 1900 2811
rect 2030 2815 2036 2816
rect 2030 2811 2031 2815
rect 2035 2811 2036 2815
rect 2030 2810 2036 2811
rect 1896 2799 1898 2810
rect 2032 2799 2034 2810
rect 1863 2798 1867 2799
rect 110 2793 116 2794
rect 110 2789 111 2793
rect 115 2789 116 2793
rect 110 2788 116 2789
rect 1822 2793 1828 2794
rect 1863 2793 1867 2794
rect 1895 2798 1899 2799
rect 1895 2793 1899 2794
rect 2031 2798 2035 2799
rect 2031 2793 2035 2794
rect 2063 2798 2067 2799
rect 2063 2793 2067 2794
rect 1822 2789 1823 2793
rect 1827 2789 1828 2793
rect 1822 2788 1828 2789
rect 362 2779 368 2780
rect 110 2776 116 2777
rect 110 2772 111 2776
rect 115 2772 116 2776
rect 362 2775 363 2779
rect 367 2775 368 2779
rect 362 2774 368 2775
rect 626 2779 632 2780
rect 626 2775 627 2779
rect 631 2775 632 2779
rect 626 2774 632 2775
rect 646 2779 652 2780
rect 646 2775 647 2779
rect 651 2775 652 2779
rect 646 2774 652 2775
rect 1822 2776 1828 2777
rect 110 2771 116 2772
rect 112 2739 114 2771
rect 174 2763 180 2764
rect 174 2759 175 2763
rect 179 2759 180 2763
rect 174 2758 180 2759
rect 302 2763 308 2764
rect 302 2759 303 2763
rect 307 2759 308 2763
rect 302 2758 308 2759
rect 176 2739 178 2758
rect 183 2756 187 2757
rect 182 2751 188 2752
rect 182 2747 183 2751
rect 187 2747 188 2751
rect 182 2746 188 2747
rect 304 2739 306 2758
rect 111 2738 115 2739
rect 111 2733 115 2734
rect 143 2738 147 2739
rect 143 2733 147 2734
rect 175 2738 179 2739
rect 175 2733 179 2734
rect 231 2738 235 2739
rect 231 2733 235 2734
rect 303 2738 307 2739
rect 303 2733 307 2734
rect 351 2738 355 2739
rect 351 2733 355 2734
rect 112 2709 114 2733
rect 144 2722 146 2733
rect 210 2731 216 2732
rect 210 2727 211 2731
rect 215 2727 216 2731
rect 210 2726 216 2727
rect 142 2721 148 2722
rect 142 2717 143 2721
rect 147 2717 148 2721
rect 142 2716 148 2717
rect 110 2708 116 2709
rect 110 2704 111 2708
rect 115 2704 116 2708
rect 212 2704 214 2726
rect 232 2722 234 2733
rect 352 2722 354 2733
rect 364 2732 366 2774
rect 430 2763 436 2764
rect 430 2759 431 2763
rect 435 2759 436 2763
rect 430 2758 436 2759
rect 566 2763 572 2764
rect 566 2759 567 2763
rect 571 2759 572 2763
rect 566 2758 572 2759
rect 432 2739 434 2758
rect 568 2739 570 2758
rect 628 2752 630 2774
rect 648 2757 650 2774
rect 1822 2772 1823 2776
rect 1827 2772 1828 2776
rect 1822 2771 1828 2772
rect 702 2763 708 2764
rect 702 2759 703 2763
rect 707 2759 708 2763
rect 702 2758 708 2759
rect 830 2763 836 2764
rect 830 2759 831 2763
rect 835 2759 836 2763
rect 830 2758 836 2759
rect 958 2763 964 2764
rect 958 2759 959 2763
rect 963 2759 964 2763
rect 958 2758 964 2759
rect 1086 2763 1092 2764
rect 1086 2759 1087 2763
rect 1091 2759 1092 2763
rect 1086 2758 1092 2759
rect 1214 2763 1220 2764
rect 1214 2759 1215 2763
rect 1219 2759 1220 2763
rect 1214 2758 1220 2759
rect 1350 2763 1356 2764
rect 1350 2759 1351 2763
rect 1355 2759 1356 2763
rect 1350 2758 1356 2759
rect 647 2756 651 2757
rect 626 2751 632 2752
rect 647 2751 651 2752
rect 626 2747 627 2751
rect 631 2747 632 2751
rect 626 2746 632 2747
rect 704 2739 706 2758
rect 832 2739 834 2758
rect 960 2739 962 2758
rect 1088 2739 1090 2758
rect 1216 2739 1218 2758
rect 1352 2739 1354 2758
rect 1824 2739 1826 2771
rect 1864 2769 1866 2793
rect 1896 2782 1898 2793
rect 2064 2782 2066 2793
rect 2092 2792 2094 2826
rect 2198 2815 2204 2816
rect 2198 2811 2199 2815
rect 2203 2811 2204 2815
rect 2198 2810 2204 2811
rect 2366 2815 2372 2816
rect 2366 2811 2367 2815
rect 2371 2811 2372 2815
rect 2366 2810 2372 2811
rect 2526 2815 2532 2816
rect 2526 2811 2527 2815
rect 2531 2811 2532 2815
rect 2526 2810 2532 2811
rect 2678 2815 2684 2816
rect 2678 2811 2679 2815
rect 2683 2811 2684 2815
rect 2678 2810 2684 2811
rect 2200 2799 2202 2810
rect 2368 2799 2370 2810
rect 2528 2799 2530 2810
rect 2680 2799 2682 2810
rect 2688 2804 2690 2858
rect 2808 2856 2810 2861
rect 2936 2856 2938 2861
rect 3056 2856 3058 2861
rect 2806 2855 2812 2856
rect 2806 2851 2807 2855
rect 2811 2851 2812 2855
rect 2806 2850 2812 2851
rect 2934 2855 2940 2856
rect 2934 2851 2935 2855
rect 2939 2851 2940 2855
rect 2934 2850 2940 2851
rect 3054 2855 3060 2856
rect 3054 2851 3055 2855
rect 3059 2851 3060 2855
rect 3054 2850 3060 2851
rect 2814 2815 2820 2816
rect 2814 2811 2815 2815
rect 2819 2811 2820 2815
rect 2814 2810 2820 2811
rect 2942 2815 2948 2816
rect 2942 2811 2943 2815
rect 2947 2811 2948 2815
rect 2942 2810 2948 2811
rect 3062 2815 3068 2816
rect 3062 2811 3063 2815
rect 3067 2811 3068 2815
rect 3062 2810 3068 2811
rect 2686 2803 2692 2804
rect 2686 2799 2687 2803
rect 2691 2799 2692 2803
rect 2816 2799 2818 2810
rect 2944 2799 2946 2810
rect 3064 2799 3066 2810
rect 3072 2804 3074 2882
rect 3158 2877 3164 2878
rect 3158 2873 3159 2877
rect 3163 2873 3164 2877
rect 3158 2872 3164 2873
rect 3478 2877 3484 2878
rect 3478 2873 3479 2877
rect 3483 2873 3484 2877
rect 3478 2872 3484 2873
rect 3160 2867 3162 2872
rect 3480 2867 3482 2872
rect 3576 2867 3578 2882
rect 3159 2866 3163 2867
rect 3159 2861 3163 2862
rect 3167 2866 3171 2867
rect 3167 2861 3171 2862
rect 3279 2866 3283 2867
rect 3279 2861 3283 2862
rect 3391 2866 3395 2867
rect 3391 2861 3395 2862
rect 3479 2866 3483 2867
rect 3479 2861 3483 2862
rect 3575 2866 3579 2867
rect 3575 2861 3579 2862
rect 3168 2856 3170 2861
rect 3280 2856 3282 2861
rect 3392 2856 3394 2861
rect 3480 2856 3482 2861
rect 3166 2855 3172 2856
rect 3166 2851 3167 2855
rect 3171 2851 3172 2855
rect 3166 2850 3172 2851
rect 3278 2855 3284 2856
rect 3278 2851 3279 2855
rect 3283 2851 3284 2855
rect 3278 2850 3284 2851
rect 3390 2855 3396 2856
rect 3390 2851 3391 2855
rect 3395 2851 3396 2855
rect 3390 2850 3396 2851
rect 3478 2855 3484 2856
rect 3478 2851 3479 2855
rect 3483 2851 3484 2855
rect 3478 2850 3484 2851
rect 3576 2846 3578 2861
rect 3574 2845 3580 2846
rect 3574 2841 3575 2845
rect 3579 2841 3580 2845
rect 3574 2840 3580 2841
rect 3234 2831 3240 2832
rect 3234 2827 3235 2831
rect 3239 2827 3240 2831
rect 3234 2826 3240 2827
rect 3346 2831 3352 2832
rect 3346 2827 3347 2831
rect 3351 2827 3352 2831
rect 3346 2826 3352 2827
rect 3470 2831 3476 2832
rect 3470 2827 3471 2831
rect 3475 2827 3476 2831
rect 3470 2826 3476 2827
rect 3574 2828 3580 2829
rect 3174 2815 3180 2816
rect 3174 2811 3175 2815
rect 3179 2811 3180 2815
rect 3174 2810 3180 2811
rect 3070 2803 3076 2804
rect 3070 2799 3071 2803
rect 3075 2799 3076 2803
rect 3176 2799 3178 2810
rect 3236 2804 3238 2826
rect 3286 2815 3292 2816
rect 3286 2811 3287 2815
rect 3291 2811 3292 2815
rect 3286 2810 3292 2811
rect 3234 2803 3240 2804
rect 3234 2799 3235 2803
rect 3239 2799 3240 2803
rect 3288 2799 3290 2810
rect 3348 2804 3350 2826
rect 3398 2815 3404 2816
rect 3398 2811 3399 2815
rect 3403 2811 3404 2815
rect 3398 2810 3404 2811
rect 3346 2803 3352 2804
rect 3346 2799 3347 2803
rect 3351 2799 3352 2803
rect 3400 2799 3402 2810
rect 3426 2803 3432 2804
rect 3426 2799 3427 2803
rect 3431 2799 3432 2803
rect 2199 2798 2203 2799
rect 2199 2793 2203 2794
rect 2255 2798 2259 2799
rect 2255 2793 2259 2794
rect 2367 2798 2371 2799
rect 2367 2793 2371 2794
rect 2439 2798 2443 2799
rect 2439 2793 2443 2794
rect 2527 2798 2531 2799
rect 2527 2793 2531 2794
rect 2615 2798 2619 2799
rect 2615 2793 2619 2794
rect 2679 2798 2683 2799
rect 2686 2798 2692 2799
rect 2783 2798 2787 2799
rect 2679 2793 2683 2794
rect 2783 2793 2787 2794
rect 2815 2798 2819 2799
rect 2815 2793 2819 2794
rect 2935 2798 2939 2799
rect 2935 2793 2939 2794
rect 2943 2798 2947 2799
rect 2943 2793 2947 2794
rect 3063 2798 3067 2799
rect 3070 2798 3076 2799
rect 3079 2798 3083 2799
rect 3063 2793 3067 2794
rect 3079 2793 3083 2794
rect 3175 2798 3179 2799
rect 3175 2793 3179 2794
rect 3223 2798 3227 2799
rect 3234 2798 3240 2799
rect 3287 2798 3291 2799
rect 3346 2798 3352 2799
rect 3367 2798 3371 2799
rect 3223 2793 3227 2794
rect 3287 2793 3291 2794
rect 3367 2793 3371 2794
rect 3399 2798 3403 2799
rect 3426 2798 3432 2799
rect 3399 2793 3403 2794
rect 2090 2791 2096 2792
rect 2090 2787 2091 2791
rect 2095 2787 2096 2791
rect 2090 2786 2096 2787
rect 2256 2782 2258 2793
rect 2338 2791 2344 2792
rect 2338 2787 2339 2791
rect 2343 2787 2344 2791
rect 2338 2786 2344 2787
rect 1894 2781 1900 2782
rect 1894 2777 1895 2781
rect 1899 2777 1900 2781
rect 1894 2776 1900 2777
rect 2062 2781 2068 2782
rect 2062 2777 2063 2781
rect 2067 2777 2068 2781
rect 2062 2776 2068 2777
rect 2254 2781 2260 2782
rect 2254 2777 2255 2781
rect 2259 2777 2260 2781
rect 2254 2776 2260 2777
rect 1862 2768 1868 2769
rect 1862 2764 1863 2768
rect 1867 2764 1868 2768
rect 2340 2764 2342 2786
rect 2440 2782 2442 2793
rect 2506 2791 2512 2792
rect 2506 2787 2507 2791
rect 2511 2787 2512 2791
rect 2506 2786 2512 2787
rect 2562 2791 2568 2792
rect 2562 2787 2563 2791
rect 2567 2787 2568 2791
rect 2562 2786 2568 2787
rect 2438 2781 2444 2782
rect 2438 2777 2439 2781
rect 2443 2777 2444 2781
rect 2438 2776 2444 2777
rect 2508 2764 2510 2786
rect 1862 2763 1868 2764
rect 2338 2763 2344 2764
rect 2338 2759 2339 2763
rect 2343 2759 2344 2763
rect 2338 2758 2344 2759
rect 2506 2763 2512 2764
rect 2506 2759 2507 2763
rect 2511 2759 2512 2763
rect 2506 2758 2512 2759
rect 1862 2751 1868 2752
rect 1862 2747 1863 2751
rect 1867 2747 1868 2751
rect 1862 2746 1868 2747
rect 431 2738 435 2739
rect 431 2733 435 2734
rect 479 2738 483 2739
rect 479 2733 483 2734
rect 567 2738 571 2739
rect 567 2733 571 2734
rect 615 2738 619 2739
rect 615 2733 619 2734
rect 703 2738 707 2739
rect 703 2733 707 2734
rect 759 2738 763 2739
rect 759 2733 763 2734
rect 831 2738 835 2739
rect 831 2733 835 2734
rect 903 2738 907 2739
rect 903 2733 907 2734
rect 959 2738 963 2739
rect 959 2733 963 2734
rect 1047 2738 1051 2739
rect 1047 2733 1051 2734
rect 1087 2738 1091 2739
rect 1087 2733 1091 2734
rect 1215 2738 1219 2739
rect 1215 2733 1219 2734
rect 1351 2738 1355 2739
rect 1351 2733 1355 2734
rect 1823 2738 1827 2739
rect 1823 2733 1827 2734
rect 362 2731 368 2732
rect 362 2727 363 2731
rect 367 2727 368 2731
rect 362 2726 368 2727
rect 480 2722 482 2733
rect 616 2722 618 2733
rect 760 2722 762 2733
rect 904 2722 906 2733
rect 1048 2722 1050 2733
rect 230 2721 236 2722
rect 230 2717 231 2721
rect 235 2717 236 2721
rect 230 2716 236 2717
rect 350 2721 356 2722
rect 350 2717 351 2721
rect 355 2717 356 2721
rect 350 2716 356 2717
rect 478 2721 484 2722
rect 478 2717 479 2721
rect 483 2717 484 2721
rect 478 2716 484 2717
rect 614 2721 620 2722
rect 614 2717 615 2721
rect 619 2717 620 2721
rect 614 2716 620 2717
rect 758 2721 764 2722
rect 758 2717 759 2721
rect 763 2717 764 2721
rect 758 2716 764 2717
rect 902 2721 908 2722
rect 902 2717 903 2721
rect 907 2717 908 2721
rect 902 2716 908 2717
rect 1046 2721 1052 2722
rect 1046 2717 1047 2721
rect 1051 2717 1052 2721
rect 1046 2716 1052 2717
rect 1824 2709 1826 2733
rect 1864 2727 1866 2746
rect 1886 2741 1892 2742
rect 1886 2737 1887 2741
rect 1891 2737 1892 2741
rect 1886 2736 1892 2737
rect 2054 2741 2060 2742
rect 2054 2737 2055 2741
rect 2059 2737 2060 2741
rect 2054 2736 2060 2737
rect 2246 2741 2252 2742
rect 2246 2737 2247 2741
rect 2251 2737 2252 2741
rect 2246 2736 2252 2737
rect 2430 2741 2436 2742
rect 2430 2737 2431 2741
rect 2435 2737 2436 2741
rect 2430 2736 2436 2737
rect 1888 2727 1890 2736
rect 2056 2727 2058 2736
rect 2248 2727 2250 2736
rect 2432 2727 2434 2736
rect 1863 2726 1867 2727
rect 1863 2721 1867 2722
rect 1887 2726 1891 2727
rect 1887 2721 1891 2722
rect 2047 2726 2051 2727
rect 2047 2721 2051 2722
rect 2055 2726 2059 2727
rect 2055 2721 2059 2722
rect 2207 2726 2211 2727
rect 2207 2721 2211 2722
rect 2247 2726 2251 2727
rect 2247 2721 2251 2722
rect 2359 2726 2363 2727
rect 2359 2721 2363 2722
rect 2431 2726 2435 2727
rect 2431 2721 2435 2722
rect 2495 2726 2499 2727
rect 2495 2721 2499 2722
rect 1822 2708 1828 2709
rect 1822 2704 1823 2708
rect 1827 2704 1828 2708
rect 1864 2706 1866 2721
rect 1888 2716 1890 2721
rect 2048 2716 2050 2721
rect 2208 2716 2210 2721
rect 2360 2716 2362 2721
rect 2496 2716 2498 2721
rect 1886 2715 1892 2716
rect 1886 2711 1887 2715
rect 1891 2711 1892 2715
rect 1886 2710 1892 2711
rect 2046 2715 2052 2716
rect 2046 2711 2047 2715
rect 2051 2711 2052 2715
rect 2046 2710 2052 2711
rect 2206 2715 2212 2716
rect 2206 2711 2207 2715
rect 2211 2711 2212 2715
rect 2206 2710 2212 2711
rect 2358 2715 2364 2716
rect 2358 2711 2359 2715
rect 2363 2711 2364 2715
rect 2358 2710 2364 2711
rect 2494 2715 2500 2716
rect 2494 2711 2495 2715
rect 2499 2711 2500 2715
rect 2494 2710 2500 2711
rect 2564 2708 2566 2786
rect 2616 2782 2618 2793
rect 2784 2782 2786 2793
rect 2846 2791 2852 2792
rect 2846 2787 2847 2791
rect 2851 2787 2852 2791
rect 2846 2786 2852 2787
rect 2614 2781 2620 2782
rect 2614 2777 2615 2781
rect 2619 2777 2620 2781
rect 2614 2776 2620 2777
rect 2782 2781 2788 2782
rect 2782 2777 2783 2781
rect 2787 2777 2788 2781
rect 2782 2776 2788 2777
rect 2606 2741 2612 2742
rect 2606 2737 2607 2741
rect 2611 2737 2612 2741
rect 2606 2736 2612 2737
rect 2774 2741 2780 2742
rect 2774 2737 2775 2741
rect 2779 2737 2780 2741
rect 2774 2736 2780 2737
rect 2608 2727 2610 2736
rect 2776 2727 2778 2736
rect 2848 2728 2850 2786
rect 2936 2782 2938 2793
rect 3080 2782 3082 2793
rect 3224 2782 3226 2793
rect 3368 2782 3370 2793
rect 2934 2781 2940 2782
rect 2934 2777 2935 2781
rect 2939 2777 2940 2781
rect 2934 2776 2940 2777
rect 3078 2781 3084 2782
rect 3078 2777 3079 2781
rect 3083 2777 3084 2781
rect 3078 2776 3084 2777
rect 3222 2781 3228 2782
rect 3222 2777 3223 2781
rect 3227 2777 3228 2781
rect 3222 2776 3228 2777
rect 3366 2781 3372 2782
rect 3366 2777 3367 2781
rect 3371 2777 3372 2781
rect 3366 2776 3372 2777
rect 3428 2768 3430 2798
rect 3472 2792 3474 2826
rect 3574 2824 3575 2828
rect 3579 2824 3580 2828
rect 3574 2823 3580 2824
rect 3486 2815 3492 2816
rect 3486 2811 3487 2815
rect 3491 2811 3492 2815
rect 3486 2810 3492 2811
rect 3488 2799 3490 2810
rect 3576 2799 3578 2823
rect 3487 2798 3491 2799
rect 3487 2793 3491 2794
rect 3575 2798 3579 2799
rect 3575 2793 3579 2794
rect 3434 2791 3440 2792
rect 3434 2787 3435 2791
rect 3439 2787 3440 2791
rect 3434 2786 3440 2787
rect 3470 2791 3476 2792
rect 3470 2787 3471 2791
rect 3475 2787 3476 2791
rect 3470 2786 3476 2787
rect 3426 2767 3432 2768
rect 3426 2763 3427 2767
rect 3431 2763 3432 2767
rect 3436 2764 3438 2786
rect 3488 2782 3490 2793
rect 3486 2781 3492 2782
rect 3486 2777 3487 2781
rect 3491 2777 3492 2781
rect 3486 2776 3492 2777
rect 3576 2769 3578 2793
rect 3574 2768 3580 2769
rect 3574 2764 3575 2768
rect 3579 2764 3580 2768
rect 3426 2762 3432 2763
rect 3434 2763 3440 2764
rect 3574 2763 3580 2764
rect 3434 2759 3435 2763
rect 3439 2759 3440 2763
rect 3434 2758 3440 2759
rect 3574 2751 3580 2752
rect 3574 2747 3575 2751
rect 3579 2747 3580 2751
rect 3574 2746 3580 2747
rect 2926 2741 2932 2742
rect 2926 2737 2927 2741
rect 2931 2737 2932 2741
rect 2926 2736 2932 2737
rect 3070 2741 3076 2742
rect 3070 2737 3071 2741
rect 3075 2737 3076 2741
rect 3070 2736 3076 2737
rect 3214 2741 3220 2742
rect 3214 2737 3215 2741
rect 3219 2737 3220 2741
rect 3214 2736 3220 2737
rect 3358 2741 3364 2742
rect 3358 2737 3359 2741
rect 3363 2737 3364 2741
rect 3358 2736 3364 2737
rect 3478 2741 3484 2742
rect 3478 2737 3479 2741
rect 3483 2737 3484 2741
rect 3478 2736 3484 2737
rect 2846 2727 2852 2728
rect 2928 2727 2930 2736
rect 2974 2735 2980 2736
rect 2974 2731 2975 2735
rect 2979 2731 2980 2735
rect 2974 2730 2980 2731
rect 2607 2726 2611 2727
rect 2607 2721 2611 2722
rect 2623 2726 2627 2727
rect 2623 2721 2627 2722
rect 2743 2726 2747 2727
rect 2743 2721 2747 2722
rect 2775 2726 2779 2727
rect 2846 2723 2847 2727
rect 2851 2723 2852 2727
rect 2846 2722 2852 2723
rect 2863 2726 2867 2727
rect 2775 2721 2779 2722
rect 2863 2721 2867 2722
rect 2927 2726 2931 2727
rect 2927 2721 2931 2722
rect 2624 2716 2626 2721
rect 2744 2716 2746 2721
rect 2864 2716 2866 2721
rect 2622 2715 2628 2716
rect 2622 2711 2623 2715
rect 2627 2711 2628 2715
rect 2622 2710 2628 2711
rect 2742 2715 2748 2716
rect 2742 2711 2743 2715
rect 2747 2711 2748 2715
rect 2742 2710 2748 2711
rect 2862 2715 2868 2716
rect 2862 2711 2863 2715
rect 2867 2711 2868 2715
rect 2862 2710 2868 2711
rect 2562 2707 2568 2708
rect 110 2703 116 2704
rect 210 2703 216 2704
rect 1822 2703 1828 2704
rect 1862 2705 1868 2706
rect 210 2699 211 2703
rect 215 2699 216 2703
rect 1862 2701 1863 2705
rect 1867 2701 1868 2705
rect 2562 2703 2563 2707
rect 2567 2703 2568 2707
rect 2562 2702 2568 2703
rect 1862 2700 1868 2701
rect 210 2698 216 2699
rect 110 2691 116 2692
rect 110 2687 111 2691
rect 115 2687 116 2691
rect 110 2686 116 2687
rect 1822 2691 1828 2692
rect 1822 2687 1823 2691
rect 1827 2687 1828 2691
rect 1954 2691 1960 2692
rect 1822 2686 1828 2687
rect 1862 2688 1868 2689
rect 112 2667 114 2686
rect 134 2681 140 2682
rect 134 2677 135 2681
rect 139 2677 140 2681
rect 134 2676 140 2677
rect 222 2681 228 2682
rect 222 2677 223 2681
rect 227 2677 228 2681
rect 222 2676 228 2677
rect 342 2681 348 2682
rect 342 2677 343 2681
rect 347 2677 348 2681
rect 342 2676 348 2677
rect 470 2681 476 2682
rect 470 2677 471 2681
rect 475 2677 476 2681
rect 470 2676 476 2677
rect 606 2681 612 2682
rect 606 2677 607 2681
rect 611 2677 612 2681
rect 606 2676 612 2677
rect 750 2681 756 2682
rect 750 2677 751 2681
rect 755 2677 756 2681
rect 750 2676 756 2677
rect 894 2681 900 2682
rect 894 2677 895 2681
rect 899 2677 900 2681
rect 894 2676 900 2677
rect 1038 2681 1044 2682
rect 1038 2677 1039 2681
rect 1043 2677 1044 2681
rect 1038 2676 1044 2677
rect 136 2667 138 2676
rect 224 2667 226 2676
rect 344 2667 346 2676
rect 472 2667 474 2676
rect 608 2667 610 2676
rect 752 2667 754 2676
rect 896 2667 898 2676
rect 1040 2667 1042 2676
rect 1824 2667 1826 2686
rect 1862 2684 1863 2688
rect 1867 2684 1868 2688
rect 1954 2687 1955 2691
rect 1959 2687 1960 2691
rect 1954 2686 1960 2687
rect 2690 2691 2696 2692
rect 2690 2687 2691 2691
rect 2695 2687 2696 2691
rect 2690 2686 2696 2687
rect 2698 2691 2704 2692
rect 2698 2687 2699 2691
rect 2703 2687 2704 2691
rect 2698 2686 2704 2687
rect 2810 2691 2816 2692
rect 2810 2687 2811 2691
rect 2815 2687 2816 2691
rect 2810 2686 2816 2687
rect 1862 2683 1868 2684
rect 111 2666 115 2667
rect 111 2661 115 2662
rect 135 2666 139 2667
rect 135 2661 139 2662
rect 223 2666 227 2667
rect 223 2661 227 2662
rect 231 2666 235 2667
rect 231 2661 235 2662
rect 343 2666 347 2667
rect 343 2661 347 2662
rect 351 2666 355 2667
rect 351 2661 355 2662
rect 471 2666 475 2667
rect 471 2661 475 2662
rect 583 2666 587 2667
rect 583 2661 587 2662
rect 607 2666 611 2667
rect 607 2661 611 2662
rect 695 2666 699 2667
rect 695 2661 699 2662
rect 751 2666 755 2667
rect 751 2661 755 2662
rect 799 2666 803 2667
rect 799 2661 803 2662
rect 895 2666 899 2667
rect 895 2661 899 2662
rect 903 2666 907 2667
rect 903 2661 907 2662
rect 999 2666 1003 2667
rect 999 2661 1003 2662
rect 1039 2666 1043 2667
rect 1039 2661 1043 2662
rect 1103 2666 1107 2667
rect 1103 2661 1107 2662
rect 1207 2666 1211 2667
rect 1207 2661 1211 2662
rect 1311 2666 1315 2667
rect 1311 2661 1315 2662
rect 1823 2666 1827 2667
rect 1823 2661 1827 2662
rect 112 2646 114 2661
rect 136 2656 138 2661
rect 232 2656 234 2661
rect 352 2656 354 2661
rect 472 2656 474 2661
rect 584 2656 586 2661
rect 696 2656 698 2661
rect 800 2656 802 2661
rect 904 2656 906 2661
rect 1000 2656 1002 2661
rect 1104 2656 1106 2661
rect 1208 2656 1210 2661
rect 1312 2656 1314 2661
rect 134 2655 140 2656
rect 134 2651 135 2655
rect 139 2651 140 2655
rect 134 2650 140 2651
rect 230 2655 236 2656
rect 230 2651 231 2655
rect 235 2651 236 2655
rect 230 2650 236 2651
rect 350 2655 356 2656
rect 350 2651 351 2655
rect 355 2651 356 2655
rect 350 2650 356 2651
rect 470 2655 476 2656
rect 470 2651 471 2655
rect 475 2651 476 2655
rect 470 2650 476 2651
rect 582 2655 588 2656
rect 582 2651 583 2655
rect 587 2651 588 2655
rect 582 2650 588 2651
rect 694 2655 700 2656
rect 694 2651 695 2655
rect 699 2651 700 2655
rect 694 2650 700 2651
rect 798 2655 804 2656
rect 798 2651 799 2655
rect 803 2651 804 2655
rect 798 2650 804 2651
rect 902 2655 908 2656
rect 902 2651 903 2655
rect 907 2651 908 2655
rect 902 2650 908 2651
rect 998 2655 1004 2656
rect 998 2651 999 2655
rect 1003 2651 1004 2655
rect 998 2650 1004 2651
rect 1102 2655 1108 2656
rect 1102 2651 1103 2655
rect 1107 2651 1108 2655
rect 1102 2650 1108 2651
rect 1206 2655 1212 2656
rect 1206 2651 1207 2655
rect 1211 2651 1212 2655
rect 1206 2650 1212 2651
rect 1310 2655 1316 2656
rect 1310 2651 1311 2655
rect 1315 2651 1316 2655
rect 1310 2650 1316 2651
rect 422 2647 428 2648
rect 110 2645 116 2646
rect 110 2641 111 2645
rect 115 2641 116 2645
rect 422 2643 423 2647
rect 427 2643 428 2647
rect 422 2642 428 2643
rect 1274 2647 1280 2648
rect 1274 2643 1275 2647
rect 1279 2643 1280 2647
rect 1824 2646 1826 2661
rect 1864 2651 1866 2683
rect 1894 2675 1900 2676
rect 1894 2671 1895 2675
rect 1899 2671 1900 2675
rect 1894 2670 1900 2671
rect 1896 2651 1898 2670
rect 1956 2664 1958 2686
rect 2054 2675 2060 2676
rect 2054 2671 2055 2675
rect 2059 2671 2060 2675
rect 2054 2670 2060 2671
rect 2214 2675 2220 2676
rect 2214 2671 2215 2675
rect 2219 2671 2220 2675
rect 2214 2670 2220 2671
rect 2366 2675 2372 2676
rect 2366 2671 2367 2675
rect 2371 2671 2372 2675
rect 2366 2670 2372 2671
rect 2502 2675 2508 2676
rect 2502 2671 2503 2675
rect 2507 2671 2508 2675
rect 2502 2670 2508 2671
rect 2630 2675 2636 2676
rect 2630 2671 2631 2675
rect 2635 2671 2636 2675
rect 2630 2670 2636 2671
rect 1954 2663 1960 2664
rect 1954 2659 1955 2663
rect 1959 2659 1960 2663
rect 1954 2658 1960 2659
rect 2056 2651 2058 2670
rect 2216 2651 2218 2670
rect 2326 2663 2332 2664
rect 2326 2659 2327 2663
rect 2331 2659 2332 2663
rect 2326 2658 2332 2659
rect 1863 2650 1867 2651
rect 1274 2642 1280 2643
rect 1822 2645 1828 2646
rect 1863 2645 1867 2646
rect 1895 2650 1899 2651
rect 1895 2645 1899 2646
rect 1999 2650 2003 2651
rect 1999 2645 2003 2646
rect 2055 2650 2059 2651
rect 2055 2645 2059 2646
rect 2119 2650 2123 2651
rect 2119 2645 2123 2646
rect 2215 2650 2219 2651
rect 2215 2645 2219 2646
rect 2239 2650 2243 2651
rect 2239 2645 2243 2646
rect 110 2640 116 2641
rect 110 2628 116 2629
rect 110 2624 111 2628
rect 115 2624 116 2628
rect 110 2623 116 2624
rect 112 2595 114 2623
rect 142 2615 148 2616
rect 142 2611 143 2615
rect 147 2611 148 2615
rect 142 2610 148 2611
rect 238 2615 244 2616
rect 238 2611 239 2615
rect 243 2611 244 2615
rect 238 2610 244 2611
rect 358 2615 364 2616
rect 358 2611 359 2615
rect 363 2611 364 2615
rect 358 2610 364 2611
rect 144 2595 146 2610
rect 240 2595 242 2610
rect 360 2595 362 2610
rect 111 2594 115 2595
rect 111 2589 115 2590
rect 143 2594 147 2595
rect 143 2589 147 2590
rect 239 2594 243 2595
rect 239 2589 243 2590
rect 271 2594 275 2595
rect 271 2589 275 2590
rect 359 2594 363 2595
rect 359 2589 363 2590
rect 415 2594 419 2595
rect 415 2589 419 2590
rect 112 2565 114 2589
rect 144 2578 146 2589
rect 210 2587 216 2588
rect 210 2583 211 2587
rect 215 2583 216 2587
rect 210 2582 216 2583
rect 142 2577 148 2578
rect 142 2573 143 2577
rect 147 2573 148 2577
rect 142 2572 148 2573
rect 110 2564 116 2565
rect 110 2560 111 2564
rect 115 2560 116 2564
rect 212 2560 214 2582
rect 272 2578 274 2589
rect 338 2587 344 2588
rect 338 2583 339 2587
rect 343 2583 344 2587
rect 338 2582 344 2583
rect 270 2577 276 2578
rect 270 2573 271 2577
rect 275 2573 276 2577
rect 270 2572 276 2573
rect 340 2560 342 2582
rect 416 2578 418 2589
rect 424 2588 426 2642
rect 478 2615 484 2616
rect 478 2611 479 2615
rect 483 2611 484 2615
rect 478 2610 484 2611
rect 590 2615 596 2616
rect 590 2611 591 2615
rect 595 2611 596 2615
rect 590 2610 596 2611
rect 702 2615 708 2616
rect 702 2611 703 2615
rect 707 2611 708 2615
rect 702 2610 708 2611
rect 806 2615 812 2616
rect 806 2611 807 2615
rect 811 2611 812 2615
rect 806 2610 812 2611
rect 910 2615 916 2616
rect 910 2611 911 2615
rect 915 2611 916 2615
rect 910 2610 916 2611
rect 1006 2615 1012 2616
rect 1006 2611 1007 2615
rect 1011 2611 1012 2615
rect 1006 2610 1012 2611
rect 1110 2615 1116 2616
rect 1110 2611 1111 2615
rect 1115 2611 1116 2615
rect 1110 2610 1116 2611
rect 1214 2615 1220 2616
rect 1214 2611 1215 2615
rect 1219 2611 1220 2615
rect 1214 2610 1220 2611
rect 480 2595 482 2610
rect 592 2595 594 2610
rect 618 2603 624 2604
rect 618 2599 619 2603
rect 623 2599 624 2603
rect 618 2598 624 2599
rect 479 2594 483 2595
rect 479 2589 483 2590
rect 551 2594 555 2595
rect 551 2589 555 2590
rect 591 2594 595 2595
rect 591 2589 595 2590
rect 422 2587 428 2588
rect 422 2583 423 2587
rect 427 2583 428 2587
rect 422 2582 428 2583
rect 552 2578 554 2589
rect 414 2577 420 2578
rect 414 2573 415 2577
rect 419 2573 420 2577
rect 414 2572 420 2573
rect 550 2577 556 2578
rect 550 2573 551 2577
rect 555 2573 556 2577
rect 550 2572 556 2573
rect 620 2564 622 2598
rect 704 2595 706 2610
rect 746 2603 752 2604
rect 746 2599 747 2603
rect 751 2599 752 2603
rect 746 2598 752 2599
rect 679 2594 683 2595
rect 679 2589 683 2590
rect 703 2594 707 2595
rect 703 2589 707 2590
rect 650 2587 656 2588
rect 650 2583 651 2587
rect 655 2583 656 2587
rect 650 2582 656 2583
rect 662 2587 668 2588
rect 662 2583 663 2587
rect 667 2583 668 2587
rect 662 2582 668 2583
rect 618 2563 624 2564
rect 110 2559 116 2560
rect 210 2559 216 2560
rect 210 2555 211 2559
rect 215 2555 216 2559
rect 210 2554 216 2555
rect 338 2559 344 2560
rect 338 2555 339 2559
rect 343 2555 344 2559
rect 618 2559 619 2563
rect 623 2559 624 2563
rect 652 2560 654 2582
rect 618 2558 624 2559
rect 650 2559 656 2560
rect 338 2554 344 2555
rect 650 2555 651 2559
rect 655 2555 656 2559
rect 650 2554 656 2555
rect 110 2547 116 2548
rect 110 2543 111 2547
rect 115 2543 116 2547
rect 110 2542 116 2543
rect 112 2527 114 2542
rect 134 2537 140 2538
rect 134 2533 135 2537
rect 139 2533 140 2537
rect 134 2532 140 2533
rect 262 2537 268 2538
rect 262 2533 263 2537
rect 267 2533 268 2537
rect 262 2532 268 2533
rect 406 2537 412 2538
rect 406 2533 407 2537
rect 411 2533 412 2537
rect 406 2532 412 2533
rect 542 2537 548 2538
rect 542 2533 543 2537
rect 547 2533 548 2537
rect 542 2532 548 2533
rect 136 2527 138 2532
rect 264 2527 266 2532
rect 408 2527 410 2532
rect 544 2527 546 2532
rect 111 2526 115 2527
rect 111 2521 115 2522
rect 135 2526 139 2527
rect 135 2521 139 2522
rect 263 2526 267 2527
rect 263 2521 267 2522
rect 279 2526 283 2527
rect 279 2521 283 2522
rect 407 2526 411 2527
rect 407 2521 411 2522
rect 439 2526 443 2527
rect 439 2521 443 2522
rect 543 2526 547 2527
rect 543 2521 547 2522
rect 591 2526 595 2527
rect 591 2521 595 2522
rect 112 2506 114 2521
rect 136 2516 138 2521
rect 280 2516 282 2521
rect 440 2516 442 2521
rect 592 2516 594 2521
rect 134 2515 140 2516
rect 134 2511 135 2515
rect 139 2511 140 2515
rect 134 2510 140 2511
rect 278 2515 284 2516
rect 278 2511 279 2515
rect 283 2511 284 2515
rect 278 2510 284 2511
rect 438 2515 444 2516
rect 438 2511 439 2515
rect 443 2511 444 2515
rect 438 2510 444 2511
rect 590 2515 596 2516
rect 590 2511 591 2515
rect 595 2511 596 2515
rect 590 2510 596 2511
rect 664 2508 666 2582
rect 680 2578 682 2589
rect 678 2577 684 2578
rect 678 2573 679 2577
rect 683 2573 684 2577
rect 678 2572 684 2573
rect 748 2560 750 2598
rect 808 2595 810 2610
rect 912 2595 914 2610
rect 1008 2595 1010 2610
rect 1112 2595 1114 2610
rect 1216 2595 1218 2610
rect 807 2594 811 2595
rect 807 2589 811 2590
rect 911 2594 915 2595
rect 911 2589 915 2590
rect 927 2594 931 2595
rect 927 2589 931 2590
rect 1007 2594 1011 2595
rect 1007 2589 1011 2590
rect 1047 2594 1051 2595
rect 1047 2589 1051 2590
rect 1111 2594 1115 2595
rect 1111 2589 1115 2590
rect 1175 2594 1179 2595
rect 1175 2589 1179 2590
rect 1215 2594 1219 2595
rect 1215 2589 1219 2590
rect 808 2578 810 2589
rect 814 2587 820 2588
rect 814 2583 815 2587
rect 819 2583 820 2587
rect 814 2582 820 2583
rect 806 2577 812 2578
rect 806 2573 807 2577
rect 811 2573 812 2577
rect 806 2572 812 2573
rect 746 2559 752 2560
rect 746 2555 747 2559
rect 751 2555 752 2559
rect 746 2554 752 2555
rect 670 2537 676 2538
rect 670 2533 671 2537
rect 675 2533 676 2537
rect 670 2532 676 2533
rect 798 2537 804 2538
rect 798 2533 799 2537
rect 803 2533 804 2537
rect 798 2532 804 2533
rect 672 2527 674 2532
rect 800 2527 802 2532
rect 671 2526 675 2527
rect 671 2521 675 2522
rect 735 2526 739 2527
rect 735 2521 739 2522
rect 799 2526 803 2527
rect 799 2521 803 2522
rect 736 2516 738 2521
rect 734 2515 740 2516
rect 734 2511 735 2515
rect 739 2511 740 2515
rect 734 2510 740 2511
rect 816 2508 818 2582
rect 928 2578 930 2589
rect 994 2587 1000 2588
rect 994 2583 995 2587
rect 999 2583 1000 2587
rect 994 2582 1000 2583
rect 926 2577 932 2578
rect 926 2573 927 2577
rect 931 2573 932 2577
rect 926 2572 932 2573
rect 996 2560 998 2582
rect 1048 2578 1050 2589
rect 1118 2587 1124 2588
rect 1118 2583 1119 2587
rect 1123 2583 1124 2587
rect 1118 2582 1124 2583
rect 1046 2577 1052 2578
rect 1046 2573 1047 2577
rect 1051 2573 1052 2577
rect 1046 2572 1052 2573
rect 1120 2560 1122 2582
rect 1176 2578 1178 2589
rect 1276 2588 1278 2642
rect 1822 2641 1823 2645
rect 1827 2641 1828 2645
rect 1822 2640 1828 2641
rect 1822 2628 1828 2629
rect 1822 2624 1823 2628
rect 1827 2624 1828 2628
rect 1822 2623 1828 2624
rect 1318 2615 1324 2616
rect 1318 2611 1319 2615
rect 1323 2611 1324 2615
rect 1318 2610 1324 2611
rect 1320 2595 1322 2610
rect 1824 2595 1826 2623
rect 1864 2621 1866 2645
rect 1896 2634 1898 2645
rect 2000 2634 2002 2645
rect 2120 2634 2122 2645
rect 2240 2634 2242 2645
rect 2314 2643 2320 2644
rect 2314 2639 2315 2643
rect 2319 2639 2320 2643
rect 2314 2638 2320 2639
rect 1894 2633 1900 2634
rect 1894 2629 1895 2633
rect 1899 2629 1900 2633
rect 1894 2628 1900 2629
rect 1998 2633 2004 2634
rect 1998 2629 1999 2633
rect 2003 2629 2004 2633
rect 1998 2628 2004 2629
rect 2118 2633 2124 2634
rect 2118 2629 2119 2633
rect 2123 2629 2124 2633
rect 2118 2628 2124 2629
rect 2238 2633 2244 2634
rect 2238 2629 2239 2633
rect 2243 2629 2244 2633
rect 2238 2628 2244 2629
rect 1862 2620 1868 2621
rect 2316 2620 2318 2638
rect 1862 2616 1863 2620
rect 1867 2616 1868 2620
rect 1862 2615 1868 2616
rect 2314 2619 2320 2620
rect 2314 2615 2315 2619
rect 2319 2615 2320 2619
rect 2328 2616 2330 2658
rect 2368 2651 2370 2670
rect 2504 2651 2506 2670
rect 2632 2651 2634 2670
rect 2351 2650 2355 2651
rect 2351 2645 2355 2646
rect 2367 2650 2371 2651
rect 2367 2645 2371 2646
rect 2455 2650 2459 2651
rect 2455 2645 2459 2646
rect 2503 2650 2507 2651
rect 2503 2645 2507 2646
rect 2551 2650 2555 2651
rect 2551 2645 2555 2646
rect 2631 2650 2635 2651
rect 2631 2645 2635 2646
rect 2655 2650 2659 2651
rect 2655 2645 2659 2646
rect 2352 2634 2354 2645
rect 2456 2634 2458 2645
rect 2522 2643 2528 2644
rect 2522 2639 2523 2643
rect 2527 2639 2528 2643
rect 2522 2638 2528 2639
rect 2350 2633 2356 2634
rect 2350 2629 2351 2633
rect 2355 2629 2356 2633
rect 2350 2628 2356 2629
rect 2454 2633 2460 2634
rect 2454 2629 2455 2633
rect 2459 2629 2460 2633
rect 2454 2628 2460 2629
rect 2524 2616 2526 2638
rect 2552 2634 2554 2645
rect 2656 2634 2658 2645
rect 2692 2644 2694 2686
rect 2700 2664 2702 2686
rect 2750 2675 2756 2676
rect 2750 2671 2751 2675
rect 2755 2671 2756 2675
rect 2750 2670 2756 2671
rect 2698 2663 2704 2664
rect 2698 2659 2699 2663
rect 2703 2659 2704 2663
rect 2698 2658 2704 2659
rect 2752 2651 2754 2670
rect 2812 2664 2814 2686
rect 2870 2675 2876 2676
rect 2870 2671 2871 2675
rect 2875 2671 2876 2675
rect 2870 2670 2876 2671
rect 2810 2663 2816 2664
rect 2810 2659 2811 2663
rect 2815 2659 2816 2663
rect 2810 2658 2816 2659
rect 2872 2651 2874 2670
rect 2976 2664 2978 2730
rect 3072 2727 3074 2736
rect 3216 2727 3218 2736
rect 3360 2727 3362 2736
rect 3480 2727 3482 2736
rect 3576 2727 3578 2746
rect 2983 2726 2987 2727
rect 2983 2721 2987 2722
rect 3071 2726 3075 2727
rect 3071 2721 3075 2722
rect 3103 2726 3107 2727
rect 3103 2721 3107 2722
rect 3215 2726 3219 2727
rect 3215 2721 3219 2722
rect 3359 2726 3363 2727
rect 3359 2721 3363 2722
rect 3479 2726 3483 2727
rect 3479 2721 3483 2722
rect 3575 2726 3579 2727
rect 3575 2721 3579 2722
rect 2984 2716 2986 2721
rect 3104 2716 3106 2721
rect 2982 2715 2988 2716
rect 2982 2711 2983 2715
rect 2987 2711 2988 2715
rect 2982 2710 2988 2711
rect 3102 2715 3108 2716
rect 3102 2711 3103 2715
rect 3107 2711 3108 2715
rect 3102 2710 3108 2711
rect 3050 2707 3056 2708
rect 3050 2703 3051 2707
rect 3055 2703 3056 2707
rect 3576 2706 3578 2721
rect 3050 2702 3056 2703
rect 3574 2705 3580 2706
rect 2990 2675 2996 2676
rect 2990 2671 2991 2675
rect 2995 2671 2996 2675
rect 2990 2670 2996 2671
rect 2974 2663 2980 2664
rect 2974 2659 2975 2663
rect 2979 2659 2980 2663
rect 2974 2658 2980 2659
rect 2992 2651 2994 2670
rect 3052 2656 3054 2702
rect 3574 2701 3575 2705
rect 3579 2701 3580 2705
rect 3574 2700 3580 2701
rect 3574 2688 3580 2689
rect 3574 2684 3575 2688
rect 3579 2684 3580 2688
rect 3574 2683 3580 2684
rect 3110 2675 3116 2676
rect 3110 2671 3111 2675
rect 3115 2671 3116 2675
rect 3110 2670 3116 2671
rect 3050 2655 3056 2656
rect 3050 2651 3051 2655
rect 3055 2651 3056 2655
rect 3112 2651 3114 2670
rect 3576 2651 3578 2683
rect 2751 2650 2755 2651
rect 2751 2645 2755 2646
rect 2759 2650 2763 2651
rect 2759 2645 2763 2646
rect 2863 2650 2867 2651
rect 2863 2645 2867 2646
rect 2871 2650 2875 2651
rect 2871 2645 2875 2646
rect 2991 2650 2995 2651
rect 3050 2650 3056 2651
rect 3111 2650 3115 2651
rect 2991 2645 2995 2646
rect 3111 2645 3115 2646
rect 3575 2650 3579 2651
rect 3575 2645 3579 2646
rect 2690 2643 2696 2644
rect 2690 2639 2691 2643
rect 2695 2639 2696 2643
rect 2690 2638 2696 2639
rect 2760 2634 2762 2645
rect 2864 2634 2866 2645
rect 2550 2633 2556 2634
rect 2550 2629 2551 2633
rect 2555 2629 2556 2633
rect 2550 2628 2556 2629
rect 2654 2633 2660 2634
rect 2654 2629 2655 2633
rect 2659 2629 2660 2633
rect 2654 2628 2660 2629
rect 2758 2633 2764 2634
rect 2758 2629 2759 2633
rect 2763 2629 2764 2633
rect 2758 2628 2764 2629
rect 2862 2633 2868 2634
rect 2862 2629 2863 2633
rect 2867 2629 2868 2633
rect 2862 2628 2868 2629
rect 3576 2621 3578 2645
rect 3574 2620 3580 2621
rect 3574 2616 3575 2620
rect 3579 2616 3580 2620
rect 2314 2614 2320 2615
rect 2326 2615 2332 2616
rect 2326 2611 2327 2615
rect 2331 2611 2332 2615
rect 2326 2610 2332 2611
rect 2522 2615 2528 2616
rect 3574 2615 3580 2616
rect 2522 2611 2523 2615
rect 2527 2611 2528 2615
rect 2522 2610 2528 2611
rect 1862 2603 1868 2604
rect 1862 2599 1863 2603
rect 1867 2599 1868 2603
rect 1862 2598 1868 2599
rect 3574 2603 3580 2604
rect 3574 2599 3575 2603
rect 3579 2599 3580 2603
rect 3574 2598 3580 2599
rect 1319 2594 1323 2595
rect 1319 2589 1323 2590
rect 1823 2594 1827 2595
rect 1823 2589 1827 2590
rect 1274 2587 1280 2588
rect 1274 2583 1275 2587
rect 1279 2583 1280 2587
rect 1274 2582 1280 2583
rect 1174 2577 1180 2578
rect 1174 2573 1175 2577
rect 1179 2573 1180 2577
rect 1174 2572 1180 2573
rect 1824 2565 1826 2589
rect 1864 2579 1866 2598
rect 1886 2593 1892 2594
rect 1886 2589 1887 2593
rect 1891 2589 1892 2593
rect 1886 2588 1892 2589
rect 1990 2593 1996 2594
rect 1990 2589 1991 2593
rect 1995 2589 1996 2593
rect 1990 2588 1996 2589
rect 2110 2593 2116 2594
rect 2110 2589 2111 2593
rect 2115 2589 2116 2593
rect 2110 2588 2116 2589
rect 2230 2593 2236 2594
rect 2230 2589 2231 2593
rect 2235 2589 2236 2593
rect 2230 2588 2236 2589
rect 2342 2593 2348 2594
rect 2342 2589 2343 2593
rect 2347 2589 2348 2593
rect 2342 2588 2348 2589
rect 2446 2593 2452 2594
rect 2446 2589 2447 2593
rect 2451 2589 2452 2593
rect 2446 2588 2452 2589
rect 2542 2593 2548 2594
rect 2542 2589 2543 2593
rect 2547 2589 2548 2593
rect 2542 2588 2548 2589
rect 2646 2593 2652 2594
rect 2646 2589 2647 2593
rect 2651 2589 2652 2593
rect 2646 2588 2652 2589
rect 2750 2593 2756 2594
rect 2750 2589 2751 2593
rect 2755 2589 2756 2593
rect 2750 2588 2756 2589
rect 2854 2593 2860 2594
rect 2854 2589 2855 2593
rect 2859 2589 2860 2593
rect 2854 2588 2860 2589
rect 1888 2579 1890 2588
rect 1992 2579 1994 2588
rect 2112 2579 2114 2588
rect 2232 2579 2234 2588
rect 2344 2579 2346 2588
rect 2448 2579 2450 2588
rect 2486 2587 2492 2588
rect 2486 2583 2487 2587
rect 2491 2583 2492 2587
rect 2486 2582 2492 2583
rect 1863 2578 1867 2579
rect 1863 2573 1867 2574
rect 1887 2578 1891 2579
rect 1887 2573 1891 2574
rect 1991 2578 1995 2579
rect 1991 2573 1995 2574
rect 2111 2578 2115 2579
rect 2111 2573 2115 2574
rect 2231 2578 2235 2579
rect 2231 2573 2235 2574
rect 2343 2578 2347 2579
rect 2343 2573 2347 2574
rect 2351 2578 2355 2579
rect 2351 2573 2355 2574
rect 2447 2578 2451 2579
rect 2447 2573 2451 2574
rect 2471 2578 2475 2579
rect 2471 2573 2475 2574
rect 1822 2564 1828 2565
rect 1822 2560 1823 2564
rect 1827 2560 1828 2564
rect 994 2559 1000 2560
rect 994 2555 995 2559
rect 999 2555 1000 2559
rect 994 2554 1000 2555
rect 1118 2559 1124 2560
rect 1822 2559 1828 2560
rect 1118 2555 1119 2559
rect 1123 2555 1124 2559
rect 1864 2558 1866 2573
rect 1888 2568 1890 2573
rect 1992 2568 1994 2573
rect 2112 2568 2114 2573
rect 2232 2568 2234 2573
rect 2352 2568 2354 2573
rect 2472 2568 2474 2573
rect 1886 2567 1892 2568
rect 1886 2563 1887 2567
rect 1891 2563 1892 2567
rect 1886 2562 1892 2563
rect 1990 2567 1996 2568
rect 1990 2563 1991 2567
rect 1995 2563 1996 2567
rect 1990 2562 1996 2563
rect 2110 2567 2116 2568
rect 2110 2563 2111 2567
rect 2115 2563 2116 2567
rect 2110 2562 2116 2563
rect 2230 2567 2236 2568
rect 2230 2563 2231 2567
rect 2235 2563 2236 2567
rect 2230 2562 2236 2563
rect 2350 2567 2356 2568
rect 2350 2563 2351 2567
rect 2355 2563 2356 2567
rect 2350 2562 2356 2563
rect 2470 2567 2476 2568
rect 2470 2563 2471 2567
rect 2475 2563 2476 2567
rect 2470 2562 2476 2563
rect 1118 2554 1124 2555
rect 1862 2557 1868 2558
rect 1862 2553 1863 2557
rect 1867 2553 1868 2557
rect 1862 2552 1868 2553
rect 886 2547 892 2548
rect 886 2543 887 2547
rect 891 2543 892 2547
rect 886 2542 892 2543
rect 1822 2547 1828 2548
rect 1822 2543 1823 2547
rect 1827 2543 1828 2547
rect 1822 2542 1828 2543
rect 1954 2543 1960 2544
rect 871 2526 875 2527
rect 871 2521 875 2522
rect 872 2516 874 2521
rect 870 2515 876 2516
rect 870 2511 871 2515
rect 875 2511 876 2515
rect 870 2510 876 2511
rect 662 2507 668 2508
rect 110 2505 116 2506
rect 110 2501 111 2505
rect 115 2501 116 2505
rect 662 2503 663 2507
rect 667 2503 668 2507
rect 662 2502 668 2503
rect 814 2507 820 2508
rect 814 2503 815 2507
rect 819 2503 820 2507
rect 814 2502 820 2503
rect 110 2500 116 2501
rect 110 2488 116 2489
rect 110 2484 111 2488
rect 115 2484 116 2488
rect 110 2483 116 2484
rect 112 2459 114 2483
rect 142 2475 148 2476
rect 142 2471 143 2475
rect 147 2471 148 2475
rect 142 2470 148 2471
rect 286 2475 292 2476
rect 286 2471 287 2475
rect 291 2471 292 2475
rect 286 2470 292 2471
rect 446 2475 452 2476
rect 446 2471 447 2475
rect 451 2471 452 2475
rect 446 2470 452 2471
rect 598 2475 604 2476
rect 598 2471 599 2475
rect 603 2471 604 2475
rect 598 2470 604 2471
rect 742 2475 748 2476
rect 742 2471 743 2475
rect 747 2471 748 2475
rect 742 2470 748 2471
rect 878 2475 884 2476
rect 878 2471 879 2475
rect 883 2471 884 2475
rect 878 2470 884 2471
rect 144 2459 146 2470
rect 288 2459 290 2470
rect 448 2459 450 2470
rect 582 2463 588 2464
rect 582 2459 583 2463
rect 587 2459 588 2463
rect 600 2459 602 2470
rect 744 2459 746 2470
rect 794 2463 800 2464
rect 794 2459 795 2463
rect 799 2459 800 2463
rect 880 2459 882 2470
rect 888 2464 890 2542
rect 918 2537 924 2538
rect 918 2533 919 2537
rect 923 2533 924 2537
rect 918 2532 924 2533
rect 1038 2537 1044 2538
rect 1038 2533 1039 2537
rect 1043 2533 1044 2537
rect 1038 2532 1044 2533
rect 1166 2537 1172 2538
rect 1166 2533 1167 2537
rect 1171 2533 1172 2537
rect 1166 2532 1172 2533
rect 920 2527 922 2532
rect 1040 2527 1042 2532
rect 1168 2527 1170 2532
rect 1824 2527 1826 2542
rect 1862 2540 1868 2541
rect 1862 2536 1863 2540
rect 1867 2536 1868 2540
rect 1954 2539 1955 2543
rect 1959 2539 1960 2543
rect 1954 2538 1960 2539
rect 2178 2543 2184 2544
rect 2178 2539 2179 2543
rect 2183 2539 2184 2543
rect 2178 2538 2184 2539
rect 2326 2543 2332 2544
rect 2326 2539 2327 2543
rect 2331 2539 2332 2543
rect 2326 2538 2332 2539
rect 1862 2535 1868 2536
rect 919 2526 923 2527
rect 919 2521 923 2522
rect 1007 2526 1011 2527
rect 1007 2521 1011 2522
rect 1039 2526 1043 2527
rect 1039 2521 1043 2522
rect 1143 2526 1147 2527
rect 1143 2521 1147 2522
rect 1167 2526 1171 2527
rect 1167 2521 1171 2522
rect 1279 2526 1283 2527
rect 1279 2521 1283 2522
rect 1823 2526 1827 2527
rect 1823 2521 1827 2522
rect 1008 2516 1010 2521
rect 1144 2516 1146 2521
rect 1280 2516 1282 2521
rect 1006 2515 1012 2516
rect 1006 2511 1007 2515
rect 1011 2511 1012 2515
rect 1006 2510 1012 2511
rect 1142 2515 1148 2516
rect 1142 2511 1143 2515
rect 1147 2511 1148 2515
rect 1142 2510 1148 2511
rect 1278 2515 1284 2516
rect 1278 2511 1279 2515
rect 1283 2511 1284 2515
rect 1278 2510 1284 2511
rect 1218 2507 1224 2508
rect 1218 2503 1219 2507
rect 1223 2503 1224 2507
rect 1824 2506 1826 2521
rect 1864 2507 1866 2535
rect 1894 2527 1900 2528
rect 1894 2523 1895 2527
rect 1899 2523 1900 2527
rect 1894 2522 1900 2523
rect 1896 2507 1898 2522
rect 1956 2516 1958 2538
rect 1998 2527 2004 2528
rect 1998 2523 1999 2527
rect 2003 2523 2004 2527
rect 1998 2522 2004 2523
rect 2118 2527 2124 2528
rect 2118 2523 2119 2527
rect 2123 2523 2124 2527
rect 2118 2522 2124 2523
rect 1954 2515 1960 2516
rect 1954 2511 1955 2515
rect 1959 2511 1960 2515
rect 1954 2510 1960 2511
rect 2000 2507 2002 2522
rect 2120 2507 2122 2522
rect 2180 2516 2182 2538
rect 2238 2527 2244 2528
rect 2238 2523 2239 2527
rect 2243 2523 2244 2527
rect 2238 2522 2244 2523
rect 2178 2515 2184 2516
rect 2178 2511 2179 2515
rect 2183 2511 2184 2515
rect 2178 2510 2184 2511
rect 2240 2507 2242 2522
rect 2328 2516 2330 2538
rect 2358 2527 2364 2528
rect 2358 2523 2359 2527
rect 2363 2523 2364 2527
rect 2358 2522 2364 2523
rect 2478 2527 2484 2528
rect 2478 2523 2479 2527
rect 2483 2523 2484 2527
rect 2478 2522 2484 2523
rect 2326 2515 2332 2516
rect 2326 2511 2327 2515
rect 2331 2511 2332 2515
rect 2326 2510 2332 2511
rect 2334 2515 2340 2516
rect 2334 2511 2335 2515
rect 2339 2511 2340 2515
rect 2334 2510 2340 2511
rect 1863 2506 1867 2507
rect 1218 2502 1224 2503
rect 1822 2505 1828 2506
rect 1014 2475 1020 2476
rect 1014 2471 1015 2475
rect 1019 2471 1020 2475
rect 1014 2470 1020 2471
rect 1150 2475 1156 2476
rect 1150 2471 1151 2475
rect 1155 2471 1156 2475
rect 1150 2470 1156 2471
rect 1007 2468 1011 2469
rect 886 2463 892 2464
rect 1007 2463 1011 2464
rect 886 2459 887 2463
rect 891 2459 892 2463
rect 111 2458 115 2459
rect 111 2453 115 2454
rect 143 2458 147 2459
rect 143 2453 147 2454
rect 191 2458 195 2459
rect 191 2453 195 2454
rect 287 2458 291 2459
rect 287 2453 291 2454
rect 319 2458 323 2459
rect 319 2453 323 2454
rect 447 2458 451 2459
rect 447 2453 451 2454
rect 455 2458 459 2459
rect 582 2458 588 2459
rect 591 2458 595 2459
rect 455 2453 459 2454
rect 112 2429 114 2453
rect 192 2442 194 2453
rect 258 2451 264 2452
rect 258 2447 259 2451
rect 263 2447 264 2451
rect 258 2446 264 2447
rect 190 2441 196 2442
rect 190 2437 191 2441
rect 195 2437 196 2441
rect 190 2436 196 2437
rect 110 2428 116 2429
rect 110 2424 111 2428
rect 115 2424 116 2428
rect 260 2424 262 2446
rect 320 2442 322 2453
rect 390 2451 396 2452
rect 390 2447 391 2451
rect 395 2447 396 2451
rect 390 2446 396 2447
rect 318 2441 324 2442
rect 318 2437 319 2441
rect 323 2437 324 2441
rect 318 2436 324 2437
rect 392 2424 394 2446
rect 456 2442 458 2453
rect 454 2441 460 2442
rect 454 2437 455 2441
rect 459 2437 460 2441
rect 454 2436 460 2437
rect 584 2424 586 2458
rect 591 2453 595 2454
rect 599 2458 603 2459
rect 599 2453 603 2454
rect 727 2458 731 2459
rect 727 2453 731 2454
rect 743 2458 747 2459
rect 794 2458 800 2459
rect 863 2458 867 2459
rect 743 2453 747 2454
rect 592 2442 594 2453
rect 678 2451 684 2452
rect 678 2447 679 2451
rect 683 2447 684 2451
rect 678 2446 684 2447
rect 590 2441 596 2442
rect 590 2437 591 2441
rect 595 2437 596 2441
rect 590 2436 596 2437
rect 680 2424 682 2446
rect 728 2442 730 2453
rect 766 2451 772 2452
rect 766 2447 767 2451
rect 771 2447 772 2451
rect 766 2446 772 2447
rect 726 2441 732 2442
rect 726 2437 727 2441
rect 731 2437 732 2441
rect 726 2436 732 2437
rect 110 2423 116 2424
rect 258 2423 264 2424
rect 258 2419 259 2423
rect 263 2419 264 2423
rect 258 2418 264 2419
rect 390 2423 396 2424
rect 390 2419 391 2423
rect 395 2419 396 2423
rect 390 2418 396 2419
rect 582 2423 588 2424
rect 582 2419 583 2423
rect 587 2419 588 2423
rect 582 2418 588 2419
rect 678 2423 684 2424
rect 678 2419 679 2423
rect 683 2419 684 2423
rect 678 2418 684 2419
rect 110 2411 116 2412
rect 110 2407 111 2411
rect 115 2407 116 2411
rect 110 2406 116 2407
rect 174 2411 180 2412
rect 174 2407 175 2411
rect 179 2407 180 2411
rect 174 2406 180 2407
rect 112 2379 114 2406
rect 111 2378 115 2379
rect 111 2373 115 2374
rect 159 2378 163 2379
rect 159 2373 163 2374
rect 112 2358 114 2373
rect 160 2368 162 2373
rect 158 2367 164 2368
rect 158 2363 159 2367
rect 163 2363 164 2367
rect 158 2362 164 2363
rect 110 2357 116 2358
rect 110 2353 111 2357
rect 115 2353 116 2357
rect 110 2352 116 2353
rect 110 2340 116 2341
rect 110 2336 111 2340
rect 115 2336 116 2340
rect 110 2335 116 2336
rect 112 2303 114 2335
rect 166 2327 172 2328
rect 166 2323 167 2327
rect 171 2323 172 2327
rect 166 2322 172 2323
rect 168 2303 170 2322
rect 176 2316 178 2406
rect 182 2401 188 2402
rect 182 2397 183 2401
rect 187 2397 188 2401
rect 182 2396 188 2397
rect 310 2401 316 2402
rect 310 2397 311 2401
rect 315 2397 316 2401
rect 310 2396 316 2397
rect 446 2401 452 2402
rect 446 2397 447 2401
rect 451 2397 452 2401
rect 446 2396 452 2397
rect 582 2401 588 2402
rect 582 2397 583 2401
rect 587 2397 588 2401
rect 582 2396 588 2397
rect 718 2401 724 2402
rect 718 2397 719 2401
rect 723 2397 724 2401
rect 718 2396 724 2397
rect 184 2379 186 2396
rect 312 2379 314 2396
rect 448 2379 450 2396
rect 584 2379 586 2396
rect 720 2379 722 2396
rect 183 2378 187 2379
rect 183 2373 187 2374
rect 247 2378 251 2379
rect 247 2373 251 2374
rect 311 2378 315 2379
rect 311 2373 315 2374
rect 335 2378 339 2379
rect 335 2373 339 2374
rect 439 2378 443 2379
rect 439 2373 443 2374
rect 447 2378 451 2379
rect 447 2373 451 2374
rect 559 2378 563 2379
rect 559 2373 563 2374
rect 583 2378 587 2379
rect 583 2373 587 2374
rect 687 2378 691 2379
rect 687 2373 691 2374
rect 719 2378 723 2379
rect 719 2373 723 2374
rect 248 2368 250 2373
rect 336 2368 338 2373
rect 440 2368 442 2373
rect 560 2368 562 2373
rect 688 2368 690 2373
rect 246 2367 252 2368
rect 246 2363 247 2367
rect 251 2363 252 2367
rect 246 2362 252 2363
rect 334 2367 340 2368
rect 334 2363 335 2367
rect 339 2363 340 2367
rect 334 2362 340 2363
rect 438 2367 444 2368
rect 438 2363 439 2367
rect 443 2363 444 2367
rect 438 2362 444 2363
rect 558 2367 564 2368
rect 558 2363 559 2367
rect 563 2363 564 2367
rect 558 2362 564 2363
rect 686 2367 692 2368
rect 686 2363 687 2367
rect 691 2363 692 2367
rect 686 2362 692 2363
rect 768 2360 770 2446
rect 796 2424 798 2458
rect 863 2453 867 2454
rect 879 2458 883 2459
rect 886 2458 892 2459
rect 999 2458 1003 2459
rect 879 2453 883 2454
rect 999 2453 1003 2454
rect 864 2442 866 2453
rect 886 2451 892 2452
rect 886 2447 887 2451
rect 891 2447 892 2451
rect 886 2446 892 2447
rect 862 2441 868 2442
rect 862 2437 863 2441
rect 867 2437 868 2441
rect 862 2436 868 2437
rect 794 2423 800 2424
rect 794 2419 795 2423
rect 799 2419 800 2423
rect 794 2418 800 2419
rect 854 2401 860 2402
rect 854 2397 855 2401
rect 859 2397 860 2401
rect 854 2396 860 2397
rect 856 2379 858 2396
rect 815 2378 819 2379
rect 815 2373 819 2374
rect 855 2378 859 2379
rect 855 2373 859 2374
rect 816 2368 818 2373
rect 814 2367 820 2368
rect 814 2363 815 2367
rect 819 2363 820 2367
rect 814 2362 820 2363
rect 888 2360 890 2446
rect 1000 2442 1002 2453
rect 1008 2452 1010 2463
rect 1016 2459 1018 2470
rect 1152 2459 1154 2470
rect 1220 2469 1222 2502
rect 1822 2501 1823 2505
rect 1827 2501 1828 2505
rect 1863 2501 1867 2502
rect 1895 2506 1899 2507
rect 1895 2501 1899 2502
rect 1999 2506 2003 2507
rect 1999 2501 2003 2502
rect 2031 2506 2035 2507
rect 2031 2501 2035 2502
rect 2119 2506 2123 2507
rect 2119 2501 2123 2502
rect 2191 2506 2195 2507
rect 2191 2501 2195 2502
rect 2239 2506 2243 2507
rect 2239 2501 2243 2502
rect 1822 2500 1828 2501
rect 1822 2488 1828 2489
rect 1822 2484 1823 2488
rect 1827 2484 1828 2488
rect 1822 2483 1828 2484
rect 1286 2475 1292 2476
rect 1286 2471 1287 2475
rect 1291 2471 1292 2475
rect 1286 2470 1292 2471
rect 1219 2468 1223 2469
rect 1219 2463 1223 2464
rect 1288 2459 1290 2470
rect 1824 2459 1826 2483
rect 1864 2477 1866 2501
rect 1896 2490 1898 2501
rect 2032 2490 2034 2501
rect 2192 2490 2194 2501
rect 1894 2489 1900 2490
rect 1894 2485 1895 2489
rect 1899 2485 1900 2489
rect 1894 2484 1900 2485
rect 2030 2489 2036 2490
rect 2030 2485 2031 2489
rect 2035 2485 2036 2489
rect 2030 2484 2036 2485
rect 2190 2489 2196 2490
rect 2190 2485 2191 2489
rect 2195 2485 2196 2489
rect 2190 2484 2196 2485
rect 1862 2476 1868 2477
rect 1862 2472 1863 2476
rect 1867 2472 1868 2476
rect 2336 2472 2338 2510
rect 2360 2507 2362 2522
rect 2480 2507 2482 2522
rect 2488 2516 2490 2582
rect 2544 2579 2546 2588
rect 2648 2579 2650 2588
rect 2752 2579 2754 2588
rect 2856 2579 2858 2588
rect 3576 2579 3578 2598
rect 2543 2578 2547 2579
rect 2543 2573 2547 2574
rect 2591 2578 2595 2579
rect 2591 2573 2595 2574
rect 2647 2578 2651 2579
rect 2647 2573 2651 2574
rect 2711 2578 2715 2579
rect 2711 2573 2715 2574
rect 2751 2578 2755 2579
rect 2751 2573 2755 2574
rect 2831 2578 2835 2579
rect 2831 2573 2835 2574
rect 2855 2578 2859 2579
rect 2855 2573 2859 2574
rect 3575 2578 3579 2579
rect 3575 2573 3579 2574
rect 2592 2568 2594 2573
rect 2712 2568 2714 2573
rect 2832 2568 2834 2573
rect 2590 2567 2596 2568
rect 2590 2563 2591 2567
rect 2595 2563 2596 2567
rect 2590 2562 2596 2563
rect 2710 2567 2716 2568
rect 2710 2563 2711 2567
rect 2715 2563 2716 2567
rect 2710 2562 2716 2563
rect 2830 2567 2836 2568
rect 2830 2563 2831 2567
rect 2835 2563 2836 2567
rect 2830 2562 2836 2563
rect 2778 2559 2784 2560
rect 2778 2555 2779 2559
rect 2783 2555 2784 2559
rect 3576 2558 3578 2573
rect 2778 2554 2784 2555
rect 3574 2557 3580 2558
rect 2598 2527 2604 2528
rect 2495 2524 2499 2525
rect 2598 2523 2599 2527
rect 2603 2523 2604 2527
rect 2598 2522 2604 2523
rect 2718 2527 2724 2528
rect 2718 2523 2719 2527
rect 2723 2523 2724 2527
rect 2780 2525 2782 2554
rect 3574 2553 3575 2557
rect 3579 2553 3580 2557
rect 3574 2552 3580 2553
rect 3574 2540 3580 2541
rect 3574 2536 3575 2540
rect 3579 2536 3580 2540
rect 3574 2535 3580 2536
rect 2838 2527 2844 2528
rect 2718 2522 2724 2523
rect 2779 2524 2783 2525
rect 2495 2519 2499 2520
rect 2486 2515 2492 2516
rect 2486 2511 2487 2515
rect 2491 2511 2492 2515
rect 2486 2510 2492 2511
rect 2343 2506 2347 2507
rect 2343 2501 2347 2502
rect 2359 2506 2363 2507
rect 2359 2501 2363 2502
rect 2479 2506 2483 2507
rect 2479 2501 2483 2502
rect 2487 2506 2491 2507
rect 2487 2501 2491 2502
rect 2344 2490 2346 2501
rect 2488 2490 2490 2501
rect 2496 2500 2498 2519
rect 2600 2507 2602 2522
rect 2720 2507 2722 2522
rect 2838 2523 2839 2527
rect 2843 2523 2844 2527
rect 2838 2522 2844 2523
rect 2779 2519 2783 2520
rect 2840 2507 2842 2522
rect 3576 2507 3578 2535
rect 2599 2506 2603 2507
rect 2599 2501 2603 2502
rect 2623 2506 2627 2507
rect 2623 2501 2627 2502
rect 2719 2506 2723 2507
rect 2719 2501 2723 2502
rect 2751 2506 2755 2507
rect 2751 2501 2755 2502
rect 2839 2506 2843 2507
rect 2839 2501 2843 2502
rect 2879 2506 2883 2507
rect 2879 2501 2883 2502
rect 3015 2506 3019 2507
rect 3015 2501 3019 2502
rect 3575 2506 3579 2507
rect 3575 2501 3579 2502
rect 2494 2499 2500 2500
rect 2494 2495 2495 2499
rect 2499 2495 2500 2499
rect 2494 2494 2500 2495
rect 2624 2490 2626 2501
rect 2752 2490 2754 2501
rect 2880 2490 2882 2501
rect 3016 2490 3018 2501
rect 2342 2489 2348 2490
rect 2342 2485 2343 2489
rect 2347 2485 2348 2489
rect 2342 2484 2348 2485
rect 2486 2489 2492 2490
rect 2486 2485 2487 2489
rect 2491 2485 2492 2489
rect 2486 2484 2492 2485
rect 2622 2489 2628 2490
rect 2622 2485 2623 2489
rect 2627 2485 2628 2489
rect 2622 2484 2628 2485
rect 2750 2489 2756 2490
rect 2750 2485 2751 2489
rect 2755 2485 2756 2489
rect 2750 2484 2756 2485
rect 2878 2489 2884 2490
rect 2878 2485 2879 2489
rect 2883 2485 2884 2489
rect 2878 2484 2884 2485
rect 3014 2489 3020 2490
rect 3014 2485 3015 2489
rect 3019 2485 3020 2489
rect 3014 2484 3020 2485
rect 3576 2477 3578 2501
rect 3574 2476 3580 2477
rect 3574 2472 3575 2476
rect 3579 2472 3580 2476
rect 1862 2471 1868 2472
rect 2334 2471 2340 2472
rect 3574 2471 3580 2472
rect 2334 2467 2335 2471
rect 2339 2467 2340 2471
rect 2334 2466 2340 2467
rect 1862 2459 1868 2460
rect 1015 2458 1019 2459
rect 1015 2453 1019 2454
rect 1135 2458 1139 2459
rect 1135 2453 1139 2454
rect 1151 2458 1155 2459
rect 1151 2453 1155 2454
rect 1271 2458 1275 2459
rect 1271 2453 1275 2454
rect 1287 2458 1291 2459
rect 1287 2453 1291 2454
rect 1407 2458 1411 2459
rect 1407 2453 1411 2454
rect 1823 2458 1827 2459
rect 1862 2455 1863 2459
rect 1867 2455 1868 2459
rect 1862 2454 1868 2455
rect 2030 2459 2036 2460
rect 2030 2455 2031 2459
rect 2035 2455 2036 2459
rect 2030 2454 2036 2455
rect 2966 2459 2972 2460
rect 2966 2455 2967 2459
rect 2971 2455 2972 2459
rect 2966 2454 2972 2455
rect 3574 2459 3580 2460
rect 3574 2455 3575 2459
rect 3579 2455 3580 2459
rect 3574 2454 3580 2455
rect 1823 2453 1827 2454
rect 1006 2451 1012 2452
rect 1006 2447 1007 2451
rect 1011 2447 1012 2451
rect 1006 2446 1012 2447
rect 1136 2442 1138 2453
rect 1272 2442 1274 2453
rect 1408 2442 1410 2453
rect 998 2441 1004 2442
rect 998 2437 999 2441
rect 1003 2437 1004 2441
rect 998 2436 1004 2437
rect 1134 2441 1140 2442
rect 1134 2437 1135 2441
rect 1139 2437 1140 2441
rect 1134 2436 1140 2437
rect 1270 2441 1276 2442
rect 1270 2437 1271 2441
rect 1275 2437 1276 2441
rect 1270 2436 1276 2437
rect 1406 2441 1412 2442
rect 1406 2437 1407 2441
rect 1411 2437 1412 2441
rect 1406 2436 1412 2437
rect 1824 2429 1826 2453
rect 1864 2439 1866 2454
rect 1886 2449 1892 2450
rect 1886 2445 1887 2449
rect 1891 2445 1892 2449
rect 1886 2444 1892 2445
rect 2022 2449 2028 2450
rect 2022 2445 2023 2449
rect 2027 2445 2028 2449
rect 2022 2444 2028 2445
rect 1888 2439 1890 2444
rect 2024 2439 2026 2444
rect 1863 2438 1867 2439
rect 1863 2433 1867 2434
rect 1887 2438 1891 2439
rect 1887 2433 1891 2434
rect 2015 2438 2019 2439
rect 2015 2433 2019 2434
rect 2023 2438 2027 2439
rect 2023 2433 2027 2434
rect 1822 2428 1828 2429
rect 1822 2424 1823 2428
rect 1827 2424 1828 2428
rect 1822 2423 1828 2424
rect 1864 2418 1866 2433
rect 1888 2428 1890 2433
rect 2016 2428 2018 2433
rect 1886 2427 1892 2428
rect 1886 2423 1887 2427
rect 1891 2423 1892 2427
rect 1886 2422 1892 2423
rect 2014 2427 2020 2428
rect 2014 2423 2015 2427
rect 2019 2423 2020 2427
rect 2014 2422 2020 2423
rect 1862 2417 1868 2418
rect 1862 2413 1863 2417
rect 1867 2413 1868 2417
rect 1862 2412 1868 2413
rect 1338 2411 1344 2412
rect 1338 2407 1339 2411
rect 1343 2407 1344 2411
rect 1338 2406 1344 2407
rect 1822 2411 1828 2412
rect 1822 2407 1823 2411
rect 1827 2407 1828 2411
rect 1822 2406 1828 2407
rect 990 2401 996 2402
rect 990 2397 991 2401
rect 995 2397 996 2401
rect 990 2396 996 2397
rect 1126 2401 1132 2402
rect 1126 2397 1127 2401
rect 1131 2397 1132 2401
rect 1126 2396 1132 2397
rect 1262 2401 1268 2402
rect 1262 2397 1263 2401
rect 1267 2397 1268 2401
rect 1262 2396 1268 2397
rect 992 2379 994 2396
rect 1128 2379 1130 2396
rect 1135 2388 1139 2389
rect 1135 2383 1139 2384
rect 951 2378 955 2379
rect 951 2373 955 2374
rect 991 2378 995 2379
rect 991 2373 995 2374
rect 1079 2378 1083 2379
rect 1079 2373 1083 2374
rect 1127 2378 1131 2379
rect 1127 2373 1131 2374
rect 952 2368 954 2373
rect 1080 2368 1082 2373
rect 950 2367 956 2368
rect 950 2363 951 2367
rect 955 2363 956 2367
rect 950 2362 956 2363
rect 1078 2367 1084 2368
rect 1078 2363 1079 2367
rect 1083 2363 1084 2367
rect 1078 2362 1084 2363
rect 766 2359 772 2360
rect 766 2355 767 2359
rect 771 2355 772 2359
rect 766 2354 772 2355
rect 886 2359 892 2360
rect 886 2355 887 2359
rect 891 2355 892 2359
rect 886 2354 892 2355
rect 226 2343 232 2344
rect 226 2339 227 2343
rect 231 2339 232 2343
rect 226 2338 232 2339
rect 314 2343 320 2344
rect 314 2339 315 2343
rect 319 2339 320 2343
rect 314 2338 320 2339
rect 402 2343 408 2344
rect 402 2339 403 2343
rect 407 2339 408 2343
rect 402 2338 408 2339
rect 654 2343 660 2344
rect 654 2339 655 2343
rect 659 2339 660 2343
rect 654 2338 660 2339
rect 762 2343 768 2344
rect 762 2339 763 2343
rect 767 2339 768 2343
rect 762 2338 768 2339
rect 228 2316 230 2338
rect 254 2327 260 2328
rect 254 2323 255 2327
rect 259 2323 260 2327
rect 254 2322 260 2323
rect 174 2315 180 2316
rect 174 2311 175 2315
rect 179 2311 180 2315
rect 174 2310 180 2311
rect 226 2315 232 2316
rect 226 2311 227 2315
rect 231 2311 232 2315
rect 226 2310 232 2311
rect 256 2303 258 2322
rect 316 2316 318 2338
rect 342 2327 348 2328
rect 342 2323 343 2327
rect 347 2323 348 2327
rect 342 2322 348 2323
rect 314 2315 320 2316
rect 314 2311 315 2315
rect 319 2311 320 2315
rect 314 2310 320 2311
rect 344 2303 346 2322
rect 404 2316 406 2338
rect 446 2327 452 2328
rect 446 2323 447 2327
rect 451 2323 452 2327
rect 446 2322 452 2323
rect 566 2327 572 2328
rect 566 2323 567 2327
rect 571 2323 572 2327
rect 566 2322 572 2323
rect 402 2315 408 2316
rect 402 2311 403 2315
rect 407 2311 408 2315
rect 402 2310 408 2311
rect 448 2303 450 2322
rect 568 2303 570 2322
rect 656 2316 658 2338
rect 694 2327 700 2328
rect 694 2323 695 2327
rect 699 2323 700 2327
rect 694 2322 700 2323
rect 654 2315 660 2316
rect 654 2311 655 2315
rect 659 2311 660 2315
rect 654 2310 660 2311
rect 696 2303 698 2322
rect 764 2316 766 2338
rect 822 2327 828 2328
rect 822 2323 823 2327
rect 827 2323 828 2327
rect 822 2322 828 2323
rect 958 2327 964 2328
rect 958 2323 959 2327
rect 963 2323 964 2327
rect 958 2322 964 2323
rect 1086 2327 1092 2328
rect 1086 2323 1087 2327
rect 1091 2323 1092 2327
rect 1086 2322 1092 2323
rect 762 2315 768 2316
rect 762 2311 763 2315
rect 767 2311 768 2315
rect 762 2310 768 2311
rect 824 2303 826 2322
rect 960 2303 962 2322
rect 1088 2303 1090 2322
rect 1136 2316 1138 2383
rect 1264 2379 1266 2396
rect 1340 2389 1342 2406
rect 1398 2401 1404 2402
rect 1398 2397 1399 2401
rect 1403 2397 1404 2401
rect 1398 2396 1404 2397
rect 1339 2388 1343 2389
rect 1339 2383 1343 2384
rect 1400 2379 1402 2396
rect 1824 2379 1826 2406
rect 1954 2403 1960 2404
rect 1862 2400 1868 2401
rect 1862 2396 1863 2400
rect 1867 2396 1868 2400
rect 1954 2399 1955 2403
rect 1959 2399 1960 2403
rect 1954 2398 1960 2399
rect 1962 2403 1968 2404
rect 1962 2399 1963 2403
rect 1967 2399 1968 2403
rect 1962 2398 1968 2399
rect 1862 2395 1868 2396
rect 1207 2378 1211 2379
rect 1207 2373 1211 2374
rect 1263 2378 1267 2379
rect 1263 2373 1267 2374
rect 1327 2378 1331 2379
rect 1327 2373 1331 2374
rect 1399 2378 1403 2379
rect 1399 2373 1403 2374
rect 1455 2378 1459 2379
rect 1455 2373 1459 2374
rect 1583 2378 1587 2379
rect 1583 2373 1587 2374
rect 1823 2378 1827 2379
rect 1823 2373 1827 2374
rect 1208 2368 1210 2373
rect 1328 2368 1330 2373
rect 1456 2368 1458 2373
rect 1584 2368 1586 2373
rect 1206 2367 1212 2368
rect 1206 2363 1207 2367
rect 1211 2363 1212 2367
rect 1206 2362 1212 2363
rect 1326 2367 1332 2368
rect 1326 2363 1327 2367
rect 1331 2363 1332 2367
rect 1326 2362 1332 2363
rect 1454 2367 1460 2368
rect 1454 2363 1455 2367
rect 1459 2363 1460 2367
rect 1454 2362 1460 2363
rect 1582 2367 1588 2368
rect 1582 2363 1583 2367
rect 1587 2363 1588 2367
rect 1582 2362 1588 2363
rect 1522 2359 1528 2360
rect 1522 2355 1523 2359
rect 1527 2355 1528 2359
rect 1824 2358 1826 2373
rect 1864 2367 1866 2395
rect 1894 2387 1900 2388
rect 1894 2383 1895 2387
rect 1899 2383 1900 2387
rect 1894 2382 1900 2383
rect 1896 2367 1898 2382
rect 1863 2366 1867 2367
rect 1863 2361 1867 2362
rect 1895 2366 1899 2367
rect 1895 2361 1899 2362
rect 1927 2366 1931 2367
rect 1927 2361 1931 2362
rect 1522 2354 1528 2355
rect 1822 2357 1828 2358
rect 1154 2343 1160 2344
rect 1154 2339 1155 2343
rect 1159 2339 1160 2343
rect 1154 2338 1160 2339
rect 1402 2343 1408 2344
rect 1402 2339 1403 2343
rect 1407 2339 1408 2343
rect 1402 2338 1408 2339
rect 1156 2316 1158 2338
rect 1214 2327 1220 2328
rect 1214 2323 1215 2327
rect 1219 2323 1220 2327
rect 1214 2322 1220 2323
rect 1334 2327 1340 2328
rect 1334 2323 1335 2327
rect 1339 2323 1340 2327
rect 1334 2322 1340 2323
rect 1183 2316 1187 2317
rect 1134 2315 1140 2316
rect 1134 2311 1135 2315
rect 1139 2311 1140 2315
rect 1134 2310 1140 2311
rect 1154 2315 1160 2316
rect 1154 2311 1155 2315
rect 1159 2311 1160 2315
rect 1183 2311 1187 2312
rect 1154 2310 1160 2311
rect 111 2302 115 2303
rect 111 2297 115 2298
rect 167 2302 171 2303
rect 167 2297 171 2298
rect 255 2302 259 2303
rect 255 2297 259 2298
rect 343 2302 347 2303
rect 343 2297 347 2298
rect 447 2302 451 2303
rect 447 2297 451 2298
rect 567 2302 571 2303
rect 567 2297 571 2298
rect 695 2302 699 2303
rect 695 2297 699 2298
rect 823 2302 827 2303
rect 823 2297 827 2298
rect 863 2302 867 2303
rect 863 2297 867 2298
rect 959 2302 963 2303
rect 959 2297 963 2298
rect 1023 2302 1027 2303
rect 1023 2297 1027 2298
rect 1087 2302 1091 2303
rect 1087 2297 1091 2298
rect 1175 2302 1179 2303
rect 1175 2297 1179 2298
rect 112 2273 114 2297
rect 696 2286 698 2297
rect 702 2295 708 2296
rect 702 2290 703 2295
rect 707 2290 708 2295
rect 703 2287 707 2288
rect 864 2286 866 2297
rect 939 2292 943 2293
rect 939 2287 943 2288
rect 694 2285 700 2286
rect 694 2281 695 2285
rect 699 2281 700 2285
rect 694 2280 700 2281
rect 862 2285 868 2286
rect 862 2281 863 2285
rect 867 2281 868 2285
rect 862 2280 868 2281
rect 110 2272 116 2273
rect 110 2268 111 2272
rect 115 2268 116 2272
rect 940 2268 942 2287
rect 1024 2286 1026 2297
rect 1030 2295 1036 2296
rect 1030 2291 1031 2295
rect 1035 2291 1036 2295
rect 1030 2290 1036 2291
rect 1022 2285 1028 2286
rect 1022 2281 1023 2285
rect 1027 2281 1028 2285
rect 1022 2280 1028 2281
rect 110 2267 116 2268
rect 938 2267 944 2268
rect 938 2263 939 2267
rect 943 2263 944 2267
rect 938 2262 944 2263
rect 110 2255 116 2256
rect 110 2251 111 2255
rect 115 2251 116 2255
rect 110 2250 116 2251
rect 112 2227 114 2250
rect 686 2245 692 2246
rect 686 2241 687 2245
rect 691 2241 692 2245
rect 686 2240 692 2241
rect 854 2245 860 2246
rect 854 2241 855 2245
rect 859 2241 860 2245
rect 854 2240 860 2241
rect 1014 2245 1020 2246
rect 1014 2241 1015 2245
rect 1019 2241 1020 2245
rect 1014 2240 1020 2241
rect 688 2227 690 2240
rect 856 2227 858 2240
rect 1016 2227 1018 2240
rect 111 2226 115 2227
rect 111 2221 115 2222
rect 535 2226 539 2227
rect 535 2221 539 2222
rect 687 2226 691 2227
rect 687 2221 691 2222
rect 719 2226 723 2227
rect 719 2221 723 2222
rect 855 2226 859 2227
rect 855 2221 859 2222
rect 895 2226 899 2227
rect 895 2221 899 2222
rect 1015 2226 1019 2227
rect 1015 2221 1019 2222
rect 112 2206 114 2221
rect 536 2216 538 2221
rect 720 2216 722 2221
rect 896 2216 898 2221
rect 534 2215 540 2216
rect 534 2211 535 2215
rect 539 2211 540 2215
rect 534 2210 540 2211
rect 718 2215 724 2216
rect 718 2211 719 2215
rect 723 2211 724 2215
rect 718 2210 724 2211
rect 894 2215 900 2216
rect 894 2211 895 2215
rect 899 2211 900 2215
rect 894 2210 900 2211
rect 1032 2208 1034 2290
rect 1176 2286 1178 2297
rect 1184 2296 1186 2311
rect 1216 2303 1218 2322
rect 1336 2303 1338 2322
rect 1404 2316 1406 2338
rect 1462 2327 1468 2328
rect 1462 2323 1463 2327
rect 1467 2323 1468 2327
rect 1462 2322 1468 2323
rect 1402 2315 1408 2316
rect 1402 2311 1403 2315
rect 1407 2311 1408 2315
rect 1402 2310 1408 2311
rect 1464 2303 1466 2322
rect 1524 2317 1526 2354
rect 1822 2353 1823 2357
rect 1827 2353 1828 2357
rect 1822 2352 1828 2353
rect 1530 2343 1536 2344
rect 1530 2339 1531 2343
rect 1535 2339 1536 2343
rect 1530 2338 1536 2339
rect 1822 2340 1828 2341
rect 1523 2316 1527 2317
rect 1532 2316 1534 2338
rect 1822 2336 1823 2340
rect 1827 2336 1828 2340
rect 1864 2337 1866 2361
rect 1928 2350 1930 2361
rect 1956 2360 1958 2398
rect 1964 2376 1966 2398
rect 2022 2387 2028 2388
rect 2022 2383 2023 2387
rect 2027 2383 2028 2387
rect 2022 2382 2028 2383
rect 1962 2375 1968 2376
rect 1962 2371 1963 2375
rect 1967 2371 1968 2375
rect 1962 2370 1968 2371
rect 2024 2367 2026 2382
rect 2032 2376 2034 2454
rect 2182 2449 2188 2450
rect 2182 2445 2183 2449
rect 2187 2445 2188 2449
rect 2182 2444 2188 2445
rect 2334 2449 2340 2450
rect 2334 2445 2335 2449
rect 2339 2445 2340 2449
rect 2334 2444 2340 2445
rect 2478 2449 2484 2450
rect 2478 2445 2479 2449
rect 2483 2445 2484 2449
rect 2478 2444 2484 2445
rect 2614 2449 2620 2450
rect 2614 2445 2615 2449
rect 2619 2445 2620 2449
rect 2614 2444 2620 2445
rect 2742 2449 2748 2450
rect 2742 2445 2743 2449
rect 2747 2445 2748 2449
rect 2742 2444 2748 2445
rect 2870 2449 2876 2450
rect 2870 2445 2871 2449
rect 2875 2445 2876 2449
rect 2870 2444 2876 2445
rect 2184 2439 2186 2444
rect 2336 2439 2338 2444
rect 2480 2439 2482 2444
rect 2616 2439 2618 2444
rect 2744 2439 2746 2444
rect 2872 2439 2874 2444
rect 2175 2438 2179 2439
rect 2175 2433 2179 2434
rect 2183 2438 2187 2439
rect 2183 2433 2187 2434
rect 2335 2438 2339 2439
rect 2335 2433 2339 2434
rect 2479 2438 2483 2439
rect 2479 2433 2483 2434
rect 2495 2438 2499 2439
rect 2495 2433 2499 2434
rect 2615 2438 2619 2439
rect 2615 2433 2619 2434
rect 2647 2438 2651 2439
rect 2647 2433 2651 2434
rect 2743 2438 2747 2439
rect 2743 2433 2747 2434
rect 2799 2438 2803 2439
rect 2799 2433 2803 2434
rect 2871 2438 2875 2439
rect 2871 2433 2875 2434
rect 2951 2438 2955 2439
rect 2951 2433 2955 2434
rect 2176 2428 2178 2433
rect 2336 2428 2338 2433
rect 2496 2428 2498 2433
rect 2648 2428 2650 2433
rect 2800 2428 2802 2433
rect 2952 2428 2954 2433
rect 2174 2427 2180 2428
rect 2174 2423 2175 2427
rect 2179 2423 2180 2427
rect 2174 2422 2180 2423
rect 2334 2427 2340 2428
rect 2334 2423 2335 2427
rect 2339 2423 2340 2427
rect 2334 2422 2340 2423
rect 2494 2427 2500 2428
rect 2494 2423 2495 2427
rect 2499 2423 2500 2427
rect 2494 2422 2500 2423
rect 2646 2427 2652 2428
rect 2646 2423 2647 2427
rect 2651 2423 2652 2427
rect 2646 2422 2652 2423
rect 2798 2427 2804 2428
rect 2798 2423 2799 2427
rect 2803 2423 2804 2427
rect 2798 2422 2804 2423
rect 2950 2427 2956 2428
rect 2950 2423 2951 2427
rect 2955 2423 2956 2427
rect 2950 2422 2956 2423
rect 2242 2403 2248 2404
rect 2242 2399 2243 2403
rect 2247 2399 2248 2403
rect 2242 2398 2248 2399
rect 2402 2403 2408 2404
rect 2402 2399 2403 2403
rect 2407 2399 2408 2403
rect 2402 2398 2408 2399
rect 2182 2387 2188 2388
rect 2182 2383 2183 2387
rect 2187 2383 2188 2387
rect 2182 2382 2188 2383
rect 2030 2375 2036 2376
rect 2030 2371 2031 2375
rect 2035 2371 2036 2375
rect 2030 2370 2036 2371
rect 2184 2367 2186 2382
rect 2244 2376 2246 2398
rect 2342 2387 2348 2388
rect 2342 2383 2343 2387
rect 2347 2383 2348 2387
rect 2342 2382 2348 2383
rect 2242 2375 2248 2376
rect 2242 2371 2243 2375
rect 2247 2371 2248 2375
rect 2242 2370 2248 2371
rect 2344 2367 2346 2382
rect 2404 2376 2406 2398
rect 2711 2396 2715 2397
rect 2711 2391 2715 2392
rect 2502 2387 2508 2388
rect 2502 2383 2503 2387
rect 2507 2383 2508 2387
rect 2502 2382 2508 2383
rect 2654 2387 2660 2388
rect 2654 2383 2655 2387
rect 2659 2383 2660 2387
rect 2654 2382 2660 2383
rect 2402 2375 2408 2376
rect 2402 2371 2403 2375
rect 2407 2371 2408 2375
rect 2402 2370 2408 2371
rect 2478 2367 2484 2368
rect 2504 2367 2506 2382
rect 2656 2367 2658 2382
rect 2663 2380 2667 2381
rect 2662 2375 2668 2376
rect 2662 2371 2663 2375
rect 2667 2371 2668 2375
rect 2662 2370 2668 2371
rect 2023 2366 2027 2367
rect 2023 2361 2027 2362
rect 2087 2366 2091 2367
rect 2087 2361 2091 2362
rect 2183 2366 2187 2367
rect 2183 2361 2187 2362
rect 2247 2366 2251 2367
rect 2247 2361 2251 2362
rect 2343 2366 2347 2367
rect 2343 2361 2347 2362
rect 2407 2366 2411 2367
rect 2478 2363 2479 2367
rect 2483 2363 2484 2367
rect 2478 2362 2484 2363
rect 2503 2366 2507 2367
rect 2407 2361 2411 2362
rect 1954 2359 1960 2360
rect 1954 2355 1955 2359
rect 1959 2355 1960 2359
rect 1954 2354 1960 2355
rect 2088 2350 2090 2361
rect 2248 2350 2250 2361
rect 2408 2350 2410 2361
rect 1926 2349 1932 2350
rect 1926 2345 1927 2349
rect 1931 2345 1932 2349
rect 1926 2344 1932 2345
rect 2086 2349 2092 2350
rect 2086 2345 2087 2349
rect 2091 2345 2092 2349
rect 2086 2344 2092 2345
rect 2246 2349 2252 2350
rect 2246 2345 2247 2349
rect 2251 2345 2252 2349
rect 2246 2344 2252 2345
rect 2406 2349 2412 2350
rect 2406 2345 2407 2349
rect 2411 2345 2412 2349
rect 2406 2344 2412 2345
rect 1822 2335 1828 2336
rect 1862 2336 1868 2337
rect 1590 2327 1596 2328
rect 1590 2323 1591 2327
rect 1595 2323 1596 2327
rect 1590 2322 1596 2323
rect 1523 2311 1527 2312
rect 1530 2315 1536 2316
rect 1530 2311 1531 2315
rect 1535 2311 1536 2315
rect 1530 2310 1536 2311
rect 1592 2303 1594 2322
rect 1824 2303 1826 2335
rect 1862 2332 1863 2336
rect 1867 2332 1868 2336
rect 1862 2331 1868 2332
rect 2480 2320 2482 2362
rect 2503 2361 2507 2362
rect 2559 2366 2563 2367
rect 2559 2361 2563 2362
rect 2655 2366 2659 2367
rect 2655 2361 2659 2362
rect 2703 2366 2707 2367
rect 2703 2361 2707 2362
rect 2560 2350 2562 2361
rect 2566 2359 2572 2360
rect 2566 2355 2567 2359
rect 2571 2355 2572 2359
rect 2566 2354 2572 2355
rect 2558 2349 2564 2350
rect 2558 2345 2559 2349
rect 2563 2345 2564 2349
rect 2558 2344 2564 2345
rect 1862 2319 1868 2320
rect 1862 2315 1863 2319
rect 1867 2315 1868 2319
rect 1862 2314 1868 2315
rect 2478 2319 2484 2320
rect 2478 2315 2479 2319
rect 2483 2315 2484 2319
rect 2478 2314 2484 2315
rect 1215 2302 1219 2303
rect 1215 2297 1219 2298
rect 1319 2302 1323 2303
rect 1319 2297 1323 2298
rect 1335 2302 1339 2303
rect 1335 2297 1339 2298
rect 1463 2302 1467 2303
rect 1463 2297 1467 2298
rect 1591 2302 1595 2303
rect 1591 2297 1595 2298
rect 1599 2302 1603 2303
rect 1599 2297 1603 2298
rect 1735 2302 1739 2303
rect 1735 2297 1739 2298
rect 1823 2302 1827 2303
rect 1823 2297 1827 2298
rect 1182 2295 1188 2296
rect 1182 2291 1183 2295
rect 1187 2291 1188 2295
rect 1182 2290 1188 2291
rect 1320 2286 1322 2297
rect 1464 2286 1466 2297
rect 1600 2286 1602 2297
rect 1736 2286 1738 2297
rect 1174 2285 1180 2286
rect 1174 2281 1175 2285
rect 1179 2281 1180 2285
rect 1174 2280 1180 2281
rect 1318 2285 1324 2286
rect 1318 2281 1319 2285
rect 1323 2281 1324 2285
rect 1318 2280 1324 2281
rect 1462 2285 1468 2286
rect 1462 2281 1463 2285
rect 1467 2281 1468 2285
rect 1462 2280 1468 2281
rect 1598 2285 1604 2286
rect 1598 2281 1599 2285
rect 1603 2281 1604 2285
rect 1598 2280 1604 2281
rect 1734 2285 1740 2286
rect 1734 2281 1735 2285
rect 1739 2281 1740 2285
rect 1734 2280 1740 2281
rect 1824 2273 1826 2297
rect 1864 2295 1866 2314
rect 1918 2309 1924 2310
rect 1918 2305 1919 2309
rect 1923 2305 1924 2309
rect 1918 2304 1924 2305
rect 2078 2309 2084 2310
rect 2078 2305 2079 2309
rect 2083 2305 2084 2309
rect 2078 2304 2084 2305
rect 2238 2309 2244 2310
rect 2238 2305 2239 2309
rect 2243 2305 2244 2309
rect 2238 2304 2244 2305
rect 2398 2309 2404 2310
rect 2398 2305 2399 2309
rect 2403 2305 2404 2309
rect 2398 2304 2404 2305
rect 2550 2309 2556 2310
rect 2550 2305 2551 2309
rect 2555 2305 2556 2309
rect 2550 2304 2556 2305
rect 1920 2295 1922 2304
rect 2080 2295 2082 2304
rect 2240 2295 2242 2304
rect 2400 2295 2402 2304
rect 2552 2295 2554 2304
rect 1863 2294 1867 2295
rect 1863 2289 1867 2290
rect 1919 2294 1923 2295
rect 1919 2289 1923 2290
rect 1975 2294 1979 2295
rect 1975 2289 1979 2290
rect 2079 2294 2083 2295
rect 2079 2289 2083 2290
rect 2143 2294 2147 2295
rect 2143 2289 2147 2290
rect 2239 2294 2243 2295
rect 2239 2289 2243 2290
rect 2311 2294 2315 2295
rect 2311 2289 2315 2290
rect 2399 2294 2403 2295
rect 2399 2289 2403 2290
rect 2479 2294 2483 2295
rect 2479 2289 2483 2290
rect 2551 2294 2555 2295
rect 2551 2289 2555 2290
rect 1864 2274 1866 2289
rect 1976 2284 1978 2289
rect 2144 2284 2146 2289
rect 2312 2284 2314 2289
rect 2480 2284 2482 2289
rect 1974 2283 1980 2284
rect 1974 2279 1975 2283
rect 1979 2279 1980 2283
rect 1974 2278 1980 2279
rect 2142 2283 2148 2284
rect 2142 2279 2143 2283
rect 2147 2279 2148 2283
rect 2142 2278 2148 2279
rect 2310 2283 2316 2284
rect 2310 2279 2311 2283
rect 2315 2279 2316 2283
rect 2310 2278 2316 2279
rect 2478 2283 2484 2284
rect 2478 2279 2479 2283
rect 2483 2279 2484 2283
rect 2478 2278 2484 2279
rect 2568 2276 2570 2354
rect 2704 2350 2706 2361
rect 2712 2360 2714 2391
rect 2806 2387 2812 2388
rect 2806 2383 2807 2387
rect 2811 2383 2812 2387
rect 2806 2382 2812 2383
rect 2958 2387 2964 2388
rect 2958 2383 2959 2387
rect 2963 2383 2964 2387
rect 2958 2382 2964 2383
rect 2808 2367 2810 2382
rect 2960 2367 2962 2382
rect 2968 2381 2970 2454
rect 3006 2449 3012 2450
rect 3006 2445 3007 2449
rect 3011 2445 3012 2449
rect 3006 2444 3012 2445
rect 3008 2439 3010 2444
rect 3576 2439 3578 2454
rect 3007 2438 3011 2439
rect 3007 2433 3011 2434
rect 3111 2438 3115 2439
rect 3111 2433 3115 2434
rect 3575 2438 3579 2439
rect 3575 2433 3579 2434
rect 3112 2428 3114 2433
rect 3110 2427 3116 2428
rect 3110 2423 3111 2427
rect 3115 2423 3116 2427
rect 3110 2422 3116 2423
rect 3018 2419 3024 2420
rect 3018 2415 3019 2419
rect 3023 2415 3024 2419
rect 3576 2418 3578 2433
rect 3018 2414 3024 2415
rect 3574 2417 3580 2418
rect 3020 2397 3022 2414
rect 3574 2413 3575 2417
rect 3579 2413 3580 2417
rect 3574 2412 3580 2413
rect 3574 2400 3580 2401
rect 3019 2396 3023 2397
rect 3574 2396 3575 2400
rect 3579 2396 3580 2400
rect 3574 2395 3580 2396
rect 3019 2391 3023 2392
rect 3118 2387 3124 2388
rect 3118 2383 3119 2387
rect 3123 2383 3124 2387
rect 3118 2382 3124 2383
rect 2967 2380 2971 2381
rect 2967 2375 2971 2376
rect 3120 2367 3122 2382
rect 3576 2367 3578 2395
rect 2807 2366 2811 2367
rect 2807 2361 2811 2362
rect 2831 2366 2835 2367
rect 2831 2361 2835 2362
rect 2951 2366 2955 2367
rect 2951 2361 2955 2362
rect 2959 2366 2963 2367
rect 2959 2361 2963 2362
rect 3071 2366 3075 2367
rect 3071 2361 3075 2362
rect 3119 2366 3123 2367
rect 3119 2361 3123 2362
rect 3183 2366 3187 2367
rect 3183 2361 3187 2362
rect 3287 2366 3291 2367
rect 3287 2361 3291 2362
rect 3399 2366 3403 2367
rect 3399 2361 3403 2362
rect 3487 2366 3491 2367
rect 3487 2361 3491 2362
rect 3575 2366 3579 2367
rect 3575 2361 3579 2362
rect 2710 2359 2716 2360
rect 2710 2355 2711 2359
rect 2715 2355 2716 2359
rect 2710 2354 2716 2355
rect 2832 2350 2834 2361
rect 2952 2350 2954 2361
rect 3072 2350 3074 2361
rect 3184 2350 3186 2361
rect 3288 2350 3290 2361
rect 3400 2350 3402 2361
rect 3488 2350 3490 2361
rect 2702 2349 2708 2350
rect 2702 2345 2703 2349
rect 2707 2345 2708 2349
rect 2702 2344 2708 2345
rect 2830 2349 2836 2350
rect 2830 2345 2831 2349
rect 2835 2345 2836 2349
rect 2830 2344 2836 2345
rect 2950 2349 2956 2350
rect 2950 2345 2951 2349
rect 2955 2345 2956 2349
rect 2950 2344 2956 2345
rect 3070 2349 3076 2350
rect 3070 2345 3071 2349
rect 3075 2345 3076 2349
rect 3070 2344 3076 2345
rect 3182 2349 3188 2350
rect 3182 2345 3183 2349
rect 3187 2345 3188 2349
rect 3182 2344 3188 2345
rect 3286 2349 3292 2350
rect 3286 2345 3287 2349
rect 3291 2345 3292 2349
rect 3286 2344 3292 2345
rect 3398 2349 3404 2350
rect 3398 2345 3399 2349
rect 3403 2345 3404 2349
rect 3398 2344 3404 2345
rect 3486 2349 3492 2350
rect 3486 2345 3487 2349
rect 3491 2345 3492 2349
rect 3486 2344 3492 2345
rect 3576 2337 3578 2361
rect 3574 2336 3580 2337
rect 3574 2332 3575 2336
rect 3579 2332 3580 2336
rect 3574 2331 3580 2332
rect 3182 2319 3188 2320
rect 3182 2315 3183 2319
rect 3187 2315 3188 2319
rect 3182 2314 3188 2315
rect 3574 2319 3580 2320
rect 3574 2315 3575 2319
rect 3579 2315 3580 2319
rect 3574 2314 3580 2315
rect 2694 2309 2700 2310
rect 2694 2305 2695 2309
rect 2699 2305 2700 2309
rect 2694 2304 2700 2305
rect 2822 2309 2828 2310
rect 2822 2305 2823 2309
rect 2827 2305 2828 2309
rect 2822 2304 2828 2305
rect 2942 2309 2948 2310
rect 2942 2305 2943 2309
rect 2947 2305 2948 2309
rect 2942 2304 2948 2305
rect 3062 2309 3068 2310
rect 3062 2305 3063 2309
rect 3067 2305 3068 2309
rect 3062 2304 3068 2305
rect 3174 2309 3180 2310
rect 3174 2305 3175 2309
rect 3179 2305 3180 2309
rect 3174 2304 3180 2305
rect 2696 2295 2698 2304
rect 2824 2295 2826 2304
rect 2944 2295 2946 2304
rect 3064 2295 3066 2304
rect 3176 2295 3178 2304
rect 2639 2294 2643 2295
rect 2639 2289 2643 2290
rect 2695 2294 2699 2295
rect 2695 2289 2699 2290
rect 2783 2294 2787 2295
rect 2783 2289 2787 2290
rect 2823 2294 2827 2295
rect 2823 2289 2827 2290
rect 2919 2294 2923 2295
rect 2919 2289 2923 2290
rect 2943 2294 2947 2295
rect 2943 2289 2947 2290
rect 3039 2294 3043 2295
rect 3039 2289 3043 2290
rect 3063 2294 3067 2295
rect 3063 2289 3067 2290
rect 3159 2294 3163 2295
rect 3159 2289 3163 2290
rect 3175 2294 3179 2295
rect 3175 2289 3179 2290
rect 2640 2284 2642 2289
rect 2784 2284 2786 2289
rect 2920 2284 2922 2289
rect 3040 2284 3042 2289
rect 3160 2284 3162 2289
rect 2638 2283 2644 2284
rect 2638 2279 2639 2283
rect 2643 2279 2644 2283
rect 2638 2278 2644 2279
rect 2782 2283 2788 2284
rect 2782 2279 2783 2283
rect 2787 2279 2788 2283
rect 2782 2278 2788 2279
rect 2918 2283 2924 2284
rect 2918 2279 2919 2283
rect 2923 2279 2924 2283
rect 2918 2278 2924 2279
rect 3038 2283 3044 2284
rect 3038 2279 3039 2283
rect 3043 2279 3044 2283
rect 3038 2278 3044 2279
rect 3158 2283 3164 2284
rect 3158 2279 3159 2283
rect 3163 2279 3164 2283
rect 3158 2278 3164 2279
rect 2566 2275 2572 2276
rect 1862 2273 1868 2274
rect 1822 2272 1828 2273
rect 1822 2268 1823 2272
rect 1827 2268 1828 2272
rect 1862 2269 1863 2273
rect 1867 2269 1868 2273
rect 2566 2271 2567 2275
rect 2571 2271 2572 2275
rect 2566 2270 2572 2271
rect 3110 2275 3116 2276
rect 3110 2271 3111 2275
rect 3115 2271 3116 2275
rect 3110 2270 3116 2271
rect 1862 2268 1868 2269
rect 1822 2267 1828 2268
rect 2042 2259 2048 2260
rect 1862 2256 1868 2257
rect 1666 2255 1672 2256
rect 1666 2251 1667 2255
rect 1671 2251 1672 2255
rect 1666 2250 1672 2251
rect 1822 2255 1828 2256
rect 1822 2251 1823 2255
rect 1827 2251 1828 2255
rect 1862 2252 1863 2256
rect 1867 2252 1868 2256
rect 2042 2255 2043 2259
rect 2047 2255 2048 2259
rect 2042 2254 2048 2255
rect 2050 2259 2056 2260
rect 2050 2255 2051 2259
rect 2055 2255 2056 2259
rect 2050 2254 2056 2255
rect 1862 2251 1868 2252
rect 1822 2250 1828 2251
rect 1166 2245 1172 2246
rect 1166 2241 1167 2245
rect 1171 2241 1172 2245
rect 1166 2240 1172 2241
rect 1310 2245 1316 2246
rect 1310 2241 1311 2245
rect 1315 2241 1316 2245
rect 1310 2240 1316 2241
rect 1454 2245 1460 2246
rect 1454 2241 1455 2245
rect 1459 2241 1460 2245
rect 1454 2240 1460 2241
rect 1590 2245 1596 2246
rect 1590 2241 1591 2245
rect 1595 2241 1596 2245
rect 1590 2240 1596 2241
rect 1168 2227 1170 2240
rect 1312 2227 1314 2240
rect 1456 2227 1458 2240
rect 1592 2227 1594 2240
rect 1071 2226 1075 2227
rect 1071 2221 1075 2222
rect 1167 2226 1171 2227
rect 1167 2221 1171 2222
rect 1239 2226 1243 2227
rect 1239 2221 1243 2222
rect 1311 2226 1315 2227
rect 1311 2221 1315 2222
rect 1407 2226 1411 2227
rect 1407 2221 1411 2222
rect 1455 2226 1459 2227
rect 1455 2221 1459 2222
rect 1575 2226 1579 2227
rect 1575 2221 1579 2222
rect 1591 2226 1595 2227
rect 1591 2221 1595 2222
rect 1072 2216 1074 2221
rect 1240 2216 1242 2221
rect 1408 2216 1410 2221
rect 1576 2216 1578 2221
rect 1070 2215 1076 2216
rect 1070 2211 1071 2215
rect 1075 2211 1076 2215
rect 1070 2210 1076 2211
rect 1238 2215 1244 2216
rect 1238 2211 1239 2215
rect 1243 2211 1244 2215
rect 1238 2210 1244 2211
rect 1406 2215 1412 2216
rect 1406 2211 1407 2215
rect 1411 2211 1412 2215
rect 1406 2210 1412 2211
rect 1574 2215 1580 2216
rect 1574 2211 1575 2215
rect 1579 2211 1580 2215
rect 1574 2210 1580 2211
rect 1030 2207 1036 2208
rect 110 2205 116 2206
rect 110 2201 111 2205
rect 115 2201 116 2205
rect 1030 2203 1031 2207
rect 1035 2203 1036 2207
rect 1030 2202 1036 2203
rect 1642 2207 1648 2208
rect 1642 2203 1643 2207
rect 1647 2203 1648 2207
rect 1642 2202 1648 2203
rect 110 2200 116 2201
rect 110 2188 116 2189
rect 110 2184 111 2188
rect 115 2184 116 2188
rect 110 2183 116 2184
rect 112 2159 114 2183
rect 1255 2180 1259 2181
rect 542 2175 548 2176
rect 542 2171 543 2175
rect 547 2171 548 2175
rect 542 2170 548 2171
rect 726 2175 732 2176
rect 726 2171 727 2175
rect 731 2171 732 2175
rect 726 2170 732 2171
rect 902 2175 908 2176
rect 902 2171 903 2175
rect 907 2171 908 2175
rect 902 2170 908 2171
rect 1078 2175 1084 2176
rect 1078 2171 1079 2175
rect 1083 2171 1084 2175
rect 1078 2170 1084 2171
rect 1246 2175 1252 2176
rect 1255 2175 1259 2176
rect 1414 2175 1420 2176
rect 1246 2171 1247 2175
rect 1251 2171 1252 2175
rect 1246 2170 1252 2171
rect 544 2159 546 2170
rect 574 2163 580 2164
rect 574 2159 575 2163
rect 579 2159 580 2163
rect 728 2159 730 2170
rect 904 2159 906 2170
rect 1080 2159 1082 2170
rect 1248 2159 1250 2170
rect 1256 2164 1258 2175
rect 1414 2171 1415 2175
rect 1419 2171 1420 2175
rect 1414 2170 1420 2171
rect 1582 2175 1588 2176
rect 1582 2171 1583 2175
rect 1587 2171 1588 2175
rect 1582 2170 1588 2171
rect 1254 2163 1260 2164
rect 1254 2159 1255 2163
rect 1259 2159 1260 2163
rect 1416 2159 1418 2170
rect 1584 2159 1586 2170
rect 111 2158 115 2159
rect 111 2153 115 2154
rect 495 2158 499 2159
rect 495 2153 499 2154
rect 543 2158 547 2159
rect 574 2158 580 2159
rect 623 2158 627 2159
rect 543 2153 547 2154
rect 112 2129 114 2153
rect 496 2142 498 2153
rect 550 2151 556 2152
rect 550 2146 551 2151
rect 555 2146 556 2151
rect 551 2143 555 2144
rect 494 2141 500 2142
rect 494 2137 495 2141
rect 499 2137 500 2141
rect 494 2136 500 2137
rect 110 2128 116 2129
rect 110 2124 111 2128
rect 115 2124 116 2128
rect 110 2123 116 2124
rect 576 2117 578 2158
rect 623 2153 627 2154
rect 727 2158 731 2159
rect 727 2153 731 2154
rect 759 2158 763 2159
rect 759 2153 763 2154
rect 895 2158 899 2159
rect 895 2153 899 2154
rect 903 2158 907 2159
rect 903 2153 907 2154
rect 1039 2158 1043 2159
rect 1039 2153 1043 2154
rect 1079 2158 1083 2159
rect 1079 2153 1083 2154
rect 1183 2158 1187 2159
rect 1183 2153 1187 2154
rect 1247 2158 1251 2159
rect 1254 2158 1260 2159
rect 1327 2158 1331 2159
rect 1247 2153 1251 2154
rect 1327 2153 1331 2154
rect 1415 2158 1419 2159
rect 1415 2153 1419 2154
rect 1471 2158 1475 2159
rect 1471 2153 1475 2154
rect 1583 2158 1587 2159
rect 1583 2153 1587 2154
rect 1623 2158 1627 2159
rect 1623 2153 1627 2154
rect 624 2142 626 2153
rect 760 2142 762 2153
rect 767 2148 771 2149
rect 767 2143 771 2144
rect 622 2141 628 2142
rect 622 2137 623 2141
rect 627 2137 628 2141
rect 622 2136 628 2137
rect 758 2141 764 2142
rect 758 2137 759 2141
rect 763 2137 764 2141
rect 758 2136 764 2137
rect 575 2116 579 2117
rect 110 2111 116 2112
rect 575 2111 579 2112
rect 110 2107 111 2111
rect 115 2107 116 2111
rect 110 2106 116 2107
rect 112 2087 114 2106
rect 486 2101 492 2102
rect 486 2097 487 2101
rect 491 2097 492 2101
rect 486 2096 492 2097
rect 614 2101 620 2102
rect 614 2097 615 2101
rect 619 2097 620 2101
rect 614 2096 620 2097
rect 750 2101 756 2102
rect 750 2097 751 2101
rect 755 2097 756 2101
rect 750 2096 756 2097
rect 488 2087 490 2096
rect 616 2087 618 2096
rect 752 2087 754 2096
rect 111 2086 115 2087
rect 111 2081 115 2082
rect 319 2086 323 2087
rect 319 2081 323 2082
rect 431 2086 435 2087
rect 431 2081 435 2082
rect 487 2086 491 2087
rect 487 2081 491 2082
rect 551 2086 555 2087
rect 551 2081 555 2082
rect 615 2086 619 2087
rect 615 2081 619 2082
rect 679 2086 683 2087
rect 679 2081 683 2082
rect 751 2086 755 2087
rect 751 2081 755 2082
rect 112 2066 114 2081
rect 320 2076 322 2081
rect 432 2076 434 2081
rect 552 2076 554 2081
rect 680 2076 682 2081
rect 318 2075 324 2076
rect 318 2071 319 2075
rect 323 2071 324 2075
rect 318 2070 324 2071
rect 430 2075 436 2076
rect 430 2071 431 2075
rect 435 2071 436 2075
rect 430 2070 436 2071
rect 550 2075 556 2076
rect 550 2071 551 2075
rect 555 2071 556 2075
rect 550 2070 556 2071
rect 678 2075 684 2076
rect 678 2071 679 2075
rect 683 2071 684 2075
rect 678 2070 684 2071
rect 768 2068 770 2143
rect 896 2142 898 2153
rect 1040 2142 1042 2153
rect 1184 2142 1186 2153
rect 1238 2151 1244 2152
rect 1238 2147 1239 2151
rect 1243 2147 1244 2151
rect 1238 2146 1244 2147
rect 894 2141 900 2142
rect 894 2137 895 2141
rect 899 2137 900 2141
rect 894 2136 900 2137
rect 1038 2141 1044 2142
rect 1038 2137 1039 2141
rect 1043 2137 1044 2141
rect 1038 2136 1044 2137
rect 1182 2141 1188 2142
rect 1182 2137 1183 2141
rect 1187 2137 1188 2141
rect 1182 2136 1188 2137
rect 1038 2111 1044 2112
rect 1038 2106 1039 2111
rect 1043 2106 1044 2111
rect 1039 2103 1043 2104
rect 886 2101 892 2102
rect 886 2097 887 2101
rect 891 2097 892 2101
rect 886 2096 892 2097
rect 1030 2101 1036 2102
rect 1030 2097 1031 2101
rect 1035 2097 1036 2101
rect 1030 2096 1036 2097
rect 1174 2101 1180 2102
rect 1174 2097 1175 2101
rect 1179 2097 1180 2101
rect 1174 2096 1180 2097
rect 1240 2096 1242 2146
rect 1328 2142 1330 2153
rect 1472 2142 1474 2153
rect 1538 2151 1544 2152
rect 1538 2147 1539 2151
rect 1543 2147 1544 2151
rect 1538 2146 1544 2147
rect 1326 2141 1332 2142
rect 1326 2137 1327 2141
rect 1331 2137 1332 2141
rect 1326 2136 1332 2137
rect 1470 2141 1476 2142
rect 1470 2137 1471 2141
rect 1475 2137 1476 2141
rect 1470 2136 1476 2137
rect 1540 2124 1542 2146
rect 1624 2142 1626 2153
rect 1644 2152 1646 2202
rect 1668 2181 1670 2250
rect 1726 2245 1732 2246
rect 1726 2241 1727 2245
rect 1731 2241 1732 2245
rect 1726 2240 1732 2241
rect 1728 2227 1730 2240
rect 1824 2227 1826 2250
rect 1864 2227 1866 2251
rect 1982 2243 1988 2244
rect 1982 2239 1983 2243
rect 1987 2239 1988 2243
rect 1982 2238 1988 2239
rect 1984 2227 1986 2238
rect 1727 2226 1731 2227
rect 1727 2221 1731 2222
rect 1823 2226 1827 2227
rect 1823 2221 1827 2222
rect 1863 2226 1867 2227
rect 1863 2221 1867 2222
rect 1983 2226 1987 2227
rect 1983 2221 1987 2222
rect 2007 2226 2011 2227
rect 2007 2221 2011 2222
rect 1728 2216 1730 2221
rect 1726 2215 1732 2216
rect 1726 2211 1727 2215
rect 1731 2211 1732 2215
rect 1726 2210 1732 2211
rect 1824 2206 1826 2221
rect 1822 2205 1828 2206
rect 1822 2201 1823 2205
rect 1827 2201 1828 2205
rect 1822 2200 1828 2201
rect 1864 2197 1866 2221
rect 2008 2210 2010 2221
rect 2044 2220 2046 2254
rect 2052 2232 2054 2254
rect 2150 2243 2156 2244
rect 2150 2239 2151 2243
rect 2155 2239 2156 2243
rect 2150 2238 2156 2239
rect 2318 2243 2324 2244
rect 2318 2239 2319 2243
rect 2323 2239 2324 2243
rect 2318 2238 2324 2239
rect 2486 2243 2492 2244
rect 2486 2239 2487 2243
rect 2491 2239 2492 2243
rect 2486 2238 2492 2239
rect 2646 2243 2652 2244
rect 2646 2239 2647 2243
rect 2651 2239 2652 2243
rect 2646 2238 2652 2239
rect 2790 2243 2796 2244
rect 2790 2239 2791 2243
rect 2795 2239 2796 2243
rect 2790 2238 2796 2239
rect 2926 2243 2932 2244
rect 2926 2239 2927 2243
rect 2931 2239 2932 2243
rect 2926 2238 2932 2239
rect 3046 2243 3052 2244
rect 3046 2239 3047 2243
rect 3051 2239 3052 2243
rect 3046 2238 3052 2239
rect 2050 2231 2056 2232
rect 2050 2227 2051 2231
rect 2055 2227 2056 2231
rect 2152 2227 2154 2238
rect 2320 2227 2322 2238
rect 2402 2231 2408 2232
rect 2402 2227 2403 2231
rect 2407 2227 2408 2231
rect 2488 2227 2490 2238
rect 2648 2227 2650 2238
rect 2792 2227 2794 2238
rect 2799 2236 2803 2237
rect 2798 2231 2804 2232
rect 2798 2227 2799 2231
rect 2803 2227 2804 2231
rect 2928 2227 2930 2238
rect 3048 2227 3050 2238
rect 2050 2226 2056 2227
rect 2151 2226 2155 2227
rect 2151 2221 2155 2222
rect 2167 2226 2171 2227
rect 2167 2221 2171 2222
rect 2319 2226 2323 2227
rect 2319 2221 2323 2222
rect 2335 2226 2339 2227
rect 2402 2226 2408 2227
rect 2487 2226 2491 2227
rect 2335 2221 2339 2222
rect 2042 2219 2048 2220
rect 2042 2215 2043 2219
rect 2047 2215 2048 2219
rect 2042 2214 2048 2215
rect 2168 2210 2170 2221
rect 2336 2210 2338 2221
rect 2006 2209 2012 2210
rect 2006 2205 2007 2209
rect 2011 2205 2012 2209
rect 2006 2204 2012 2205
rect 2166 2209 2172 2210
rect 2166 2205 2167 2209
rect 2171 2205 2172 2209
rect 2166 2204 2172 2205
rect 2334 2209 2340 2210
rect 2334 2205 2335 2209
rect 2339 2205 2340 2209
rect 2334 2204 2340 2205
rect 1862 2196 1868 2197
rect 1862 2192 1863 2196
rect 1867 2192 1868 2196
rect 2404 2192 2406 2226
rect 2487 2221 2491 2222
rect 2519 2226 2523 2227
rect 2519 2221 2523 2222
rect 2647 2226 2651 2227
rect 2647 2221 2651 2222
rect 2711 2226 2715 2227
rect 2711 2221 2715 2222
rect 2791 2226 2795 2227
rect 2798 2226 2804 2227
rect 2903 2226 2907 2227
rect 2791 2221 2795 2222
rect 2903 2221 2907 2222
rect 2927 2226 2931 2227
rect 2927 2221 2931 2222
rect 3047 2226 3051 2227
rect 3047 2221 3051 2222
rect 3103 2226 3107 2227
rect 3103 2221 3107 2222
rect 2520 2210 2522 2221
rect 2586 2219 2592 2220
rect 2586 2215 2587 2219
rect 2591 2215 2592 2219
rect 2586 2214 2592 2215
rect 2518 2209 2524 2210
rect 2518 2205 2519 2209
rect 2523 2205 2524 2209
rect 2518 2204 2524 2205
rect 2588 2192 2590 2214
rect 2712 2210 2714 2221
rect 2838 2219 2844 2220
rect 2838 2215 2839 2219
rect 2843 2215 2844 2219
rect 2838 2214 2844 2215
rect 2710 2209 2716 2210
rect 2710 2205 2711 2209
rect 2715 2205 2716 2209
rect 2710 2204 2716 2205
rect 1862 2191 1868 2192
rect 2402 2191 2408 2192
rect 1822 2188 1828 2189
rect 1822 2184 1823 2188
rect 1827 2184 1828 2188
rect 2402 2187 2403 2191
rect 2407 2187 2408 2191
rect 2402 2186 2408 2187
rect 2586 2191 2592 2192
rect 2586 2187 2587 2191
rect 2591 2187 2592 2191
rect 2586 2186 2592 2187
rect 1822 2183 1828 2184
rect 1667 2180 1671 2181
rect 1667 2175 1671 2176
rect 1734 2175 1740 2176
rect 1734 2171 1735 2175
rect 1739 2171 1740 2175
rect 1734 2170 1740 2171
rect 1736 2159 1738 2170
rect 1824 2159 1826 2183
rect 1862 2179 1868 2180
rect 1862 2175 1863 2179
rect 1867 2175 1868 2179
rect 1862 2174 1868 2175
rect 2234 2179 2240 2180
rect 2234 2175 2235 2179
rect 2239 2175 2240 2179
rect 2234 2174 2240 2175
rect 1735 2158 1739 2159
rect 1735 2153 1739 2154
rect 1823 2158 1827 2159
rect 1823 2153 1827 2154
rect 1642 2151 1648 2152
rect 1642 2147 1643 2151
rect 1647 2147 1648 2151
rect 1642 2146 1648 2147
rect 1622 2141 1628 2142
rect 1622 2137 1623 2141
rect 1627 2137 1628 2141
rect 1622 2136 1628 2137
rect 1824 2129 1826 2153
rect 1864 2151 1866 2174
rect 1998 2169 2004 2170
rect 1998 2165 1999 2169
rect 2003 2165 2004 2169
rect 1998 2164 2004 2165
rect 2158 2169 2164 2170
rect 2158 2165 2159 2169
rect 2163 2165 2164 2169
rect 2158 2164 2164 2165
rect 2000 2151 2002 2164
rect 2160 2151 2162 2164
rect 1863 2150 1867 2151
rect 1863 2145 1867 2146
rect 1999 2150 2003 2151
rect 1999 2145 2003 2146
rect 2023 2150 2027 2151
rect 2023 2145 2027 2146
rect 2159 2150 2163 2151
rect 2159 2145 2163 2146
rect 2167 2150 2171 2151
rect 2167 2145 2171 2146
rect 1864 2130 1866 2145
rect 2024 2140 2026 2145
rect 2168 2140 2170 2145
rect 2022 2139 2028 2140
rect 2022 2135 2023 2139
rect 2027 2135 2028 2139
rect 2022 2134 2028 2135
rect 2166 2139 2172 2140
rect 2166 2135 2167 2139
rect 2171 2135 2172 2139
rect 2166 2134 2172 2135
rect 1862 2129 1868 2130
rect 1822 2128 1828 2129
rect 1822 2124 1823 2128
rect 1827 2124 1828 2128
rect 1862 2125 1863 2129
rect 1867 2125 1868 2129
rect 1862 2124 1868 2125
rect 1538 2123 1544 2124
rect 1822 2123 1828 2124
rect 1538 2119 1539 2123
rect 1543 2119 1544 2123
rect 1538 2118 1544 2119
rect 2106 2115 2112 2116
rect 1862 2112 1868 2113
rect 1398 2111 1404 2112
rect 1398 2107 1399 2111
rect 1403 2107 1404 2111
rect 1398 2106 1404 2107
rect 1822 2111 1828 2112
rect 1822 2107 1823 2111
rect 1827 2107 1828 2111
rect 1862 2108 1863 2112
rect 1867 2108 1868 2112
rect 2106 2111 2107 2115
rect 2111 2111 2112 2115
rect 2106 2110 2112 2111
rect 1862 2107 1868 2108
rect 1822 2106 1828 2107
rect 1318 2101 1324 2102
rect 1318 2097 1319 2101
rect 1323 2097 1324 2101
rect 1318 2096 1324 2097
rect 888 2087 890 2096
rect 1032 2087 1034 2096
rect 1176 2087 1178 2096
rect 1238 2095 1244 2096
rect 1238 2091 1239 2095
rect 1243 2091 1244 2095
rect 1238 2090 1244 2091
rect 1320 2087 1322 2096
rect 799 2086 803 2087
rect 799 2081 803 2082
rect 887 2086 891 2087
rect 887 2081 891 2082
rect 919 2086 923 2087
rect 919 2081 923 2082
rect 1031 2086 1035 2087
rect 1031 2081 1035 2082
rect 1039 2086 1043 2087
rect 1039 2081 1043 2082
rect 1159 2086 1163 2087
rect 1159 2081 1163 2082
rect 1175 2086 1179 2087
rect 1175 2081 1179 2082
rect 1279 2086 1283 2087
rect 1279 2081 1283 2082
rect 1319 2086 1323 2087
rect 1319 2081 1323 2082
rect 800 2076 802 2081
rect 920 2076 922 2081
rect 1040 2076 1042 2081
rect 1160 2076 1162 2081
rect 1280 2076 1282 2081
rect 798 2075 804 2076
rect 798 2071 799 2075
rect 803 2071 804 2075
rect 798 2070 804 2071
rect 918 2075 924 2076
rect 918 2071 919 2075
rect 923 2071 924 2075
rect 918 2070 924 2071
rect 1038 2075 1044 2076
rect 1038 2071 1039 2075
rect 1043 2071 1044 2075
rect 1038 2070 1044 2071
rect 1158 2075 1164 2076
rect 1158 2071 1159 2075
rect 1163 2071 1164 2075
rect 1158 2070 1164 2071
rect 1278 2075 1284 2076
rect 1278 2071 1279 2075
rect 1283 2071 1284 2075
rect 1278 2070 1284 2071
rect 766 2067 772 2068
rect 110 2065 116 2066
rect 110 2061 111 2065
rect 115 2061 116 2065
rect 766 2063 767 2067
rect 771 2063 772 2067
rect 766 2062 772 2063
rect 110 2060 116 2061
rect 1126 2051 1132 2052
rect 110 2048 116 2049
rect 110 2044 111 2048
rect 115 2044 116 2048
rect 1126 2047 1127 2051
rect 1131 2047 1132 2051
rect 1126 2046 1132 2047
rect 1226 2051 1232 2052
rect 1226 2047 1227 2051
rect 1231 2047 1232 2051
rect 1226 2046 1232 2047
rect 1346 2051 1352 2052
rect 1346 2047 1347 2051
rect 1351 2047 1352 2051
rect 1346 2046 1352 2047
rect 110 2043 116 2044
rect 112 2015 114 2043
rect 326 2035 332 2036
rect 326 2031 327 2035
rect 331 2031 332 2035
rect 326 2030 332 2031
rect 438 2035 444 2036
rect 438 2031 439 2035
rect 443 2031 444 2035
rect 438 2030 444 2031
rect 558 2035 564 2036
rect 558 2031 559 2035
rect 563 2031 564 2035
rect 558 2030 564 2031
rect 686 2035 692 2036
rect 686 2031 687 2035
rect 691 2031 692 2035
rect 686 2030 692 2031
rect 806 2035 812 2036
rect 806 2031 807 2035
rect 811 2031 812 2035
rect 806 2030 812 2031
rect 926 2035 932 2036
rect 926 2031 927 2035
rect 931 2031 932 2035
rect 926 2030 932 2031
rect 1046 2035 1052 2036
rect 1046 2031 1047 2035
rect 1051 2031 1052 2035
rect 1046 2030 1052 2031
rect 328 2015 330 2030
rect 440 2015 442 2030
rect 560 2015 562 2030
rect 688 2015 690 2030
rect 808 2015 810 2030
rect 928 2015 930 2030
rect 1048 2015 1050 2030
rect 111 2014 115 2015
rect 111 2009 115 2010
rect 183 2014 187 2015
rect 183 2009 187 2010
rect 295 2014 299 2015
rect 295 2009 299 2010
rect 327 2014 331 2015
rect 327 2009 331 2010
rect 415 2014 419 2015
rect 415 2009 419 2010
rect 439 2014 443 2015
rect 439 2009 443 2010
rect 535 2014 539 2015
rect 535 2009 539 2010
rect 559 2014 563 2015
rect 559 2009 563 2010
rect 655 2014 659 2015
rect 655 2009 659 2010
rect 687 2014 691 2015
rect 687 2009 691 2010
rect 775 2014 779 2015
rect 775 2009 779 2010
rect 807 2014 811 2015
rect 807 2009 811 2010
rect 895 2014 899 2015
rect 895 2009 899 2010
rect 927 2014 931 2015
rect 927 2009 931 2010
rect 1015 2014 1019 2015
rect 1015 2009 1019 2010
rect 1047 2014 1051 2015
rect 1047 2009 1051 2010
rect 112 1985 114 2009
rect 184 1998 186 2009
rect 238 2007 244 2008
rect 238 2003 239 2007
rect 243 2003 244 2007
rect 238 2002 244 2003
rect 182 1997 188 1998
rect 182 1993 183 1997
rect 187 1993 188 1997
rect 182 1992 188 1993
rect 110 1984 116 1985
rect 110 1980 111 1984
rect 115 1980 116 1984
rect 110 1979 116 1980
rect 110 1967 116 1968
rect 110 1963 111 1967
rect 115 1963 116 1967
rect 240 1965 242 2002
rect 296 1998 298 2009
rect 416 1998 418 2009
rect 536 1998 538 2009
rect 656 1998 658 2009
rect 776 1998 778 2009
rect 842 2007 848 2008
rect 842 2003 843 2007
rect 847 2003 848 2007
rect 842 2002 848 2003
rect 294 1997 300 1998
rect 294 1993 295 1997
rect 299 1993 300 1997
rect 294 1992 300 1993
rect 414 1997 420 1998
rect 414 1993 415 1997
rect 419 1993 420 1997
rect 414 1992 420 1993
rect 534 1997 540 1998
rect 534 1993 535 1997
rect 539 1993 540 1997
rect 534 1992 540 1993
rect 654 1997 660 1998
rect 654 1993 655 1997
rect 659 1993 660 1997
rect 654 1992 660 1993
rect 774 1997 780 1998
rect 774 1993 775 1997
rect 779 1993 780 1997
rect 774 1992 780 1993
rect 844 1980 846 2002
rect 896 1998 898 2009
rect 962 2007 968 2008
rect 962 2003 963 2007
rect 967 2003 968 2007
rect 962 2002 968 2003
rect 894 1997 900 1998
rect 894 1993 895 1997
rect 899 1993 900 1997
rect 894 1992 900 1993
rect 964 1980 966 2002
rect 1016 1998 1018 2009
rect 1128 2008 1130 2046
rect 1166 2035 1172 2036
rect 1166 2031 1167 2035
rect 1171 2031 1172 2035
rect 1166 2030 1172 2031
rect 1168 2015 1170 2030
rect 1228 2024 1230 2046
rect 1286 2035 1292 2036
rect 1286 2031 1287 2035
rect 1291 2031 1292 2035
rect 1286 2030 1292 2031
rect 1226 2023 1232 2024
rect 1226 2019 1227 2023
rect 1231 2019 1232 2023
rect 1226 2018 1232 2019
rect 1288 2015 1290 2030
rect 1348 2024 1350 2046
rect 1400 2024 1402 2106
rect 1462 2101 1468 2102
rect 1462 2097 1463 2101
rect 1467 2097 1468 2101
rect 1462 2096 1468 2097
rect 1614 2101 1620 2102
rect 1614 2097 1615 2101
rect 1619 2097 1620 2101
rect 1614 2096 1620 2097
rect 1464 2087 1466 2096
rect 1616 2087 1618 2096
rect 1824 2087 1826 2106
rect 1407 2086 1411 2087
rect 1407 2081 1411 2082
rect 1463 2086 1467 2087
rect 1463 2081 1467 2082
rect 1615 2086 1619 2087
rect 1615 2081 1619 2082
rect 1823 2086 1827 2087
rect 1823 2081 1827 2082
rect 1408 2076 1410 2081
rect 1406 2075 1412 2076
rect 1406 2071 1407 2075
rect 1411 2071 1412 2075
rect 1406 2070 1412 2071
rect 1824 2066 1826 2081
rect 1864 2079 1866 2107
rect 2030 2099 2036 2100
rect 2030 2095 2031 2099
rect 2035 2095 2036 2099
rect 2030 2094 2036 2095
rect 2032 2079 2034 2094
rect 2108 2088 2110 2110
rect 2174 2099 2180 2100
rect 2174 2095 2175 2099
rect 2179 2095 2180 2099
rect 2174 2094 2180 2095
rect 2106 2087 2112 2088
rect 2106 2083 2107 2087
rect 2111 2083 2112 2087
rect 2106 2082 2112 2083
rect 2176 2079 2178 2094
rect 2236 2088 2238 2174
rect 2326 2169 2332 2170
rect 2326 2165 2327 2169
rect 2331 2165 2332 2169
rect 2326 2164 2332 2165
rect 2510 2169 2516 2170
rect 2510 2165 2511 2169
rect 2515 2165 2516 2169
rect 2510 2164 2516 2165
rect 2702 2169 2708 2170
rect 2702 2165 2703 2169
rect 2707 2165 2708 2169
rect 2702 2164 2708 2165
rect 2328 2151 2330 2164
rect 2512 2151 2514 2164
rect 2704 2151 2706 2164
rect 2319 2150 2323 2151
rect 2319 2145 2323 2146
rect 2327 2150 2331 2151
rect 2327 2145 2331 2146
rect 2471 2150 2475 2151
rect 2471 2145 2475 2146
rect 2511 2150 2515 2151
rect 2511 2145 2515 2146
rect 2615 2150 2619 2151
rect 2615 2145 2619 2146
rect 2703 2150 2707 2151
rect 2703 2145 2707 2146
rect 2759 2150 2763 2151
rect 2759 2145 2763 2146
rect 2320 2140 2322 2145
rect 2472 2140 2474 2145
rect 2616 2140 2618 2145
rect 2760 2140 2762 2145
rect 2318 2139 2324 2140
rect 2318 2135 2319 2139
rect 2323 2135 2324 2139
rect 2318 2134 2324 2135
rect 2470 2139 2476 2140
rect 2470 2135 2471 2139
rect 2475 2135 2476 2139
rect 2470 2134 2476 2135
rect 2614 2139 2620 2140
rect 2614 2135 2615 2139
rect 2619 2135 2620 2139
rect 2614 2134 2620 2135
rect 2758 2139 2764 2140
rect 2758 2135 2759 2139
rect 2763 2135 2764 2139
rect 2758 2134 2764 2135
rect 2840 2132 2842 2214
rect 2904 2210 2906 2221
rect 3104 2210 3106 2221
rect 3112 2220 3114 2270
rect 3150 2259 3156 2260
rect 3150 2255 3151 2259
rect 3155 2255 3156 2259
rect 3150 2254 3156 2255
rect 3152 2232 3154 2254
rect 3166 2243 3172 2244
rect 3166 2239 3167 2243
rect 3171 2239 3172 2243
rect 3166 2238 3172 2239
rect 3150 2231 3156 2232
rect 3150 2227 3151 2231
rect 3155 2227 3156 2231
rect 3168 2227 3170 2238
rect 3184 2237 3186 2314
rect 3278 2309 3284 2310
rect 3278 2305 3279 2309
rect 3283 2305 3284 2309
rect 3278 2304 3284 2305
rect 3390 2309 3396 2310
rect 3390 2305 3391 2309
rect 3395 2305 3396 2309
rect 3390 2304 3396 2305
rect 3478 2309 3484 2310
rect 3478 2305 3479 2309
rect 3483 2305 3484 2309
rect 3478 2304 3484 2305
rect 3280 2295 3282 2304
rect 3392 2295 3394 2304
rect 3480 2295 3482 2304
rect 3576 2295 3578 2314
rect 3271 2294 3275 2295
rect 3271 2289 3275 2290
rect 3279 2294 3283 2295
rect 3279 2289 3283 2290
rect 3383 2294 3387 2295
rect 3383 2289 3387 2290
rect 3391 2294 3395 2295
rect 3391 2289 3395 2290
rect 3479 2294 3483 2295
rect 3479 2289 3483 2290
rect 3575 2294 3579 2295
rect 3575 2289 3579 2290
rect 3272 2284 3274 2289
rect 3384 2284 3386 2289
rect 3480 2284 3482 2289
rect 3270 2283 3276 2284
rect 3270 2279 3271 2283
rect 3275 2279 3276 2283
rect 3270 2278 3276 2279
rect 3382 2283 3388 2284
rect 3382 2279 3383 2283
rect 3387 2279 3388 2283
rect 3382 2278 3388 2279
rect 3478 2283 3484 2284
rect 3478 2279 3479 2283
rect 3483 2279 3484 2283
rect 3478 2278 3484 2279
rect 3576 2274 3578 2289
rect 3574 2273 3580 2274
rect 3574 2269 3575 2273
rect 3579 2269 3580 2273
rect 3574 2268 3580 2269
rect 3338 2259 3344 2260
rect 3338 2255 3339 2259
rect 3343 2255 3344 2259
rect 3338 2254 3344 2255
rect 3470 2259 3476 2260
rect 3470 2255 3471 2259
rect 3475 2255 3476 2259
rect 3470 2254 3476 2255
rect 3574 2256 3580 2257
rect 3278 2243 3284 2244
rect 3278 2239 3279 2243
rect 3283 2239 3284 2243
rect 3278 2238 3284 2239
rect 3183 2236 3187 2237
rect 3183 2231 3187 2232
rect 3280 2227 3282 2238
rect 3340 2232 3342 2254
rect 3390 2243 3396 2244
rect 3390 2239 3391 2243
rect 3395 2239 3396 2243
rect 3390 2238 3396 2239
rect 3338 2231 3344 2232
rect 3338 2227 3339 2231
rect 3343 2227 3344 2231
rect 3392 2227 3394 2238
rect 3150 2226 3156 2227
rect 3167 2226 3171 2227
rect 3167 2221 3171 2222
rect 3279 2226 3283 2227
rect 3279 2221 3283 2222
rect 3303 2226 3307 2227
rect 3338 2226 3344 2227
rect 3391 2226 3395 2227
rect 3303 2221 3307 2222
rect 3391 2221 3395 2222
rect 3110 2219 3116 2220
rect 3110 2215 3111 2219
rect 3115 2215 3116 2219
rect 3110 2214 3116 2215
rect 3304 2210 3306 2221
rect 3472 2220 3474 2254
rect 3574 2252 3575 2256
rect 3579 2252 3580 2256
rect 3574 2251 3580 2252
rect 3486 2243 3492 2244
rect 3486 2239 3487 2243
rect 3491 2239 3492 2243
rect 3486 2238 3492 2239
rect 3488 2227 3490 2238
rect 3576 2227 3578 2251
rect 3487 2226 3491 2227
rect 3487 2221 3491 2222
rect 3575 2226 3579 2227
rect 3575 2221 3579 2222
rect 3470 2219 3476 2220
rect 3470 2215 3471 2219
rect 3475 2215 3476 2219
rect 3470 2214 3476 2215
rect 3488 2210 3490 2221
rect 2902 2209 2908 2210
rect 2902 2205 2903 2209
rect 2907 2205 2908 2209
rect 2902 2204 2908 2205
rect 3102 2209 3108 2210
rect 3102 2205 3103 2209
rect 3107 2205 3108 2209
rect 3102 2204 3108 2205
rect 3302 2209 3308 2210
rect 3302 2205 3303 2209
rect 3307 2205 3308 2209
rect 3302 2204 3308 2205
rect 3486 2209 3492 2210
rect 3486 2205 3487 2209
rect 3491 2205 3492 2209
rect 3486 2204 3492 2205
rect 3576 2197 3578 2221
rect 3574 2196 3580 2197
rect 3574 2192 3575 2196
rect 3579 2192 3580 2196
rect 3574 2191 3580 2192
rect 3574 2179 3580 2180
rect 3574 2175 3575 2179
rect 3579 2175 3580 2179
rect 3574 2174 3580 2175
rect 2894 2169 2900 2170
rect 2894 2165 2895 2169
rect 2899 2165 2900 2169
rect 2894 2164 2900 2165
rect 3094 2169 3100 2170
rect 3094 2165 3095 2169
rect 3099 2165 3100 2169
rect 3094 2164 3100 2165
rect 3294 2169 3300 2170
rect 3294 2165 3295 2169
rect 3299 2165 3300 2169
rect 3294 2164 3300 2165
rect 3478 2169 3484 2170
rect 3478 2165 3479 2169
rect 3483 2165 3484 2169
rect 3478 2164 3484 2165
rect 2896 2151 2898 2164
rect 3096 2151 3098 2164
rect 3296 2151 3298 2164
rect 3480 2151 3482 2164
rect 3576 2151 3578 2174
rect 2895 2150 2899 2151
rect 2895 2145 2899 2146
rect 3023 2150 3027 2151
rect 3023 2145 3027 2146
rect 3095 2150 3099 2151
rect 3095 2145 3099 2146
rect 3143 2150 3147 2151
rect 3143 2145 3147 2146
rect 3263 2150 3267 2151
rect 3263 2145 3267 2146
rect 3295 2150 3299 2151
rect 3295 2145 3299 2146
rect 3383 2150 3387 2151
rect 3383 2145 3387 2146
rect 3479 2150 3483 2151
rect 3479 2145 3483 2146
rect 3575 2150 3579 2151
rect 3575 2145 3579 2146
rect 2896 2140 2898 2145
rect 3024 2140 3026 2145
rect 3144 2140 3146 2145
rect 3264 2140 3266 2145
rect 3384 2140 3386 2145
rect 3480 2140 3482 2145
rect 2894 2139 2900 2140
rect 2894 2135 2895 2139
rect 2899 2135 2900 2139
rect 2894 2134 2900 2135
rect 3022 2139 3028 2140
rect 3022 2135 3023 2139
rect 3027 2135 3028 2139
rect 3022 2134 3028 2135
rect 3142 2139 3148 2140
rect 3142 2135 3143 2139
rect 3147 2135 3148 2139
rect 3142 2134 3148 2135
rect 3262 2139 3268 2140
rect 3262 2135 3263 2139
rect 3267 2135 3268 2139
rect 3262 2134 3268 2135
rect 3382 2139 3388 2140
rect 3382 2135 3383 2139
rect 3387 2135 3388 2139
rect 3382 2134 3388 2135
rect 3478 2139 3484 2140
rect 3478 2135 3479 2139
rect 3483 2135 3484 2139
rect 3478 2134 3484 2135
rect 2838 2131 2844 2132
rect 2838 2127 2839 2131
rect 2843 2127 2844 2131
rect 2838 2126 2844 2127
rect 3450 2131 3456 2132
rect 3450 2127 3451 2131
rect 3455 2127 3456 2131
rect 3576 2130 3578 2145
rect 3450 2126 3456 2127
rect 3574 2129 3580 2130
rect 2826 2115 2832 2116
rect 2826 2111 2827 2115
rect 2831 2111 2832 2115
rect 2826 2110 2832 2111
rect 2962 2115 2968 2116
rect 2962 2111 2963 2115
rect 2967 2111 2968 2115
rect 2962 2110 2968 2111
rect 3090 2115 3096 2116
rect 3090 2111 3091 2115
rect 3095 2111 3096 2115
rect 3090 2110 3096 2111
rect 3210 2115 3216 2116
rect 3210 2111 3211 2115
rect 3215 2111 3216 2115
rect 3210 2110 3216 2111
rect 2326 2099 2332 2100
rect 2326 2095 2327 2099
rect 2331 2095 2332 2099
rect 2326 2094 2332 2095
rect 2478 2099 2484 2100
rect 2478 2095 2479 2099
rect 2483 2095 2484 2099
rect 2478 2094 2484 2095
rect 2622 2099 2628 2100
rect 2622 2095 2623 2099
rect 2627 2095 2628 2099
rect 2622 2094 2628 2095
rect 2766 2099 2772 2100
rect 2766 2095 2767 2099
rect 2771 2095 2772 2099
rect 2766 2094 2772 2095
rect 2234 2087 2240 2088
rect 2234 2083 2235 2087
rect 2239 2083 2240 2087
rect 2234 2082 2240 2083
rect 2302 2087 2308 2088
rect 2302 2083 2303 2087
rect 2307 2083 2308 2087
rect 2302 2082 2308 2083
rect 1863 2078 1867 2079
rect 1863 2073 1867 2074
rect 1983 2078 1987 2079
rect 1983 2073 1987 2074
rect 2031 2078 2035 2079
rect 2031 2073 2035 2074
rect 2143 2078 2147 2079
rect 2143 2073 2147 2074
rect 2175 2078 2179 2079
rect 2175 2073 2179 2074
rect 1822 2065 1828 2066
rect 1822 2061 1823 2065
rect 1827 2061 1828 2065
rect 1822 2060 1828 2061
rect 1864 2049 1866 2073
rect 1984 2062 1986 2073
rect 2144 2062 2146 2073
rect 1982 2061 1988 2062
rect 1982 2057 1983 2061
rect 1987 2057 1988 2061
rect 1982 2056 1988 2057
rect 2142 2061 2148 2062
rect 2142 2057 2143 2061
rect 2147 2057 2148 2061
rect 2142 2056 2148 2057
rect 1822 2048 1828 2049
rect 1822 2044 1823 2048
rect 1827 2044 1828 2048
rect 1822 2043 1828 2044
rect 1862 2048 1868 2049
rect 1862 2044 1863 2048
rect 1867 2044 1868 2048
rect 2304 2044 2306 2082
rect 2328 2079 2330 2094
rect 2480 2079 2482 2094
rect 2624 2079 2626 2094
rect 2768 2079 2770 2094
rect 2311 2078 2315 2079
rect 2311 2073 2315 2074
rect 2327 2078 2331 2079
rect 2327 2073 2331 2074
rect 2471 2078 2475 2079
rect 2471 2073 2475 2074
rect 2479 2078 2483 2079
rect 2479 2073 2483 2074
rect 2623 2078 2627 2079
rect 2623 2073 2627 2074
rect 2631 2078 2635 2079
rect 2631 2073 2635 2074
rect 2767 2078 2771 2079
rect 2767 2073 2771 2074
rect 2775 2078 2779 2079
rect 2775 2073 2779 2074
rect 2312 2062 2314 2073
rect 2472 2062 2474 2073
rect 2610 2071 2616 2072
rect 2610 2067 2611 2071
rect 2615 2067 2616 2071
rect 2610 2066 2616 2067
rect 2310 2061 2316 2062
rect 2310 2057 2311 2061
rect 2315 2057 2316 2061
rect 2310 2056 2316 2057
rect 2470 2061 2476 2062
rect 2470 2057 2471 2061
rect 2475 2057 2476 2061
rect 2470 2056 2476 2057
rect 1862 2043 1868 2044
rect 2302 2043 2308 2044
rect 1414 2035 1420 2036
rect 1414 2031 1415 2035
rect 1419 2031 1420 2035
rect 1414 2030 1420 2031
rect 1346 2023 1352 2024
rect 1346 2019 1347 2023
rect 1351 2019 1352 2023
rect 1346 2018 1352 2019
rect 1398 2023 1404 2024
rect 1398 2019 1399 2023
rect 1403 2019 1404 2023
rect 1398 2018 1404 2019
rect 1416 2015 1418 2030
rect 1824 2015 1826 2043
rect 2302 2039 2303 2043
rect 2307 2039 2308 2043
rect 2302 2038 2308 2039
rect 1862 2031 1868 2032
rect 1862 2027 1863 2031
rect 1867 2027 1868 2031
rect 1862 2026 1868 2027
rect 1135 2014 1139 2015
rect 1135 2009 1139 2010
rect 1167 2014 1171 2015
rect 1167 2009 1171 2010
rect 1255 2014 1259 2015
rect 1255 2009 1259 2010
rect 1287 2014 1291 2015
rect 1287 2009 1291 2010
rect 1415 2014 1419 2015
rect 1415 2009 1419 2010
rect 1823 2014 1827 2015
rect 1864 2011 1866 2026
rect 1974 2021 1980 2022
rect 1974 2017 1975 2021
rect 1979 2017 1980 2021
rect 1974 2016 1980 2017
rect 2134 2021 2140 2022
rect 2134 2017 2135 2021
rect 2139 2017 2140 2021
rect 2134 2016 2140 2017
rect 2302 2021 2308 2022
rect 2302 2017 2303 2021
rect 2307 2017 2308 2021
rect 2302 2016 2308 2017
rect 2462 2021 2468 2022
rect 2462 2017 2463 2021
rect 2467 2017 2468 2021
rect 2462 2016 2468 2017
rect 1976 2011 1978 2016
rect 2136 2011 2138 2016
rect 2304 2011 2306 2016
rect 2464 2011 2466 2016
rect 1823 2009 1827 2010
rect 1863 2010 1867 2011
rect 1118 2007 1124 2008
rect 1118 2003 1119 2007
rect 1123 2003 1124 2007
rect 1118 2002 1124 2003
rect 1126 2007 1132 2008
rect 1126 2003 1127 2007
rect 1131 2003 1132 2007
rect 1126 2002 1132 2003
rect 1014 1997 1020 1998
rect 1014 1993 1015 1997
rect 1019 1993 1020 1997
rect 1014 1992 1020 1993
rect 842 1979 848 1980
rect 842 1975 843 1979
rect 847 1975 848 1979
rect 842 1974 848 1975
rect 962 1979 968 1980
rect 962 1975 963 1979
rect 967 1975 968 1979
rect 962 1974 968 1975
rect 110 1962 116 1963
rect 239 1964 243 1965
rect 112 1943 114 1962
rect 239 1959 243 1960
rect 563 1964 567 1965
rect 563 1959 567 1960
rect 174 1957 180 1958
rect 174 1953 175 1957
rect 179 1953 180 1957
rect 174 1952 180 1953
rect 286 1957 292 1958
rect 286 1953 287 1957
rect 291 1953 292 1957
rect 286 1952 292 1953
rect 406 1957 412 1958
rect 406 1953 407 1957
rect 411 1953 412 1957
rect 406 1952 412 1953
rect 526 1957 532 1958
rect 526 1953 527 1957
rect 531 1953 532 1957
rect 526 1952 532 1953
rect 176 1943 178 1952
rect 288 1943 290 1952
rect 408 1943 410 1952
rect 528 1943 530 1952
rect 111 1942 115 1943
rect 111 1937 115 1938
rect 135 1942 139 1943
rect 135 1937 139 1938
rect 175 1942 179 1943
rect 175 1937 179 1938
rect 223 1942 227 1943
rect 223 1937 227 1938
rect 287 1942 291 1943
rect 287 1937 291 1938
rect 351 1942 355 1943
rect 351 1937 355 1938
rect 407 1942 411 1943
rect 407 1937 411 1938
rect 495 1942 499 1943
rect 495 1937 499 1938
rect 527 1942 531 1943
rect 527 1937 531 1938
rect 112 1922 114 1937
rect 136 1932 138 1937
rect 224 1932 226 1937
rect 352 1932 354 1937
rect 496 1932 498 1937
rect 134 1931 140 1932
rect 134 1927 135 1931
rect 139 1927 140 1931
rect 134 1926 140 1927
rect 222 1931 228 1932
rect 222 1927 223 1931
rect 227 1927 228 1931
rect 222 1926 228 1927
rect 350 1931 356 1932
rect 350 1927 351 1931
rect 355 1927 356 1931
rect 350 1926 356 1927
rect 494 1931 500 1932
rect 494 1927 495 1931
rect 499 1927 500 1931
rect 494 1926 500 1927
rect 564 1924 566 1959
rect 646 1957 652 1958
rect 646 1953 647 1957
rect 651 1953 652 1957
rect 646 1952 652 1953
rect 766 1957 772 1958
rect 766 1953 767 1957
rect 771 1953 772 1957
rect 766 1952 772 1953
rect 886 1957 892 1958
rect 886 1953 887 1957
rect 891 1953 892 1957
rect 886 1952 892 1953
rect 1006 1957 1012 1958
rect 1006 1953 1007 1957
rect 1011 1953 1012 1957
rect 1006 1952 1012 1953
rect 1120 1952 1122 2002
rect 1136 1998 1138 2009
rect 1256 1998 1258 2009
rect 1134 1997 1140 1998
rect 1134 1993 1135 1997
rect 1139 1993 1140 1997
rect 1134 1992 1140 1993
rect 1254 1997 1260 1998
rect 1254 1993 1255 1997
rect 1259 1993 1260 1997
rect 1254 1992 1260 1993
rect 1824 1985 1826 2009
rect 1863 2005 1867 2006
rect 1887 2010 1891 2011
rect 1887 2005 1891 2006
rect 1975 2010 1979 2011
rect 1975 2005 1979 2006
rect 2031 2010 2035 2011
rect 2031 2005 2035 2006
rect 2135 2010 2139 2011
rect 2135 2005 2139 2006
rect 2199 2010 2203 2011
rect 2199 2005 2203 2006
rect 2303 2010 2307 2011
rect 2303 2005 2307 2006
rect 2375 2010 2379 2011
rect 2375 2005 2379 2006
rect 2463 2010 2467 2011
rect 2463 2005 2467 2006
rect 2543 2010 2547 2011
rect 2543 2005 2547 2006
rect 1864 1990 1866 2005
rect 1888 2000 1890 2005
rect 2032 2000 2034 2005
rect 2200 2000 2202 2005
rect 2376 2000 2378 2005
rect 2544 2000 2546 2005
rect 1886 1999 1892 2000
rect 1886 1995 1887 1999
rect 1891 1995 1892 1999
rect 1886 1994 1892 1995
rect 2030 1999 2036 2000
rect 2030 1995 2031 1999
rect 2035 1995 2036 1999
rect 2030 1994 2036 1995
rect 2198 1999 2204 2000
rect 2198 1995 2199 1999
rect 2203 1995 2204 1999
rect 2198 1994 2204 1995
rect 2374 1999 2380 2000
rect 2374 1995 2375 1999
rect 2379 1995 2380 1999
rect 2374 1994 2380 1995
rect 2542 1999 2548 2000
rect 2542 1995 2543 1999
rect 2547 1995 2548 1999
rect 2542 1994 2548 1995
rect 2612 1992 2614 2066
rect 2632 2062 2634 2073
rect 2776 2062 2778 2073
rect 2828 2072 2830 2110
rect 2902 2099 2908 2100
rect 2902 2095 2903 2099
rect 2907 2095 2908 2099
rect 2902 2094 2908 2095
rect 2904 2079 2906 2094
rect 2964 2088 2966 2110
rect 3030 2099 3036 2100
rect 3030 2095 3031 2099
rect 3035 2095 3036 2099
rect 3030 2094 3036 2095
rect 2962 2087 2968 2088
rect 2962 2083 2963 2087
rect 2967 2083 2968 2087
rect 2962 2082 2968 2083
rect 3032 2079 3034 2094
rect 3092 2088 3094 2110
rect 3150 2099 3156 2100
rect 3150 2095 3151 2099
rect 3155 2095 3156 2099
rect 3150 2094 3156 2095
rect 3090 2087 3096 2088
rect 3090 2083 3091 2087
rect 3095 2083 3096 2087
rect 3090 2082 3096 2083
rect 3152 2079 3154 2094
rect 3212 2088 3214 2110
rect 3270 2099 3276 2100
rect 3270 2095 3271 2099
rect 3275 2095 3276 2099
rect 3270 2094 3276 2095
rect 3390 2099 3396 2100
rect 3390 2095 3391 2099
rect 3395 2095 3396 2099
rect 3390 2094 3396 2095
rect 3210 2087 3216 2088
rect 3210 2083 3211 2087
rect 3215 2083 3216 2087
rect 3210 2082 3216 2083
rect 3272 2079 3274 2094
rect 3392 2079 3394 2094
rect 3452 2088 3454 2126
rect 3574 2125 3575 2129
rect 3579 2125 3580 2129
rect 3574 2124 3580 2125
rect 3470 2115 3476 2116
rect 3470 2111 3471 2115
rect 3475 2111 3476 2115
rect 3470 2110 3476 2111
rect 3574 2112 3580 2113
rect 3450 2087 3456 2088
rect 3450 2083 3451 2087
rect 3455 2083 3456 2087
rect 3450 2082 3456 2083
rect 2903 2078 2907 2079
rect 2903 2073 2907 2074
rect 2911 2078 2915 2079
rect 2911 2073 2915 2074
rect 3031 2078 3035 2079
rect 3031 2073 3035 2074
rect 3039 2078 3043 2079
rect 3039 2073 3043 2074
rect 3151 2078 3155 2079
rect 3151 2073 3155 2074
rect 3159 2078 3163 2079
rect 3159 2073 3163 2074
rect 3271 2078 3275 2079
rect 3271 2073 3275 2074
rect 3279 2078 3283 2079
rect 3279 2073 3283 2074
rect 3391 2078 3395 2079
rect 3391 2073 3395 2074
rect 2826 2071 2832 2072
rect 2826 2067 2827 2071
rect 2831 2067 2832 2071
rect 2826 2066 2832 2067
rect 2912 2062 2914 2073
rect 3040 2062 3042 2073
rect 3160 2062 3162 2073
rect 3280 2062 3282 2073
rect 3346 2071 3352 2072
rect 3346 2067 3347 2071
rect 3351 2067 3352 2071
rect 3346 2066 3352 2067
rect 2630 2061 2636 2062
rect 2630 2057 2631 2061
rect 2635 2057 2636 2061
rect 2630 2056 2636 2057
rect 2774 2061 2780 2062
rect 2774 2057 2775 2061
rect 2779 2057 2780 2061
rect 2774 2056 2780 2057
rect 2910 2061 2916 2062
rect 2910 2057 2911 2061
rect 2915 2057 2916 2061
rect 2910 2056 2916 2057
rect 3038 2061 3044 2062
rect 3038 2057 3039 2061
rect 3043 2057 3044 2061
rect 3038 2056 3044 2057
rect 3158 2061 3164 2062
rect 3158 2057 3159 2061
rect 3163 2057 3164 2061
rect 3158 2056 3164 2057
rect 3278 2061 3284 2062
rect 3278 2057 3279 2061
rect 3283 2057 3284 2061
rect 3278 2056 3284 2057
rect 3348 2044 3350 2066
rect 3392 2062 3394 2073
rect 3472 2072 3474 2110
rect 3574 2108 3575 2112
rect 3579 2108 3580 2112
rect 3574 2107 3580 2108
rect 3486 2099 3492 2100
rect 3486 2095 3487 2099
rect 3491 2095 3492 2099
rect 3486 2094 3492 2095
rect 3488 2079 3490 2094
rect 3576 2079 3578 2107
rect 3487 2078 3491 2079
rect 3487 2073 3491 2074
rect 3575 2078 3579 2079
rect 3575 2073 3579 2074
rect 3458 2071 3464 2072
rect 3458 2067 3459 2071
rect 3463 2067 3464 2071
rect 3458 2066 3464 2067
rect 3470 2071 3476 2072
rect 3470 2067 3471 2071
rect 3475 2067 3476 2071
rect 3470 2066 3476 2067
rect 3390 2061 3396 2062
rect 3390 2057 3391 2061
rect 3395 2057 3396 2061
rect 3390 2056 3396 2057
rect 3460 2044 3462 2066
rect 3488 2062 3490 2073
rect 3486 2061 3492 2062
rect 3486 2057 3487 2061
rect 3491 2057 3492 2061
rect 3486 2056 3492 2057
rect 3576 2049 3578 2073
rect 3574 2048 3580 2049
rect 3574 2044 3575 2048
rect 3579 2044 3580 2048
rect 3346 2043 3352 2044
rect 3346 2039 3347 2043
rect 3351 2039 3352 2043
rect 3346 2038 3352 2039
rect 3458 2043 3464 2044
rect 3574 2043 3580 2044
rect 3458 2039 3459 2043
rect 3463 2039 3464 2043
rect 3458 2038 3464 2039
rect 3574 2031 3580 2032
rect 3574 2027 3575 2031
rect 3579 2027 3580 2031
rect 3574 2026 3580 2027
rect 2622 2021 2628 2022
rect 2622 2017 2623 2021
rect 2627 2017 2628 2021
rect 2622 2016 2628 2017
rect 2766 2021 2772 2022
rect 2766 2017 2767 2021
rect 2771 2017 2772 2021
rect 2766 2016 2772 2017
rect 2902 2021 2908 2022
rect 2902 2017 2903 2021
rect 2907 2017 2908 2021
rect 2902 2016 2908 2017
rect 3030 2021 3036 2022
rect 3030 2017 3031 2021
rect 3035 2017 3036 2021
rect 3030 2016 3036 2017
rect 3150 2021 3156 2022
rect 3150 2017 3151 2021
rect 3155 2017 3156 2021
rect 3150 2016 3156 2017
rect 3270 2021 3276 2022
rect 3270 2017 3271 2021
rect 3275 2017 3276 2021
rect 3270 2016 3276 2017
rect 3382 2021 3388 2022
rect 3382 2017 3383 2021
rect 3387 2017 3388 2021
rect 3382 2016 3388 2017
rect 3478 2021 3484 2022
rect 3478 2017 3479 2021
rect 3483 2017 3484 2021
rect 3478 2016 3484 2017
rect 2624 2011 2626 2016
rect 2768 2011 2770 2016
rect 2904 2011 2906 2016
rect 3032 2011 3034 2016
rect 3152 2011 3154 2016
rect 3272 2011 3274 2016
rect 3384 2011 3386 2016
rect 3480 2011 3482 2016
rect 3576 2011 3578 2026
rect 2623 2010 2627 2011
rect 2623 2005 2627 2006
rect 2711 2010 2715 2011
rect 2711 2005 2715 2006
rect 2767 2010 2771 2011
rect 2767 2005 2771 2006
rect 2871 2010 2875 2011
rect 2871 2005 2875 2006
rect 2903 2010 2907 2011
rect 2903 2005 2907 2006
rect 3031 2010 3035 2011
rect 3031 2005 3035 2006
rect 3039 2010 3043 2011
rect 3039 2005 3043 2006
rect 3151 2010 3155 2011
rect 3151 2005 3155 2006
rect 3207 2010 3211 2011
rect 3207 2005 3211 2006
rect 3271 2010 3275 2011
rect 3271 2005 3275 2006
rect 3383 2010 3387 2011
rect 3383 2005 3387 2006
rect 3479 2010 3483 2011
rect 3479 2005 3483 2006
rect 3575 2010 3579 2011
rect 3575 2005 3579 2006
rect 2712 2000 2714 2005
rect 2872 2000 2874 2005
rect 3040 2000 3042 2005
rect 3208 2000 3210 2005
rect 2710 1999 2716 2000
rect 2710 1995 2711 1999
rect 2715 1995 2716 1999
rect 2710 1994 2716 1995
rect 2870 1999 2876 2000
rect 2870 1995 2871 1999
rect 2875 1995 2876 1999
rect 2870 1994 2876 1995
rect 3038 1999 3044 2000
rect 3038 1995 3039 1999
rect 3043 1995 3044 1999
rect 3038 1994 3044 1995
rect 3206 1999 3212 2000
rect 3206 1995 3207 1999
rect 3211 1995 3212 1999
rect 3206 1994 3212 1995
rect 2610 1991 2616 1992
rect 1862 1989 1868 1990
rect 1862 1985 1863 1989
rect 1867 1985 1868 1989
rect 2610 1987 2611 1991
rect 2615 1987 2616 1991
rect 3576 1990 3578 2005
rect 2610 1986 2616 1987
rect 3574 1989 3580 1990
rect 1822 1984 1828 1985
rect 1862 1984 1868 1985
rect 3574 1985 3575 1989
rect 3579 1985 3580 1989
rect 3574 1984 3580 1985
rect 1822 1980 1823 1984
rect 1827 1980 1828 1984
rect 1822 1979 1828 1980
rect 1982 1975 1988 1976
rect 1862 1972 1868 1973
rect 1862 1968 1863 1972
rect 1867 1968 1868 1972
rect 1982 1971 1983 1975
rect 1987 1971 1988 1975
rect 1982 1970 1988 1971
rect 1990 1975 1996 1976
rect 1990 1971 1991 1975
rect 1995 1971 1996 1975
rect 1990 1970 1996 1971
rect 2098 1975 2104 1976
rect 2098 1971 2099 1975
rect 2103 1971 2104 1975
rect 2098 1970 2104 1971
rect 2998 1975 3004 1976
rect 2998 1971 2999 1975
rect 3003 1971 3004 1975
rect 2998 1970 3004 1971
rect 3150 1975 3156 1976
rect 3150 1971 3151 1975
rect 3155 1971 3156 1975
rect 3150 1970 3156 1971
rect 3158 1975 3164 1976
rect 3158 1971 3159 1975
rect 3163 1971 3164 1975
rect 3158 1970 3164 1971
rect 3574 1972 3580 1973
rect 1822 1967 1828 1968
rect 1862 1967 1868 1968
rect 1822 1963 1823 1967
rect 1827 1963 1828 1967
rect 1822 1962 1828 1963
rect 1126 1957 1132 1958
rect 1126 1953 1127 1957
rect 1131 1953 1132 1957
rect 1126 1952 1132 1953
rect 1246 1957 1252 1958
rect 1246 1953 1247 1957
rect 1251 1953 1252 1957
rect 1246 1952 1252 1953
rect 648 1943 650 1952
rect 768 1943 770 1952
rect 888 1943 890 1952
rect 1008 1943 1010 1952
rect 1118 1951 1124 1952
rect 1118 1947 1119 1951
rect 1123 1947 1124 1951
rect 1118 1946 1124 1947
rect 1128 1943 1130 1952
rect 1248 1943 1250 1952
rect 1824 1943 1826 1962
rect 647 1942 651 1943
rect 647 1937 651 1938
rect 655 1942 659 1943
rect 655 1937 659 1938
rect 767 1942 771 1943
rect 767 1937 771 1938
rect 839 1942 843 1943
rect 839 1937 843 1938
rect 887 1942 891 1943
rect 887 1937 891 1938
rect 1007 1942 1011 1943
rect 1007 1937 1011 1938
rect 1039 1942 1043 1943
rect 1039 1937 1043 1938
rect 1127 1942 1131 1943
rect 1127 1937 1131 1938
rect 1247 1942 1251 1943
rect 1247 1937 1251 1938
rect 1463 1942 1467 1943
rect 1463 1937 1467 1938
rect 1823 1942 1827 1943
rect 1823 1937 1827 1938
rect 656 1932 658 1937
rect 840 1932 842 1937
rect 1040 1932 1042 1937
rect 1248 1932 1250 1937
rect 1464 1932 1466 1937
rect 654 1931 660 1932
rect 654 1927 655 1931
rect 659 1927 660 1931
rect 654 1926 660 1927
rect 838 1931 844 1932
rect 838 1927 839 1931
rect 843 1927 844 1931
rect 838 1926 844 1927
rect 1038 1931 1044 1932
rect 1038 1927 1039 1931
rect 1043 1927 1044 1931
rect 1038 1926 1044 1927
rect 1246 1931 1252 1932
rect 1246 1927 1247 1931
rect 1251 1927 1252 1931
rect 1246 1926 1252 1927
rect 1462 1931 1468 1932
rect 1462 1927 1463 1931
rect 1467 1927 1468 1931
rect 1462 1926 1468 1927
rect 562 1923 568 1924
rect 110 1921 116 1922
rect 110 1917 111 1921
rect 115 1917 116 1921
rect 562 1919 563 1923
rect 567 1919 568 1923
rect 562 1918 568 1919
rect 1158 1923 1164 1924
rect 1158 1919 1159 1923
rect 1163 1919 1164 1923
rect 1824 1922 1826 1937
rect 1864 1935 1866 1967
rect 1894 1959 1900 1960
rect 1894 1955 1895 1959
rect 1899 1955 1900 1959
rect 1894 1954 1900 1955
rect 1896 1935 1898 1954
rect 1863 1934 1867 1935
rect 1863 1929 1867 1930
rect 1895 1934 1899 1935
rect 1895 1929 1899 1930
rect 1158 1918 1164 1919
rect 1822 1921 1828 1922
rect 110 1916 116 1917
rect 110 1904 116 1905
rect 110 1900 111 1904
rect 115 1900 116 1904
rect 110 1899 116 1900
rect 112 1867 114 1899
rect 142 1891 148 1892
rect 142 1887 143 1891
rect 147 1887 148 1891
rect 142 1886 148 1887
rect 230 1891 236 1892
rect 230 1887 231 1891
rect 235 1887 236 1891
rect 230 1886 236 1887
rect 358 1891 364 1892
rect 358 1887 359 1891
rect 363 1887 364 1891
rect 358 1886 364 1887
rect 502 1891 508 1892
rect 502 1887 503 1891
rect 507 1887 508 1891
rect 502 1886 508 1887
rect 662 1891 668 1892
rect 662 1887 663 1891
rect 667 1887 668 1891
rect 662 1886 668 1887
rect 846 1891 852 1892
rect 846 1887 847 1891
rect 851 1887 852 1891
rect 846 1886 852 1887
rect 1046 1891 1052 1892
rect 1046 1887 1047 1891
rect 1051 1887 1052 1891
rect 1046 1886 1052 1887
rect 134 1879 140 1880
rect 134 1875 135 1879
rect 139 1875 140 1879
rect 134 1874 140 1875
rect 111 1866 115 1867
rect 111 1861 115 1862
rect 112 1837 114 1861
rect 110 1836 116 1837
rect 110 1832 111 1836
rect 115 1832 116 1836
rect 136 1832 138 1874
rect 144 1867 146 1886
rect 232 1867 234 1886
rect 360 1867 362 1886
rect 504 1867 506 1886
rect 664 1867 666 1886
rect 848 1867 850 1886
rect 951 1884 955 1885
rect 951 1879 955 1880
rect 143 1866 147 1867
rect 143 1861 147 1862
rect 231 1866 235 1867
rect 231 1861 235 1862
rect 271 1866 275 1867
rect 271 1861 275 1862
rect 359 1866 363 1867
rect 359 1861 363 1862
rect 415 1866 419 1867
rect 415 1861 419 1862
rect 503 1866 507 1867
rect 503 1861 507 1862
rect 559 1866 563 1867
rect 559 1861 563 1862
rect 663 1866 667 1867
rect 663 1861 667 1862
rect 695 1866 699 1867
rect 695 1861 699 1862
rect 823 1866 827 1867
rect 823 1861 827 1862
rect 847 1866 851 1867
rect 847 1861 851 1862
rect 943 1866 947 1867
rect 943 1861 947 1862
rect 144 1850 146 1861
rect 210 1859 216 1860
rect 210 1855 211 1859
rect 215 1855 216 1859
rect 210 1854 216 1855
rect 142 1849 148 1850
rect 142 1845 143 1849
rect 147 1845 148 1849
rect 142 1844 148 1845
rect 212 1832 214 1854
rect 272 1850 274 1861
rect 338 1859 344 1860
rect 338 1855 339 1859
rect 343 1855 344 1859
rect 338 1854 344 1855
rect 370 1859 376 1860
rect 370 1855 371 1859
rect 375 1855 376 1859
rect 370 1854 376 1855
rect 270 1849 276 1850
rect 270 1845 271 1849
rect 275 1845 276 1849
rect 270 1844 276 1845
rect 340 1832 342 1854
rect 110 1831 116 1832
rect 134 1831 140 1832
rect 134 1827 135 1831
rect 139 1827 140 1831
rect 134 1826 140 1827
rect 210 1831 216 1832
rect 210 1827 211 1831
rect 215 1827 216 1831
rect 210 1826 216 1827
rect 338 1831 344 1832
rect 338 1827 339 1831
rect 343 1827 344 1831
rect 338 1826 344 1827
rect 110 1819 116 1820
rect 110 1815 111 1819
rect 115 1815 116 1819
rect 110 1814 116 1815
rect 112 1787 114 1814
rect 134 1809 140 1810
rect 134 1805 135 1809
rect 139 1805 140 1809
rect 134 1804 140 1805
rect 262 1809 268 1810
rect 262 1805 263 1809
rect 267 1805 268 1809
rect 262 1804 268 1805
rect 136 1787 138 1804
rect 264 1787 266 1804
rect 111 1786 115 1787
rect 111 1781 115 1782
rect 135 1786 139 1787
rect 135 1781 139 1782
rect 263 1786 267 1787
rect 263 1781 267 1782
rect 303 1786 307 1787
rect 303 1781 307 1782
rect 112 1766 114 1781
rect 136 1776 138 1781
rect 304 1776 306 1781
rect 134 1775 140 1776
rect 134 1771 135 1775
rect 139 1771 140 1775
rect 134 1770 140 1771
rect 302 1775 308 1776
rect 302 1771 303 1775
rect 307 1771 308 1775
rect 302 1770 308 1771
rect 372 1768 374 1854
rect 416 1850 418 1861
rect 560 1850 562 1861
rect 696 1850 698 1861
rect 762 1859 768 1860
rect 762 1855 763 1859
rect 767 1855 768 1859
rect 762 1854 768 1855
rect 414 1849 420 1850
rect 414 1845 415 1849
rect 419 1845 420 1849
rect 414 1844 420 1845
rect 558 1849 564 1850
rect 558 1845 559 1849
rect 563 1845 564 1849
rect 558 1844 564 1845
rect 694 1849 700 1850
rect 694 1845 695 1849
rect 699 1845 700 1849
rect 694 1844 700 1845
rect 764 1832 766 1854
rect 824 1850 826 1861
rect 890 1859 896 1860
rect 890 1855 891 1859
rect 895 1855 896 1859
rect 890 1854 896 1855
rect 822 1849 828 1850
rect 822 1845 823 1849
rect 827 1845 828 1849
rect 822 1844 828 1845
rect 892 1832 894 1854
rect 944 1850 946 1861
rect 952 1860 954 1879
rect 1048 1867 1050 1886
rect 1160 1885 1162 1918
rect 1822 1917 1823 1921
rect 1827 1917 1828 1921
rect 1822 1916 1828 1917
rect 1864 1905 1866 1929
rect 1896 1918 1898 1929
rect 1984 1928 1986 1970
rect 1992 1948 1994 1970
rect 2038 1959 2044 1960
rect 2038 1955 2039 1959
rect 2043 1955 2044 1959
rect 2038 1954 2044 1955
rect 1990 1947 1996 1948
rect 1990 1943 1991 1947
rect 1995 1943 1996 1947
rect 1990 1942 1996 1943
rect 2040 1935 2042 1954
rect 2100 1948 2102 1970
rect 2206 1959 2212 1960
rect 2206 1955 2207 1959
rect 2211 1955 2212 1959
rect 2206 1954 2212 1955
rect 2382 1959 2388 1960
rect 2382 1955 2383 1959
rect 2387 1955 2388 1959
rect 2382 1954 2388 1955
rect 2550 1959 2556 1960
rect 2550 1955 2551 1959
rect 2555 1955 2556 1959
rect 2550 1954 2556 1955
rect 2718 1959 2724 1960
rect 2718 1955 2719 1959
rect 2723 1955 2724 1959
rect 2878 1959 2884 1960
rect 2718 1954 2724 1955
rect 2727 1956 2731 1957
rect 2098 1947 2104 1948
rect 2098 1943 2099 1947
rect 2103 1943 2104 1947
rect 2098 1942 2104 1943
rect 2208 1935 2210 1954
rect 2338 1947 2344 1948
rect 2338 1943 2339 1947
rect 2343 1943 2344 1947
rect 2338 1942 2344 1943
rect 1991 1934 1995 1935
rect 1991 1929 1995 1930
rect 2039 1934 2043 1935
rect 2039 1929 2043 1930
rect 2119 1934 2123 1935
rect 2119 1929 2123 1930
rect 2207 1934 2211 1935
rect 2207 1929 2211 1930
rect 2255 1934 2259 1935
rect 2255 1929 2259 1930
rect 1982 1927 1988 1928
rect 1982 1923 1983 1927
rect 1987 1923 1988 1927
rect 1982 1922 1988 1923
rect 1992 1918 1994 1929
rect 2120 1918 2122 1929
rect 2256 1918 2258 1929
rect 1894 1917 1900 1918
rect 1894 1913 1895 1917
rect 1899 1913 1900 1917
rect 1894 1912 1900 1913
rect 1990 1917 1996 1918
rect 1990 1913 1991 1917
rect 1995 1913 1996 1917
rect 1990 1912 1996 1913
rect 2118 1917 2124 1918
rect 2118 1913 2119 1917
rect 2123 1913 2124 1917
rect 2118 1912 2124 1913
rect 2254 1917 2260 1918
rect 2254 1913 2255 1917
rect 2259 1913 2260 1917
rect 2254 1912 2260 1913
rect 1822 1904 1828 1905
rect 1822 1900 1823 1904
rect 1827 1900 1828 1904
rect 1822 1899 1828 1900
rect 1862 1904 1868 1905
rect 2340 1904 2342 1942
rect 2384 1935 2386 1954
rect 2552 1935 2554 1954
rect 2720 1935 2722 1954
rect 2878 1955 2879 1959
rect 2883 1955 2884 1959
rect 2878 1954 2884 1955
rect 2727 1951 2731 1952
rect 2728 1948 2730 1951
rect 2726 1947 2732 1948
rect 2726 1943 2727 1947
rect 2731 1943 2732 1947
rect 2726 1942 2732 1943
rect 2880 1935 2882 1954
rect 2383 1934 2387 1935
rect 2383 1929 2387 1930
rect 2511 1934 2515 1935
rect 2511 1929 2515 1930
rect 2551 1934 2555 1935
rect 2551 1929 2555 1930
rect 2631 1934 2635 1935
rect 2631 1929 2635 1930
rect 2719 1934 2723 1935
rect 2719 1929 2723 1930
rect 2751 1934 2755 1935
rect 2751 1929 2755 1930
rect 2879 1934 2883 1935
rect 2879 1929 2883 1930
rect 2346 1927 2352 1928
rect 2346 1923 2347 1927
rect 2351 1923 2352 1927
rect 2346 1922 2352 1923
rect 2366 1927 2372 1928
rect 2366 1923 2367 1927
rect 2371 1923 2372 1927
rect 2366 1922 2372 1923
rect 1862 1900 1863 1904
rect 1867 1900 1868 1904
rect 1862 1899 1868 1900
rect 2338 1903 2344 1904
rect 2338 1899 2339 1903
rect 2343 1899 2344 1903
rect 2348 1900 2350 1922
rect 1254 1891 1260 1892
rect 1254 1887 1255 1891
rect 1259 1887 1260 1891
rect 1254 1886 1260 1887
rect 1470 1891 1476 1892
rect 1470 1887 1471 1891
rect 1475 1887 1476 1891
rect 1470 1886 1476 1887
rect 1159 1884 1163 1885
rect 1159 1879 1163 1880
rect 1256 1867 1258 1886
rect 1426 1867 1432 1868
rect 1472 1867 1474 1886
rect 1824 1867 1826 1899
rect 2338 1898 2344 1899
rect 2346 1899 2352 1900
rect 2346 1895 2347 1899
rect 2351 1895 2352 1899
rect 2346 1894 2352 1895
rect 1862 1887 1868 1888
rect 1862 1883 1863 1887
rect 1867 1883 1868 1887
rect 1862 1882 1868 1883
rect 1870 1887 1876 1888
rect 1870 1883 1871 1887
rect 1875 1883 1876 1887
rect 1870 1882 1876 1883
rect 1047 1866 1051 1867
rect 1047 1861 1051 1862
rect 1055 1866 1059 1867
rect 1055 1861 1059 1862
rect 1159 1866 1163 1867
rect 1159 1861 1163 1862
rect 1255 1866 1259 1867
rect 1255 1861 1259 1862
rect 1263 1866 1267 1867
rect 1263 1861 1267 1862
rect 1359 1866 1363 1867
rect 1426 1863 1427 1867
rect 1431 1863 1432 1867
rect 1426 1862 1432 1863
rect 1455 1866 1459 1867
rect 1359 1861 1363 1862
rect 950 1859 956 1860
rect 950 1855 951 1859
rect 955 1855 956 1859
rect 950 1854 956 1855
rect 1056 1850 1058 1861
rect 1110 1859 1116 1860
rect 1110 1855 1111 1859
rect 1115 1855 1116 1859
rect 1110 1854 1116 1855
rect 1112 1851 1114 1854
rect 942 1849 948 1850
rect 942 1845 943 1849
rect 947 1845 948 1849
rect 942 1844 948 1845
rect 1054 1849 1060 1850
rect 1112 1849 1118 1851
rect 1160 1850 1162 1861
rect 1264 1850 1266 1861
rect 1360 1850 1362 1861
rect 1054 1845 1055 1849
rect 1059 1845 1060 1849
rect 1054 1844 1060 1845
rect 762 1831 768 1832
rect 762 1827 763 1831
rect 767 1827 768 1831
rect 762 1826 768 1827
rect 890 1831 896 1832
rect 890 1827 891 1831
rect 895 1827 896 1831
rect 890 1826 896 1827
rect 510 1819 516 1820
rect 510 1815 511 1819
rect 515 1815 516 1819
rect 510 1814 516 1815
rect 406 1809 412 1810
rect 406 1805 407 1809
rect 411 1805 412 1809
rect 406 1804 412 1805
rect 408 1787 410 1804
rect 407 1786 411 1787
rect 407 1781 411 1782
rect 495 1786 499 1787
rect 495 1781 499 1782
rect 496 1776 498 1781
rect 494 1775 500 1776
rect 494 1771 495 1775
rect 499 1771 500 1775
rect 494 1770 500 1771
rect 370 1767 376 1768
rect 110 1765 116 1766
rect 110 1761 111 1765
rect 115 1761 116 1765
rect 370 1763 371 1767
rect 375 1763 376 1767
rect 370 1762 376 1763
rect 110 1760 116 1761
rect 110 1748 116 1749
rect 110 1744 111 1748
rect 115 1744 116 1748
rect 110 1743 116 1744
rect 112 1715 114 1743
rect 142 1735 148 1736
rect 142 1731 143 1735
rect 147 1731 148 1735
rect 142 1730 148 1731
rect 310 1735 316 1736
rect 310 1731 311 1735
rect 315 1731 316 1735
rect 310 1730 316 1731
rect 502 1735 508 1736
rect 502 1731 503 1735
rect 507 1731 508 1735
rect 502 1730 508 1731
rect 134 1723 140 1724
rect 134 1719 135 1723
rect 139 1719 140 1723
rect 134 1718 140 1719
rect 111 1714 115 1715
rect 111 1709 115 1710
rect 112 1685 114 1709
rect 110 1684 116 1685
rect 110 1680 111 1684
rect 115 1680 116 1684
rect 136 1680 138 1718
rect 144 1715 146 1730
rect 312 1715 314 1730
rect 504 1715 506 1730
rect 512 1724 514 1814
rect 550 1809 556 1810
rect 550 1805 551 1809
rect 555 1805 556 1809
rect 550 1804 556 1805
rect 686 1809 692 1810
rect 686 1805 687 1809
rect 691 1805 692 1809
rect 686 1804 692 1805
rect 814 1809 820 1810
rect 814 1805 815 1809
rect 819 1805 820 1809
rect 814 1804 820 1805
rect 934 1809 940 1810
rect 934 1805 935 1809
rect 939 1805 940 1809
rect 934 1804 940 1805
rect 1046 1809 1052 1810
rect 1046 1805 1047 1809
rect 1051 1805 1052 1809
rect 1046 1804 1052 1805
rect 552 1787 554 1804
rect 688 1787 690 1804
rect 816 1787 818 1804
rect 936 1787 938 1804
rect 1048 1787 1050 1804
rect 551 1786 555 1787
rect 551 1781 555 1782
rect 687 1786 691 1787
rect 687 1781 691 1782
rect 815 1786 819 1787
rect 815 1781 819 1782
rect 871 1786 875 1787
rect 871 1781 875 1782
rect 935 1786 939 1787
rect 935 1781 939 1782
rect 1047 1786 1051 1787
rect 1047 1781 1051 1782
rect 688 1776 690 1781
rect 872 1776 874 1781
rect 1048 1776 1050 1781
rect 686 1775 692 1776
rect 686 1771 687 1775
rect 691 1771 692 1775
rect 686 1770 692 1771
rect 870 1775 876 1776
rect 870 1771 871 1775
rect 875 1771 876 1775
rect 870 1770 876 1771
rect 1046 1775 1052 1776
rect 1046 1771 1047 1775
rect 1051 1771 1052 1775
rect 1046 1770 1052 1771
rect 1116 1768 1118 1849
rect 1158 1849 1164 1850
rect 1158 1845 1159 1849
rect 1163 1845 1164 1849
rect 1158 1844 1164 1845
rect 1262 1849 1268 1850
rect 1262 1845 1263 1849
rect 1267 1845 1268 1849
rect 1262 1844 1268 1845
rect 1358 1849 1364 1850
rect 1358 1845 1359 1849
rect 1363 1845 1364 1849
rect 1358 1844 1364 1845
rect 1428 1832 1430 1862
rect 1455 1861 1459 1862
rect 1471 1866 1475 1867
rect 1471 1861 1475 1862
rect 1551 1866 1555 1867
rect 1551 1861 1555 1862
rect 1647 1866 1651 1867
rect 1647 1861 1651 1862
rect 1735 1866 1739 1867
rect 1735 1861 1739 1862
rect 1823 1866 1827 1867
rect 1823 1861 1827 1862
rect 1456 1850 1458 1861
rect 1552 1850 1554 1861
rect 1618 1859 1624 1860
rect 1618 1855 1619 1859
rect 1623 1855 1624 1859
rect 1618 1854 1624 1855
rect 1454 1849 1460 1850
rect 1454 1845 1455 1849
rect 1459 1845 1460 1849
rect 1454 1844 1460 1845
rect 1550 1849 1556 1850
rect 1550 1845 1551 1849
rect 1555 1845 1556 1849
rect 1550 1844 1556 1845
rect 1620 1832 1622 1854
rect 1648 1850 1650 1861
rect 1714 1859 1720 1860
rect 1714 1855 1715 1859
rect 1719 1855 1720 1859
rect 1714 1854 1720 1855
rect 1646 1849 1652 1850
rect 1646 1845 1647 1849
rect 1651 1845 1652 1849
rect 1646 1844 1652 1845
rect 1716 1832 1718 1854
rect 1736 1850 1738 1861
rect 1734 1849 1740 1850
rect 1734 1845 1735 1849
rect 1739 1845 1740 1849
rect 1734 1844 1740 1845
rect 1824 1837 1826 1861
rect 1864 1859 1866 1882
rect 1872 1860 1874 1882
rect 1886 1877 1892 1878
rect 1886 1873 1887 1877
rect 1891 1873 1892 1877
rect 1886 1872 1892 1873
rect 1982 1877 1988 1878
rect 1982 1873 1983 1877
rect 1987 1873 1988 1877
rect 1982 1872 1988 1873
rect 2110 1877 2116 1878
rect 2110 1873 2111 1877
rect 2115 1873 2116 1877
rect 2110 1872 2116 1873
rect 2246 1877 2252 1878
rect 2246 1873 2247 1877
rect 2251 1873 2252 1877
rect 2246 1872 2252 1873
rect 1870 1859 1876 1860
rect 1888 1859 1890 1872
rect 1984 1859 1986 1872
rect 2112 1859 2114 1872
rect 2248 1859 2250 1872
rect 1863 1858 1867 1859
rect 1870 1855 1871 1859
rect 1875 1855 1876 1859
rect 1870 1854 1876 1855
rect 1887 1858 1891 1859
rect 1863 1853 1867 1854
rect 1887 1853 1891 1854
rect 1983 1858 1987 1859
rect 1983 1853 1987 1854
rect 2111 1858 2115 1859
rect 2111 1853 2115 1854
rect 2223 1858 2227 1859
rect 2223 1853 2227 1854
rect 2247 1858 2251 1859
rect 2247 1853 2251 1854
rect 2359 1858 2363 1859
rect 2359 1853 2363 1854
rect 1864 1838 1866 1853
rect 2224 1848 2226 1853
rect 2360 1848 2362 1853
rect 2222 1847 2228 1848
rect 2222 1843 2223 1847
rect 2227 1843 2228 1847
rect 2222 1842 2228 1843
rect 2358 1847 2364 1848
rect 2358 1843 2359 1847
rect 2363 1843 2364 1847
rect 2358 1842 2364 1843
rect 1862 1837 1868 1838
rect 1822 1836 1828 1837
rect 1822 1832 1823 1836
rect 1827 1832 1828 1836
rect 1862 1833 1863 1837
rect 1867 1833 1868 1837
rect 2368 1836 2370 1922
rect 2384 1918 2386 1929
rect 2512 1918 2514 1929
rect 2578 1927 2584 1928
rect 2578 1923 2579 1927
rect 2583 1923 2584 1927
rect 2578 1922 2584 1923
rect 2382 1917 2388 1918
rect 2382 1913 2383 1917
rect 2387 1913 2388 1917
rect 2382 1912 2388 1913
rect 2510 1917 2516 1918
rect 2510 1913 2511 1917
rect 2515 1913 2516 1917
rect 2510 1912 2516 1913
rect 2580 1900 2582 1922
rect 2632 1918 2634 1929
rect 2698 1927 2704 1928
rect 2698 1923 2699 1927
rect 2703 1923 2704 1927
rect 2698 1922 2704 1923
rect 2630 1917 2636 1918
rect 2630 1913 2631 1917
rect 2635 1913 2636 1917
rect 2630 1912 2636 1913
rect 2700 1900 2702 1922
rect 2752 1918 2754 1929
rect 2818 1927 2824 1928
rect 2818 1923 2819 1927
rect 2823 1923 2824 1927
rect 2818 1922 2824 1923
rect 2750 1917 2756 1918
rect 2750 1913 2751 1917
rect 2755 1913 2756 1917
rect 2750 1912 2756 1913
rect 2820 1900 2822 1922
rect 2880 1918 2882 1929
rect 3000 1928 3002 1970
rect 3046 1959 3052 1960
rect 3046 1955 3047 1959
rect 3051 1955 3052 1959
rect 3046 1954 3052 1955
rect 3048 1935 3050 1954
rect 3152 1948 3154 1970
rect 3160 1957 3162 1970
rect 3574 1968 3575 1972
rect 3579 1968 3580 1972
rect 3574 1967 3580 1968
rect 3214 1959 3220 1960
rect 3159 1956 3163 1957
rect 3214 1955 3215 1959
rect 3219 1955 3220 1959
rect 3214 1954 3220 1955
rect 3159 1951 3163 1952
rect 3150 1947 3156 1948
rect 3150 1943 3151 1947
rect 3155 1943 3156 1947
rect 3150 1942 3156 1943
rect 3216 1935 3218 1954
rect 3576 1935 3578 1967
rect 3007 1934 3011 1935
rect 3007 1929 3011 1930
rect 3047 1934 3051 1935
rect 3047 1929 3051 1930
rect 3215 1934 3219 1935
rect 3215 1929 3219 1930
rect 3575 1934 3579 1935
rect 3575 1929 3579 1930
rect 2946 1927 2952 1928
rect 2946 1923 2947 1927
rect 2951 1923 2952 1927
rect 2946 1922 2952 1923
rect 2998 1927 3004 1928
rect 2998 1923 2999 1927
rect 3003 1923 3004 1927
rect 2998 1922 3004 1923
rect 2878 1917 2884 1918
rect 2878 1913 2879 1917
rect 2883 1913 2884 1917
rect 2878 1912 2884 1913
rect 2948 1900 2950 1922
rect 3008 1918 3010 1929
rect 3006 1917 3012 1918
rect 3006 1913 3007 1917
rect 3011 1913 3012 1917
rect 3006 1912 3012 1913
rect 3576 1905 3578 1929
rect 3574 1904 3580 1905
rect 3574 1900 3575 1904
rect 3579 1900 3580 1904
rect 2578 1899 2584 1900
rect 2578 1895 2579 1899
rect 2583 1895 2584 1899
rect 2578 1894 2584 1895
rect 2698 1899 2704 1900
rect 2698 1895 2699 1899
rect 2703 1895 2704 1899
rect 2698 1894 2704 1895
rect 2818 1899 2824 1900
rect 2818 1895 2819 1899
rect 2823 1895 2824 1899
rect 2818 1894 2824 1895
rect 2946 1899 2952 1900
rect 3574 1899 3580 1900
rect 2946 1895 2947 1899
rect 2951 1895 2952 1899
rect 2946 1894 2952 1895
rect 2510 1887 2516 1888
rect 2510 1883 2511 1887
rect 2515 1883 2516 1887
rect 2510 1882 2516 1883
rect 3574 1887 3580 1888
rect 3574 1883 3575 1887
rect 3579 1883 3580 1887
rect 3574 1882 3580 1883
rect 2374 1877 2380 1878
rect 2374 1873 2375 1877
rect 2379 1873 2380 1877
rect 2374 1872 2380 1873
rect 2502 1877 2508 1878
rect 2502 1873 2503 1877
rect 2507 1873 2508 1877
rect 2502 1872 2508 1873
rect 2376 1859 2378 1872
rect 2504 1859 2506 1872
rect 2375 1858 2379 1859
rect 2375 1853 2379 1854
rect 2495 1858 2499 1859
rect 2495 1853 2499 1854
rect 2503 1858 2507 1859
rect 2503 1853 2507 1854
rect 2496 1848 2498 1853
rect 2494 1847 2500 1848
rect 2494 1843 2495 1847
rect 2499 1843 2500 1847
rect 2494 1842 2500 1843
rect 1862 1832 1868 1833
rect 2366 1835 2372 1836
rect 1426 1831 1432 1832
rect 1426 1827 1427 1831
rect 1431 1827 1432 1831
rect 1426 1826 1432 1827
rect 1618 1831 1624 1832
rect 1618 1827 1619 1831
rect 1623 1827 1624 1831
rect 1618 1826 1624 1827
rect 1714 1831 1720 1832
rect 1822 1831 1828 1832
rect 2366 1831 2367 1835
rect 2371 1831 2372 1835
rect 1714 1827 1715 1831
rect 1719 1827 1720 1831
rect 2366 1830 2372 1831
rect 1714 1826 1720 1827
rect 1862 1820 1868 1821
rect 1550 1819 1556 1820
rect 1550 1815 1551 1819
rect 1555 1815 1556 1819
rect 1550 1814 1556 1815
rect 1822 1819 1828 1820
rect 1822 1815 1823 1819
rect 1827 1815 1828 1819
rect 1862 1816 1863 1820
rect 1867 1816 1868 1820
rect 1862 1815 1868 1816
rect 1822 1814 1828 1815
rect 1150 1809 1156 1810
rect 1150 1805 1151 1809
rect 1155 1805 1156 1809
rect 1150 1804 1156 1805
rect 1254 1809 1260 1810
rect 1254 1805 1255 1809
rect 1259 1805 1260 1809
rect 1254 1804 1260 1805
rect 1350 1809 1356 1810
rect 1350 1805 1351 1809
rect 1355 1805 1356 1809
rect 1350 1804 1356 1805
rect 1446 1809 1452 1810
rect 1446 1805 1447 1809
rect 1451 1805 1452 1809
rect 1446 1804 1452 1805
rect 1542 1809 1548 1810
rect 1542 1805 1543 1809
rect 1547 1805 1548 1809
rect 1542 1804 1548 1805
rect 1152 1787 1154 1804
rect 1256 1787 1258 1804
rect 1352 1787 1354 1804
rect 1390 1803 1396 1804
rect 1390 1799 1391 1803
rect 1395 1799 1396 1803
rect 1390 1798 1396 1799
rect 1151 1786 1155 1787
rect 1151 1781 1155 1782
rect 1215 1786 1219 1787
rect 1215 1781 1219 1782
rect 1255 1786 1259 1787
rect 1255 1781 1259 1782
rect 1351 1786 1355 1787
rect 1351 1781 1355 1782
rect 1375 1786 1379 1787
rect 1375 1781 1379 1782
rect 1216 1776 1218 1781
rect 1376 1776 1378 1781
rect 1214 1775 1220 1776
rect 1214 1771 1215 1775
rect 1219 1771 1220 1775
rect 1214 1770 1220 1771
rect 1374 1775 1380 1776
rect 1374 1771 1375 1775
rect 1379 1771 1380 1775
rect 1374 1770 1380 1771
rect 1114 1767 1120 1768
rect 1114 1763 1115 1767
rect 1119 1763 1120 1767
rect 1114 1762 1120 1763
rect 694 1735 700 1736
rect 694 1731 695 1735
rect 699 1731 700 1735
rect 694 1730 700 1731
rect 878 1735 884 1736
rect 878 1731 879 1735
rect 883 1731 884 1735
rect 878 1730 884 1731
rect 1054 1735 1060 1736
rect 1054 1731 1055 1735
rect 1059 1731 1060 1735
rect 1054 1730 1060 1731
rect 1222 1735 1228 1736
rect 1222 1731 1223 1735
rect 1227 1731 1228 1735
rect 1222 1730 1228 1731
rect 1382 1735 1388 1736
rect 1382 1731 1383 1735
rect 1387 1731 1388 1735
rect 1382 1730 1388 1731
rect 510 1723 516 1724
rect 510 1719 511 1723
rect 515 1719 516 1723
rect 510 1718 516 1719
rect 696 1715 698 1730
rect 880 1715 882 1730
rect 1056 1715 1058 1730
rect 1082 1723 1088 1724
rect 1082 1719 1083 1723
rect 1087 1719 1088 1723
rect 1082 1718 1088 1719
rect 143 1714 147 1715
rect 143 1709 147 1710
rect 287 1714 291 1715
rect 287 1709 291 1710
rect 311 1714 315 1715
rect 311 1709 315 1710
rect 471 1714 475 1715
rect 471 1709 475 1710
rect 503 1714 507 1715
rect 503 1709 507 1710
rect 655 1714 659 1715
rect 655 1709 659 1710
rect 695 1714 699 1715
rect 695 1709 699 1710
rect 839 1714 843 1715
rect 839 1709 843 1710
rect 879 1714 883 1715
rect 879 1709 883 1710
rect 1023 1714 1027 1715
rect 1023 1709 1027 1710
rect 1055 1714 1059 1715
rect 1055 1709 1059 1710
rect 144 1698 146 1709
rect 288 1698 290 1709
rect 382 1707 388 1708
rect 382 1703 383 1707
rect 387 1703 388 1707
rect 382 1702 388 1703
rect 142 1697 148 1698
rect 142 1693 143 1697
rect 147 1693 148 1697
rect 142 1692 148 1693
rect 286 1697 292 1698
rect 286 1693 287 1697
rect 291 1693 292 1697
rect 286 1692 292 1693
rect 384 1680 386 1702
rect 472 1698 474 1709
rect 656 1698 658 1709
rect 750 1707 756 1708
rect 750 1703 751 1707
rect 755 1703 756 1707
rect 750 1702 756 1703
rect 470 1697 476 1698
rect 470 1693 471 1697
rect 475 1693 476 1697
rect 470 1692 476 1693
rect 654 1697 660 1698
rect 654 1693 655 1697
rect 659 1693 660 1697
rect 654 1692 660 1693
rect 752 1680 754 1702
rect 840 1698 842 1709
rect 998 1707 1004 1708
rect 998 1703 999 1707
rect 1003 1703 1004 1707
rect 998 1702 1004 1703
rect 838 1697 844 1698
rect 838 1693 839 1697
rect 843 1693 844 1697
rect 838 1692 844 1693
rect 110 1679 116 1680
rect 134 1679 140 1680
rect 134 1675 135 1679
rect 139 1675 140 1679
rect 134 1674 140 1675
rect 382 1679 388 1680
rect 382 1675 383 1679
rect 387 1675 388 1679
rect 382 1674 388 1675
rect 750 1679 756 1680
rect 750 1675 751 1679
rect 755 1675 756 1679
rect 750 1674 756 1675
rect 110 1667 116 1668
rect 110 1663 111 1667
rect 115 1663 116 1667
rect 110 1662 116 1663
rect 286 1667 292 1668
rect 286 1663 287 1667
rect 291 1663 292 1667
rect 286 1662 292 1663
rect 112 1639 114 1662
rect 134 1657 140 1658
rect 134 1653 135 1657
rect 139 1653 140 1657
rect 134 1652 140 1653
rect 278 1657 284 1658
rect 278 1653 279 1657
rect 283 1653 284 1657
rect 278 1652 284 1653
rect 136 1639 138 1652
rect 280 1639 282 1652
rect 111 1638 115 1639
rect 111 1633 115 1634
rect 135 1638 139 1639
rect 135 1633 139 1634
rect 271 1638 275 1639
rect 271 1633 275 1634
rect 279 1638 283 1639
rect 279 1633 283 1634
rect 112 1618 114 1633
rect 136 1628 138 1633
rect 272 1628 274 1633
rect 134 1627 140 1628
rect 134 1623 135 1627
rect 139 1623 140 1627
rect 134 1622 140 1623
rect 270 1627 276 1628
rect 270 1623 271 1627
rect 275 1623 276 1627
rect 270 1622 276 1623
rect 110 1617 116 1618
rect 110 1613 111 1617
rect 115 1613 116 1617
rect 110 1612 116 1613
rect 110 1600 116 1601
rect 110 1596 111 1600
rect 115 1596 116 1600
rect 110 1595 116 1596
rect 112 1571 114 1595
rect 142 1587 148 1588
rect 142 1583 143 1587
rect 147 1583 148 1587
rect 142 1582 148 1583
rect 278 1587 284 1588
rect 278 1583 279 1587
rect 283 1583 284 1587
rect 278 1582 284 1583
rect 134 1575 140 1576
rect 134 1571 135 1575
rect 139 1571 140 1575
rect 144 1571 146 1582
rect 280 1571 282 1582
rect 288 1576 290 1662
rect 462 1657 468 1658
rect 462 1653 463 1657
rect 467 1653 468 1657
rect 462 1652 468 1653
rect 646 1657 652 1658
rect 646 1653 647 1657
rect 651 1653 652 1657
rect 646 1652 652 1653
rect 830 1657 836 1658
rect 830 1653 831 1657
rect 835 1653 836 1657
rect 830 1652 836 1653
rect 464 1639 466 1652
rect 648 1639 650 1652
rect 832 1639 834 1652
rect 447 1638 451 1639
rect 447 1633 451 1634
rect 463 1638 467 1639
rect 463 1633 467 1634
rect 631 1638 635 1639
rect 631 1633 635 1634
rect 647 1638 651 1639
rect 647 1633 651 1634
rect 815 1638 819 1639
rect 815 1633 819 1634
rect 831 1638 835 1639
rect 831 1633 835 1634
rect 991 1638 995 1639
rect 991 1633 995 1634
rect 448 1628 450 1633
rect 632 1628 634 1633
rect 816 1628 818 1633
rect 992 1628 994 1633
rect 446 1627 452 1628
rect 446 1623 447 1627
rect 451 1623 452 1627
rect 446 1622 452 1623
rect 630 1627 636 1628
rect 630 1623 631 1627
rect 635 1623 636 1627
rect 630 1622 636 1623
rect 814 1627 820 1628
rect 814 1623 815 1627
rect 819 1623 820 1627
rect 814 1622 820 1623
rect 990 1627 996 1628
rect 990 1623 991 1627
rect 995 1623 996 1627
rect 990 1622 996 1623
rect 1000 1616 1002 1702
rect 1024 1698 1026 1709
rect 1022 1697 1028 1698
rect 1022 1693 1023 1697
rect 1027 1693 1028 1697
rect 1022 1692 1028 1693
rect 1084 1684 1086 1718
rect 1224 1715 1226 1730
rect 1384 1715 1386 1730
rect 1392 1724 1394 1798
rect 1448 1787 1450 1804
rect 1544 1787 1546 1804
rect 1447 1786 1451 1787
rect 1447 1781 1451 1782
rect 1535 1786 1539 1787
rect 1535 1781 1539 1782
rect 1543 1786 1547 1787
rect 1543 1781 1547 1782
rect 1536 1776 1538 1781
rect 1534 1775 1540 1776
rect 1534 1771 1535 1775
rect 1539 1771 1540 1775
rect 1534 1770 1540 1771
rect 1542 1735 1548 1736
rect 1542 1731 1543 1735
rect 1547 1731 1548 1735
rect 1542 1730 1548 1731
rect 1390 1723 1396 1724
rect 1390 1719 1391 1723
rect 1395 1719 1396 1723
rect 1390 1718 1396 1719
rect 1544 1715 1546 1730
rect 1552 1724 1554 1814
rect 1638 1809 1644 1810
rect 1638 1805 1639 1809
rect 1643 1805 1644 1809
rect 1638 1804 1644 1805
rect 1726 1809 1732 1810
rect 1726 1805 1727 1809
rect 1731 1805 1732 1809
rect 1726 1804 1732 1805
rect 1640 1787 1642 1804
rect 1728 1787 1730 1804
rect 1824 1787 1826 1814
rect 1864 1787 1866 1815
rect 2230 1807 2236 1808
rect 2230 1803 2231 1807
rect 2235 1803 2236 1807
rect 2230 1802 2236 1803
rect 2366 1807 2372 1808
rect 2366 1803 2367 1807
rect 2371 1803 2372 1807
rect 2366 1802 2372 1803
rect 2502 1807 2508 1808
rect 2502 1803 2503 1807
rect 2507 1803 2508 1807
rect 2502 1802 2508 1803
rect 2232 1787 2234 1802
rect 2330 1795 2336 1796
rect 2330 1791 2331 1795
rect 2335 1791 2336 1795
rect 2330 1790 2336 1791
rect 1639 1786 1643 1787
rect 1639 1781 1643 1782
rect 1703 1786 1707 1787
rect 1703 1781 1707 1782
rect 1727 1786 1731 1787
rect 1727 1781 1731 1782
rect 1823 1786 1827 1787
rect 1823 1781 1827 1782
rect 1863 1786 1867 1787
rect 1863 1781 1867 1782
rect 2231 1786 2235 1787
rect 2231 1781 2235 1782
rect 2271 1786 2275 1787
rect 2271 1781 2275 1782
rect 1704 1776 1706 1781
rect 1702 1775 1708 1776
rect 1702 1771 1703 1775
rect 1707 1771 1708 1775
rect 1702 1770 1708 1771
rect 1824 1766 1826 1781
rect 1822 1765 1828 1766
rect 1822 1761 1823 1765
rect 1827 1761 1828 1765
rect 1822 1760 1828 1761
rect 1864 1757 1866 1781
rect 2272 1770 2274 1781
rect 2270 1769 2276 1770
rect 2270 1765 2271 1769
rect 2275 1765 2276 1769
rect 2270 1764 2276 1765
rect 1862 1756 1868 1757
rect 2332 1756 2334 1790
rect 2368 1787 2370 1802
rect 2504 1787 2506 1802
rect 2512 1796 2514 1882
rect 2622 1877 2628 1878
rect 2622 1873 2623 1877
rect 2627 1873 2628 1877
rect 2622 1872 2628 1873
rect 2742 1877 2748 1878
rect 2742 1873 2743 1877
rect 2747 1873 2748 1877
rect 2742 1872 2748 1873
rect 2870 1877 2876 1878
rect 2870 1873 2871 1877
rect 2875 1873 2876 1877
rect 2870 1872 2876 1873
rect 2998 1877 3004 1878
rect 2998 1873 2999 1877
rect 3003 1873 3004 1877
rect 2998 1872 3004 1873
rect 2624 1859 2626 1872
rect 2744 1859 2746 1872
rect 2872 1859 2874 1872
rect 3000 1859 3002 1872
rect 3576 1859 3578 1882
rect 2623 1858 2627 1859
rect 2623 1853 2627 1854
rect 2743 1858 2747 1859
rect 2743 1853 2747 1854
rect 2863 1858 2867 1859
rect 2863 1853 2867 1854
rect 2871 1858 2875 1859
rect 2871 1853 2875 1854
rect 2991 1858 2995 1859
rect 2991 1853 2995 1854
rect 2999 1858 3003 1859
rect 2999 1853 3003 1854
rect 3575 1858 3579 1859
rect 3575 1853 3579 1854
rect 2624 1848 2626 1853
rect 2744 1848 2746 1853
rect 2864 1848 2866 1853
rect 2992 1848 2994 1853
rect 2622 1847 2628 1848
rect 2622 1843 2623 1847
rect 2627 1843 2628 1847
rect 2622 1842 2628 1843
rect 2742 1847 2748 1848
rect 2742 1843 2743 1847
rect 2747 1843 2748 1847
rect 2742 1842 2748 1843
rect 2862 1847 2868 1848
rect 2862 1843 2863 1847
rect 2867 1843 2868 1847
rect 2862 1842 2868 1843
rect 2990 1847 2996 1848
rect 2990 1843 2991 1847
rect 2995 1843 2996 1847
rect 2990 1842 2996 1843
rect 2930 1839 2936 1840
rect 2930 1835 2931 1839
rect 2935 1835 2936 1839
rect 3576 1838 3578 1853
rect 2930 1834 2936 1835
rect 3574 1837 3580 1838
rect 2630 1807 2636 1808
rect 2630 1803 2631 1807
rect 2635 1803 2636 1807
rect 2630 1802 2636 1803
rect 2750 1807 2756 1808
rect 2750 1803 2751 1807
rect 2755 1803 2756 1807
rect 2750 1802 2756 1803
rect 2870 1807 2876 1808
rect 2870 1803 2871 1807
rect 2875 1803 2876 1807
rect 2870 1802 2876 1803
rect 2510 1795 2516 1796
rect 2510 1791 2511 1795
rect 2515 1791 2516 1795
rect 2510 1790 2516 1791
rect 2632 1787 2634 1802
rect 2752 1787 2754 1802
rect 2872 1787 2874 1802
rect 2932 1788 2934 1834
rect 3574 1833 3575 1837
rect 3579 1833 3580 1837
rect 3574 1832 3580 1833
rect 3574 1820 3580 1821
rect 3574 1816 3575 1820
rect 3579 1816 3580 1820
rect 3574 1815 3580 1816
rect 2998 1807 3004 1808
rect 2998 1803 2999 1807
rect 3003 1803 3004 1807
rect 2998 1802 3004 1803
rect 2930 1787 2936 1788
rect 3000 1787 3002 1802
rect 3576 1787 3578 1815
rect 2359 1786 2363 1787
rect 2359 1781 2363 1782
rect 2367 1786 2371 1787
rect 2367 1781 2371 1782
rect 2455 1786 2459 1787
rect 2455 1781 2459 1782
rect 2503 1786 2507 1787
rect 2503 1781 2507 1782
rect 2559 1786 2563 1787
rect 2559 1781 2563 1782
rect 2631 1786 2635 1787
rect 2631 1781 2635 1782
rect 2663 1786 2667 1787
rect 2663 1781 2667 1782
rect 2751 1786 2755 1787
rect 2751 1781 2755 1782
rect 2759 1786 2763 1787
rect 2759 1781 2763 1782
rect 2863 1786 2867 1787
rect 2863 1781 2867 1782
rect 2871 1786 2875 1787
rect 2930 1783 2931 1787
rect 2935 1783 2936 1787
rect 2930 1782 2936 1783
rect 2967 1786 2971 1787
rect 2871 1781 2875 1782
rect 2967 1781 2971 1782
rect 2999 1786 3003 1787
rect 2999 1781 3003 1782
rect 3071 1786 3075 1787
rect 3071 1781 3075 1782
rect 3175 1786 3179 1787
rect 3175 1781 3179 1782
rect 3575 1786 3579 1787
rect 3575 1781 3579 1782
rect 2338 1779 2344 1780
rect 2338 1775 2339 1779
rect 2343 1775 2344 1779
rect 2338 1774 2344 1775
rect 1862 1752 1863 1756
rect 1867 1752 1868 1756
rect 1862 1751 1868 1752
rect 2330 1755 2336 1756
rect 2330 1751 2331 1755
rect 2335 1751 2336 1755
rect 2340 1752 2342 1774
rect 2360 1770 2362 1781
rect 2426 1779 2432 1780
rect 2426 1775 2427 1779
rect 2431 1775 2432 1779
rect 2426 1774 2432 1775
rect 2358 1769 2364 1770
rect 2358 1765 2359 1769
rect 2363 1765 2364 1769
rect 2358 1764 2364 1765
rect 2428 1752 2430 1774
rect 2456 1770 2458 1781
rect 2522 1779 2528 1780
rect 2522 1775 2523 1779
rect 2527 1775 2528 1779
rect 2522 1774 2528 1775
rect 2454 1769 2460 1770
rect 2454 1765 2455 1769
rect 2459 1765 2460 1769
rect 2454 1764 2460 1765
rect 2524 1752 2526 1774
rect 2560 1770 2562 1781
rect 2664 1770 2666 1781
rect 2722 1779 2728 1780
rect 2722 1775 2723 1779
rect 2727 1775 2728 1779
rect 2722 1774 2728 1775
rect 2558 1769 2564 1770
rect 2558 1765 2559 1769
rect 2563 1765 2564 1769
rect 2558 1764 2564 1765
rect 2662 1769 2668 1770
rect 2662 1765 2663 1769
rect 2667 1765 2668 1769
rect 2662 1764 2668 1765
rect 2330 1750 2336 1751
rect 2338 1751 2344 1752
rect 1822 1748 1828 1749
rect 1822 1744 1823 1748
rect 1827 1744 1828 1748
rect 2338 1747 2339 1751
rect 2343 1747 2344 1751
rect 2338 1746 2344 1747
rect 2426 1751 2432 1752
rect 2426 1747 2427 1751
rect 2431 1747 2432 1751
rect 2426 1746 2432 1747
rect 2522 1751 2528 1752
rect 2522 1747 2523 1751
rect 2527 1747 2528 1751
rect 2522 1746 2528 1747
rect 1822 1743 1828 1744
rect 1710 1735 1716 1736
rect 1710 1731 1711 1735
rect 1715 1731 1716 1735
rect 1710 1730 1716 1731
rect 1550 1723 1556 1724
rect 1550 1719 1551 1723
rect 1555 1719 1556 1723
rect 1550 1718 1556 1719
rect 1712 1715 1714 1730
rect 1824 1715 1826 1743
rect 1862 1739 1868 1740
rect 1862 1735 1863 1739
rect 1867 1735 1868 1739
rect 1862 1734 1868 1735
rect 1864 1715 1866 1734
rect 2262 1729 2268 1730
rect 2262 1725 2263 1729
rect 2267 1725 2268 1729
rect 2262 1724 2268 1725
rect 2350 1729 2356 1730
rect 2350 1725 2351 1729
rect 2355 1725 2356 1729
rect 2350 1724 2356 1725
rect 2446 1729 2452 1730
rect 2446 1725 2447 1729
rect 2451 1725 2452 1729
rect 2446 1724 2452 1725
rect 2550 1729 2556 1730
rect 2550 1725 2551 1729
rect 2555 1725 2556 1729
rect 2550 1724 2556 1725
rect 2654 1729 2660 1730
rect 2654 1725 2655 1729
rect 2659 1725 2660 1729
rect 2654 1724 2660 1725
rect 2264 1715 2266 1724
rect 2352 1715 2354 1724
rect 2448 1715 2450 1724
rect 2552 1715 2554 1724
rect 2656 1715 2658 1724
rect 1191 1714 1195 1715
rect 1191 1709 1195 1710
rect 1223 1714 1227 1715
rect 1223 1709 1227 1710
rect 1359 1714 1363 1715
rect 1359 1709 1363 1710
rect 1383 1714 1387 1715
rect 1383 1709 1387 1710
rect 1527 1714 1531 1715
rect 1527 1709 1531 1710
rect 1543 1714 1547 1715
rect 1543 1709 1547 1710
rect 1695 1714 1699 1715
rect 1695 1709 1699 1710
rect 1711 1714 1715 1715
rect 1711 1709 1715 1710
rect 1823 1714 1827 1715
rect 1823 1709 1827 1710
rect 1863 1714 1867 1715
rect 1863 1709 1867 1710
rect 2247 1714 2251 1715
rect 2247 1709 2251 1710
rect 2263 1714 2267 1715
rect 2263 1709 2267 1710
rect 2351 1714 2355 1715
rect 2351 1709 2355 1710
rect 2367 1714 2371 1715
rect 2367 1709 2371 1710
rect 2447 1714 2451 1715
rect 2447 1709 2451 1710
rect 2495 1714 2499 1715
rect 2495 1709 2499 1710
rect 2551 1714 2555 1715
rect 2551 1709 2555 1710
rect 2623 1714 2627 1715
rect 2623 1709 2627 1710
rect 2655 1714 2659 1715
rect 2655 1709 2659 1710
rect 1192 1698 1194 1709
rect 1360 1698 1362 1709
rect 1426 1707 1432 1708
rect 1426 1703 1427 1707
rect 1431 1703 1432 1707
rect 1426 1702 1432 1703
rect 1190 1697 1196 1698
rect 1190 1693 1191 1697
rect 1195 1693 1196 1697
rect 1190 1692 1196 1693
rect 1358 1697 1364 1698
rect 1358 1693 1359 1697
rect 1363 1693 1364 1697
rect 1358 1692 1364 1693
rect 1082 1683 1088 1684
rect 1082 1679 1083 1683
rect 1087 1679 1088 1683
rect 1428 1680 1430 1702
rect 1528 1698 1530 1709
rect 1696 1698 1698 1709
rect 1526 1697 1532 1698
rect 1526 1693 1527 1697
rect 1531 1693 1532 1697
rect 1526 1692 1532 1693
rect 1694 1697 1700 1698
rect 1694 1693 1695 1697
rect 1699 1693 1700 1697
rect 1694 1692 1700 1693
rect 1824 1685 1826 1709
rect 1864 1694 1866 1709
rect 2248 1704 2250 1709
rect 2368 1704 2370 1709
rect 2496 1704 2498 1709
rect 2624 1704 2626 1709
rect 2246 1703 2252 1704
rect 2246 1699 2247 1703
rect 2251 1699 2252 1703
rect 2246 1698 2252 1699
rect 2366 1703 2372 1704
rect 2366 1699 2367 1703
rect 2371 1699 2372 1703
rect 2366 1698 2372 1699
rect 2494 1703 2500 1704
rect 2494 1699 2495 1703
rect 2499 1699 2500 1703
rect 2494 1698 2500 1699
rect 2622 1703 2628 1704
rect 2622 1699 2623 1703
rect 2627 1699 2628 1703
rect 2622 1698 2628 1699
rect 2724 1696 2726 1774
rect 2760 1770 2762 1781
rect 2864 1770 2866 1781
rect 2968 1770 2970 1781
rect 3072 1770 3074 1781
rect 3176 1770 3178 1781
rect 2758 1769 2764 1770
rect 2758 1765 2759 1769
rect 2763 1765 2764 1769
rect 2758 1764 2764 1765
rect 2862 1769 2868 1770
rect 2862 1765 2863 1769
rect 2867 1765 2868 1769
rect 2862 1764 2868 1765
rect 2966 1769 2972 1770
rect 2966 1765 2967 1769
rect 2971 1765 2972 1769
rect 2966 1764 2972 1765
rect 3070 1769 3076 1770
rect 3070 1765 3071 1769
rect 3075 1765 3076 1769
rect 3070 1764 3076 1765
rect 3174 1769 3180 1770
rect 3174 1765 3175 1769
rect 3179 1765 3180 1769
rect 3174 1764 3180 1765
rect 3576 1757 3578 1781
rect 3574 1756 3580 1757
rect 3574 1752 3575 1756
rect 3579 1752 3580 1756
rect 3574 1751 3580 1752
rect 3574 1739 3580 1740
rect 3574 1735 3575 1739
rect 3579 1735 3580 1739
rect 3574 1734 3580 1735
rect 2750 1729 2756 1730
rect 2750 1725 2751 1729
rect 2755 1725 2756 1729
rect 2750 1724 2756 1725
rect 2854 1729 2860 1730
rect 2854 1725 2855 1729
rect 2859 1725 2860 1729
rect 2854 1724 2860 1725
rect 2958 1729 2964 1730
rect 2958 1725 2959 1729
rect 2963 1725 2964 1729
rect 2958 1724 2964 1725
rect 3062 1729 3068 1730
rect 3062 1725 3063 1729
rect 3067 1725 3068 1729
rect 3062 1724 3068 1725
rect 3166 1729 3172 1730
rect 3166 1725 3167 1729
rect 3171 1725 3172 1729
rect 3166 1724 3172 1725
rect 2752 1715 2754 1724
rect 2856 1715 2858 1724
rect 2902 1723 2908 1724
rect 2902 1719 2903 1723
rect 2907 1719 2908 1723
rect 2902 1718 2908 1719
rect 2751 1714 2755 1715
rect 2751 1709 2755 1710
rect 2759 1714 2763 1715
rect 2759 1709 2763 1710
rect 2855 1714 2859 1715
rect 2855 1709 2859 1710
rect 2887 1714 2891 1715
rect 2887 1709 2891 1710
rect 2760 1704 2762 1709
rect 2888 1704 2890 1709
rect 2758 1703 2764 1704
rect 2758 1699 2759 1703
rect 2763 1699 2764 1703
rect 2758 1698 2764 1699
rect 2886 1703 2892 1704
rect 2886 1699 2887 1703
rect 2891 1699 2892 1703
rect 2886 1698 2892 1699
rect 2722 1695 2728 1696
rect 1862 1693 1868 1694
rect 1862 1689 1863 1693
rect 1867 1689 1868 1693
rect 2722 1691 2723 1695
rect 2727 1691 2728 1695
rect 2722 1690 2728 1691
rect 1862 1688 1868 1689
rect 1822 1684 1828 1685
rect 1822 1680 1823 1684
rect 1827 1680 1828 1684
rect 1082 1678 1088 1679
rect 1426 1679 1432 1680
rect 1822 1679 1828 1680
rect 1426 1675 1427 1679
rect 1431 1675 1432 1679
rect 1426 1674 1432 1675
rect 1862 1676 1868 1677
rect 1862 1672 1863 1676
rect 1867 1672 1868 1676
rect 1862 1671 1868 1672
rect 1166 1667 1172 1668
rect 1166 1663 1167 1667
rect 1171 1663 1172 1667
rect 1166 1662 1172 1663
rect 1822 1667 1828 1668
rect 1822 1663 1823 1667
rect 1827 1663 1828 1667
rect 1822 1662 1828 1663
rect 1014 1657 1020 1658
rect 1014 1653 1015 1657
rect 1019 1653 1020 1657
rect 1014 1652 1020 1653
rect 1016 1639 1018 1652
rect 1015 1638 1019 1639
rect 1015 1633 1019 1634
rect 1151 1638 1155 1639
rect 1151 1633 1155 1634
rect 1152 1628 1154 1633
rect 1150 1627 1156 1628
rect 1150 1623 1151 1627
rect 1155 1623 1156 1627
rect 1150 1622 1156 1623
rect 998 1615 1004 1616
rect 998 1611 999 1615
rect 1003 1611 1004 1615
rect 998 1610 1004 1611
rect 454 1587 460 1588
rect 454 1583 455 1587
rect 459 1583 460 1587
rect 454 1582 460 1583
rect 638 1587 644 1588
rect 638 1583 639 1587
rect 643 1583 644 1587
rect 638 1582 644 1583
rect 822 1587 828 1588
rect 822 1583 823 1587
rect 827 1583 828 1587
rect 822 1582 828 1583
rect 998 1587 1004 1588
rect 998 1583 999 1587
rect 1003 1583 1004 1587
rect 998 1582 1004 1583
rect 1158 1587 1164 1588
rect 1158 1583 1159 1587
rect 1163 1583 1164 1587
rect 1158 1582 1164 1583
rect 286 1575 292 1576
rect 286 1571 287 1575
rect 291 1571 292 1575
rect 456 1571 458 1582
rect 640 1571 642 1582
rect 824 1571 826 1582
rect 1000 1571 1002 1582
rect 1026 1575 1032 1576
rect 1026 1571 1027 1575
rect 1031 1571 1032 1575
rect 1160 1571 1162 1582
rect 1168 1576 1170 1662
rect 1182 1657 1188 1658
rect 1182 1653 1183 1657
rect 1187 1653 1188 1657
rect 1182 1652 1188 1653
rect 1350 1657 1356 1658
rect 1350 1653 1351 1657
rect 1355 1653 1356 1657
rect 1350 1652 1356 1653
rect 1518 1657 1524 1658
rect 1518 1653 1519 1657
rect 1523 1653 1524 1657
rect 1518 1652 1524 1653
rect 1686 1657 1692 1658
rect 1686 1653 1687 1657
rect 1691 1653 1692 1657
rect 1686 1652 1692 1653
rect 1184 1639 1186 1652
rect 1352 1639 1354 1652
rect 1520 1639 1522 1652
rect 1688 1639 1690 1652
rect 1824 1639 1826 1662
rect 1864 1643 1866 1671
rect 2254 1663 2260 1664
rect 2254 1659 2255 1663
rect 2259 1659 2260 1663
rect 2254 1658 2260 1659
rect 2374 1663 2380 1664
rect 2374 1659 2375 1663
rect 2379 1659 2380 1663
rect 2374 1658 2380 1659
rect 2502 1663 2508 1664
rect 2502 1659 2503 1663
rect 2507 1659 2508 1663
rect 2502 1658 2508 1659
rect 2630 1663 2636 1664
rect 2630 1659 2631 1663
rect 2635 1659 2636 1663
rect 2630 1658 2636 1659
rect 2766 1663 2772 1664
rect 2766 1659 2767 1663
rect 2771 1659 2772 1663
rect 2766 1658 2772 1659
rect 2894 1663 2900 1664
rect 2894 1659 2895 1663
rect 2899 1659 2900 1663
rect 2894 1658 2900 1659
rect 2256 1643 2258 1658
rect 2376 1643 2378 1658
rect 2504 1643 2506 1658
rect 2632 1643 2634 1658
rect 2768 1643 2770 1658
rect 2896 1643 2898 1658
rect 2904 1652 2906 1718
rect 2960 1715 2962 1724
rect 3064 1715 3066 1724
rect 3168 1715 3170 1724
rect 3576 1715 3578 1734
rect 2959 1714 2963 1715
rect 2959 1709 2963 1710
rect 3015 1714 3019 1715
rect 3015 1709 3019 1710
rect 3063 1714 3067 1715
rect 3063 1709 3067 1710
rect 3135 1714 3139 1715
rect 3135 1709 3139 1710
rect 3167 1714 3171 1715
rect 3167 1709 3171 1710
rect 3247 1714 3251 1715
rect 3247 1709 3251 1710
rect 3367 1714 3371 1715
rect 3367 1709 3371 1710
rect 3479 1714 3483 1715
rect 3479 1709 3483 1710
rect 3575 1714 3579 1715
rect 3575 1709 3579 1710
rect 3016 1704 3018 1709
rect 3136 1704 3138 1709
rect 3248 1704 3250 1709
rect 3368 1704 3370 1709
rect 3480 1704 3482 1709
rect 3014 1703 3020 1704
rect 3014 1699 3015 1703
rect 3019 1699 3020 1703
rect 3014 1698 3020 1699
rect 3134 1703 3140 1704
rect 3134 1699 3135 1703
rect 3139 1699 3140 1703
rect 3134 1698 3140 1699
rect 3246 1703 3252 1704
rect 3246 1699 3247 1703
rect 3251 1699 3252 1703
rect 3246 1698 3252 1699
rect 3366 1703 3372 1704
rect 3366 1699 3367 1703
rect 3371 1699 3372 1703
rect 3366 1698 3372 1699
rect 3478 1703 3484 1704
rect 3478 1699 3479 1703
rect 3483 1699 3484 1703
rect 3478 1698 3484 1699
rect 3576 1694 3578 1709
rect 3574 1693 3580 1694
rect 3574 1689 3575 1693
rect 3579 1689 3580 1693
rect 3574 1688 3580 1689
rect 3126 1679 3132 1680
rect 3126 1675 3127 1679
rect 3131 1675 3132 1679
rect 3126 1674 3132 1675
rect 3574 1676 3580 1677
rect 3022 1663 3028 1664
rect 3022 1659 3023 1663
rect 3027 1659 3028 1663
rect 3022 1658 3028 1659
rect 2902 1651 2908 1652
rect 2902 1647 2903 1651
rect 2907 1647 2908 1651
rect 2902 1646 2908 1647
rect 3024 1643 3026 1658
rect 3128 1652 3130 1674
rect 3574 1672 3575 1676
rect 3579 1672 3580 1676
rect 3574 1671 3580 1672
rect 3142 1663 3148 1664
rect 3142 1659 3143 1663
rect 3147 1659 3148 1663
rect 3142 1658 3148 1659
rect 3254 1663 3260 1664
rect 3254 1659 3255 1663
rect 3259 1659 3260 1663
rect 3254 1658 3260 1659
rect 3374 1663 3380 1664
rect 3374 1659 3375 1663
rect 3379 1659 3380 1663
rect 3374 1658 3380 1659
rect 3486 1663 3492 1664
rect 3486 1659 3487 1663
rect 3491 1659 3492 1663
rect 3486 1658 3492 1659
rect 3126 1651 3132 1652
rect 3126 1647 3127 1651
rect 3131 1647 3132 1651
rect 3126 1646 3132 1647
rect 3098 1643 3104 1644
rect 3144 1643 3146 1658
rect 3256 1643 3258 1658
rect 3376 1643 3378 1658
rect 3488 1643 3490 1658
rect 3498 1651 3504 1652
rect 3498 1647 3499 1651
rect 3503 1647 3504 1651
rect 3498 1646 3504 1647
rect 1863 1642 1867 1643
rect 1183 1638 1187 1639
rect 1183 1633 1187 1634
rect 1303 1638 1307 1639
rect 1303 1633 1307 1634
rect 1351 1638 1355 1639
rect 1351 1633 1355 1634
rect 1455 1638 1459 1639
rect 1455 1633 1459 1634
rect 1519 1638 1523 1639
rect 1519 1633 1523 1634
rect 1599 1638 1603 1639
rect 1599 1633 1603 1634
rect 1687 1638 1691 1639
rect 1687 1633 1691 1634
rect 1727 1638 1731 1639
rect 1727 1633 1731 1634
rect 1823 1638 1827 1639
rect 1863 1637 1867 1638
rect 2151 1642 2155 1643
rect 2151 1637 2155 1638
rect 2255 1642 2259 1643
rect 2255 1637 2259 1638
rect 2343 1642 2347 1643
rect 2343 1637 2347 1638
rect 2375 1642 2379 1643
rect 2375 1637 2379 1638
rect 2503 1642 2507 1643
rect 2503 1637 2507 1638
rect 2527 1642 2531 1643
rect 2527 1637 2531 1638
rect 2631 1642 2635 1643
rect 2631 1637 2635 1638
rect 2703 1642 2707 1643
rect 2703 1637 2707 1638
rect 2767 1642 2771 1643
rect 2767 1637 2771 1638
rect 2871 1642 2875 1643
rect 2871 1637 2875 1638
rect 2895 1642 2899 1643
rect 2895 1637 2899 1638
rect 3023 1642 3027 1643
rect 3023 1637 3027 1638
rect 3031 1642 3035 1643
rect 3098 1639 3099 1643
rect 3103 1639 3104 1643
rect 3098 1638 3104 1639
rect 3143 1642 3147 1643
rect 3031 1637 3035 1638
rect 1823 1633 1827 1634
rect 1304 1628 1306 1633
rect 1456 1628 1458 1633
rect 1600 1628 1602 1633
rect 1728 1628 1730 1633
rect 1302 1627 1308 1628
rect 1302 1623 1303 1627
rect 1307 1623 1308 1627
rect 1302 1622 1308 1623
rect 1454 1627 1460 1628
rect 1454 1623 1455 1627
rect 1459 1623 1460 1627
rect 1454 1622 1460 1623
rect 1598 1627 1604 1628
rect 1598 1623 1599 1627
rect 1603 1623 1604 1627
rect 1598 1622 1604 1623
rect 1726 1627 1732 1628
rect 1726 1623 1727 1627
rect 1731 1623 1732 1627
rect 1726 1622 1732 1623
rect 1824 1618 1826 1633
rect 1822 1617 1828 1618
rect 1822 1613 1823 1617
rect 1827 1613 1828 1617
rect 1864 1613 1866 1637
rect 2152 1626 2154 1637
rect 2158 1635 2164 1636
rect 2158 1631 2159 1635
rect 2163 1631 2164 1635
rect 2158 1630 2164 1631
rect 2150 1625 2156 1626
rect 2150 1621 2151 1625
rect 2155 1621 2156 1625
rect 2150 1620 2156 1621
rect 1822 1612 1828 1613
rect 1862 1612 1868 1613
rect 1862 1608 1863 1612
rect 1867 1608 1868 1612
rect 1862 1607 1868 1608
rect 1582 1603 1588 1604
rect 1582 1599 1583 1603
rect 1587 1599 1588 1603
rect 1582 1598 1588 1599
rect 1666 1603 1672 1604
rect 1666 1599 1667 1603
rect 1671 1599 1672 1603
rect 1666 1598 1672 1599
rect 1822 1600 1828 1601
rect 1310 1587 1316 1588
rect 1310 1583 1311 1587
rect 1315 1583 1316 1587
rect 1310 1582 1316 1583
rect 1462 1587 1468 1588
rect 1462 1583 1463 1587
rect 1467 1583 1468 1587
rect 1462 1582 1468 1583
rect 1166 1575 1172 1576
rect 1166 1571 1167 1575
rect 1171 1571 1172 1575
rect 1312 1571 1314 1582
rect 1464 1571 1466 1582
rect 111 1570 115 1571
rect 134 1570 140 1571
rect 143 1570 147 1571
rect 111 1565 115 1566
rect 112 1541 114 1565
rect 110 1540 116 1541
rect 110 1536 111 1540
rect 115 1536 116 1540
rect 136 1536 138 1570
rect 143 1565 147 1566
rect 271 1570 275 1571
rect 271 1565 275 1566
rect 279 1570 283 1571
rect 286 1570 292 1571
rect 431 1570 435 1571
rect 279 1565 283 1566
rect 431 1565 435 1566
rect 455 1570 459 1571
rect 455 1565 459 1566
rect 599 1570 603 1571
rect 599 1565 603 1566
rect 639 1570 643 1571
rect 639 1565 643 1566
rect 767 1570 771 1571
rect 767 1565 771 1566
rect 823 1570 827 1571
rect 823 1565 827 1566
rect 935 1570 939 1571
rect 935 1565 939 1566
rect 999 1570 1003 1571
rect 1026 1570 1032 1571
rect 1103 1570 1107 1571
rect 999 1565 1003 1566
rect 144 1554 146 1565
rect 210 1563 216 1564
rect 210 1559 211 1563
rect 215 1559 216 1563
rect 210 1558 216 1559
rect 250 1563 256 1564
rect 250 1559 251 1563
rect 255 1559 256 1563
rect 250 1558 256 1559
rect 142 1553 148 1554
rect 142 1549 143 1553
rect 147 1549 148 1553
rect 142 1548 148 1549
rect 212 1536 214 1558
rect 110 1535 116 1536
rect 134 1535 140 1536
rect 134 1531 135 1535
rect 139 1531 140 1535
rect 134 1530 140 1531
rect 210 1535 216 1536
rect 210 1531 211 1535
rect 215 1531 216 1535
rect 210 1530 216 1531
rect 110 1523 116 1524
rect 110 1519 111 1523
rect 115 1519 116 1523
rect 110 1518 116 1519
rect 112 1499 114 1518
rect 134 1513 140 1514
rect 134 1509 135 1513
rect 139 1509 140 1513
rect 134 1508 140 1509
rect 136 1499 138 1508
rect 111 1498 115 1499
rect 111 1493 115 1494
rect 135 1498 139 1499
rect 135 1493 139 1494
rect 183 1498 187 1499
rect 183 1493 187 1494
rect 112 1478 114 1493
rect 184 1488 186 1493
rect 182 1487 188 1488
rect 182 1483 183 1487
rect 187 1483 188 1487
rect 182 1482 188 1483
rect 252 1480 254 1558
rect 272 1554 274 1565
rect 432 1554 434 1565
rect 514 1563 520 1564
rect 514 1559 515 1563
rect 519 1559 520 1563
rect 514 1558 520 1559
rect 270 1553 276 1554
rect 270 1549 271 1553
rect 275 1549 276 1553
rect 270 1548 276 1549
rect 430 1553 436 1554
rect 430 1549 431 1553
rect 435 1549 436 1553
rect 430 1548 436 1549
rect 516 1536 518 1558
rect 600 1554 602 1565
rect 666 1563 672 1564
rect 666 1559 667 1563
rect 671 1559 672 1563
rect 666 1558 672 1559
rect 598 1553 604 1554
rect 598 1549 599 1553
rect 603 1549 604 1553
rect 598 1548 604 1549
rect 668 1536 670 1558
rect 768 1554 770 1565
rect 936 1554 938 1565
rect 942 1563 948 1564
rect 942 1559 943 1563
rect 947 1559 948 1563
rect 942 1558 948 1559
rect 1018 1563 1024 1564
rect 1018 1559 1019 1563
rect 1023 1559 1024 1563
rect 1018 1558 1024 1559
rect 766 1553 772 1554
rect 766 1549 767 1553
rect 771 1549 772 1553
rect 766 1548 772 1549
rect 934 1553 940 1554
rect 934 1549 935 1553
rect 939 1549 940 1553
rect 934 1548 940 1549
rect 514 1535 520 1536
rect 514 1531 515 1535
rect 519 1531 520 1535
rect 514 1530 520 1531
rect 666 1535 672 1536
rect 666 1531 667 1535
rect 671 1531 672 1535
rect 666 1530 672 1531
rect 350 1523 356 1524
rect 350 1519 351 1523
rect 355 1519 356 1523
rect 350 1518 356 1519
rect 262 1513 268 1514
rect 262 1509 263 1513
rect 267 1509 268 1513
rect 262 1508 268 1509
rect 264 1499 266 1508
rect 263 1498 267 1499
rect 263 1493 267 1494
rect 327 1498 331 1499
rect 327 1493 331 1494
rect 328 1488 330 1493
rect 326 1487 332 1488
rect 326 1483 327 1487
rect 331 1483 332 1487
rect 326 1482 332 1483
rect 250 1479 256 1480
rect 110 1477 116 1478
rect 110 1473 111 1477
rect 115 1473 116 1477
rect 250 1475 251 1479
rect 255 1475 256 1479
rect 250 1474 256 1475
rect 110 1472 116 1473
rect 110 1460 116 1461
rect 110 1456 111 1460
rect 115 1456 116 1460
rect 110 1455 116 1456
rect 112 1423 114 1455
rect 190 1447 196 1448
rect 190 1443 191 1447
rect 195 1443 196 1447
rect 190 1442 196 1443
rect 334 1447 340 1448
rect 334 1443 335 1447
rect 339 1443 340 1447
rect 334 1442 340 1443
rect 182 1435 188 1436
rect 182 1431 183 1435
rect 187 1431 188 1435
rect 182 1430 188 1431
rect 111 1422 115 1423
rect 111 1417 115 1418
rect 112 1393 114 1417
rect 110 1392 116 1393
rect 110 1388 111 1392
rect 115 1388 116 1392
rect 184 1388 186 1430
rect 192 1423 194 1442
rect 336 1423 338 1442
rect 352 1436 354 1518
rect 422 1513 428 1514
rect 422 1509 423 1513
rect 427 1509 428 1513
rect 422 1508 428 1509
rect 590 1513 596 1514
rect 590 1509 591 1513
rect 595 1509 596 1513
rect 590 1508 596 1509
rect 758 1513 764 1514
rect 758 1509 759 1513
rect 763 1509 764 1513
rect 758 1508 764 1509
rect 926 1513 932 1514
rect 926 1509 927 1513
rect 931 1509 932 1513
rect 926 1508 932 1509
rect 424 1499 426 1508
rect 592 1499 594 1508
rect 760 1499 762 1508
rect 928 1499 930 1508
rect 423 1498 427 1499
rect 423 1493 427 1494
rect 471 1498 475 1499
rect 471 1493 475 1494
rect 591 1498 595 1499
rect 591 1493 595 1494
rect 607 1498 611 1499
rect 607 1493 611 1494
rect 743 1498 747 1499
rect 743 1493 747 1494
rect 759 1498 763 1499
rect 759 1493 763 1494
rect 871 1498 875 1499
rect 871 1493 875 1494
rect 927 1498 931 1499
rect 927 1493 931 1494
rect 472 1488 474 1493
rect 608 1488 610 1493
rect 744 1488 746 1493
rect 872 1488 874 1493
rect 470 1487 476 1488
rect 470 1483 471 1487
rect 475 1483 476 1487
rect 470 1482 476 1483
rect 606 1487 612 1488
rect 606 1483 607 1487
rect 611 1483 612 1487
rect 606 1482 612 1483
rect 742 1487 748 1488
rect 742 1483 743 1487
rect 747 1483 748 1487
rect 742 1482 748 1483
rect 870 1487 876 1488
rect 870 1483 871 1487
rect 875 1483 876 1487
rect 870 1482 876 1483
rect 944 1480 946 1558
rect 1020 1540 1022 1558
rect 1018 1539 1024 1540
rect 1018 1535 1019 1539
rect 1023 1535 1024 1539
rect 1028 1536 1030 1570
rect 1103 1565 1107 1566
rect 1159 1570 1163 1571
rect 1166 1570 1172 1571
rect 1263 1570 1267 1571
rect 1159 1565 1163 1566
rect 1263 1565 1267 1566
rect 1311 1570 1315 1571
rect 1311 1565 1315 1566
rect 1423 1570 1427 1571
rect 1423 1565 1427 1566
rect 1463 1570 1467 1571
rect 1463 1565 1467 1566
rect 1104 1554 1106 1565
rect 1264 1554 1266 1565
rect 1342 1563 1348 1564
rect 1342 1559 1343 1563
rect 1347 1559 1348 1563
rect 1342 1558 1348 1559
rect 1102 1553 1108 1554
rect 1102 1549 1103 1553
rect 1107 1549 1108 1553
rect 1102 1548 1108 1549
rect 1262 1553 1268 1554
rect 1262 1549 1263 1553
rect 1267 1549 1268 1553
rect 1262 1548 1268 1549
rect 1344 1540 1346 1558
rect 1424 1554 1426 1565
rect 1584 1564 1586 1598
rect 1606 1587 1612 1588
rect 1606 1583 1607 1587
rect 1611 1583 1612 1587
rect 1606 1582 1612 1583
rect 1608 1571 1610 1582
rect 1668 1576 1670 1598
rect 1822 1596 1823 1600
rect 1827 1596 1828 1600
rect 1822 1595 1828 1596
rect 1862 1595 1868 1596
rect 1734 1587 1740 1588
rect 1734 1583 1735 1587
rect 1739 1583 1740 1587
rect 1734 1582 1740 1583
rect 1666 1575 1672 1576
rect 1666 1571 1667 1575
rect 1671 1571 1672 1575
rect 1736 1571 1738 1582
rect 1824 1571 1826 1595
rect 1862 1591 1863 1595
rect 1867 1591 1868 1595
rect 1862 1590 1868 1591
rect 1864 1575 1866 1590
rect 2142 1585 2148 1586
rect 2142 1581 2143 1585
rect 2147 1581 2148 1585
rect 2142 1580 2148 1581
rect 2144 1575 2146 1580
rect 1863 1574 1867 1575
rect 1591 1570 1595 1571
rect 1591 1565 1595 1566
rect 1607 1570 1611 1571
rect 1666 1570 1672 1571
rect 1735 1570 1739 1571
rect 1607 1565 1611 1566
rect 1735 1565 1739 1566
rect 1823 1570 1827 1571
rect 1863 1569 1867 1570
rect 2087 1574 2091 1575
rect 2143 1574 2147 1575
rect 2087 1569 2091 1570
rect 2102 1571 2108 1572
rect 1823 1565 1827 1566
rect 1582 1563 1588 1564
rect 1582 1559 1583 1563
rect 1587 1559 1588 1563
rect 1582 1558 1588 1559
rect 1592 1554 1594 1565
rect 1662 1563 1668 1564
rect 1662 1559 1663 1563
rect 1667 1559 1668 1563
rect 1662 1558 1668 1559
rect 1422 1553 1428 1554
rect 1422 1549 1423 1553
rect 1427 1549 1428 1553
rect 1422 1548 1428 1549
rect 1590 1553 1596 1554
rect 1590 1549 1591 1553
rect 1595 1549 1596 1553
rect 1590 1548 1596 1549
rect 1664 1540 1666 1558
rect 1736 1554 1738 1565
rect 1734 1553 1740 1554
rect 1734 1549 1735 1553
rect 1739 1549 1740 1553
rect 1734 1548 1740 1549
rect 1824 1541 1826 1565
rect 1864 1554 1866 1569
rect 2088 1564 2090 1569
rect 2102 1567 2103 1571
rect 2107 1567 2108 1571
rect 2143 1569 2147 1570
rect 2102 1566 2108 1567
rect 2086 1563 2092 1564
rect 2086 1559 2087 1563
rect 2091 1559 2092 1563
rect 2086 1558 2092 1559
rect 1862 1553 1868 1554
rect 1862 1549 1863 1553
rect 1867 1549 1868 1553
rect 1862 1548 1868 1549
rect 1822 1540 1828 1541
rect 1342 1539 1348 1540
rect 1018 1534 1024 1535
rect 1026 1535 1032 1536
rect 1026 1531 1027 1535
rect 1031 1531 1032 1535
rect 1342 1535 1343 1539
rect 1347 1535 1348 1539
rect 1342 1534 1348 1535
rect 1662 1539 1668 1540
rect 1662 1535 1663 1539
rect 1667 1535 1668 1539
rect 1822 1536 1823 1540
rect 1827 1536 1828 1540
rect 1822 1535 1828 1536
rect 1862 1536 1868 1537
rect 1662 1534 1668 1535
rect 1862 1532 1863 1536
rect 1867 1532 1868 1536
rect 1862 1531 1868 1532
rect 1026 1530 1032 1531
rect 1390 1523 1396 1524
rect 1390 1519 1391 1523
rect 1395 1519 1396 1523
rect 1390 1518 1396 1519
rect 1814 1523 1820 1524
rect 1814 1519 1815 1523
rect 1819 1519 1820 1523
rect 1814 1518 1820 1519
rect 1822 1523 1828 1524
rect 1822 1519 1823 1523
rect 1827 1519 1828 1523
rect 1822 1518 1828 1519
rect 1094 1513 1100 1514
rect 1094 1509 1095 1513
rect 1099 1509 1100 1513
rect 1094 1508 1100 1509
rect 1254 1513 1260 1514
rect 1254 1509 1255 1513
rect 1259 1509 1260 1513
rect 1254 1508 1260 1509
rect 1096 1499 1098 1508
rect 1256 1499 1258 1508
rect 991 1498 995 1499
rect 991 1493 995 1494
rect 1095 1498 1099 1499
rect 1095 1493 1099 1494
rect 1119 1498 1123 1499
rect 1119 1493 1123 1494
rect 1247 1498 1251 1499
rect 1247 1493 1251 1494
rect 1255 1498 1259 1499
rect 1255 1493 1259 1494
rect 1375 1498 1379 1499
rect 1375 1493 1379 1494
rect 992 1488 994 1493
rect 1120 1488 1122 1493
rect 1248 1488 1250 1493
rect 1376 1488 1378 1493
rect 990 1487 996 1488
rect 990 1483 991 1487
rect 995 1483 996 1487
rect 990 1482 996 1483
rect 1118 1487 1124 1488
rect 1118 1483 1119 1487
rect 1123 1483 1124 1487
rect 1118 1482 1124 1483
rect 1246 1487 1252 1488
rect 1246 1483 1247 1487
rect 1251 1483 1252 1487
rect 1246 1482 1252 1483
rect 1374 1487 1380 1488
rect 1374 1483 1375 1487
rect 1379 1483 1380 1487
rect 1374 1482 1380 1483
rect 942 1479 948 1480
rect 942 1475 943 1479
rect 947 1475 948 1479
rect 942 1474 948 1475
rect 938 1463 944 1464
rect 938 1459 939 1463
rect 943 1459 944 1463
rect 938 1458 944 1459
rect 1058 1463 1064 1464
rect 1058 1459 1059 1463
rect 1063 1459 1064 1463
rect 1058 1458 1064 1459
rect 1314 1463 1320 1464
rect 1314 1459 1315 1463
rect 1319 1459 1320 1463
rect 1314 1458 1320 1459
rect 478 1447 484 1448
rect 478 1443 479 1447
rect 483 1443 484 1447
rect 478 1442 484 1443
rect 614 1447 620 1448
rect 614 1443 615 1447
rect 619 1443 620 1447
rect 614 1442 620 1443
rect 750 1447 756 1448
rect 750 1443 751 1447
rect 755 1443 756 1447
rect 750 1442 756 1443
rect 878 1447 884 1448
rect 878 1443 879 1447
rect 883 1443 884 1447
rect 878 1442 884 1443
rect 350 1435 356 1436
rect 350 1431 351 1435
rect 355 1431 356 1435
rect 350 1430 356 1431
rect 480 1423 482 1442
rect 616 1423 618 1442
rect 658 1423 664 1424
rect 752 1423 754 1442
rect 880 1423 882 1442
rect 940 1436 942 1458
rect 998 1447 1004 1448
rect 998 1443 999 1447
rect 1003 1443 1004 1447
rect 998 1442 1004 1443
rect 938 1435 944 1436
rect 938 1431 939 1435
rect 943 1431 944 1435
rect 938 1430 944 1431
rect 1000 1423 1002 1442
rect 1060 1436 1062 1458
rect 1126 1447 1132 1448
rect 1126 1443 1127 1447
rect 1131 1443 1132 1447
rect 1126 1442 1132 1443
rect 1254 1447 1260 1448
rect 1254 1443 1255 1447
rect 1259 1443 1260 1447
rect 1254 1442 1260 1443
rect 1058 1435 1064 1436
rect 1058 1431 1059 1435
rect 1063 1431 1064 1435
rect 1058 1430 1064 1431
rect 1110 1435 1116 1436
rect 1110 1431 1111 1435
rect 1115 1431 1116 1435
rect 1110 1430 1116 1431
rect 191 1422 195 1423
rect 191 1417 195 1418
rect 199 1422 203 1423
rect 199 1417 203 1418
rect 335 1422 339 1423
rect 335 1417 339 1418
rect 463 1422 467 1423
rect 463 1417 467 1418
rect 479 1422 483 1423
rect 479 1417 483 1418
rect 583 1422 587 1423
rect 583 1417 587 1418
rect 615 1422 619 1423
rect 658 1419 659 1423
rect 663 1419 664 1423
rect 658 1418 664 1419
rect 703 1422 707 1423
rect 615 1417 619 1418
rect 200 1406 202 1417
rect 270 1415 276 1416
rect 270 1411 271 1415
rect 275 1411 276 1415
rect 270 1410 276 1411
rect 298 1415 304 1416
rect 298 1411 299 1415
rect 303 1411 304 1415
rect 298 1410 304 1411
rect 198 1405 204 1406
rect 198 1401 199 1405
rect 203 1401 204 1405
rect 198 1400 204 1401
rect 272 1388 274 1410
rect 110 1387 116 1388
rect 182 1387 188 1388
rect 182 1383 183 1387
rect 187 1383 188 1387
rect 182 1382 188 1383
rect 270 1387 276 1388
rect 270 1383 271 1387
rect 275 1383 276 1387
rect 270 1382 276 1383
rect 110 1375 116 1376
rect 110 1371 111 1375
rect 115 1371 116 1375
rect 110 1370 116 1371
rect 112 1351 114 1370
rect 190 1365 196 1366
rect 190 1361 191 1365
rect 195 1361 196 1365
rect 190 1360 196 1361
rect 192 1351 194 1360
rect 111 1350 115 1351
rect 111 1345 115 1346
rect 191 1350 195 1351
rect 191 1345 195 1346
rect 231 1350 235 1351
rect 231 1345 235 1346
rect 112 1330 114 1345
rect 232 1340 234 1345
rect 230 1339 236 1340
rect 230 1335 231 1339
rect 235 1335 236 1339
rect 230 1334 236 1335
rect 300 1332 302 1410
rect 336 1406 338 1417
rect 464 1406 466 1417
rect 584 1406 586 1417
rect 334 1405 340 1406
rect 334 1401 335 1405
rect 339 1401 340 1405
rect 334 1400 340 1401
rect 462 1405 468 1406
rect 462 1401 463 1405
rect 467 1401 468 1405
rect 462 1400 468 1401
rect 582 1405 588 1406
rect 582 1401 583 1405
rect 587 1401 588 1405
rect 582 1400 588 1401
rect 660 1388 662 1418
rect 703 1417 707 1418
rect 751 1422 755 1423
rect 751 1417 755 1418
rect 815 1422 819 1423
rect 815 1417 819 1418
rect 879 1422 883 1423
rect 879 1417 883 1418
rect 919 1422 923 1423
rect 919 1417 923 1418
rect 999 1422 1003 1423
rect 999 1417 1003 1418
rect 1015 1422 1019 1423
rect 1015 1417 1019 1418
rect 704 1406 706 1417
rect 770 1415 776 1416
rect 770 1411 771 1415
rect 775 1411 776 1415
rect 770 1410 776 1411
rect 702 1405 708 1406
rect 702 1401 703 1405
rect 707 1401 708 1405
rect 702 1400 708 1401
rect 658 1387 664 1388
rect 658 1383 659 1387
rect 663 1383 664 1387
rect 658 1382 664 1383
rect 326 1365 332 1366
rect 326 1361 327 1365
rect 331 1361 332 1365
rect 326 1360 332 1361
rect 454 1365 460 1366
rect 454 1361 455 1365
rect 459 1361 460 1365
rect 454 1360 460 1361
rect 574 1365 580 1366
rect 574 1361 575 1365
rect 579 1361 580 1365
rect 574 1360 580 1361
rect 694 1365 700 1366
rect 694 1361 695 1365
rect 699 1361 700 1365
rect 694 1360 700 1361
rect 328 1351 330 1360
rect 456 1351 458 1360
rect 576 1351 578 1360
rect 696 1351 698 1360
rect 327 1350 331 1351
rect 327 1345 331 1346
rect 383 1350 387 1351
rect 383 1345 387 1346
rect 455 1350 459 1351
rect 455 1345 459 1346
rect 543 1350 547 1351
rect 543 1345 547 1346
rect 575 1350 579 1351
rect 575 1345 579 1346
rect 695 1350 699 1351
rect 695 1345 699 1346
rect 703 1350 707 1351
rect 703 1345 707 1346
rect 384 1340 386 1345
rect 544 1340 546 1345
rect 704 1340 706 1345
rect 382 1339 388 1340
rect 382 1335 383 1339
rect 387 1335 388 1339
rect 382 1334 388 1335
rect 542 1339 548 1340
rect 542 1335 543 1339
rect 547 1335 548 1339
rect 542 1334 548 1335
rect 702 1339 708 1340
rect 702 1335 703 1339
rect 707 1335 708 1339
rect 702 1334 708 1335
rect 772 1332 774 1410
rect 816 1406 818 1417
rect 920 1406 922 1417
rect 1016 1406 1018 1417
rect 814 1405 820 1406
rect 814 1401 815 1405
rect 819 1401 820 1405
rect 814 1400 820 1401
rect 918 1405 924 1406
rect 918 1401 919 1405
rect 923 1401 924 1405
rect 918 1400 924 1401
rect 1014 1405 1020 1406
rect 1014 1401 1015 1405
rect 1019 1401 1020 1405
rect 1014 1400 1020 1401
rect 1112 1388 1114 1430
rect 1128 1423 1130 1442
rect 1256 1423 1258 1442
rect 1316 1436 1318 1458
rect 1382 1447 1388 1448
rect 1382 1443 1383 1447
rect 1387 1443 1388 1447
rect 1382 1442 1388 1443
rect 1314 1435 1320 1436
rect 1314 1431 1315 1435
rect 1319 1431 1320 1435
rect 1314 1430 1320 1431
rect 1384 1423 1386 1442
rect 1392 1436 1394 1518
rect 1414 1513 1420 1514
rect 1414 1509 1415 1513
rect 1419 1509 1420 1513
rect 1414 1508 1420 1509
rect 1582 1513 1588 1514
rect 1582 1509 1583 1513
rect 1587 1509 1588 1513
rect 1582 1508 1588 1509
rect 1726 1513 1732 1514
rect 1726 1509 1727 1513
rect 1731 1509 1732 1513
rect 1726 1508 1732 1509
rect 1416 1499 1418 1508
rect 1584 1499 1586 1508
rect 1728 1499 1730 1508
rect 1415 1498 1419 1499
rect 1415 1493 1419 1494
rect 1583 1498 1587 1499
rect 1583 1493 1587 1494
rect 1727 1498 1731 1499
rect 1727 1493 1731 1494
rect 1816 1492 1818 1518
rect 1824 1499 1826 1518
rect 1864 1499 1866 1531
rect 2094 1523 2100 1524
rect 2094 1519 2095 1523
rect 2099 1519 2100 1523
rect 2094 1518 2100 1519
rect 2096 1499 2098 1518
rect 2104 1512 2106 1566
rect 2160 1556 2162 1630
rect 2344 1626 2346 1637
rect 2528 1626 2530 1637
rect 2704 1626 2706 1637
rect 2872 1626 2874 1637
rect 3032 1626 3034 1637
rect 2342 1625 2348 1626
rect 2342 1621 2343 1625
rect 2347 1621 2348 1625
rect 2342 1620 2348 1621
rect 2526 1625 2532 1626
rect 2526 1621 2527 1625
rect 2531 1621 2532 1625
rect 2526 1620 2532 1621
rect 2702 1625 2708 1626
rect 2702 1621 2703 1625
rect 2707 1621 2708 1625
rect 2702 1620 2708 1621
rect 2870 1625 2876 1626
rect 2870 1621 2871 1625
rect 2875 1621 2876 1625
rect 2870 1620 2876 1621
rect 3030 1625 3036 1626
rect 3030 1621 3031 1625
rect 3035 1621 3036 1625
rect 3030 1620 3036 1621
rect 3100 1608 3102 1638
rect 3143 1637 3147 1638
rect 3191 1642 3195 1643
rect 3191 1637 3195 1638
rect 3255 1642 3259 1643
rect 3255 1637 3259 1638
rect 3351 1642 3355 1643
rect 3351 1637 3355 1638
rect 3375 1642 3379 1643
rect 3375 1637 3379 1638
rect 3487 1642 3491 1643
rect 3487 1637 3491 1638
rect 3192 1626 3194 1637
rect 3352 1626 3354 1637
rect 3488 1626 3490 1637
rect 3190 1625 3196 1626
rect 3190 1621 3191 1625
rect 3195 1621 3196 1625
rect 3190 1620 3196 1621
rect 3350 1625 3356 1626
rect 3350 1621 3351 1625
rect 3355 1621 3356 1625
rect 3350 1620 3356 1621
rect 3486 1625 3492 1626
rect 3486 1621 3487 1625
rect 3491 1621 3492 1625
rect 3486 1620 3492 1621
rect 3098 1607 3104 1608
rect 3098 1603 3099 1607
rect 3103 1603 3104 1607
rect 3098 1602 3104 1603
rect 3470 1595 3476 1596
rect 3470 1591 3471 1595
rect 3475 1591 3476 1595
rect 3470 1590 3476 1591
rect 2334 1585 2340 1586
rect 2334 1581 2335 1585
rect 2339 1581 2340 1585
rect 2334 1580 2340 1581
rect 2518 1585 2524 1586
rect 2518 1581 2519 1585
rect 2523 1581 2524 1585
rect 2518 1580 2524 1581
rect 2694 1585 2700 1586
rect 2694 1581 2695 1585
rect 2699 1581 2700 1585
rect 2694 1580 2700 1581
rect 2862 1585 2868 1586
rect 2862 1581 2863 1585
rect 2867 1581 2868 1585
rect 2862 1580 2868 1581
rect 3022 1585 3028 1586
rect 3022 1581 3023 1585
rect 3027 1581 3028 1585
rect 3022 1580 3028 1581
rect 3182 1585 3188 1586
rect 3182 1581 3183 1585
rect 3187 1581 3188 1585
rect 3182 1580 3188 1581
rect 3342 1585 3348 1586
rect 3342 1581 3343 1585
rect 3347 1581 3348 1585
rect 3342 1580 3348 1581
rect 2336 1575 2338 1580
rect 2520 1575 2522 1580
rect 2696 1575 2698 1580
rect 2864 1575 2866 1580
rect 3024 1575 3026 1580
rect 3184 1575 3186 1580
rect 3344 1575 3346 1580
rect 2279 1574 2283 1575
rect 2279 1569 2283 1570
rect 2335 1574 2339 1575
rect 2335 1569 2339 1570
rect 2455 1574 2459 1575
rect 2455 1569 2459 1570
rect 2519 1574 2523 1575
rect 2519 1569 2523 1570
rect 2623 1574 2627 1575
rect 2623 1569 2627 1570
rect 2695 1574 2699 1575
rect 2695 1569 2699 1570
rect 2791 1574 2795 1575
rect 2791 1569 2795 1570
rect 2863 1574 2867 1575
rect 2863 1569 2867 1570
rect 2951 1574 2955 1575
rect 2951 1569 2955 1570
rect 3023 1574 3027 1575
rect 3023 1569 3027 1570
rect 3111 1574 3115 1575
rect 3111 1569 3115 1570
rect 3183 1574 3187 1575
rect 3183 1569 3187 1570
rect 3271 1574 3275 1575
rect 3271 1569 3275 1570
rect 3343 1574 3347 1575
rect 3343 1569 3347 1570
rect 3431 1574 3435 1575
rect 3431 1569 3435 1570
rect 2280 1564 2282 1569
rect 2456 1564 2458 1569
rect 2624 1564 2626 1569
rect 2792 1564 2794 1569
rect 2952 1564 2954 1569
rect 3112 1564 3114 1569
rect 3272 1564 3274 1569
rect 3432 1564 3434 1569
rect 2278 1563 2284 1564
rect 2278 1559 2279 1563
rect 2283 1559 2284 1563
rect 2278 1558 2284 1559
rect 2454 1563 2460 1564
rect 2454 1559 2455 1563
rect 2459 1559 2460 1563
rect 2454 1558 2460 1559
rect 2622 1563 2628 1564
rect 2622 1559 2623 1563
rect 2627 1559 2628 1563
rect 2622 1558 2628 1559
rect 2790 1563 2796 1564
rect 2790 1559 2791 1563
rect 2795 1559 2796 1563
rect 2790 1558 2796 1559
rect 2950 1563 2956 1564
rect 2950 1559 2951 1563
rect 2955 1559 2956 1563
rect 2950 1558 2956 1559
rect 3110 1563 3116 1564
rect 3110 1559 3111 1563
rect 3115 1559 3116 1563
rect 3110 1558 3116 1559
rect 3270 1563 3276 1564
rect 3270 1559 3271 1563
rect 3275 1559 3276 1563
rect 3270 1558 3276 1559
rect 3430 1563 3436 1564
rect 3430 1559 3431 1563
rect 3435 1559 3436 1563
rect 3430 1558 3436 1559
rect 2158 1555 2164 1556
rect 2158 1551 2159 1555
rect 2163 1551 2164 1555
rect 2158 1550 2164 1551
rect 3214 1555 3220 1556
rect 3214 1551 3215 1555
rect 3219 1551 3220 1555
rect 3214 1550 3220 1551
rect 3078 1539 3084 1540
rect 3078 1535 3079 1539
rect 3083 1535 3084 1539
rect 3078 1534 3084 1535
rect 2286 1523 2292 1524
rect 2286 1519 2287 1523
rect 2291 1519 2292 1523
rect 2286 1518 2292 1519
rect 2462 1523 2468 1524
rect 2462 1519 2463 1523
rect 2467 1519 2468 1523
rect 2462 1518 2468 1519
rect 2630 1523 2636 1524
rect 2630 1519 2631 1523
rect 2635 1519 2636 1523
rect 2630 1518 2636 1519
rect 2798 1523 2804 1524
rect 2798 1519 2799 1523
rect 2803 1519 2804 1523
rect 2798 1518 2804 1519
rect 2958 1523 2964 1524
rect 2958 1519 2959 1523
rect 2963 1519 2964 1523
rect 2958 1518 2964 1519
rect 2102 1511 2108 1512
rect 2102 1507 2103 1511
rect 2107 1507 2108 1511
rect 2102 1506 2108 1507
rect 2178 1511 2184 1512
rect 2178 1507 2179 1511
rect 2183 1507 2184 1511
rect 2178 1506 2184 1507
rect 1823 1498 1827 1499
rect 1823 1493 1827 1494
rect 1863 1498 1867 1499
rect 1863 1493 1867 1494
rect 1895 1498 1899 1499
rect 1895 1493 1899 1494
rect 1991 1498 1995 1499
rect 1991 1493 1995 1494
rect 2095 1498 2099 1499
rect 2095 1493 2099 1494
rect 2119 1498 2123 1499
rect 2119 1493 2123 1494
rect 1814 1491 1820 1492
rect 1814 1487 1815 1491
rect 1819 1487 1820 1491
rect 1814 1486 1820 1487
rect 1824 1478 1826 1493
rect 1822 1477 1828 1478
rect 1822 1473 1823 1477
rect 1827 1473 1828 1477
rect 1822 1472 1828 1473
rect 1864 1469 1866 1493
rect 1896 1482 1898 1493
rect 1992 1482 1994 1493
rect 2120 1482 2122 1493
rect 1894 1481 1900 1482
rect 1894 1477 1895 1481
rect 1899 1477 1900 1481
rect 1894 1476 1900 1477
rect 1990 1481 1996 1482
rect 1990 1477 1991 1481
rect 1995 1477 1996 1481
rect 1990 1476 1996 1477
rect 2118 1481 2124 1482
rect 2118 1477 2119 1481
rect 2123 1477 2124 1481
rect 2118 1476 2124 1477
rect 1862 1468 1868 1469
rect 2180 1468 2182 1506
rect 2288 1499 2290 1518
rect 2464 1499 2466 1518
rect 2632 1499 2634 1518
rect 2639 1516 2643 1517
rect 2638 1511 2644 1512
rect 2638 1507 2639 1511
rect 2643 1507 2644 1511
rect 2638 1506 2644 1507
rect 2778 1499 2784 1500
rect 2800 1499 2802 1518
rect 2960 1499 2962 1518
rect 2247 1498 2251 1499
rect 2247 1493 2251 1494
rect 2287 1498 2291 1499
rect 2287 1493 2291 1494
rect 2383 1498 2387 1499
rect 2383 1493 2387 1494
rect 2463 1498 2467 1499
rect 2463 1493 2467 1494
rect 2535 1498 2539 1499
rect 2535 1493 2539 1494
rect 2631 1498 2635 1499
rect 2631 1493 2635 1494
rect 2703 1498 2707 1499
rect 2778 1495 2779 1499
rect 2783 1495 2784 1499
rect 2778 1494 2784 1495
rect 2799 1498 2803 1499
rect 2703 1493 2707 1494
rect 2186 1491 2192 1492
rect 2186 1487 2187 1491
rect 2191 1487 2192 1491
rect 2186 1486 2192 1487
rect 1862 1464 1863 1468
rect 1867 1464 1868 1468
rect 1862 1463 1868 1464
rect 2178 1467 2184 1468
rect 2178 1463 2179 1467
rect 2183 1463 2184 1467
rect 2188 1464 2190 1486
rect 2248 1482 2250 1493
rect 2384 1482 2386 1493
rect 2390 1491 2396 1492
rect 2390 1487 2391 1491
rect 2395 1487 2396 1491
rect 2390 1486 2396 1487
rect 2246 1481 2252 1482
rect 2246 1477 2247 1481
rect 2251 1477 2252 1481
rect 2246 1476 2252 1477
rect 2382 1481 2388 1482
rect 2382 1477 2383 1481
rect 2387 1477 2388 1481
rect 2382 1476 2388 1477
rect 2178 1462 2184 1463
rect 2186 1463 2192 1464
rect 1822 1460 1828 1461
rect 1822 1456 1823 1460
rect 1827 1456 1828 1460
rect 2186 1459 2187 1463
rect 2191 1459 2192 1463
rect 2186 1458 2192 1459
rect 1822 1455 1828 1456
rect 1390 1435 1396 1436
rect 1390 1431 1391 1435
rect 1395 1431 1396 1435
rect 1390 1430 1396 1431
rect 1824 1423 1826 1455
rect 1862 1451 1868 1452
rect 1862 1447 1863 1451
rect 1867 1447 1868 1451
rect 1862 1446 1868 1447
rect 1864 1427 1866 1446
rect 1886 1441 1892 1442
rect 1886 1437 1887 1441
rect 1891 1437 1892 1441
rect 1886 1436 1892 1437
rect 1982 1441 1988 1442
rect 1982 1437 1983 1441
rect 1987 1437 1988 1441
rect 1982 1436 1988 1437
rect 2110 1441 2116 1442
rect 2110 1437 2111 1441
rect 2115 1437 2116 1441
rect 2110 1436 2116 1437
rect 2238 1441 2244 1442
rect 2238 1437 2239 1441
rect 2243 1437 2244 1441
rect 2238 1436 2244 1437
rect 2374 1441 2380 1442
rect 2374 1437 2375 1441
rect 2379 1437 2380 1441
rect 2374 1436 2380 1437
rect 1888 1427 1890 1436
rect 1984 1427 1986 1436
rect 2112 1427 2114 1436
rect 2240 1427 2242 1436
rect 2376 1427 2378 1436
rect 1863 1426 1867 1427
rect 1119 1422 1123 1423
rect 1119 1417 1123 1418
rect 1127 1422 1131 1423
rect 1127 1417 1131 1418
rect 1223 1422 1227 1423
rect 1223 1417 1227 1418
rect 1255 1422 1259 1423
rect 1255 1417 1259 1418
rect 1327 1422 1331 1423
rect 1327 1417 1331 1418
rect 1383 1422 1387 1423
rect 1383 1417 1387 1418
rect 1823 1422 1827 1423
rect 1863 1421 1867 1422
rect 1887 1426 1891 1427
rect 1887 1421 1891 1422
rect 1975 1426 1979 1427
rect 1975 1421 1979 1422
rect 1983 1426 1987 1427
rect 1983 1421 1987 1422
rect 2071 1426 2075 1427
rect 2071 1421 2075 1422
rect 2111 1426 2115 1427
rect 2111 1421 2115 1422
rect 2183 1426 2187 1427
rect 2183 1421 2187 1422
rect 2239 1426 2243 1427
rect 2239 1421 2243 1422
rect 2303 1426 2307 1427
rect 2303 1421 2307 1422
rect 2375 1426 2379 1427
rect 2375 1421 2379 1422
rect 1823 1417 1827 1418
rect 1120 1406 1122 1417
rect 1224 1406 1226 1417
rect 1328 1406 1330 1417
rect 1118 1405 1124 1406
rect 1118 1401 1119 1405
rect 1123 1401 1124 1405
rect 1118 1400 1124 1401
rect 1222 1405 1228 1406
rect 1222 1401 1223 1405
rect 1227 1401 1228 1405
rect 1222 1400 1228 1401
rect 1326 1405 1332 1406
rect 1326 1401 1327 1405
rect 1331 1401 1332 1405
rect 1326 1400 1332 1401
rect 1824 1393 1826 1417
rect 1864 1406 1866 1421
rect 1888 1416 1890 1421
rect 1976 1416 1978 1421
rect 2072 1416 2074 1421
rect 2184 1416 2186 1421
rect 2304 1416 2306 1421
rect 1886 1415 1892 1416
rect 1886 1411 1887 1415
rect 1891 1411 1892 1415
rect 1886 1410 1892 1411
rect 1974 1415 1980 1416
rect 1974 1411 1975 1415
rect 1979 1411 1980 1415
rect 1974 1410 1980 1411
rect 2070 1415 2076 1416
rect 2070 1411 2071 1415
rect 2075 1411 2076 1415
rect 2070 1410 2076 1411
rect 2182 1415 2188 1416
rect 2182 1411 2183 1415
rect 2187 1411 2188 1415
rect 2182 1410 2188 1411
rect 2302 1415 2308 1416
rect 2302 1411 2303 1415
rect 2307 1411 2308 1415
rect 2302 1410 2308 1411
rect 2392 1408 2394 1486
rect 2536 1482 2538 1493
rect 2704 1482 2706 1493
rect 2534 1481 2540 1482
rect 2534 1477 2535 1481
rect 2539 1477 2540 1481
rect 2534 1476 2540 1477
rect 2702 1481 2708 1482
rect 2702 1477 2703 1481
rect 2707 1477 2708 1481
rect 2702 1476 2708 1477
rect 2780 1464 2782 1494
rect 2799 1493 2803 1494
rect 2887 1498 2891 1499
rect 2887 1493 2891 1494
rect 2959 1498 2963 1499
rect 2959 1493 2963 1494
rect 2888 1482 2890 1493
rect 3080 1492 3082 1534
rect 3118 1523 3124 1524
rect 3118 1519 3119 1523
rect 3123 1519 3124 1523
rect 3118 1518 3124 1519
rect 3120 1499 3122 1518
rect 3216 1517 3218 1550
rect 3278 1523 3284 1524
rect 3278 1519 3279 1523
rect 3283 1519 3284 1523
rect 3278 1518 3284 1519
rect 3438 1523 3444 1524
rect 3438 1519 3439 1523
rect 3443 1519 3444 1523
rect 3438 1518 3444 1519
rect 3215 1516 3219 1517
rect 3215 1511 3219 1512
rect 3218 1499 3224 1500
rect 3280 1499 3282 1518
rect 3440 1499 3442 1518
rect 3087 1498 3091 1499
rect 3087 1493 3091 1494
rect 3119 1498 3123 1499
rect 3218 1495 3219 1499
rect 3223 1495 3224 1499
rect 3218 1494 3224 1495
rect 3279 1498 3283 1499
rect 3119 1493 3123 1494
rect 3078 1491 3084 1492
rect 3078 1487 3079 1491
rect 3083 1487 3084 1491
rect 3078 1486 3084 1487
rect 3088 1482 3090 1493
rect 2886 1481 2892 1482
rect 2886 1477 2887 1481
rect 2891 1477 2892 1481
rect 2886 1476 2892 1477
rect 3086 1481 3092 1482
rect 3086 1477 3087 1481
rect 3091 1477 3092 1481
rect 3086 1476 3092 1477
rect 3220 1464 3222 1494
rect 3279 1493 3283 1494
rect 3295 1498 3299 1499
rect 3295 1493 3299 1494
rect 3439 1498 3443 1499
rect 3439 1493 3443 1494
rect 3296 1482 3298 1493
rect 3472 1492 3474 1590
rect 3478 1585 3484 1586
rect 3478 1581 3479 1585
rect 3483 1581 3484 1585
rect 3478 1580 3484 1581
rect 3480 1575 3482 1580
rect 3479 1574 3483 1575
rect 3479 1569 3483 1570
rect 3500 1556 3502 1646
rect 3576 1643 3578 1671
rect 3575 1642 3579 1643
rect 3575 1637 3579 1638
rect 3576 1613 3578 1637
rect 3574 1612 3580 1613
rect 3574 1608 3575 1612
rect 3579 1608 3580 1612
rect 3574 1607 3580 1608
rect 3574 1595 3580 1596
rect 3574 1591 3575 1595
rect 3579 1591 3580 1595
rect 3574 1590 3580 1591
rect 3576 1575 3578 1590
rect 3575 1574 3579 1575
rect 3575 1569 3579 1570
rect 3498 1555 3504 1556
rect 3498 1551 3499 1555
rect 3503 1551 3504 1555
rect 3576 1554 3578 1569
rect 3498 1550 3504 1551
rect 3574 1553 3580 1554
rect 3574 1549 3575 1553
rect 3579 1549 3580 1553
rect 3574 1548 3580 1549
rect 3574 1536 3580 1537
rect 3574 1532 3575 1536
rect 3579 1532 3580 1536
rect 3574 1531 3580 1532
rect 3576 1499 3578 1531
rect 3487 1498 3491 1499
rect 3487 1493 3491 1494
rect 3575 1498 3579 1499
rect 3575 1493 3579 1494
rect 3470 1491 3476 1492
rect 3470 1487 3471 1491
rect 3475 1487 3476 1491
rect 3470 1486 3476 1487
rect 3488 1482 3490 1493
rect 3294 1481 3300 1482
rect 3294 1477 3295 1481
rect 3299 1477 3300 1481
rect 3294 1476 3300 1477
rect 3486 1481 3492 1482
rect 3486 1477 3487 1481
rect 3491 1477 3492 1481
rect 3486 1476 3492 1477
rect 3576 1469 3578 1493
rect 3574 1468 3580 1469
rect 3574 1464 3575 1468
rect 3579 1464 3580 1468
rect 2778 1463 2784 1464
rect 2778 1459 2779 1463
rect 2783 1459 2784 1463
rect 2778 1458 2784 1459
rect 3218 1463 3224 1464
rect 3574 1463 3580 1464
rect 3218 1459 3219 1463
rect 3223 1459 3224 1463
rect 3218 1458 3224 1459
rect 3574 1451 3580 1452
rect 3574 1447 3575 1451
rect 3579 1447 3580 1451
rect 3574 1446 3580 1447
rect 2526 1441 2532 1442
rect 2526 1437 2527 1441
rect 2531 1437 2532 1441
rect 2526 1436 2532 1437
rect 2694 1441 2700 1442
rect 2694 1437 2695 1441
rect 2699 1437 2700 1441
rect 2694 1436 2700 1437
rect 2878 1441 2884 1442
rect 2878 1437 2879 1441
rect 2883 1437 2884 1441
rect 2878 1436 2884 1437
rect 3078 1441 3084 1442
rect 3078 1437 3079 1441
rect 3083 1437 3084 1441
rect 3078 1436 3084 1437
rect 3286 1441 3292 1442
rect 3286 1437 3287 1441
rect 3291 1437 3292 1441
rect 3286 1436 3292 1437
rect 3478 1441 3484 1442
rect 3478 1437 3479 1441
rect 3483 1437 3484 1441
rect 3478 1436 3484 1437
rect 2528 1427 2530 1436
rect 2696 1427 2698 1436
rect 2880 1427 2882 1436
rect 3080 1427 3082 1436
rect 3288 1427 3290 1436
rect 3480 1427 3482 1436
rect 3576 1427 3578 1446
rect 2439 1426 2443 1427
rect 2439 1421 2443 1422
rect 2527 1426 2531 1427
rect 2527 1421 2531 1422
rect 2607 1426 2611 1427
rect 2607 1421 2611 1422
rect 2695 1426 2699 1427
rect 2695 1421 2699 1422
rect 2807 1426 2811 1427
rect 2807 1421 2811 1422
rect 2879 1426 2883 1427
rect 2879 1421 2883 1422
rect 3031 1426 3035 1427
rect 3031 1421 3035 1422
rect 3079 1426 3083 1427
rect 3079 1421 3083 1422
rect 3263 1426 3267 1427
rect 3263 1421 3267 1422
rect 3287 1426 3291 1427
rect 3287 1421 3291 1422
rect 3479 1426 3483 1427
rect 3479 1421 3483 1422
rect 3575 1426 3579 1427
rect 3575 1421 3579 1422
rect 2440 1416 2442 1421
rect 2608 1416 2610 1421
rect 2808 1416 2810 1421
rect 3032 1416 3034 1421
rect 3264 1416 3266 1421
rect 3480 1416 3482 1421
rect 2438 1415 2444 1416
rect 2438 1411 2439 1415
rect 2443 1411 2444 1415
rect 2438 1410 2444 1411
rect 2606 1415 2612 1416
rect 2606 1411 2607 1415
rect 2611 1411 2612 1415
rect 2606 1410 2612 1411
rect 2806 1415 2812 1416
rect 2806 1411 2807 1415
rect 2811 1411 2812 1415
rect 2806 1410 2812 1411
rect 3030 1415 3036 1416
rect 3030 1411 3031 1415
rect 3035 1411 3036 1415
rect 3030 1410 3036 1411
rect 3262 1415 3268 1416
rect 3262 1411 3263 1415
rect 3267 1411 3268 1415
rect 3262 1410 3268 1411
rect 3478 1415 3484 1416
rect 3478 1411 3479 1415
rect 3483 1411 3484 1415
rect 3478 1410 3484 1411
rect 2390 1407 2396 1408
rect 1862 1405 1868 1406
rect 1862 1401 1863 1405
rect 1867 1401 1868 1405
rect 2390 1403 2391 1407
rect 2395 1403 2396 1407
rect 2390 1402 2396 1403
rect 3210 1407 3216 1408
rect 3210 1403 3211 1407
rect 3215 1403 3216 1407
rect 3576 1406 3578 1421
rect 3210 1402 3216 1403
rect 3574 1405 3580 1406
rect 1862 1400 1868 1401
rect 1822 1392 1828 1393
rect 1822 1388 1823 1392
rect 1827 1388 1828 1392
rect 1954 1391 1960 1392
rect 1110 1387 1116 1388
rect 1822 1387 1828 1388
rect 1862 1388 1868 1389
rect 1110 1383 1111 1387
rect 1115 1383 1116 1387
rect 1862 1384 1863 1388
rect 1867 1384 1868 1388
rect 1954 1387 1955 1391
rect 1959 1387 1960 1391
rect 1954 1386 1960 1387
rect 2042 1391 2048 1392
rect 2042 1387 2043 1391
rect 2047 1387 2048 1391
rect 2042 1386 2048 1387
rect 2250 1391 2256 1392
rect 2250 1387 2251 1391
rect 2255 1387 2256 1391
rect 2250 1386 2256 1387
rect 2370 1391 2376 1392
rect 2370 1387 2371 1391
rect 2375 1387 2376 1391
rect 2370 1386 2376 1387
rect 2506 1391 2512 1392
rect 2506 1387 2507 1391
rect 2511 1387 2512 1391
rect 2506 1386 2512 1387
rect 1862 1383 1868 1384
rect 1110 1382 1116 1383
rect 1822 1375 1828 1376
rect 1822 1371 1823 1375
rect 1827 1371 1828 1375
rect 1822 1370 1828 1371
rect 806 1365 812 1366
rect 806 1361 807 1365
rect 811 1361 812 1365
rect 806 1360 812 1361
rect 910 1365 916 1366
rect 910 1361 911 1365
rect 915 1361 916 1365
rect 910 1360 916 1361
rect 1006 1365 1012 1366
rect 1006 1361 1007 1365
rect 1011 1361 1012 1365
rect 1006 1360 1012 1361
rect 1110 1365 1116 1366
rect 1110 1361 1111 1365
rect 1115 1361 1116 1365
rect 1110 1360 1116 1361
rect 1214 1365 1220 1366
rect 1214 1361 1215 1365
rect 1219 1361 1220 1365
rect 1214 1360 1220 1361
rect 1318 1365 1324 1366
rect 1318 1361 1319 1365
rect 1323 1361 1324 1365
rect 1318 1360 1324 1361
rect 808 1351 810 1360
rect 912 1351 914 1360
rect 1008 1351 1010 1360
rect 1112 1351 1114 1360
rect 1216 1351 1218 1360
rect 1320 1351 1322 1360
rect 1366 1359 1372 1360
rect 1366 1355 1367 1359
rect 1371 1355 1372 1359
rect 1366 1354 1372 1355
rect 807 1350 811 1351
rect 807 1345 811 1346
rect 871 1350 875 1351
rect 871 1345 875 1346
rect 911 1350 915 1351
rect 911 1345 915 1346
rect 1007 1350 1011 1351
rect 1007 1345 1011 1346
rect 1039 1350 1043 1351
rect 1039 1345 1043 1346
rect 1111 1350 1115 1351
rect 1111 1345 1115 1346
rect 1207 1350 1211 1351
rect 1207 1345 1211 1346
rect 1215 1350 1219 1351
rect 1215 1345 1219 1346
rect 1319 1350 1323 1351
rect 1319 1345 1323 1346
rect 872 1340 874 1345
rect 1040 1340 1042 1345
rect 1208 1340 1210 1345
rect 870 1339 876 1340
rect 870 1335 871 1339
rect 875 1335 876 1339
rect 870 1334 876 1335
rect 1038 1339 1044 1340
rect 1038 1335 1039 1339
rect 1043 1335 1044 1339
rect 1038 1334 1044 1335
rect 1206 1339 1212 1340
rect 1206 1335 1207 1339
rect 1211 1335 1212 1339
rect 1206 1334 1212 1335
rect 298 1331 304 1332
rect 110 1329 116 1330
rect 110 1325 111 1329
rect 115 1325 116 1329
rect 298 1327 299 1331
rect 303 1327 304 1331
rect 298 1326 304 1327
rect 770 1331 776 1332
rect 770 1327 771 1331
rect 775 1327 776 1331
rect 770 1326 776 1327
rect 110 1324 116 1325
rect 450 1315 456 1316
rect 110 1312 116 1313
rect 110 1308 111 1312
rect 115 1308 116 1312
rect 450 1311 451 1315
rect 455 1311 456 1315
rect 450 1310 456 1311
rect 798 1315 804 1316
rect 798 1311 799 1315
rect 803 1311 804 1315
rect 798 1310 804 1311
rect 1106 1315 1112 1316
rect 1106 1311 1107 1315
rect 1111 1311 1112 1315
rect 1106 1310 1112 1311
rect 1274 1315 1280 1316
rect 1274 1311 1275 1315
rect 1279 1311 1280 1315
rect 1274 1310 1280 1311
rect 110 1307 116 1308
rect 112 1283 114 1307
rect 238 1299 244 1300
rect 238 1295 239 1299
rect 243 1295 244 1299
rect 238 1294 244 1295
rect 390 1299 396 1300
rect 390 1295 391 1299
rect 395 1295 396 1299
rect 390 1294 396 1295
rect 240 1283 242 1294
rect 392 1283 394 1294
rect 452 1288 454 1310
rect 550 1299 556 1300
rect 550 1295 551 1299
rect 555 1295 556 1299
rect 550 1294 556 1295
rect 710 1299 716 1300
rect 710 1295 711 1299
rect 715 1295 716 1299
rect 710 1294 716 1295
rect 450 1287 456 1288
rect 450 1283 451 1287
rect 455 1283 456 1287
rect 552 1283 554 1294
rect 559 1292 563 1293
rect 558 1287 564 1288
rect 558 1283 559 1287
rect 563 1283 564 1287
rect 712 1283 714 1294
rect 800 1293 802 1310
rect 878 1299 884 1300
rect 878 1295 879 1299
rect 883 1295 884 1299
rect 878 1294 884 1295
rect 1046 1299 1052 1300
rect 1046 1295 1047 1299
rect 1051 1295 1052 1299
rect 1046 1294 1052 1295
rect 799 1292 803 1293
rect 799 1287 803 1288
rect 880 1283 882 1294
rect 898 1287 904 1288
rect 898 1283 899 1287
rect 903 1283 904 1287
rect 1048 1283 1050 1294
rect 1108 1288 1110 1310
rect 1214 1299 1220 1300
rect 1214 1295 1215 1299
rect 1219 1295 1220 1299
rect 1214 1294 1220 1295
rect 1106 1287 1112 1288
rect 1106 1283 1107 1287
rect 1111 1283 1112 1287
rect 1216 1283 1218 1294
rect 1276 1288 1278 1310
rect 1368 1288 1370 1354
rect 1824 1351 1826 1370
rect 1864 1355 1866 1383
rect 1894 1375 1900 1376
rect 1894 1371 1895 1375
rect 1899 1371 1900 1375
rect 1894 1370 1900 1371
rect 1896 1355 1898 1370
rect 1956 1364 1958 1386
rect 1982 1375 1988 1376
rect 1982 1371 1983 1375
rect 1987 1371 1988 1375
rect 1982 1370 1988 1371
rect 1954 1363 1960 1364
rect 1954 1359 1955 1363
rect 1959 1359 1960 1363
rect 1954 1358 1960 1359
rect 1984 1355 1986 1370
rect 2044 1364 2046 1386
rect 2078 1375 2084 1376
rect 2078 1371 2079 1375
rect 2083 1371 2084 1375
rect 2078 1370 2084 1371
rect 2190 1375 2196 1376
rect 2190 1371 2191 1375
rect 2195 1371 2196 1375
rect 2190 1370 2196 1371
rect 2042 1363 2048 1364
rect 2042 1359 2043 1363
rect 2047 1359 2048 1363
rect 2042 1358 2048 1359
rect 2080 1355 2082 1370
rect 2192 1355 2194 1370
rect 2252 1364 2254 1386
rect 2310 1375 2316 1376
rect 2310 1371 2311 1375
rect 2315 1371 2316 1375
rect 2310 1370 2316 1371
rect 2250 1363 2256 1364
rect 2250 1359 2251 1363
rect 2255 1359 2256 1363
rect 2250 1358 2256 1359
rect 2312 1355 2314 1370
rect 1863 1354 1867 1355
rect 1375 1350 1379 1351
rect 1375 1345 1379 1346
rect 1823 1350 1827 1351
rect 1863 1349 1867 1350
rect 1895 1354 1899 1355
rect 1895 1349 1899 1350
rect 1983 1354 1987 1355
rect 1983 1349 1987 1350
rect 2079 1354 2083 1355
rect 2079 1349 2083 1350
rect 2103 1354 2107 1355
rect 2103 1349 2107 1350
rect 2191 1354 2195 1355
rect 2191 1349 2195 1350
rect 2223 1354 2227 1355
rect 2223 1349 2227 1350
rect 2311 1354 2315 1355
rect 2311 1349 2315 1350
rect 2359 1354 2363 1355
rect 2359 1349 2363 1350
rect 1823 1345 1827 1346
rect 1376 1340 1378 1345
rect 1374 1339 1380 1340
rect 1374 1335 1375 1339
rect 1379 1335 1380 1339
rect 1374 1334 1380 1335
rect 1824 1330 1826 1345
rect 1822 1329 1828 1330
rect 1822 1325 1823 1329
rect 1827 1325 1828 1329
rect 1864 1325 1866 1349
rect 1896 1338 1898 1349
rect 1984 1338 1986 1349
rect 2104 1338 2106 1349
rect 2224 1338 2226 1349
rect 2360 1338 2362 1349
rect 2372 1348 2374 1386
rect 2446 1375 2452 1376
rect 2446 1371 2447 1375
rect 2451 1371 2452 1375
rect 2446 1370 2452 1371
rect 2448 1355 2450 1370
rect 2508 1364 2510 1386
rect 2614 1375 2620 1376
rect 2614 1371 2615 1375
rect 2619 1371 2620 1375
rect 2614 1370 2620 1371
rect 2814 1375 2820 1376
rect 2814 1371 2815 1375
rect 2819 1371 2820 1375
rect 2814 1370 2820 1371
rect 3038 1375 3044 1376
rect 3038 1371 3039 1375
rect 3043 1371 3044 1375
rect 3038 1370 3044 1371
rect 2506 1363 2512 1364
rect 2506 1359 2507 1363
rect 2511 1359 2512 1363
rect 2506 1358 2512 1359
rect 2616 1355 2618 1370
rect 2775 1364 2779 1365
rect 2774 1359 2775 1364
rect 2779 1359 2780 1364
rect 2774 1358 2780 1359
rect 2816 1355 2818 1370
rect 3040 1355 3042 1370
rect 3212 1365 3214 1402
rect 3574 1401 3575 1405
rect 3579 1401 3580 1405
rect 3574 1400 3580 1401
rect 3254 1391 3260 1392
rect 3254 1387 3255 1391
rect 3259 1387 3260 1391
rect 3254 1386 3260 1387
rect 3470 1391 3476 1392
rect 3470 1387 3471 1391
rect 3475 1387 3476 1391
rect 3470 1386 3476 1387
rect 3574 1388 3580 1389
rect 3211 1364 3215 1365
rect 3256 1364 3258 1386
rect 3270 1375 3276 1376
rect 3270 1371 3271 1375
rect 3275 1371 3276 1375
rect 3270 1370 3276 1371
rect 3211 1359 3215 1360
rect 3254 1363 3260 1364
rect 3254 1359 3255 1363
rect 3259 1359 3260 1363
rect 3254 1358 3260 1359
rect 3272 1355 3274 1370
rect 2447 1354 2451 1355
rect 2447 1349 2451 1350
rect 2511 1354 2515 1355
rect 2511 1349 2515 1350
rect 2615 1354 2619 1355
rect 2615 1349 2619 1350
rect 2687 1354 2691 1355
rect 2687 1349 2691 1350
rect 2815 1354 2819 1355
rect 2815 1349 2819 1350
rect 2871 1354 2875 1355
rect 2871 1349 2875 1350
rect 3039 1354 3043 1355
rect 3039 1349 3043 1350
rect 3071 1354 3075 1355
rect 3071 1349 3075 1350
rect 3271 1354 3275 1355
rect 3271 1349 3275 1350
rect 3279 1354 3283 1355
rect 3279 1349 3283 1350
rect 2370 1347 2376 1348
rect 2370 1343 2371 1347
rect 2375 1343 2376 1347
rect 2370 1342 2376 1343
rect 2512 1338 2514 1349
rect 2688 1338 2690 1349
rect 2872 1338 2874 1349
rect 3072 1338 3074 1349
rect 3254 1347 3260 1348
rect 3254 1343 3255 1347
rect 3259 1343 3260 1347
rect 3254 1342 3260 1343
rect 1894 1337 1900 1338
rect 1894 1333 1895 1337
rect 1899 1333 1900 1337
rect 1894 1332 1900 1333
rect 1982 1337 1988 1338
rect 1982 1333 1983 1337
rect 1987 1333 1988 1337
rect 1982 1332 1988 1333
rect 2102 1337 2108 1338
rect 2102 1333 2103 1337
rect 2107 1333 2108 1337
rect 2102 1332 2108 1333
rect 2222 1337 2228 1338
rect 2222 1333 2223 1337
rect 2227 1333 2228 1337
rect 2222 1332 2228 1333
rect 2358 1337 2364 1338
rect 2358 1333 2359 1337
rect 2363 1333 2364 1337
rect 2358 1332 2364 1333
rect 2510 1337 2516 1338
rect 2510 1333 2511 1337
rect 2515 1333 2516 1337
rect 2510 1332 2516 1333
rect 2686 1337 2692 1338
rect 2686 1333 2687 1337
rect 2691 1333 2692 1337
rect 2686 1332 2692 1333
rect 2870 1337 2876 1338
rect 2870 1333 2871 1337
rect 2875 1333 2876 1337
rect 2870 1332 2876 1333
rect 3070 1337 3076 1338
rect 3070 1333 3071 1337
rect 3075 1333 3076 1337
rect 3070 1332 3076 1333
rect 1822 1324 1828 1325
rect 1862 1324 1868 1325
rect 1862 1320 1863 1324
rect 1867 1320 1868 1324
rect 1862 1319 1868 1320
rect 1822 1312 1828 1313
rect 1822 1308 1823 1312
rect 1827 1308 1828 1312
rect 1822 1307 1828 1308
rect 1862 1307 1868 1308
rect 1382 1299 1388 1300
rect 1382 1295 1383 1299
rect 1387 1295 1388 1299
rect 1382 1294 1388 1295
rect 1274 1287 1280 1288
rect 1274 1283 1275 1287
rect 1279 1283 1280 1287
rect 1366 1287 1372 1288
rect 1366 1283 1367 1287
rect 1371 1283 1372 1287
rect 1384 1283 1386 1294
rect 1824 1283 1826 1307
rect 1862 1303 1863 1307
rect 1867 1303 1868 1307
rect 1862 1302 1868 1303
rect 2958 1307 2964 1308
rect 2958 1303 2959 1307
rect 2963 1303 2964 1307
rect 2958 1302 2964 1303
rect 111 1282 115 1283
rect 111 1277 115 1278
rect 215 1282 219 1283
rect 215 1277 219 1278
rect 239 1282 243 1283
rect 239 1277 243 1278
rect 359 1282 363 1283
rect 359 1277 363 1278
rect 391 1282 395 1283
rect 450 1282 456 1283
rect 519 1282 523 1283
rect 391 1277 395 1278
rect 519 1277 523 1278
rect 551 1282 555 1283
rect 558 1282 564 1283
rect 679 1282 683 1283
rect 551 1277 555 1278
rect 679 1277 683 1278
rect 711 1282 715 1283
rect 711 1277 715 1278
rect 839 1282 843 1283
rect 839 1277 843 1278
rect 879 1282 883 1283
rect 898 1282 904 1283
rect 999 1282 1003 1283
rect 879 1277 883 1278
rect 112 1253 114 1277
rect 198 1275 204 1276
rect 198 1271 199 1275
rect 203 1271 204 1275
rect 198 1270 204 1271
rect 110 1252 116 1253
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 110 1247 116 1248
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 110 1230 116 1231
rect 112 1207 114 1230
rect 111 1206 115 1207
rect 111 1201 115 1202
rect 135 1206 139 1207
rect 135 1201 139 1202
rect 112 1186 114 1201
rect 136 1196 138 1201
rect 134 1195 140 1196
rect 134 1191 135 1195
rect 139 1191 140 1195
rect 134 1190 140 1191
rect 200 1188 202 1270
rect 216 1266 218 1277
rect 360 1266 362 1277
rect 520 1266 522 1277
rect 680 1266 682 1277
rect 840 1266 842 1277
rect 214 1265 220 1266
rect 214 1261 215 1265
rect 219 1261 220 1265
rect 214 1260 220 1261
rect 358 1265 364 1266
rect 358 1261 359 1265
rect 363 1261 364 1265
rect 358 1260 364 1261
rect 518 1265 524 1266
rect 518 1261 519 1265
rect 523 1261 524 1265
rect 518 1260 524 1261
rect 678 1265 684 1266
rect 678 1261 679 1265
rect 683 1261 684 1265
rect 678 1260 684 1261
rect 838 1265 844 1266
rect 838 1261 839 1265
rect 843 1261 844 1265
rect 838 1260 844 1261
rect 900 1252 902 1282
rect 999 1277 1003 1278
rect 1047 1282 1051 1283
rect 1106 1282 1112 1283
rect 1151 1282 1155 1283
rect 1047 1277 1051 1278
rect 1151 1277 1155 1278
rect 1215 1282 1219 1283
rect 1274 1282 1280 1283
rect 1295 1282 1299 1283
rect 1366 1282 1372 1283
rect 1383 1282 1387 1283
rect 1215 1277 1219 1278
rect 1295 1277 1299 1278
rect 1383 1277 1387 1278
rect 1439 1282 1443 1283
rect 1439 1277 1443 1278
rect 1591 1282 1595 1283
rect 1591 1277 1595 1278
rect 1823 1282 1827 1283
rect 1823 1277 1827 1278
rect 1000 1266 1002 1277
rect 1152 1266 1154 1277
rect 1296 1266 1298 1277
rect 1440 1266 1442 1277
rect 1592 1266 1594 1277
rect 998 1265 1004 1266
rect 998 1261 999 1265
rect 1003 1261 1004 1265
rect 998 1260 1004 1261
rect 1150 1265 1156 1266
rect 1150 1261 1151 1265
rect 1155 1261 1156 1265
rect 1150 1260 1156 1261
rect 1294 1265 1300 1266
rect 1294 1261 1295 1265
rect 1299 1261 1300 1265
rect 1294 1260 1300 1261
rect 1438 1265 1444 1266
rect 1438 1261 1439 1265
rect 1443 1261 1444 1265
rect 1438 1260 1444 1261
rect 1590 1265 1596 1266
rect 1590 1261 1591 1265
rect 1595 1261 1596 1265
rect 1590 1260 1596 1261
rect 1824 1253 1826 1277
rect 1864 1275 1866 1302
rect 1886 1297 1892 1298
rect 1886 1293 1887 1297
rect 1891 1293 1892 1297
rect 1886 1292 1892 1293
rect 1974 1297 1980 1298
rect 1974 1293 1975 1297
rect 1979 1293 1980 1297
rect 1974 1292 1980 1293
rect 2094 1297 2100 1298
rect 2094 1293 2095 1297
rect 2099 1293 2100 1297
rect 2094 1292 2100 1293
rect 2214 1297 2220 1298
rect 2214 1293 2215 1297
rect 2219 1293 2220 1297
rect 2214 1292 2220 1293
rect 2350 1297 2356 1298
rect 2350 1293 2351 1297
rect 2355 1293 2356 1297
rect 2350 1292 2356 1293
rect 2502 1297 2508 1298
rect 2502 1293 2503 1297
rect 2507 1293 2508 1297
rect 2502 1292 2508 1293
rect 2678 1297 2684 1298
rect 2678 1293 2679 1297
rect 2683 1293 2684 1297
rect 2678 1292 2684 1293
rect 2862 1297 2868 1298
rect 2862 1293 2863 1297
rect 2867 1293 2868 1297
rect 2862 1292 2868 1293
rect 1888 1275 1890 1292
rect 1976 1275 1978 1292
rect 2096 1275 2098 1292
rect 2216 1275 2218 1292
rect 2352 1275 2354 1292
rect 2504 1275 2506 1292
rect 2680 1275 2682 1292
rect 2864 1275 2866 1292
rect 1863 1274 1867 1275
rect 1863 1269 1867 1270
rect 1887 1274 1891 1275
rect 1887 1269 1891 1270
rect 1975 1274 1979 1275
rect 1975 1269 1979 1270
rect 2055 1274 2059 1275
rect 2055 1269 2059 1270
rect 2095 1274 2099 1275
rect 2095 1269 2099 1270
rect 2143 1274 2147 1275
rect 2143 1269 2147 1270
rect 2215 1274 2219 1275
rect 2215 1269 2219 1270
rect 2239 1274 2243 1275
rect 2239 1269 2243 1270
rect 2335 1274 2339 1275
rect 2335 1269 2339 1270
rect 2351 1274 2355 1275
rect 2351 1269 2355 1270
rect 2431 1274 2435 1275
rect 2431 1269 2435 1270
rect 2503 1274 2507 1275
rect 2503 1269 2507 1270
rect 2551 1274 2555 1275
rect 2551 1269 2555 1270
rect 2679 1274 2683 1275
rect 2679 1269 2683 1270
rect 2687 1274 2691 1275
rect 2687 1269 2691 1270
rect 2855 1274 2859 1275
rect 2855 1269 2859 1270
rect 2863 1274 2867 1275
rect 2863 1269 2867 1270
rect 1864 1254 1866 1269
rect 2056 1264 2058 1269
rect 2144 1264 2146 1269
rect 2240 1264 2242 1269
rect 2336 1264 2338 1269
rect 2432 1264 2434 1269
rect 2552 1264 2554 1269
rect 2688 1264 2690 1269
rect 2856 1264 2858 1269
rect 2054 1263 2060 1264
rect 2054 1259 2055 1263
rect 2059 1259 2060 1263
rect 2054 1258 2060 1259
rect 2142 1263 2148 1264
rect 2142 1259 2143 1263
rect 2147 1259 2148 1263
rect 2142 1258 2148 1259
rect 2238 1263 2244 1264
rect 2238 1259 2239 1263
rect 2243 1259 2244 1263
rect 2238 1258 2244 1259
rect 2334 1263 2340 1264
rect 2334 1259 2335 1263
rect 2339 1259 2340 1263
rect 2334 1258 2340 1259
rect 2430 1263 2436 1264
rect 2430 1259 2431 1263
rect 2435 1259 2436 1263
rect 2430 1258 2436 1259
rect 2550 1263 2556 1264
rect 2550 1259 2551 1263
rect 2555 1259 2556 1263
rect 2686 1263 2692 1264
rect 2550 1258 2556 1259
rect 2567 1260 2571 1261
rect 2686 1259 2687 1263
rect 2691 1259 2692 1263
rect 2686 1258 2692 1259
rect 2854 1263 2860 1264
rect 2854 1259 2855 1263
rect 2859 1259 2860 1263
rect 2960 1261 2962 1302
rect 3062 1297 3068 1298
rect 3062 1293 3063 1297
rect 3067 1293 3068 1297
rect 3062 1292 3068 1293
rect 3064 1275 3066 1292
rect 3039 1274 3043 1275
rect 3039 1269 3043 1270
rect 3063 1274 3067 1275
rect 3063 1269 3067 1270
rect 3231 1274 3235 1275
rect 3231 1269 3235 1270
rect 3040 1264 3042 1269
rect 3232 1264 3234 1269
rect 3038 1263 3044 1264
rect 2854 1258 2860 1259
rect 2959 1260 2963 1261
rect 2122 1255 2128 1256
rect 2567 1255 2571 1256
rect 3038 1259 3039 1263
rect 3043 1259 3044 1263
rect 3038 1258 3044 1259
rect 3230 1263 3236 1264
rect 3230 1259 3231 1263
rect 3235 1259 3236 1263
rect 3230 1258 3236 1259
rect 2959 1255 2963 1256
rect 3106 1255 3112 1256
rect 1862 1253 1868 1254
rect 1822 1252 1828 1253
rect 898 1251 904 1252
rect 898 1247 899 1251
rect 903 1247 904 1251
rect 1822 1248 1823 1252
rect 1827 1248 1828 1252
rect 1862 1249 1863 1253
rect 1867 1249 1868 1253
rect 2122 1251 2123 1255
rect 2127 1251 2128 1255
rect 2122 1250 2128 1251
rect 1862 1248 1868 1249
rect 1822 1247 1828 1248
rect 898 1246 904 1247
rect 1862 1236 1868 1237
rect 1590 1235 1596 1236
rect 1590 1231 1591 1235
rect 1595 1231 1596 1235
rect 1590 1230 1596 1231
rect 1822 1235 1828 1236
rect 1822 1231 1823 1235
rect 1827 1231 1828 1235
rect 1862 1232 1863 1236
rect 1867 1232 1868 1236
rect 1862 1231 1868 1232
rect 1822 1230 1828 1231
rect 206 1225 212 1226
rect 206 1221 207 1225
rect 211 1221 212 1225
rect 206 1220 212 1221
rect 350 1225 356 1226
rect 350 1221 351 1225
rect 355 1221 356 1225
rect 350 1220 356 1221
rect 510 1225 516 1226
rect 510 1221 511 1225
rect 515 1221 516 1225
rect 510 1220 516 1221
rect 670 1225 676 1226
rect 670 1221 671 1225
rect 675 1221 676 1225
rect 670 1220 676 1221
rect 830 1225 836 1226
rect 830 1221 831 1225
rect 835 1221 836 1225
rect 830 1220 836 1221
rect 990 1225 996 1226
rect 990 1221 991 1225
rect 995 1221 996 1225
rect 990 1220 996 1221
rect 1142 1225 1148 1226
rect 1142 1221 1143 1225
rect 1147 1221 1148 1225
rect 1142 1220 1148 1221
rect 1286 1225 1292 1226
rect 1286 1221 1287 1225
rect 1291 1221 1292 1225
rect 1286 1220 1292 1221
rect 1430 1225 1436 1226
rect 1430 1221 1431 1225
rect 1435 1221 1436 1225
rect 1430 1220 1436 1221
rect 1582 1225 1588 1226
rect 1582 1221 1583 1225
rect 1587 1221 1588 1225
rect 1582 1220 1588 1221
rect 208 1207 210 1220
rect 352 1207 354 1220
rect 512 1207 514 1220
rect 672 1207 674 1220
rect 832 1207 834 1220
rect 992 1207 994 1220
rect 1144 1207 1146 1220
rect 1288 1207 1290 1220
rect 1432 1207 1434 1220
rect 1584 1207 1586 1220
rect 207 1206 211 1207
rect 207 1201 211 1202
rect 271 1206 275 1207
rect 271 1201 275 1202
rect 351 1206 355 1207
rect 351 1201 355 1202
rect 423 1206 427 1207
rect 423 1201 427 1202
rect 511 1206 515 1207
rect 511 1201 515 1202
rect 575 1206 579 1207
rect 575 1201 579 1202
rect 671 1206 675 1207
rect 671 1201 675 1202
rect 727 1206 731 1207
rect 727 1201 731 1202
rect 831 1206 835 1207
rect 831 1201 835 1202
rect 887 1206 891 1207
rect 887 1201 891 1202
rect 991 1206 995 1207
rect 991 1201 995 1202
rect 1055 1206 1059 1207
rect 1055 1201 1059 1202
rect 1143 1206 1147 1207
rect 1143 1201 1147 1202
rect 1231 1206 1235 1207
rect 1231 1201 1235 1202
rect 1287 1206 1291 1207
rect 1287 1201 1291 1202
rect 1415 1206 1419 1207
rect 1415 1201 1419 1202
rect 1431 1206 1435 1207
rect 1431 1201 1435 1202
rect 1583 1206 1587 1207
rect 1583 1201 1587 1202
rect 272 1196 274 1201
rect 424 1196 426 1201
rect 576 1196 578 1201
rect 728 1196 730 1201
rect 888 1196 890 1201
rect 1056 1196 1058 1201
rect 1232 1196 1234 1201
rect 1416 1196 1418 1201
rect 270 1195 276 1196
rect 270 1191 271 1195
rect 275 1191 276 1195
rect 270 1190 276 1191
rect 422 1195 428 1196
rect 422 1191 423 1195
rect 427 1191 428 1195
rect 422 1190 428 1191
rect 574 1195 580 1196
rect 574 1191 575 1195
rect 579 1191 580 1195
rect 574 1190 580 1191
rect 726 1195 732 1196
rect 726 1191 727 1195
rect 731 1191 732 1195
rect 726 1190 732 1191
rect 886 1195 892 1196
rect 886 1191 887 1195
rect 891 1191 892 1195
rect 886 1190 892 1191
rect 1054 1195 1060 1196
rect 1054 1191 1055 1195
rect 1059 1191 1060 1195
rect 1054 1190 1060 1191
rect 1230 1195 1236 1196
rect 1230 1191 1231 1195
rect 1235 1191 1236 1195
rect 1230 1190 1236 1191
rect 1414 1195 1420 1196
rect 1414 1191 1415 1195
rect 1419 1191 1420 1195
rect 1414 1190 1420 1191
rect 200 1187 208 1188
rect 110 1185 116 1186
rect 200 1185 203 1187
rect 110 1181 111 1185
rect 115 1181 116 1185
rect 202 1183 203 1185
rect 207 1183 208 1187
rect 202 1182 208 1183
rect 110 1180 116 1181
rect 202 1171 208 1172
rect 110 1168 116 1169
rect 110 1164 111 1168
rect 115 1164 116 1168
rect 202 1167 203 1171
rect 207 1167 208 1171
rect 202 1166 208 1167
rect 338 1171 344 1172
rect 338 1167 339 1171
rect 343 1167 344 1171
rect 338 1166 344 1167
rect 654 1171 660 1172
rect 654 1167 655 1171
rect 659 1167 660 1171
rect 654 1166 660 1167
rect 794 1171 800 1172
rect 794 1167 795 1171
rect 799 1167 800 1171
rect 794 1166 800 1167
rect 954 1171 960 1172
rect 954 1167 955 1171
rect 959 1167 960 1171
rect 954 1166 960 1167
rect 1122 1171 1128 1172
rect 1122 1167 1123 1171
rect 1127 1167 1128 1171
rect 1122 1166 1128 1167
rect 1538 1171 1544 1172
rect 1538 1167 1539 1171
rect 1543 1167 1544 1171
rect 1538 1166 1544 1167
rect 110 1163 116 1164
rect 112 1139 114 1163
rect 142 1155 148 1156
rect 142 1151 143 1155
rect 147 1151 148 1155
rect 142 1150 148 1151
rect 144 1139 146 1150
rect 204 1144 206 1166
rect 278 1155 284 1156
rect 278 1151 279 1155
rect 283 1151 284 1155
rect 278 1150 284 1151
rect 202 1143 208 1144
rect 202 1139 203 1143
rect 207 1139 208 1143
rect 280 1139 282 1150
rect 340 1144 342 1166
rect 430 1155 436 1156
rect 430 1151 431 1155
rect 435 1151 436 1155
rect 430 1150 436 1151
rect 582 1155 588 1156
rect 582 1151 583 1155
rect 587 1151 588 1155
rect 582 1150 588 1151
rect 338 1143 344 1144
rect 338 1139 339 1143
rect 343 1139 344 1143
rect 432 1139 434 1150
rect 584 1139 586 1150
rect 111 1138 115 1139
rect 111 1133 115 1134
rect 143 1138 147 1139
rect 202 1138 208 1139
rect 279 1138 283 1139
rect 143 1133 147 1134
rect 279 1133 283 1134
rect 295 1138 299 1139
rect 338 1138 344 1139
rect 431 1138 435 1139
rect 295 1133 299 1134
rect 431 1133 435 1134
rect 479 1138 483 1139
rect 479 1133 483 1134
rect 583 1138 587 1139
rect 583 1133 587 1134
rect 112 1109 114 1133
rect 144 1122 146 1133
rect 296 1122 298 1133
rect 480 1122 482 1133
rect 656 1132 658 1166
rect 734 1155 740 1156
rect 734 1151 735 1155
rect 739 1151 740 1155
rect 734 1150 740 1151
rect 736 1139 738 1150
rect 796 1144 798 1166
rect 894 1155 900 1156
rect 894 1151 895 1155
rect 899 1151 900 1155
rect 894 1150 900 1151
rect 794 1143 800 1144
rect 794 1139 795 1143
rect 799 1139 800 1143
rect 896 1139 898 1150
rect 956 1144 958 1166
rect 1062 1155 1068 1156
rect 1062 1151 1063 1155
rect 1067 1151 1068 1155
rect 1062 1150 1068 1151
rect 954 1143 960 1144
rect 954 1139 955 1143
rect 959 1139 960 1143
rect 1064 1139 1066 1150
rect 1124 1144 1126 1166
rect 1238 1155 1244 1156
rect 1238 1151 1239 1155
rect 1243 1151 1244 1155
rect 1238 1150 1244 1151
rect 1422 1155 1428 1156
rect 1422 1151 1423 1155
rect 1427 1151 1428 1155
rect 1422 1150 1428 1151
rect 1122 1143 1128 1144
rect 1122 1139 1123 1143
rect 1127 1139 1128 1143
rect 1240 1139 1242 1150
rect 1266 1143 1272 1144
rect 1266 1139 1267 1143
rect 1271 1139 1272 1143
rect 1424 1139 1426 1150
rect 1540 1144 1542 1166
rect 1592 1144 1594 1230
rect 1824 1207 1826 1230
rect 1599 1206 1603 1207
rect 1599 1201 1603 1202
rect 1823 1206 1827 1207
rect 1864 1203 1866 1231
rect 2062 1223 2068 1224
rect 2062 1219 2063 1223
rect 2067 1219 2068 1223
rect 2062 1218 2068 1219
rect 2064 1203 2066 1218
rect 2124 1212 2126 1250
rect 2210 1239 2216 1240
rect 2210 1235 2211 1239
rect 2215 1235 2216 1239
rect 2210 1234 2216 1235
rect 2402 1239 2408 1240
rect 2402 1235 2403 1239
rect 2407 1235 2408 1239
rect 2402 1234 2408 1235
rect 2150 1223 2156 1224
rect 2150 1219 2151 1223
rect 2155 1219 2156 1223
rect 2150 1218 2156 1219
rect 2122 1211 2128 1212
rect 2122 1207 2123 1211
rect 2127 1207 2128 1211
rect 2122 1206 2128 1207
rect 2152 1203 2154 1218
rect 2212 1212 2214 1234
rect 2246 1223 2252 1224
rect 2246 1219 2247 1223
rect 2251 1219 2252 1223
rect 2246 1218 2252 1219
rect 2342 1223 2348 1224
rect 2342 1219 2343 1223
rect 2347 1219 2348 1223
rect 2342 1218 2348 1219
rect 2210 1211 2216 1212
rect 2210 1207 2211 1211
rect 2215 1207 2216 1211
rect 2210 1206 2216 1207
rect 2248 1203 2250 1218
rect 2344 1203 2346 1218
rect 2404 1212 2406 1234
rect 2438 1223 2444 1224
rect 2438 1219 2439 1223
rect 2443 1219 2444 1223
rect 2438 1218 2444 1219
rect 2558 1223 2564 1224
rect 2558 1219 2559 1223
rect 2563 1219 2564 1223
rect 2558 1218 2564 1219
rect 2402 1211 2408 1212
rect 2402 1207 2403 1211
rect 2407 1207 2408 1211
rect 2402 1206 2408 1207
rect 2440 1203 2442 1218
rect 2474 1211 2480 1212
rect 2474 1207 2475 1211
rect 2479 1207 2480 1211
rect 2474 1206 2480 1207
rect 1823 1201 1827 1202
rect 1863 1202 1867 1203
rect 1600 1196 1602 1201
rect 1598 1195 1604 1196
rect 1598 1191 1599 1195
rect 1603 1191 1604 1195
rect 1598 1190 1604 1191
rect 1824 1186 1826 1201
rect 1863 1197 1867 1198
rect 2039 1202 2043 1203
rect 2039 1197 2043 1198
rect 2063 1202 2067 1203
rect 2063 1197 2067 1198
rect 2151 1202 2155 1203
rect 2151 1197 2155 1198
rect 2247 1202 2251 1203
rect 2247 1197 2251 1198
rect 2279 1202 2283 1203
rect 2279 1197 2283 1198
rect 2343 1202 2347 1203
rect 2343 1197 2347 1198
rect 2415 1202 2419 1203
rect 2415 1197 2419 1198
rect 2439 1202 2443 1203
rect 2439 1197 2443 1198
rect 1822 1185 1828 1186
rect 1822 1181 1823 1185
rect 1827 1181 1828 1185
rect 1822 1180 1828 1181
rect 1864 1173 1866 1197
rect 2040 1186 2042 1197
rect 2152 1186 2154 1197
rect 2280 1186 2282 1197
rect 2416 1186 2418 1197
rect 2038 1185 2044 1186
rect 2038 1181 2039 1185
rect 2043 1181 2044 1185
rect 2038 1180 2044 1181
rect 2150 1185 2156 1186
rect 2150 1181 2151 1185
rect 2155 1181 2156 1185
rect 2150 1180 2156 1181
rect 2278 1185 2284 1186
rect 2278 1181 2279 1185
rect 2283 1181 2284 1185
rect 2278 1180 2284 1181
rect 2414 1185 2420 1186
rect 2414 1181 2415 1185
rect 2419 1181 2420 1185
rect 2414 1180 2420 1181
rect 1862 1172 1868 1173
rect 2476 1172 2478 1206
rect 2560 1203 2562 1218
rect 2568 1212 2570 1255
rect 3106 1251 3107 1255
rect 3111 1251 3112 1255
rect 3106 1250 3112 1251
rect 2694 1223 2700 1224
rect 2694 1219 2695 1223
rect 2699 1219 2700 1223
rect 2694 1218 2700 1219
rect 2862 1223 2868 1224
rect 2862 1219 2863 1223
rect 2867 1219 2868 1223
rect 2862 1218 2868 1219
rect 3046 1223 3052 1224
rect 3046 1219 3047 1223
rect 3051 1219 3052 1223
rect 3046 1218 3052 1219
rect 2566 1211 2572 1212
rect 2566 1207 2567 1211
rect 2571 1207 2572 1211
rect 2566 1206 2572 1207
rect 2696 1203 2698 1218
rect 2864 1203 2866 1218
rect 3048 1203 3050 1218
rect 2559 1202 2563 1203
rect 2559 1197 2563 1198
rect 2695 1202 2699 1203
rect 2695 1197 2699 1198
rect 2711 1202 2715 1203
rect 2711 1197 2715 1198
rect 2863 1202 2867 1203
rect 2863 1197 2867 1198
rect 3015 1202 3019 1203
rect 3015 1197 3019 1198
rect 3047 1202 3051 1203
rect 3047 1197 3051 1198
rect 2482 1195 2488 1196
rect 2482 1191 2483 1195
rect 2487 1191 2488 1195
rect 2482 1190 2488 1191
rect 2542 1195 2548 1196
rect 2542 1191 2543 1195
rect 2547 1191 2548 1195
rect 2542 1190 2548 1191
rect 1822 1168 1828 1169
rect 1822 1164 1823 1168
rect 1827 1164 1828 1168
rect 1862 1168 1863 1172
rect 1867 1168 1868 1172
rect 1862 1167 1868 1168
rect 2474 1171 2480 1172
rect 2474 1167 2475 1171
rect 2479 1167 2480 1171
rect 2484 1168 2486 1190
rect 2474 1166 2480 1167
rect 2482 1167 2488 1168
rect 1822 1163 1828 1164
rect 2482 1163 2483 1167
rect 2487 1163 2488 1167
rect 1606 1155 1612 1156
rect 1606 1151 1607 1155
rect 1611 1151 1612 1155
rect 1606 1150 1612 1151
rect 1538 1143 1544 1144
rect 1538 1139 1539 1143
rect 1543 1139 1544 1143
rect 1590 1143 1596 1144
rect 1590 1139 1591 1143
rect 1595 1139 1596 1143
rect 1608 1139 1610 1150
rect 1824 1139 1826 1163
rect 2482 1162 2488 1163
rect 1862 1155 1868 1156
rect 1862 1151 1863 1155
rect 1867 1151 1868 1155
rect 1862 1150 1868 1151
rect 1958 1155 1964 1156
rect 1958 1151 1959 1155
rect 1963 1151 1964 1155
rect 1958 1150 1964 1151
rect 663 1138 667 1139
rect 663 1133 667 1134
rect 735 1138 739 1139
rect 794 1138 800 1139
rect 847 1138 851 1139
rect 735 1133 739 1134
rect 847 1133 851 1134
rect 895 1138 899 1139
rect 954 1138 960 1139
rect 1031 1138 1035 1139
rect 895 1133 899 1134
rect 1031 1133 1035 1134
rect 1063 1138 1067 1139
rect 1122 1138 1128 1139
rect 1207 1138 1211 1139
rect 1063 1133 1067 1134
rect 1207 1133 1211 1134
rect 1239 1138 1243 1139
rect 1266 1138 1272 1139
rect 1391 1138 1395 1139
rect 1239 1133 1243 1134
rect 594 1131 600 1132
rect 594 1127 595 1131
rect 599 1127 600 1131
rect 594 1126 600 1127
rect 654 1131 660 1132
rect 654 1127 655 1131
rect 659 1127 660 1131
rect 654 1126 660 1127
rect 142 1121 148 1122
rect 142 1117 143 1121
rect 147 1117 148 1121
rect 142 1116 148 1117
rect 294 1121 300 1122
rect 294 1117 295 1121
rect 299 1117 300 1121
rect 294 1116 300 1117
rect 478 1121 484 1122
rect 478 1117 479 1121
rect 483 1117 484 1121
rect 478 1116 484 1117
rect 110 1108 116 1109
rect 110 1104 111 1108
rect 115 1104 116 1108
rect 110 1103 116 1104
rect 110 1091 116 1092
rect 110 1087 111 1091
rect 115 1087 116 1091
rect 110 1086 116 1087
rect 362 1091 368 1092
rect 362 1087 363 1091
rect 367 1087 368 1091
rect 362 1086 368 1087
rect 112 1071 114 1086
rect 134 1081 140 1082
rect 134 1077 135 1081
rect 139 1077 140 1081
rect 134 1076 140 1077
rect 286 1081 292 1082
rect 286 1077 287 1081
rect 291 1077 292 1081
rect 286 1076 292 1077
rect 136 1071 138 1076
rect 288 1071 290 1076
rect 111 1070 115 1071
rect 111 1065 115 1066
rect 135 1070 139 1071
rect 135 1065 139 1066
rect 271 1070 275 1071
rect 271 1065 275 1066
rect 287 1070 291 1071
rect 287 1065 291 1066
rect 112 1050 114 1065
rect 136 1060 138 1065
rect 272 1060 274 1065
rect 134 1059 140 1060
rect 134 1055 135 1059
rect 139 1055 140 1059
rect 134 1054 140 1055
rect 270 1059 276 1060
rect 270 1055 271 1059
rect 275 1055 276 1059
rect 270 1054 276 1055
rect 110 1049 116 1050
rect 110 1045 111 1049
rect 115 1045 116 1049
rect 110 1044 116 1045
rect 110 1032 116 1033
rect 110 1028 111 1032
rect 115 1028 116 1032
rect 110 1027 116 1028
rect 112 999 114 1027
rect 142 1019 148 1020
rect 142 1015 143 1019
rect 147 1015 148 1019
rect 142 1014 148 1015
rect 278 1019 284 1020
rect 278 1015 279 1019
rect 283 1015 284 1019
rect 278 1014 284 1015
rect 144 999 146 1014
rect 280 999 282 1014
rect 364 1008 366 1086
rect 470 1081 476 1082
rect 470 1077 471 1081
rect 475 1077 476 1081
rect 470 1076 476 1077
rect 596 1076 598 1126
rect 664 1122 666 1133
rect 848 1122 850 1133
rect 966 1131 972 1132
rect 966 1127 967 1131
rect 971 1127 972 1131
rect 966 1126 972 1127
rect 662 1121 668 1122
rect 662 1117 663 1121
rect 667 1117 668 1121
rect 662 1116 668 1117
rect 846 1121 852 1122
rect 846 1117 847 1121
rect 851 1117 852 1121
rect 846 1116 852 1117
rect 654 1081 660 1082
rect 654 1077 655 1081
rect 659 1077 660 1081
rect 654 1076 660 1077
rect 838 1081 844 1082
rect 838 1077 839 1081
rect 843 1077 844 1081
rect 838 1076 844 1077
rect 472 1071 474 1076
rect 594 1075 600 1076
rect 594 1071 595 1075
rect 599 1071 600 1075
rect 656 1071 658 1076
rect 840 1071 842 1076
rect 431 1070 435 1071
rect 431 1065 435 1066
rect 471 1070 475 1071
rect 471 1065 475 1066
rect 583 1070 587 1071
rect 594 1070 600 1071
rect 655 1070 659 1071
rect 583 1065 587 1066
rect 655 1065 659 1066
rect 735 1070 739 1071
rect 735 1065 739 1066
rect 839 1070 843 1071
rect 839 1065 843 1066
rect 887 1070 891 1071
rect 887 1065 891 1066
rect 432 1060 434 1065
rect 584 1060 586 1065
rect 736 1060 738 1065
rect 888 1060 890 1065
rect 430 1059 436 1060
rect 430 1055 431 1059
rect 435 1055 436 1059
rect 430 1054 436 1055
rect 582 1059 588 1060
rect 582 1055 583 1059
rect 587 1055 588 1059
rect 582 1054 588 1055
rect 734 1059 740 1060
rect 734 1055 735 1059
rect 739 1055 740 1059
rect 734 1054 740 1055
rect 886 1059 892 1060
rect 886 1055 887 1059
rect 891 1055 892 1059
rect 886 1054 892 1055
rect 968 1052 970 1126
rect 1032 1122 1034 1133
rect 1208 1122 1210 1133
rect 1030 1121 1036 1122
rect 1030 1117 1031 1121
rect 1035 1117 1036 1121
rect 1030 1116 1036 1117
rect 1206 1121 1212 1122
rect 1206 1117 1207 1121
rect 1211 1117 1212 1121
rect 1206 1116 1212 1117
rect 1268 1108 1270 1138
rect 1391 1133 1395 1134
rect 1423 1138 1427 1139
rect 1538 1138 1544 1139
rect 1575 1138 1579 1139
rect 1590 1138 1596 1139
rect 1607 1138 1611 1139
rect 1423 1133 1427 1134
rect 1575 1133 1579 1134
rect 1607 1133 1611 1134
rect 1735 1138 1739 1139
rect 1735 1133 1739 1134
rect 1823 1138 1827 1139
rect 1823 1133 1827 1134
rect 1392 1122 1394 1133
rect 1576 1122 1578 1133
rect 1736 1122 1738 1133
rect 1390 1121 1396 1122
rect 1390 1117 1391 1121
rect 1395 1117 1396 1121
rect 1390 1116 1396 1117
rect 1574 1121 1580 1122
rect 1574 1117 1575 1121
rect 1579 1117 1580 1121
rect 1574 1116 1580 1117
rect 1734 1121 1740 1122
rect 1734 1117 1735 1121
rect 1739 1117 1740 1121
rect 1734 1116 1740 1117
rect 1824 1109 1826 1133
rect 1864 1123 1866 1150
rect 1863 1122 1867 1123
rect 1863 1117 1867 1118
rect 1943 1122 1947 1123
rect 1943 1117 1947 1118
rect 1822 1108 1828 1109
rect 1266 1107 1272 1108
rect 1266 1103 1267 1107
rect 1271 1103 1272 1107
rect 1822 1104 1823 1108
rect 1827 1104 1828 1108
rect 1822 1103 1828 1104
rect 1266 1102 1272 1103
rect 1864 1102 1866 1117
rect 1944 1112 1946 1117
rect 1942 1111 1948 1112
rect 1942 1107 1943 1111
rect 1947 1107 1948 1111
rect 1942 1106 1948 1107
rect 1862 1101 1868 1102
rect 1862 1097 1863 1101
rect 1867 1097 1868 1101
rect 1862 1096 1868 1097
rect 1822 1091 1828 1092
rect 1822 1087 1823 1091
rect 1827 1087 1828 1091
rect 1822 1086 1828 1087
rect 1022 1081 1028 1082
rect 1022 1077 1023 1081
rect 1027 1077 1028 1081
rect 1022 1076 1028 1077
rect 1198 1081 1204 1082
rect 1198 1077 1199 1081
rect 1203 1077 1204 1081
rect 1198 1076 1204 1077
rect 1382 1081 1388 1082
rect 1382 1077 1383 1081
rect 1387 1077 1388 1081
rect 1382 1076 1388 1077
rect 1566 1081 1572 1082
rect 1566 1077 1567 1081
rect 1571 1077 1572 1081
rect 1566 1076 1572 1077
rect 1726 1081 1732 1082
rect 1726 1077 1727 1081
rect 1731 1077 1732 1081
rect 1726 1076 1732 1077
rect 1024 1071 1026 1076
rect 1200 1071 1202 1076
rect 1384 1071 1386 1076
rect 1568 1071 1570 1076
rect 1728 1071 1730 1076
rect 1824 1071 1826 1086
rect 1862 1084 1868 1085
rect 1862 1080 1863 1084
rect 1867 1080 1868 1084
rect 1862 1079 1868 1080
rect 1023 1070 1027 1071
rect 1023 1065 1027 1066
rect 1047 1070 1051 1071
rect 1047 1065 1051 1066
rect 1199 1070 1203 1071
rect 1199 1065 1203 1066
rect 1215 1070 1219 1071
rect 1215 1065 1219 1066
rect 1383 1070 1387 1071
rect 1383 1065 1387 1066
rect 1559 1070 1563 1071
rect 1559 1065 1563 1066
rect 1567 1070 1571 1071
rect 1567 1065 1571 1066
rect 1727 1070 1731 1071
rect 1727 1065 1731 1066
rect 1823 1070 1827 1071
rect 1823 1065 1827 1066
rect 1048 1060 1050 1065
rect 1216 1060 1218 1065
rect 1384 1060 1386 1065
rect 1560 1060 1562 1065
rect 1728 1060 1730 1065
rect 1046 1059 1052 1060
rect 1046 1055 1047 1059
rect 1051 1055 1052 1059
rect 1046 1054 1052 1055
rect 1214 1059 1220 1060
rect 1214 1055 1215 1059
rect 1219 1055 1220 1059
rect 1214 1054 1220 1055
rect 1382 1059 1388 1060
rect 1382 1055 1383 1059
rect 1387 1055 1388 1059
rect 1382 1054 1388 1055
rect 1558 1059 1564 1060
rect 1558 1055 1559 1059
rect 1563 1055 1564 1059
rect 1558 1054 1564 1055
rect 1726 1059 1732 1060
rect 1726 1055 1727 1059
rect 1731 1055 1732 1059
rect 1726 1054 1732 1055
rect 966 1051 972 1052
rect 966 1047 967 1051
rect 971 1047 972 1051
rect 966 1046 972 1047
rect 1282 1051 1288 1052
rect 1282 1047 1283 1051
rect 1287 1047 1288 1051
rect 1824 1050 1826 1065
rect 1282 1046 1288 1047
rect 1822 1049 1828 1050
rect 814 1035 820 1036
rect 814 1031 815 1035
rect 819 1031 820 1035
rect 814 1030 820 1031
rect 954 1035 960 1036
rect 954 1031 955 1035
rect 959 1031 960 1035
rect 954 1030 960 1031
rect 438 1019 444 1020
rect 438 1015 439 1019
rect 443 1015 444 1019
rect 438 1014 444 1015
rect 590 1019 596 1020
rect 590 1015 591 1019
rect 595 1015 596 1019
rect 590 1014 596 1015
rect 742 1019 748 1020
rect 742 1015 743 1019
rect 747 1015 748 1019
rect 742 1014 748 1015
rect 362 1007 368 1008
rect 362 1003 363 1007
rect 367 1003 368 1007
rect 362 1002 368 1003
rect 440 999 442 1014
rect 592 999 594 1014
rect 744 999 746 1014
rect 111 998 115 999
rect 111 993 115 994
rect 143 998 147 999
rect 143 993 147 994
rect 279 998 283 999
rect 279 993 283 994
rect 287 998 291 999
rect 287 993 291 994
rect 439 998 443 999
rect 439 993 443 994
rect 463 998 467 999
rect 463 993 467 994
rect 591 998 595 999
rect 591 993 595 994
rect 647 998 651 999
rect 647 993 651 994
rect 743 998 747 999
rect 743 993 747 994
rect 112 969 114 993
rect 144 982 146 993
rect 288 982 290 993
rect 464 982 466 993
rect 648 982 650 993
rect 816 992 818 1030
rect 894 1019 900 1020
rect 894 1015 895 1019
rect 899 1015 900 1019
rect 894 1014 900 1015
rect 896 999 898 1014
rect 956 1008 958 1030
rect 1054 1019 1060 1020
rect 1054 1015 1055 1019
rect 1059 1015 1060 1019
rect 1054 1014 1060 1015
rect 1222 1019 1228 1020
rect 1222 1015 1223 1019
rect 1227 1015 1228 1019
rect 1222 1014 1228 1015
rect 954 1007 960 1008
rect 954 1003 955 1007
rect 959 1003 960 1007
rect 954 1002 960 1003
rect 1056 999 1058 1014
rect 1063 1012 1067 1013
rect 1062 1007 1068 1008
rect 1062 1003 1063 1007
rect 1067 1003 1068 1007
rect 1062 1002 1068 1003
rect 1224 999 1226 1014
rect 1284 1013 1286 1046
rect 1822 1045 1823 1049
rect 1827 1045 1828 1049
rect 1822 1044 1828 1045
rect 1864 1043 1866 1079
rect 1950 1071 1956 1072
rect 1950 1067 1951 1071
rect 1955 1067 1956 1071
rect 1950 1066 1956 1067
rect 1952 1043 1954 1066
rect 1960 1060 1962 1150
rect 2030 1145 2036 1146
rect 2030 1141 2031 1145
rect 2035 1141 2036 1145
rect 2030 1140 2036 1141
rect 2142 1145 2148 1146
rect 2142 1141 2143 1145
rect 2147 1141 2148 1145
rect 2142 1140 2148 1141
rect 2270 1145 2276 1146
rect 2270 1141 2271 1145
rect 2275 1141 2276 1145
rect 2270 1140 2276 1141
rect 2406 1145 2412 1146
rect 2406 1141 2407 1145
rect 2411 1141 2412 1145
rect 2406 1140 2412 1141
rect 2032 1123 2034 1140
rect 2144 1123 2146 1140
rect 2272 1123 2274 1140
rect 2408 1123 2410 1140
rect 2031 1122 2035 1123
rect 2031 1117 2035 1118
rect 2087 1122 2091 1123
rect 2087 1117 2091 1118
rect 2143 1122 2147 1123
rect 2143 1117 2147 1118
rect 2231 1122 2235 1123
rect 2231 1117 2235 1118
rect 2271 1122 2275 1123
rect 2271 1117 2275 1118
rect 2383 1122 2387 1123
rect 2383 1117 2387 1118
rect 2407 1122 2411 1123
rect 2407 1117 2411 1118
rect 2535 1122 2539 1123
rect 2535 1117 2539 1118
rect 2088 1112 2090 1117
rect 2232 1112 2234 1117
rect 2384 1112 2386 1117
rect 2536 1112 2538 1117
rect 2086 1111 2092 1112
rect 2086 1107 2087 1111
rect 2091 1107 2092 1111
rect 2086 1106 2092 1107
rect 2230 1111 2236 1112
rect 2230 1107 2231 1111
rect 2235 1107 2236 1111
rect 2230 1106 2236 1107
rect 2382 1111 2388 1112
rect 2382 1107 2383 1111
rect 2387 1107 2388 1111
rect 2382 1106 2388 1107
rect 2534 1111 2540 1112
rect 2534 1107 2535 1111
rect 2539 1107 2540 1111
rect 2534 1106 2540 1107
rect 2154 1103 2160 1104
rect 2154 1099 2155 1103
rect 2159 1099 2160 1103
rect 2544 1100 2546 1190
rect 2560 1186 2562 1197
rect 2712 1186 2714 1197
rect 2778 1195 2784 1196
rect 2778 1191 2779 1195
rect 2783 1191 2784 1195
rect 2778 1190 2784 1191
rect 2558 1185 2564 1186
rect 2558 1181 2559 1185
rect 2563 1181 2564 1185
rect 2558 1180 2564 1181
rect 2710 1185 2716 1186
rect 2710 1181 2711 1185
rect 2715 1181 2716 1185
rect 2710 1180 2716 1181
rect 2780 1168 2782 1190
rect 2864 1186 2866 1197
rect 2934 1195 2940 1196
rect 2934 1191 2935 1195
rect 2939 1191 2940 1195
rect 2934 1190 2940 1191
rect 2862 1185 2868 1186
rect 2862 1181 2863 1185
rect 2867 1181 2868 1185
rect 2862 1180 2868 1181
rect 2936 1168 2938 1190
rect 3016 1186 3018 1197
rect 3108 1196 3110 1250
rect 3238 1223 3244 1224
rect 3238 1219 3239 1223
rect 3243 1219 3244 1223
rect 3238 1218 3244 1219
rect 3240 1203 3242 1218
rect 3167 1202 3171 1203
rect 3167 1197 3171 1198
rect 3239 1202 3243 1203
rect 3239 1197 3243 1198
rect 3106 1195 3112 1196
rect 3106 1191 3107 1195
rect 3111 1191 3112 1195
rect 3106 1190 3112 1191
rect 3168 1186 3170 1197
rect 3246 1195 3252 1196
rect 3246 1191 3247 1195
rect 3251 1191 3252 1195
rect 3246 1190 3252 1191
rect 3014 1185 3020 1186
rect 3014 1181 3015 1185
rect 3019 1181 3020 1185
rect 3014 1180 3020 1181
rect 3166 1185 3172 1186
rect 3166 1181 3167 1185
rect 3171 1181 3172 1185
rect 3166 1180 3172 1181
rect 3248 1168 3250 1190
rect 3256 1176 3258 1342
rect 3280 1338 3282 1349
rect 3472 1348 3474 1386
rect 3574 1384 3575 1388
rect 3579 1384 3580 1388
rect 3574 1383 3580 1384
rect 3486 1375 3492 1376
rect 3486 1371 3487 1375
rect 3491 1371 3492 1375
rect 3486 1370 3492 1371
rect 3488 1355 3490 1370
rect 3576 1355 3578 1383
rect 3487 1354 3491 1355
rect 3487 1349 3491 1350
rect 3575 1354 3579 1355
rect 3575 1349 3579 1350
rect 3470 1347 3476 1348
rect 3470 1343 3471 1347
rect 3475 1343 3476 1347
rect 3470 1342 3476 1343
rect 3488 1338 3490 1349
rect 3278 1337 3284 1338
rect 3278 1333 3279 1337
rect 3283 1333 3284 1337
rect 3278 1332 3284 1333
rect 3486 1337 3492 1338
rect 3486 1333 3487 1337
rect 3491 1333 3492 1337
rect 3486 1332 3492 1333
rect 3576 1325 3578 1349
rect 3574 1324 3580 1325
rect 3574 1320 3575 1324
rect 3579 1320 3580 1324
rect 3574 1319 3580 1320
rect 3454 1307 3460 1308
rect 3454 1303 3455 1307
rect 3459 1303 3460 1307
rect 3454 1302 3460 1303
rect 3574 1307 3580 1308
rect 3574 1303 3575 1307
rect 3579 1303 3580 1307
rect 3574 1302 3580 1303
rect 3270 1297 3276 1298
rect 3270 1293 3271 1297
rect 3275 1293 3276 1297
rect 3270 1292 3276 1293
rect 3272 1275 3274 1292
rect 3271 1274 3275 1275
rect 3271 1269 3275 1270
rect 3431 1274 3435 1275
rect 3431 1269 3435 1270
rect 3432 1264 3434 1269
rect 3430 1263 3436 1264
rect 3430 1259 3431 1263
rect 3435 1259 3436 1263
rect 3430 1258 3436 1259
rect 3438 1223 3444 1224
rect 3438 1219 3439 1223
rect 3443 1219 3444 1223
rect 3438 1218 3444 1219
rect 3440 1203 3442 1218
rect 3456 1212 3458 1302
rect 3478 1297 3484 1298
rect 3478 1293 3479 1297
rect 3483 1293 3484 1297
rect 3478 1292 3484 1293
rect 3480 1275 3482 1292
rect 3576 1275 3578 1302
rect 3479 1274 3483 1275
rect 3479 1269 3483 1270
rect 3575 1274 3579 1275
rect 3575 1269 3579 1270
rect 3576 1254 3578 1269
rect 3574 1253 3580 1254
rect 3574 1249 3575 1253
rect 3579 1249 3580 1253
rect 3574 1248 3580 1249
rect 3498 1239 3504 1240
rect 3498 1235 3499 1239
rect 3503 1235 3504 1239
rect 3498 1234 3504 1235
rect 3574 1236 3580 1237
rect 3454 1211 3460 1212
rect 3454 1207 3455 1211
rect 3459 1207 3460 1211
rect 3454 1206 3460 1207
rect 3327 1202 3331 1203
rect 3327 1197 3331 1198
rect 3439 1202 3443 1203
rect 3439 1197 3443 1198
rect 3487 1202 3491 1203
rect 3487 1197 3491 1198
rect 3328 1186 3330 1197
rect 3488 1186 3490 1197
rect 3500 1196 3502 1234
rect 3574 1232 3575 1236
rect 3579 1232 3580 1236
rect 3574 1231 3580 1232
rect 3576 1203 3578 1231
rect 3575 1202 3579 1203
rect 3575 1197 3579 1198
rect 3498 1195 3504 1196
rect 3498 1191 3499 1195
rect 3503 1191 3504 1195
rect 3498 1190 3504 1191
rect 3326 1185 3332 1186
rect 3326 1181 3327 1185
rect 3331 1181 3332 1185
rect 3326 1180 3332 1181
rect 3486 1185 3492 1186
rect 3486 1181 3487 1185
rect 3491 1181 3492 1185
rect 3486 1180 3492 1181
rect 3254 1175 3260 1176
rect 3254 1171 3255 1175
rect 3259 1171 3260 1175
rect 3576 1173 3578 1197
rect 3254 1170 3260 1171
rect 3574 1172 3580 1173
rect 3574 1168 3575 1172
rect 3579 1168 3580 1172
rect 2778 1167 2784 1168
rect 2778 1163 2779 1167
rect 2783 1163 2784 1167
rect 2778 1162 2784 1163
rect 2934 1167 2940 1168
rect 2934 1163 2935 1167
rect 2939 1163 2940 1167
rect 2934 1162 2940 1163
rect 3246 1167 3252 1168
rect 3574 1167 3580 1168
rect 3246 1163 3247 1167
rect 3251 1163 3252 1167
rect 3246 1162 3252 1163
rect 2710 1155 2716 1156
rect 2710 1151 2711 1155
rect 2715 1151 2716 1155
rect 2710 1150 2716 1151
rect 3574 1155 3580 1156
rect 3574 1151 3575 1155
rect 3579 1151 3580 1155
rect 3574 1150 3580 1151
rect 2550 1145 2556 1146
rect 2550 1141 2551 1145
rect 2555 1141 2556 1145
rect 2550 1140 2556 1141
rect 2702 1145 2708 1146
rect 2702 1141 2703 1145
rect 2707 1141 2708 1145
rect 2702 1140 2708 1141
rect 2552 1123 2554 1140
rect 2704 1123 2706 1140
rect 2551 1122 2555 1123
rect 2551 1117 2555 1118
rect 2687 1122 2691 1123
rect 2687 1117 2691 1118
rect 2703 1122 2707 1123
rect 2703 1117 2707 1118
rect 2688 1112 2690 1117
rect 2686 1111 2692 1112
rect 2686 1107 2687 1111
rect 2691 1107 2692 1111
rect 2686 1106 2692 1107
rect 2154 1098 2160 1099
rect 2542 1099 2548 1100
rect 2094 1071 2100 1072
rect 2094 1067 2095 1071
rect 2099 1067 2100 1071
rect 2094 1066 2100 1067
rect 1958 1059 1964 1060
rect 1958 1055 1959 1059
rect 1963 1055 1964 1059
rect 1958 1054 1964 1055
rect 2096 1043 2098 1066
rect 1863 1042 1867 1043
rect 1863 1037 1867 1038
rect 1919 1042 1923 1043
rect 1919 1037 1923 1038
rect 1951 1042 1955 1043
rect 1951 1037 1955 1038
rect 2095 1042 2099 1043
rect 2095 1037 2099 1038
rect 2127 1042 2131 1043
rect 2127 1037 2131 1038
rect 1646 1035 1652 1036
rect 1646 1031 1647 1035
rect 1651 1031 1652 1035
rect 1646 1030 1652 1031
rect 1822 1032 1828 1033
rect 1390 1019 1396 1020
rect 1390 1015 1391 1019
rect 1395 1015 1396 1019
rect 1390 1014 1396 1015
rect 1566 1019 1572 1020
rect 1566 1015 1567 1019
rect 1571 1015 1572 1019
rect 1566 1014 1572 1015
rect 1283 1012 1287 1013
rect 1230 1007 1236 1008
rect 1283 1007 1287 1008
rect 1230 1003 1231 1007
rect 1235 1003 1236 1007
rect 1230 1002 1236 1003
rect 823 998 827 999
rect 823 993 827 994
rect 895 998 899 999
rect 895 993 899 994
rect 999 998 1003 999
rect 999 993 1003 994
rect 1055 998 1059 999
rect 1055 993 1059 994
rect 1167 998 1171 999
rect 1167 993 1171 994
rect 1223 998 1227 999
rect 1223 993 1227 994
rect 814 991 820 992
rect 814 987 815 991
rect 819 987 820 991
rect 814 986 820 987
rect 824 982 826 993
rect 1000 982 1002 993
rect 1006 991 1012 992
rect 1006 987 1007 991
rect 1011 987 1012 991
rect 1006 986 1012 987
rect 142 981 148 982
rect 142 977 143 981
rect 147 977 148 981
rect 142 976 148 977
rect 286 981 292 982
rect 286 977 287 981
rect 291 977 292 981
rect 286 976 292 977
rect 462 981 468 982
rect 462 977 463 981
rect 467 977 468 981
rect 462 976 468 977
rect 646 981 652 982
rect 646 977 647 981
rect 651 977 652 981
rect 646 976 652 977
rect 822 981 828 982
rect 822 977 823 981
rect 827 977 828 981
rect 822 976 828 977
rect 998 981 1004 982
rect 998 977 999 981
rect 1003 977 1004 981
rect 998 976 1004 977
rect 110 968 116 969
rect 110 964 111 968
rect 115 964 116 968
rect 110 963 116 964
rect 110 951 116 952
rect 110 947 111 951
rect 115 947 116 951
rect 110 946 116 947
rect 112 923 114 946
rect 134 941 140 942
rect 134 937 135 941
rect 139 937 140 941
rect 134 936 140 937
rect 278 941 284 942
rect 278 937 279 941
rect 283 937 284 941
rect 278 936 284 937
rect 454 941 460 942
rect 454 937 455 941
rect 459 937 460 941
rect 454 936 460 937
rect 638 941 644 942
rect 638 937 639 941
rect 643 937 644 941
rect 638 936 644 937
rect 814 941 820 942
rect 814 937 815 941
rect 819 937 820 941
rect 814 936 820 937
rect 990 941 996 942
rect 990 937 991 941
rect 995 937 996 941
rect 990 936 996 937
rect 136 923 138 936
rect 280 923 282 936
rect 456 923 458 936
rect 640 923 642 936
rect 816 923 818 936
rect 992 923 994 936
rect 111 922 115 923
rect 111 917 115 918
rect 135 922 139 923
rect 135 917 139 918
rect 271 922 275 923
rect 271 917 275 918
rect 279 922 283 923
rect 279 917 283 918
rect 439 922 443 923
rect 439 917 443 918
rect 455 922 459 923
rect 455 917 459 918
rect 607 922 611 923
rect 607 917 611 918
rect 639 922 643 923
rect 639 917 643 918
rect 775 922 779 923
rect 775 917 779 918
rect 815 922 819 923
rect 815 917 819 918
rect 935 922 939 923
rect 935 917 939 918
rect 991 922 995 923
rect 991 917 995 918
rect 112 902 114 917
rect 136 912 138 917
rect 272 912 274 917
rect 440 912 442 917
rect 608 912 610 917
rect 776 912 778 917
rect 936 912 938 917
rect 134 911 140 912
rect 134 907 135 911
rect 139 907 140 911
rect 134 906 140 907
rect 270 911 276 912
rect 270 907 271 911
rect 275 907 276 911
rect 270 906 276 907
rect 438 911 444 912
rect 438 907 439 911
rect 443 907 444 911
rect 438 906 444 907
rect 606 911 612 912
rect 606 907 607 911
rect 611 907 612 911
rect 606 906 612 907
rect 774 911 780 912
rect 774 907 775 911
rect 779 907 780 911
rect 774 906 780 907
rect 934 911 940 912
rect 934 907 935 911
rect 939 907 940 911
rect 934 906 940 907
rect 1008 904 1010 986
rect 1168 982 1170 993
rect 1166 981 1172 982
rect 1166 977 1167 981
rect 1171 977 1172 981
rect 1166 976 1172 977
rect 1232 968 1234 1002
rect 1392 999 1394 1014
rect 1568 999 1570 1014
rect 1578 999 1584 1000
rect 1327 998 1331 999
rect 1327 993 1331 994
rect 1391 998 1395 999
rect 1391 993 1395 994
rect 1487 998 1491 999
rect 1487 993 1491 994
rect 1567 998 1571 999
rect 1578 995 1579 999
rect 1583 995 1584 999
rect 1578 994 1584 995
rect 1567 993 1571 994
rect 1328 982 1330 993
rect 1488 982 1490 993
rect 1326 981 1332 982
rect 1326 977 1327 981
rect 1331 977 1332 981
rect 1326 976 1332 977
rect 1486 981 1492 982
rect 1486 977 1487 981
rect 1491 977 1492 981
rect 1486 976 1492 977
rect 1230 967 1236 968
rect 1230 963 1231 967
rect 1235 963 1236 967
rect 1580 964 1582 994
rect 1648 992 1650 1030
rect 1822 1028 1823 1032
rect 1827 1028 1828 1032
rect 1822 1027 1828 1028
rect 1734 1019 1740 1020
rect 1734 1015 1735 1019
rect 1739 1015 1740 1019
rect 1734 1014 1740 1015
rect 1736 999 1738 1014
rect 1824 999 1826 1027
rect 1864 1013 1866 1037
rect 1920 1026 1922 1037
rect 1986 1035 1992 1036
rect 1986 1031 1987 1035
rect 1991 1031 1992 1035
rect 1986 1030 1992 1031
rect 1918 1025 1924 1026
rect 1918 1021 1919 1025
rect 1923 1021 1924 1025
rect 1918 1020 1924 1021
rect 1862 1012 1868 1013
rect 1862 1008 1863 1012
rect 1867 1008 1868 1012
rect 1988 1008 1990 1030
rect 2128 1026 2130 1037
rect 2156 1036 2158 1098
rect 2542 1095 2543 1099
rect 2547 1095 2548 1099
rect 2542 1094 2548 1095
rect 2238 1071 2244 1072
rect 2238 1067 2239 1071
rect 2243 1067 2244 1071
rect 2238 1066 2244 1067
rect 2390 1071 2396 1072
rect 2390 1067 2391 1071
rect 2395 1067 2396 1071
rect 2390 1066 2396 1067
rect 2542 1071 2548 1072
rect 2542 1067 2543 1071
rect 2547 1067 2548 1071
rect 2542 1066 2548 1067
rect 2694 1071 2700 1072
rect 2694 1067 2695 1071
rect 2699 1067 2700 1071
rect 2694 1066 2700 1067
rect 2240 1043 2242 1066
rect 2392 1043 2394 1066
rect 2544 1043 2546 1066
rect 2696 1043 2698 1066
rect 2712 1060 2714 1150
rect 2854 1145 2860 1146
rect 2854 1141 2855 1145
rect 2859 1141 2860 1145
rect 2854 1140 2860 1141
rect 3006 1145 3012 1146
rect 3006 1141 3007 1145
rect 3011 1141 3012 1145
rect 3006 1140 3012 1141
rect 3158 1145 3164 1146
rect 3158 1141 3159 1145
rect 3163 1141 3164 1145
rect 3158 1140 3164 1141
rect 3318 1145 3324 1146
rect 3318 1141 3319 1145
rect 3323 1141 3324 1145
rect 3318 1140 3324 1141
rect 3478 1145 3484 1146
rect 3478 1141 3479 1145
rect 3483 1141 3484 1145
rect 3478 1140 3484 1141
rect 2856 1123 2858 1140
rect 3008 1123 3010 1140
rect 3160 1123 3162 1140
rect 3320 1123 3322 1140
rect 3480 1123 3482 1140
rect 3576 1123 3578 1150
rect 2839 1122 2843 1123
rect 2839 1117 2843 1118
rect 2855 1122 2859 1123
rect 2855 1117 2859 1118
rect 2991 1122 2995 1123
rect 2991 1117 2995 1118
rect 3007 1122 3011 1123
rect 3007 1117 3011 1118
rect 3151 1122 3155 1123
rect 3151 1117 3155 1118
rect 3159 1122 3163 1123
rect 3159 1117 3163 1118
rect 3319 1122 3323 1123
rect 3319 1117 3323 1118
rect 3479 1122 3483 1123
rect 3479 1117 3483 1118
rect 3575 1122 3579 1123
rect 3575 1117 3579 1118
rect 2840 1112 2842 1117
rect 2992 1112 2994 1117
rect 3152 1112 3154 1117
rect 3320 1112 3322 1117
rect 3480 1112 3482 1117
rect 2838 1111 2844 1112
rect 2838 1107 2839 1111
rect 2843 1107 2844 1111
rect 2838 1106 2844 1107
rect 2990 1111 2996 1112
rect 2990 1107 2991 1111
rect 2995 1107 2996 1111
rect 2990 1106 2996 1107
rect 3150 1111 3156 1112
rect 3150 1107 3151 1111
rect 3155 1107 3156 1111
rect 3150 1106 3156 1107
rect 3318 1111 3324 1112
rect 3318 1107 3319 1111
rect 3323 1107 3324 1111
rect 3318 1106 3324 1107
rect 3478 1111 3484 1112
rect 3478 1107 3479 1111
rect 3483 1107 3484 1111
rect 3478 1106 3484 1107
rect 3078 1103 3084 1104
rect 3078 1099 3079 1103
rect 3083 1099 3084 1103
rect 3576 1102 3578 1117
rect 3078 1098 3084 1099
rect 3574 1101 3580 1102
rect 2846 1071 2852 1072
rect 2846 1067 2847 1071
rect 2851 1067 2852 1071
rect 2846 1066 2852 1067
rect 2998 1071 3004 1072
rect 2998 1067 2999 1071
rect 3003 1067 3004 1071
rect 2998 1066 3004 1067
rect 2710 1059 2716 1060
rect 2710 1055 2711 1059
rect 2715 1055 2716 1059
rect 2710 1054 2716 1055
rect 2703 1052 2707 1053
rect 2703 1047 2707 1048
rect 2239 1042 2243 1043
rect 2239 1037 2243 1038
rect 2327 1042 2331 1043
rect 2327 1037 2331 1038
rect 2391 1042 2395 1043
rect 2391 1037 2395 1038
rect 2519 1042 2523 1043
rect 2519 1037 2523 1038
rect 2543 1042 2547 1043
rect 2543 1037 2547 1038
rect 2695 1042 2699 1043
rect 2695 1037 2699 1038
rect 2154 1035 2160 1036
rect 2154 1031 2155 1035
rect 2159 1031 2160 1035
rect 2154 1030 2160 1031
rect 2328 1026 2330 1037
rect 2520 1026 2522 1037
rect 2526 1035 2532 1036
rect 2526 1031 2527 1035
rect 2531 1031 2532 1035
rect 2526 1030 2532 1031
rect 2126 1025 2132 1026
rect 2126 1021 2127 1025
rect 2131 1021 2132 1025
rect 2126 1020 2132 1021
rect 2326 1025 2332 1026
rect 2326 1021 2327 1025
rect 2331 1021 2332 1025
rect 2326 1020 2332 1021
rect 2518 1025 2524 1026
rect 2518 1021 2519 1025
rect 2523 1021 2524 1025
rect 2518 1020 2524 1021
rect 1862 1007 1868 1008
rect 1986 1007 1992 1008
rect 1986 1003 1987 1007
rect 1991 1003 1992 1007
rect 1986 1002 1992 1003
rect 1655 998 1659 999
rect 1655 993 1659 994
rect 1735 998 1739 999
rect 1735 993 1739 994
rect 1823 998 1827 999
rect 1823 993 1827 994
rect 1862 995 1868 996
rect 1646 991 1652 992
rect 1646 987 1647 991
rect 1651 987 1652 991
rect 1646 986 1652 987
rect 1656 982 1658 993
rect 1654 981 1660 982
rect 1654 977 1655 981
rect 1659 977 1660 981
rect 1654 976 1660 977
rect 1824 969 1826 993
rect 1862 991 1863 995
rect 1867 991 1868 995
rect 1862 990 1868 991
rect 1902 995 1908 996
rect 1902 991 1903 995
rect 1907 991 1908 995
rect 1902 990 1908 991
rect 1864 971 1866 990
rect 1863 970 1867 971
rect 1822 968 1828 969
rect 1822 964 1823 968
rect 1827 964 1828 968
rect 1863 965 1867 966
rect 1887 970 1891 971
rect 1887 965 1891 966
rect 1230 962 1236 963
rect 1578 963 1584 964
rect 1822 963 1828 964
rect 1578 959 1579 963
rect 1583 959 1584 963
rect 1578 958 1584 959
rect 1822 951 1828 952
rect 1822 947 1823 951
rect 1827 947 1828 951
rect 1864 950 1866 965
rect 1888 960 1890 965
rect 1886 959 1892 960
rect 1886 955 1887 959
rect 1891 955 1892 959
rect 1886 954 1892 955
rect 1822 946 1828 947
rect 1862 949 1868 950
rect 1158 941 1164 942
rect 1158 937 1159 941
rect 1163 937 1164 941
rect 1158 936 1164 937
rect 1318 941 1324 942
rect 1318 937 1319 941
rect 1323 937 1324 941
rect 1318 936 1324 937
rect 1478 941 1484 942
rect 1478 937 1479 941
rect 1483 937 1484 941
rect 1478 936 1484 937
rect 1646 941 1652 942
rect 1646 937 1647 941
rect 1651 937 1652 941
rect 1646 936 1652 937
rect 1160 923 1162 936
rect 1320 923 1322 936
rect 1480 923 1482 936
rect 1648 923 1650 936
rect 1824 923 1826 946
rect 1862 945 1863 949
rect 1867 945 1868 949
rect 1862 944 1868 945
rect 1862 932 1868 933
rect 1862 928 1863 932
rect 1867 928 1868 932
rect 1862 927 1868 928
rect 1095 922 1099 923
rect 1095 917 1099 918
rect 1159 922 1163 923
rect 1159 917 1163 918
rect 1247 922 1251 923
rect 1247 917 1251 918
rect 1319 922 1323 923
rect 1319 917 1323 918
rect 1399 922 1403 923
rect 1399 917 1403 918
rect 1479 922 1483 923
rect 1479 917 1483 918
rect 1551 922 1555 923
rect 1551 917 1555 918
rect 1647 922 1651 923
rect 1647 917 1651 918
rect 1823 922 1827 923
rect 1823 917 1827 918
rect 1096 912 1098 917
rect 1248 912 1250 917
rect 1400 912 1402 917
rect 1552 912 1554 917
rect 1094 911 1100 912
rect 1094 907 1095 911
rect 1099 907 1100 911
rect 1094 906 1100 907
rect 1246 911 1252 912
rect 1246 907 1247 911
rect 1251 907 1252 911
rect 1246 906 1252 907
rect 1398 911 1404 912
rect 1398 907 1399 911
rect 1403 907 1404 911
rect 1398 906 1404 907
rect 1550 911 1556 912
rect 1550 907 1551 911
rect 1555 907 1556 911
rect 1550 906 1556 907
rect 706 903 712 904
rect 110 901 116 902
rect 110 897 111 901
rect 115 897 116 901
rect 706 899 707 903
rect 711 899 712 903
rect 706 898 712 899
rect 1006 903 1012 904
rect 1006 899 1007 903
rect 1011 899 1012 903
rect 1824 902 1826 917
rect 1006 898 1012 899
rect 1822 901 1828 902
rect 110 896 116 897
rect 202 887 208 888
rect 110 884 116 885
rect 110 880 111 884
rect 115 880 116 884
rect 202 883 203 887
rect 207 883 208 887
rect 202 882 208 883
rect 338 887 344 888
rect 338 883 339 887
rect 343 883 344 887
rect 338 882 344 883
rect 110 879 116 880
rect 112 855 114 879
rect 142 871 148 872
rect 142 867 143 871
rect 147 867 148 871
rect 142 866 148 867
rect 144 855 146 866
rect 204 860 206 882
rect 278 871 284 872
rect 278 867 279 871
rect 283 867 284 871
rect 278 866 284 867
rect 198 859 206 860
rect 198 855 199 859
rect 203 857 206 859
rect 203 855 204 857
rect 280 855 282 866
rect 111 854 115 855
rect 111 849 115 850
rect 143 854 147 855
rect 198 854 204 855
rect 279 854 283 855
rect 143 849 147 850
rect 279 849 283 850
rect 287 854 291 855
rect 287 849 291 850
rect 112 825 114 849
rect 144 838 146 849
rect 288 838 290 849
rect 340 848 342 882
rect 446 871 452 872
rect 446 867 447 871
rect 451 867 452 871
rect 614 871 620 872
rect 446 866 452 867
rect 455 868 459 869
rect 448 855 450 866
rect 614 867 615 871
rect 619 867 620 871
rect 708 869 710 898
rect 1822 897 1823 901
rect 1827 897 1828 901
rect 1822 896 1828 897
rect 1864 895 1866 927
rect 1894 919 1900 920
rect 1894 915 1895 919
rect 1899 915 1900 919
rect 1894 914 1900 915
rect 1896 895 1898 914
rect 1904 908 1906 990
rect 1910 985 1916 986
rect 1910 981 1911 985
rect 1915 981 1916 985
rect 1910 980 1916 981
rect 2118 985 2124 986
rect 2118 981 2119 985
rect 2123 981 2124 985
rect 2118 980 2124 981
rect 2318 985 2324 986
rect 2318 981 2319 985
rect 2323 981 2324 985
rect 2318 980 2324 981
rect 2510 985 2516 986
rect 2510 981 2511 985
rect 2515 981 2516 985
rect 2510 980 2516 981
rect 1912 971 1914 980
rect 2120 971 2122 980
rect 2320 971 2322 980
rect 2512 971 2514 980
rect 1911 970 1915 971
rect 1911 965 1915 966
rect 2071 970 2075 971
rect 2071 965 2075 966
rect 2119 970 2123 971
rect 2119 965 2123 966
rect 2263 970 2267 971
rect 2263 965 2267 966
rect 2319 970 2323 971
rect 2319 965 2323 966
rect 2455 970 2459 971
rect 2455 965 2459 966
rect 2511 970 2515 971
rect 2511 965 2515 966
rect 2072 960 2074 965
rect 2264 960 2266 965
rect 2456 960 2458 965
rect 2070 959 2076 960
rect 2070 955 2071 959
rect 2075 955 2076 959
rect 2070 954 2076 955
rect 2262 959 2268 960
rect 2262 955 2263 959
rect 2267 955 2268 959
rect 2262 954 2268 955
rect 2454 959 2460 960
rect 2454 955 2455 959
rect 2459 955 2460 959
rect 2454 954 2460 955
rect 2528 952 2530 1030
rect 2696 1026 2698 1037
rect 2704 1036 2706 1047
rect 2848 1043 2850 1066
rect 3000 1043 3002 1066
rect 3080 1053 3082 1098
rect 3574 1097 3575 1101
rect 3579 1097 3580 1101
rect 3574 1096 3580 1097
rect 3470 1087 3476 1088
rect 3470 1083 3471 1087
rect 3475 1083 3476 1087
rect 3470 1082 3476 1083
rect 3574 1084 3580 1085
rect 3158 1071 3164 1072
rect 3158 1067 3159 1071
rect 3163 1067 3164 1071
rect 3158 1066 3164 1067
rect 3326 1071 3332 1072
rect 3326 1067 3327 1071
rect 3331 1067 3332 1071
rect 3326 1066 3332 1067
rect 3079 1052 3083 1053
rect 3079 1047 3083 1048
rect 3160 1043 3162 1066
rect 3328 1043 3330 1066
rect 2847 1042 2851 1043
rect 2847 1037 2851 1038
rect 2863 1042 2867 1043
rect 2863 1037 2867 1038
rect 2999 1042 3003 1043
rect 2999 1037 3003 1038
rect 3023 1042 3027 1043
rect 3023 1037 3027 1038
rect 3159 1042 3163 1043
rect 3159 1037 3163 1038
rect 3183 1042 3187 1043
rect 3183 1037 3187 1038
rect 3327 1042 3331 1043
rect 3327 1037 3331 1038
rect 3343 1042 3347 1043
rect 3343 1037 3347 1038
rect 2702 1035 2708 1036
rect 2702 1031 2703 1035
rect 2707 1031 2708 1035
rect 2702 1030 2708 1031
rect 2864 1026 2866 1037
rect 3024 1026 3026 1037
rect 3184 1026 3186 1037
rect 3344 1026 3346 1037
rect 3472 1036 3474 1082
rect 3574 1080 3575 1084
rect 3579 1080 3580 1084
rect 3574 1079 3580 1080
rect 3486 1071 3492 1072
rect 3486 1067 3487 1071
rect 3491 1067 3492 1071
rect 3486 1066 3492 1067
rect 3488 1043 3490 1066
rect 3576 1043 3578 1079
rect 3487 1042 3491 1043
rect 3487 1037 3491 1038
rect 3575 1042 3579 1043
rect 3575 1037 3579 1038
rect 3350 1035 3356 1036
rect 3350 1031 3351 1035
rect 3355 1031 3356 1035
rect 3350 1030 3356 1031
rect 3470 1035 3476 1036
rect 3470 1031 3471 1035
rect 3475 1031 3476 1035
rect 3470 1030 3476 1031
rect 2694 1025 2700 1026
rect 2694 1021 2695 1025
rect 2699 1021 2700 1025
rect 2694 1020 2700 1021
rect 2862 1025 2868 1026
rect 2862 1021 2863 1025
rect 2867 1021 2868 1025
rect 2862 1020 2868 1021
rect 3022 1025 3028 1026
rect 3022 1021 3023 1025
rect 3027 1021 3028 1025
rect 3022 1020 3028 1021
rect 3182 1025 3188 1026
rect 3182 1021 3183 1025
rect 3187 1021 3188 1025
rect 3182 1020 3188 1021
rect 3342 1025 3348 1026
rect 3342 1021 3343 1025
rect 3347 1021 3348 1025
rect 3342 1020 3348 1021
rect 3110 995 3116 996
rect 3110 991 3111 995
rect 3115 991 3116 995
rect 3110 990 3116 991
rect 2686 985 2692 986
rect 2686 981 2687 985
rect 2691 981 2692 985
rect 2686 980 2692 981
rect 2854 985 2860 986
rect 2854 981 2855 985
rect 2859 981 2860 985
rect 2854 980 2860 981
rect 3014 985 3020 986
rect 3014 981 3015 985
rect 3019 981 3020 985
rect 3014 980 3020 981
rect 2688 971 2690 980
rect 2856 971 2858 980
rect 3016 971 3018 980
rect 2631 970 2635 971
rect 2631 965 2635 966
rect 2687 970 2691 971
rect 2687 965 2691 966
rect 2799 970 2803 971
rect 2799 965 2803 966
rect 2855 970 2859 971
rect 2855 965 2859 966
rect 2951 970 2955 971
rect 2951 965 2955 966
rect 3015 970 3019 971
rect 3015 965 3019 966
rect 3095 970 3099 971
rect 3095 965 3099 966
rect 2632 960 2634 965
rect 2800 960 2802 965
rect 2952 960 2954 965
rect 3096 960 3098 965
rect 2630 959 2636 960
rect 2630 955 2631 959
rect 2635 955 2636 959
rect 2630 954 2636 955
rect 2798 959 2804 960
rect 2798 955 2799 959
rect 2803 955 2804 959
rect 2798 954 2804 955
rect 2950 959 2956 960
rect 2950 955 2951 959
rect 2955 955 2956 959
rect 2950 954 2956 955
rect 3094 959 3100 960
rect 3094 955 3095 959
rect 3099 955 3100 959
rect 3094 954 3100 955
rect 2526 951 2532 952
rect 2526 947 2527 951
rect 2531 947 2532 951
rect 2526 946 2532 947
rect 2174 935 2180 936
rect 2174 931 2175 935
rect 2179 931 2180 935
rect 2174 930 2180 931
rect 2078 919 2084 920
rect 2078 915 2079 919
rect 2083 915 2084 919
rect 2078 914 2084 915
rect 1902 907 1908 908
rect 1902 903 1903 907
rect 1907 903 1908 907
rect 1902 902 1908 903
rect 2080 895 2082 914
rect 1863 894 1867 895
rect 1863 889 1867 890
rect 1895 894 1899 895
rect 1895 889 1899 890
rect 2023 894 2027 895
rect 2023 889 2027 890
rect 2079 894 2083 895
rect 2079 889 2083 890
rect 1002 887 1008 888
rect 1002 883 1003 887
rect 1007 883 1008 887
rect 1002 882 1008 883
rect 1494 887 1500 888
rect 1494 883 1495 887
rect 1499 883 1500 887
rect 1494 882 1500 883
rect 1822 884 1828 885
rect 782 871 788 872
rect 614 866 620 867
rect 707 868 711 869
rect 455 863 459 864
rect 456 860 458 863
rect 454 859 460 860
rect 454 855 455 859
rect 459 855 460 859
rect 616 855 618 866
rect 782 867 783 871
rect 787 867 788 871
rect 782 866 788 867
rect 942 871 948 872
rect 942 867 943 871
rect 947 867 948 871
rect 942 866 948 867
rect 707 863 711 864
rect 784 855 786 866
rect 944 855 946 866
rect 1004 860 1006 882
rect 1102 871 1108 872
rect 1102 867 1103 871
rect 1107 867 1108 871
rect 1102 866 1108 867
rect 1254 871 1260 872
rect 1254 867 1255 871
rect 1259 867 1260 871
rect 1406 871 1412 872
rect 1254 866 1260 867
rect 1263 868 1267 869
rect 1002 859 1008 860
rect 1002 855 1003 859
rect 1007 855 1008 859
rect 1104 855 1106 866
rect 1256 855 1258 866
rect 1406 867 1407 871
rect 1411 867 1412 871
rect 1496 869 1498 882
rect 1822 880 1823 884
rect 1827 880 1828 884
rect 1822 879 1828 880
rect 1558 871 1564 872
rect 1406 866 1412 867
rect 1495 868 1499 869
rect 1263 863 1267 864
rect 1264 860 1266 863
rect 1262 859 1268 860
rect 1262 855 1263 859
rect 1267 855 1268 859
rect 1408 855 1410 866
rect 1558 867 1559 871
rect 1563 867 1564 871
rect 1558 866 1564 867
rect 1495 863 1499 864
rect 1560 855 1562 866
rect 1824 855 1826 879
rect 1864 865 1866 889
rect 1896 878 1898 889
rect 1962 887 1968 888
rect 1962 883 1963 887
rect 1967 883 1968 887
rect 1962 882 1968 883
rect 1894 877 1900 878
rect 1894 873 1895 877
rect 1899 873 1900 877
rect 1894 872 1900 873
rect 1862 864 1868 865
rect 1862 860 1863 864
rect 1867 860 1868 864
rect 1964 860 1966 882
rect 2024 878 2026 889
rect 2176 888 2178 930
rect 2270 919 2276 920
rect 2270 915 2271 919
rect 2275 915 2276 919
rect 2270 914 2276 915
rect 2462 919 2468 920
rect 2462 915 2463 919
rect 2467 915 2468 919
rect 2462 914 2468 915
rect 2638 919 2644 920
rect 2638 915 2639 919
rect 2643 915 2644 919
rect 2638 914 2644 915
rect 2806 919 2812 920
rect 2806 915 2807 919
rect 2811 915 2812 919
rect 2958 919 2964 920
rect 2806 914 2812 915
rect 2815 916 2819 917
rect 2272 895 2274 914
rect 2464 895 2466 914
rect 2640 895 2642 914
rect 2808 895 2810 914
rect 2958 915 2959 919
rect 2963 915 2964 919
rect 2958 914 2964 915
rect 3102 919 3108 920
rect 3102 915 3103 919
rect 3107 915 3108 919
rect 3112 917 3114 990
rect 3174 985 3180 986
rect 3174 981 3175 985
rect 3179 981 3180 985
rect 3174 980 3180 981
rect 3334 985 3340 986
rect 3334 981 3335 985
rect 3339 981 3340 985
rect 3334 980 3340 981
rect 3176 971 3178 980
rect 3336 971 3338 980
rect 3175 970 3179 971
rect 3175 965 3179 966
rect 3231 970 3235 971
rect 3231 965 3235 966
rect 3335 970 3339 971
rect 3335 965 3339 966
rect 3232 960 3234 965
rect 3230 959 3236 960
rect 3230 955 3231 959
rect 3235 955 3236 959
rect 3230 954 3236 955
rect 3352 952 3354 1030
rect 3488 1026 3490 1037
rect 3486 1025 3492 1026
rect 3486 1021 3487 1025
rect 3491 1021 3492 1025
rect 3486 1020 3492 1021
rect 3576 1013 3578 1037
rect 3574 1012 3580 1013
rect 3574 1008 3575 1012
rect 3579 1008 3580 1012
rect 3574 1007 3580 1008
rect 3574 995 3580 996
rect 3574 991 3575 995
rect 3579 991 3580 995
rect 3574 990 3580 991
rect 3478 985 3484 986
rect 3478 981 3479 985
rect 3483 981 3484 985
rect 3478 980 3484 981
rect 3480 971 3482 980
rect 3576 971 3578 990
rect 3367 970 3371 971
rect 3367 965 3371 966
rect 3479 970 3483 971
rect 3479 965 3483 966
rect 3575 970 3579 971
rect 3575 965 3579 966
rect 3368 960 3370 965
rect 3480 960 3482 965
rect 3366 959 3372 960
rect 3366 955 3367 959
rect 3371 955 3372 959
rect 3366 954 3372 955
rect 3478 959 3484 960
rect 3478 955 3479 959
rect 3483 955 3484 959
rect 3478 954 3484 955
rect 3350 951 3356 952
rect 3350 947 3351 951
rect 3355 947 3356 951
rect 3576 950 3578 965
rect 3350 946 3356 947
rect 3574 949 3580 950
rect 3574 945 3575 949
rect 3579 945 3580 949
rect 3574 944 3580 945
rect 3470 935 3476 936
rect 3470 931 3471 935
rect 3475 931 3476 935
rect 3470 930 3476 931
rect 3574 932 3580 933
rect 3238 919 3244 920
rect 3102 914 3108 915
rect 3111 916 3115 917
rect 2815 911 2819 912
rect 2816 908 2818 911
rect 2814 907 2820 908
rect 2814 903 2815 907
rect 2819 903 2820 907
rect 2814 902 2820 903
rect 2960 895 2962 914
rect 3104 895 3106 914
rect 3238 915 3239 919
rect 3243 915 3244 919
rect 3238 914 3244 915
rect 3374 919 3380 920
rect 3374 915 3375 919
rect 3379 915 3380 919
rect 3374 914 3380 915
rect 3111 911 3115 912
rect 3240 895 3242 914
rect 3376 895 3378 914
rect 2183 894 2187 895
rect 2183 889 2187 890
rect 2271 894 2275 895
rect 2271 889 2275 890
rect 2351 894 2355 895
rect 2351 889 2355 890
rect 2463 894 2467 895
rect 2463 889 2467 890
rect 2519 894 2523 895
rect 2519 889 2523 890
rect 2639 894 2643 895
rect 2639 889 2643 890
rect 2687 894 2691 895
rect 2687 889 2691 890
rect 2807 894 2811 895
rect 2807 889 2811 890
rect 2839 894 2843 895
rect 2839 889 2843 890
rect 2959 894 2963 895
rect 2959 889 2963 890
rect 2983 894 2987 895
rect 2983 889 2987 890
rect 3103 894 3107 895
rect 3103 889 3107 890
rect 3119 894 3123 895
rect 3119 889 3123 890
rect 3239 894 3243 895
rect 3239 889 3243 890
rect 3247 894 3251 895
rect 3247 889 3251 890
rect 3375 894 3379 895
rect 3375 889 3379 890
rect 2174 887 2180 888
rect 2174 883 2175 887
rect 2179 883 2180 887
rect 2174 882 2180 883
rect 2184 878 2186 889
rect 2352 878 2354 889
rect 2438 887 2444 888
rect 2438 883 2439 887
rect 2443 883 2444 887
rect 2438 882 2444 883
rect 2022 877 2028 878
rect 2022 873 2023 877
rect 2027 873 2028 877
rect 2022 872 2028 873
rect 2182 877 2188 878
rect 2182 873 2183 877
rect 2187 873 2188 877
rect 2182 872 2188 873
rect 2350 877 2356 878
rect 2350 873 2351 877
rect 2355 873 2356 877
rect 2350 872 2356 873
rect 2440 860 2442 882
rect 2520 878 2522 889
rect 2606 887 2612 888
rect 2606 883 2607 887
rect 2611 883 2612 887
rect 2606 882 2612 883
rect 2518 877 2524 878
rect 2518 873 2519 877
rect 2523 873 2524 877
rect 2518 872 2524 873
rect 2608 860 2610 882
rect 2688 878 2690 889
rect 2694 887 2700 888
rect 2694 883 2695 887
rect 2699 883 2700 887
rect 2694 882 2700 883
rect 2686 877 2692 878
rect 2686 873 2687 877
rect 2691 873 2692 877
rect 2686 872 2692 873
rect 1862 859 1868 860
rect 1962 859 1968 860
rect 1962 855 1963 859
rect 1967 855 1968 859
rect 447 854 451 855
rect 454 854 460 855
rect 463 854 467 855
rect 447 849 451 850
rect 463 849 467 850
rect 615 854 619 855
rect 615 849 619 850
rect 639 854 643 855
rect 639 849 643 850
rect 783 854 787 855
rect 783 849 787 850
rect 807 854 811 855
rect 807 849 811 850
rect 943 854 947 855
rect 943 849 947 850
rect 983 854 987 855
rect 1002 854 1008 855
rect 1103 854 1107 855
rect 983 849 987 850
rect 1103 849 1107 850
rect 1159 854 1163 855
rect 1159 849 1163 850
rect 1255 854 1259 855
rect 1262 854 1268 855
rect 1335 854 1339 855
rect 1255 849 1259 850
rect 1335 849 1339 850
rect 1407 854 1411 855
rect 1407 849 1411 850
rect 1511 854 1515 855
rect 1511 849 1515 850
rect 1559 854 1563 855
rect 1559 849 1563 850
rect 1823 854 1827 855
rect 1962 854 1968 855
rect 2438 859 2444 860
rect 2438 855 2439 859
rect 2443 855 2444 859
rect 2438 854 2444 855
rect 2606 859 2612 860
rect 2606 855 2607 859
rect 2611 855 2612 859
rect 2606 854 2612 855
rect 1823 849 1827 850
rect 338 847 344 848
rect 338 843 339 847
rect 343 843 344 847
rect 338 842 344 843
rect 464 838 466 849
rect 640 838 642 849
rect 808 838 810 849
rect 984 838 986 849
rect 1058 847 1064 848
rect 1058 843 1059 847
rect 1063 843 1064 847
rect 1058 842 1064 843
rect 142 837 148 838
rect 142 833 143 837
rect 147 833 148 837
rect 142 832 148 833
rect 286 837 292 838
rect 286 833 287 837
rect 291 833 292 837
rect 286 832 292 833
rect 462 837 468 838
rect 462 833 463 837
rect 467 833 468 837
rect 462 832 468 833
rect 638 837 644 838
rect 638 833 639 837
rect 643 833 644 837
rect 638 832 644 833
rect 806 837 812 838
rect 806 833 807 837
rect 811 833 812 837
rect 806 832 812 833
rect 982 837 988 838
rect 982 833 983 837
rect 987 833 988 837
rect 982 832 988 833
rect 110 824 116 825
rect 110 820 111 824
rect 115 820 116 824
rect 1060 820 1062 842
rect 1160 838 1162 849
rect 1166 847 1172 848
rect 1166 843 1167 847
rect 1171 843 1172 847
rect 1166 842 1172 843
rect 1158 837 1164 838
rect 1158 833 1159 837
rect 1163 833 1164 837
rect 1158 832 1164 833
rect 110 819 116 820
rect 1058 819 1064 820
rect 1058 815 1059 819
rect 1063 815 1064 819
rect 1058 814 1064 815
rect 110 807 116 808
rect 110 803 111 807
rect 115 803 116 807
rect 110 802 116 803
rect 790 807 796 808
rect 790 803 791 807
rect 795 803 796 807
rect 790 802 796 803
rect 112 783 114 802
rect 134 797 140 798
rect 134 793 135 797
rect 139 793 140 797
rect 134 792 140 793
rect 278 797 284 798
rect 278 793 279 797
rect 283 793 284 797
rect 278 792 284 793
rect 454 797 460 798
rect 454 793 455 797
rect 459 793 460 797
rect 454 792 460 793
rect 630 797 636 798
rect 630 793 631 797
rect 635 793 636 797
rect 630 792 636 793
rect 136 783 138 792
rect 280 783 282 792
rect 456 783 458 792
rect 632 783 634 792
rect 111 782 115 783
rect 111 777 115 778
rect 135 782 139 783
rect 135 777 139 778
rect 271 782 275 783
rect 271 777 275 778
rect 279 782 283 783
rect 279 777 283 778
rect 439 782 443 783
rect 439 777 443 778
rect 455 782 459 783
rect 455 777 459 778
rect 607 782 611 783
rect 607 777 611 778
rect 631 782 635 783
rect 631 777 635 778
rect 775 782 779 783
rect 775 777 779 778
rect 112 762 114 777
rect 136 772 138 777
rect 272 772 274 777
rect 440 772 442 777
rect 608 772 610 777
rect 776 772 778 777
rect 134 771 140 772
rect 134 767 135 771
rect 139 767 140 771
rect 134 766 140 767
rect 270 771 276 772
rect 270 767 271 771
rect 275 767 276 771
rect 270 766 276 767
rect 438 771 444 772
rect 438 767 439 771
rect 443 767 444 771
rect 438 766 444 767
rect 606 771 612 772
rect 606 767 607 771
rect 611 767 612 771
rect 606 766 612 767
rect 774 771 780 772
rect 774 767 775 771
rect 779 767 780 771
rect 774 766 780 767
rect 110 761 116 762
rect 110 757 111 761
rect 115 757 116 761
rect 110 756 116 757
rect 202 747 208 748
rect 110 744 116 745
rect 110 740 111 744
rect 115 740 116 744
rect 202 743 203 747
rect 207 743 208 747
rect 202 742 208 743
rect 506 747 512 748
rect 506 743 507 747
rect 511 743 512 747
rect 506 742 512 743
rect 674 747 680 748
rect 674 743 675 747
rect 679 743 680 747
rect 674 742 680 743
rect 110 739 116 740
rect 112 711 114 739
rect 142 731 148 732
rect 142 727 143 731
rect 147 727 148 731
rect 142 726 148 727
rect 144 711 146 726
rect 204 720 206 742
rect 278 731 284 732
rect 278 727 279 731
rect 283 727 284 731
rect 278 726 284 727
rect 446 731 452 732
rect 446 727 447 731
rect 451 727 452 731
rect 446 726 452 727
rect 202 719 208 720
rect 202 715 203 719
rect 207 715 208 719
rect 202 714 208 715
rect 270 719 276 720
rect 270 715 271 719
rect 275 715 276 719
rect 270 714 276 715
rect 111 710 115 711
rect 111 705 115 706
rect 143 710 147 711
rect 143 705 147 706
rect 112 681 114 705
rect 144 694 146 705
rect 214 703 220 704
rect 214 699 215 703
rect 219 699 220 703
rect 214 698 220 699
rect 142 693 148 694
rect 142 689 143 693
rect 147 689 148 693
rect 142 688 148 689
rect 110 680 116 681
rect 216 680 218 698
rect 110 676 111 680
rect 115 676 116 680
rect 110 675 116 676
rect 214 679 220 680
rect 214 675 215 679
rect 219 675 220 679
rect 272 676 274 714
rect 280 711 282 726
rect 448 711 450 726
rect 508 720 510 742
rect 614 731 620 732
rect 614 727 615 731
rect 619 727 620 731
rect 614 726 620 727
rect 506 719 512 720
rect 506 715 507 719
rect 511 715 512 719
rect 506 714 512 715
rect 616 711 618 726
rect 676 720 678 742
rect 782 731 788 732
rect 782 727 783 731
rect 787 727 788 731
rect 782 726 788 727
rect 674 719 680 720
rect 674 715 675 719
rect 679 715 680 719
rect 674 714 680 715
rect 784 711 786 726
rect 792 720 794 802
rect 798 797 804 798
rect 798 793 799 797
rect 803 793 804 797
rect 798 792 804 793
rect 974 797 980 798
rect 974 793 975 797
rect 979 793 980 797
rect 974 792 980 793
rect 1150 797 1156 798
rect 1150 793 1151 797
rect 1155 793 1156 797
rect 1150 792 1156 793
rect 800 783 802 792
rect 976 783 978 792
rect 1152 783 1154 792
rect 799 782 803 783
rect 799 777 803 778
rect 935 782 939 783
rect 935 777 939 778
rect 975 782 979 783
rect 975 777 979 778
rect 1087 782 1091 783
rect 1087 777 1091 778
rect 1151 782 1155 783
rect 1151 777 1155 778
rect 936 772 938 777
rect 1088 772 1090 777
rect 934 771 940 772
rect 934 767 935 771
rect 939 767 940 771
rect 934 766 940 767
rect 1086 771 1092 772
rect 1086 767 1087 771
rect 1091 767 1092 771
rect 1086 766 1092 767
rect 1168 764 1170 842
rect 1336 838 1338 849
rect 1512 838 1514 849
rect 1334 837 1340 838
rect 1334 833 1335 837
rect 1339 833 1340 837
rect 1334 832 1340 833
rect 1510 837 1516 838
rect 1510 833 1511 837
rect 1515 833 1516 837
rect 1510 832 1516 833
rect 1824 825 1826 849
rect 1862 847 1868 848
rect 1862 843 1863 847
rect 1867 843 1868 847
rect 1862 842 1868 843
rect 1822 824 1828 825
rect 1822 820 1823 824
rect 1827 820 1828 824
rect 1822 819 1828 820
rect 1864 819 1866 842
rect 1886 837 1892 838
rect 1886 833 1887 837
rect 1891 833 1892 837
rect 1886 832 1892 833
rect 2014 837 2020 838
rect 2014 833 2015 837
rect 2019 833 2020 837
rect 2014 832 2020 833
rect 2174 837 2180 838
rect 2174 833 2175 837
rect 2179 833 2180 837
rect 2174 832 2180 833
rect 2342 837 2348 838
rect 2342 833 2343 837
rect 2347 833 2348 837
rect 2342 832 2348 833
rect 2510 837 2516 838
rect 2510 833 2511 837
rect 2515 833 2516 837
rect 2510 832 2516 833
rect 2678 837 2684 838
rect 2678 833 2679 837
rect 2683 833 2684 837
rect 2678 832 2684 833
rect 1888 819 1890 832
rect 2016 819 2018 832
rect 2176 819 2178 832
rect 2344 819 2346 832
rect 2512 819 2514 832
rect 2680 819 2682 832
rect 1863 818 1867 819
rect 1863 813 1867 814
rect 1887 818 1891 819
rect 1887 813 1891 814
rect 2015 818 2019 819
rect 2015 813 2019 814
rect 2071 818 2075 819
rect 2071 813 2075 814
rect 2175 818 2179 819
rect 2175 813 2179 814
rect 2263 818 2267 819
rect 2263 813 2267 814
rect 2343 818 2347 819
rect 2343 813 2347 814
rect 2447 818 2451 819
rect 2447 813 2451 814
rect 2511 818 2515 819
rect 2511 813 2515 814
rect 2623 818 2627 819
rect 2623 813 2627 814
rect 2679 818 2683 819
rect 2679 813 2683 814
rect 1294 807 1300 808
rect 1294 803 1295 807
rect 1299 803 1300 807
rect 1294 802 1300 803
rect 1822 807 1828 808
rect 1822 803 1823 807
rect 1827 803 1828 807
rect 1822 802 1828 803
rect 1239 782 1243 783
rect 1239 777 1243 778
rect 1240 772 1242 777
rect 1238 771 1244 772
rect 1238 767 1239 771
rect 1243 767 1244 771
rect 1238 766 1244 767
rect 1166 763 1172 764
rect 1166 759 1167 763
rect 1171 759 1172 763
rect 1166 758 1172 759
rect 942 731 948 732
rect 942 727 943 731
rect 947 727 948 731
rect 942 726 948 727
rect 1094 731 1100 732
rect 1094 727 1095 731
rect 1099 727 1100 731
rect 1094 726 1100 727
rect 1246 731 1252 732
rect 1246 727 1247 731
rect 1251 727 1252 731
rect 1246 726 1252 727
rect 790 719 796 720
rect 790 715 791 719
rect 795 715 796 719
rect 790 714 796 715
rect 944 711 946 726
rect 1096 711 1098 726
rect 1248 711 1250 726
rect 1296 720 1298 802
rect 1326 797 1332 798
rect 1326 793 1327 797
rect 1331 793 1332 797
rect 1326 792 1332 793
rect 1502 797 1508 798
rect 1502 793 1503 797
rect 1507 793 1508 797
rect 1502 792 1508 793
rect 1328 783 1330 792
rect 1504 783 1506 792
rect 1824 783 1826 802
rect 1864 798 1866 813
rect 1888 808 1890 813
rect 2072 808 2074 813
rect 2264 808 2266 813
rect 2448 808 2450 813
rect 2624 808 2626 813
rect 1886 807 1892 808
rect 1886 803 1887 807
rect 1891 803 1892 807
rect 1886 802 1892 803
rect 2070 807 2076 808
rect 2070 803 2071 807
rect 2075 803 2076 807
rect 2070 802 2076 803
rect 2262 807 2268 808
rect 2262 803 2263 807
rect 2267 803 2268 807
rect 2262 802 2268 803
rect 2446 807 2452 808
rect 2446 803 2447 807
rect 2451 803 2452 807
rect 2446 802 2452 803
rect 2622 807 2628 808
rect 2622 803 2623 807
rect 2627 803 2628 807
rect 2622 802 2628 803
rect 2696 800 2698 882
rect 2840 878 2842 889
rect 2906 887 2912 888
rect 2906 883 2907 887
rect 2911 883 2912 887
rect 2906 882 2912 883
rect 2838 877 2844 878
rect 2838 873 2839 877
rect 2843 873 2844 877
rect 2838 872 2844 873
rect 2908 860 2910 882
rect 2984 878 2986 889
rect 3050 887 3056 888
rect 3050 883 3051 887
rect 3055 883 3056 887
rect 3050 882 3056 883
rect 2982 877 2988 878
rect 2982 873 2983 877
rect 2987 873 2988 877
rect 2982 872 2988 873
rect 3052 860 3054 882
rect 3120 878 3122 889
rect 3198 887 3204 888
rect 3198 883 3199 887
rect 3203 883 3204 887
rect 3198 882 3204 883
rect 3118 877 3124 878
rect 3118 873 3119 877
rect 3123 873 3124 877
rect 3118 872 3124 873
rect 3200 860 3202 882
rect 3248 878 3250 889
rect 3314 887 3320 888
rect 3314 883 3315 887
rect 3319 883 3320 887
rect 3314 882 3320 883
rect 3246 877 3252 878
rect 3246 873 3247 877
rect 3251 873 3252 877
rect 3246 872 3252 873
rect 3316 860 3318 882
rect 3376 878 3378 889
rect 3472 888 3474 930
rect 3574 928 3575 932
rect 3579 928 3580 932
rect 3574 927 3580 928
rect 3486 919 3492 920
rect 3486 915 3487 919
rect 3491 915 3492 919
rect 3486 914 3492 915
rect 3488 895 3490 914
rect 3576 895 3578 927
rect 3487 894 3491 895
rect 3487 889 3491 890
rect 3575 894 3579 895
rect 3575 889 3579 890
rect 3470 887 3476 888
rect 3470 883 3471 887
rect 3475 883 3476 887
rect 3470 882 3476 883
rect 3488 878 3490 889
rect 3374 877 3380 878
rect 3374 873 3375 877
rect 3379 873 3380 877
rect 3374 872 3380 873
rect 3486 877 3492 878
rect 3486 873 3487 877
rect 3491 873 3492 877
rect 3486 872 3492 873
rect 3576 865 3578 889
rect 3574 864 3580 865
rect 3574 860 3575 864
rect 3579 860 3580 864
rect 2906 859 2912 860
rect 2906 855 2907 859
rect 2911 855 2912 859
rect 2906 854 2912 855
rect 3050 859 3056 860
rect 3050 855 3051 859
rect 3055 855 3056 859
rect 3050 854 3056 855
rect 3198 859 3204 860
rect 3198 855 3199 859
rect 3203 855 3204 859
rect 3198 854 3204 855
rect 3314 859 3320 860
rect 3574 859 3580 860
rect 3314 855 3315 859
rect 3319 855 3320 859
rect 3314 854 3320 855
rect 2806 847 2812 848
rect 2806 843 2807 847
rect 2811 843 2812 847
rect 2806 842 2812 843
rect 3574 847 3580 848
rect 3574 843 3575 847
rect 3579 843 3580 847
rect 3574 842 3580 843
rect 2791 818 2795 819
rect 2791 813 2795 814
rect 2792 808 2794 813
rect 2790 807 2796 808
rect 2790 803 2791 807
rect 2795 803 2796 807
rect 2790 802 2796 803
rect 1954 799 1960 800
rect 1862 797 1868 798
rect 1862 793 1863 797
rect 1867 793 1868 797
rect 1954 795 1955 799
rect 1959 795 1960 799
rect 1954 794 1960 795
rect 2694 799 2700 800
rect 2694 795 2695 799
rect 2699 795 2700 799
rect 2694 794 2700 795
rect 1862 792 1868 793
rect 1327 782 1331 783
rect 1327 777 1331 778
rect 1391 782 1395 783
rect 1391 777 1395 778
rect 1503 782 1507 783
rect 1503 777 1507 778
rect 1551 782 1555 783
rect 1551 777 1555 778
rect 1823 782 1827 783
rect 1823 777 1827 778
rect 1862 780 1868 781
rect 1392 772 1394 777
rect 1552 772 1554 777
rect 1390 771 1396 772
rect 1390 767 1391 771
rect 1395 767 1396 771
rect 1390 766 1396 767
rect 1550 771 1556 772
rect 1550 767 1551 771
rect 1555 767 1556 771
rect 1550 766 1556 767
rect 1824 762 1826 777
rect 1862 776 1863 780
rect 1867 776 1868 780
rect 1862 775 1868 776
rect 1822 761 1828 762
rect 1822 757 1823 761
rect 1827 757 1828 761
rect 1822 756 1828 757
rect 1864 751 1866 775
rect 1894 767 1900 768
rect 1894 763 1895 767
rect 1899 763 1900 767
rect 1894 762 1900 763
rect 1896 751 1898 762
rect 1863 750 1867 751
rect 1618 747 1624 748
rect 1618 743 1619 747
rect 1623 743 1624 747
rect 1863 745 1867 746
rect 1895 750 1899 751
rect 1895 745 1899 746
rect 1618 742 1624 743
rect 1822 744 1828 745
rect 1398 731 1404 732
rect 1398 727 1399 731
rect 1403 727 1404 731
rect 1398 726 1404 727
rect 1558 731 1564 732
rect 1558 727 1559 731
rect 1563 727 1564 731
rect 1558 726 1564 727
rect 1294 719 1300 720
rect 1294 715 1295 719
rect 1299 715 1300 719
rect 1294 714 1300 715
rect 1400 711 1402 726
rect 1560 711 1562 726
rect 279 710 283 711
rect 279 705 283 706
rect 287 710 291 711
rect 287 705 291 706
rect 447 710 451 711
rect 447 705 451 706
rect 455 710 459 711
rect 455 705 459 706
rect 615 710 619 711
rect 615 705 619 706
rect 623 710 627 711
rect 623 705 627 706
rect 783 710 787 711
rect 783 705 787 706
rect 791 710 795 711
rect 791 705 795 706
rect 943 710 947 711
rect 943 705 947 706
rect 959 710 963 711
rect 959 705 963 706
rect 1095 710 1099 711
rect 1095 705 1099 706
rect 1119 710 1123 711
rect 1119 705 1123 706
rect 1247 710 1251 711
rect 1247 705 1251 706
rect 1279 710 1283 711
rect 1279 705 1283 706
rect 1399 710 1403 711
rect 1399 705 1403 706
rect 1439 710 1443 711
rect 1439 705 1443 706
rect 1559 710 1563 711
rect 1559 705 1563 706
rect 1599 710 1603 711
rect 1599 705 1603 706
rect 288 694 290 705
rect 456 694 458 705
rect 526 703 532 704
rect 526 699 527 703
rect 531 699 532 703
rect 526 698 532 699
rect 286 693 292 694
rect 286 689 287 693
rect 291 689 292 693
rect 286 688 292 689
rect 454 693 460 694
rect 454 689 455 693
rect 459 689 460 693
rect 454 688 460 689
rect 528 680 530 698
rect 624 694 626 705
rect 710 703 716 704
rect 710 699 711 703
rect 715 699 716 703
rect 710 698 716 699
rect 622 693 628 694
rect 622 689 623 693
rect 627 689 628 693
rect 622 688 628 689
rect 712 680 714 698
rect 792 694 794 705
rect 960 694 962 705
rect 1026 703 1032 704
rect 1026 699 1027 703
rect 1031 699 1032 703
rect 1026 698 1032 699
rect 790 693 796 694
rect 790 689 791 693
rect 795 689 796 693
rect 790 688 796 689
rect 958 693 964 694
rect 958 689 959 693
rect 963 689 964 693
rect 958 688 964 689
rect 526 679 532 680
rect 214 674 220 675
rect 270 675 276 676
rect 270 671 271 675
rect 275 671 276 675
rect 526 675 527 679
rect 531 675 532 679
rect 526 674 532 675
rect 710 679 716 680
rect 710 675 711 679
rect 715 675 716 679
rect 1028 676 1030 698
rect 1120 694 1122 705
rect 1280 694 1282 705
rect 1362 703 1368 704
rect 1362 699 1363 703
rect 1367 699 1368 703
rect 1362 698 1368 699
rect 1118 693 1124 694
rect 1118 689 1119 693
rect 1123 689 1124 693
rect 1118 688 1124 689
rect 1278 693 1284 694
rect 1278 689 1279 693
rect 1283 689 1284 693
rect 1278 688 1284 689
rect 1364 676 1366 698
rect 1440 694 1442 705
rect 1514 703 1520 704
rect 1514 699 1515 703
rect 1519 699 1520 703
rect 1514 698 1520 699
rect 1438 693 1444 694
rect 1438 689 1439 693
rect 1443 689 1444 693
rect 1438 688 1444 689
rect 1516 676 1518 698
rect 1600 694 1602 705
rect 1620 704 1622 742
rect 1822 740 1823 744
rect 1827 740 1828 744
rect 1822 739 1828 740
rect 1824 711 1826 739
rect 1864 721 1866 745
rect 1896 734 1898 745
rect 1956 744 1958 794
rect 2078 767 2084 768
rect 2078 763 2079 767
rect 2083 763 2084 767
rect 2078 762 2084 763
rect 2270 767 2276 768
rect 2270 763 2271 767
rect 2275 763 2276 767
rect 2270 762 2276 763
rect 2454 767 2460 768
rect 2454 763 2455 767
rect 2459 763 2460 767
rect 2454 762 2460 763
rect 2630 767 2636 768
rect 2630 763 2631 767
rect 2635 763 2636 767
rect 2630 762 2636 763
rect 2798 767 2804 768
rect 2798 763 2799 767
rect 2803 763 2804 767
rect 2798 762 2804 763
rect 2080 751 2082 762
rect 2254 755 2260 756
rect 2254 751 2255 755
rect 2259 751 2260 755
rect 2272 751 2274 762
rect 2456 751 2458 762
rect 2632 751 2634 762
rect 2800 751 2802 762
rect 2808 756 2810 842
rect 2830 837 2836 838
rect 2830 833 2831 837
rect 2835 833 2836 837
rect 2830 832 2836 833
rect 2974 837 2980 838
rect 2974 833 2975 837
rect 2979 833 2980 837
rect 2974 832 2980 833
rect 3110 837 3116 838
rect 3110 833 3111 837
rect 3115 833 3116 837
rect 3110 832 3116 833
rect 3238 837 3244 838
rect 3238 833 3239 837
rect 3243 833 3244 837
rect 3238 832 3244 833
rect 3366 837 3372 838
rect 3366 833 3367 837
rect 3371 833 3372 837
rect 3366 832 3372 833
rect 3478 837 3484 838
rect 3478 833 3479 837
rect 3483 833 3484 837
rect 3478 832 3484 833
rect 2832 819 2834 832
rect 2976 819 2978 832
rect 3112 819 3114 832
rect 3240 819 3242 832
rect 3368 819 3370 832
rect 3480 819 3482 832
rect 3576 819 3578 842
rect 2831 818 2835 819
rect 2831 813 2835 814
rect 2943 818 2947 819
rect 2943 813 2947 814
rect 2975 818 2979 819
rect 2975 813 2979 814
rect 3087 818 3091 819
rect 3087 813 3091 814
rect 3111 818 3115 819
rect 3111 813 3115 814
rect 3223 818 3227 819
rect 3223 813 3227 814
rect 3239 818 3243 819
rect 3239 813 3243 814
rect 3359 818 3363 819
rect 3359 813 3363 814
rect 3367 818 3371 819
rect 3367 813 3371 814
rect 3479 818 3483 819
rect 3479 813 3483 814
rect 3575 818 3579 819
rect 3575 813 3579 814
rect 2944 808 2946 813
rect 3088 808 3090 813
rect 3224 808 3226 813
rect 3360 808 3362 813
rect 3480 808 3482 813
rect 2942 807 2948 808
rect 2942 803 2943 807
rect 2947 803 2948 807
rect 2942 802 2948 803
rect 3086 807 3092 808
rect 3086 803 3087 807
rect 3091 803 3092 807
rect 3086 802 3092 803
rect 3222 807 3228 808
rect 3222 803 3223 807
rect 3227 803 3228 807
rect 3222 802 3228 803
rect 3358 807 3364 808
rect 3358 803 3359 807
rect 3363 803 3364 807
rect 3358 802 3364 803
rect 3478 807 3484 808
rect 3478 803 3479 807
rect 3483 803 3484 807
rect 3478 802 3484 803
rect 3576 798 3578 813
rect 3574 797 3580 798
rect 3574 793 3575 797
rect 3579 793 3580 797
rect 3574 792 3580 793
rect 3158 783 3164 784
rect 3158 779 3159 783
rect 3163 779 3164 783
rect 3158 778 3164 779
rect 3426 783 3432 784
rect 3426 779 3427 783
rect 3431 779 3432 783
rect 3426 778 3432 779
rect 3574 780 3580 781
rect 2950 767 2956 768
rect 2950 763 2951 767
rect 2955 763 2956 767
rect 2950 762 2956 763
rect 3094 767 3100 768
rect 3094 763 3095 767
rect 3099 763 3100 767
rect 3094 762 3100 763
rect 2806 755 2812 756
rect 2806 751 2807 755
rect 2811 751 2812 755
rect 2952 751 2954 762
rect 3096 751 3098 762
rect 2071 750 2075 751
rect 2071 745 2075 746
rect 2079 750 2083 751
rect 2254 750 2260 751
rect 2263 750 2267 751
rect 2079 745 2083 746
rect 1954 743 1960 744
rect 1954 739 1955 743
rect 1959 739 1960 743
rect 1954 738 1960 739
rect 2072 734 2074 745
rect 1894 733 1900 734
rect 1894 729 1895 733
rect 1899 729 1900 733
rect 1894 728 1900 729
rect 2070 733 2076 734
rect 2070 729 2071 733
rect 2075 729 2076 733
rect 2070 728 2076 729
rect 1862 720 1868 721
rect 1862 716 1863 720
rect 1867 716 1868 720
rect 2256 716 2258 750
rect 2263 745 2267 746
rect 2271 750 2275 751
rect 2271 745 2275 746
rect 2447 750 2451 751
rect 2447 745 2451 746
rect 2455 750 2459 751
rect 2455 745 2459 746
rect 2623 750 2627 751
rect 2623 745 2627 746
rect 2631 750 2635 751
rect 2631 745 2635 746
rect 2799 750 2803 751
rect 2806 750 2812 751
rect 2951 750 2955 751
rect 2799 745 2803 746
rect 2951 745 2955 746
rect 2975 750 2979 751
rect 2975 745 2979 746
rect 3095 750 3099 751
rect 3095 745 3099 746
rect 3151 750 3155 751
rect 3151 745 3155 746
rect 2264 734 2266 745
rect 2374 743 2380 744
rect 2374 739 2375 743
rect 2379 739 2380 743
rect 2374 738 2380 739
rect 2262 733 2268 734
rect 2262 729 2263 733
rect 2267 729 2268 733
rect 2262 728 2268 729
rect 2376 716 2378 738
rect 2448 734 2450 745
rect 2462 743 2468 744
rect 2462 739 2463 743
rect 2467 739 2468 743
rect 2462 738 2468 739
rect 2446 733 2452 734
rect 2446 729 2447 733
rect 2451 729 2452 733
rect 2446 728 2452 729
rect 1862 715 1868 716
rect 2254 715 2260 716
rect 2254 711 2255 715
rect 2259 711 2260 715
rect 1823 710 1827 711
rect 2254 710 2260 711
rect 2374 715 2380 716
rect 2374 711 2375 715
rect 2379 711 2380 715
rect 2374 710 2380 711
rect 1823 705 1827 706
rect 1618 703 1624 704
rect 1618 699 1619 703
rect 1623 699 1624 703
rect 1618 698 1624 699
rect 1598 693 1604 694
rect 1598 689 1599 693
rect 1603 689 1604 693
rect 1598 688 1604 689
rect 1824 681 1826 705
rect 1862 703 1868 704
rect 1862 699 1863 703
rect 1867 699 1868 703
rect 1862 698 1868 699
rect 1822 680 1828 681
rect 1822 676 1823 680
rect 1827 676 1828 680
rect 1864 679 1866 698
rect 1886 693 1892 694
rect 1886 689 1887 693
rect 1891 689 1892 693
rect 1886 688 1892 689
rect 2062 693 2068 694
rect 2062 689 2063 693
rect 2067 689 2068 693
rect 2062 688 2068 689
rect 2254 693 2260 694
rect 2254 689 2255 693
rect 2259 689 2260 693
rect 2254 688 2260 689
rect 2438 693 2444 694
rect 2438 689 2439 693
rect 2443 689 2444 693
rect 2438 688 2444 689
rect 1888 679 1890 688
rect 2064 679 2066 688
rect 2110 687 2116 688
rect 2110 683 2111 687
rect 2115 683 2116 687
rect 2110 682 2116 683
rect 710 674 716 675
rect 1026 675 1032 676
rect 270 670 276 671
rect 1026 671 1027 675
rect 1031 671 1032 675
rect 1026 670 1032 671
rect 1362 675 1368 676
rect 1362 671 1363 675
rect 1367 671 1368 675
rect 1362 670 1368 671
rect 1514 675 1520 676
rect 1822 675 1828 676
rect 1863 678 1867 679
rect 1514 671 1515 675
rect 1519 671 1520 675
rect 1863 673 1867 674
rect 1887 678 1891 679
rect 1887 673 1891 674
rect 1975 678 1979 679
rect 1975 673 1979 674
rect 2063 678 2067 679
rect 2063 673 2067 674
rect 2095 678 2099 679
rect 2095 673 2099 674
rect 1514 670 1520 671
rect 110 663 116 664
rect 110 659 111 663
rect 115 659 116 663
rect 110 658 116 659
rect 790 663 796 664
rect 790 659 791 663
rect 795 659 796 663
rect 790 658 796 659
rect 1822 663 1828 664
rect 1822 659 1823 663
rect 1827 659 1828 663
rect 1822 658 1828 659
rect 1864 658 1866 673
rect 1888 668 1890 673
rect 1976 668 1978 673
rect 2096 668 2098 673
rect 1886 667 1892 668
rect 1886 663 1887 667
rect 1891 663 1892 667
rect 1886 662 1892 663
rect 1974 667 1980 668
rect 1974 663 1975 667
rect 1979 663 1980 667
rect 1974 662 1980 663
rect 2094 667 2100 668
rect 2094 663 2095 667
rect 2099 663 2100 667
rect 2094 662 2100 663
rect 112 635 114 658
rect 134 653 140 654
rect 134 649 135 653
rect 139 649 140 653
rect 134 648 140 649
rect 278 653 284 654
rect 278 649 279 653
rect 283 649 284 653
rect 278 648 284 649
rect 446 653 452 654
rect 446 649 447 653
rect 451 649 452 653
rect 446 648 452 649
rect 614 653 620 654
rect 614 649 615 653
rect 619 649 620 653
rect 614 648 620 649
rect 782 653 788 654
rect 782 649 783 653
rect 787 649 788 653
rect 782 648 788 649
rect 136 635 138 648
rect 280 635 282 648
rect 448 635 450 648
rect 616 635 618 648
rect 784 635 786 648
rect 111 634 115 635
rect 111 629 115 630
rect 135 634 139 635
rect 135 629 139 630
rect 279 634 283 635
rect 279 629 283 630
rect 287 634 291 635
rect 287 629 291 630
rect 447 634 451 635
rect 447 629 451 630
rect 455 634 459 635
rect 455 629 459 630
rect 615 634 619 635
rect 615 629 619 630
rect 631 634 635 635
rect 631 629 635 630
rect 783 634 787 635
rect 783 629 787 630
rect 112 614 114 629
rect 136 624 138 629
rect 288 624 290 629
rect 456 624 458 629
rect 632 624 634 629
rect 134 623 140 624
rect 134 619 135 623
rect 139 619 140 623
rect 134 618 140 619
rect 286 623 292 624
rect 286 619 287 623
rect 291 619 292 623
rect 286 618 292 619
rect 454 623 460 624
rect 454 619 455 623
rect 459 619 460 623
rect 454 618 460 619
rect 630 623 636 624
rect 630 619 631 623
rect 635 619 636 623
rect 630 618 636 619
rect 110 613 116 614
rect 110 609 111 613
rect 115 609 116 613
rect 110 608 116 609
rect 202 599 208 600
rect 110 596 116 597
rect 110 592 111 596
rect 115 592 116 596
rect 202 595 203 599
rect 207 595 208 599
rect 202 594 208 595
rect 522 599 528 600
rect 522 595 523 599
rect 527 595 528 599
rect 522 594 528 595
rect 698 599 704 600
rect 698 595 699 599
rect 703 595 704 599
rect 698 594 704 595
rect 110 591 116 592
rect 112 563 114 591
rect 142 583 148 584
rect 142 579 143 583
rect 147 579 148 583
rect 142 578 148 579
rect 144 563 146 578
rect 204 572 206 594
rect 294 583 300 584
rect 294 579 295 583
rect 299 579 300 583
rect 294 578 300 579
rect 462 583 468 584
rect 462 579 463 583
rect 467 579 468 583
rect 462 578 468 579
rect 202 571 208 572
rect 202 567 203 571
rect 207 567 208 571
rect 202 566 208 567
rect 296 563 298 578
rect 464 563 466 578
rect 524 572 526 594
rect 638 583 644 584
rect 638 579 639 583
rect 643 579 644 583
rect 638 578 644 579
rect 522 571 528 572
rect 522 567 523 571
rect 527 567 528 571
rect 522 566 528 567
rect 640 563 642 578
rect 700 572 702 594
rect 792 572 794 658
rect 950 653 956 654
rect 950 649 951 653
rect 955 649 956 653
rect 950 648 956 649
rect 1110 653 1116 654
rect 1110 649 1111 653
rect 1115 649 1116 653
rect 1110 648 1116 649
rect 1270 653 1276 654
rect 1270 649 1271 653
rect 1275 649 1276 653
rect 1270 648 1276 649
rect 1430 653 1436 654
rect 1430 649 1431 653
rect 1435 649 1436 653
rect 1430 648 1436 649
rect 1590 653 1596 654
rect 1590 649 1591 653
rect 1595 649 1596 653
rect 1590 648 1596 649
rect 952 635 954 648
rect 1112 635 1114 648
rect 1272 635 1274 648
rect 1432 635 1434 648
rect 1592 635 1594 648
rect 1824 635 1826 658
rect 1862 657 1868 658
rect 1862 653 1863 657
rect 1867 653 1868 657
rect 1862 652 1868 653
rect 1954 643 1960 644
rect 1862 640 1868 641
rect 1862 636 1863 640
rect 1867 636 1868 640
rect 1954 639 1955 643
rect 1959 639 1960 643
rect 1954 638 1960 639
rect 2042 643 2048 644
rect 2042 639 2043 643
rect 2047 639 2048 643
rect 2042 638 2048 639
rect 1862 635 1868 636
rect 799 634 803 635
rect 799 629 803 630
rect 951 634 955 635
rect 951 629 955 630
rect 967 634 971 635
rect 967 629 971 630
rect 1111 634 1115 635
rect 1111 629 1115 630
rect 1119 634 1123 635
rect 1119 629 1123 630
rect 1271 634 1275 635
rect 1271 629 1275 630
rect 1415 634 1419 635
rect 1415 629 1419 630
rect 1431 634 1435 635
rect 1431 629 1435 630
rect 1559 634 1563 635
rect 1559 629 1563 630
rect 1591 634 1595 635
rect 1591 629 1595 630
rect 1711 634 1715 635
rect 1711 629 1715 630
rect 1823 634 1827 635
rect 1823 629 1827 630
rect 800 624 802 629
rect 968 624 970 629
rect 1120 624 1122 629
rect 1272 624 1274 629
rect 1416 624 1418 629
rect 1560 624 1562 629
rect 1712 624 1714 629
rect 798 623 804 624
rect 798 619 799 623
rect 803 619 804 623
rect 798 618 804 619
rect 966 623 972 624
rect 966 619 967 623
rect 971 619 972 623
rect 966 618 972 619
rect 1118 623 1124 624
rect 1118 619 1119 623
rect 1123 619 1124 623
rect 1118 618 1124 619
rect 1270 623 1276 624
rect 1270 619 1271 623
rect 1275 619 1276 623
rect 1270 618 1276 619
rect 1414 623 1420 624
rect 1414 619 1415 623
rect 1419 619 1420 623
rect 1414 618 1420 619
rect 1558 623 1564 624
rect 1558 619 1559 623
rect 1563 619 1564 623
rect 1558 618 1564 619
rect 1710 623 1716 624
rect 1710 619 1711 623
rect 1715 619 1716 623
rect 1710 618 1716 619
rect 1638 615 1644 616
rect 1638 611 1639 615
rect 1643 611 1644 615
rect 1824 614 1826 629
rect 1638 610 1644 611
rect 1822 613 1828 614
rect 1640 589 1642 610
rect 1822 609 1823 613
rect 1827 609 1828 613
rect 1822 608 1828 609
rect 1864 607 1866 635
rect 1894 627 1900 628
rect 1894 623 1895 627
rect 1899 623 1900 627
rect 1894 622 1900 623
rect 1896 607 1898 622
rect 1956 616 1958 638
rect 1982 627 1988 628
rect 1982 623 1983 627
rect 1987 623 1988 627
rect 1982 622 1988 623
rect 1954 615 1960 616
rect 1954 611 1955 615
rect 1959 611 1960 615
rect 1954 610 1960 611
rect 1984 607 1986 622
rect 2044 616 2046 638
rect 2102 627 2108 628
rect 2102 623 2103 627
rect 2107 623 2108 627
rect 2102 622 2108 623
rect 2042 615 2048 616
rect 2042 611 2043 615
rect 2047 611 2048 615
rect 2042 610 2048 611
rect 2104 607 2106 622
rect 2112 616 2114 682
rect 2256 679 2258 688
rect 2440 679 2442 688
rect 2223 678 2227 679
rect 2223 673 2227 674
rect 2255 678 2259 679
rect 2255 673 2259 674
rect 2351 678 2355 679
rect 2351 673 2355 674
rect 2439 678 2443 679
rect 2439 673 2443 674
rect 2224 668 2226 673
rect 2352 668 2354 673
rect 2222 667 2228 668
rect 2222 663 2223 667
rect 2227 663 2228 667
rect 2222 662 2228 663
rect 2350 667 2356 668
rect 2350 663 2351 667
rect 2355 663 2356 667
rect 2350 662 2356 663
rect 2464 660 2466 738
rect 2624 734 2626 745
rect 2646 743 2652 744
rect 2646 739 2647 743
rect 2651 739 2652 743
rect 2646 738 2652 739
rect 2622 733 2628 734
rect 2622 729 2623 733
rect 2627 729 2628 733
rect 2622 728 2628 729
rect 2614 693 2620 694
rect 2614 689 2615 693
rect 2619 689 2620 693
rect 2614 688 2620 689
rect 2648 688 2650 738
rect 2800 734 2802 745
rect 2976 734 2978 745
rect 3054 743 3060 744
rect 3054 738 3055 743
rect 3059 738 3060 743
rect 3055 735 3059 736
rect 3152 734 3154 745
rect 3160 744 3162 778
rect 3230 767 3236 768
rect 3230 763 3231 767
rect 3235 763 3236 767
rect 3230 762 3236 763
rect 3366 767 3372 768
rect 3366 763 3367 767
rect 3371 763 3372 767
rect 3366 762 3372 763
rect 3232 751 3234 762
rect 3368 751 3370 762
rect 3231 750 3235 751
rect 3231 745 3235 746
rect 3327 750 3331 751
rect 3327 745 3331 746
rect 3367 750 3371 751
rect 3428 748 3430 778
rect 3574 776 3575 780
rect 3579 776 3580 780
rect 3574 775 3580 776
rect 3486 767 3492 768
rect 3486 763 3487 767
rect 3491 763 3492 767
rect 3486 762 3492 763
rect 3488 751 3490 762
rect 3576 751 3578 775
rect 3487 750 3491 751
rect 3367 745 3371 746
rect 3426 747 3432 748
rect 3158 743 3164 744
rect 3158 739 3159 743
rect 3163 739 3164 743
rect 3158 738 3164 739
rect 3259 740 3263 741
rect 3259 735 3263 736
rect 2798 733 2804 734
rect 2798 729 2799 733
rect 2803 729 2804 733
rect 2798 728 2804 729
rect 2974 733 2980 734
rect 2974 729 2975 733
rect 2979 729 2980 733
rect 2974 728 2980 729
rect 3150 733 3156 734
rect 3150 729 3151 733
rect 3155 729 3156 733
rect 3150 728 3156 729
rect 3260 716 3262 735
rect 3328 734 3330 745
rect 3426 743 3427 747
rect 3431 743 3432 747
rect 3487 745 3491 746
rect 3575 750 3579 751
rect 3575 745 3579 746
rect 3426 742 3432 743
rect 3488 734 3490 745
rect 3326 733 3332 734
rect 3326 729 3327 733
rect 3331 729 3332 733
rect 3326 728 3332 729
rect 3486 733 3492 734
rect 3486 729 3487 733
rect 3491 729 3492 733
rect 3486 728 3492 729
rect 3576 721 3578 745
rect 3574 720 3580 721
rect 3574 716 3575 720
rect 3579 716 3580 720
rect 3258 715 3264 716
rect 3574 715 3580 716
rect 3258 711 3259 715
rect 3263 711 3264 715
rect 3258 710 3264 711
rect 3574 703 3580 704
rect 3574 699 3575 703
rect 3579 699 3580 703
rect 3574 698 3580 699
rect 2790 693 2796 694
rect 2790 689 2791 693
rect 2795 689 2796 693
rect 2790 688 2796 689
rect 2966 693 2972 694
rect 2966 689 2967 693
rect 2971 689 2972 693
rect 2966 688 2972 689
rect 3142 693 3148 694
rect 3142 689 3143 693
rect 3147 689 3148 693
rect 3142 688 3148 689
rect 3318 693 3324 694
rect 3318 689 3319 693
rect 3323 689 3324 693
rect 3318 688 3324 689
rect 3478 693 3484 694
rect 3478 689 3479 693
rect 3483 689 3484 693
rect 3478 688 3484 689
rect 2616 679 2618 688
rect 2646 687 2652 688
rect 2646 683 2647 687
rect 2651 683 2652 687
rect 2646 682 2652 683
rect 2792 679 2794 688
rect 2968 679 2970 688
rect 3144 679 3146 688
rect 3320 679 3322 688
rect 3480 679 3482 688
rect 3576 679 3578 698
rect 2479 678 2483 679
rect 2479 673 2483 674
rect 2615 678 2619 679
rect 2615 673 2619 674
rect 2767 678 2771 679
rect 2767 673 2771 674
rect 2791 678 2795 679
rect 2791 673 2795 674
rect 2935 678 2939 679
rect 2935 673 2939 674
rect 2967 678 2971 679
rect 2967 673 2971 674
rect 3119 678 3123 679
rect 3119 673 3123 674
rect 3143 678 3147 679
rect 3143 673 3147 674
rect 3311 678 3315 679
rect 3311 673 3315 674
rect 3319 678 3323 679
rect 3319 673 3323 674
rect 3479 678 3483 679
rect 3479 673 3483 674
rect 3575 678 3579 679
rect 3575 673 3579 674
rect 2480 668 2482 673
rect 2616 668 2618 673
rect 2768 668 2770 673
rect 2936 668 2938 673
rect 3120 668 3122 673
rect 3312 668 3314 673
rect 3480 668 3482 673
rect 2478 667 2484 668
rect 2478 663 2479 667
rect 2483 663 2484 667
rect 2478 662 2484 663
rect 2614 667 2620 668
rect 2614 663 2615 667
rect 2619 663 2620 667
rect 2614 662 2620 663
rect 2766 667 2772 668
rect 2766 663 2767 667
rect 2771 663 2772 667
rect 2766 662 2772 663
rect 2934 667 2940 668
rect 2934 663 2935 667
rect 2939 663 2940 667
rect 2934 662 2940 663
rect 3118 667 3124 668
rect 3118 663 3119 667
rect 3123 663 3124 667
rect 3118 662 3124 663
rect 3310 667 3316 668
rect 3310 663 3311 667
rect 3315 663 3316 667
rect 3310 662 3316 663
rect 3478 667 3484 668
rect 3478 663 3479 667
rect 3483 663 3484 667
rect 3478 662 3484 663
rect 2462 659 2468 660
rect 2462 655 2463 659
rect 2467 655 2468 659
rect 3576 658 3578 673
rect 2462 654 2468 655
rect 3574 657 3580 658
rect 3574 653 3575 657
rect 3579 653 3580 657
rect 3574 652 3580 653
rect 2834 643 2840 644
rect 2834 639 2835 643
rect 2839 639 2840 643
rect 2834 638 2840 639
rect 3226 643 3232 644
rect 3226 639 3227 643
rect 3231 639 3232 643
rect 3226 638 3232 639
rect 3234 643 3240 644
rect 3234 639 3235 643
rect 3239 639 3240 643
rect 3234 638 3240 639
rect 3470 643 3476 644
rect 3470 639 3471 643
rect 3475 639 3476 643
rect 3470 638 3476 639
rect 3574 640 3580 641
rect 2230 627 2236 628
rect 2230 623 2231 627
rect 2235 623 2236 627
rect 2230 622 2236 623
rect 2358 627 2364 628
rect 2358 623 2359 627
rect 2363 623 2364 627
rect 2358 622 2364 623
rect 2486 627 2492 628
rect 2486 623 2487 627
rect 2491 623 2492 627
rect 2486 622 2492 623
rect 2622 627 2628 628
rect 2622 623 2623 627
rect 2627 623 2628 627
rect 2622 622 2628 623
rect 2774 627 2780 628
rect 2774 623 2775 627
rect 2779 623 2780 627
rect 2774 622 2780 623
rect 2110 615 2116 616
rect 2110 611 2111 615
rect 2115 611 2116 615
rect 2110 610 2116 611
rect 2206 615 2212 616
rect 2206 611 2207 615
rect 2211 611 2212 615
rect 2206 610 2212 611
rect 1863 606 1867 607
rect 1863 601 1867 602
rect 1895 606 1899 607
rect 1895 601 1899 602
rect 1983 606 1987 607
rect 1983 601 1987 602
rect 2047 606 2051 607
rect 2047 601 2051 602
rect 2103 606 2107 607
rect 2103 601 2107 602
rect 1822 596 1828 597
rect 1822 592 1823 596
rect 1827 592 1828 596
rect 1822 591 1828 592
rect 1199 588 1203 589
rect 1639 588 1643 589
rect 806 583 812 584
rect 806 579 807 583
rect 811 579 812 583
rect 806 578 812 579
rect 974 583 980 584
rect 974 579 975 583
rect 979 579 980 583
rect 974 578 980 579
rect 1126 583 1132 584
rect 1199 583 1203 584
rect 1278 583 1284 584
rect 1126 579 1127 583
rect 1131 579 1132 583
rect 1126 578 1132 579
rect 698 571 704 572
rect 698 567 699 571
rect 703 567 704 571
rect 698 566 704 567
rect 790 571 796 572
rect 790 567 791 571
rect 795 567 796 571
rect 790 566 796 567
rect 808 563 810 578
rect 976 563 978 578
rect 986 571 992 572
rect 986 567 987 571
rect 991 567 992 571
rect 986 566 992 567
rect 111 562 115 563
rect 111 557 115 558
rect 143 562 147 563
rect 143 557 147 558
rect 151 562 155 563
rect 151 557 155 558
rect 295 562 299 563
rect 295 557 299 558
rect 311 562 315 563
rect 311 557 315 558
rect 463 562 467 563
rect 463 557 467 558
rect 471 562 475 563
rect 471 557 475 558
rect 631 562 635 563
rect 631 557 635 558
rect 639 562 643 563
rect 639 557 643 558
rect 783 562 787 563
rect 783 557 787 558
rect 807 562 811 563
rect 807 557 811 558
rect 927 562 931 563
rect 927 557 931 558
rect 975 562 979 563
rect 975 557 979 558
rect 112 533 114 557
rect 152 546 154 557
rect 312 546 314 557
rect 472 546 474 557
rect 632 546 634 557
rect 784 546 786 557
rect 928 546 930 557
rect 150 545 156 546
rect 150 541 151 545
rect 155 541 156 545
rect 150 540 156 541
rect 310 545 316 546
rect 310 541 311 545
rect 315 541 316 545
rect 310 540 316 541
rect 470 545 476 546
rect 470 541 471 545
rect 475 541 476 545
rect 470 540 476 541
rect 630 545 636 546
rect 630 541 631 545
rect 635 541 636 545
rect 630 540 636 541
rect 782 545 788 546
rect 782 541 783 545
rect 787 541 788 545
rect 782 540 788 541
rect 926 545 932 546
rect 926 541 927 545
rect 931 541 932 545
rect 926 540 932 541
rect 110 532 116 533
rect 988 532 990 566
rect 1128 563 1130 578
rect 1063 562 1067 563
rect 1063 557 1067 558
rect 1127 562 1131 563
rect 1127 557 1131 558
rect 1191 562 1195 563
rect 1191 557 1195 558
rect 994 555 1000 556
rect 994 551 995 555
rect 999 551 1000 555
rect 994 550 1000 551
rect 110 528 111 532
rect 115 528 116 532
rect 110 527 116 528
rect 986 531 992 532
rect 986 527 987 531
rect 991 527 992 531
rect 996 528 998 550
rect 1064 546 1066 557
rect 1074 555 1080 556
rect 1074 551 1075 555
rect 1079 551 1080 555
rect 1074 550 1080 551
rect 1062 545 1068 546
rect 1062 541 1063 545
rect 1067 541 1068 545
rect 1062 540 1068 541
rect 986 526 992 527
rect 994 527 1000 528
rect 994 523 995 527
rect 999 523 1000 527
rect 994 522 1000 523
rect 110 515 116 516
rect 110 511 111 515
rect 115 511 116 515
rect 110 510 116 511
rect 782 515 788 516
rect 782 511 783 515
rect 787 511 788 515
rect 782 510 788 511
rect 112 487 114 510
rect 142 505 148 506
rect 142 501 143 505
rect 147 501 148 505
rect 142 500 148 501
rect 302 505 308 506
rect 302 501 303 505
rect 307 501 308 505
rect 302 500 308 501
rect 462 505 468 506
rect 462 501 463 505
rect 467 501 468 505
rect 462 500 468 501
rect 622 505 628 506
rect 622 501 623 505
rect 627 501 628 505
rect 622 500 628 501
rect 774 505 780 506
rect 774 501 775 505
rect 779 501 780 505
rect 774 500 780 501
rect 144 487 146 500
rect 304 487 306 500
rect 464 487 466 500
rect 624 487 626 500
rect 776 487 778 500
rect 111 486 115 487
rect 111 481 115 482
rect 143 486 147 487
rect 143 481 147 482
rect 159 486 163 487
rect 159 481 163 482
rect 303 486 307 487
rect 303 481 307 482
rect 311 486 315 487
rect 311 481 315 482
rect 463 486 467 487
rect 463 481 467 482
rect 615 486 619 487
rect 615 481 619 482
rect 623 486 627 487
rect 623 481 627 482
rect 759 486 763 487
rect 759 481 763 482
rect 775 486 779 487
rect 775 481 779 482
rect 112 466 114 481
rect 160 476 162 481
rect 312 476 314 481
rect 464 476 466 481
rect 616 476 618 481
rect 760 476 762 481
rect 158 475 164 476
rect 158 471 159 475
rect 163 471 164 475
rect 158 470 164 471
rect 310 475 316 476
rect 310 471 311 475
rect 315 471 316 475
rect 310 470 316 471
rect 462 475 468 476
rect 462 471 463 475
rect 467 471 468 475
rect 462 470 468 471
rect 614 475 620 476
rect 614 471 615 475
rect 619 471 620 475
rect 614 470 620 471
rect 758 475 764 476
rect 758 471 759 475
rect 763 471 764 475
rect 758 470 764 471
rect 110 465 116 466
rect 110 461 111 465
rect 115 461 116 465
rect 110 460 116 461
rect 542 451 548 452
rect 110 448 116 449
rect 110 444 111 448
rect 115 444 116 448
rect 542 447 543 451
rect 547 447 548 451
rect 542 446 548 447
rect 698 451 704 452
rect 698 447 699 451
rect 703 447 704 451
rect 698 446 704 447
rect 110 443 116 444
rect 112 419 114 443
rect 166 435 172 436
rect 166 431 167 435
rect 171 431 172 435
rect 166 430 172 431
rect 318 435 324 436
rect 318 431 319 435
rect 323 431 324 435
rect 318 430 324 431
rect 470 435 476 436
rect 470 431 471 435
rect 475 431 476 435
rect 470 430 476 431
rect 168 419 170 430
rect 320 419 322 430
rect 330 423 336 424
rect 330 419 331 423
rect 335 419 336 423
rect 472 419 474 430
rect 111 418 115 419
rect 111 413 115 414
rect 151 418 155 419
rect 151 413 155 414
rect 167 418 171 419
rect 167 413 171 414
rect 271 418 275 419
rect 271 413 275 414
rect 319 418 323 419
rect 330 418 336 419
rect 407 418 411 419
rect 319 413 323 414
rect 112 389 114 413
rect 152 402 154 413
rect 158 411 164 412
rect 158 407 159 411
rect 163 407 164 411
rect 158 406 164 407
rect 150 401 156 402
rect 150 397 151 401
rect 155 397 156 401
rect 150 396 156 397
rect 160 389 162 406
rect 272 402 274 413
rect 270 401 276 402
rect 270 397 271 401
rect 275 397 276 401
rect 270 396 276 397
rect 110 388 116 389
rect 110 384 111 388
rect 115 384 116 388
rect 110 383 116 384
rect 159 388 163 389
rect 332 388 334 418
rect 407 413 411 414
rect 471 418 475 419
rect 471 413 475 414
rect 408 402 410 413
rect 544 412 546 446
rect 622 435 628 436
rect 622 431 623 435
rect 627 431 628 435
rect 622 430 628 431
rect 624 419 626 430
rect 700 424 702 446
rect 766 435 772 436
rect 766 431 767 435
rect 771 431 772 435
rect 766 430 772 431
rect 698 423 704 424
rect 698 419 699 423
rect 703 419 704 423
rect 768 419 770 430
rect 784 424 786 510
rect 918 505 924 506
rect 918 501 919 505
rect 923 501 924 505
rect 918 500 924 501
rect 1054 505 1060 506
rect 1054 501 1055 505
rect 1059 501 1060 505
rect 1054 500 1060 501
rect 920 487 922 500
rect 1056 487 1058 500
rect 887 486 891 487
rect 887 481 891 482
rect 919 486 923 487
rect 919 481 923 482
rect 1007 486 1011 487
rect 1007 481 1011 482
rect 1055 486 1059 487
rect 1055 481 1059 482
rect 888 476 890 481
rect 1008 476 1010 481
rect 886 475 892 476
rect 886 471 887 475
rect 891 471 892 475
rect 886 470 892 471
rect 1006 475 1012 476
rect 1006 471 1007 475
rect 1011 471 1012 475
rect 1006 470 1012 471
rect 1076 468 1078 550
rect 1192 546 1194 557
rect 1200 556 1202 583
rect 1278 579 1279 583
rect 1283 579 1284 583
rect 1278 578 1284 579
rect 1422 583 1428 584
rect 1422 579 1423 583
rect 1427 579 1428 583
rect 1422 578 1428 579
rect 1566 583 1572 584
rect 1639 583 1643 584
rect 1718 583 1724 584
rect 1566 579 1567 583
rect 1571 579 1572 583
rect 1566 578 1572 579
rect 1718 579 1719 583
rect 1723 579 1724 583
rect 1718 578 1724 579
rect 1280 563 1282 578
rect 1424 563 1426 578
rect 1568 563 1570 578
rect 1720 563 1722 578
rect 1824 563 1826 591
rect 1864 577 1866 601
rect 1896 590 1898 601
rect 2048 590 2050 601
rect 2054 599 2060 600
rect 2054 595 2055 599
rect 2059 595 2060 599
rect 2054 594 2060 595
rect 1894 589 1900 590
rect 1894 585 1895 589
rect 1899 585 1900 589
rect 1894 584 1900 585
rect 2046 589 2052 590
rect 2046 585 2047 589
rect 2051 585 2052 589
rect 2046 584 2052 585
rect 1862 576 1868 577
rect 1862 572 1863 576
rect 1867 572 1868 576
rect 1862 571 1868 572
rect 1279 562 1283 563
rect 1279 557 1283 558
rect 1311 562 1315 563
rect 1311 557 1315 558
rect 1423 562 1427 563
rect 1423 557 1427 558
rect 1535 562 1539 563
rect 1535 557 1539 558
rect 1567 562 1571 563
rect 1567 557 1571 558
rect 1647 562 1651 563
rect 1647 557 1651 558
rect 1719 562 1723 563
rect 1719 557 1723 558
rect 1735 562 1739 563
rect 1735 557 1739 558
rect 1823 562 1827 563
rect 1823 557 1827 558
rect 1862 559 1868 560
rect 1198 555 1204 556
rect 1198 551 1199 555
rect 1203 551 1204 555
rect 1198 550 1204 551
rect 1312 546 1314 557
rect 1424 546 1426 557
rect 1536 546 1538 557
rect 1602 555 1608 556
rect 1602 551 1603 555
rect 1607 551 1608 555
rect 1602 550 1608 551
rect 1190 545 1196 546
rect 1190 541 1191 545
rect 1195 541 1196 545
rect 1190 540 1196 541
rect 1310 545 1316 546
rect 1310 541 1311 545
rect 1315 541 1316 545
rect 1310 540 1316 541
rect 1422 545 1428 546
rect 1422 541 1423 545
rect 1427 541 1428 545
rect 1422 540 1428 541
rect 1534 545 1540 546
rect 1534 541 1535 545
rect 1539 541 1540 545
rect 1534 540 1540 541
rect 1604 528 1606 550
rect 1648 546 1650 557
rect 1670 555 1676 556
rect 1670 551 1671 555
rect 1675 551 1676 555
rect 1670 550 1676 551
rect 1646 545 1652 546
rect 1646 541 1647 545
rect 1651 541 1652 545
rect 1646 540 1652 541
rect 1602 527 1608 528
rect 1602 523 1603 527
rect 1607 523 1608 527
rect 1602 522 1608 523
rect 1490 515 1496 516
rect 1490 511 1491 515
rect 1495 511 1496 515
rect 1490 510 1496 511
rect 1182 505 1188 506
rect 1182 501 1183 505
rect 1187 501 1188 505
rect 1182 500 1188 501
rect 1302 505 1308 506
rect 1302 501 1303 505
rect 1307 501 1308 505
rect 1302 500 1308 501
rect 1414 505 1420 506
rect 1414 501 1415 505
rect 1419 501 1420 505
rect 1414 500 1420 501
rect 1184 487 1186 500
rect 1304 487 1306 500
rect 1416 487 1418 500
rect 1454 499 1460 500
rect 1454 495 1455 499
rect 1459 495 1460 499
rect 1454 494 1460 495
rect 1127 486 1131 487
rect 1127 481 1131 482
rect 1183 486 1187 487
rect 1183 481 1187 482
rect 1239 486 1243 487
rect 1239 481 1243 482
rect 1303 486 1307 487
rect 1303 481 1307 482
rect 1343 486 1347 487
rect 1343 481 1347 482
rect 1415 486 1419 487
rect 1415 481 1419 482
rect 1439 486 1443 487
rect 1439 481 1443 482
rect 1128 476 1130 481
rect 1240 476 1242 481
rect 1344 476 1346 481
rect 1440 476 1442 481
rect 1126 475 1132 476
rect 1126 471 1127 475
rect 1131 471 1132 475
rect 1126 470 1132 471
rect 1238 475 1244 476
rect 1238 471 1239 475
rect 1243 471 1244 475
rect 1238 470 1244 471
rect 1342 475 1348 476
rect 1342 471 1343 475
rect 1347 471 1348 475
rect 1342 470 1348 471
rect 1438 475 1444 476
rect 1438 471 1439 475
rect 1443 471 1444 475
rect 1438 470 1444 471
rect 1074 467 1080 468
rect 1074 463 1075 467
rect 1079 463 1080 467
rect 1074 462 1080 463
rect 1430 451 1436 452
rect 1430 447 1431 451
rect 1435 447 1436 451
rect 1430 446 1436 447
rect 894 435 900 436
rect 894 431 895 435
rect 899 431 900 435
rect 894 430 900 431
rect 1014 435 1020 436
rect 1014 431 1015 435
rect 1019 431 1020 435
rect 1014 430 1020 431
rect 1134 435 1140 436
rect 1134 431 1135 435
rect 1139 431 1140 435
rect 1134 430 1140 431
rect 1246 435 1252 436
rect 1246 431 1247 435
rect 1251 431 1252 435
rect 1246 430 1252 431
rect 1350 435 1356 436
rect 1350 431 1351 435
rect 1355 431 1356 435
rect 1350 430 1356 431
rect 782 423 788 424
rect 782 419 783 423
rect 787 419 788 423
rect 896 419 898 430
rect 902 423 908 424
rect 902 419 903 423
rect 907 419 908 423
rect 1016 419 1018 430
rect 1136 419 1138 430
rect 1143 428 1147 429
rect 1142 423 1148 424
rect 1142 419 1143 423
rect 1147 419 1148 423
rect 1248 419 1250 430
rect 1352 419 1354 430
rect 551 418 555 419
rect 551 413 555 414
rect 623 418 627 419
rect 698 418 704 419
rect 711 418 715 419
rect 623 413 627 414
rect 711 413 715 414
rect 767 418 771 419
rect 782 418 788 419
rect 887 418 891 419
rect 767 413 771 414
rect 887 413 891 414
rect 895 418 899 419
rect 902 418 908 419
rect 1015 418 1019 419
rect 895 413 899 414
rect 542 411 548 412
rect 542 407 543 411
rect 547 407 548 411
rect 542 406 548 407
rect 552 402 554 413
rect 646 411 652 412
rect 646 407 647 411
rect 651 407 652 411
rect 646 406 652 407
rect 406 401 412 402
rect 406 397 407 401
rect 411 397 412 401
rect 406 396 412 397
rect 550 401 556 402
rect 550 397 551 401
rect 555 397 556 401
rect 550 396 556 397
rect 339 388 343 389
rect 648 388 650 406
rect 712 402 714 413
rect 888 402 890 413
rect 710 401 716 402
rect 710 397 711 401
rect 715 397 716 401
rect 710 396 716 397
rect 886 401 892 402
rect 886 397 887 401
rect 891 397 892 401
rect 904 397 906 418
rect 1015 413 1019 414
rect 1063 418 1067 419
rect 1063 413 1067 414
rect 1135 418 1139 419
rect 1142 418 1148 419
rect 1247 418 1251 419
rect 1135 413 1139 414
rect 1247 413 1251 414
rect 1351 418 1355 419
rect 1351 413 1355 414
rect 1064 402 1066 413
rect 1082 411 1088 412
rect 1082 407 1083 411
rect 1087 407 1088 411
rect 1082 406 1088 407
rect 1062 401 1068 402
rect 1062 397 1063 401
rect 1067 397 1068 401
rect 886 396 892 397
rect 903 396 907 397
rect 1062 396 1068 397
rect 903 391 907 392
rect 159 383 163 384
rect 330 387 336 388
rect 330 383 331 387
rect 335 383 336 387
rect 646 387 652 388
rect 330 382 336 383
rect 338 383 344 384
rect 338 379 339 383
rect 343 379 344 383
rect 646 383 647 387
rect 651 383 652 387
rect 646 382 652 383
rect 338 378 344 379
rect 110 371 116 372
rect 110 367 111 371
rect 115 367 116 371
rect 110 366 116 367
rect 854 371 860 372
rect 854 367 855 371
rect 859 367 860 371
rect 854 366 860 367
rect 112 335 114 366
rect 142 361 148 362
rect 142 357 143 361
rect 147 357 148 361
rect 142 356 148 357
rect 262 361 268 362
rect 262 357 263 361
rect 267 357 268 361
rect 262 356 268 357
rect 398 361 404 362
rect 398 357 399 361
rect 403 357 404 361
rect 398 356 404 357
rect 542 361 548 362
rect 542 357 543 361
rect 547 357 548 361
rect 542 356 548 357
rect 702 361 708 362
rect 702 357 703 361
rect 707 357 708 361
rect 702 356 708 357
rect 144 335 146 356
rect 264 335 266 356
rect 400 335 402 356
rect 544 335 546 356
rect 704 335 706 356
rect 111 334 115 335
rect 111 329 115 330
rect 135 334 139 335
rect 135 329 139 330
rect 143 334 147 335
rect 143 329 147 330
rect 223 334 227 335
rect 223 329 227 330
rect 263 334 267 335
rect 263 329 267 330
rect 311 334 315 335
rect 311 329 315 330
rect 399 334 403 335
rect 399 329 403 330
rect 487 334 491 335
rect 487 329 491 330
rect 543 334 547 335
rect 543 329 547 330
rect 575 334 579 335
rect 575 329 579 330
rect 663 334 667 335
rect 663 329 667 330
rect 703 334 707 335
rect 703 329 707 330
rect 751 334 755 335
rect 751 329 755 330
rect 839 334 843 335
rect 839 329 843 330
rect 112 314 114 329
rect 136 324 138 329
rect 224 324 226 329
rect 312 324 314 329
rect 400 324 402 329
rect 488 324 490 329
rect 576 324 578 329
rect 664 324 666 329
rect 752 324 754 329
rect 840 324 842 329
rect 134 323 140 324
rect 134 319 135 323
rect 139 319 140 323
rect 134 318 140 319
rect 222 323 228 324
rect 222 319 223 323
rect 227 319 228 323
rect 222 318 228 319
rect 310 323 316 324
rect 310 319 311 323
rect 315 319 316 323
rect 310 318 316 319
rect 398 323 404 324
rect 398 319 399 323
rect 403 319 404 323
rect 398 318 404 319
rect 486 323 492 324
rect 486 319 487 323
rect 491 319 492 323
rect 486 318 492 319
rect 574 323 580 324
rect 574 319 575 323
rect 579 319 580 323
rect 574 318 580 319
rect 662 323 668 324
rect 662 319 663 323
rect 667 319 668 323
rect 662 318 668 319
rect 750 323 756 324
rect 750 319 751 323
rect 755 319 756 323
rect 750 318 756 319
rect 838 323 844 324
rect 838 319 839 323
rect 843 319 844 323
rect 838 318 844 319
rect 730 315 736 316
rect 110 313 116 314
rect 110 309 111 313
rect 115 309 116 313
rect 730 311 731 315
rect 735 311 736 315
rect 730 310 736 311
rect 110 308 116 309
rect 110 296 116 297
rect 110 292 111 296
rect 115 292 116 296
rect 110 291 116 292
rect 112 263 114 291
rect 142 283 148 284
rect 142 279 143 283
rect 147 279 148 283
rect 142 278 148 279
rect 230 283 236 284
rect 230 279 231 283
rect 235 279 236 283
rect 230 278 236 279
rect 318 283 324 284
rect 318 279 319 283
rect 323 279 324 283
rect 318 278 324 279
rect 406 283 412 284
rect 406 279 407 283
rect 411 279 412 283
rect 406 278 412 279
rect 494 283 500 284
rect 494 279 495 283
rect 499 279 500 283
rect 494 278 500 279
rect 582 283 588 284
rect 582 279 583 283
rect 587 279 588 283
rect 582 278 588 279
rect 670 283 676 284
rect 670 279 671 283
rect 675 279 676 283
rect 670 278 676 279
rect 134 271 140 272
rect 134 267 135 271
rect 139 267 140 271
rect 134 266 140 267
rect 111 262 115 263
rect 111 257 115 258
rect 112 233 114 257
rect 110 232 116 233
rect 110 228 111 232
rect 115 228 116 232
rect 136 228 138 266
rect 144 263 146 278
rect 232 263 234 278
rect 320 263 322 278
rect 408 263 410 278
rect 496 263 498 278
rect 584 263 586 278
rect 672 263 674 278
rect 732 264 734 310
rect 818 299 824 300
rect 818 295 819 299
rect 823 295 824 299
rect 818 294 824 295
rect 758 283 764 284
rect 758 279 759 283
rect 763 279 764 283
rect 758 278 764 279
rect 730 263 736 264
rect 143 262 147 263
rect 143 257 147 258
rect 231 262 235 263
rect 231 257 235 258
rect 319 262 323 263
rect 319 257 323 258
rect 407 262 411 263
rect 407 257 411 258
rect 495 262 499 263
rect 495 257 499 258
rect 583 262 587 263
rect 583 257 587 258
rect 671 262 675 263
rect 730 259 731 263
rect 735 259 736 263
rect 730 258 736 259
rect 738 263 744 264
rect 760 263 762 278
rect 820 272 822 294
rect 846 283 852 284
rect 846 279 847 283
rect 851 279 852 283
rect 846 278 852 279
rect 818 271 824 272
rect 818 267 819 271
rect 823 267 824 271
rect 818 266 824 267
rect 848 263 850 278
rect 856 272 858 366
rect 878 361 884 362
rect 878 357 879 361
rect 883 357 884 361
rect 878 356 884 357
rect 1054 361 1060 362
rect 1054 357 1055 361
rect 1059 357 1060 361
rect 1054 356 1060 357
rect 880 335 882 356
rect 1056 335 1058 356
rect 879 334 883 335
rect 879 329 883 330
rect 927 334 931 335
rect 927 329 931 330
rect 1015 334 1019 335
rect 1015 329 1019 330
rect 1055 334 1059 335
rect 1055 329 1059 330
rect 928 324 930 329
rect 1016 324 1018 329
rect 926 323 932 324
rect 926 319 927 323
rect 931 319 932 323
rect 926 318 932 319
rect 1014 323 1020 324
rect 1014 319 1015 323
rect 1019 319 1020 323
rect 1014 318 1020 319
rect 1084 316 1086 406
rect 1248 402 1250 413
rect 1432 412 1434 446
rect 1446 435 1452 436
rect 1446 431 1447 435
rect 1451 431 1452 435
rect 1446 430 1452 431
rect 1448 419 1450 430
rect 1456 424 1458 494
rect 1492 429 1494 510
rect 1526 505 1532 506
rect 1526 501 1527 505
rect 1531 501 1532 505
rect 1526 500 1532 501
rect 1638 505 1644 506
rect 1638 501 1639 505
rect 1643 501 1644 505
rect 1638 500 1644 501
rect 1528 487 1530 500
rect 1640 487 1642 500
rect 1672 492 1674 550
rect 1736 546 1738 557
rect 1734 545 1740 546
rect 1734 541 1735 545
rect 1739 541 1740 545
rect 1734 540 1740 541
rect 1824 533 1826 557
rect 1862 555 1863 559
rect 1867 555 1868 559
rect 1862 554 1868 555
rect 1822 532 1828 533
rect 1822 528 1823 532
rect 1827 528 1828 532
rect 1864 531 1866 554
rect 1886 549 1892 550
rect 1886 545 1887 549
rect 1891 545 1892 549
rect 1886 544 1892 545
rect 2038 549 2044 550
rect 2038 545 2039 549
rect 2043 545 2044 549
rect 2038 544 2044 545
rect 1888 531 1890 544
rect 2040 531 2042 544
rect 1822 527 1828 528
rect 1863 530 1867 531
rect 1863 525 1867 526
rect 1887 530 1891 531
rect 1887 525 1891 526
rect 2039 530 2043 531
rect 2056 528 2058 594
rect 2208 572 2210 610
rect 2232 607 2234 622
rect 2360 607 2362 622
rect 2488 607 2490 622
rect 2624 607 2626 622
rect 2631 620 2635 621
rect 2630 615 2636 616
rect 2630 611 2631 615
rect 2635 611 2636 615
rect 2630 610 2636 611
rect 2776 607 2778 622
rect 2215 606 2219 607
rect 2215 601 2219 602
rect 2231 606 2235 607
rect 2231 601 2235 602
rect 2359 606 2363 607
rect 2359 601 2363 602
rect 2391 606 2395 607
rect 2391 601 2395 602
rect 2487 606 2491 607
rect 2487 601 2491 602
rect 2583 606 2587 607
rect 2583 601 2587 602
rect 2623 606 2627 607
rect 2623 601 2627 602
rect 2775 606 2779 607
rect 2775 601 2779 602
rect 2799 606 2803 607
rect 2799 601 2803 602
rect 2216 590 2218 601
rect 2392 590 2394 601
rect 2584 590 2586 601
rect 2800 590 2802 601
rect 2836 600 2838 638
rect 2942 627 2948 628
rect 2942 623 2943 627
rect 2947 623 2948 627
rect 2942 622 2948 623
rect 3126 627 3132 628
rect 3126 623 3127 627
rect 3131 623 3132 627
rect 3126 622 3132 623
rect 2944 607 2946 622
rect 3128 607 3130 622
rect 3228 616 3230 638
rect 3236 621 3238 638
rect 3318 627 3324 628
rect 3318 623 3319 627
rect 3323 623 3324 627
rect 3318 622 3324 623
rect 3235 620 3239 621
rect 3226 615 3232 616
rect 3235 615 3239 616
rect 3226 611 3227 615
rect 3231 611 3232 615
rect 3226 610 3232 611
rect 3320 607 3322 622
rect 2943 606 2947 607
rect 2943 601 2947 602
rect 3023 606 3027 607
rect 3023 601 3027 602
rect 3127 606 3131 607
rect 3127 601 3131 602
rect 3255 606 3259 607
rect 3255 601 3259 602
rect 3319 606 3323 607
rect 3319 601 3323 602
rect 2834 599 2840 600
rect 2834 595 2835 599
rect 2839 595 2840 599
rect 2834 594 2840 595
rect 3024 590 3026 601
rect 3256 590 3258 601
rect 3472 600 3474 638
rect 3574 636 3575 640
rect 3579 636 3580 640
rect 3574 635 3580 636
rect 3486 627 3492 628
rect 3486 623 3487 627
rect 3491 623 3492 627
rect 3486 622 3492 623
rect 3488 607 3490 622
rect 3576 607 3578 635
rect 3487 606 3491 607
rect 3487 601 3491 602
rect 3575 606 3579 607
rect 3575 601 3579 602
rect 3470 599 3476 600
rect 3470 595 3471 599
rect 3475 595 3476 599
rect 3470 594 3476 595
rect 3488 590 3490 601
rect 2214 589 2220 590
rect 2214 585 2215 589
rect 2219 585 2220 589
rect 2214 584 2220 585
rect 2390 589 2396 590
rect 2390 585 2391 589
rect 2395 585 2396 589
rect 2390 584 2396 585
rect 2582 589 2588 590
rect 2582 585 2583 589
rect 2587 585 2588 589
rect 2582 584 2588 585
rect 2798 589 2804 590
rect 2798 585 2799 589
rect 2803 585 2804 589
rect 2798 584 2804 585
rect 3022 589 3028 590
rect 3022 585 3023 589
rect 3027 585 3028 589
rect 3022 584 3028 585
rect 3254 589 3260 590
rect 3254 585 3255 589
rect 3259 585 3260 589
rect 3254 584 3260 585
rect 3486 589 3492 590
rect 3486 585 3487 589
rect 3491 585 3492 589
rect 3486 584 3492 585
rect 3576 577 3578 601
rect 3574 576 3580 577
rect 3574 572 3575 576
rect 3579 572 3580 576
rect 2206 571 2212 572
rect 3574 571 3580 572
rect 2206 567 2207 571
rect 2211 567 2212 571
rect 2206 566 2212 567
rect 3574 559 3580 560
rect 3574 555 3575 559
rect 3579 555 3580 559
rect 3574 554 3580 555
rect 2206 549 2212 550
rect 2206 545 2207 549
rect 2211 545 2212 549
rect 2206 544 2212 545
rect 2382 549 2388 550
rect 2382 545 2383 549
rect 2387 545 2388 549
rect 2382 544 2388 545
rect 2574 549 2580 550
rect 2574 545 2575 549
rect 2579 545 2580 549
rect 2574 544 2580 545
rect 2790 549 2796 550
rect 2790 545 2791 549
rect 2795 545 2796 549
rect 2790 544 2796 545
rect 3014 549 3020 550
rect 3014 545 3015 549
rect 3019 545 3020 549
rect 3014 544 3020 545
rect 3246 549 3252 550
rect 3246 545 3247 549
rect 3251 545 3252 549
rect 3246 544 3252 545
rect 3478 549 3484 550
rect 3478 545 3479 549
rect 3483 545 3484 549
rect 3478 544 3484 545
rect 2208 531 2210 544
rect 2384 531 2386 544
rect 2576 531 2578 544
rect 2792 531 2794 544
rect 3016 531 3018 544
rect 3248 531 3250 544
rect 3480 531 3482 544
rect 3576 531 3578 554
rect 2191 530 2195 531
rect 2039 525 2043 526
rect 2054 527 2060 528
rect 1822 515 1828 516
rect 1822 511 1823 515
rect 1827 511 1828 515
rect 1822 510 1828 511
rect 1864 510 1866 525
rect 2054 523 2055 527
rect 2059 523 2060 527
rect 2191 525 2195 526
rect 2207 530 2211 531
rect 2207 525 2211 526
rect 2279 530 2283 531
rect 2279 525 2283 526
rect 2375 530 2379 531
rect 2375 525 2379 526
rect 2383 530 2387 531
rect 2383 525 2387 526
rect 2487 530 2491 531
rect 2487 525 2491 526
rect 2575 530 2579 531
rect 2575 525 2579 526
rect 2631 530 2635 531
rect 2631 525 2635 526
rect 2791 530 2795 531
rect 2791 525 2795 526
rect 2807 530 2811 531
rect 2807 525 2811 526
rect 3007 530 3011 531
rect 3007 525 3011 526
rect 3015 530 3019 531
rect 3015 525 3019 526
rect 3215 530 3219 531
rect 3215 525 3219 526
rect 3247 530 3251 531
rect 3247 525 3251 526
rect 3431 530 3435 531
rect 3431 525 3435 526
rect 3479 530 3483 531
rect 3479 525 3483 526
rect 3575 530 3579 531
rect 3575 525 3579 526
rect 2054 522 2060 523
rect 2192 520 2194 525
rect 2280 520 2282 525
rect 2376 520 2378 525
rect 2488 520 2490 525
rect 2632 520 2634 525
rect 2808 520 2810 525
rect 3008 520 3010 525
rect 3216 520 3218 525
rect 3432 520 3434 525
rect 2190 519 2196 520
rect 2190 515 2191 519
rect 2195 515 2196 519
rect 2190 514 2196 515
rect 2278 519 2284 520
rect 2278 515 2279 519
rect 2283 515 2284 519
rect 2278 514 2284 515
rect 2374 519 2380 520
rect 2374 515 2375 519
rect 2379 515 2380 519
rect 2374 514 2380 515
rect 2486 519 2492 520
rect 2486 515 2487 519
rect 2491 515 2492 519
rect 2486 514 2492 515
rect 2630 519 2636 520
rect 2630 515 2631 519
rect 2635 515 2636 519
rect 2630 514 2636 515
rect 2806 519 2812 520
rect 2806 515 2807 519
rect 2811 515 2812 519
rect 2806 514 2812 515
rect 3006 519 3012 520
rect 3006 515 3007 519
rect 3011 515 3012 519
rect 3006 514 3012 515
rect 3214 519 3220 520
rect 3214 515 3215 519
rect 3219 515 3220 519
rect 3214 514 3220 515
rect 3430 519 3436 520
rect 3430 515 3431 519
rect 3435 515 3436 519
rect 3430 514 3436 515
rect 3576 510 3578 525
rect 1726 505 1732 506
rect 1726 501 1727 505
rect 1731 501 1732 505
rect 1726 500 1732 501
rect 1670 491 1676 492
rect 1670 487 1671 491
rect 1675 487 1676 491
rect 1728 487 1730 500
rect 1824 487 1826 510
rect 1862 509 1868 510
rect 1862 505 1863 509
rect 1867 505 1868 509
rect 1862 504 1868 505
rect 3574 509 3580 510
rect 3574 505 3575 509
rect 3579 505 3580 509
rect 3574 504 3580 505
rect 2346 495 2352 496
rect 1862 492 1868 493
rect 1862 488 1863 492
rect 1867 488 1868 492
rect 2346 491 2347 495
rect 2351 491 2352 495
rect 3186 495 3192 496
rect 2346 490 2352 491
rect 2391 492 2395 493
rect 1862 487 1868 488
rect 1527 486 1531 487
rect 1527 481 1531 482
rect 1543 486 1547 487
rect 1543 481 1547 482
rect 1639 486 1643 487
rect 1670 486 1676 487
rect 1727 486 1731 487
rect 1639 481 1643 482
rect 1727 481 1731 482
rect 1823 486 1827 487
rect 1823 481 1827 482
rect 1544 476 1546 481
rect 1640 476 1642 481
rect 1728 476 1730 481
rect 1542 475 1548 476
rect 1542 471 1543 475
rect 1547 471 1548 475
rect 1542 470 1548 471
rect 1638 475 1644 476
rect 1638 471 1639 475
rect 1643 471 1644 475
rect 1638 470 1644 471
rect 1726 475 1732 476
rect 1726 471 1727 475
rect 1731 471 1732 475
rect 1726 470 1732 471
rect 1824 466 1826 481
rect 1822 465 1828 466
rect 1822 461 1823 465
rect 1827 461 1828 465
rect 1822 460 1828 461
rect 1864 455 1866 487
rect 2198 479 2204 480
rect 2198 475 2199 479
rect 2203 475 2204 479
rect 2198 474 2204 475
rect 2286 479 2292 480
rect 2286 475 2287 479
rect 2291 475 2292 479
rect 2286 474 2292 475
rect 2200 455 2202 474
rect 2288 455 2290 474
rect 2348 468 2350 490
rect 3186 490 3187 495
rect 2391 487 2395 488
rect 3191 490 3192 495
rect 3498 495 3504 496
rect 3498 491 3499 495
rect 3503 491 3504 495
rect 3498 490 3504 491
rect 3574 492 3580 493
rect 3187 487 3191 488
rect 2382 479 2388 480
rect 2382 475 2383 479
rect 2387 475 2388 479
rect 2382 474 2388 475
rect 2346 467 2352 468
rect 2346 463 2347 467
rect 2351 463 2352 467
rect 2346 462 2352 463
rect 2384 455 2386 474
rect 1863 454 1867 455
rect 1863 449 1867 450
rect 1895 454 1899 455
rect 1895 449 1899 450
rect 2039 454 2043 455
rect 2039 449 2043 450
rect 2199 454 2203 455
rect 2199 449 2203 450
rect 2207 454 2211 455
rect 2207 449 2211 450
rect 2287 454 2291 455
rect 2287 449 2291 450
rect 2383 454 2387 455
rect 2383 449 2387 450
rect 1822 448 1828 449
rect 1822 444 1823 448
rect 1827 444 1828 448
rect 1822 443 1828 444
rect 1550 435 1556 436
rect 1550 431 1551 435
rect 1555 431 1556 435
rect 1550 430 1556 431
rect 1646 435 1652 436
rect 1646 431 1647 435
rect 1651 431 1652 435
rect 1646 430 1652 431
rect 1734 435 1740 436
rect 1734 431 1735 435
rect 1739 431 1740 435
rect 1734 430 1740 431
rect 1491 428 1495 429
rect 1454 423 1460 424
rect 1491 423 1495 424
rect 1454 419 1455 423
rect 1459 419 1460 423
rect 1552 419 1554 430
rect 1648 419 1650 430
rect 1736 419 1738 430
rect 1824 419 1826 443
rect 1864 425 1866 449
rect 1896 438 1898 449
rect 2040 438 2042 449
rect 2208 438 2210 449
rect 2218 447 2224 448
rect 2218 443 2219 447
rect 2223 443 2224 447
rect 2218 442 2224 443
rect 1894 437 1900 438
rect 1894 433 1895 437
rect 1899 433 1900 437
rect 1894 432 1900 433
rect 2038 437 2044 438
rect 2038 433 2039 437
rect 2043 433 2044 437
rect 2038 432 2044 433
rect 2206 437 2212 438
rect 2206 433 2207 437
rect 2211 433 2212 437
rect 2206 432 2212 433
rect 1862 424 1868 425
rect 1862 420 1863 424
rect 1867 420 1868 424
rect 1862 419 1868 420
rect 1439 418 1443 419
rect 1439 413 1443 414
rect 1447 418 1451 419
rect 1454 418 1460 419
rect 1551 418 1555 419
rect 1447 413 1451 414
rect 1551 413 1555 414
rect 1639 418 1643 419
rect 1639 413 1643 414
rect 1647 418 1651 419
rect 1647 413 1651 414
rect 1735 418 1739 419
rect 1735 413 1739 414
rect 1823 418 1827 419
rect 1823 413 1827 414
rect 1430 411 1436 412
rect 1430 407 1431 411
rect 1435 407 1436 411
rect 1430 406 1436 407
rect 1440 402 1442 413
rect 1640 402 1642 413
rect 1246 401 1252 402
rect 1246 397 1247 401
rect 1251 397 1252 401
rect 1163 396 1167 397
rect 1246 396 1252 397
rect 1438 401 1444 402
rect 1438 397 1439 401
rect 1443 397 1444 401
rect 1438 396 1444 397
rect 1638 401 1644 402
rect 1638 397 1639 401
rect 1643 397 1644 401
rect 1638 396 1644 397
rect 1163 391 1167 392
rect 1164 384 1166 391
rect 1824 389 1826 413
rect 1862 407 1868 408
rect 1862 403 1863 407
rect 1867 403 1868 407
rect 1862 402 1868 403
rect 1822 388 1828 389
rect 1822 384 1823 388
rect 1827 384 1828 388
rect 1864 387 1866 402
rect 1886 397 1892 398
rect 1886 393 1887 397
rect 1891 393 1892 397
rect 1886 392 1892 393
rect 2030 397 2036 398
rect 2030 393 2031 397
rect 2035 393 2036 397
rect 2030 392 2036 393
rect 2198 397 2204 398
rect 2198 393 2199 397
rect 2203 393 2204 397
rect 2198 392 2204 393
rect 1888 387 1890 392
rect 2032 387 2034 392
rect 2200 387 2202 392
rect 1162 383 1168 384
rect 1822 383 1828 384
rect 1863 386 1867 387
rect 1162 379 1163 383
rect 1167 379 1168 383
rect 1863 381 1867 382
rect 1887 386 1891 387
rect 1975 386 1979 387
rect 1887 381 1891 382
rect 1902 383 1908 384
rect 1162 378 1168 379
rect 1822 371 1828 372
rect 1822 367 1823 371
rect 1827 367 1828 371
rect 1822 366 1828 367
rect 1864 366 1866 381
rect 1888 376 1890 381
rect 1902 379 1903 383
rect 1907 379 1908 383
rect 1975 381 1979 382
rect 2031 386 2035 387
rect 2031 381 2035 382
rect 2063 386 2067 387
rect 2063 381 2067 382
rect 2151 386 2155 387
rect 2151 381 2155 382
rect 2199 386 2203 387
rect 2199 381 2203 382
rect 1902 378 1908 379
rect 1886 375 1892 376
rect 1886 371 1887 375
rect 1891 371 1892 375
rect 1886 370 1892 371
rect 1238 361 1244 362
rect 1238 357 1239 361
rect 1243 357 1244 361
rect 1238 356 1244 357
rect 1430 361 1436 362
rect 1430 357 1431 361
rect 1435 357 1436 361
rect 1430 356 1436 357
rect 1630 361 1636 362
rect 1630 357 1631 361
rect 1635 357 1636 361
rect 1630 356 1636 357
rect 1240 335 1242 356
rect 1432 335 1434 356
rect 1632 335 1634 356
rect 1824 335 1826 366
rect 1862 365 1868 366
rect 1862 361 1863 365
rect 1867 361 1868 365
rect 1862 360 1868 361
rect 1862 348 1868 349
rect 1862 344 1863 348
rect 1867 344 1868 348
rect 1862 343 1868 344
rect 1103 334 1107 335
rect 1103 329 1107 330
rect 1191 334 1195 335
rect 1191 329 1195 330
rect 1239 334 1243 335
rect 1239 329 1243 330
rect 1287 334 1291 335
rect 1287 329 1291 330
rect 1383 334 1387 335
rect 1383 329 1387 330
rect 1431 334 1435 335
rect 1431 329 1435 330
rect 1479 334 1483 335
rect 1479 329 1483 330
rect 1575 334 1579 335
rect 1575 329 1579 330
rect 1631 334 1635 335
rect 1631 329 1635 330
rect 1671 334 1675 335
rect 1671 329 1675 330
rect 1823 334 1827 335
rect 1823 329 1827 330
rect 1104 324 1106 329
rect 1192 324 1194 329
rect 1288 324 1290 329
rect 1384 324 1386 329
rect 1480 324 1482 329
rect 1576 324 1578 329
rect 1672 324 1674 329
rect 1102 323 1108 324
rect 1102 319 1103 323
rect 1107 319 1108 323
rect 1102 318 1108 319
rect 1190 323 1196 324
rect 1190 319 1191 323
rect 1195 319 1196 323
rect 1190 318 1196 319
rect 1286 323 1292 324
rect 1286 319 1287 323
rect 1291 319 1292 323
rect 1286 318 1292 319
rect 1382 323 1388 324
rect 1382 319 1383 323
rect 1387 319 1388 323
rect 1382 318 1388 319
rect 1478 323 1484 324
rect 1478 319 1479 323
rect 1483 319 1484 323
rect 1478 318 1484 319
rect 1574 323 1580 324
rect 1574 319 1575 323
rect 1579 319 1580 323
rect 1574 318 1580 319
rect 1670 323 1676 324
rect 1670 319 1671 323
rect 1675 319 1676 323
rect 1670 318 1676 319
rect 1082 315 1088 316
rect 1082 311 1083 315
rect 1087 311 1088 315
rect 1824 314 1826 329
rect 1864 319 1866 343
rect 1894 335 1900 336
rect 1894 331 1895 335
rect 1899 331 1900 335
rect 1894 330 1900 331
rect 1896 319 1898 330
rect 1863 318 1867 319
rect 1082 310 1088 311
rect 1822 313 1828 314
rect 1863 313 1867 314
rect 1895 318 1899 319
rect 1895 313 1899 314
rect 1822 309 1823 313
rect 1827 309 1828 313
rect 1822 308 1828 309
rect 1082 299 1088 300
rect 1082 295 1083 299
rect 1087 295 1088 299
rect 1082 294 1088 295
rect 1170 299 1176 300
rect 1170 295 1171 299
rect 1175 295 1176 299
rect 1170 294 1176 295
rect 1562 299 1568 300
rect 1562 295 1563 299
rect 1567 295 1568 299
rect 1562 294 1568 295
rect 1642 299 1648 300
rect 1642 295 1643 299
rect 1647 295 1648 299
rect 1642 294 1648 295
rect 1822 296 1828 297
rect 934 283 940 284
rect 934 279 935 283
rect 939 279 940 283
rect 934 278 940 279
rect 1022 283 1028 284
rect 1022 279 1023 283
rect 1027 279 1028 283
rect 1022 278 1028 279
rect 854 271 860 272
rect 854 267 855 271
rect 859 267 860 271
rect 854 266 860 267
rect 936 263 938 278
rect 1024 263 1026 278
rect 1084 264 1086 294
rect 1110 283 1116 284
rect 1110 279 1111 283
rect 1115 279 1116 283
rect 1110 278 1116 279
rect 1082 263 1088 264
rect 1112 263 1114 278
rect 1172 272 1174 294
rect 1198 283 1204 284
rect 1198 279 1199 283
rect 1203 279 1204 283
rect 1198 278 1204 279
rect 1294 283 1300 284
rect 1294 279 1295 283
rect 1299 279 1300 283
rect 1294 278 1300 279
rect 1390 283 1396 284
rect 1390 279 1391 283
rect 1395 279 1396 283
rect 1390 278 1396 279
rect 1486 283 1492 284
rect 1486 279 1487 283
rect 1491 279 1492 283
rect 1486 278 1492 279
rect 1170 271 1176 272
rect 1170 267 1171 271
rect 1175 267 1176 271
rect 1170 266 1176 267
rect 1190 271 1196 272
rect 1190 267 1191 271
rect 1195 267 1196 271
rect 1190 266 1196 267
rect 738 259 739 263
rect 743 259 744 263
rect 738 258 744 259
rect 759 262 763 263
rect 671 257 675 258
rect 144 246 146 257
rect 210 255 216 256
rect 210 251 211 255
rect 215 251 216 255
rect 210 250 216 251
rect 142 245 148 246
rect 142 241 143 245
rect 147 241 148 245
rect 142 240 148 241
rect 212 228 214 250
rect 232 246 234 257
rect 298 255 304 256
rect 298 251 299 255
rect 303 251 304 255
rect 298 250 304 251
rect 230 245 236 246
rect 230 241 231 245
rect 235 241 236 245
rect 230 240 236 241
rect 300 228 302 250
rect 320 246 322 257
rect 386 255 392 256
rect 386 251 387 255
rect 391 251 392 255
rect 386 250 392 251
rect 318 245 324 246
rect 318 241 319 245
rect 323 241 324 245
rect 318 240 324 241
rect 388 228 390 250
rect 408 246 410 257
rect 474 255 480 256
rect 474 251 475 255
rect 479 251 480 255
rect 474 250 480 251
rect 406 245 412 246
rect 406 241 407 245
rect 411 241 412 245
rect 406 240 412 241
rect 476 228 478 250
rect 496 246 498 257
rect 562 255 568 256
rect 562 251 563 255
rect 567 251 568 255
rect 562 250 568 251
rect 494 245 500 246
rect 494 241 495 245
rect 499 241 500 245
rect 494 240 500 241
rect 564 228 566 250
rect 584 246 586 257
rect 650 255 656 256
rect 650 251 651 255
rect 655 251 656 255
rect 650 250 656 251
rect 582 245 588 246
rect 582 241 583 245
rect 587 241 588 245
rect 582 240 588 241
rect 652 228 654 250
rect 672 246 674 257
rect 740 256 742 258
rect 759 257 763 258
rect 847 262 851 263
rect 847 257 851 258
rect 935 262 939 263
rect 935 257 939 258
rect 1023 262 1027 263
rect 1082 259 1083 263
rect 1087 259 1088 263
rect 1082 258 1088 259
rect 1111 262 1115 263
rect 1023 257 1027 258
rect 1111 257 1115 258
rect 734 255 742 256
rect 734 251 735 255
rect 739 251 742 255
rect 734 250 742 251
rect 736 249 742 250
rect 760 246 762 257
rect 848 246 850 257
rect 936 246 938 257
rect 1024 246 1026 257
rect 1030 255 1036 256
rect 1030 250 1031 255
rect 1035 250 1036 255
rect 1031 247 1035 248
rect 1112 246 1114 257
rect 670 245 676 246
rect 670 241 671 245
rect 675 241 676 245
rect 670 240 676 241
rect 758 245 764 246
rect 758 241 759 245
rect 763 241 764 245
rect 758 240 764 241
rect 846 245 852 246
rect 846 241 847 245
rect 851 241 852 245
rect 846 240 852 241
rect 934 245 940 246
rect 934 241 935 245
rect 939 241 940 245
rect 934 240 940 241
rect 1022 245 1028 246
rect 1022 241 1023 245
rect 1027 241 1028 245
rect 1022 240 1028 241
rect 1110 245 1116 246
rect 1110 241 1111 245
rect 1115 241 1116 245
rect 1110 240 1116 241
rect 1192 228 1194 266
rect 1200 263 1202 278
rect 1296 263 1298 278
rect 1303 276 1307 277
rect 1302 271 1308 272
rect 1302 267 1303 271
rect 1307 267 1308 271
rect 1302 266 1308 267
rect 1392 263 1394 278
rect 1488 263 1490 278
rect 1564 277 1566 294
rect 1582 283 1588 284
rect 1582 279 1583 283
rect 1587 279 1588 283
rect 1582 278 1588 279
rect 1563 276 1567 277
rect 1563 271 1567 272
rect 1584 263 1586 278
rect 1644 272 1646 294
rect 1822 292 1823 296
rect 1827 292 1828 296
rect 1822 291 1828 292
rect 1678 283 1684 284
rect 1678 279 1679 283
rect 1683 279 1684 283
rect 1678 278 1684 279
rect 1642 271 1648 272
rect 1642 267 1643 271
rect 1647 267 1648 271
rect 1642 266 1648 267
rect 1680 263 1682 278
rect 1824 263 1826 291
rect 1864 289 1866 313
rect 1896 302 1898 313
rect 1904 312 1906 378
rect 1976 376 1978 381
rect 2064 376 2066 381
rect 2152 376 2154 381
rect 1974 375 1980 376
rect 1974 371 1975 375
rect 1979 371 1980 375
rect 1974 370 1980 371
rect 2062 375 2068 376
rect 2062 371 2063 375
rect 2067 371 2068 375
rect 2062 370 2068 371
rect 2150 375 2156 376
rect 2150 371 2151 375
rect 2155 371 2156 375
rect 2150 370 2156 371
rect 2220 368 2222 442
rect 2384 438 2386 449
rect 2392 448 2394 487
rect 2494 479 2500 480
rect 2494 475 2495 479
rect 2499 475 2500 479
rect 2494 474 2500 475
rect 2638 479 2644 480
rect 2638 475 2639 479
rect 2643 475 2644 479
rect 2638 474 2644 475
rect 2814 479 2820 480
rect 2814 475 2815 479
rect 2819 475 2820 479
rect 2814 474 2820 475
rect 3014 479 3020 480
rect 3014 475 3015 479
rect 3019 475 3020 479
rect 3014 474 3020 475
rect 3222 479 3228 480
rect 3222 475 3223 479
rect 3227 475 3228 479
rect 3222 474 3228 475
rect 3438 479 3444 480
rect 3438 475 3439 479
rect 3443 475 3444 479
rect 3438 474 3444 475
rect 2496 455 2498 474
rect 2640 455 2642 474
rect 2816 455 2818 474
rect 3016 455 3018 474
rect 3224 455 3226 474
rect 3440 455 3442 474
rect 2495 454 2499 455
rect 2495 449 2499 450
rect 2575 454 2579 455
rect 2575 449 2579 450
rect 2639 454 2643 455
rect 2639 449 2643 450
rect 2783 454 2787 455
rect 2783 449 2787 450
rect 2815 454 2819 455
rect 2815 449 2819 450
rect 3007 454 3011 455
rect 3007 449 3011 450
rect 3015 454 3019 455
rect 3015 449 3019 450
rect 3223 454 3227 455
rect 3223 449 3227 450
rect 3239 454 3243 455
rect 3239 449 3243 450
rect 3439 454 3443 455
rect 3439 449 3443 450
rect 3471 454 3475 455
rect 3471 449 3475 450
rect 2390 447 2396 448
rect 2390 443 2391 447
rect 2395 443 2396 447
rect 2390 442 2396 443
rect 2576 438 2578 449
rect 2784 438 2786 449
rect 3008 438 3010 449
rect 3240 438 3242 449
rect 3472 438 3474 449
rect 3500 448 3502 490
rect 3574 488 3575 492
rect 3579 488 3580 492
rect 3574 487 3580 488
rect 3576 455 3578 487
rect 3575 454 3579 455
rect 3575 449 3579 450
rect 3498 447 3504 448
rect 3498 443 3499 447
rect 3503 443 3504 447
rect 3498 442 3504 443
rect 2382 437 2388 438
rect 2382 433 2383 437
rect 2387 433 2388 437
rect 2382 432 2388 433
rect 2574 437 2580 438
rect 2574 433 2575 437
rect 2579 433 2580 437
rect 2574 432 2580 433
rect 2782 437 2788 438
rect 2782 433 2783 437
rect 2787 433 2788 437
rect 2782 432 2788 433
rect 3006 437 3012 438
rect 3006 433 3007 437
rect 3011 433 3012 437
rect 3006 432 3012 433
rect 3238 437 3244 438
rect 3238 433 3239 437
rect 3243 433 3244 437
rect 3238 432 3244 433
rect 3470 437 3476 438
rect 3470 433 3471 437
rect 3475 433 3476 437
rect 3470 432 3476 433
rect 3576 425 3578 449
rect 3574 424 3580 425
rect 3574 420 3575 424
rect 3579 420 3580 424
rect 3574 419 3580 420
rect 3178 407 3184 408
rect 3178 403 3179 407
rect 3183 403 3184 407
rect 3178 402 3184 403
rect 3470 407 3476 408
rect 3470 403 3471 407
rect 3475 403 3476 407
rect 3470 402 3476 403
rect 3574 407 3580 408
rect 3574 403 3575 407
rect 3579 403 3580 407
rect 3574 402 3580 403
rect 2374 397 2380 398
rect 2374 393 2375 397
rect 2379 393 2380 397
rect 2374 392 2380 393
rect 2566 397 2572 398
rect 2566 393 2567 397
rect 2571 393 2572 397
rect 2566 392 2572 393
rect 2774 397 2780 398
rect 2774 393 2775 397
rect 2779 393 2780 397
rect 2774 392 2780 393
rect 2998 397 3004 398
rect 2998 393 2999 397
rect 3003 393 3004 397
rect 2998 392 3004 393
rect 2376 387 2378 392
rect 2568 387 2570 392
rect 2776 387 2778 392
rect 3000 387 3002 392
rect 2263 386 2267 387
rect 2263 381 2267 382
rect 2375 386 2379 387
rect 2375 381 2379 382
rect 2383 386 2387 387
rect 2383 381 2387 382
rect 2519 386 2523 387
rect 2519 381 2523 382
rect 2567 386 2571 387
rect 2567 381 2571 382
rect 2671 386 2675 387
rect 2671 381 2675 382
rect 2775 386 2779 387
rect 2775 381 2779 382
rect 2847 386 2851 387
rect 2847 381 2851 382
rect 2999 386 3003 387
rect 2999 381 3003 382
rect 3031 386 3035 387
rect 3031 381 3035 382
rect 2264 376 2266 381
rect 2384 376 2386 381
rect 2520 376 2522 381
rect 2672 376 2674 381
rect 2848 376 2850 381
rect 3032 376 3034 381
rect 2262 375 2268 376
rect 2262 371 2263 375
rect 2267 371 2268 375
rect 2262 370 2268 371
rect 2382 375 2388 376
rect 2382 371 2383 375
rect 2387 371 2388 375
rect 2382 370 2388 371
rect 2518 375 2524 376
rect 2518 371 2519 375
rect 2523 371 2524 375
rect 2518 370 2524 371
rect 2670 375 2676 376
rect 2670 371 2671 375
rect 2675 371 2676 375
rect 2670 370 2676 371
rect 2846 375 2852 376
rect 2846 371 2847 375
rect 2851 371 2852 375
rect 2846 370 2852 371
rect 3030 375 3036 376
rect 3030 371 3031 375
rect 3035 371 3036 375
rect 3030 370 3036 371
rect 2218 367 2224 368
rect 2218 363 2219 367
rect 2223 363 2224 367
rect 2218 362 2224 363
rect 2450 351 2456 352
rect 2450 347 2451 351
rect 2455 347 2456 351
rect 3150 351 3156 352
rect 2450 346 2456 347
rect 2703 348 2707 349
rect 1982 335 1988 336
rect 1982 331 1983 335
rect 1987 331 1988 335
rect 1982 330 1988 331
rect 2070 335 2076 336
rect 2070 331 2071 335
rect 2075 331 2076 335
rect 2070 330 2076 331
rect 2158 335 2164 336
rect 2158 331 2159 335
rect 2163 331 2164 335
rect 2158 330 2164 331
rect 2270 335 2276 336
rect 2270 331 2271 335
rect 2275 331 2276 335
rect 2270 330 2276 331
rect 2390 335 2396 336
rect 2390 331 2391 335
rect 2395 331 2396 335
rect 2390 330 2396 331
rect 1984 319 1986 330
rect 2072 319 2074 330
rect 2160 319 2162 330
rect 2272 319 2274 330
rect 2392 319 2394 330
rect 2452 324 2454 346
rect 3150 347 3151 351
rect 3155 347 3156 351
rect 3150 346 3156 347
rect 3158 351 3164 352
rect 3158 346 3159 351
rect 2703 343 2707 344
rect 2526 335 2532 336
rect 2526 331 2527 335
rect 2531 331 2532 335
rect 2526 330 2532 331
rect 2678 335 2684 336
rect 2678 331 2679 335
rect 2683 331 2684 335
rect 2678 330 2684 331
rect 2687 332 2691 333
rect 2450 323 2456 324
rect 2450 319 2451 323
rect 2455 319 2456 323
rect 2528 319 2530 330
rect 2534 323 2540 324
rect 2534 319 2535 323
rect 2539 319 2540 323
rect 2680 319 2682 330
rect 2687 327 2691 328
rect 2688 324 2690 327
rect 2686 323 2692 324
rect 2686 319 2687 323
rect 2691 319 2692 323
rect 1983 318 1987 319
rect 1983 313 1987 314
rect 2071 318 2075 319
rect 2071 313 2075 314
rect 2159 318 2163 319
rect 2159 313 2163 314
rect 2247 318 2251 319
rect 2247 313 2251 314
rect 2271 318 2275 319
rect 2271 313 2275 314
rect 2359 318 2363 319
rect 2359 313 2363 314
rect 2391 318 2395 319
rect 2450 318 2456 319
rect 2471 318 2475 319
rect 2391 313 2395 314
rect 2471 313 2475 314
rect 2527 318 2531 319
rect 2534 318 2540 319
rect 2583 318 2587 319
rect 2527 313 2531 314
rect 1902 311 1908 312
rect 1902 307 1903 311
rect 1907 307 1908 311
rect 1902 306 1908 307
rect 1984 302 1986 313
rect 2072 302 2074 313
rect 2160 302 2162 313
rect 2248 302 2250 313
rect 2360 302 2362 313
rect 2366 311 2372 312
rect 2366 306 2367 311
rect 2371 306 2372 311
rect 2367 303 2371 304
rect 2472 302 2474 313
rect 1894 301 1900 302
rect 1894 297 1895 301
rect 1899 297 1900 301
rect 1894 296 1900 297
rect 1982 301 1988 302
rect 1982 297 1983 301
rect 1987 297 1988 301
rect 1982 296 1988 297
rect 2070 301 2076 302
rect 2070 297 2071 301
rect 2075 297 2076 301
rect 2070 296 2076 297
rect 2158 301 2164 302
rect 2158 297 2159 301
rect 2163 297 2164 301
rect 2158 296 2164 297
rect 2246 301 2252 302
rect 2246 297 2247 301
rect 2251 297 2252 301
rect 2246 296 2252 297
rect 2358 301 2364 302
rect 2358 297 2359 301
rect 2363 297 2364 301
rect 2358 296 2364 297
rect 2470 301 2476 302
rect 2470 297 2471 301
rect 2475 297 2476 301
rect 2470 296 2476 297
rect 1862 288 1868 289
rect 2536 288 2538 318
rect 2583 313 2587 314
rect 2679 318 2683 319
rect 2686 318 2692 319
rect 2695 318 2699 319
rect 2679 313 2683 314
rect 2695 313 2699 314
rect 2543 308 2547 309
rect 2543 303 2547 304
rect 1862 284 1863 288
rect 1867 284 1868 288
rect 1862 283 1868 284
rect 2534 287 2540 288
rect 2534 283 2535 287
rect 2539 283 2540 287
rect 2544 284 2546 303
rect 2584 302 2586 313
rect 2602 311 2608 312
rect 2602 307 2603 311
rect 2607 307 2608 311
rect 2602 306 2608 307
rect 2582 301 2588 302
rect 2582 297 2583 301
rect 2587 297 2588 301
rect 2582 296 2588 297
rect 2534 282 2540 283
rect 2542 283 2548 284
rect 2542 279 2543 283
rect 2547 279 2548 283
rect 2542 278 2548 279
rect 1862 271 1868 272
rect 1862 267 1863 271
rect 1867 267 1868 271
rect 1862 266 1868 267
rect 2226 271 2232 272
rect 2226 267 2227 271
rect 2231 267 2232 271
rect 2226 266 2232 267
rect 1199 262 1203 263
rect 1199 257 1203 258
rect 1287 262 1291 263
rect 1287 257 1291 258
rect 1295 262 1299 263
rect 1295 257 1299 258
rect 1375 262 1379 263
rect 1375 257 1379 258
rect 1391 262 1395 263
rect 1391 257 1395 258
rect 1463 262 1467 263
rect 1463 257 1467 258
rect 1487 262 1491 263
rect 1487 257 1491 258
rect 1551 262 1555 263
rect 1551 257 1555 258
rect 1583 262 1587 263
rect 1583 257 1587 258
rect 1639 262 1643 263
rect 1639 257 1643 258
rect 1679 262 1683 263
rect 1679 257 1683 258
rect 1727 262 1731 263
rect 1727 257 1731 258
rect 1823 262 1827 263
rect 1823 257 1827 258
rect 1200 246 1202 257
rect 1267 252 1271 253
rect 1267 247 1271 248
rect 1198 245 1204 246
rect 1198 241 1199 245
rect 1203 241 1204 245
rect 1198 240 1204 241
rect 1268 228 1270 247
rect 1288 246 1290 257
rect 1354 255 1360 256
rect 1354 251 1355 255
rect 1359 251 1360 255
rect 1354 250 1360 251
rect 1286 245 1292 246
rect 1286 241 1287 245
rect 1291 241 1292 245
rect 1286 240 1292 241
rect 1356 228 1358 250
rect 1376 246 1378 257
rect 1442 255 1448 256
rect 1442 251 1443 255
rect 1447 251 1448 255
rect 1442 250 1448 251
rect 1374 245 1380 246
rect 1374 241 1375 245
rect 1379 241 1380 245
rect 1374 240 1380 241
rect 1444 228 1446 250
rect 1464 246 1466 257
rect 1534 255 1540 256
rect 1534 251 1535 255
rect 1539 251 1540 255
rect 1534 250 1540 251
rect 1462 245 1468 246
rect 1462 241 1463 245
rect 1467 241 1468 245
rect 1462 240 1468 241
rect 110 227 116 228
rect 134 227 140 228
rect 134 223 135 227
rect 139 223 140 227
rect 134 222 140 223
rect 210 227 216 228
rect 210 223 211 227
rect 215 223 216 227
rect 210 222 216 223
rect 298 227 304 228
rect 298 223 299 227
rect 303 223 304 227
rect 298 222 304 223
rect 386 227 392 228
rect 386 223 387 227
rect 391 223 392 227
rect 386 222 392 223
rect 474 227 480 228
rect 474 223 475 227
rect 479 223 480 227
rect 474 222 480 223
rect 562 227 568 228
rect 562 223 563 227
rect 567 223 568 227
rect 562 222 568 223
rect 650 227 656 228
rect 650 223 651 227
rect 655 223 656 227
rect 650 222 656 223
rect 1190 227 1196 228
rect 1190 223 1191 227
rect 1195 223 1196 227
rect 1190 222 1196 223
rect 1266 227 1272 228
rect 1266 223 1267 227
rect 1271 223 1272 227
rect 1266 222 1272 223
rect 1354 227 1360 228
rect 1354 223 1355 227
rect 1359 223 1360 227
rect 1354 222 1360 223
rect 1442 227 1448 228
rect 1442 223 1443 227
rect 1447 223 1448 227
rect 1442 222 1448 223
rect 110 215 116 216
rect 110 211 111 215
rect 115 211 116 215
rect 110 210 116 211
rect 112 195 114 210
rect 134 205 140 206
rect 134 201 135 205
rect 139 201 140 205
rect 134 200 140 201
rect 222 205 228 206
rect 222 201 223 205
rect 227 201 228 205
rect 222 200 228 201
rect 310 205 316 206
rect 310 201 311 205
rect 315 201 316 205
rect 310 200 316 201
rect 398 205 404 206
rect 398 201 399 205
rect 403 201 404 205
rect 398 200 404 201
rect 486 205 492 206
rect 486 201 487 205
rect 491 201 492 205
rect 486 200 492 201
rect 574 205 580 206
rect 574 201 575 205
rect 579 201 580 205
rect 574 200 580 201
rect 662 205 668 206
rect 662 201 663 205
rect 667 201 668 205
rect 662 200 668 201
rect 750 205 756 206
rect 750 201 751 205
rect 755 201 756 205
rect 750 200 756 201
rect 838 205 844 206
rect 838 201 839 205
rect 843 201 844 205
rect 838 200 844 201
rect 926 205 932 206
rect 926 201 927 205
rect 931 201 932 205
rect 926 200 932 201
rect 1014 205 1020 206
rect 1014 201 1015 205
rect 1019 201 1020 205
rect 1014 200 1020 201
rect 1102 205 1108 206
rect 1102 201 1103 205
rect 1107 201 1108 205
rect 1102 200 1108 201
rect 1190 205 1196 206
rect 1190 201 1191 205
rect 1195 201 1196 205
rect 1190 200 1196 201
rect 1278 205 1284 206
rect 1278 201 1279 205
rect 1283 201 1284 205
rect 1278 200 1284 201
rect 1366 205 1372 206
rect 1366 201 1367 205
rect 1371 201 1372 205
rect 1366 200 1372 201
rect 1454 205 1460 206
rect 1454 201 1455 205
rect 1459 201 1460 205
rect 1454 200 1460 201
rect 1536 200 1538 250
rect 1552 246 1554 257
rect 1640 246 1642 257
rect 1706 255 1712 256
rect 1706 251 1707 255
rect 1711 251 1712 255
rect 1706 250 1712 251
rect 1550 245 1556 246
rect 1550 241 1551 245
rect 1555 241 1556 245
rect 1550 240 1556 241
rect 1638 245 1644 246
rect 1638 241 1639 245
rect 1643 241 1644 245
rect 1638 240 1644 241
rect 1708 216 1710 250
rect 1728 246 1730 257
rect 1726 245 1732 246
rect 1726 241 1727 245
rect 1731 241 1732 245
rect 1726 240 1732 241
rect 1824 233 1826 257
rect 1864 251 1866 266
rect 1886 261 1892 262
rect 1886 257 1887 261
rect 1891 257 1892 261
rect 1886 256 1892 257
rect 1974 261 1980 262
rect 1974 257 1975 261
rect 1979 257 1980 261
rect 1974 256 1980 257
rect 2062 261 2068 262
rect 2062 257 2063 261
rect 2067 257 2068 261
rect 2062 256 2068 257
rect 2150 261 2156 262
rect 2150 257 2151 261
rect 2155 257 2156 261
rect 2150 256 2156 257
rect 1888 251 1890 256
rect 1976 251 1978 256
rect 2064 251 2066 256
rect 2152 251 2154 256
rect 1863 250 1867 251
rect 1863 245 1867 246
rect 1887 250 1891 251
rect 1887 245 1891 246
rect 1975 250 1979 251
rect 1975 245 1979 246
rect 2063 250 2067 251
rect 2063 245 2067 246
rect 2151 250 2155 251
rect 2151 245 2155 246
rect 1822 232 1828 233
rect 1822 228 1823 232
rect 1827 228 1828 232
rect 1864 230 1866 245
rect 1888 240 1890 245
rect 1976 240 1978 245
rect 2064 240 2066 245
rect 2152 240 2154 245
rect 1886 239 1892 240
rect 1886 235 1887 239
rect 1891 235 1892 239
rect 1886 234 1892 235
rect 1974 239 1980 240
rect 1974 235 1975 239
rect 1979 235 1980 239
rect 1974 234 1980 235
rect 2062 239 2068 240
rect 2062 235 2063 239
rect 2067 235 2068 239
rect 2062 234 2068 235
rect 2150 239 2156 240
rect 2150 235 2151 239
rect 2155 235 2156 239
rect 2150 234 2156 235
rect 1822 227 1828 228
rect 1862 229 1868 230
rect 2228 229 2230 266
rect 2238 261 2244 262
rect 2238 257 2239 261
rect 2243 257 2244 261
rect 2238 256 2244 257
rect 2350 261 2356 262
rect 2350 257 2351 261
rect 2355 257 2356 261
rect 2350 256 2356 257
rect 2462 261 2468 262
rect 2462 257 2463 261
rect 2467 257 2468 261
rect 2462 256 2468 257
rect 2574 261 2580 262
rect 2574 257 2575 261
rect 2579 257 2580 261
rect 2574 256 2580 257
rect 2240 251 2242 256
rect 2352 251 2354 256
rect 2464 251 2466 256
rect 2576 251 2578 256
rect 2239 250 2243 251
rect 2239 245 2243 246
rect 2263 250 2267 251
rect 2263 245 2267 246
rect 2351 250 2355 251
rect 2351 245 2355 246
rect 2399 250 2403 251
rect 2399 245 2403 246
rect 2463 250 2467 251
rect 2463 245 2467 246
rect 2535 250 2539 251
rect 2535 245 2539 246
rect 2575 250 2579 251
rect 2575 245 2579 246
rect 2264 240 2266 245
rect 2400 240 2402 245
rect 2536 240 2538 245
rect 2262 239 2268 240
rect 2262 235 2263 239
rect 2267 235 2268 239
rect 2262 234 2268 235
rect 2398 239 2404 240
rect 2398 235 2399 239
rect 2403 235 2404 239
rect 2398 234 2404 235
rect 2534 239 2540 240
rect 2534 235 2535 239
rect 2539 235 2540 239
rect 2534 234 2540 235
rect 2604 232 2606 306
rect 2696 302 2698 313
rect 2704 312 2706 343
rect 2854 335 2860 336
rect 2854 331 2855 335
rect 2859 331 2860 335
rect 2854 330 2860 331
rect 3038 335 3044 336
rect 3038 331 3039 335
rect 3043 331 3044 335
rect 3038 330 3044 331
rect 2856 319 2858 330
rect 3040 319 3042 330
rect 3152 324 3154 346
rect 3163 346 3164 351
rect 3159 343 3163 344
rect 3180 333 3182 402
rect 3230 397 3236 398
rect 3230 393 3231 397
rect 3235 393 3236 397
rect 3230 392 3236 393
rect 3462 397 3468 398
rect 3462 393 3463 397
rect 3467 393 3468 397
rect 3462 392 3468 393
rect 3232 387 3234 392
rect 3464 387 3466 392
rect 3231 386 3235 387
rect 3231 381 3235 382
rect 3431 386 3435 387
rect 3431 381 3435 382
rect 3463 386 3467 387
rect 3463 381 3467 382
rect 3232 376 3234 381
rect 3432 376 3434 381
rect 3230 375 3236 376
rect 3230 371 3231 375
rect 3235 371 3236 375
rect 3230 370 3236 371
rect 3430 375 3436 376
rect 3430 371 3431 375
rect 3435 371 3436 375
rect 3430 370 3436 371
rect 3238 335 3244 336
rect 3179 332 3183 333
rect 3238 331 3239 335
rect 3243 331 3244 335
rect 3238 330 3244 331
rect 3438 335 3444 336
rect 3438 331 3439 335
rect 3443 331 3444 335
rect 3438 330 3444 331
rect 3179 327 3183 328
rect 3150 323 3156 324
rect 3150 319 3151 323
rect 3155 319 3156 323
rect 3240 319 3242 330
rect 3426 323 3432 324
rect 3426 319 3427 323
rect 3431 319 3432 323
rect 3440 319 3442 330
rect 2807 318 2811 319
rect 2807 313 2811 314
rect 2855 318 2859 319
rect 2855 313 2859 314
rect 2919 318 2923 319
rect 2919 313 2923 314
rect 3039 318 3043 319
rect 3150 318 3156 319
rect 3159 318 3163 319
rect 3039 313 3043 314
rect 3159 313 3163 314
rect 3239 318 3243 319
rect 3426 318 3432 319
rect 3439 318 3443 319
rect 3239 313 3243 314
rect 2702 311 2708 312
rect 2702 307 2703 311
rect 2707 307 2708 311
rect 2702 306 2708 307
rect 2808 302 2810 313
rect 2920 302 2922 313
rect 3040 302 3042 313
rect 3160 302 3162 313
rect 2694 301 2700 302
rect 2694 297 2695 301
rect 2699 297 2700 301
rect 2694 296 2700 297
rect 2806 301 2812 302
rect 2806 297 2807 301
rect 2811 297 2812 301
rect 2806 296 2812 297
rect 2918 301 2924 302
rect 2918 297 2919 301
rect 2923 297 2924 301
rect 2918 296 2924 297
rect 3038 301 3044 302
rect 3038 297 3039 301
rect 3043 297 3044 301
rect 3038 296 3044 297
rect 3158 301 3164 302
rect 3158 297 3159 301
rect 3163 297 3164 301
rect 3158 296 3164 297
rect 3106 271 3112 272
rect 3106 267 3107 271
rect 3111 267 3112 271
rect 3106 266 3112 267
rect 2686 261 2692 262
rect 2686 257 2687 261
rect 2691 257 2692 261
rect 2686 256 2692 257
rect 2798 261 2804 262
rect 2798 257 2799 261
rect 2803 257 2804 261
rect 2798 256 2804 257
rect 2910 261 2916 262
rect 2910 257 2911 261
rect 2915 257 2916 261
rect 2910 256 2916 257
rect 3030 261 3036 262
rect 3030 257 3031 261
rect 3035 257 3036 261
rect 3030 256 3036 257
rect 2688 251 2690 256
rect 2800 251 2802 256
rect 2912 251 2914 256
rect 3032 251 3034 256
rect 2679 250 2683 251
rect 2679 245 2683 246
rect 2687 250 2691 251
rect 2687 245 2691 246
rect 2799 250 2803 251
rect 2799 245 2803 246
rect 2815 250 2819 251
rect 2815 245 2819 246
rect 2911 250 2915 251
rect 2911 245 2915 246
rect 2951 250 2955 251
rect 2951 245 2955 246
rect 3031 250 3035 251
rect 3031 245 3035 246
rect 3087 250 3091 251
rect 3087 245 3091 246
rect 2680 240 2682 245
rect 2816 240 2818 245
rect 2952 240 2954 245
rect 3088 240 3090 245
rect 2678 239 2684 240
rect 2678 235 2679 239
rect 2683 235 2684 239
rect 2678 234 2684 235
rect 2814 239 2820 240
rect 2814 235 2815 239
rect 2819 235 2820 239
rect 2814 234 2820 235
rect 2950 239 2956 240
rect 2950 235 2951 239
rect 2955 235 2956 239
rect 2950 234 2956 235
rect 3086 239 3092 240
rect 3086 235 3087 239
rect 3091 235 3092 239
rect 3086 234 3092 235
rect 2602 231 2608 232
rect 1862 225 1863 229
rect 1867 225 1868 229
rect 1862 224 1868 225
rect 1903 228 1907 229
rect 1903 223 1907 224
rect 2227 228 2231 229
rect 2602 227 2603 231
rect 2607 227 2608 231
rect 2602 226 2608 227
rect 2227 223 2231 224
rect 1706 215 1712 216
rect 1706 211 1707 215
rect 1711 211 1712 215
rect 1706 210 1712 211
rect 1726 215 1732 216
rect 1726 211 1727 215
rect 1731 211 1732 215
rect 1726 210 1732 211
rect 1822 215 1828 216
rect 1822 211 1823 215
rect 1827 211 1828 215
rect 1822 210 1828 211
rect 1862 212 1868 213
rect 1542 205 1548 206
rect 1542 201 1543 205
rect 1547 201 1548 205
rect 1542 200 1548 201
rect 1630 205 1636 206
rect 1630 201 1631 205
rect 1635 201 1636 205
rect 1630 200 1636 201
rect 1718 205 1724 206
rect 1718 201 1719 205
rect 1723 201 1724 205
rect 1718 200 1724 201
rect 1728 200 1730 210
rect 136 195 138 200
rect 224 195 226 200
rect 312 195 314 200
rect 400 195 402 200
rect 488 195 490 200
rect 576 195 578 200
rect 664 195 666 200
rect 752 195 754 200
rect 840 195 842 200
rect 928 195 930 200
rect 1016 195 1018 200
rect 1104 195 1106 200
rect 1192 195 1194 200
rect 1280 195 1282 200
rect 1368 195 1370 200
rect 1456 195 1458 200
rect 1534 199 1540 200
rect 1534 195 1535 199
rect 1539 195 1540 199
rect 1544 195 1546 200
rect 1632 195 1634 200
rect 1720 195 1722 200
rect 1726 199 1732 200
rect 1726 195 1727 199
rect 1731 195 1732 199
rect 1824 195 1826 210
rect 1862 208 1863 212
rect 1867 208 1868 212
rect 1862 207 1868 208
rect 111 194 115 195
rect 111 189 115 190
rect 135 194 139 195
rect 135 189 139 190
rect 223 194 227 195
rect 223 189 227 190
rect 311 194 315 195
rect 311 189 315 190
rect 399 194 403 195
rect 399 189 403 190
rect 487 194 491 195
rect 487 189 491 190
rect 575 194 579 195
rect 575 189 579 190
rect 663 194 667 195
rect 663 189 667 190
rect 751 194 755 195
rect 751 189 755 190
rect 839 194 843 195
rect 839 189 843 190
rect 927 194 931 195
rect 927 189 931 190
rect 1015 194 1019 195
rect 1015 189 1019 190
rect 1103 194 1107 195
rect 1103 189 1107 190
rect 1191 194 1195 195
rect 1191 189 1195 190
rect 1279 194 1283 195
rect 1279 189 1283 190
rect 1367 194 1371 195
rect 1367 189 1371 190
rect 1455 194 1459 195
rect 1534 194 1540 195
rect 1543 194 1547 195
rect 1455 189 1459 190
rect 1543 189 1547 190
rect 1631 194 1635 195
rect 1631 189 1635 190
rect 1719 194 1723 195
rect 1726 194 1732 195
rect 1823 194 1827 195
rect 1719 189 1723 190
rect 1823 189 1827 190
rect 1864 151 1866 207
rect 1894 199 1900 200
rect 1894 195 1895 199
rect 1899 195 1900 199
rect 1894 194 1900 195
rect 1896 151 1898 194
rect 1904 188 1906 223
rect 1982 199 1988 200
rect 1982 195 1983 199
rect 1987 195 1988 199
rect 1982 194 1988 195
rect 2070 199 2076 200
rect 2070 195 2071 199
rect 2075 195 2076 199
rect 2070 194 2076 195
rect 2158 199 2164 200
rect 2158 195 2159 199
rect 2163 195 2164 199
rect 2158 194 2164 195
rect 2270 199 2276 200
rect 2270 195 2271 199
rect 2275 195 2276 199
rect 2270 194 2276 195
rect 2406 199 2412 200
rect 2406 195 2407 199
rect 2411 195 2412 199
rect 2406 194 2412 195
rect 2542 199 2548 200
rect 2542 195 2543 199
rect 2547 195 2548 199
rect 2542 194 2548 195
rect 2686 199 2692 200
rect 2686 195 2687 199
rect 2691 195 2692 199
rect 2686 194 2692 195
rect 2822 199 2828 200
rect 2822 195 2823 199
rect 2827 195 2828 199
rect 2958 199 2964 200
rect 2822 194 2828 195
rect 2831 196 2835 197
rect 1902 187 1908 188
rect 1902 183 1903 187
rect 1907 183 1908 187
rect 1902 182 1908 183
rect 1984 151 1986 194
rect 2072 151 2074 194
rect 2160 151 2162 194
rect 2272 151 2274 194
rect 2408 151 2410 194
rect 2544 151 2546 194
rect 2688 151 2690 194
rect 2791 180 2795 181
rect 2791 175 2795 176
rect 1863 150 1867 151
rect 1863 145 1867 146
rect 1895 150 1899 151
rect 1895 145 1899 146
rect 1983 150 1987 151
rect 1983 145 1987 146
rect 2071 150 2075 151
rect 2071 145 2075 146
rect 2159 150 2163 151
rect 2159 145 2163 146
rect 2271 150 2275 151
rect 2271 145 2275 146
rect 2407 150 2411 151
rect 2407 145 2411 146
rect 2543 150 2547 151
rect 2543 145 2547 146
rect 2687 150 2691 151
rect 2687 145 2691 146
rect 2783 150 2787 151
rect 2783 145 2787 146
rect 1864 121 1866 145
rect 2784 134 2786 145
rect 2792 144 2794 175
rect 2824 151 2826 194
rect 2958 195 2959 199
rect 2963 195 2964 199
rect 2958 194 2964 195
rect 3094 199 3100 200
rect 3094 195 3095 199
rect 3099 195 3100 199
rect 3108 197 3110 266
rect 3150 261 3156 262
rect 3150 257 3151 261
rect 3155 257 3156 261
rect 3150 256 3156 257
rect 3152 251 3154 256
rect 3151 250 3155 251
rect 3151 245 3155 246
rect 3223 250 3227 251
rect 3223 245 3227 246
rect 3359 250 3363 251
rect 3359 245 3363 246
rect 3224 240 3226 245
rect 3360 240 3362 245
rect 3222 239 3228 240
rect 3222 235 3223 239
rect 3227 235 3228 239
rect 3222 234 3228 235
rect 3358 239 3364 240
rect 3358 235 3359 239
rect 3363 235 3364 239
rect 3358 234 3364 235
rect 3428 232 3430 318
rect 3439 313 3443 314
rect 3190 231 3196 232
rect 3190 227 3191 231
rect 3195 227 3196 231
rect 3190 226 3196 227
rect 3426 231 3432 232
rect 3426 227 3427 231
rect 3431 227 3432 231
rect 3426 226 3432 227
rect 3094 194 3100 195
rect 3107 196 3111 197
rect 2831 191 2835 192
rect 2832 188 2834 191
rect 2830 187 2836 188
rect 2830 183 2831 187
rect 2835 183 2836 187
rect 2830 182 2836 183
rect 2960 151 2962 194
rect 3096 151 3098 194
rect 3107 191 3111 192
rect 3192 181 3194 226
rect 3230 199 3236 200
rect 3230 195 3231 199
rect 3235 195 3236 199
rect 3230 194 3236 195
rect 3366 199 3372 200
rect 3366 195 3367 199
rect 3371 195 3372 199
rect 3366 194 3372 195
rect 3191 180 3195 181
rect 3191 175 3195 176
rect 3232 151 3234 194
rect 3368 151 3370 194
rect 3472 188 3474 402
rect 3576 387 3578 402
rect 3575 386 3579 387
rect 3575 381 3579 382
rect 3576 366 3578 381
rect 3574 365 3580 366
rect 3574 361 3575 365
rect 3579 361 3580 365
rect 3574 360 3580 361
rect 3574 348 3580 349
rect 3574 344 3575 348
rect 3579 344 3580 348
rect 3574 343 3580 344
rect 3576 319 3578 343
rect 3575 318 3579 319
rect 3575 313 3579 314
rect 3576 289 3578 313
rect 3574 288 3580 289
rect 3574 284 3575 288
rect 3579 284 3580 288
rect 3574 283 3580 284
rect 3574 271 3580 272
rect 3574 267 3575 271
rect 3579 267 3580 271
rect 3574 266 3580 267
rect 3576 251 3578 266
rect 3479 250 3483 251
rect 3479 245 3483 246
rect 3575 250 3579 251
rect 3575 245 3579 246
rect 3480 240 3482 245
rect 3478 239 3484 240
rect 3478 235 3479 239
rect 3483 235 3484 239
rect 3478 234 3484 235
rect 3576 230 3578 245
rect 3574 229 3580 230
rect 3574 225 3575 229
rect 3579 225 3580 229
rect 3574 224 3580 225
rect 3574 212 3580 213
rect 3574 208 3575 212
rect 3579 208 3580 212
rect 3574 207 3580 208
rect 3486 199 3492 200
rect 3486 195 3487 199
rect 3491 195 3492 199
rect 3486 194 3492 195
rect 3374 187 3380 188
rect 3374 183 3375 187
rect 3379 183 3380 187
rect 3374 182 3380 183
rect 3470 187 3476 188
rect 3470 183 3471 187
rect 3475 183 3476 187
rect 3470 182 3476 183
rect 2823 150 2827 151
rect 2823 145 2827 146
rect 2871 150 2875 151
rect 2871 145 2875 146
rect 2959 150 2963 151
rect 2959 145 2963 146
rect 3047 150 3051 151
rect 3047 145 3051 146
rect 3095 150 3099 151
rect 3095 145 3099 146
rect 3135 150 3139 151
rect 3135 145 3139 146
rect 3223 150 3227 151
rect 3223 145 3227 146
rect 3231 150 3235 151
rect 3231 145 3235 146
rect 3311 150 3315 151
rect 3311 145 3315 146
rect 3367 150 3371 151
rect 3367 145 3371 146
rect 2790 143 2796 144
rect 2790 139 2791 143
rect 2795 139 2796 143
rect 2790 138 2796 139
rect 2872 134 2874 145
rect 2960 134 2962 145
rect 3048 134 3050 145
rect 3136 134 3138 145
rect 3224 134 3226 145
rect 3312 134 3314 145
rect 2782 133 2788 134
rect 2782 129 2783 133
rect 2787 129 2788 133
rect 2782 128 2788 129
rect 2870 133 2876 134
rect 2870 129 2871 133
rect 2875 129 2876 133
rect 2870 128 2876 129
rect 2958 133 2964 134
rect 2958 129 2959 133
rect 2963 129 2964 133
rect 2958 128 2964 129
rect 3046 133 3052 134
rect 3046 129 3047 133
rect 3051 129 3052 133
rect 3046 128 3052 129
rect 3134 133 3140 134
rect 3134 129 3135 133
rect 3139 129 3140 133
rect 3134 128 3140 129
rect 3222 133 3228 134
rect 3222 129 3223 133
rect 3227 129 3228 133
rect 3222 128 3228 129
rect 3310 133 3316 134
rect 3310 129 3311 133
rect 3315 129 3316 133
rect 3310 128 3316 129
rect 1862 120 1868 121
rect 3376 120 3378 182
rect 3488 151 3490 194
rect 3576 151 3578 207
rect 3399 150 3403 151
rect 3399 145 3403 146
rect 3487 150 3491 151
rect 3487 145 3491 146
rect 3575 150 3579 151
rect 3575 145 3579 146
rect 3400 134 3402 145
rect 3458 143 3464 144
rect 3458 139 3459 143
rect 3463 139 3464 143
rect 3458 138 3464 139
rect 3398 133 3404 134
rect 3398 129 3399 133
rect 3403 129 3404 133
rect 3398 128 3404 129
rect 3460 120 3462 138
rect 3488 134 3490 145
rect 3486 133 3492 134
rect 3486 129 3487 133
rect 3491 129 3492 133
rect 3486 128 3492 129
rect 3576 121 3578 145
rect 3574 120 3580 121
rect 1862 116 1863 120
rect 1867 116 1868 120
rect 1862 115 1868 116
rect 3374 119 3380 120
rect 3374 115 3375 119
rect 3379 115 3380 119
rect 3374 114 3380 115
rect 3458 119 3464 120
rect 3458 115 3459 119
rect 3463 115 3464 119
rect 3574 116 3575 120
rect 3579 116 3580 120
rect 3574 115 3580 116
rect 3458 114 3464 115
rect 1862 103 1868 104
rect 1862 99 1863 103
rect 1867 99 1868 103
rect 1862 98 1868 99
rect 3574 103 3580 104
rect 3574 99 3575 103
rect 3579 99 3580 103
rect 3574 98 3580 99
rect 1864 83 1866 98
rect 2774 93 2780 94
rect 2774 89 2775 93
rect 2779 89 2780 93
rect 2774 88 2780 89
rect 2862 93 2868 94
rect 2862 89 2863 93
rect 2867 89 2868 93
rect 2862 88 2868 89
rect 2950 93 2956 94
rect 2950 89 2951 93
rect 2955 89 2956 93
rect 2950 88 2956 89
rect 3038 93 3044 94
rect 3038 89 3039 93
rect 3043 89 3044 93
rect 3038 88 3044 89
rect 3126 93 3132 94
rect 3126 89 3127 93
rect 3131 89 3132 93
rect 3126 88 3132 89
rect 3214 93 3220 94
rect 3214 89 3215 93
rect 3219 89 3220 93
rect 3214 88 3220 89
rect 3302 93 3308 94
rect 3302 89 3303 93
rect 3307 89 3308 93
rect 3302 88 3308 89
rect 3390 93 3396 94
rect 3390 89 3391 93
rect 3395 89 3396 93
rect 3390 88 3396 89
rect 3478 93 3484 94
rect 3478 89 3479 93
rect 3483 89 3484 93
rect 3478 88 3484 89
rect 2776 83 2778 88
rect 2864 83 2866 88
rect 2952 83 2954 88
rect 3040 83 3042 88
rect 3128 83 3130 88
rect 3216 83 3218 88
rect 3304 83 3306 88
rect 3392 83 3394 88
rect 3480 83 3482 88
rect 3576 83 3578 98
rect 1863 82 1867 83
rect 1863 77 1867 78
rect 2775 82 2779 83
rect 2775 77 2779 78
rect 2863 82 2867 83
rect 2863 77 2867 78
rect 2951 82 2955 83
rect 2951 77 2955 78
rect 3039 82 3043 83
rect 3039 77 3043 78
rect 3127 82 3131 83
rect 3127 77 3131 78
rect 3215 82 3219 83
rect 3215 77 3219 78
rect 3303 82 3307 83
rect 3303 77 3307 78
rect 3391 82 3395 83
rect 3391 77 3395 78
rect 3479 82 3483 83
rect 3479 77 3483 78
rect 3575 82 3579 83
rect 3575 77 3579 78
<< m4c >>
rect 111 3666 115 3670
rect 135 3666 139 3670
rect 223 3666 227 3670
rect 1823 3666 1827 3670
rect 111 3598 115 3602
rect 143 3598 147 3602
rect 231 3598 235 3602
rect 319 3598 323 3602
rect 407 3598 411 3602
rect 495 3598 499 3602
rect 1823 3598 1827 3602
rect 1863 3590 1867 3594
rect 1887 3590 1891 3594
rect 1975 3590 1979 3594
rect 2063 3590 2067 3594
rect 2151 3590 2155 3594
rect 2239 3590 2243 3594
rect 2327 3590 2331 3594
rect 2431 3590 2435 3594
rect 2535 3590 2539 3594
rect 2631 3590 2635 3594
rect 2727 3590 2731 3594
rect 2823 3590 2827 3594
rect 2919 3590 2923 3594
rect 3015 3590 3019 3594
rect 3119 3590 3123 3594
rect 3223 3590 3227 3594
rect 3575 3590 3579 3594
rect 2111 3552 2115 3556
rect 2499 3552 2503 3556
rect 111 3530 115 3534
rect 135 3530 139 3534
rect 223 3530 227 3534
rect 247 3530 251 3534
rect 311 3530 315 3534
rect 375 3530 379 3534
rect 399 3530 403 3534
rect 487 3530 491 3534
rect 503 3530 507 3534
rect 623 3530 627 3534
rect 743 3530 747 3534
rect 863 3530 867 3534
rect 975 3530 979 3534
rect 1079 3530 1083 3534
rect 1175 3530 1179 3534
rect 1271 3530 1275 3534
rect 1367 3530 1371 3534
rect 1471 3530 1475 3534
rect 1575 3530 1579 3534
rect 1823 3530 1827 3534
rect 1863 3522 1867 3526
rect 111 3462 115 3466
rect 175 3462 179 3466
rect 255 3462 259 3466
rect 303 3462 307 3466
rect 383 3462 387 3466
rect 447 3462 451 3466
rect 511 3462 515 3466
rect 591 3462 595 3466
rect 631 3462 635 3466
rect 743 3462 747 3466
rect 751 3462 755 3466
rect 871 3462 875 3466
rect 895 3462 899 3466
rect 983 3462 987 3466
rect 1039 3462 1043 3466
rect 1087 3462 1091 3466
rect 1183 3462 1187 3466
rect 1279 3462 1283 3466
rect 1327 3462 1331 3466
rect 1375 3462 1379 3466
rect 1479 3462 1483 3466
rect 1895 3522 1899 3526
rect 1983 3522 1987 3526
rect 2071 3522 2075 3526
rect 2103 3522 2107 3526
rect 1583 3462 1587 3466
rect 1823 3462 1827 3466
rect 1863 3446 1867 3450
rect 1887 3446 1891 3450
rect 1975 3446 1979 3450
rect 1439 3432 1443 3436
rect 1471 3432 1475 3436
rect 2159 3522 2163 3526
rect 2231 3522 2235 3526
rect 2247 3522 2251 3526
rect 2335 3522 2339 3526
rect 2367 3522 2371 3526
rect 2439 3522 2443 3526
rect 2511 3522 2515 3526
rect 2543 3522 2547 3526
rect 2639 3522 2643 3526
rect 2655 3522 2659 3526
rect 2735 3522 2739 3526
rect 2791 3522 2795 3526
rect 2831 3522 2835 3526
rect 2927 3522 2931 3526
rect 2935 3522 2939 3526
rect 3023 3522 3027 3526
rect 3079 3522 3083 3526
rect 3127 3522 3131 3526
rect 2023 3446 2027 3450
rect 2095 3446 2099 3450
rect 2191 3446 2195 3450
rect 2223 3446 2227 3450
rect 2359 3446 2363 3450
rect 2367 3446 2371 3450
rect 2503 3446 2507 3450
rect 2543 3446 2547 3450
rect 2647 3446 2651 3450
rect 2711 3446 2715 3450
rect 2783 3446 2787 3450
rect 3223 3522 3227 3526
rect 3231 3522 3235 3526
rect 3575 3522 3579 3526
rect 2871 3446 2875 3450
rect 111 3394 115 3398
rect 135 3394 139 3398
rect 167 3394 171 3398
rect 263 3394 267 3398
rect 295 3394 299 3398
rect 407 3394 411 3398
rect 439 3394 443 3398
rect 567 3394 571 3398
rect 583 3394 587 3398
rect 727 3394 731 3398
rect 735 3394 739 3398
rect 887 3394 891 3398
rect 1031 3394 1035 3398
rect 1047 3394 1051 3398
rect 1175 3394 1179 3398
rect 1207 3394 1211 3398
rect 215 3336 219 3340
rect 111 3322 115 3326
rect 143 3322 147 3326
rect 207 3322 211 3326
rect 683 3336 687 3340
rect 1319 3394 1323 3398
rect 1367 3394 1371 3398
rect 1471 3394 1475 3398
rect 1527 3394 1531 3398
rect 1823 3394 1827 3398
rect 1863 3370 1867 3374
rect 1895 3370 1899 3374
rect 2031 3370 2035 3374
rect 2199 3370 2203 3374
rect 2375 3370 2379 3374
rect 2551 3370 2555 3374
rect 2927 3446 2931 3450
rect 3031 3446 3035 3450
rect 3071 3446 3075 3450
rect 3191 3446 3195 3450
rect 3215 3446 3219 3450
rect 3359 3446 3363 3450
rect 3575 3446 3579 3450
rect 3047 3392 3051 3396
rect 2719 3370 2723 3374
rect 2879 3370 2883 3374
rect 3039 3370 3043 3374
rect 271 3322 275 3326
rect 335 3322 339 3326
rect 415 3322 419 3326
rect 479 3322 483 3326
rect 575 3322 579 3326
rect 639 3322 643 3326
rect 735 3322 739 3326
rect 807 3322 811 3326
rect 895 3322 899 3326
rect 983 3322 987 3326
rect 1055 3322 1059 3326
rect 1167 3322 1171 3326
rect 1215 3322 1219 3326
rect 1351 3322 1355 3326
rect 1375 3322 1379 3326
rect 1535 3322 1539 3326
rect 1543 3322 1547 3326
rect 1823 3322 1827 3326
rect 111 3250 115 3254
rect 199 3250 203 3254
rect 327 3250 331 3254
rect 367 3250 371 3254
rect 471 3250 475 3254
rect 503 3250 507 3254
rect 631 3250 635 3254
rect 639 3250 643 3254
rect 783 3250 787 3254
rect 799 3250 803 3254
rect 935 3250 939 3254
rect 975 3250 979 3254
rect 1095 3250 1099 3254
rect 1159 3250 1163 3254
rect 1863 3302 1867 3306
rect 1887 3302 1891 3306
rect 2007 3302 2011 3306
rect 2023 3302 2027 3306
rect 2151 3302 2155 3306
rect 2191 3302 2195 3306
rect 2303 3302 2307 3306
rect 2367 3302 2371 3306
rect 2463 3302 2467 3306
rect 2183 3272 2187 3276
rect 1255 3250 1259 3254
rect 1343 3250 1347 3254
rect 1415 3250 1419 3254
rect 1535 3250 1539 3254
rect 1575 3250 1579 3254
rect 1823 3250 1827 3254
rect 487 3192 491 3196
rect 111 3174 115 3178
rect 375 3174 379 3178
rect 447 3174 451 3178
rect 1863 3226 1867 3230
rect 1895 3226 1899 3230
rect 951 3200 955 3204
rect 1163 3200 1167 3204
rect 711 3192 715 3196
rect 511 3174 515 3178
rect 559 3174 563 3178
rect 647 3174 651 3178
rect 687 3174 691 3178
rect 791 3174 795 3178
rect 823 3174 827 3178
rect 943 3174 947 3178
rect 975 3174 979 3178
rect 1103 3174 1107 3178
rect 1135 3174 1139 3178
rect 1263 3174 1267 3178
rect 1295 3174 1299 3178
rect 1423 3174 1427 3178
rect 1463 3174 1467 3178
rect 1583 3174 1587 3178
rect 1639 3174 1643 3178
rect 111 3098 115 3102
rect 439 3098 443 3102
rect 551 3098 555 3102
rect 663 3098 667 3102
rect 679 3098 683 3102
rect 783 3098 787 3102
rect 815 3098 819 3102
rect 903 3098 907 3102
rect 967 3098 971 3102
rect 1031 3098 1035 3102
rect 1127 3098 1131 3102
rect 1159 3098 1163 3102
rect 1287 3098 1291 3102
rect 2167 3248 2171 3252
rect 2015 3226 2019 3230
rect 2023 3226 2027 3230
rect 2159 3226 2163 3230
rect 2175 3226 2179 3230
rect 1823 3174 1827 3178
rect 1863 3154 1867 3158
rect 1887 3154 1891 3158
rect 2015 3154 2019 3158
rect 2543 3302 2547 3306
rect 2631 3302 2635 3306
rect 2711 3302 2715 3306
rect 2799 3302 2803 3306
rect 2871 3302 2875 3306
rect 3259 3392 3263 3396
rect 3191 3370 3195 3374
rect 3199 3370 3203 3374
rect 3343 3370 3347 3374
rect 3367 3370 3371 3374
rect 3487 3370 3491 3374
rect 3575 3370 3579 3374
rect 2967 3302 2971 3306
rect 3031 3302 3035 3306
rect 3135 3302 3139 3306
rect 3183 3302 3187 3306
rect 3311 3302 3315 3306
rect 3335 3302 3339 3306
rect 2539 3272 2543 3276
rect 2479 3248 2483 3252
rect 2311 3226 2315 3230
rect 2327 3226 2331 3230
rect 2463 3226 2467 3230
rect 2471 3226 2475 3230
rect 2599 3226 2603 3230
rect 2639 3226 2643 3230
rect 2735 3226 2739 3230
rect 2807 3226 2811 3230
rect 2871 3226 2875 3230
rect 2975 3226 2979 3230
rect 3015 3226 3019 3230
rect 3143 3226 3147 3230
rect 3167 3226 3171 3230
rect 2047 3154 2051 3158
rect 2167 3154 2171 3158
rect 2199 3154 2203 3158
rect 2319 3154 2323 3158
rect 2351 3154 2355 3158
rect 2455 3154 2459 3158
rect 2511 3154 2515 3158
rect 1423 3098 1427 3102
rect 1455 3098 1459 3102
rect 1559 3098 1563 3102
rect 1631 3098 1635 3102
rect 1695 3098 1699 3102
rect 1823 3098 1827 3102
rect 2215 3096 2219 3100
rect 2591 3154 2595 3158
rect 2679 3154 2683 3158
rect 2727 3154 2731 3158
rect 3479 3302 3483 3306
rect 3575 3302 3579 3306
rect 3319 3226 3323 3230
rect 3327 3226 3331 3230
rect 3487 3226 3491 3230
rect 3575 3226 3579 3230
rect 2863 3154 2867 3158
rect 2871 3154 2875 3158
rect 3007 3154 3011 3158
rect 3071 3154 3075 3158
rect 3159 3154 3163 3158
rect 3287 3154 3291 3158
rect 3319 3154 3323 3158
rect 3479 3154 3483 3158
rect 3575 3154 3579 3158
rect 2531 3096 2535 3100
rect 1863 3078 1867 3082
rect 1895 3078 1899 3082
rect 1919 3078 1923 3082
rect 2055 3078 2059 3082
rect 2087 3078 2091 3082
rect 2207 3078 2211 3082
rect 2279 3078 2283 3082
rect 2359 3078 2363 3082
rect 2487 3078 2491 3082
rect 2519 3078 2523 3082
rect 2687 3078 2691 3082
rect 2719 3078 2723 3082
rect 567 3072 571 3076
rect 891 3072 895 3076
rect 111 3026 115 3030
rect 559 3026 563 3030
rect 575 3026 579 3030
rect 671 3026 675 3030
rect 703 3026 707 3030
rect 791 3026 795 3030
rect 831 3026 835 3030
rect 911 3026 915 3030
rect 967 3026 971 3030
rect 1039 3026 1043 3030
rect 1103 3026 1107 3030
rect 1167 3026 1171 3030
rect 1239 3026 1243 3030
rect 1295 3026 1299 3030
rect 1367 3026 1371 3030
rect 1431 3026 1435 3030
rect 1495 3026 1499 3030
rect 1567 3026 1571 3030
rect 1623 3026 1627 3030
rect 1703 3026 1707 3030
rect 1735 3026 1739 3030
rect 111 2958 115 2962
rect 495 2958 499 2962
rect 567 2958 571 2962
rect 639 2958 643 2962
rect 695 2958 699 2962
rect 783 2958 787 2962
rect 823 2958 827 2962
rect 919 2958 923 2962
rect 959 2958 963 2962
rect 1055 2958 1059 2962
rect 1095 2958 1099 2962
rect 1183 2958 1187 2962
rect 1231 2958 1235 2962
rect 1303 2958 1307 2962
rect 1359 2958 1363 2962
rect 1415 2958 1419 2962
rect 1487 2958 1491 2962
rect 1527 2958 1531 2962
rect 2879 3078 2883 3082
rect 2975 3078 2979 3082
rect 3079 3078 3083 3082
rect 3239 3078 3243 3082
rect 3295 3078 3299 3082
rect 2503 3048 2507 3052
rect 2899 3048 2903 3052
rect 1823 3026 1827 3030
rect 1863 3006 1867 3010
rect 1911 3006 1915 3010
rect 2023 3006 2027 3010
rect 2079 3006 2083 3010
rect 2159 3006 2163 3010
rect 2271 3006 2275 3010
rect 2287 3006 2291 3010
rect 2415 3006 2419 3010
rect 1615 2958 1619 2962
rect 1639 2958 1643 2962
rect 111 2886 115 2890
rect 327 2886 331 2890
rect 455 2886 459 2890
rect 503 2886 507 2890
rect 591 2886 595 2890
rect 647 2886 651 2890
rect 727 2886 731 2890
rect 791 2886 795 2890
rect 871 2886 875 2890
rect 927 2886 931 2890
rect 1007 2886 1011 2890
rect 1063 2886 1067 2890
rect 1143 2886 1147 2890
rect 111 2810 115 2814
rect 167 2810 171 2814
rect 295 2810 299 2814
rect 319 2810 323 2814
rect 423 2810 427 2814
rect 447 2810 451 2814
rect 559 2810 563 2814
rect 583 2810 587 2814
rect 695 2810 699 2814
rect 719 2810 723 2814
rect 823 2810 827 2814
rect 863 2810 867 2814
rect 951 2810 955 2814
rect 999 2810 1003 2814
rect 1727 2958 1731 2962
rect 1823 2958 1827 2962
rect 2479 3006 2483 3010
rect 2535 3006 2539 3010
rect 2663 3006 2667 3010
rect 2711 3006 2715 3010
rect 2807 3006 2811 3010
rect 2967 3006 2971 3010
rect 3143 3006 3147 3010
rect 3231 3006 3235 3010
rect 3487 3078 3491 3082
rect 3575 3078 3579 3082
rect 3319 3006 3323 3010
rect 3479 3006 3483 3010
rect 3575 3006 3579 3010
rect 1863 2930 1867 2934
rect 1895 2930 1899 2934
rect 2031 2930 2035 2934
rect 2167 2930 2171 2934
rect 2175 2930 2179 2934
rect 2295 2930 2299 2934
rect 2423 2930 2427 2934
rect 2495 2930 2499 2934
rect 2543 2930 2547 2934
rect 2671 2930 2675 2934
rect 2815 2930 2819 2934
rect 2823 2930 2827 2934
rect 2975 2930 2979 2934
rect 3151 2930 3155 2934
rect 3167 2930 3171 2934
rect 3327 2930 3331 2934
rect 3487 2930 3491 2934
rect 3575 2930 3579 2934
rect 1191 2886 1195 2890
rect 1279 2886 1283 2890
rect 1311 2886 1315 2890
rect 1415 2886 1419 2890
rect 1423 2886 1427 2890
rect 1535 2886 1539 2890
rect 1551 2886 1555 2890
rect 1647 2886 1651 2890
rect 1735 2886 1739 2890
rect 1823 2886 1827 2890
rect 1167 2864 1171 2868
rect 1511 2864 1515 2868
rect 1863 2862 1867 2866
rect 1887 2862 1891 2866
rect 2023 2862 2027 2866
rect 2167 2862 2171 2866
rect 2191 2862 2195 2866
rect 2359 2862 2363 2866
rect 2487 2862 2491 2866
rect 2519 2862 2523 2866
rect 2671 2862 2675 2866
rect 2807 2862 2811 2866
rect 2815 2862 2819 2866
rect 2935 2862 2939 2866
rect 3055 2862 3059 2866
rect 1079 2810 1083 2814
rect 1135 2810 1139 2814
rect 1207 2810 1211 2814
rect 1271 2810 1275 2814
rect 1343 2810 1347 2814
rect 1407 2810 1411 2814
rect 1543 2810 1547 2814
rect 1823 2810 1827 2814
rect 1863 2794 1867 2798
rect 1895 2794 1899 2798
rect 2031 2794 2035 2798
rect 2063 2794 2067 2798
rect 183 2752 187 2756
rect 111 2734 115 2738
rect 143 2734 147 2738
rect 175 2734 179 2738
rect 231 2734 235 2738
rect 303 2734 307 2738
rect 351 2734 355 2738
rect 647 2752 651 2756
rect 3159 2862 3163 2866
rect 3167 2862 3171 2866
rect 3279 2862 3283 2866
rect 3391 2862 3395 2866
rect 3479 2862 3483 2866
rect 3575 2862 3579 2866
rect 2199 2794 2203 2798
rect 2255 2794 2259 2798
rect 2367 2794 2371 2798
rect 2439 2794 2443 2798
rect 2527 2794 2531 2798
rect 2615 2794 2619 2798
rect 2679 2794 2683 2798
rect 2783 2794 2787 2798
rect 2815 2794 2819 2798
rect 2935 2794 2939 2798
rect 2943 2794 2947 2798
rect 3063 2794 3067 2798
rect 3079 2794 3083 2798
rect 3175 2794 3179 2798
rect 3223 2794 3227 2798
rect 3287 2794 3291 2798
rect 3367 2794 3371 2798
rect 3399 2794 3403 2798
rect 431 2734 435 2738
rect 479 2734 483 2738
rect 567 2734 571 2738
rect 615 2734 619 2738
rect 703 2734 707 2738
rect 759 2734 763 2738
rect 831 2734 835 2738
rect 903 2734 907 2738
rect 959 2734 963 2738
rect 1047 2734 1051 2738
rect 1087 2734 1091 2738
rect 1215 2734 1219 2738
rect 1351 2734 1355 2738
rect 1823 2734 1827 2738
rect 1863 2722 1867 2726
rect 1887 2722 1891 2726
rect 2047 2722 2051 2726
rect 2055 2722 2059 2726
rect 2207 2722 2211 2726
rect 2247 2722 2251 2726
rect 2359 2722 2363 2726
rect 2431 2722 2435 2726
rect 2495 2722 2499 2726
rect 3487 2794 3491 2798
rect 3575 2794 3579 2798
rect 2607 2722 2611 2726
rect 2623 2722 2627 2726
rect 2743 2722 2747 2726
rect 2775 2722 2779 2726
rect 2863 2722 2867 2726
rect 2927 2722 2931 2726
rect 111 2662 115 2666
rect 135 2662 139 2666
rect 223 2662 227 2666
rect 231 2662 235 2666
rect 343 2662 347 2666
rect 351 2662 355 2666
rect 471 2662 475 2666
rect 583 2662 587 2666
rect 607 2662 611 2666
rect 695 2662 699 2666
rect 751 2662 755 2666
rect 799 2662 803 2666
rect 895 2662 899 2666
rect 903 2662 907 2666
rect 999 2662 1003 2666
rect 1039 2662 1043 2666
rect 1103 2662 1107 2666
rect 1207 2662 1211 2666
rect 1311 2662 1315 2666
rect 1823 2662 1827 2666
rect 1863 2646 1867 2650
rect 1895 2646 1899 2650
rect 1999 2646 2003 2650
rect 2055 2646 2059 2650
rect 2119 2646 2123 2650
rect 2215 2646 2219 2650
rect 2239 2646 2243 2650
rect 111 2590 115 2594
rect 143 2590 147 2594
rect 239 2590 243 2594
rect 271 2590 275 2594
rect 359 2590 363 2594
rect 415 2590 419 2594
rect 479 2590 483 2594
rect 551 2590 555 2594
rect 591 2590 595 2594
rect 679 2590 683 2594
rect 703 2590 707 2594
rect 111 2522 115 2526
rect 135 2522 139 2526
rect 263 2522 267 2526
rect 279 2522 283 2526
rect 407 2522 411 2526
rect 439 2522 443 2526
rect 543 2522 547 2526
rect 591 2522 595 2526
rect 807 2590 811 2594
rect 911 2590 915 2594
rect 927 2590 931 2594
rect 1007 2590 1011 2594
rect 1047 2590 1051 2594
rect 1111 2590 1115 2594
rect 1175 2590 1179 2594
rect 1215 2590 1219 2594
rect 671 2522 675 2526
rect 735 2522 739 2526
rect 799 2522 803 2526
rect 2351 2646 2355 2650
rect 2367 2646 2371 2650
rect 2455 2646 2459 2650
rect 2503 2646 2507 2650
rect 2551 2646 2555 2650
rect 2631 2646 2635 2650
rect 2655 2646 2659 2650
rect 2983 2722 2987 2726
rect 3071 2722 3075 2726
rect 3103 2722 3107 2726
rect 3215 2722 3219 2726
rect 3359 2722 3363 2726
rect 3479 2722 3483 2726
rect 3575 2722 3579 2726
rect 2751 2646 2755 2650
rect 2759 2646 2763 2650
rect 2863 2646 2867 2650
rect 2871 2646 2875 2650
rect 2991 2646 2995 2650
rect 3111 2646 3115 2650
rect 3575 2646 3579 2650
rect 1319 2590 1323 2594
rect 1823 2590 1827 2594
rect 1863 2574 1867 2578
rect 1887 2574 1891 2578
rect 1991 2574 1995 2578
rect 2111 2574 2115 2578
rect 2231 2574 2235 2578
rect 2343 2574 2347 2578
rect 2351 2574 2355 2578
rect 2447 2574 2451 2578
rect 2471 2574 2475 2578
rect 871 2522 875 2526
rect 919 2522 923 2526
rect 1007 2522 1011 2526
rect 1039 2522 1043 2526
rect 1143 2522 1147 2526
rect 1167 2522 1171 2526
rect 1279 2522 1283 2526
rect 1823 2522 1827 2526
rect 1007 2464 1011 2468
rect 111 2454 115 2458
rect 143 2454 147 2458
rect 191 2454 195 2458
rect 287 2454 291 2458
rect 319 2454 323 2458
rect 447 2454 451 2458
rect 455 2454 459 2458
rect 591 2454 595 2458
rect 599 2454 603 2458
rect 727 2454 731 2458
rect 743 2454 747 2458
rect 111 2374 115 2378
rect 159 2374 163 2378
rect 183 2374 187 2378
rect 247 2374 251 2378
rect 311 2374 315 2378
rect 335 2374 339 2378
rect 439 2374 443 2378
rect 447 2374 451 2378
rect 559 2374 563 2378
rect 583 2374 587 2378
rect 687 2374 691 2378
rect 719 2374 723 2378
rect 863 2454 867 2458
rect 879 2454 883 2458
rect 999 2454 1003 2458
rect 815 2374 819 2378
rect 855 2374 859 2378
rect 1863 2502 1867 2506
rect 1895 2502 1899 2506
rect 1999 2502 2003 2506
rect 2031 2502 2035 2506
rect 2119 2502 2123 2506
rect 2191 2502 2195 2506
rect 2239 2502 2243 2506
rect 1219 2464 1223 2468
rect 2543 2574 2547 2578
rect 2591 2574 2595 2578
rect 2647 2574 2651 2578
rect 2711 2574 2715 2578
rect 2751 2574 2755 2578
rect 2831 2574 2835 2578
rect 2855 2574 2859 2578
rect 3575 2574 3579 2578
rect 2495 2520 2499 2524
rect 2343 2502 2347 2506
rect 2359 2502 2363 2506
rect 2479 2502 2483 2506
rect 2487 2502 2491 2506
rect 2779 2520 2783 2524
rect 2599 2502 2603 2506
rect 2623 2502 2627 2506
rect 2719 2502 2723 2506
rect 2751 2502 2755 2506
rect 2839 2502 2843 2506
rect 2879 2502 2883 2506
rect 3015 2502 3019 2506
rect 3575 2502 3579 2506
rect 1015 2454 1019 2458
rect 1135 2454 1139 2458
rect 1151 2454 1155 2458
rect 1271 2454 1275 2458
rect 1287 2454 1291 2458
rect 1407 2454 1411 2458
rect 1823 2454 1827 2458
rect 1863 2434 1867 2438
rect 1887 2434 1891 2438
rect 2015 2434 2019 2438
rect 2023 2434 2027 2438
rect 1135 2384 1139 2388
rect 951 2374 955 2378
rect 991 2374 995 2378
rect 1079 2374 1083 2378
rect 1127 2374 1131 2378
rect 1339 2384 1343 2388
rect 1207 2374 1211 2378
rect 1263 2374 1267 2378
rect 1327 2374 1331 2378
rect 1399 2374 1403 2378
rect 1455 2374 1459 2378
rect 1583 2374 1587 2378
rect 1823 2374 1827 2378
rect 1863 2362 1867 2366
rect 1895 2362 1899 2366
rect 1927 2362 1931 2366
rect 1183 2312 1187 2316
rect 111 2298 115 2302
rect 167 2298 171 2302
rect 255 2298 259 2302
rect 343 2298 347 2302
rect 447 2298 451 2302
rect 567 2298 571 2302
rect 695 2298 699 2302
rect 823 2298 827 2302
rect 863 2298 867 2302
rect 959 2298 963 2302
rect 1023 2298 1027 2302
rect 1087 2298 1091 2302
rect 1175 2298 1179 2302
rect 703 2291 707 2292
rect 703 2288 707 2291
rect 939 2288 943 2292
rect 111 2222 115 2226
rect 535 2222 539 2226
rect 687 2222 691 2226
rect 719 2222 723 2226
rect 855 2222 859 2226
rect 895 2222 899 2226
rect 1015 2222 1019 2226
rect 2175 2434 2179 2438
rect 2183 2434 2187 2438
rect 2335 2434 2339 2438
rect 2479 2434 2483 2438
rect 2495 2434 2499 2438
rect 2615 2434 2619 2438
rect 2647 2434 2651 2438
rect 2743 2434 2747 2438
rect 2799 2434 2803 2438
rect 2871 2434 2875 2438
rect 2951 2434 2955 2438
rect 2711 2392 2715 2396
rect 2663 2376 2667 2380
rect 2023 2362 2027 2366
rect 2087 2362 2091 2366
rect 2183 2362 2187 2366
rect 2247 2362 2251 2366
rect 2343 2362 2347 2366
rect 2407 2362 2411 2366
rect 2503 2362 2507 2366
rect 1523 2312 1527 2316
rect 2559 2362 2563 2366
rect 2655 2362 2659 2366
rect 2703 2362 2707 2366
rect 1215 2298 1219 2302
rect 1319 2298 1323 2302
rect 1335 2298 1339 2302
rect 1463 2298 1467 2302
rect 1591 2298 1595 2302
rect 1599 2298 1603 2302
rect 1735 2298 1739 2302
rect 1823 2298 1827 2302
rect 1863 2290 1867 2294
rect 1919 2290 1923 2294
rect 1975 2290 1979 2294
rect 2079 2290 2083 2294
rect 2143 2290 2147 2294
rect 2239 2290 2243 2294
rect 2311 2290 2315 2294
rect 2399 2290 2403 2294
rect 2479 2290 2483 2294
rect 2551 2290 2555 2294
rect 3007 2434 3011 2438
rect 3111 2434 3115 2438
rect 3575 2434 3579 2438
rect 3019 2392 3023 2396
rect 2967 2376 2971 2380
rect 2807 2362 2811 2366
rect 2831 2362 2835 2366
rect 2951 2362 2955 2366
rect 2959 2362 2963 2366
rect 3071 2362 3075 2366
rect 3119 2362 3123 2366
rect 3183 2362 3187 2366
rect 3287 2362 3291 2366
rect 3399 2362 3403 2366
rect 3487 2362 3491 2366
rect 3575 2362 3579 2366
rect 2639 2290 2643 2294
rect 2695 2290 2699 2294
rect 2783 2290 2787 2294
rect 2823 2290 2827 2294
rect 2919 2290 2923 2294
rect 2943 2290 2947 2294
rect 3039 2290 3043 2294
rect 3063 2290 3067 2294
rect 3159 2290 3163 2294
rect 3175 2290 3179 2294
rect 1071 2222 1075 2226
rect 1167 2222 1171 2226
rect 1239 2222 1243 2226
rect 1311 2222 1315 2226
rect 1407 2222 1411 2226
rect 1455 2222 1459 2226
rect 1575 2222 1579 2226
rect 1591 2222 1595 2226
rect 1255 2176 1259 2180
rect 111 2154 115 2158
rect 495 2154 499 2158
rect 543 2154 547 2158
rect 551 2147 555 2148
rect 551 2144 555 2147
rect 623 2154 627 2158
rect 727 2154 731 2158
rect 759 2154 763 2158
rect 895 2154 899 2158
rect 903 2154 907 2158
rect 1039 2154 1043 2158
rect 1079 2154 1083 2158
rect 1183 2154 1187 2158
rect 1247 2154 1251 2158
rect 1327 2154 1331 2158
rect 1415 2154 1419 2158
rect 1471 2154 1475 2158
rect 1583 2154 1587 2158
rect 1623 2154 1627 2158
rect 767 2144 771 2148
rect 575 2112 579 2116
rect 111 2082 115 2086
rect 319 2082 323 2086
rect 431 2082 435 2086
rect 487 2082 491 2086
rect 551 2082 555 2086
rect 615 2082 619 2086
rect 679 2082 683 2086
rect 751 2082 755 2086
rect 1039 2107 1043 2108
rect 1039 2104 1043 2107
rect 1727 2222 1731 2226
rect 1823 2222 1827 2226
rect 1863 2222 1867 2226
rect 1983 2222 1987 2226
rect 2007 2222 2011 2226
rect 2799 2232 2803 2236
rect 2151 2222 2155 2226
rect 2167 2222 2171 2226
rect 2319 2222 2323 2226
rect 2335 2222 2339 2226
rect 2487 2222 2491 2226
rect 2519 2222 2523 2226
rect 2647 2222 2651 2226
rect 2711 2222 2715 2226
rect 2791 2222 2795 2226
rect 2903 2222 2907 2226
rect 2927 2222 2931 2226
rect 3047 2222 3051 2226
rect 3103 2222 3107 2226
rect 1667 2176 1671 2180
rect 1735 2154 1739 2158
rect 1823 2154 1827 2158
rect 1863 2146 1867 2150
rect 1999 2146 2003 2150
rect 2023 2146 2027 2150
rect 2159 2146 2163 2150
rect 2167 2146 2171 2150
rect 799 2082 803 2086
rect 887 2082 891 2086
rect 919 2082 923 2086
rect 1031 2082 1035 2086
rect 1039 2082 1043 2086
rect 1159 2082 1163 2086
rect 1175 2082 1179 2086
rect 1279 2082 1283 2086
rect 1319 2082 1323 2086
rect 111 2010 115 2014
rect 183 2010 187 2014
rect 295 2010 299 2014
rect 327 2010 331 2014
rect 415 2010 419 2014
rect 439 2010 443 2014
rect 535 2010 539 2014
rect 559 2010 563 2014
rect 655 2010 659 2014
rect 687 2010 691 2014
rect 775 2010 779 2014
rect 807 2010 811 2014
rect 895 2010 899 2014
rect 927 2010 931 2014
rect 1015 2010 1019 2014
rect 1047 2010 1051 2014
rect 1407 2082 1411 2086
rect 1463 2082 1467 2086
rect 1615 2082 1619 2086
rect 1823 2082 1827 2086
rect 2319 2146 2323 2150
rect 2327 2146 2331 2150
rect 2471 2146 2475 2150
rect 2511 2146 2515 2150
rect 2615 2146 2619 2150
rect 2703 2146 2707 2150
rect 2759 2146 2763 2150
rect 3271 2290 3275 2294
rect 3279 2290 3283 2294
rect 3383 2290 3387 2294
rect 3391 2290 3395 2294
rect 3479 2290 3483 2294
rect 3575 2290 3579 2294
rect 3183 2232 3187 2236
rect 3167 2222 3171 2226
rect 3279 2222 3283 2226
rect 3303 2222 3307 2226
rect 3391 2222 3395 2226
rect 3487 2222 3491 2226
rect 3575 2222 3579 2226
rect 2895 2146 2899 2150
rect 3023 2146 3027 2150
rect 3095 2146 3099 2150
rect 3143 2146 3147 2150
rect 3263 2146 3267 2150
rect 3295 2146 3299 2150
rect 3383 2146 3387 2150
rect 3479 2146 3483 2150
rect 3575 2146 3579 2150
rect 1863 2074 1867 2078
rect 1983 2074 1987 2078
rect 2031 2074 2035 2078
rect 2143 2074 2147 2078
rect 2175 2074 2179 2078
rect 2311 2074 2315 2078
rect 2327 2074 2331 2078
rect 2471 2074 2475 2078
rect 2479 2074 2483 2078
rect 2623 2074 2627 2078
rect 2631 2074 2635 2078
rect 2767 2074 2771 2078
rect 2775 2074 2779 2078
rect 1135 2010 1139 2014
rect 1167 2010 1171 2014
rect 1255 2010 1259 2014
rect 1287 2010 1291 2014
rect 1415 2010 1419 2014
rect 1823 2010 1827 2014
rect 239 1960 243 1964
rect 563 1960 567 1964
rect 111 1938 115 1942
rect 135 1938 139 1942
rect 175 1938 179 1942
rect 223 1938 227 1942
rect 287 1938 291 1942
rect 351 1938 355 1942
rect 407 1938 411 1942
rect 495 1938 499 1942
rect 527 1938 531 1942
rect 1863 2006 1867 2010
rect 1887 2006 1891 2010
rect 1975 2006 1979 2010
rect 2031 2006 2035 2010
rect 2135 2006 2139 2010
rect 2199 2006 2203 2010
rect 2303 2006 2307 2010
rect 2375 2006 2379 2010
rect 2463 2006 2467 2010
rect 2543 2006 2547 2010
rect 2903 2074 2907 2078
rect 2911 2074 2915 2078
rect 3031 2074 3035 2078
rect 3039 2074 3043 2078
rect 3151 2074 3155 2078
rect 3159 2074 3163 2078
rect 3271 2074 3275 2078
rect 3279 2074 3283 2078
rect 3391 2074 3395 2078
rect 3487 2074 3491 2078
rect 3575 2074 3579 2078
rect 2623 2006 2627 2010
rect 2711 2006 2715 2010
rect 2767 2006 2771 2010
rect 2871 2006 2875 2010
rect 2903 2006 2907 2010
rect 3031 2006 3035 2010
rect 3039 2006 3043 2010
rect 3151 2006 3155 2010
rect 3207 2006 3211 2010
rect 3271 2006 3275 2010
rect 3383 2006 3387 2010
rect 3479 2006 3483 2010
rect 3575 2006 3579 2010
rect 647 1938 651 1942
rect 655 1938 659 1942
rect 767 1938 771 1942
rect 839 1938 843 1942
rect 887 1938 891 1942
rect 1007 1938 1011 1942
rect 1039 1938 1043 1942
rect 1127 1938 1131 1942
rect 1247 1938 1251 1942
rect 1463 1938 1467 1942
rect 1823 1938 1827 1942
rect 1863 1930 1867 1934
rect 1895 1930 1899 1934
rect 111 1862 115 1866
rect 951 1880 955 1884
rect 143 1862 147 1866
rect 231 1862 235 1866
rect 271 1862 275 1866
rect 359 1862 363 1866
rect 415 1862 419 1866
rect 503 1862 507 1866
rect 559 1862 563 1866
rect 663 1862 667 1866
rect 695 1862 699 1866
rect 823 1862 827 1866
rect 847 1862 851 1866
rect 943 1862 947 1866
rect 111 1782 115 1786
rect 135 1782 139 1786
rect 263 1782 267 1786
rect 303 1782 307 1786
rect 1991 1930 1995 1934
rect 2039 1930 2043 1934
rect 2119 1930 2123 1934
rect 2207 1930 2211 1934
rect 2255 1930 2259 1934
rect 2727 1952 2731 1956
rect 2383 1930 2387 1934
rect 2511 1930 2515 1934
rect 2551 1930 2555 1934
rect 2631 1930 2635 1934
rect 2719 1930 2723 1934
rect 2751 1930 2755 1934
rect 2879 1930 2883 1934
rect 1159 1880 1163 1884
rect 1047 1862 1051 1866
rect 1055 1862 1059 1866
rect 1159 1862 1163 1866
rect 1255 1862 1259 1866
rect 1263 1862 1267 1866
rect 1359 1862 1363 1866
rect 1455 1862 1459 1866
rect 407 1782 411 1786
rect 495 1782 499 1786
rect 111 1710 115 1714
rect 551 1782 555 1786
rect 687 1782 691 1786
rect 815 1782 819 1786
rect 871 1782 875 1786
rect 935 1782 939 1786
rect 1047 1782 1051 1786
rect 1471 1862 1475 1866
rect 1551 1862 1555 1866
rect 1647 1862 1651 1866
rect 1735 1862 1739 1866
rect 1823 1862 1827 1866
rect 1863 1854 1867 1858
rect 1887 1854 1891 1858
rect 1983 1854 1987 1858
rect 2111 1854 2115 1858
rect 2223 1854 2227 1858
rect 2247 1854 2251 1858
rect 2359 1854 2363 1858
rect 3159 1952 3163 1956
rect 3007 1930 3011 1934
rect 3047 1930 3051 1934
rect 3215 1930 3219 1934
rect 3575 1930 3579 1934
rect 2375 1854 2379 1858
rect 2495 1854 2499 1858
rect 2503 1854 2507 1858
rect 1151 1782 1155 1786
rect 1215 1782 1219 1786
rect 1255 1782 1259 1786
rect 1351 1782 1355 1786
rect 1375 1782 1379 1786
rect 143 1710 147 1714
rect 287 1710 291 1714
rect 311 1710 315 1714
rect 471 1710 475 1714
rect 503 1710 507 1714
rect 655 1710 659 1714
rect 695 1710 699 1714
rect 839 1710 843 1714
rect 879 1710 883 1714
rect 1023 1710 1027 1714
rect 1055 1710 1059 1714
rect 111 1634 115 1638
rect 135 1634 139 1638
rect 271 1634 275 1638
rect 279 1634 283 1638
rect 447 1634 451 1638
rect 463 1634 467 1638
rect 631 1634 635 1638
rect 647 1634 651 1638
rect 815 1634 819 1638
rect 831 1634 835 1638
rect 991 1634 995 1638
rect 1447 1782 1451 1786
rect 1535 1782 1539 1786
rect 1543 1782 1547 1786
rect 1639 1782 1643 1786
rect 1703 1782 1707 1786
rect 1727 1782 1731 1786
rect 1823 1782 1827 1786
rect 1863 1782 1867 1786
rect 2231 1782 2235 1786
rect 2271 1782 2275 1786
rect 2623 1854 2627 1858
rect 2743 1854 2747 1858
rect 2863 1854 2867 1858
rect 2871 1854 2875 1858
rect 2991 1854 2995 1858
rect 2999 1854 3003 1858
rect 3575 1854 3579 1858
rect 2359 1782 2363 1786
rect 2367 1782 2371 1786
rect 2455 1782 2459 1786
rect 2503 1782 2507 1786
rect 2559 1782 2563 1786
rect 2631 1782 2635 1786
rect 2663 1782 2667 1786
rect 2751 1782 2755 1786
rect 2759 1782 2763 1786
rect 2863 1782 2867 1786
rect 2871 1782 2875 1786
rect 2967 1782 2971 1786
rect 2999 1782 3003 1786
rect 3071 1782 3075 1786
rect 3175 1782 3179 1786
rect 3575 1782 3579 1786
rect 1191 1710 1195 1714
rect 1223 1710 1227 1714
rect 1359 1710 1363 1714
rect 1383 1710 1387 1714
rect 1527 1710 1531 1714
rect 1543 1710 1547 1714
rect 1695 1710 1699 1714
rect 1711 1710 1715 1714
rect 1823 1710 1827 1714
rect 1863 1710 1867 1714
rect 2247 1710 2251 1714
rect 2263 1710 2267 1714
rect 2351 1710 2355 1714
rect 2367 1710 2371 1714
rect 2447 1710 2451 1714
rect 2495 1710 2499 1714
rect 2551 1710 2555 1714
rect 2623 1710 2627 1714
rect 2655 1710 2659 1714
rect 2751 1710 2755 1714
rect 2759 1710 2763 1714
rect 2855 1710 2859 1714
rect 2887 1710 2891 1714
rect 1015 1634 1019 1638
rect 1151 1634 1155 1638
rect 2959 1710 2963 1714
rect 3015 1710 3019 1714
rect 3063 1710 3067 1714
rect 3135 1710 3139 1714
rect 3167 1710 3171 1714
rect 3247 1710 3251 1714
rect 3367 1710 3371 1714
rect 3479 1710 3483 1714
rect 3575 1710 3579 1714
rect 1183 1634 1187 1638
rect 1303 1634 1307 1638
rect 1351 1634 1355 1638
rect 1455 1634 1459 1638
rect 1519 1634 1523 1638
rect 1599 1634 1603 1638
rect 1687 1634 1691 1638
rect 1727 1634 1731 1638
rect 1823 1634 1827 1638
rect 1863 1638 1867 1642
rect 2151 1638 2155 1642
rect 2255 1638 2259 1642
rect 2343 1638 2347 1642
rect 2375 1638 2379 1642
rect 2503 1638 2507 1642
rect 2527 1638 2531 1642
rect 2631 1638 2635 1642
rect 2703 1638 2707 1642
rect 2767 1638 2771 1642
rect 2871 1638 2875 1642
rect 2895 1638 2899 1642
rect 3023 1638 3027 1642
rect 3031 1638 3035 1642
rect 3143 1638 3147 1642
rect 111 1566 115 1570
rect 143 1566 147 1570
rect 271 1566 275 1570
rect 279 1566 283 1570
rect 431 1566 435 1570
rect 455 1566 459 1570
rect 599 1566 603 1570
rect 639 1566 643 1570
rect 767 1566 771 1570
rect 823 1566 827 1570
rect 935 1566 939 1570
rect 999 1566 1003 1570
rect 111 1494 115 1498
rect 135 1494 139 1498
rect 183 1494 187 1498
rect 263 1494 267 1498
rect 327 1494 331 1498
rect 111 1418 115 1422
rect 423 1494 427 1498
rect 471 1494 475 1498
rect 591 1494 595 1498
rect 607 1494 611 1498
rect 743 1494 747 1498
rect 759 1494 763 1498
rect 871 1494 875 1498
rect 927 1494 931 1498
rect 1103 1566 1107 1570
rect 1159 1566 1163 1570
rect 1263 1566 1267 1570
rect 1311 1566 1315 1570
rect 1423 1566 1427 1570
rect 1463 1566 1467 1570
rect 1591 1566 1595 1570
rect 1607 1566 1611 1570
rect 1735 1566 1739 1570
rect 1823 1566 1827 1570
rect 1863 1570 1867 1574
rect 2087 1570 2091 1574
rect 2143 1570 2147 1574
rect 991 1494 995 1498
rect 1095 1494 1099 1498
rect 1119 1494 1123 1498
rect 1247 1494 1251 1498
rect 1255 1494 1259 1498
rect 1375 1494 1379 1498
rect 191 1418 195 1422
rect 199 1418 203 1422
rect 335 1418 339 1422
rect 463 1418 467 1422
rect 479 1418 483 1422
rect 583 1418 587 1422
rect 615 1418 619 1422
rect 703 1418 707 1422
rect 111 1346 115 1350
rect 191 1346 195 1350
rect 231 1346 235 1350
rect 751 1418 755 1422
rect 815 1418 819 1422
rect 879 1418 883 1422
rect 919 1418 923 1422
rect 999 1418 1003 1422
rect 1015 1418 1019 1422
rect 327 1346 331 1350
rect 383 1346 387 1350
rect 455 1346 459 1350
rect 543 1346 547 1350
rect 575 1346 579 1350
rect 695 1346 699 1350
rect 703 1346 707 1350
rect 1415 1494 1419 1498
rect 1583 1494 1587 1498
rect 1727 1494 1731 1498
rect 3191 1638 3195 1642
rect 3255 1638 3259 1642
rect 3351 1638 3355 1642
rect 3375 1638 3379 1642
rect 3487 1638 3491 1642
rect 2279 1570 2283 1574
rect 2335 1570 2339 1574
rect 2455 1570 2459 1574
rect 2519 1570 2523 1574
rect 2623 1570 2627 1574
rect 2695 1570 2699 1574
rect 2791 1570 2795 1574
rect 2863 1570 2867 1574
rect 2951 1570 2955 1574
rect 3023 1570 3027 1574
rect 3111 1570 3115 1574
rect 3183 1570 3187 1574
rect 3271 1570 3275 1574
rect 3343 1570 3347 1574
rect 3431 1570 3435 1574
rect 1823 1494 1827 1498
rect 1863 1494 1867 1498
rect 1895 1494 1899 1498
rect 1991 1494 1995 1498
rect 2095 1494 2099 1498
rect 2119 1494 2123 1498
rect 2639 1512 2643 1516
rect 2247 1494 2251 1498
rect 2287 1494 2291 1498
rect 2383 1494 2387 1498
rect 2463 1494 2467 1498
rect 2535 1494 2539 1498
rect 2631 1494 2635 1498
rect 2703 1494 2707 1498
rect 2799 1494 2803 1498
rect 1119 1418 1123 1422
rect 1127 1418 1131 1422
rect 1223 1418 1227 1422
rect 1255 1418 1259 1422
rect 1327 1418 1331 1422
rect 1383 1418 1387 1422
rect 1823 1418 1827 1422
rect 1863 1422 1867 1426
rect 1887 1422 1891 1426
rect 1975 1422 1979 1426
rect 1983 1422 1987 1426
rect 2071 1422 2075 1426
rect 2111 1422 2115 1426
rect 2183 1422 2187 1426
rect 2239 1422 2243 1426
rect 2303 1422 2307 1426
rect 2375 1422 2379 1426
rect 2887 1494 2891 1498
rect 2959 1494 2963 1498
rect 3215 1512 3219 1516
rect 3087 1494 3091 1498
rect 3119 1494 3123 1498
rect 3279 1494 3283 1498
rect 3295 1494 3299 1498
rect 3439 1494 3443 1498
rect 3479 1570 3483 1574
rect 3575 1638 3579 1642
rect 3575 1570 3579 1574
rect 3487 1494 3491 1498
rect 3575 1494 3579 1498
rect 2439 1422 2443 1426
rect 2527 1422 2531 1426
rect 2607 1422 2611 1426
rect 2695 1422 2699 1426
rect 2807 1422 2811 1426
rect 2879 1422 2883 1426
rect 3031 1422 3035 1426
rect 3079 1422 3083 1426
rect 3263 1422 3267 1426
rect 3287 1422 3291 1426
rect 3479 1422 3483 1426
rect 3575 1422 3579 1426
rect 807 1346 811 1350
rect 871 1346 875 1350
rect 911 1346 915 1350
rect 1007 1346 1011 1350
rect 1039 1346 1043 1350
rect 1111 1346 1115 1350
rect 1207 1346 1211 1350
rect 1215 1346 1219 1350
rect 1319 1346 1323 1350
rect 559 1288 563 1292
rect 799 1288 803 1292
rect 1375 1346 1379 1350
rect 1823 1346 1827 1350
rect 1863 1350 1867 1354
rect 1895 1350 1899 1354
rect 1983 1350 1987 1354
rect 2079 1350 2083 1354
rect 2103 1350 2107 1354
rect 2191 1350 2195 1354
rect 2223 1350 2227 1354
rect 2311 1350 2315 1354
rect 2359 1350 2363 1354
rect 2775 1363 2779 1364
rect 2775 1360 2779 1363
rect 3211 1360 3215 1364
rect 2447 1350 2451 1354
rect 2511 1350 2515 1354
rect 2615 1350 2619 1354
rect 2687 1350 2691 1354
rect 2815 1350 2819 1354
rect 2871 1350 2875 1354
rect 3039 1350 3043 1354
rect 3071 1350 3075 1354
rect 3271 1350 3275 1354
rect 3279 1350 3283 1354
rect 111 1278 115 1282
rect 215 1278 219 1282
rect 239 1278 243 1282
rect 359 1278 363 1282
rect 391 1278 395 1282
rect 519 1278 523 1282
rect 551 1278 555 1282
rect 679 1278 683 1282
rect 711 1278 715 1282
rect 839 1278 843 1282
rect 879 1278 883 1282
rect 111 1202 115 1206
rect 135 1202 139 1206
rect 999 1278 1003 1282
rect 1047 1278 1051 1282
rect 1151 1278 1155 1282
rect 1215 1278 1219 1282
rect 1295 1278 1299 1282
rect 1383 1278 1387 1282
rect 1439 1278 1443 1282
rect 1591 1278 1595 1282
rect 1823 1278 1827 1282
rect 1863 1270 1867 1274
rect 1887 1270 1891 1274
rect 1975 1270 1979 1274
rect 2055 1270 2059 1274
rect 2095 1270 2099 1274
rect 2143 1270 2147 1274
rect 2215 1270 2219 1274
rect 2239 1270 2243 1274
rect 2335 1270 2339 1274
rect 2351 1270 2355 1274
rect 2431 1270 2435 1274
rect 2503 1270 2507 1274
rect 2551 1270 2555 1274
rect 2679 1270 2683 1274
rect 2687 1270 2691 1274
rect 2855 1270 2859 1274
rect 2863 1270 2867 1274
rect 2567 1256 2571 1260
rect 3039 1270 3043 1274
rect 3063 1270 3067 1274
rect 3231 1270 3235 1274
rect 2959 1256 2963 1260
rect 207 1202 211 1206
rect 271 1202 275 1206
rect 351 1202 355 1206
rect 423 1202 427 1206
rect 511 1202 515 1206
rect 575 1202 579 1206
rect 671 1202 675 1206
rect 727 1202 731 1206
rect 831 1202 835 1206
rect 887 1202 891 1206
rect 991 1202 995 1206
rect 1055 1202 1059 1206
rect 1143 1202 1147 1206
rect 1231 1202 1235 1206
rect 1287 1202 1291 1206
rect 1415 1202 1419 1206
rect 1431 1202 1435 1206
rect 1583 1202 1587 1206
rect 111 1134 115 1138
rect 143 1134 147 1138
rect 279 1134 283 1138
rect 295 1134 299 1138
rect 431 1134 435 1138
rect 479 1134 483 1138
rect 583 1134 587 1138
rect 1599 1202 1603 1206
rect 1823 1202 1827 1206
rect 1863 1198 1867 1202
rect 2039 1198 2043 1202
rect 2063 1198 2067 1202
rect 2151 1198 2155 1202
rect 2247 1198 2251 1202
rect 2279 1198 2283 1202
rect 2343 1198 2347 1202
rect 2415 1198 2419 1202
rect 2439 1198 2443 1202
rect 2559 1198 2563 1202
rect 2695 1198 2699 1202
rect 2711 1198 2715 1202
rect 2863 1198 2867 1202
rect 3015 1198 3019 1202
rect 3047 1198 3051 1202
rect 663 1134 667 1138
rect 735 1134 739 1138
rect 847 1134 851 1138
rect 895 1134 899 1138
rect 1031 1134 1035 1138
rect 1063 1134 1067 1138
rect 1207 1134 1211 1138
rect 1239 1134 1243 1138
rect 111 1066 115 1070
rect 135 1066 139 1070
rect 271 1066 275 1070
rect 287 1066 291 1070
rect 431 1066 435 1070
rect 471 1066 475 1070
rect 583 1066 587 1070
rect 655 1066 659 1070
rect 735 1066 739 1070
rect 839 1066 843 1070
rect 887 1066 891 1070
rect 1391 1134 1395 1138
rect 1423 1134 1427 1138
rect 1575 1134 1579 1138
rect 1607 1134 1611 1138
rect 1735 1134 1739 1138
rect 1823 1134 1827 1138
rect 1863 1118 1867 1122
rect 1943 1118 1947 1122
rect 1023 1066 1027 1070
rect 1047 1066 1051 1070
rect 1199 1066 1203 1070
rect 1215 1066 1219 1070
rect 1383 1066 1387 1070
rect 1559 1066 1563 1070
rect 1567 1066 1571 1070
rect 1727 1066 1731 1070
rect 1823 1066 1827 1070
rect 111 994 115 998
rect 143 994 147 998
rect 279 994 283 998
rect 287 994 291 998
rect 439 994 443 998
rect 463 994 467 998
rect 591 994 595 998
rect 647 994 651 998
rect 743 994 747 998
rect 1063 1008 1067 1012
rect 2031 1118 2035 1122
rect 2087 1118 2091 1122
rect 2143 1118 2147 1122
rect 2231 1118 2235 1122
rect 2271 1118 2275 1122
rect 2383 1118 2387 1122
rect 2407 1118 2411 1122
rect 2535 1118 2539 1122
rect 3167 1198 3171 1202
rect 3239 1198 3243 1202
rect 3487 1350 3491 1354
rect 3575 1350 3579 1354
rect 3271 1270 3275 1274
rect 3431 1270 3435 1274
rect 3479 1270 3483 1274
rect 3575 1270 3579 1274
rect 3327 1198 3331 1202
rect 3439 1198 3443 1202
rect 3487 1198 3491 1202
rect 3575 1198 3579 1202
rect 2551 1118 2555 1122
rect 2687 1118 2691 1122
rect 2703 1118 2707 1122
rect 1863 1038 1867 1042
rect 1919 1038 1923 1042
rect 1951 1038 1955 1042
rect 2095 1038 2099 1042
rect 2127 1038 2131 1042
rect 1283 1008 1287 1012
rect 823 994 827 998
rect 895 994 899 998
rect 999 994 1003 998
rect 1055 994 1059 998
rect 1167 994 1171 998
rect 1223 994 1227 998
rect 111 918 115 922
rect 135 918 139 922
rect 271 918 275 922
rect 279 918 283 922
rect 439 918 443 922
rect 455 918 459 922
rect 607 918 611 922
rect 639 918 643 922
rect 775 918 779 922
rect 815 918 819 922
rect 935 918 939 922
rect 991 918 995 922
rect 1327 994 1331 998
rect 1391 994 1395 998
rect 1487 994 1491 998
rect 1567 994 1571 998
rect 2839 1118 2843 1122
rect 2855 1118 2859 1122
rect 2991 1118 2995 1122
rect 3007 1118 3011 1122
rect 3151 1118 3155 1122
rect 3159 1118 3163 1122
rect 3319 1118 3323 1122
rect 3479 1118 3483 1122
rect 3575 1118 3579 1122
rect 2703 1048 2707 1052
rect 2239 1038 2243 1042
rect 2327 1038 2331 1042
rect 2391 1038 2395 1042
rect 2519 1038 2523 1042
rect 2543 1038 2547 1042
rect 2695 1038 2699 1042
rect 1655 994 1659 998
rect 1735 994 1739 998
rect 1823 994 1827 998
rect 1863 966 1867 970
rect 1887 966 1891 970
rect 1095 918 1099 922
rect 1159 918 1163 922
rect 1247 918 1251 922
rect 1319 918 1323 922
rect 1399 918 1403 922
rect 1479 918 1483 922
rect 1551 918 1555 922
rect 1647 918 1651 922
rect 1823 918 1827 922
rect 111 850 115 854
rect 143 850 147 854
rect 279 850 283 854
rect 287 850 291 854
rect 455 864 459 868
rect 1911 966 1915 970
rect 2071 966 2075 970
rect 2119 966 2123 970
rect 2263 966 2267 970
rect 2319 966 2323 970
rect 2455 966 2459 970
rect 2511 966 2515 970
rect 3079 1048 3083 1052
rect 2847 1038 2851 1042
rect 2863 1038 2867 1042
rect 2999 1038 3003 1042
rect 3023 1038 3027 1042
rect 3159 1038 3163 1042
rect 3183 1038 3187 1042
rect 3327 1038 3331 1042
rect 3343 1038 3347 1042
rect 3487 1038 3491 1042
rect 3575 1038 3579 1042
rect 2631 966 2635 970
rect 2687 966 2691 970
rect 2799 966 2803 970
rect 2855 966 2859 970
rect 2951 966 2955 970
rect 3015 966 3019 970
rect 3095 966 3099 970
rect 1863 890 1867 894
rect 1895 890 1899 894
rect 2023 890 2027 894
rect 2079 890 2083 894
rect 707 864 711 868
rect 1263 864 1267 868
rect 1495 864 1499 868
rect 2815 912 2819 916
rect 3175 966 3179 970
rect 3231 966 3235 970
rect 3335 966 3339 970
rect 3367 966 3371 970
rect 3479 966 3483 970
rect 3575 966 3579 970
rect 3111 912 3115 916
rect 2183 890 2187 894
rect 2271 890 2275 894
rect 2351 890 2355 894
rect 2463 890 2467 894
rect 2519 890 2523 894
rect 2639 890 2643 894
rect 2687 890 2691 894
rect 2807 890 2811 894
rect 2839 890 2843 894
rect 2959 890 2963 894
rect 2983 890 2987 894
rect 3103 890 3107 894
rect 3119 890 3123 894
rect 3239 890 3243 894
rect 3247 890 3251 894
rect 3375 890 3379 894
rect 447 850 451 854
rect 463 850 467 854
rect 615 850 619 854
rect 639 850 643 854
rect 783 850 787 854
rect 807 850 811 854
rect 943 850 947 854
rect 983 850 987 854
rect 1103 850 1107 854
rect 1159 850 1163 854
rect 1255 850 1259 854
rect 1335 850 1339 854
rect 1407 850 1411 854
rect 1511 850 1515 854
rect 1559 850 1563 854
rect 1823 850 1827 854
rect 111 778 115 782
rect 135 778 139 782
rect 271 778 275 782
rect 279 778 283 782
rect 439 778 443 782
rect 455 778 459 782
rect 607 778 611 782
rect 631 778 635 782
rect 775 778 779 782
rect 111 706 115 710
rect 143 706 147 710
rect 799 778 803 782
rect 935 778 939 782
rect 975 778 979 782
rect 1087 778 1091 782
rect 1151 778 1155 782
rect 1863 814 1867 818
rect 1887 814 1891 818
rect 2015 814 2019 818
rect 2071 814 2075 818
rect 2175 814 2179 818
rect 2263 814 2267 818
rect 2343 814 2347 818
rect 2447 814 2451 818
rect 2511 814 2515 818
rect 2623 814 2627 818
rect 2679 814 2683 818
rect 1239 778 1243 782
rect 3487 890 3491 894
rect 3575 890 3579 894
rect 2791 814 2795 818
rect 1327 778 1331 782
rect 1391 778 1395 782
rect 1503 778 1507 782
rect 1551 778 1555 782
rect 1823 778 1827 782
rect 1863 746 1867 750
rect 1895 746 1899 750
rect 279 706 283 710
rect 287 706 291 710
rect 447 706 451 710
rect 455 706 459 710
rect 615 706 619 710
rect 623 706 627 710
rect 783 706 787 710
rect 791 706 795 710
rect 943 706 947 710
rect 959 706 963 710
rect 1095 706 1099 710
rect 1119 706 1123 710
rect 1247 706 1251 710
rect 1279 706 1283 710
rect 1399 706 1403 710
rect 1439 706 1443 710
rect 1559 706 1563 710
rect 1599 706 1603 710
rect 2831 814 2835 818
rect 2943 814 2947 818
rect 2975 814 2979 818
rect 3087 814 3091 818
rect 3111 814 3115 818
rect 3223 814 3227 818
rect 3239 814 3243 818
rect 3359 814 3363 818
rect 3367 814 3371 818
rect 3479 814 3483 818
rect 3575 814 3579 818
rect 2071 746 2075 750
rect 2079 746 2083 750
rect 2263 746 2267 750
rect 2271 746 2275 750
rect 2447 746 2451 750
rect 2455 746 2459 750
rect 2623 746 2627 750
rect 2631 746 2635 750
rect 2799 746 2803 750
rect 2951 746 2955 750
rect 2975 746 2979 750
rect 3095 746 3099 750
rect 3151 746 3155 750
rect 1823 706 1827 710
rect 1863 674 1867 678
rect 1887 674 1891 678
rect 1975 674 1979 678
rect 2063 674 2067 678
rect 2095 674 2099 678
rect 111 630 115 634
rect 135 630 139 634
rect 279 630 283 634
rect 287 630 291 634
rect 447 630 451 634
rect 455 630 459 634
rect 615 630 619 634
rect 631 630 635 634
rect 783 630 787 634
rect 799 630 803 634
rect 951 630 955 634
rect 967 630 971 634
rect 1111 630 1115 634
rect 1119 630 1123 634
rect 1271 630 1275 634
rect 1415 630 1419 634
rect 1431 630 1435 634
rect 1559 630 1563 634
rect 1591 630 1595 634
rect 1711 630 1715 634
rect 1823 630 1827 634
rect 2223 674 2227 678
rect 2255 674 2259 678
rect 2351 674 2355 678
rect 2439 674 2443 678
rect 3055 739 3059 740
rect 3055 736 3059 739
rect 3231 746 3235 750
rect 3327 746 3331 750
rect 3367 746 3371 750
rect 3259 736 3263 740
rect 3487 746 3491 750
rect 3575 746 3579 750
rect 2479 674 2483 678
rect 2615 674 2619 678
rect 2767 674 2771 678
rect 2791 674 2795 678
rect 2935 674 2939 678
rect 2967 674 2971 678
rect 3119 674 3123 678
rect 3143 674 3147 678
rect 3311 674 3315 678
rect 3319 674 3323 678
rect 3479 674 3483 678
rect 3575 674 3579 678
rect 1863 602 1867 606
rect 1895 602 1899 606
rect 1983 602 1987 606
rect 2047 602 2051 606
rect 2103 602 2107 606
rect 1199 584 1203 588
rect 1639 584 1643 588
rect 111 558 115 562
rect 143 558 147 562
rect 151 558 155 562
rect 295 558 299 562
rect 311 558 315 562
rect 463 558 467 562
rect 471 558 475 562
rect 631 558 635 562
rect 639 558 643 562
rect 783 558 787 562
rect 807 558 811 562
rect 927 558 931 562
rect 975 558 979 562
rect 1063 558 1067 562
rect 1127 558 1131 562
rect 1191 558 1195 562
rect 111 482 115 486
rect 143 482 147 486
rect 159 482 163 486
rect 303 482 307 486
rect 311 482 315 486
rect 463 482 467 486
rect 615 482 619 486
rect 623 482 627 486
rect 759 482 763 486
rect 775 482 779 486
rect 111 414 115 418
rect 151 414 155 418
rect 167 414 171 418
rect 271 414 275 418
rect 319 414 323 418
rect 407 414 411 418
rect 471 414 475 418
rect 887 482 891 486
rect 919 482 923 486
rect 1007 482 1011 486
rect 1055 482 1059 486
rect 1279 558 1283 562
rect 1311 558 1315 562
rect 1423 558 1427 562
rect 1535 558 1539 562
rect 1567 558 1571 562
rect 1647 558 1651 562
rect 1719 558 1723 562
rect 1735 558 1739 562
rect 1823 558 1827 562
rect 1127 482 1131 486
rect 1183 482 1187 486
rect 1239 482 1243 486
rect 1303 482 1307 486
rect 1343 482 1347 486
rect 1415 482 1419 486
rect 1439 482 1443 486
rect 1143 424 1147 428
rect 551 414 555 418
rect 623 414 627 418
rect 711 414 715 418
rect 767 414 771 418
rect 887 414 891 418
rect 895 414 899 418
rect 1015 414 1019 418
rect 1063 414 1067 418
rect 1135 414 1139 418
rect 1247 414 1251 418
rect 1351 414 1355 418
rect 903 392 907 396
rect 159 384 163 388
rect 339 384 343 388
rect 111 330 115 334
rect 135 330 139 334
rect 143 330 147 334
rect 223 330 227 334
rect 263 330 267 334
rect 311 330 315 334
rect 399 330 403 334
rect 487 330 491 334
rect 543 330 547 334
rect 575 330 579 334
rect 663 330 667 334
rect 703 330 707 334
rect 751 330 755 334
rect 839 330 843 334
rect 111 258 115 262
rect 143 258 147 262
rect 231 258 235 262
rect 319 258 323 262
rect 407 258 411 262
rect 495 258 499 262
rect 583 258 587 262
rect 671 258 675 262
rect 879 330 883 334
rect 927 330 931 334
rect 1015 330 1019 334
rect 1055 330 1059 334
rect 1863 526 1867 530
rect 1887 526 1891 530
rect 2039 526 2043 530
rect 2631 616 2635 620
rect 2215 602 2219 606
rect 2231 602 2235 606
rect 2359 602 2363 606
rect 2391 602 2395 606
rect 2487 602 2491 606
rect 2583 602 2587 606
rect 2623 602 2627 606
rect 2775 602 2779 606
rect 2799 602 2803 606
rect 3235 616 3239 620
rect 2943 602 2947 606
rect 3023 602 3027 606
rect 3127 602 3131 606
rect 3255 602 3259 606
rect 3319 602 3323 606
rect 3487 602 3491 606
rect 3575 602 3579 606
rect 2191 526 2195 530
rect 2207 526 2211 530
rect 2279 526 2283 530
rect 2375 526 2379 530
rect 2383 526 2387 530
rect 2487 526 2491 530
rect 2575 526 2579 530
rect 2631 526 2635 530
rect 2791 526 2795 530
rect 2807 526 2811 530
rect 3007 526 3011 530
rect 3015 526 3019 530
rect 3215 526 3219 530
rect 3247 526 3251 530
rect 3431 526 3435 530
rect 3479 526 3483 530
rect 3575 526 3579 530
rect 1527 482 1531 486
rect 1543 482 1547 486
rect 1639 482 1643 486
rect 1727 482 1731 486
rect 1823 482 1827 486
rect 2391 488 2395 492
rect 3187 491 3191 492
rect 3187 488 3191 491
rect 1863 450 1867 454
rect 1895 450 1899 454
rect 2039 450 2043 454
rect 2199 450 2203 454
rect 2207 450 2211 454
rect 2287 450 2291 454
rect 2383 450 2387 454
rect 1491 424 1495 428
rect 1439 414 1443 418
rect 1447 414 1451 418
rect 1551 414 1555 418
rect 1639 414 1643 418
rect 1647 414 1651 418
rect 1735 414 1739 418
rect 1823 414 1827 418
rect 1163 392 1167 396
rect 1863 382 1867 386
rect 1887 382 1891 386
rect 1975 382 1979 386
rect 2031 382 2035 386
rect 2063 382 2067 386
rect 2151 382 2155 386
rect 2199 382 2203 386
rect 1103 330 1107 334
rect 1191 330 1195 334
rect 1239 330 1243 334
rect 1287 330 1291 334
rect 1383 330 1387 334
rect 1431 330 1435 334
rect 1479 330 1483 334
rect 1575 330 1579 334
rect 1631 330 1635 334
rect 1671 330 1675 334
rect 1823 330 1827 334
rect 1863 314 1867 318
rect 1895 314 1899 318
rect 759 258 763 262
rect 847 258 851 262
rect 935 258 939 262
rect 1023 258 1027 262
rect 1111 258 1115 262
rect 1031 251 1035 252
rect 1031 248 1035 251
rect 1303 272 1307 276
rect 1563 272 1567 276
rect 2495 450 2499 454
rect 2575 450 2579 454
rect 2639 450 2643 454
rect 2783 450 2787 454
rect 2815 450 2819 454
rect 3007 450 3011 454
rect 3015 450 3019 454
rect 3223 450 3227 454
rect 3239 450 3243 454
rect 3439 450 3443 454
rect 3471 450 3475 454
rect 3575 450 3579 454
rect 2263 382 2267 386
rect 2375 382 2379 386
rect 2383 382 2387 386
rect 2519 382 2523 386
rect 2567 382 2571 386
rect 2671 382 2675 386
rect 2775 382 2779 386
rect 2847 382 2851 386
rect 2999 382 3003 386
rect 3031 382 3035 386
rect 2703 344 2707 348
rect 3159 347 3163 348
rect 2687 328 2691 332
rect 1983 314 1987 318
rect 2071 314 2075 318
rect 2159 314 2163 318
rect 2247 314 2251 318
rect 2271 314 2275 318
rect 2359 314 2363 318
rect 2391 314 2395 318
rect 2471 314 2475 318
rect 2527 314 2531 318
rect 2367 307 2371 308
rect 2367 304 2371 307
rect 2583 314 2587 318
rect 2679 314 2683 318
rect 2695 314 2699 318
rect 2543 304 2547 308
rect 1199 258 1203 262
rect 1287 258 1291 262
rect 1295 258 1299 262
rect 1375 258 1379 262
rect 1391 258 1395 262
rect 1463 258 1467 262
rect 1487 258 1491 262
rect 1551 258 1555 262
rect 1583 258 1587 262
rect 1639 258 1643 262
rect 1679 258 1683 262
rect 1727 258 1731 262
rect 1823 258 1827 262
rect 1267 248 1271 252
rect 1863 246 1867 250
rect 1887 246 1891 250
rect 1975 246 1979 250
rect 2063 246 2067 250
rect 2151 246 2155 250
rect 2239 246 2243 250
rect 2263 246 2267 250
rect 2351 246 2355 250
rect 2399 246 2403 250
rect 2463 246 2467 250
rect 2535 246 2539 250
rect 2575 246 2579 250
rect 3159 344 3163 347
rect 3231 382 3235 386
rect 3431 382 3435 386
rect 3463 382 3467 386
rect 3179 328 3183 332
rect 2807 314 2811 318
rect 2855 314 2859 318
rect 2919 314 2923 318
rect 3039 314 3043 318
rect 3159 314 3163 318
rect 3239 314 3243 318
rect 2679 246 2683 250
rect 2687 246 2691 250
rect 2799 246 2803 250
rect 2815 246 2819 250
rect 2911 246 2915 250
rect 2951 246 2955 250
rect 3031 246 3035 250
rect 3087 246 3091 250
rect 1903 224 1907 228
rect 2227 224 2231 228
rect 111 190 115 194
rect 135 190 139 194
rect 223 190 227 194
rect 311 190 315 194
rect 399 190 403 194
rect 487 190 491 194
rect 575 190 579 194
rect 663 190 667 194
rect 751 190 755 194
rect 839 190 843 194
rect 927 190 931 194
rect 1015 190 1019 194
rect 1103 190 1107 194
rect 1191 190 1195 194
rect 1279 190 1283 194
rect 1367 190 1371 194
rect 1455 190 1459 194
rect 1543 190 1547 194
rect 1631 190 1635 194
rect 1719 190 1723 194
rect 1823 190 1827 194
rect 2791 176 2795 180
rect 1863 146 1867 150
rect 1895 146 1899 150
rect 1983 146 1987 150
rect 2071 146 2075 150
rect 2159 146 2163 150
rect 2271 146 2275 150
rect 2407 146 2411 150
rect 2543 146 2547 150
rect 2687 146 2691 150
rect 2783 146 2787 150
rect 2831 192 2835 196
rect 3151 246 3155 250
rect 3223 246 3227 250
rect 3359 246 3363 250
rect 3439 314 3443 318
rect 3107 192 3111 196
rect 3191 176 3195 180
rect 3575 382 3579 386
rect 3575 314 3579 318
rect 3479 246 3483 250
rect 3575 246 3579 250
rect 2823 146 2827 150
rect 2871 146 2875 150
rect 2959 146 2963 150
rect 3047 146 3051 150
rect 3095 146 3099 150
rect 3135 146 3139 150
rect 3223 146 3227 150
rect 3231 146 3235 150
rect 3311 146 3315 150
rect 3367 146 3371 150
rect 3399 146 3403 150
rect 3487 146 3491 150
rect 3575 146 3579 150
rect 1863 78 1867 82
rect 2775 78 2779 82
rect 2863 78 2867 82
rect 2951 78 2955 82
rect 3039 78 3043 82
rect 3127 78 3131 82
rect 3215 78 3219 82
rect 3303 78 3307 82
rect 3391 78 3395 82
rect 3479 78 3483 82
rect 3575 78 3579 82
<< m4 >>
rect 84 3665 85 3671
rect 91 3670 1835 3671
rect 91 3666 111 3670
rect 115 3666 135 3670
rect 139 3666 223 3670
rect 227 3666 1823 3670
rect 1827 3666 1835 3670
rect 91 3665 1835 3666
rect 1841 3665 1842 3671
rect 1834 3607 1835 3613
rect 1841 3607 1866 3613
rect 96 3597 97 3603
rect 103 3602 1847 3603
rect 103 3598 111 3602
rect 115 3598 143 3602
rect 147 3598 231 3602
rect 235 3598 319 3602
rect 323 3598 407 3602
rect 411 3598 495 3602
rect 499 3598 1823 3602
rect 1827 3598 1847 3602
rect 103 3597 1847 3598
rect 1853 3597 1854 3603
rect 1860 3595 1866 3607
rect 1860 3594 3599 3595
rect 1860 3590 1863 3594
rect 1867 3590 1887 3594
rect 1891 3590 1975 3594
rect 1979 3590 2063 3594
rect 2067 3590 2151 3594
rect 2155 3590 2239 3594
rect 2243 3590 2327 3594
rect 2331 3590 2431 3594
rect 2435 3590 2535 3594
rect 2539 3590 2631 3594
rect 2635 3590 2727 3594
rect 2731 3590 2823 3594
rect 2827 3590 2919 3594
rect 2923 3590 3015 3594
rect 3019 3590 3119 3594
rect 3123 3590 3223 3594
rect 3227 3590 3575 3594
rect 3579 3590 3599 3594
rect 1860 3589 3599 3590
rect 3605 3589 3606 3595
rect 2110 3556 2116 3557
rect 2498 3556 2504 3557
rect 2110 3552 2111 3556
rect 2115 3552 2499 3556
rect 2503 3552 2504 3556
rect 2110 3551 2116 3552
rect 2498 3551 2504 3552
rect 84 3529 85 3535
rect 91 3534 1835 3535
rect 91 3530 111 3534
rect 115 3530 135 3534
rect 139 3530 223 3534
rect 227 3530 247 3534
rect 251 3530 311 3534
rect 315 3530 375 3534
rect 379 3530 399 3534
rect 403 3530 487 3534
rect 491 3530 503 3534
rect 507 3530 623 3534
rect 627 3530 743 3534
rect 747 3530 863 3534
rect 867 3530 975 3534
rect 979 3530 1079 3534
rect 1083 3530 1175 3534
rect 1179 3530 1271 3534
rect 1275 3530 1367 3534
rect 1371 3530 1471 3534
rect 1475 3530 1575 3534
rect 1579 3530 1823 3534
rect 1827 3530 1835 3534
rect 91 3529 1835 3530
rect 1841 3529 1842 3535
rect 1846 3521 1847 3527
rect 1853 3526 3611 3527
rect 1853 3522 1863 3526
rect 1867 3522 1895 3526
rect 1899 3522 1983 3526
rect 1987 3522 2071 3526
rect 2075 3522 2103 3526
rect 2107 3522 2159 3526
rect 2163 3522 2231 3526
rect 2235 3522 2247 3526
rect 2251 3522 2335 3526
rect 2339 3522 2367 3526
rect 2371 3522 2439 3526
rect 2443 3522 2511 3526
rect 2515 3522 2543 3526
rect 2547 3522 2639 3526
rect 2643 3522 2655 3526
rect 2659 3522 2735 3526
rect 2739 3522 2791 3526
rect 2795 3522 2831 3526
rect 2835 3522 2927 3526
rect 2931 3522 2935 3526
rect 2939 3522 3023 3526
rect 3027 3522 3079 3526
rect 3083 3522 3127 3526
rect 3131 3522 3223 3526
rect 3227 3522 3231 3526
rect 3235 3522 3575 3526
rect 3579 3522 3611 3526
rect 1853 3521 3611 3522
rect 3617 3521 3618 3527
rect 96 3461 97 3467
rect 103 3466 1847 3467
rect 103 3462 111 3466
rect 115 3462 175 3466
rect 179 3462 255 3466
rect 259 3462 303 3466
rect 307 3462 383 3466
rect 387 3462 447 3466
rect 451 3462 511 3466
rect 515 3462 591 3466
rect 595 3462 631 3466
rect 635 3462 743 3466
rect 747 3462 751 3466
rect 755 3462 871 3466
rect 875 3462 895 3466
rect 899 3462 983 3466
rect 987 3462 1039 3466
rect 1043 3462 1087 3466
rect 1091 3462 1183 3466
rect 1187 3462 1279 3466
rect 1283 3462 1327 3466
rect 1331 3462 1375 3466
rect 1379 3462 1479 3466
rect 1483 3462 1583 3466
rect 1587 3462 1823 3466
rect 1827 3462 1847 3466
rect 103 3461 1847 3462
rect 1853 3461 1854 3467
rect 1834 3445 1835 3451
rect 1841 3450 3599 3451
rect 1841 3446 1863 3450
rect 1867 3446 1887 3450
rect 1891 3446 1975 3450
rect 1979 3446 2023 3450
rect 2027 3446 2095 3450
rect 2099 3446 2191 3450
rect 2195 3446 2223 3450
rect 2227 3446 2359 3450
rect 2363 3446 2367 3450
rect 2371 3446 2503 3450
rect 2507 3446 2543 3450
rect 2547 3446 2647 3450
rect 2651 3446 2711 3450
rect 2715 3446 2783 3450
rect 2787 3446 2871 3450
rect 2875 3446 2927 3450
rect 2931 3446 3031 3450
rect 3035 3446 3071 3450
rect 3075 3446 3191 3450
rect 3195 3446 3215 3450
rect 3219 3446 3359 3450
rect 3363 3446 3575 3450
rect 3579 3446 3599 3450
rect 1841 3445 3599 3446
rect 3605 3445 3606 3451
rect 1438 3436 1444 3437
rect 1470 3436 1476 3437
rect 1438 3432 1439 3436
rect 1443 3432 1471 3436
rect 1475 3432 1476 3436
rect 1438 3431 1444 3432
rect 1470 3431 1476 3432
rect 84 3393 85 3399
rect 91 3398 1835 3399
rect 91 3394 111 3398
rect 115 3394 135 3398
rect 139 3394 167 3398
rect 171 3394 263 3398
rect 267 3394 295 3398
rect 299 3394 407 3398
rect 411 3394 439 3398
rect 443 3394 567 3398
rect 571 3394 583 3398
rect 587 3394 727 3398
rect 731 3394 735 3398
rect 739 3394 887 3398
rect 891 3394 1031 3398
rect 1035 3394 1047 3398
rect 1051 3394 1175 3398
rect 1179 3394 1207 3398
rect 1211 3394 1319 3398
rect 1323 3394 1367 3398
rect 1371 3394 1471 3398
rect 1475 3394 1527 3398
rect 1531 3394 1823 3398
rect 1827 3394 1835 3398
rect 91 3393 1835 3394
rect 1841 3393 1842 3399
rect 3046 3396 3052 3397
rect 3258 3396 3264 3397
rect 3046 3392 3047 3396
rect 3051 3392 3259 3396
rect 3263 3392 3264 3396
rect 3046 3391 3052 3392
rect 3258 3391 3264 3392
rect 1846 3369 1847 3375
rect 1853 3374 3611 3375
rect 1853 3370 1863 3374
rect 1867 3370 1895 3374
rect 1899 3370 2031 3374
rect 2035 3370 2199 3374
rect 2203 3370 2375 3374
rect 2379 3370 2551 3374
rect 2555 3370 2719 3374
rect 2723 3370 2879 3374
rect 2883 3370 3039 3374
rect 3043 3370 3191 3374
rect 3195 3370 3199 3374
rect 3203 3370 3343 3374
rect 3347 3370 3367 3374
rect 3371 3370 3487 3374
rect 3491 3370 3575 3374
rect 3579 3370 3611 3374
rect 1853 3369 3611 3370
rect 3617 3369 3618 3375
rect 214 3340 220 3341
rect 682 3340 688 3341
rect 214 3336 215 3340
rect 219 3336 683 3340
rect 687 3336 688 3340
rect 214 3335 220 3336
rect 682 3335 688 3336
rect 96 3321 97 3327
rect 103 3326 1847 3327
rect 103 3322 111 3326
rect 115 3322 143 3326
rect 147 3322 207 3326
rect 211 3322 271 3326
rect 275 3322 335 3326
rect 339 3322 415 3326
rect 419 3322 479 3326
rect 483 3322 575 3326
rect 579 3322 639 3326
rect 643 3322 735 3326
rect 739 3322 807 3326
rect 811 3322 895 3326
rect 899 3322 983 3326
rect 987 3322 1055 3326
rect 1059 3322 1167 3326
rect 1171 3322 1215 3326
rect 1219 3322 1351 3326
rect 1355 3322 1375 3326
rect 1379 3322 1535 3326
rect 1539 3322 1543 3326
rect 1547 3322 1823 3326
rect 1827 3322 1847 3326
rect 103 3321 1847 3322
rect 1853 3321 1854 3327
rect 1834 3301 1835 3307
rect 1841 3306 3599 3307
rect 1841 3302 1863 3306
rect 1867 3302 1887 3306
rect 1891 3302 2007 3306
rect 2011 3302 2023 3306
rect 2027 3302 2151 3306
rect 2155 3302 2191 3306
rect 2195 3302 2303 3306
rect 2307 3302 2367 3306
rect 2371 3302 2463 3306
rect 2467 3302 2543 3306
rect 2547 3302 2631 3306
rect 2635 3302 2711 3306
rect 2715 3302 2799 3306
rect 2803 3302 2871 3306
rect 2875 3302 2967 3306
rect 2971 3302 3031 3306
rect 3035 3302 3135 3306
rect 3139 3302 3183 3306
rect 3187 3302 3311 3306
rect 3315 3302 3335 3306
rect 3339 3302 3479 3306
rect 3483 3302 3575 3306
rect 3579 3302 3599 3306
rect 1841 3301 3599 3302
rect 3605 3301 3606 3307
rect 2182 3276 2188 3277
rect 2538 3276 2544 3277
rect 2182 3272 2183 3276
rect 2187 3272 2539 3276
rect 2543 3272 2544 3276
rect 2182 3271 2188 3272
rect 2538 3271 2544 3272
rect 84 3249 85 3255
rect 91 3254 1835 3255
rect 91 3250 111 3254
rect 115 3250 199 3254
rect 203 3250 327 3254
rect 331 3250 367 3254
rect 371 3250 471 3254
rect 475 3250 503 3254
rect 507 3250 631 3254
rect 635 3250 639 3254
rect 643 3250 783 3254
rect 787 3250 799 3254
rect 803 3250 935 3254
rect 939 3250 975 3254
rect 979 3250 1095 3254
rect 1099 3250 1159 3254
rect 1163 3250 1255 3254
rect 1259 3250 1343 3254
rect 1347 3250 1415 3254
rect 1419 3250 1535 3254
rect 1539 3250 1575 3254
rect 1579 3250 1823 3254
rect 1827 3250 1835 3254
rect 91 3249 1835 3250
rect 1841 3249 1842 3255
rect 2166 3252 2172 3253
rect 2478 3252 2484 3253
rect 2166 3248 2167 3252
rect 2171 3248 2479 3252
rect 2483 3248 2484 3252
rect 2166 3247 2172 3248
rect 2478 3247 2484 3248
rect 1846 3225 1847 3231
rect 1853 3230 3611 3231
rect 1853 3226 1863 3230
rect 1867 3226 1895 3230
rect 1899 3226 2015 3230
rect 2019 3226 2023 3230
rect 2027 3226 2159 3230
rect 2163 3226 2175 3230
rect 2179 3226 2311 3230
rect 2315 3226 2327 3230
rect 2331 3226 2463 3230
rect 2467 3226 2471 3230
rect 2475 3226 2599 3230
rect 2603 3226 2639 3230
rect 2643 3226 2735 3230
rect 2739 3226 2807 3230
rect 2811 3226 2871 3230
rect 2875 3226 2975 3230
rect 2979 3226 3015 3230
rect 3019 3226 3143 3230
rect 3147 3226 3167 3230
rect 3171 3226 3319 3230
rect 3323 3226 3327 3230
rect 3331 3226 3487 3230
rect 3491 3226 3575 3230
rect 3579 3226 3611 3230
rect 1853 3225 3611 3226
rect 3617 3225 3618 3231
rect 950 3204 956 3205
rect 1162 3204 1168 3205
rect 950 3200 951 3204
rect 955 3200 1163 3204
rect 1167 3200 1168 3204
rect 950 3199 956 3200
rect 1162 3199 1168 3200
rect 486 3196 492 3197
rect 710 3196 716 3197
rect 486 3192 487 3196
rect 491 3192 711 3196
rect 715 3192 716 3196
rect 486 3191 492 3192
rect 710 3191 716 3192
rect 96 3173 97 3179
rect 103 3178 1847 3179
rect 103 3174 111 3178
rect 115 3174 375 3178
rect 379 3174 447 3178
rect 451 3174 511 3178
rect 515 3174 559 3178
rect 563 3174 647 3178
rect 651 3174 687 3178
rect 691 3174 791 3178
rect 795 3174 823 3178
rect 827 3174 943 3178
rect 947 3174 975 3178
rect 979 3174 1103 3178
rect 1107 3174 1135 3178
rect 1139 3174 1263 3178
rect 1267 3174 1295 3178
rect 1299 3174 1423 3178
rect 1427 3174 1463 3178
rect 1467 3174 1583 3178
rect 1587 3174 1639 3178
rect 1643 3174 1823 3178
rect 1827 3174 1847 3178
rect 103 3173 1847 3174
rect 1853 3173 1854 3179
rect 1834 3153 1835 3159
rect 1841 3158 3599 3159
rect 1841 3154 1863 3158
rect 1867 3154 1887 3158
rect 1891 3154 2015 3158
rect 2019 3154 2047 3158
rect 2051 3154 2167 3158
rect 2171 3154 2199 3158
rect 2203 3154 2319 3158
rect 2323 3154 2351 3158
rect 2355 3154 2455 3158
rect 2459 3154 2511 3158
rect 2515 3154 2591 3158
rect 2595 3154 2679 3158
rect 2683 3154 2727 3158
rect 2731 3154 2863 3158
rect 2867 3154 2871 3158
rect 2875 3154 3007 3158
rect 3011 3154 3071 3158
rect 3075 3154 3159 3158
rect 3163 3154 3287 3158
rect 3291 3154 3319 3158
rect 3323 3154 3479 3158
rect 3483 3154 3575 3158
rect 3579 3154 3599 3158
rect 1841 3153 3599 3154
rect 3605 3153 3606 3159
rect 84 3097 85 3103
rect 91 3102 1835 3103
rect 91 3098 111 3102
rect 115 3098 439 3102
rect 443 3098 551 3102
rect 555 3098 663 3102
rect 667 3098 679 3102
rect 683 3098 783 3102
rect 787 3098 815 3102
rect 819 3098 903 3102
rect 907 3098 967 3102
rect 971 3098 1031 3102
rect 1035 3098 1127 3102
rect 1131 3098 1159 3102
rect 1163 3098 1287 3102
rect 1291 3098 1423 3102
rect 1427 3098 1455 3102
rect 1459 3098 1559 3102
rect 1563 3098 1631 3102
rect 1635 3098 1695 3102
rect 1699 3098 1823 3102
rect 1827 3098 1835 3102
rect 91 3097 1835 3098
rect 1841 3097 1842 3103
rect 2214 3100 2220 3101
rect 2530 3100 2536 3101
rect 2214 3096 2215 3100
rect 2219 3096 2531 3100
rect 2535 3096 2536 3100
rect 2214 3095 2220 3096
rect 2530 3095 2536 3096
rect 1846 3077 1847 3083
rect 1853 3082 3611 3083
rect 1853 3078 1863 3082
rect 1867 3078 1895 3082
rect 1899 3078 1919 3082
rect 1923 3078 2055 3082
rect 2059 3078 2087 3082
rect 2091 3078 2207 3082
rect 2211 3078 2279 3082
rect 2283 3078 2359 3082
rect 2363 3078 2487 3082
rect 2491 3078 2519 3082
rect 2523 3078 2687 3082
rect 2691 3078 2719 3082
rect 2723 3078 2879 3082
rect 2883 3078 2975 3082
rect 2979 3078 3079 3082
rect 3083 3078 3239 3082
rect 3243 3078 3295 3082
rect 3299 3078 3487 3082
rect 3491 3078 3575 3082
rect 3579 3078 3611 3082
rect 1853 3077 3611 3078
rect 3617 3077 3618 3083
rect 566 3076 572 3077
rect 890 3076 896 3077
rect 566 3072 567 3076
rect 571 3072 891 3076
rect 895 3072 896 3076
rect 566 3071 572 3072
rect 890 3071 896 3072
rect 2502 3052 2508 3053
rect 2898 3052 2904 3053
rect 2502 3048 2503 3052
rect 2507 3048 2899 3052
rect 2903 3048 2904 3052
rect 2502 3047 2508 3048
rect 2898 3047 2904 3048
rect 96 3025 97 3031
rect 103 3030 1847 3031
rect 103 3026 111 3030
rect 115 3026 559 3030
rect 563 3026 575 3030
rect 579 3026 671 3030
rect 675 3026 703 3030
rect 707 3026 791 3030
rect 795 3026 831 3030
rect 835 3026 911 3030
rect 915 3026 967 3030
rect 971 3026 1039 3030
rect 1043 3026 1103 3030
rect 1107 3026 1167 3030
rect 1171 3026 1239 3030
rect 1243 3026 1295 3030
rect 1299 3026 1367 3030
rect 1371 3026 1431 3030
rect 1435 3026 1495 3030
rect 1499 3026 1567 3030
rect 1571 3026 1623 3030
rect 1627 3026 1703 3030
rect 1707 3026 1735 3030
rect 1739 3026 1823 3030
rect 1827 3026 1847 3030
rect 103 3025 1847 3026
rect 1853 3025 1854 3031
rect 1834 3005 1835 3011
rect 1841 3010 3599 3011
rect 1841 3006 1863 3010
rect 1867 3006 1911 3010
rect 1915 3006 2023 3010
rect 2027 3006 2079 3010
rect 2083 3006 2159 3010
rect 2163 3006 2271 3010
rect 2275 3006 2287 3010
rect 2291 3006 2415 3010
rect 2419 3006 2479 3010
rect 2483 3006 2535 3010
rect 2539 3006 2663 3010
rect 2667 3006 2711 3010
rect 2715 3006 2807 3010
rect 2811 3006 2967 3010
rect 2971 3006 3143 3010
rect 3147 3006 3231 3010
rect 3235 3006 3319 3010
rect 3323 3006 3479 3010
rect 3483 3006 3575 3010
rect 3579 3006 3599 3010
rect 1841 3005 3599 3006
rect 3605 3005 3606 3011
rect 84 2957 85 2963
rect 91 2962 1835 2963
rect 91 2958 111 2962
rect 115 2958 495 2962
rect 499 2958 567 2962
rect 571 2958 639 2962
rect 643 2958 695 2962
rect 699 2958 783 2962
rect 787 2958 823 2962
rect 827 2958 919 2962
rect 923 2958 959 2962
rect 963 2958 1055 2962
rect 1059 2958 1095 2962
rect 1099 2958 1183 2962
rect 1187 2958 1231 2962
rect 1235 2958 1303 2962
rect 1307 2958 1359 2962
rect 1363 2958 1415 2962
rect 1419 2958 1487 2962
rect 1491 2958 1527 2962
rect 1531 2958 1615 2962
rect 1619 2958 1639 2962
rect 1643 2958 1727 2962
rect 1731 2958 1823 2962
rect 1827 2958 1835 2962
rect 91 2957 1835 2958
rect 1841 2957 1842 2963
rect 1846 2929 1847 2935
rect 1853 2934 3611 2935
rect 1853 2930 1863 2934
rect 1867 2930 1895 2934
rect 1899 2930 2031 2934
rect 2035 2930 2167 2934
rect 2171 2930 2175 2934
rect 2179 2930 2295 2934
rect 2299 2930 2423 2934
rect 2427 2930 2495 2934
rect 2499 2930 2543 2934
rect 2547 2930 2671 2934
rect 2675 2930 2815 2934
rect 2819 2930 2823 2934
rect 2827 2930 2975 2934
rect 2979 2930 3151 2934
rect 3155 2930 3167 2934
rect 3171 2930 3327 2934
rect 3331 2930 3487 2934
rect 3491 2930 3575 2934
rect 3579 2930 3611 2934
rect 1853 2929 3611 2930
rect 3617 2929 3618 2935
rect 96 2885 97 2891
rect 103 2890 1847 2891
rect 103 2886 111 2890
rect 115 2886 327 2890
rect 331 2886 455 2890
rect 459 2886 503 2890
rect 507 2886 591 2890
rect 595 2886 647 2890
rect 651 2886 727 2890
rect 731 2886 791 2890
rect 795 2886 871 2890
rect 875 2886 927 2890
rect 931 2886 1007 2890
rect 1011 2886 1063 2890
rect 1067 2886 1143 2890
rect 1147 2886 1191 2890
rect 1195 2886 1279 2890
rect 1283 2886 1311 2890
rect 1315 2886 1415 2890
rect 1419 2886 1423 2890
rect 1427 2886 1535 2890
rect 1539 2886 1551 2890
rect 1555 2886 1647 2890
rect 1651 2886 1735 2890
rect 1739 2886 1823 2890
rect 1827 2886 1847 2890
rect 103 2885 1847 2886
rect 1853 2885 1854 2891
rect 1166 2868 1172 2869
rect 1510 2868 1516 2869
rect 1166 2864 1167 2868
rect 1171 2864 1511 2868
rect 1515 2864 1516 2868
rect 1166 2863 1172 2864
rect 1510 2863 1516 2864
rect 1834 2861 1835 2867
rect 1841 2866 3599 2867
rect 1841 2862 1863 2866
rect 1867 2862 1887 2866
rect 1891 2862 2023 2866
rect 2027 2862 2167 2866
rect 2171 2862 2191 2866
rect 2195 2862 2359 2866
rect 2363 2862 2487 2866
rect 2491 2862 2519 2866
rect 2523 2862 2671 2866
rect 2675 2862 2807 2866
rect 2811 2862 2815 2866
rect 2819 2862 2935 2866
rect 2939 2862 3055 2866
rect 3059 2862 3159 2866
rect 3163 2862 3167 2866
rect 3171 2862 3279 2866
rect 3283 2862 3391 2866
rect 3395 2862 3479 2866
rect 3483 2862 3575 2866
rect 3579 2862 3599 2866
rect 1841 2861 3599 2862
rect 3605 2861 3606 2867
rect 84 2809 85 2815
rect 91 2814 1835 2815
rect 91 2810 111 2814
rect 115 2810 167 2814
rect 171 2810 295 2814
rect 299 2810 319 2814
rect 323 2810 423 2814
rect 427 2810 447 2814
rect 451 2810 559 2814
rect 563 2810 583 2814
rect 587 2810 695 2814
rect 699 2810 719 2814
rect 723 2810 823 2814
rect 827 2810 863 2814
rect 867 2810 951 2814
rect 955 2810 999 2814
rect 1003 2810 1079 2814
rect 1083 2810 1135 2814
rect 1139 2810 1207 2814
rect 1211 2810 1271 2814
rect 1275 2810 1343 2814
rect 1347 2810 1407 2814
rect 1411 2810 1543 2814
rect 1547 2810 1823 2814
rect 1827 2810 1835 2814
rect 91 2809 1835 2810
rect 1841 2809 1842 2815
rect 1846 2793 1847 2799
rect 1853 2798 3611 2799
rect 1853 2794 1863 2798
rect 1867 2794 1895 2798
rect 1899 2794 2031 2798
rect 2035 2794 2063 2798
rect 2067 2794 2199 2798
rect 2203 2794 2255 2798
rect 2259 2794 2367 2798
rect 2371 2794 2439 2798
rect 2443 2794 2527 2798
rect 2531 2794 2615 2798
rect 2619 2794 2679 2798
rect 2683 2794 2783 2798
rect 2787 2794 2815 2798
rect 2819 2794 2935 2798
rect 2939 2794 2943 2798
rect 2947 2794 3063 2798
rect 3067 2794 3079 2798
rect 3083 2794 3175 2798
rect 3179 2794 3223 2798
rect 3227 2794 3287 2798
rect 3291 2794 3367 2798
rect 3371 2794 3399 2798
rect 3403 2794 3487 2798
rect 3491 2794 3575 2798
rect 3579 2794 3611 2798
rect 1853 2793 3611 2794
rect 3617 2793 3618 2799
rect 182 2756 188 2757
rect 646 2756 652 2757
rect 182 2752 183 2756
rect 187 2752 647 2756
rect 651 2752 652 2756
rect 182 2751 188 2752
rect 646 2751 652 2752
rect 96 2733 97 2739
rect 103 2738 1847 2739
rect 103 2734 111 2738
rect 115 2734 143 2738
rect 147 2734 175 2738
rect 179 2734 231 2738
rect 235 2734 303 2738
rect 307 2734 351 2738
rect 355 2734 431 2738
rect 435 2734 479 2738
rect 483 2734 567 2738
rect 571 2734 615 2738
rect 619 2734 703 2738
rect 707 2734 759 2738
rect 763 2734 831 2738
rect 835 2734 903 2738
rect 907 2734 959 2738
rect 963 2734 1047 2738
rect 1051 2734 1087 2738
rect 1091 2734 1215 2738
rect 1219 2734 1351 2738
rect 1355 2734 1823 2738
rect 1827 2734 1847 2738
rect 103 2733 1847 2734
rect 1853 2733 1854 2739
rect 1834 2721 1835 2727
rect 1841 2726 3599 2727
rect 1841 2722 1863 2726
rect 1867 2722 1887 2726
rect 1891 2722 2047 2726
rect 2051 2722 2055 2726
rect 2059 2722 2207 2726
rect 2211 2722 2247 2726
rect 2251 2722 2359 2726
rect 2363 2722 2431 2726
rect 2435 2722 2495 2726
rect 2499 2722 2607 2726
rect 2611 2722 2623 2726
rect 2627 2722 2743 2726
rect 2747 2722 2775 2726
rect 2779 2722 2863 2726
rect 2867 2722 2927 2726
rect 2931 2722 2983 2726
rect 2987 2722 3071 2726
rect 3075 2722 3103 2726
rect 3107 2722 3215 2726
rect 3219 2722 3359 2726
rect 3363 2722 3479 2726
rect 3483 2722 3575 2726
rect 3579 2722 3599 2726
rect 1841 2721 3599 2722
rect 3605 2721 3606 2727
rect 84 2661 85 2667
rect 91 2666 1835 2667
rect 91 2662 111 2666
rect 115 2662 135 2666
rect 139 2662 223 2666
rect 227 2662 231 2666
rect 235 2662 343 2666
rect 347 2662 351 2666
rect 355 2662 471 2666
rect 475 2662 583 2666
rect 587 2662 607 2666
rect 611 2662 695 2666
rect 699 2662 751 2666
rect 755 2662 799 2666
rect 803 2662 895 2666
rect 899 2662 903 2666
rect 907 2662 999 2666
rect 1003 2662 1039 2666
rect 1043 2662 1103 2666
rect 1107 2662 1207 2666
rect 1211 2662 1311 2666
rect 1315 2662 1823 2666
rect 1827 2662 1835 2666
rect 91 2661 1835 2662
rect 1841 2661 1842 2667
rect 1846 2645 1847 2651
rect 1853 2650 3611 2651
rect 1853 2646 1863 2650
rect 1867 2646 1895 2650
rect 1899 2646 1999 2650
rect 2003 2646 2055 2650
rect 2059 2646 2119 2650
rect 2123 2646 2215 2650
rect 2219 2646 2239 2650
rect 2243 2646 2351 2650
rect 2355 2646 2367 2650
rect 2371 2646 2455 2650
rect 2459 2646 2503 2650
rect 2507 2646 2551 2650
rect 2555 2646 2631 2650
rect 2635 2646 2655 2650
rect 2659 2646 2751 2650
rect 2755 2646 2759 2650
rect 2763 2646 2863 2650
rect 2867 2646 2871 2650
rect 2875 2646 2991 2650
rect 2995 2646 3111 2650
rect 3115 2646 3575 2650
rect 3579 2646 3611 2650
rect 1853 2645 3611 2646
rect 3617 2645 3618 2651
rect 96 2589 97 2595
rect 103 2594 1847 2595
rect 103 2590 111 2594
rect 115 2590 143 2594
rect 147 2590 239 2594
rect 243 2590 271 2594
rect 275 2590 359 2594
rect 363 2590 415 2594
rect 419 2590 479 2594
rect 483 2590 551 2594
rect 555 2590 591 2594
rect 595 2590 679 2594
rect 683 2590 703 2594
rect 707 2590 807 2594
rect 811 2590 911 2594
rect 915 2590 927 2594
rect 931 2590 1007 2594
rect 1011 2590 1047 2594
rect 1051 2590 1111 2594
rect 1115 2590 1175 2594
rect 1179 2590 1215 2594
rect 1219 2590 1319 2594
rect 1323 2590 1823 2594
rect 1827 2590 1847 2594
rect 103 2589 1847 2590
rect 1853 2589 1854 2595
rect 1834 2573 1835 2579
rect 1841 2578 3599 2579
rect 1841 2574 1863 2578
rect 1867 2574 1887 2578
rect 1891 2574 1991 2578
rect 1995 2574 2111 2578
rect 2115 2574 2231 2578
rect 2235 2574 2343 2578
rect 2347 2574 2351 2578
rect 2355 2574 2447 2578
rect 2451 2574 2471 2578
rect 2475 2574 2543 2578
rect 2547 2574 2591 2578
rect 2595 2574 2647 2578
rect 2651 2574 2711 2578
rect 2715 2574 2751 2578
rect 2755 2574 2831 2578
rect 2835 2574 2855 2578
rect 2859 2574 3575 2578
rect 3579 2574 3599 2578
rect 1841 2573 3599 2574
rect 3605 2573 3606 2579
rect 84 2521 85 2527
rect 91 2526 1835 2527
rect 91 2522 111 2526
rect 115 2522 135 2526
rect 139 2522 263 2526
rect 267 2522 279 2526
rect 283 2522 407 2526
rect 411 2522 439 2526
rect 443 2522 543 2526
rect 547 2522 591 2526
rect 595 2522 671 2526
rect 675 2522 735 2526
rect 739 2522 799 2526
rect 803 2522 871 2526
rect 875 2522 919 2526
rect 923 2522 1007 2526
rect 1011 2522 1039 2526
rect 1043 2522 1143 2526
rect 1147 2522 1167 2526
rect 1171 2522 1279 2526
rect 1283 2522 1823 2526
rect 1827 2522 1835 2526
rect 91 2521 1835 2522
rect 1841 2521 1842 2527
rect 2494 2524 2500 2525
rect 2778 2524 2784 2525
rect 2494 2520 2495 2524
rect 2499 2520 2779 2524
rect 2783 2520 2784 2524
rect 2494 2519 2500 2520
rect 2778 2519 2784 2520
rect 1846 2501 1847 2507
rect 1853 2506 3611 2507
rect 1853 2502 1863 2506
rect 1867 2502 1895 2506
rect 1899 2502 1999 2506
rect 2003 2502 2031 2506
rect 2035 2502 2119 2506
rect 2123 2502 2191 2506
rect 2195 2502 2239 2506
rect 2243 2502 2343 2506
rect 2347 2502 2359 2506
rect 2363 2502 2479 2506
rect 2483 2502 2487 2506
rect 2491 2502 2599 2506
rect 2603 2502 2623 2506
rect 2627 2502 2719 2506
rect 2723 2502 2751 2506
rect 2755 2502 2839 2506
rect 2843 2502 2879 2506
rect 2883 2502 3015 2506
rect 3019 2502 3575 2506
rect 3579 2502 3611 2506
rect 1853 2501 3611 2502
rect 3617 2501 3618 2507
rect 1006 2468 1012 2469
rect 1218 2468 1224 2469
rect 1006 2464 1007 2468
rect 1011 2464 1219 2468
rect 1223 2464 1224 2468
rect 1006 2463 1012 2464
rect 1218 2463 1224 2464
rect 96 2453 97 2459
rect 103 2458 1847 2459
rect 103 2454 111 2458
rect 115 2454 143 2458
rect 147 2454 191 2458
rect 195 2454 287 2458
rect 291 2454 319 2458
rect 323 2454 447 2458
rect 451 2454 455 2458
rect 459 2454 591 2458
rect 595 2454 599 2458
rect 603 2454 727 2458
rect 731 2454 743 2458
rect 747 2454 863 2458
rect 867 2454 879 2458
rect 883 2454 999 2458
rect 1003 2454 1015 2458
rect 1019 2454 1135 2458
rect 1139 2454 1151 2458
rect 1155 2454 1271 2458
rect 1275 2454 1287 2458
rect 1291 2454 1407 2458
rect 1411 2454 1823 2458
rect 1827 2454 1847 2458
rect 103 2453 1847 2454
rect 1853 2453 1854 2459
rect 1834 2433 1835 2439
rect 1841 2438 3599 2439
rect 1841 2434 1863 2438
rect 1867 2434 1887 2438
rect 1891 2434 2015 2438
rect 2019 2434 2023 2438
rect 2027 2434 2175 2438
rect 2179 2434 2183 2438
rect 2187 2434 2335 2438
rect 2339 2434 2479 2438
rect 2483 2434 2495 2438
rect 2499 2434 2615 2438
rect 2619 2434 2647 2438
rect 2651 2434 2743 2438
rect 2747 2434 2799 2438
rect 2803 2434 2871 2438
rect 2875 2434 2951 2438
rect 2955 2434 3007 2438
rect 3011 2434 3111 2438
rect 3115 2434 3575 2438
rect 3579 2434 3599 2438
rect 1841 2433 3599 2434
rect 3605 2433 3606 2439
rect 2710 2396 2716 2397
rect 3018 2396 3024 2397
rect 2710 2392 2711 2396
rect 2715 2392 3019 2396
rect 3023 2392 3024 2396
rect 2710 2391 2716 2392
rect 3018 2391 3024 2392
rect 1134 2388 1140 2389
rect 1338 2388 1344 2389
rect 1134 2384 1135 2388
rect 1139 2384 1339 2388
rect 1343 2384 1344 2388
rect 1134 2383 1140 2384
rect 1338 2383 1344 2384
rect 2662 2380 2668 2381
rect 2966 2380 2972 2381
rect 84 2373 85 2379
rect 91 2378 1835 2379
rect 91 2374 111 2378
rect 115 2374 159 2378
rect 163 2374 183 2378
rect 187 2374 247 2378
rect 251 2374 311 2378
rect 315 2374 335 2378
rect 339 2374 439 2378
rect 443 2374 447 2378
rect 451 2374 559 2378
rect 563 2374 583 2378
rect 587 2374 687 2378
rect 691 2374 719 2378
rect 723 2374 815 2378
rect 819 2374 855 2378
rect 859 2374 951 2378
rect 955 2374 991 2378
rect 995 2374 1079 2378
rect 1083 2374 1127 2378
rect 1131 2374 1207 2378
rect 1211 2374 1263 2378
rect 1267 2374 1327 2378
rect 1331 2374 1399 2378
rect 1403 2374 1455 2378
rect 1459 2374 1583 2378
rect 1587 2374 1823 2378
rect 1827 2374 1835 2378
rect 91 2373 1835 2374
rect 1841 2373 1842 2379
rect 2662 2376 2663 2380
rect 2667 2376 2967 2380
rect 2971 2376 2972 2380
rect 2662 2375 2668 2376
rect 2966 2375 2972 2376
rect 1846 2361 1847 2367
rect 1853 2366 3611 2367
rect 1853 2362 1863 2366
rect 1867 2362 1895 2366
rect 1899 2362 1927 2366
rect 1931 2362 2023 2366
rect 2027 2362 2087 2366
rect 2091 2362 2183 2366
rect 2187 2362 2247 2366
rect 2251 2362 2343 2366
rect 2347 2362 2407 2366
rect 2411 2362 2503 2366
rect 2507 2362 2559 2366
rect 2563 2362 2655 2366
rect 2659 2362 2703 2366
rect 2707 2362 2807 2366
rect 2811 2362 2831 2366
rect 2835 2362 2951 2366
rect 2955 2362 2959 2366
rect 2963 2362 3071 2366
rect 3075 2362 3119 2366
rect 3123 2362 3183 2366
rect 3187 2362 3287 2366
rect 3291 2362 3399 2366
rect 3403 2362 3487 2366
rect 3491 2362 3575 2366
rect 3579 2362 3611 2366
rect 1853 2361 3611 2362
rect 3617 2361 3618 2367
rect 1182 2316 1188 2317
rect 1522 2316 1528 2317
rect 1182 2312 1183 2316
rect 1187 2312 1523 2316
rect 1527 2312 1528 2316
rect 1182 2311 1188 2312
rect 1522 2311 1528 2312
rect 1834 2307 1835 2313
rect 1841 2307 1866 2313
rect 96 2297 97 2303
rect 103 2302 1847 2303
rect 103 2298 111 2302
rect 115 2298 167 2302
rect 171 2298 255 2302
rect 259 2298 343 2302
rect 347 2298 447 2302
rect 451 2298 567 2302
rect 571 2298 695 2302
rect 699 2298 823 2302
rect 827 2298 863 2302
rect 867 2298 959 2302
rect 963 2298 1023 2302
rect 1027 2298 1087 2302
rect 1091 2298 1175 2302
rect 1179 2298 1215 2302
rect 1219 2298 1319 2302
rect 1323 2298 1335 2302
rect 1339 2298 1463 2302
rect 1467 2298 1591 2302
rect 1595 2298 1599 2302
rect 1603 2298 1735 2302
rect 1739 2298 1823 2302
rect 1827 2298 1847 2302
rect 103 2297 1847 2298
rect 1853 2297 1854 2303
rect 1860 2295 1866 2307
rect 1860 2294 3599 2295
rect 702 2292 708 2293
rect 938 2292 944 2293
rect 702 2288 703 2292
rect 707 2288 939 2292
rect 943 2288 944 2292
rect 1860 2290 1863 2294
rect 1867 2290 1919 2294
rect 1923 2290 1975 2294
rect 1979 2290 2079 2294
rect 2083 2290 2143 2294
rect 2147 2290 2239 2294
rect 2243 2290 2311 2294
rect 2315 2290 2399 2294
rect 2403 2290 2479 2294
rect 2483 2290 2551 2294
rect 2555 2290 2639 2294
rect 2643 2290 2695 2294
rect 2699 2290 2783 2294
rect 2787 2290 2823 2294
rect 2827 2290 2919 2294
rect 2923 2290 2943 2294
rect 2947 2290 3039 2294
rect 3043 2290 3063 2294
rect 3067 2290 3159 2294
rect 3163 2290 3175 2294
rect 3179 2290 3271 2294
rect 3275 2290 3279 2294
rect 3283 2290 3383 2294
rect 3387 2290 3391 2294
rect 3395 2290 3479 2294
rect 3483 2290 3575 2294
rect 3579 2290 3599 2294
rect 1860 2289 3599 2290
rect 3605 2289 3606 2295
rect 702 2287 708 2288
rect 938 2287 944 2288
rect 2798 2236 2804 2237
rect 3182 2236 3188 2237
rect 2798 2232 2799 2236
rect 2803 2232 3183 2236
rect 3187 2232 3188 2236
rect 2798 2231 2804 2232
rect 3182 2231 3188 2232
rect 84 2221 85 2227
rect 91 2226 1835 2227
rect 91 2222 111 2226
rect 115 2222 535 2226
rect 539 2222 687 2226
rect 691 2222 719 2226
rect 723 2222 855 2226
rect 859 2222 895 2226
rect 899 2222 1015 2226
rect 1019 2222 1071 2226
rect 1075 2222 1167 2226
rect 1171 2222 1239 2226
rect 1243 2222 1311 2226
rect 1315 2222 1407 2226
rect 1411 2222 1455 2226
rect 1459 2222 1575 2226
rect 1579 2222 1591 2226
rect 1595 2222 1727 2226
rect 1731 2222 1823 2226
rect 1827 2222 1835 2226
rect 91 2221 1835 2222
rect 1841 2221 1842 2227
rect 1846 2221 1847 2227
rect 1853 2226 3611 2227
rect 1853 2222 1863 2226
rect 1867 2222 1983 2226
rect 1987 2222 2007 2226
rect 2011 2222 2151 2226
rect 2155 2222 2167 2226
rect 2171 2222 2319 2226
rect 2323 2222 2335 2226
rect 2339 2222 2487 2226
rect 2491 2222 2519 2226
rect 2523 2222 2647 2226
rect 2651 2222 2711 2226
rect 2715 2222 2791 2226
rect 2795 2222 2903 2226
rect 2907 2222 2927 2226
rect 2931 2222 3047 2226
rect 3051 2222 3103 2226
rect 3107 2222 3167 2226
rect 3171 2222 3279 2226
rect 3283 2222 3303 2226
rect 3307 2222 3391 2226
rect 3395 2222 3487 2226
rect 3491 2222 3575 2226
rect 3579 2222 3611 2226
rect 1853 2221 3611 2222
rect 3617 2221 3618 2227
rect 1254 2180 1260 2181
rect 1666 2180 1672 2181
rect 1254 2176 1255 2180
rect 1259 2176 1667 2180
rect 1671 2176 1672 2180
rect 1254 2175 1260 2176
rect 1666 2175 1672 2176
rect 1834 2163 1835 2169
rect 1841 2163 1866 2169
rect 96 2153 97 2159
rect 103 2158 1847 2159
rect 103 2154 111 2158
rect 115 2154 495 2158
rect 499 2154 543 2158
rect 547 2154 623 2158
rect 627 2154 727 2158
rect 731 2154 759 2158
rect 763 2154 895 2158
rect 899 2154 903 2158
rect 907 2154 1039 2158
rect 1043 2154 1079 2158
rect 1083 2154 1183 2158
rect 1187 2154 1247 2158
rect 1251 2154 1327 2158
rect 1331 2154 1415 2158
rect 1419 2154 1471 2158
rect 1475 2154 1583 2158
rect 1587 2154 1623 2158
rect 1627 2154 1735 2158
rect 1739 2154 1823 2158
rect 1827 2154 1847 2158
rect 103 2153 1847 2154
rect 1853 2153 1854 2159
rect 1860 2151 1866 2163
rect 1860 2150 3599 2151
rect 550 2148 556 2149
rect 766 2148 772 2149
rect 550 2144 551 2148
rect 555 2144 767 2148
rect 771 2144 772 2148
rect 1860 2146 1863 2150
rect 1867 2146 1999 2150
rect 2003 2146 2023 2150
rect 2027 2146 2159 2150
rect 2163 2146 2167 2150
rect 2171 2146 2319 2150
rect 2323 2146 2327 2150
rect 2331 2146 2471 2150
rect 2475 2146 2511 2150
rect 2515 2146 2615 2150
rect 2619 2146 2703 2150
rect 2707 2146 2759 2150
rect 2763 2146 2895 2150
rect 2899 2146 3023 2150
rect 3027 2146 3095 2150
rect 3099 2146 3143 2150
rect 3147 2146 3263 2150
rect 3267 2146 3295 2150
rect 3299 2146 3383 2150
rect 3387 2146 3479 2150
rect 3483 2146 3575 2150
rect 3579 2146 3599 2150
rect 1860 2145 3599 2146
rect 3605 2145 3606 2151
rect 550 2143 556 2144
rect 766 2143 772 2144
rect 574 2111 575 2117
rect 581 2111 582 2117
rect 1038 2103 1039 2109
rect 1045 2103 1046 2109
rect 84 2081 85 2087
rect 91 2086 1835 2087
rect 91 2082 111 2086
rect 115 2082 319 2086
rect 323 2082 431 2086
rect 435 2082 487 2086
rect 491 2082 551 2086
rect 555 2082 615 2086
rect 619 2082 679 2086
rect 683 2082 751 2086
rect 755 2082 799 2086
rect 803 2082 887 2086
rect 891 2082 919 2086
rect 923 2082 1031 2086
rect 1035 2082 1039 2086
rect 1043 2082 1159 2086
rect 1163 2082 1175 2086
rect 1179 2082 1279 2086
rect 1283 2082 1319 2086
rect 1323 2082 1407 2086
rect 1411 2082 1463 2086
rect 1467 2082 1615 2086
rect 1619 2082 1823 2086
rect 1827 2082 1835 2086
rect 91 2081 1835 2082
rect 1841 2081 1842 2087
rect 1846 2073 1847 2079
rect 1853 2078 3611 2079
rect 1853 2074 1863 2078
rect 1867 2074 1983 2078
rect 1987 2074 2031 2078
rect 2035 2074 2143 2078
rect 2147 2074 2175 2078
rect 2179 2074 2311 2078
rect 2315 2074 2327 2078
rect 2331 2074 2471 2078
rect 2475 2074 2479 2078
rect 2483 2074 2623 2078
rect 2627 2074 2631 2078
rect 2635 2074 2767 2078
rect 2771 2074 2775 2078
rect 2779 2074 2903 2078
rect 2907 2074 2911 2078
rect 2915 2074 3031 2078
rect 3035 2074 3039 2078
rect 3043 2074 3151 2078
rect 3155 2074 3159 2078
rect 3163 2074 3271 2078
rect 3275 2074 3279 2078
rect 3283 2074 3391 2078
rect 3395 2074 3487 2078
rect 3491 2074 3575 2078
rect 3579 2074 3611 2078
rect 1853 2073 3611 2074
rect 3617 2073 3618 2079
rect 1834 2019 1835 2025
rect 1841 2019 1866 2025
rect 96 2009 97 2015
rect 103 2014 1847 2015
rect 103 2010 111 2014
rect 115 2010 183 2014
rect 187 2010 295 2014
rect 299 2010 327 2014
rect 331 2010 415 2014
rect 419 2010 439 2014
rect 443 2010 535 2014
rect 539 2010 559 2014
rect 563 2010 655 2014
rect 659 2010 687 2014
rect 691 2010 775 2014
rect 779 2010 807 2014
rect 811 2010 895 2014
rect 899 2010 927 2014
rect 931 2010 1015 2014
rect 1019 2010 1047 2014
rect 1051 2010 1135 2014
rect 1139 2010 1167 2014
rect 1171 2010 1255 2014
rect 1259 2010 1287 2014
rect 1291 2010 1415 2014
rect 1419 2010 1823 2014
rect 1827 2010 1847 2014
rect 103 2009 1847 2010
rect 1853 2009 1854 2015
rect 1860 2011 1866 2019
rect 1860 2010 3599 2011
rect 1860 2006 1863 2010
rect 1867 2006 1887 2010
rect 1891 2006 1975 2010
rect 1979 2006 2031 2010
rect 2035 2006 2135 2010
rect 2139 2006 2199 2010
rect 2203 2006 2303 2010
rect 2307 2006 2375 2010
rect 2379 2006 2463 2010
rect 2467 2006 2543 2010
rect 2547 2006 2623 2010
rect 2627 2006 2711 2010
rect 2715 2006 2767 2010
rect 2771 2006 2871 2010
rect 2875 2006 2903 2010
rect 2907 2006 3031 2010
rect 3035 2006 3039 2010
rect 3043 2006 3151 2010
rect 3155 2006 3207 2010
rect 3211 2006 3271 2010
rect 3275 2006 3383 2010
rect 3387 2006 3479 2010
rect 3483 2006 3575 2010
rect 3579 2006 3599 2010
rect 1860 2005 3599 2006
rect 3605 2005 3606 2011
rect 238 1964 244 1965
rect 562 1964 568 1965
rect 238 1960 239 1964
rect 243 1960 563 1964
rect 567 1960 568 1964
rect 238 1959 244 1960
rect 562 1959 568 1960
rect 2726 1956 2732 1957
rect 3158 1956 3164 1957
rect 2726 1952 2727 1956
rect 2731 1952 3159 1956
rect 3163 1952 3164 1956
rect 2726 1951 2732 1952
rect 3158 1951 3164 1952
rect 84 1937 85 1943
rect 91 1942 1835 1943
rect 91 1938 111 1942
rect 115 1938 135 1942
rect 139 1938 175 1942
rect 179 1938 223 1942
rect 227 1938 287 1942
rect 291 1938 351 1942
rect 355 1938 407 1942
rect 411 1938 495 1942
rect 499 1938 527 1942
rect 531 1938 647 1942
rect 651 1938 655 1942
rect 659 1938 767 1942
rect 771 1938 839 1942
rect 843 1938 887 1942
rect 891 1938 1007 1942
rect 1011 1938 1039 1942
rect 1043 1938 1127 1942
rect 1131 1938 1247 1942
rect 1251 1938 1463 1942
rect 1467 1938 1823 1942
rect 1827 1938 1835 1942
rect 91 1937 1835 1938
rect 1841 1937 1842 1943
rect 1846 1929 1847 1935
rect 1853 1934 3611 1935
rect 1853 1930 1863 1934
rect 1867 1930 1895 1934
rect 1899 1930 1991 1934
rect 1995 1930 2039 1934
rect 2043 1930 2119 1934
rect 2123 1930 2207 1934
rect 2211 1930 2255 1934
rect 2259 1930 2383 1934
rect 2387 1930 2511 1934
rect 2515 1930 2551 1934
rect 2555 1930 2631 1934
rect 2635 1930 2719 1934
rect 2723 1930 2751 1934
rect 2755 1930 2879 1934
rect 2883 1930 3007 1934
rect 3011 1930 3047 1934
rect 3051 1930 3215 1934
rect 3219 1930 3575 1934
rect 3579 1930 3611 1934
rect 1853 1929 3611 1930
rect 3617 1929 3618 1935
rect 950 1884 956 1885
rect 1158 1884 1164 1885
rect 950 1880 951 1884
rect 955 1880 1159 1884
rect 1163 1880 1164 1884
rect 950 1879 956 1880
rect 1158 1879 1164 1880
rect 1834 1871 1835 1877
rect 1841 1871 1866 1877
rect 96 1861 97 1867
rect 103 1866 1847 1867
rect 103 1862 111 1866
rect 115 1862 143 1866
rect 147 1862 231 1866
rect 235 1862 271 1866
rect 275 1862 359 1866
rect 363 1862 415 1866
rect 419 1862 503 1866
rect 507 1862 559 1866
rect 563 1862 663 1866
rect 667 1862 695 1866
rect 699 1862 823 1866
rect 827 1862 847 1866
rect 851 1862 943 1866
rect 947 1862 1047 1866
rect 1051 1862 1055 1866
rect 1059 1862 1159 1866
rect 1163 1862 1255 1866
rect 1259 1862 1263 1866
rect 1267 1862 1359 1866
rect 1363 1862 1455 1866
rect 1459 1862 1471 1866
rect 1475 1862 1551 1866
rect 1555 1862 1647 1866
rect 1651 1862 1735 1866
rect 1739 1862 1823 1866
rect 1827 1862 1847 1866
rect 103 1861 1847 1862
rect 1853 1861 1854 1867
rect 1860 1859 1866 1871
rect 1860 1858 3599 1859
rect 1860 1854 1863 1858
rect 1867 1854 1887 1858
rect 1891 1854 1983 1858
rect 1987 1854 2111 1858
rect 2115 1854 2223 1858
rect 2227 1854 2247 1858
rect 2251 1854 2359 1858
rect 2363 1854 2375 1858
rect 2379 1854 2495 1858
rect 2499 1854 2503 1858
rect 2507 1854 2623 1858
rect 2627 1854 2743 1858
rect 2747 1854 2863 1858
rect 2867 1854 2871 1858
rect 2875 1854 2991 1858
rect 2995 1854 2999 1858
rect 3003 1854 3575 1858
rect 3579 1854 3599 1858
rect 1860 1853 3599 1854
rect 3605 1853 3606 1859
rect 84 1781 85 1787
rect 91 1786 1835 1787
rect 91 1782 111 1786
rect 115 1782 135 1786
rect 139 1782 263 1786
rect 267 1782 303 1786
rect 307 1782 407 1786
rect 411 1782 495 1786
rect 499 1782 551 1786
rect 555 1782 687 1786
rect 691 1782 815 1786
rect 819 1782 871 1786
rect 875 1782 935 1786
rect 939 1782 1047 1786
rect 1051 1782 1151 1786
rect 1155 1782 1215 1786
rect 1219 1782 1255 1786
rect 1259 1782 1351 1786
rect 1355 1782 1375 1786
rect 1379 1782 1447 1786
rect 1451 1782 1535 1786
rect 1539 1782 1543 1786
rect 1547 1782 1639 1786
rect 1643 1782 1703 1786
rect 1707 1782 1727 1786
rect 1731 1782 1823 1786
rect 1827 1782 1835 1786
rect 91 1781 1835 1782
rect 1841 1781 1842 1787
rect 1846 1781 1847 1787
rect 1853 1786 3611 1787
rect 1853 1782 1863 1786
rect 1867 1782 2231 1786
rect 2235 1782 2271 1786
rect 2275 1782 2359 1786
rect 2363 1782 2367 1786
rect 2371 1782 2455 1786
rect 2459 1782 2503 1786
rect 2507 1782 2559 1786
rect 2563 1782 2631 1786
rect 2635 1782 2663 1786
rect 2667 1782 2751 1786
rect 2755 1782 2759 1786
rect 2763 1782 2863 1786
rect 2867 1782 2871 1786
rect 2875 1782 2967 1786
rect 2971 1782 2999 1786
rect 3003 1782 3071 1786
rect 3075 1782 3175 1786
rect 3179 1782 3575 1786
rect 3579 1782 3611 1786
rect 1853 1781 3611 1782
rect 3617 1781 3618 1787
rect 1834 1719 1835 1725
rect 1841 1719 1866 1725
rect 1860 1715 1866 1719
rect 96 1709 97 1715
rect 103 1714 1847 1715
rect 103 1710 111 1714
rect 115 1710 143 1714
rect 147 1710 287 1714
rect 291 1710 311 1714
rect 315 1710 471 1714
rect 475 1710 503 1714
rect 507 1710 655 1714
rect 659 1710 695 1714
rect 699 1710 839 1714
rect 843 1710 879 1714
rect 883 1710 1023 1714
rect 1027 1710 1055 1714
rect 1059 1710 1191 1714
rect 1195 1710 1223 1714
rect 1227 1710 1359 1714
rect 1363 1710 1383 1714
rect 1387 1710 1527 1714
rect 1531 1710 1543 1714
rect 1547 1710 1695 1714
rect 1699 1710 1711 1714
rect 1715 1710 1823 1714
rect 1827 1710 1847 1714
rect 103 1709 1847 1710
rect 1853 1709 1854 1715
rect 1860 1714 3599 1715
rect 1860 1710 1863 1714
rect 1867 1710 2247 1714
rect 2251 1710 2263 1714
rect 2267 1710 2351 1714
rect 2355 1710 2367 1714
rect 2371 1710 2447 1714
rect 2451 1710 2495 1714
rect 2499 1710 2551 1714
rect 2555 1710 2623 1714
rect 2627 1710 2655 1714
rect 2659 1710 2751 1714
rect 2755 1710 2759 1714
rect 2763 1710 2855 1714
rect 2859 1710 2887 1714
rect 2891 1710 2959 1714
rect 2963 1710 3015 1714
rect 3019 1710 3063 1714
rect 3067 1710 3135 1714
rect 3139 1710 3167 1714
rect 3171 1710 3247 1714
rect 3251 1710 3367 1714
rect 3371 1710 3479 1714
rect 3483 1710 3575 1714
rect 3579 1710 3599 1714
rect 1860 1709 3599 1710
rect 3605 1709 3606 1715
rect 84 1633 85 1639
rect 91 1638 1835 1639
rect 91 1634 111 1638
rect 115 1634 135 1638
rect 139 1634 271 1638
rect 275 1634 279 1638
rect 283 1634 447 1638
rect 451 1634 463 1638
rect 467 1634 631 1638
rect 635 1634 647 1638
rect 651 1634 815 1638
rect 819 1634 831 1638
rect 835 1634 991 1638
rect 995 1634 1015 1638
rect 1019 1634 1151 1638
rect 1155 1634 1183 1638
rect 1187 1634 1303 1638
rect 1307 1634 1351 1638
rect 1355 1634 1455 1638
rect 1459 1634 1519 1638
rect 1523 1634 1599 1638
rect 1603 1634 1687 1638
rect 1691 1634 1727 1638
rect 1731 1634 1823 1638
rect 1827 1634 1835 1638
rect 91 1633 1835 1634
rect 1841 1633 1842 1639
rect 1846 1637 1847 1643
rect 1853 1642 3611 1643
rect 1853 1638 1863 1642
rect 1867 1638 2151 1642
rect 2155 1638 2255 1642
rect 2259 1638 2343 1642
rect 2347 1638 2375 1642
rect 2379 1638 2503 1642
rect 2507 1638 2527 1642
rect 2531 1638 2631 1642
rect 2635 1638 2703 1642
rect 2707 1638 2767 1642
rect 2771 1638 2871 1642
rect 2875 1638 2895 1642
rect 2899 1638 3023 1642
rect 3027 1638 3031 1642
rect 3035 1638 3143 1642
rect 3147 1638 3191 1642
rect 3195 1638 3255 1642
rect 3259 1638 3351 1642
rect 3355 1638 3375 1642
rect 3379 1638 3487 1642
rect 3491 1638 3575 1642
rect 3579 1638 3611 1642
rect 1853 1637 3611 1638
rect 3617 1637 3618 1643
rect 1834 1575 1835 1581
rect 1841 1575 1866 1581
rect 1860 1574 3599 1575
rect 96 1565 97 1571
rect 103 1570 1847 1571
rect 103 1566 111 1570
rect 115 1566 143 1570
rect 147 1566 271 1570
rect 275 1566 279 1570
rect 283 1566 431 1570
rect 435 1566 455 1570
rect 459 1566 599 1570
rect 603 1566 639 1570
rect 643 1566 767 1570
rect 771 1566 823 1570
rect 827 1566 935 1570
rect 939 1566 999 1570
rect 1003 1566 1103 1570
rect 1107 1566 1159 1570
rect 1163 1566 1263 1570
rect 1267 1566 1311 1570
rect 1315 1566 1423 1570
rect 1427 1566 1463 1570
rect 1467 1566 1591 1570
rect 1595 1566 1607 1570
rect 1611 1566 1735 1570
rect 1739 1566 1823 1570
rect 1827 1566 1847 1570
rect 103 1565 1847 1566
rect 1853 1565 1854 1571
rect 1860 1570 1863 1574
rect 1867 1570 2087 1574
rect 2091 1570 2143 1574
rect 2147 1570 2279 1574
rect 2283 1570 2335 1574
rect 2339 1570 2455 1574
rect 2459 1570 2519 1574
rect 2523 1570 2623 1574
rect 2627 1570 2695 1574
rect 2699 1570 2791 1574
rect 2795 1570 2863 1574
rect 2867 1570 2951 1574
rect 2955 1570 3023 1574
rect 3027 1570 3111 1574
rect 3115 1570 3183 1574
rect 3187 1570 3271 1574
rect 3275 1570 3343 1574
rect 3347 1570 3431 1574
rect 3435 1570 3479 1574
rect 3483 1570 3575 1574
rect 3579 1570 3599 1574
rect 1860 1569 3599 1570
rect 3605 1569 3606 1575
rect 2638 1516 2644 1517
rect 3214 1516 3220 1517
rect 2638 1512 2639 1516
rect 2643 1512 3215 1516
rect 3219 1512 3220 1516
rect 2638 1511 2644 1512
rect 3214 1511 3220 1512
rect 84 1493 85 1499
rect 91 1498 1835 1499
rect 91 1494 111 1498
rect 115 1494 135 1498
rect 139 1494 183 1498
rect 187 1494 263 1498
rect 267 1494 327 1498
rect 331 1494 423 1498
rect 427 1494 471 1498
rect 475 1494 591 1498
rect 595 1494 607 1498
rect 611 1494 743 1498
rect 747 1494 759 1498
rect 763 1494 871 1498
rect 875 1494 927 1498
rect 931 1494 991 1498
rect 995 1494 1095 1498
rect 1099 1494 1119 1498
rect 1123 1494 1247 1498
rect 1251 1494 1255 1498
rect 1259 1494 1375 1498
rect 1379 1494 1415 1498
rect 1419 1494 1583 1498
rect 1587 1494 1727 1498
rect 1731 1494 1823 1498
rect 1827 1494 1835 1498
rect 91 1493 1835 1494
rect 1841 1493 1842 1499
rect 1846 1493 1847 1499
rect 1853 1498 3611 1499
rect 1853 1494 1863 1498
rect 1867 1494 1895 1498
rect 1899 1494 1991 1498
rect 1995 1494 2095 1498
rect 2099 1494 2119 1498
rect 2123 1494 2247 1498
rect 2251 1494 2287 1498
rect 2291 1494 2383 1498
rect 2387 1494 2463 1498
rect 2467 1494 2535 1498
rect 2539 1494 2631 1498
rect 2635 1494 2703 1498
rect 2707 1494 2799 1498
rect 2803 1494 2887 1498
rect 2891 1494 2959 1498
rect 2963 1494 3087 1498
rect 3091 1494 3119 1498
rect 3123 1494 3279 1498
rect 3283 1494 3295 1498
rect 3299 1494 3439 1498
rect 3443 1494 3487 1498
rect 3491 1494 3575 1498
rect 3579 1494 3611 1498
rect 1853 1493 3611 1494
rect 3617 1493 3618 1499
rect 1834 1427 1835 1433
rect 1841 1427 1866 1433
rect 1860 1426 3599 1427
rect 96 1417 97 1423
rect 103 1422 1847 1423
rect 103 1418 111 1422
rect 115 1418 191 1422
rect 195 1418 199 1422
rect 203 1418 335 1422
rect 339 1418 463 1422
rect 467 1418 479 1422
rect 483 1418 583 1422
rect 587 1418 615 1422
rect 619 1418 703 1422
rect 707 1418 751 1422
rect 755 1418 815 1422
rect 819 1418 879 1422
rect 883 1418 919 1422
rect 923 1418 999 1422
rect 1003 1418 1015 1422
rect 1019 1418 1119 1422
rect 1123 1418 1127 1422
rect 1131 1418 1223 1422
rect 1227 1418 1255 1422
rect 1259 1418 1327 1422
rect 1331 1418 1383 1422
rect 1387 1418 1823 1422
rect 1827 1418 1847 1422
rect 103 1417 1847 1418
rect 1853 1417 1854 1423
rect 1860 1422 1863 1426
rect 1867 1422 1887 1426
rect 1891 1422 1975 1426
rect 1979 1422 1983 1426
rect 1987 1422 2071 1426
rect 2075 1422 2111 1426
rect 2115 1422 2183 1426
rect 2187 1422 2239 1426
rect 2243 1422 2303 1426
rect 2307 1422 2375 1426
rect 2379 1422 2439 1426
rect 2443 1422 2527 1426
rect 2531 1422 2607 1426
rect 2611 1422 2695 1426
rect 2699 1422 2807 1426
rect 2811 1422 2879 1426
rect 2883 1422 3031 1426
rect 3035 1422 3079 1426
rect 3083 1422 3263 1426
rect 3267 1422 3287 1426
rect 3291 1422 3479 1426
rect 3483 1422 3575 1426
rect 3579 1422 3599 1426
rect 1860 1421 3599 1422
rect 3605 1421 3606 1427
rect 2774 1364 2780 1365
rect 3210 1364 3216 1365
rect 2774 1360 2775 1364
rect 2779 1360 3211 1364
rect 3215 1360 3216 1364
rect 2774 1359 2780 1360
rect 3210 1359 3216 1360
rect 84 1345 85 1351
rect 91 1350 1835 1351
rect 91 1346 111 1350
rect 115 1346 191 1350
rect 195 1346 231 1350
rect 235 1346 327 1350
rect 331 1346 383 1350
rect 387 1346 455 1350
rect 459 1346 543 1350
rect 547 1346 575 1350
rect 579 1346 695 1350
rect 699 1346 703 1350
rect 707 1346 807 1350
rect 811 1346 871 1350
rect 875 1346 911 1350
rect 915 1346 1007 1350
rect 1011 1346 1039 1350
rect 1043 1346 1111 1350
rect 1115 1346 1207 1350
rect 1211 1346 1215 1350
rect 1219 1346 1319 1350
rect 1323 1346 1375 1350
rect 1379 1346 1823 1350
rect 1827 1346 1835 1350
rect 91 1345 1835 1346
rect 1841 1345 1842 1351
rect 1846 1349 1847 1355
rect 1853 1354 3611 1355
rect 1853 1350 1863 1354
rect 1867 1350 1895 1354
rect 1899 1350 1983 1354
rect 1987 1350 2079 1354
rect 2083 1350 2103 1354
rect 2107 1350 2191 1354
rect 2195 1350 2223 1354
rect 2227 1350 2311 1354
rect 2315 1350 2359 1354
rect 2363 1350 2447 1354
rect 2451 1350 2511 1354
rect 2515 1350 2615 1354
rect 2619 1350 2687 1354
rect 2691 1350 2815 1354
rect 2819 1350 2871 1354
rect 2875 1350 3039 1354
rect 3043 1350 3071 1354
rect 3075 1350 3271 1354
rect 3275 1350 3279 1354
rect 3283 1350 3487 1354
rect 3491 1350 3575 1354
rect 3579 1350 3611 1354
rect 1853 1349 3611 1350
rect 3617 1349 3618 1355
rect 558 1292 564 1293
rect 798 1292 804 1293
rect 558 1288 559 1292
rect 563 1288 799 1292
rect 803 1288 804 1292
rect 558 1287 564 1288
rect 798 1287 804 1288
rect 1834 1287 1835 1293
rect 1841 1287 1866 1293
rect 96 1277 97 1283
rect 103 1282 1847 1283
rect 103 1278 111 1282
rect 115 1278 215 1282
rect 219 1278 239 1282
rect 243 1278 359 1282
rect 363 1278 391 1282
rect 395 1278 519 1282
rect 523 1278 551 1282
rect 555 1278 679 1282
rect 683 1278 711 1282
rect 715 1278 839 1282
rect 843 1278 879 1282
rect 883 1278 999 1282
rect 1003 1278 1047 1282
rect 1051 1278 1151 1282
rect 1155 1278 1215 1282
rect 1219 1278 1295 1282
rect 1299 1278 1383 1282
rect 1387 1278 1439 1282
rect 1443 1278 1591 1282
rect 1595 1278 1823 1282
rect 1827 1278 1847 1282
rect 103 1277 1847 1278
rect 1853 1277 1854 1283
rect 1860 1275 1866 1287
rect 1860 1274 3599 1275
rect 1860 1270 1863 1274
rect 1867 1270 1887 1274
rect 1891 1270 1975 1274
rect 1979 1270 2055 1274
rect 2059 1270 2095 1274
rect 2099 1270 2143 1274
rect 2147 1270 2215 1274
rect 2219 1270 2239 1274
rect 2243 1270 2335 1274
rect 2339 1270 2351 1274
rect 2355 1270 2431 1274
rect 2435 1270 2503 1274
rect 2507 1270 2551 1274
rect 2555 1270 2679 1274
rect 2683 1270 2687 1274
rect 2691 1270 2855 1274
rect 2859 1270 2863 1274
rect 2867 1270 3039 1274
rect 3043 1270 3063 1274
rect 3067 1270 3231 1274
rect 3235 1270 3271 1274
rect 3275 1270 3431 1274
rect 3435 1270 3479 1274
rect 3483 1270 3575 1274
rect 3579 1270 3599 1274
rect 1860 1269 3599 1270
rect 3605 1269 3606 1275
rect 2566 1260 2572 1261
rect 2958 1260 2964 1261
rect 2566 1256 2567 1260
rect 2571 1256 2959 1260
rect 2963 1256 2964 1260
rect 2566 1255 2572 1256
rect 2958 1255 2964 1256
rect 84 1201 85 1207
rect 91 1206 1835 1207
rect 91 1202 111 1206
rect 115 1202 135 1206
rect 139 1202 207 1206
rect 211 1202 271 1206
rect 275 1202 351 1206
rect 355 1202 423 1206
rect 427 1202 511 1206
rect 515 1202 575 1206
rect 579 1202 671 1206
rect 675 1202 727 1206
rect 731 1202 831 1206
rect 835 1202 887 1206
rect 891 1202 991 1206
rect 995 1202 1055 1206
rect 1059 1202 1143 1206
rect 1147 1202 1231 1206
rect 1235 1202 1287 1206
rect 1291 1202 1415 1206
rect 1419 1202 1431 1206
rect 1435 1202 1583 1206
rect 1587 1202 1599 1206
rect 1603 1202 1823 1206
rect 1827 1202 1835 1206
rect 91 1201 1835 1202
rect 1841 1201 1842 1207
rect 1846 1197 1847 1203
rect 1853 1202 3611 1203
rect 1853 1198 1863 1202
rect 1867 1198 2039 1202
rect 2043 1198 2063 1202
rect 2067 1198 2151 1202
rect 2155 1198 2247 1202
rect 2251 1198 2279 1202
rect 2283 1198 2343 1202
rect 2347 1198 2415 1202
rect 2419 1198 2439 1202
rect 2443 1198 2559 1202
rect 2563 1198 2695 1202
rect 2699 1198 2711 1202
rect 2715 1198 2863 1202
rect 2867 1198 3015 1202
rect 3019 1198 3047 1202
rect 3051 1198 3167 1202
rect 3171 1198 3239 1202
rect 3243 1198 3327 1202
rect 3331 1198 3439 1202
rect 3443 1198 3487 1202
rect 3491 1198 3575 1202
rect 3579 1198 3611 1202
rect 1853 1197 3611 1198
rect 3617 1197 3618 1203
rect 96 1133 97 1139
rect 103 1138 1847 1139
rect 103 1134 111 1138
rect 115 1134 143 1138
rect 147 1134 279 1138
rect 283 1134 295 1138
rect 299 1134 431 1138
rect 435 1134 479 1138
rect 483 1134 583 1138
rect 587 1134 663 1138
rect 667 1134 735 1138
rect 739 1134 847 1138
rect 851 1134 895 1138
rect 899 1134 1031 1138
rect 1035 1134 1063 1138
rect 1067 1134 1207 1138
rect 1211 1134 1239 1138
rect 1243 1134 1391 1138
rect 1395 1134 1423 1138
rect 1427 1134 1575 1138
rect 1579 1134 1607 1138
rect 1611 1134 1735 1138
rect 1739 1134 1823 1138
rect 1827 1134 1847 1138
rect 103 1133 1847 1134
rect 1853 1133 1854 1139
rect 1834 1117 1835 1123
rect 1841 1122 3599 1123
rect 1841 1118 1863 1122
rect 1867 1118 1943 1122
rect 1947 1118 2031 1122
rect 2035 1118 2087 1122
rect 2091 1118 2143 1122
rect 2147 1118 2231 1122
rect 2235 1118 2271 1122
rect 2275 1118 2383 1122
rect 2387 1118 2407 1122
rect 2411 1118 2535 1122
rect 2539 1118 2551 1122
rect 2555 1118 2687 1122
rect 2691 1118 2703 1122
rect 2707 1118 2839 1122
rect 2843 1118 2855 1122
rect 2859 1118 2991 1122
rect 2995 1118 3007 1122
rect 3011 1118 3151 1122
rect 3155 1118 3159 1122
rect 3163 1118 3319 1122
rect 3323 1118 3479 1122
rect 3483 1118 3575 1122
rect 3579 1118 3599 1122
rect 1841 1117 3599 1118
rect 3605 1117 3606 1123
rect 84 1065 85 1071
rect 91 1070 1835 1071
rect 91 1066 111 1070
rect 115 1066 135 1070
rect 139 1066 271 1070
rect 275 1066 287 1070
rect 291 1066 431 1070
rect 435 1066 471 1070
rect 475 1066 583 1070
rect 587 1066 655 1070
rect 659 1066 735 1070
rect 739 1066 839 1070
rect 843 1066 887 1070
rect 891 1066 1023 1070
rect 1027 1066 1047 1070
rect 1051 1066 1199 1070
rect 1203 1066 1215 1070
rect 1219 1066 1383 1070
rect 1387 1066 1559 1070
rect 1563 1066 1567 1070
rect 1571 1066 1727 1070
rect 1731 1066 1823 1070
rect 1827 1066 1835 1070
rect 91 1065 1835 1066
rect 1841 1065 1842 1071
rect 2702 1052 2708 1053
rect 3078 1052 3084 1053
rect 2702 1048 2703 1052
rect 2707 1048 3079 1052
rect 3083 1048 3084 1052
rect 2702 1047 2708 1048
rect 3078 1047 3084 1048
rect 1846 1037 1847 1043
rect 1853 1042 3611 1043
rect 1853 1038 1863 1042
rect 1867 1038 1919 1042
rect 1923 1038 1951 1042
rect 1955 1038 2095 1042
rect 2099 1038 2127 1042
rect 2131 1038 2239 1042
rect 2243 1038 2327 1042
rect 2331 1038 2391 1042
rect 2395 1038 2519 1042
rect 2523 1038 2543 1042
rect 2547 1038 2695 1042
rect 2699 1038 2847 1042
rect 2851 1038 2863 1042
rect 2867 1038 2999 1042
rect 3003 1038 3023 1042
rect 3027 1038 3159 1042
rect 3163 1038 3183 1042
rect 3187 1038 3327 1042
rect 3331 1038 3343 1042
rect 3347 1038 3487 1042
rect 3491 1038 3575 1042
rect 3579 1038 3611 1042
rect 1853 1037 3611 1038
rect 3617 1037 3618 1043
rect 1062 1012 1068 1013
rect 1282 1012 1288 1013
rect 1062 1008 1063 1012
rect 1067 1008 1283 1012
rect 1287 1008 1288 1012
rect 1062 1007 1068 1008
rect 1282 1007 1288 1008
rect 96 993 97 999
rect 103 998 1847 999
rect 103 994 111 998
rect 115 994 143 998
rect 147 994 279 998
rect 283 994 287 998
rect 291 994 439 998
rect 443 994 463 998
rect 467 994 591 998
rect 595 994 647 998
rect 651 994 743 998
rect 747 994 823 998
rect 827 994 895 998
rect 899 994 999 998
rect 1003 994 1055 998
rect 1059 994 1167 998
rect 1171 994 1223 998
rect 1227 994 1327 998
rect 1331 994 1391 998
rect 1395 994 1487 998
rect 1491 994 1567 998
rect 1571 994 1655 998
rect 1659 994 1735 998
rect 1739 994 1823 998
rect 1827 994 1847 998
rect 103 993 1847 994
rect 1853 993 1854 999
rect 1834 965 1835 971
rect 1841 970 3599 971
rect 1841 966 1863 970
rect 1867 966 1887 970
rect 1891 966 1911 970
rect 1915 966 2071 970
rect 2075 966 2119 970
rect 2123 966 2263 970
rect 2267 966 2319 970
rect 2323 966 2455 970
rect 2459 966 2511 970
rect 2515 966 2631 970
rect 2635 966 2687 970
rect 2691 966 2799 970
rect 2803 966 2855 970
rect 2859 966 2951 970
rect 2955 966 3015 970
rect 3019 966 3095 970
rect 3099 966 3175 970
rect 3179 966 3231 970
rect 3235 966 3335 970
rect 3339 966 3367 970
rect 3371 966 3479 970
rect 3483 966 3575 970
rect 3579 966 3599 970
rect 1841 965 3599 966
rect 3605 965 3606 971
rect 84 917 85 923
rect 91 922 1835 923
rect 91 918 111 922
rect 115 918 135 922
rect 139 918 271 922
rect 275 918 279 922
rect 283 918 439 922
rect 443 918 455 922
rect 459 918 607 922
rect 611 918 639 922
rect 643 918 775 922
rect 779 918 815 922
rect 819 918 935 922
rect 939 918 991 922
rect 995 918 1095 922
rect 1099 918 1159 922
rect 1163 918 1247 922
rect 1251 918 1319 922
rect 1323 918 1399 922
rect 1403 918 1479 922
rect 1483 918 1551 922
rect 1555 918 1647 922
rect 1651 918 1823 922
rect 1827 918 1835 922
rect 91 917 1835 918
rect 1841 917 1842 923
rect 2814 916 2820 917
rect 3110 916 3116 917
rect 2814 912 2815 916
rect 2819 912 3111 916
rect 3115 912 3116 916
rect 2814 911 2820 912
rect 3110 911 3116 912
rect 1846 889 1847 895
rect 1853 894 3611 895
rect 1853 890 1863 894
rect 1867 890 1895 894
rect 1899 890 2023 894
rect 2027 890 2079 894
rect 2083 890 2183 894
rect 2187 890 2271 894
rect 2275 890 2351 894
rect 2355 890 2463 894
rect 2467 890 2519 894
rect 2523 890 2639 894
rect 2643 890 2687 894
rect 2691 890 2807 894
rect 2811 890 2839 894
rect 2843 890 2959 894
rect 2963 890 2983 894
rect 2987 890 3103 894
rect 3107 890 3119 894
rect 3123 890 3239 894
rect 3243 890 3247 894
rect 3251 890 3375 894
rect 3379 890 3487 894
rect 3491 890 3575 894
rect 3579 890 3611 894
rect 1853 889 3611 890
rect 3617 889 3618 895
rect 454 868 460 869
rect 706 868 712 869
rect 454 864 455 868
rect 459 864 707 868
rect 711 864 712 868
rect 454 863 460 864
rect 706 863 712 864
rect 1262 868 1268 869
rect 1494 868 1500 869
rect 1262 864 1263 868
rect 1267 864 1495 868
rect 1499 864 1500 868
rect 1262 863 1268 864
rect 1494 863 1500 864
rect 96 849 97 855
rect 103 854 1847 855
rect 103 850 111 854
rect 115 850 143 854
rect 147 850 279 854
rect 283 850 287 854
rect 291 850 447 854
rect 451 850 463 854
rect 467 850 615 854
rect 619 850 639 854
rect 643 850 783 854
rect 787 850 807 854
rect 811 850 943 854
rect 947 850 983 854
rect 987 850 1103 854
rect 1107 850 1159 854
rect 1163 850 1255 854
rect 1259 850 1335 854
rect 1339 850 1407 854
rect 1411 850 1511 854
rect 1515 850 1559 854
rect 1563 850 1823 854
rect 1827 850 1847 854
rect 103 849 1847 850
rect 1853 849 1854 855
rect 1834 813 1835 819
rect 1841 818 3599 819
rect 1841 814 1863 818
rect 1867 814 1887 818
rect 1891 814 2015 818
rect 2019 814 2071 818
rect 2075 814 2175 818
rect 2179 814 2263 818
rect 2267 814 2343 818
rect 2347 814 2447 818
rect 2451 814 2511 818
rect 2515 814 2623 818
rect 2627 814 2679 818
rect 2683 814 2791 818
rect 2795 814 2831 818
rect 2835 814 2943 818
rect 2947 814 2975 818
rect 2979 814 3087 818
rect 3091 814 3111 818
rect 3115 814 3223 818
rect 3227 814 3239 818
rect 3243 814 3359 818
rect 3363 814 3367 818
rect 3371 814 3479 818
rect 3483 814 3575 818
rect 3579 814 3599 818
rect 1841 813 3599 814
rect 3605 813 3606 819
rect 84 777 85 783
rect 91 782 1835 783
rect 91 778 111 782
rect 115 778 135 782
rect 139 778 271 782
rect 275 778 279 782
rect 283 778 439 782
rect 443 778 455 782
rect 459 778 607 782
rect 611 778 631 782
rect 635 778 775 782
rect 779 778 799 782
rect 803 778 935 782
rect 939 778 975 782
rect 979 778 1087 782
rect 1091 778 1151 782
rect 1155 778 1239 782
rect 1243 778 1327 782
rect 1331 778 1391 782
rect 1395 778 1503 782
rect 1507 778 1551 782
rect 1555 778 1823 782
rect 1827 778 1835 782
rect 91 777 1835 778
rect 1841 777 1842 783
rect 1846 745 1847 751
rect 1853 750 3611 751
rect 1853 746 1863 750
rect 1867 746 1895 750
rect 1899 746 2071 750
rect 2075 746 2079 750
rect 2083 746 2263 750
rect 2267 746 2271 750
rect 2275 746 2447 750
rect 2451 746 2455 750
rect 2459 746 2623 750
rect 2627 746 2631 750
rect 2635 746 2799 750
rect 2803 746 2951 750
rect 2955 746 2975 750
rect 2979 746 3095 750
rect 3099 746 3151 750
rect 3155 746 3231 750
rect 3235 746 3327 750
rect 3331 746 3367 750
rect 3371 746 3487 750
rect 3491 746 3575 750
rect 3579 746 3611 750
rect 1853 745 3611 746
rect 3617 745 3618 751
rect 3054 740 3060 741
rect 3258 740 3264 741
rect 3054 736 3055 740
rect 3059 736 3259 740
rect 3263 736 3264 740
rect 3054 735 3060 736
rect 3258 735 3264 736
rect 96 705 97 711
rect 103 710 1847 711
rect 103 706 111 710
rect 115 706 143 710
rect 147 706 279 710
rect 283 706 287 710
rect 291 706 447 710
rect 451 706 455 710
rect 459 706 615 710
rect 619 706 623 710
rect 627 706 783 710
rect 787 706 791 710
rect 795 706 943 710
rect 947 706 959 710
rect 963 706 1095 710
rect 1099 706 1119 710
rect 1123 706 1247 710
rect 1251 706 1279 710
rect 1283 706 1399 710
rect 1403 706 1439 710
rect 1443 706 1559 710
rect 1563 706 1599 710
rect 1603 706 1823 710
rect 1827 706 1847 710
rect 103 705 1847 706
rect 1853 705 1854 711
rect 1834 673 1835 679
rect 1841 678 3599 679
rect 1841 674 1863 678
rect 1867 674 1887 678
rect 1891 674 1975 678
rect 1979 674 2063 678
rect 2067 674 2095 678
rect 2099 674 2223 678
rect 2227 674 2255 678
rect 2259 674 2351 678
rect 2355 674 2439 678
rect 2443 674 2479 678
rect 2483 674 2615 678
rect 2619 674 2767 678
rect 2771 674 2791 678
rect 2795 674 2935 678
rect 2939 674 2967 678
rect 2971 674 3119 678
rect 3123 674 3143 678
rect 3147 674 3311 678
rect 3315 674 3319 678
rect 3323 674 3479 678
rect 3483 674 3575 678
rect 3579 674 3599 678
rect 1841 673 3599 674
rect 3605 673 3606 679
rect 84 629 85 635
rect 91 634 1835 635
rect 91 630 111 634
rect 115 630 135 634
rect 139 630 279 634
rect 283 630 287 634
rect 291 630 447 634
rect 451 630 455 634
rect 459 630 615 634
rect 619 630 631 634
rect 635 630 783 634
rect 787 630 799 634
rect 803 630 951 634
rect 955 630 967 634
rect 971 630 1111 634
rect 1115 630 1119 634
rect 1123 630 1271 634
rect 1275 630 1415 634
rect 1419 630 1431 634
rect 1435 630 1559 634
rect 1563 630 1591 634
rect 1595 630 1711 634
rect 1715 630 1823 634
rect 1827 630 1835 634
rect 91 629 1835 630
rect 1841 629 1842 635
rect 2630 620 2636 621
rect 3234 620 3240 621
rect 2630 616 2631 620
rect 2635 616 3235 620
rect 3239 616 3240 620
rect 2630 615 2636 616
rect 3234 615 3240 616
rect 1846 601 1847 607
rect 1853 606 3611 607
rect 1853 602 1863 606
rect 1867 602 1895 606
rect 1899 602 1983 606
rect 1987 602 2047 606
rect 2051 602 2103 606
rect 2107 602 2215 606
rect 2219 602 2231 606
rect 2235 602 2359 606
rect 2363 602 2391 606
rect 2395 602 2487 606
rect 2491 602 2583 606
rect 2587 602 2623 606
rect 2627 602 2775 606
rect 2779 602 2799 606
rect 2803 602 2943 606
rect 2947 602 3023 606
rect 3027 602 3127 606
rect 3131 602 3255 606
rect 3259 602 3319 606
rect 3323 602 3487 606
rect 3491 602 3575 606
rect 3579 602 3611 606
rect 1853 601 3611 602
rect 3617 601 3618 607
rect 1198 588 1204 589
rect 1638 588 1644 589
rect 1198 584 1199 588
rect 1203 584 1639 588
rect 1643 584 1644 588
rect 1198 583 1204 584
rect 1638 583 1644 584
rect 96 557 97 563
rect 103 562 1847 563
rect 103 558 111 562
rect 115 558 143 562
rect 147 558 151 562
rect 155 558 295 562
rect 299 558 311 562
rect 315 558 463 562
rect 467 558 471 562
rect 475 558 631 562
rect 635 558 639 562
rect 643 558 783 562
rect 787 558 807 562
rect 811 558 927 562
rect 931 558 975 562
rect 979 558 1063 562
rect 1067 558 1127 562
rect 1131 558 1191 562
rect 1195 558 1279 562
rect 1283 558 1311 562
rect 1315 558 1423 562
rect 1427 558 1535 562
rect 1539 558 1567 562
rect 1571 558 1647 562
rect 1651 558 1719 562
rect 1723 558 1735 562
rect 1739 558 1823 562
rect 1827 558 1847 562
rect 103 557 1847 558
rect 1853 557 1854 563
rect 1834 525 1835 531
rect 1841 530 3599 531
rect 1841 526 1863 530
rect 1867 526 1887 530
rect 1891 526 2039 530
rect 2043 526 2191 530
rect 2195 526 2207 530
rect 2211 526 2279 530
rect 2283 526 2375 530
rect 2379 526 2383 530
rect 2387 526 2487 530
rect 2491 526 2575 530
rect 2579 526 2631 530
rect 2635 526 2791 530
rect 2795 526 2807 530
rect 2811 526 3007 530
rect 3011 526 3015 530
rect 3019 526 3215 530
rect 3219 526 3247 530
rect 3251 526 3431 530
rect 3435 526 3479 530
rect 3483 526 3575 530
rect 3579 526 3599 530
rect 1841 525 3599 526
rect 3605 525 3606 531
rect 2390 492 2396 493
rect 3186 492 3192 493
rect 2390 488 2391 492
rect 2395 488 3187 492
rect 3191 488 3192 492
rect 2390 487 2396 488
rect 3186 487 3192 488
rect 84 481 85 487
rect 91 486 1835 487
rect 91 482 111 486
rect 115 482 143 486
rect 147 482 159 486
rect 163 482 303 486
rect 307 482 311 486
rect 315 482 463 486
rect 467 482 615 486
rect 619 482 623 486
rect 627 482 759 486
rect 763 482 775 486
rect 779 482 887 486
rect 891 482 919 486
rect 923 482 1007 486
rect 1011 482 1055 486
rect 1059 482 1127 486
rect 1131 482 1183 486
rect 1187 482 1239 486
rect 1243 482 1303 486
rect 1307 482 1343 486
rect 1347 482 1415 486
rect 1419 482 1439 486
rect 1443 482 1527 486
rect 1531 482 1543 486
rect 1547 482 1639 486
rect 1643 482 1727 486
rect 1731 482 1823 486
rect 1827 482 1835 486
rect 91 481 1835 482
rect 1841 481 1842 487
rect 1846 449 1847 455
rect 1853 454 3611 455
rect 1853 450 1863 454
rect 1867 450 1895 454
rect 1899 450 2039 454
rect 2043 450 2199 454
rect 2203 450 2207 454
rect 2211 450 2287 454
rect 2291 450 2383 454
rect 2387 450 2495 454
rect 2499 450 2575 454
rect 2579 450 2639 454
rect 2643 450 2783 454
rect 2787 450 2815 454
rect 2819 450 3007 454
rect 3011 450 3015 454
rect 3019 450 3223 454
rect 3227 450 3239 454
rect 3243 450 3439 454
rect 3443 450 3471 454
rect 3475 450 3575 454
rect 3579 450 3611 454
rect 1853 449 3611 450
rect 3617 449 3618 455
rect 1142 428 1148 429
rect 1490 428 1496 429
rect 1142 424 1143 428
rect 1147 424 1491 428
rect 1495 424 1496 428
rect 1142 423 1148 424
rect 1490 423 1496 424
rect 96 413 97 419
rect 103 418 1847 419
rect 103 414 111 418
rect 115 414 151 418
rect 155 414 167 418
rect 171 414 271 418
rect 275 414 319 418
rect 323 414 407 418
rect 411 414 471 418
rect 475 414 551 418
rect 555 414 623 418
rect 627 414 711 418
rect 715 414 767 418
rect 771 414 887 418
rect 891 414 895 418
rect 899 414 1015 418
rect 1019 414 1063 418
rect 1067 414 1135 418
rect 1139 414 1247 418
rect 1251 414 1351 418
rect 1355 414 1439 418
rect 1443 414 1447 418
rect 1451 414 1551 418
rect 1555 414 1639 418
rect 1643 414 1647 418
rect 1651 414 1735 418
rect 1739 414 1823 418
rect 1827 414 1847 418
rect 103 413 1847 414
rect 1853 413 1854 419
rect 902 396 908 397
rect 1162 396 1168 397
rect 902 392 903 396
rect 907 392 1163 396
rect 1167 392 1168 396
rect 902 391 908 392
rect 1162 391 1168 392
rect 158 388 164 389
rect 338 388 344 389
rect 158 384 159 388
rect 163 384 339 388
rect 343 384 344 388
rect 158 383 164 384
rect 338 383 344 384
rect 1834 381 1835 387
rect 1841 386 3599 387
rect 1841 382 1863 386
rect 1867 382 1887 386
rect 1891 382 1975 386
rect 1979 382 2031 386
rect 2035 382 2063 386
rect 2067 382 2151 386
rect 2155 382 2199 386
rect 2203 382 2263 386
rect 2267 382 2375 386
rect 2379 382 2383 386
rect 2387 382 2519 386
rect 2523 382 2567 386
rect 2571 382 2671 386
rect 2675 382 2775 386
rect 2779 382 2847 386
rect 2851 382 2999 386
rect 3003 382 3031 386
rect 3035 382 3231 386
rect 3235 382 3431 386
rect 3435 382 3463 386
rect 3467 382 3575 386
rect 3579 382 3599 386
rect 1841 381 3599 382
rect 3605 381 3606 387
rect 2702 348 2708 349
rect 3158 348 3164 349
rect 2702 344 2703 348
rect 2707 344 3159 348
rect 3163 344 3164 348
rect 2702 343 2708 344
rect 3158 343 3164 344
rect 84 329 85 335
rect 91 334 1835 335
rect 91 330 111 334
rect 115 330 135 334
rect 139 330 143 334
rect 147 330 223 334
rect 227 330 263 334
rect 267 330 311 334
rect 315 330 399 334
rect 403 330 487 334
rect 491 330 543 334
rect 547 330 575 334
rect 579 330 663 334
rect 667 330 703 334
rect 707 330 751 334
rect 755 330 839 334
rect 843 330 879 334
rect 883 330 927 334
rect 931 330 1015 334
rect 1019 330 1055 334
rect 1059 330 1103 334
rect 1107 330 1191 334
rect 1195 330 1239 334
rect 1243 330 1287 334
rect 1291 330 1383 334
rect 1387 330 1431 334
rect 1435 330 1479 334
rect 1483 330 1575 334
rect 1579 330 1631 334
rect 1635 330 1671 334
rect 1675 330 1823 334
rect 1827 330 1835 334
rect 91 329 1835 330
rect 1841 329 1842 335
rect 2686 332 2692 333
rect 3178 332 3184 333
rect 2686 328 2687 332
rect 2691 328 3179 332
rect 3183 328 3184 332
rect 2686 327 2692 328
rect 3178 327 3184 328
rect 1846 313 1847 319
rect 1853 318 3611 319
rect 1853 314 1863 318
rect 1867 314 1895 318
rect 1899 314 1983 318
rect 1987 314 2071 318
rect 2075 314 2159 318
rect 2163 314 2247 318
rect 2251 314 2271 318
rect 2275 314 2359 318
rect 2363 314 2391 318
rect 2395 314 2471 318
rect 2475 314 2527 318
rect 2531 314 2583 318
rect 2587 314 2679 318
rect 2683 314 2695 318
rect 2699 314 2807 318
rect 2811 314 2855 318
rect 2859 314 2919 318
rect 2923 314 3039 318
rect 3043 314 3159 318
rect 3163 314 3239 318
rect 3243 314 3439 318
rect 3443 314 3575 318
rect 3579 314 3611 318
rect 1853 313 3611 314
rect 3617 313 3618 319
rect 2366 308 2372 309
rect 2542 308 2548 309
rect 2366 304 2367 308
rect 2371 304 2543 308
rect 2547 304 2548 308
rect 2366 303 2372 304
rect 2542 303 2548 304
rect 1302 276 1308 277
rect 1562 276 1568 277
rect 1302 272 1303 276
rect 1307 272 1563 276
rect 1567 272 1568 276
rect 1302 271 1308 272
rect 1562 271 1568 272
rect 96 257 97 263
rect 103 262 1847 263
rect 103 258 111 262
rect 115 258 143 262
rect 147 258 231 262
rect 235 258 319 262
rect 323 258 407 262
rect 411 258 495 262
rect 499 258 583 262
rect 587 258 671 262
rect 675 258 759 262
rect 763 258 847 262
rect 851 258 935 262
rect 939 258 1023 262
rect 1027 258 1111 262
rect 1115 258 1199 262
rect 1203 258 1287 262
rect 1291 258 1295 262
rect 1299 258 1375 262
rect 1379 258 1391 262
rect 1395 258 1463 262
rect 1467 258 1487 262
rect 1491 258 1551 262
rect 1555 258 1583 262
rect 1587 258 1639 262
rect 1643 258 1679 262
rect 1683 258 1727 262
rect 1731 258 1823 262
rect 1827 258 1847 262
rect 103 257 1847 258
rect 1853 257 1854 263
rect 1030 252 1036 253
rect 1266 252 1272 253
rect 1030 248 1031 252
rect 1035 248 1267 252
rect 1271 248 1272 252
rect 1030 247 1036 248
rect 1266 247 1272 248
rect 1834 245 1835 251
rect 1841 250 3599 251
rect 1841 246 1863 250
rect 1867 246 1887 250
rect 1891 246 1975 250
rect 1979 246 2063 250
rect 2067 246 2151 250
rect 2155 246 2239 250
rect 2243 246 2263 250
rect 2267 246 2351 250
rect 2355 246 2399 250
rect 2403 246 2463 250
rect 2467 246 2535 250
rect 2539 246 2575 250
rect 2579 246 2679 250
rect 2683 246 2687 250
rect 2691 246 2799 250
rect 2803 246 2815 250
rect 2819 246 2911 250
rect 2915 246 2951 250
rect 2955 246 3031 250
rect 3035 246 3087 250
rect 3091 246 3151 250
rect 3155 246 3223 250
rect 3227 246 3359 250
rect 3363 246 3479 250
rect 3483 246 3575 250
rect 3579 246 3599 250
rect 1841 245 3599 246
rect 3605 245 3606 251
rect 1902 228 1908 229
rect 2226 228 2232 229
rect 1902 224 1903 228
rect 1907 224 2227 228
rect 2231 224 2232 228
rect 1902 223 1908 224
rect 2226 223 2232 224
rect 2830 196 2836 197
rect 3106 196 3112 197
rect 84 189 85 195
rect 91 194 1835 195
rect 91 190 111 194
rect 115 190 135 194
rect 139 190 223 194
rect 227 190 311 194
rect 315 190 399 194
rect 403 190 487 194
rect 491 190 575 194
rect 579 190 663 194
rect 667 190 751 194
rect 755 190 839 194
rect 843 190 927 194
rect 931 190 1015 194
rect 1019 190 1103 194
rect 1107 190 1191 194
rect 1195 190 1279 194
rect 1283 190 1367 194
rect 1371 190 1455 194
rect 1459 190 1543 194
rect 1547 190 1631 194
rect 1635 190 1719 194
rect 1723 190 1823 194
rect 1827 190 1835 194
rect 91 189 1835 190
rect 1841 189 1842 195
rect 2830 192 2831 196
rect 2835 192 3107 196
rect 3111 192 3112 196
rect 2830 191 2836 192
rect 3106 191 3112 192
rect 2790 180 2796 181
rect 3190 180 3196 181
rect 2790 176 2791 180
rect 2795 176 3191 180
rect 3195 176 3196 180
rect 2790 175 2796 176
rect 3190 175 3196 176
rect 1846 145 1847 151
rect 1853 150 3611 151
rect 1853 146 1863 150
rect 1867 146 1895 150
rect 1899 146 1983 150
rect 1987 146 2071 150
rect 2075 146 2159 150
rect 2163 146 2271 150
rect 2275 146 2407 150
rect 2411 146 2543 150
rect 2547 146 2687 150
rect 2691 146 2783 150
rect 2787 146 2823 150
rect 2827 146 2871 150
rect 2875 146 2959 150
rect 2963 146 3047 150
rect 3051 146 3095 150
rect 3099 146 3135 150
rect 3139 146 3223 150
rect 3227 146 3231 150
rect 3235 146 3311 150
rect 3315 146 3367 150
rect 3371 146 3399 150
rect 3403 146 3487 150
rect 3491 146 3575 150
rect 3579 146 3611 150
rect 1853 145 3611 146
rect 3617 145 3618 151
rect 1834 77 1835 83
rect 1841 82 3599 83
rect 1841 78 1863 82
rect 1867 78 2775 82
rect 2779 78 2863 82
rect 2867 78 2951 82
rect 2955 78 3039 82
rect 3043 78 3127 82
rect 3131 78 3215 82
rect 3219 78 3303 82
rect 3307 78 3391 82
rect 3395 78 3479 82
rect 3483 78 3575 82
rect 3579 78 3599 82
rect 1841 77 3599 78
rect 3605 77 3606 83
<< m5c >>
rect 85 3665 91 3671
rect 1835 3665 1841 3671
rect 1835 3607 1841 3613
rect 97 3597 103 3603
rect 1847 3597 1853 3603
rect 3599 3589 3605 3595
rect 85 3529 91 3535
rect 1835 3529 1841 3535
rect 1847 3521 1853 3527
rect 3611 3521 3617 3527
rect 97 3461 103 3467
rect 1847 3461 1853 3467
rect 1835 3445 1841 3451
rect 3599 3445 3605 3451
rect 85 3393 91 3399
rect 1835 3393 1841 3399
rect 1847 3369 1853 3375
rect 3611 3369 3617 3375
rect 97 3321 103 3327
rect 1847 3321 1853 3327
rect 1835 3301 1841 3307
rect 3599 3301 3605 3307
rect 85 3249 91 3255
rect 1835 3249 1841 3255
rect 1847 3225 1853 3231
rect 3611 3225 3617 3231
rect 97 3173 103 3179
rect 1847 3173 1853 3179
rect 1835 3153 1841 3159
rect 3599 3153 3605 3159
rect 85 3097 91 3103
rect 1835 3097 1841 3103
rect 1847 3077 1853 3083
rect 3611 3077 3617 3083
rect 97 3025 103 3031
rect 1847 3025 1853 3031
rect 1835 3005 1841 3011
rect 3599 3005 3605 3011
rect 85 2957 91 2963
rect 1835 2957 1841 2963
rect 1847 2929 1853 2935
rect 3611 2929 3617 2935
rect 97 2885 103 2891
rect 1847 2885 1853 2891
rect 1835 2861 1841 2867
rect 3599 2861 3605 2867
rect 85 2809 91 2815
rect 1835 2809 1841 2815
rect 1847 2793 1853 2799
rect 3611 2793 3617 2799
rect 97 2733 103 2739
rect 1847 2733 1853 2739
rect 1835 2721 1841 2727
rect 3599 2721 3605 2727
rect 85 2661 91 2667
rect 1835 2661 1841 2667
rect 1847 2645 1853 2651
rect 3611 2645 3617 2651
rect 97 2589 103 2595
rect 1847 2589 1853 2595
rect 1835 2573 1841 2579
rect 3599 2573 3605 2579
rect 85 2521 91 2527
rect 1835 2521 1841 2527
rect 1847 2501 1853 2507
rect 3611 2501 3617 2507
rect 97 2453 103 2459
rect 1847 2453 1853 2459
rect 1835 2433 1841 2439
rect 3599 2433 3605 2439
rect 85 2373 91 2379
rect 1835 2373 1841 2379
rect 1847 2361 1853 2367
rect 3611 2361 3617 2367
rect 1835 2307 1841 2313
rect 97 2297 103 2303
rect 1847 2297 1853 2303
rect 3599 2289 3605 2295
rect 85 2221 91 2227
rect 1835 2221 1841 2227
rect 1847 2221 1853 2227
rect 3611 2221 3617 2227
rect 1835 2163 1841 2169
rect 97 2153 103 2159
rect 1847 2153 1853 2159
rect 3599 2145 3605 2151
rect 575 2116 581 2117
rect 575 2112 579 2116
rect 579 2112 581 2116
rect 575 2111 581 2112
rect 1039 2108 1045 2109
rect 1039 2104 1043 2108
rect 1043 2104 1045 2108
rect 1039 2103 1045 2104
rect 85 2081 91 2087
rect 1835 2081 1841 2087
rect 1847 2073 1853 2079
rect 3611 2073 3617 2079
rect 1835 2019 1841 2025
rect 97 2009 103 2015
rect 1847 2009 1853 2015
rect 3599 2005 3605 2011
rect 85 1937 91 1943
rect 1835 1937 1841 1943
rect 1847 1929 1853 1935
rect 3611 1929 3617 1935
rect 1835 1871 1841 1877
rect 97 1861 103 1867
rect 1847 1861 1853 1867
rect 3599 1853 3605 1859
rect 85 1781 91 1787
rect 1835 1781 1841 1787
rect 1847 1781 1853 1787
rect 3611 1781 3617 1787
rect 1835 1719 1841 1725
rect 97 1709 103 1715
rect 1847 1709 1853 1715
rect 3599 1709 3605 1715
rect 85 1633 91 1639
rect 1835 1633 1841 1639
rect 1847 1637 1853 1643
rect 3611 1637 3617 1643
rect 1835 1575 1841 1581
rect 97 1565 103 1571
rect 1847 1565 1853 1571
rect 3599 1569 3605 1575
rect 85 1493 91 1499
rect 1835 1493 1841 1499
rect 1847 1493 1853 1499
rect 3611 1493 3617 1499
rect 1835 1427 1841 1433
rect 97 1417 103 1423
rect 1847 1417 1853 1423
rect 3599 1421 3605 1427
rect 85 1345 91 1351
rect 1835 1345 1841 1351
rect 1847 1349 1853 1355
rect 3611 1349 3617 1355
rect 1835 1287 1841 1293
rect 97 1277 103 1283
rect 1847 1277 1853 1283
rect 3599 1269 3605 1275
rect 85 1201 91 1207
rect 1835 1201 1841 1207
rect 1847 1197 1853 1203
rect 3611 1197 3617 1203
rect 97 1133 103 1139
rect 1847 1133 1853 1139
rect 1835 1117 1841 1123
rect 3599 1117 3605 1123
rect 85 1065 91 1071
rect 1835 1065 1841 1071
rect 1847 1037 1853 1043
rect 3611 1037 3617 1043
rect 97 993 103 999
rect 1847 993 1853 999
rect 1835 965 1841 971
rect 3599 965 3605 971
rect 85 917 91 923
rect 1835 917 1841 923
rect 1847 889 1853 895
rect 3611 889 3617 895
rect 97 849 103 855
rect 1847 849 1853 855
rect 1835 813 1841 819
rect 3599 813 3605 819
rect 85 777 91 783
rect 1835 777 1841 783
rect 1847 745 1853 751
rect 3611 745 3617 751
rect 97 705 103 711
rect 1847 705 1853 711
rect 1835 673 1841 679
rect 3599 673 3605 679
rect 85 629 91 635
rect 1835 629 1841 635
rect 1847 601 1853 607
rect 3611 601 3617 607
rect 97 557 103 563
rect 1847 557 1853 563
rect 1835 525 1841 531
rect 3599 525 3605 531
rect 85 481 91 487
rect 1835 481 1841 487
rect 1847 449 1853 455
rect 3611 449 3617 455
rect 97 413 103 419
rect 1847 413 1853 419
rect 1835 381 1841 387
rect 3599 381 3605 387
rect 85 329 91 335
rect 1835 329 1841 335
rect 1847 313 1853 319
rect 3611 313 3617 319
rect 97 257 103 263
rect 1847 257 1853 263
rect 1835 245 1841 251
rect 3599 245 3605 251
rect 85 189 91 195
rect 1835 189 1841 195
rect 1847 145 1853 151
rect 3611 145 3617 151
rect 1835 77 1841 83
rect 3599 77 3605 83
<< m5 >>
rect 84 3671 92 3672
rect 84 3665 85 3671
rect 91 3665 92 3671
rect 84 3535 92 3665
rect 84 3529 85 3535
rect 91 3529 92 3535
rect 84 3399 92 3529
rect 84 3393 85 3399
rect 91 3393 92 3399
rect 84 3255 92 3393
rect 84 3249 85 3255
rect 91 3249 92 3255
rect 84 3103 92 3249
rect 84 3097 85 3103
rect 91 3097 92 3103
rect 84 2963 92 3097
rect 84 2957 85 2963
rect 91 2957 92 2963
rect 84 2815 92 2957
rect 84 2809 85 2815
rect 91 2809 92 2815
rect 84 2667 92 2809
rect 84 2661 85 2667
rect 91 2661 92 2667
rect 84 2527 92 2661
rect 84 2521 85 2527
rect 91 2521 92 2527
rect 84 2379 92 2521
rect 84 2373 85 2379
rect 91 2373 92 2379
rect 84 2227 92 2373
rect 84 2221 85 2227
rect 91 2221 92 2227
rect 84 2087 92 2221
rect 84 2081 85 2087
rect 91 2081 92 2087
rect 84 1943 92 2081
rect 84 1937 85 1943
rect 91 1937 92 1943
rect 84 1787 92 1937
rect 84 1781 85 1787
rect 91 1781 92 1787
rect 84 1639 92 1781
rect 84 1633 85 1639
rect 91 1633 92 1639
rect 84 1499 92 1633
rect 84 1493 85 1499
rect 91 1493 92 1499
rect 84 1351 92 1493
rect 84 1345 85 1351
rect 91 1345 92 1351
rect 84 1207 92 1345
rect 84 1201 85 1207
rect 91 1201 92 1207
rect 84 1071 92 1201
rect 84 1065 85 1071
rect 91 1065 92 1071
rect 84 923 92 1065
rect 84 917 85 923
rect 91 917 92 923
rect 84 783 92 917
rect 84 777 85 783
rect 91 777 92 783
rect 84 635 92 777
rect 84 629 85 635
rect 91 629 92 635
rect 84 487 92 629
rect 84 481 85 487
rect 91 481 92 487
rect 84 335 92 481
rect 84 329 85 335
rect 91 329 92 335
rect 84 195 92 329
rect 84 189 85 195
rect 91 189 92 195
rect 84 72 92 189
rect 96 3603 104 3672
rect 96 3597 97 3603
rect 103 3597 104 3603
rect 96 3467 104 3597
rect 96 3461 97 3467
rect 103 3461 104 3467
rect 96 3327 104 3461
rect 96 3321 97 3327
rect 103 3321 104 3327
rect 96 3179 104 3321
rect 96 3173 97 3179
rect 103 3173 104 3179
rect 96 3031 104 3173
rect 96 3025 97 3031
rect 103 3025 104 3031
rect 96 2891 104 3025
rect 96 2885 97 2891
rect 103 2885 104 2891
rect 96 2739 104 2885
rect 96 2733 97 2739
rect 103 2733 104 2739
rect 96 2595 104 2733
rect 96 2589 97 2595
rect 103 2589 104 2595
rect 96 2459 104 2589
rect 96 2453 97 2459
rect 103 2453 104 2459
rect 96 2303 104 2453
rect 96 2297 97 2303
rect 103 2297 104 2303
rect 96 2159 104 2297
rect 96 2153 97 2159
rect 103 2153 104 2159
rect 96 2015 104 2153
rect 1834 3671 1842 3672
rect 1834 3665 1835 3671
rect 1841 3665 1842 3671
rect 1834 3613 1842 3665
rect 1834 3607 1835 3613
rect 1841 3607 1842 3613
rect 1834 3535 1842 3607
rect 1834 3529 1835 3535
rect 1841 3529 1842 3535
rect 1834 3451 1842 3529
rect 1834 3445 1835 3451
rect 1841 3445 1842 3451
rect 1834 3399 1842 3445
rect 1834 3393 1835 3399
rect 1841 3393 1842 3399
rect 1834 3307 1842 3393
rect 1834 3301 1835 3307
rect 1841 3301 1842 3307
rect 1834 3255 1842 3301
rect 1834 3249 1835 3255
rect 1841 3249 1842 3255
rect 1834 3159 1842 3249
rect 1834 3153 1835 3159
rect 1841 3153 1842 3159
rect 1834 3103 1842 3153
rect 1834 3097 1835 3103
rect 1841 3097 1842 3103
rect 1834 3011 1842 3097
rect 1834 3005 1835 3011
rect 1841 3005 1842 3011
rect 1834 2963 1842 3005
rect 1834 2957 1835 2963
rect 1841 2957 1842 2963
rect 1834 2867 1842 2957
rect 1834 2861 1835 2867
rect 1841 2861 1842 2867
rect 1834 2815 1842 2861
rect 1834 2809 1835 2815
rect 1841 2809 1842 2815
rect 1834 2727 1842 2809
rect 1834 2721 1835 2727
rect 1841 2721 1842 2727
rect 1834 2667 1842 2721
rect 1834 2661 1835 2667
rect 1841 2661 1842 2667
rect 1834 2579 1842 2661
rect 1834 2573 1835 2579
rect 1841 2573 1842 2579
rect 1834 2527 1842 2573
rect 1834 2521 1835 2527
rect 1841 2521 1842 2527
rect 1834 2439 1842 2521
rect 1834 2433 1835 2439
rect 1841 2433 1842 2439
rect 1834 2379 1842 2433
rect 1834 2373 1835 2379
rect 1841 2373 1842 2379
rect 1834 2313 1842 2373
rect 1834 2307 1835 2313
rect 1841 2307 1842 2313
rect 1834 2227 1842 2307
rect 1834 2221 1835 2227
rect 1841 2221 1842 2227
rect 1834 2169 1842 2221
rect 1834 2163 1835 2169
rect 1841 2163 1842 2169
rect 574 2117 582 2118
rect 574 2115 575 2117
rect 581 2115 582 2117
rect 96 2009 97 2015
rect 103 2009 104 2015
rect 96 1867 104 2009
rect 96 1861 97 1867
rect 103 1861 104 1867
rect 96 1715 104 1861
rect 96 1709 97 1715
rect 103 1709 104 1715
rect 96 1571 104 1709
rect 96 1565 97 1571
rect 103 1565 104 1571
rect 96 1423 104 1565
rect 96 1417 97 1423
rect 103 1417 104 1423
rect 96 1283 104 1417
rect 96 1277 97 1283
rect 103 1277 104 1283
rect 96 1139 104 1277
rect 96 1133 97 1139
rect 103 1133 104 1139
rect 96 999 104 1133
rect 96 993 97 999
rect 103 993 104 999
rect 96 855 104 993
rect 96 849 97 855
rect 103 849 104 855
rect 96 711 104 849
rect 96 705 97 711
rect 103 705 104 711
rect 96 563 104 705
rect 96 557 97 563
rect 103 557 104 563
rect 96 419 104 557
rect 96 413 97 419
rect 103 413 104 419
rect 96 263 104 413
rect 96 257 97 263
rect 103 257 104 263
rect 96 72 104 257
rect 1834 2087 1842 2163
rect 1834 2081 1835 2087
rect 1841 2081 1842 2087
rect 1834 2025 1842 2081
rect 1834 2019 1835 2025
rect 1841 2019 1842 2025
rect 1834 1943 1842 2019
rect 1834 1937 1835 1943
rect 1841 1937 1842 1943
rect 1834 1877 1842 1937
rect 1834 1871 1835 1877
rect 1841 1871 1842 1877
rect 1834 1787 1842 1871
rect 1834 1781 1835 1787
rect 1841 1781 1842 1787
rect 1834 1725 1842 1781
rect 1834 1719 1835 1725
rect 1841 1719 1842 1725
rect 1834 1639 1842 1719
rect 1834 1633 1835 1639
rect 1841 1633 1842 1639
rect 1834 1581 1842 1633
rect 1834 1575 1835 1581
rect 1841 1575 1842 1581
rect 1834 1499 1842 1575
rect 1834 1493 1835 1499
rect 1841 1493 1842 1499
rect 1834 1433 1842 1493
rect 1834 1427 1835 1433
rect 1841 1427 1842 1433
rect 1834 1351 1842 1427
rect 1834 1345 1835 1351
rect 1841 1345 1842 1351
rect 1834 1293 1842 1345
rect 1834 1287 1835 1293
rect 1841 1287 1842 1293
rect 1834 1207 1842 1287
rect 1834 1201 1835 1207
rect 1841 1201 1842 1207
rect 1834 1123 1842 1201
rect 1834 1117 1835 1123
rect 1841 1117 1842 1123
rect 1834 1071 1842 1117
rect 1834 1065 1835 1071
rect 1841 1065 1842 1071
rect 1834 971 1842 1065
rect 1834 965 1835 971
rect 1841 965 1842 971
rect 1834 923 1842 965
rect 1834 917 1835 923
rect 1841 917 1842 923
rect 1834 819 1842 917
rect 1834 813 1835 819
rect 1841 813 1842 819
rect 1834 783 1842 813
rect 1834 777 1835 783
rect 1841 777 1842 783
rect 1834 679 1842 777
rect 1834 673 1835 679
rect 1841 673 1842 679
rect 1834 635 1842 673
rect 1834 629 1835 635
rect 1841 629 1842 635
rect 1834 531 1842 629
rect 1834 525 1835 531
rect 1841 525 1842 531
rect 1834 487 1842 525
rect 1834 481 1835 487
rect 1841 481 1842 487
rect 1834 387 1842 481
rect 1834 381 1835 387
rect 1841 381 1842 387
rect 1834 335 1842 381
rect 1834 329 1835 335
rect 1841 329 1842 335
rect 1834 251 1842 329
rect 1834 245 1835 251
rect 1841 245 1842 251
rect 1834 195 1842 245
rect 1834 189 1835 195
rect 1841 189 1842 195
rect 1834 83 1842 189
rect 1834 77 1835 83
rect 1841 77 1842 83
rect 1834 72 1842 77
rect 1846 3603 1854 3672
rect 1846 3597 1847 3603
rect 1853 3597 1854 3603
rect 1846 3527 1854 3597
rect 1846 3521 1847 3527
rect 1853 3521 1854 3527
rect 1846 3467 1854 3521
rect 1846 3461 1847 3467
rect 1853 3461 1854 3467
rect 1846 3375 1854 3461
rect 1846 3369 1847 3375
rect 1853 3369 1854 3375
rect 1846 3327 1854 3369
rect 1846 3321 1847 3327
rect 1853 3321 1854 3327
rect 1846 3231 1854 3321
rect 1846 3225 1847 3231
rect 1853 3225 1854 3231
rect 1846 3179 1854 3225
rect 1846 3173 1847 3179
rect 1853 3173 1854 3179
rect 1846 3083 1854 3173
rect 1846 3077 1847 3083
rect 1853 3077 1854 3083
rect 1846 3031 1854 3077
rect 1846 3025 1847 3031
rect 1853 3025 1854 3031
rect 1846 2935 1854 3025
rect 1846 2929 1847 2935
rect 1853 2929 1854 2935
rect 1846 2891 1854 2929
rect 1846 2885 1847 2891
rect 1853 2885 1854 2891
rect 1846 2799 1854 2885
rect 1846 2793 1847 2799
rect 1853 2793 1854 2799
rect 1846 2739 1854 2793
rect 1846 2733 1847 2739
rect 1853 2733 1854 2739
rect 1846 2651 1854 2733
rect 1846 2645 1847 2651
rect 1853 2645 1854 2651
rect 1846 2595 1854 2645
rect 1846 2589 1847 2595
rect 1853 2589 1854 2595
rect 1846 2507 1854 2589
rect 1846 2501 1847 2507
rect 1853 2501 1854 2507
rect 1846 2459 1854 2501
rect 1846 2453 1847 2459
rect 1853 2453 1854 2459
rect 1846 2367 1854 2453
rect 1846 2361 1847 2367
rect 1853 2361 1854 2367
rect 1846 2303 1854 2361
rect 1846 2297 1847 2303
rect 1853 2297 1854 2303
rect 1846 2227 1854 2297
rect 1846 2221 1847 2227
rect 1853 2221 1854 2227
rect 1846 2159 1854 2221
rect 1846 2153 1847 2159
rect 1853 2153 1854 2159
rect 1846 2079 1854 2153
rect 1846 2073 1847 2079
rect 1853 2073 1854 2079
rect 1846 2015 1854 2073
rect 1846 2009 1847 2015
rect 1853 2009 1854 2015
rect 1846 1935 1854 2009
rect 1846 1929 1847 1935
rect 1853 1929 1854 1935
rect 1846 1867 1854 1929
rect 1846 1861 1847 1867
rect 1853 1861 1854 1867
rect 1846 1787 1854 1861
rect 1846 1781 1847 1787
rect 1853 1781 1854 1787
rect 1846 1715 1854 1781
rect 1846 1709 1847 1715
rect 1853 1709 1854 1715
rect 1846 1643 1854 1709
rect 1846 1637 1847 1643
rect 1853 1637 1854 1643
rect 1846 1571 1854 1637
rect 1846 1565 1847 1571
rect 1853 1565 1854 1571
rect 1846 1499 1854 1565
rect 1846 1493 1847 1499
rect 1853 1493 1854 1499
rect 1846 1423 1854 1493
rect 1846 1417 1847 1423
rect 1853 1417 1854 1423
rect 1846 1355 1854 1417
rect 1846 1349 1847 1355
rect 1853 1349 1854 1355
rect 1846 1283 1854 1349
rect 1846 1277 1847 1283
rect 1853 1277 1854 1283
rect 1846 1203 1854 1277
rect 1846 1197 1847 1203
rect 1853 1197 1854 1203
rect 1846 1139 1854 1197
rect 1846 1133 1847 1139
rect 1853 1133 1854 1139
rect 1846 1043 1854 1133
rect 1846 1037 1847 1043
rect 1853 1037 1854 1043
rect 1846 999 1854 1037
rect 1846 993 1847 999
rect 1853 993 1854 999
rect 1846 895 1854 993
rect 1846 889 1847 895
rect 1853 889 1854 895
rect 1846 855 1854 889
rect 1846 849 1847 855
rect 1853 849 1854 855
rect 1846 751 1854 849
rect 1846 745 1847 751
rect 1853 745 1854 751
rect 1846 711 1854 745
rect 1846 705 1847 711
rect 1853 705 1854 711
rect 1846 607 1854 705
rect 1846 601 1847 607
rect 1853 601 1854 607
rect 1846 563 1854 601
rect 1846 557 1847 563
rect 1853 557 1854 563
rect 1846 455 1854 557
rect 1846 449 1847 455
rect 1853 449 1854 455
rect 1846 419 1854 449
rect 1846 413 1847 419
rect 1853 413 1854 419
rect 1846 319 1854 413
rect 1846 313 1847 319
rect 1853 313 1854 319
rect 1846 263 1854 313
rect 1846 257 1847 263
rect 1853 257 1854 263
rect 1846 151 1854 257
rect 1846 145 1847 151
rect 1853 145 1854 151
rect 1846 72 1854 145
rect 3598 3595 3606 3672
rect 3598 3589 3599 3595
rect 3605 3589 3606 3595
rect 3598 3451 3606 3589
rect 3598 3445 3599 3451
rect 3605 3445 3606 3451
rect 3598 3307 3606 3445
rect 3598 3301 3599 3307
rect 3605 3301 3606 3307
rect 3598 3159 3606 3301
rect 3598 3153 3599 3159
rect 3605 3153 3606 3159
rect 3598 3011 3606 3153
rect 3598 3005 3599 3011
rect 3605 3005 3606 3011
rect 3598 2867 3606 3005
rect 3598 2861 3599 2867
rect 3605 2861 3606 2867
rect 3598 2727 3606 2861
rect 3598 2721 3599 2727
rect 3605 2721 3606 2727
rect 3598 2579 3606 2721
rect 3598 2573 3599 2579
rect 3605 2573 3606 2579
rect 3598 2439 3606 2573
rect 3598 2433 3599 2439
rect 3605 2433 3606 2439
rect 3598 2295 3606 2433
rect 3598 2289 3599 2295
rect 3605 2289 3606 2295
rect 3598 2151 3606 2289
rect 3598 2145 3599 2151
rect 3605 2145 3606 2151
rect 3598 2011 3606 2145
rect 3598 2005 3599 2011
rect 3605 2005 3606 2011
rect 3598 1859 3606 2005
rect 3598 1853 3599 1859
rect 3605 1853 3606 1859
rect 3598 1715 3606 1853
rect 3598 1709 3599 1715
rect 3605 1709 3606 1715
rect 3598 1575 3606 1709
rect 3598 1569 3599 1575
rect 3605 1569 3606 1575
rect 3598 1427 3606 1569
rect 3598 1421 3599 1427
rect 3605 1421 3606 1427
rect 3598 1275 3606 1421
rect 3598 1269 3599 1275
rect 3605 1269 3606 1275
rect 3598 1123 3606 1269
rect 3598 1117 3599 1123
rect 3605 1117 3606 1123
rect 3598 971 3606 1117
rect 3598 965 3599 971
rect 3605 965 3606 971
rect 3598 819 3606 965
rect 3598 813 3599 819
rect 3605 813 3606 819
rect 3598 679 3606 813
rect 3598 673 3599 679
rect 3605 673 3606 679
rect 3598 531 3606 673
rect 3598 525 3599 531
rect 3605 525 3606 531
rect 3598 387 3606 525
rect 3598 381 3599 387
rect 3605 381 3606 387
rect 3598 251 3606 381
rect 3598 245 3599 251
rect 3605 245 3606 251
rect 3598 83 3606 245
rect 3598 77 3599 83
rect 3605 77 3606 83
rect 3598 72 3606 77
rect 3610 3527 3618 3672
rect 3610 3521 3611 3527
rect 3617 3521 3618 3527
rect 3610 3375 3618 3521
rect 3610 3369 3611 3375
rect 3617 3369 3618 3375
rect 3610 3231 3618 3369
rect 3610 3225 3611 3231
rect 3617 3225 3618 3231
rect 3610 3083 3618 3225
rect 3610 3077 3611 3083
rect 3617 3077 3618 3083
rect 3610 2935 3618 3077
rect 3610 2929 3611 2935
rect 3617 2929 3618 2935
rect 3610 2799 3618 2929
rect 3610 2793 3611 2799
rect 3617 2793 3618 2799
rect 3610 2651 3618 2793
rect 3610 2645 3611 2651
rect 3617 2645 3618 2651
rect 3610 2507 3618 2645
rect 3610 2501 3611 2507
rect 3617 2501 3618 2507
rect 3610 2367 3618 2501
rect 3610 2361 3611 2367
rect 3617 2361 3618 2367
rect 3610 2227 3618 2361
rect 3610 2221 3611 2227
rect 3617 2221 3618 2227
rect 3610 2079 3618 2221
rect 3610 2073 3611 2079
rect 3617 2073 3618 2079
rect 3610 1935 3618 2073
rect 3610 1929 3611 1935
rect 3617 1929 3618 1935
rect 3610 1787 3618 1929
rect 3610 1781 3611 1787
rect 3617 1781 3618 1787
rect 3610 1643 3618 1781
rect 3610 1637 3611 1643
rect 3617 1637 3618 1643
rect 3610 1499 3618 1637
rect 3610 1493 3611 1499
rect 3617 1493 3618 1499
rect 3610 1355 3618 1493
rect 3610 1349 3611 1355
rect 3617 1349 3618 1355
rect 3610 1203 3618 1349
rect 3610 1197 3611 1203
rect 3617 1197 3618 1203
rect 3610 1043 3618 1197
rect 3610 1037 3611 1043
rect 3617 1037 3618 1043
rect 3610 895 3618 1037
rect 3610 889 3611 895
rect 3617 889 3618 895
rect 3610 751 3618 889
rect 3610 745 3611 751
rect 3617 745 3618 751
rect 3610 607 3618 745
rect 3610 601 3611 607
rect 3617 601 3618 607
rect 3610 455 3618 601
rect 3610 449 3611 455
rect 3617 449 3618 455
rect 3610 319 3618 449
rect 3610 313 3611 319
rect 3617 313 3618 319
rect 3610 151 3618 313
rect 3610 145 3611 151
rect 3617 145 3618 151
rect 3610 72 3618 145
<< m6c >>
rect 570 2111 575 2115
rect 575 2111 581 2115
rect 581 2111 586 2115
rect 570 2099 586 2111
rect 1034 2109 1050 2115
rect 1034 2103 1039 2109
rect 1039 2103 1045 2109
rect 1045 2103 1050 2109
rect 1034 2099 1050 2103
<< m6 >>
rect 567 2115 1053 2118
rect 567 2099 570 2115
rect 586 2099 1034 2115
rect 1050 2099 1053 2115
rect 567 2096 1053 2099
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__191
timestamp 1731220596
transform 1 0 3568 0 -1 3576
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220596
transform 1 0 1856 0 -1 3576
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220596
transform 1 0 3568 0 1 3472
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220596
transform 1 0 1856 0 1 3472
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220596
transform 1 0 3568 0 -1 3432
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220596
transform 1 0 1856 0 -1 3432
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220596
transform 1 0 3568 0 1 3320
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220596
transform 1 0 1856 0 1 3320
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220596
transform 1 0 3568 0 -1 3288
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220596
transform 1 0 1856 0 -1 3288
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220596
transform 1 0 3568 0 1 3176
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220596
transform 1 0 1856 0 1 3176
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220596
transform 1 0 3568 0 -1 3140
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220596
transform 1 0 1856 0 -1 3140
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220596
transform 1 0 3568 0 1 3028
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220596
transform 1 0 1856 0 1 3028
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220596
transform 1 0 3568 0 -1 2992
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220596
transform 1 0 1856 0 -1 2992
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220596
transform 1 0 3568 0 1 2880
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220596
transform 1 0 1856 0 1 2880
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220596
transform 1 0 3568 0 -1 2848
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220596
transform 1 0 1856 0 -1 2848
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220596
transform 1 0 3568 0 1 2744
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220596
transform 1 0 1856 0 1 2744
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220596
transform 1 0 3568 0 -1 2708
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220596
transform 1 0 1856 0 -1 2708
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220596
transform 1 0 3568 0 1 2596
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220596
transform 1 0 1856 0 1 2596
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220596
transform 1 0 3568 0 -1 2560
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220596
transform 1 0 1856 0 -1 2560
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220596
transform 1 0 3568 0 1 2452
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220596
transform 1 0 1856 0 1 2452
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220596
transform 1 0 3568 0 -1 2420
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220596
transform 1 0 1856 0 -1 2420
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220596
transform 1 0 3568 0 1 2312
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220596
transform 1 0 1856 0 1 2312
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220596
transform 1 0 3568 0 -1 2276
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220596
transform 1 0 1856 0 -1 2276
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220596
transform 1 0 3568 0 1 2172
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220596
transform 1 0 1856 0 1 2172
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220596
transform 1 0 3568 0 -1 2132
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220596
transform 1 0 1856 0 -1 2132
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220596
transform 1 0 3568 0 1 2024
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220596
transform 1 0 1856 0 1 2024
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220596
transform 1 0 3568 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220596
transform 1 0 1856 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220596
transform 1 0 3568 0 1 1880
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220596
transform 1 0 1856 0 1 1880
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220596
transform 1 0 3568 0 -1 1840
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220596
transform 1 0 1856 0 -1 1840
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220596
transform 1 0 3568 0 1 1732
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220596
transform 1 0 1856 0 1 1732
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220596
transform 1 0 3568 0 -1 1696
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220596
transform 1 0 1856 0 -1 1696
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220596
transform 1 0 3568 0 1 1588
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220596
transform 1 0 1856 0 1 1588
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220596
transform 1 0 3568 0 -1 1556
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220596
transform 1 0 1856 0 -1 1556
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220596
transform 1 0 3568 0 1 1444
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220596
transform 1 0 1856 0 1 1444
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220596
transform 1 0 3568 0 -1 1408
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220596
transform 1 0 1856 0 -1 1408
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220596
transform 1 0 3568 0 1 1300
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220596
transform 1 0 1856 0 1 1300
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220596
transform 1 0 3568 0 -1 1256
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220596
transform 1 0 1856 0 -1 1256
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220596
transform 1 0 3568 0 1 1148
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220596
transform 1 0 1856 0 1 1148
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220596
transform 1 0 3568 0 -1 1104
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220596
transform 1 0 1856 0 -1 1104
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220596
transform 1 0 3568 0 1 988
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220596
transform 1 0 1856 0 1 988
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220596
transform 1 0 3568 0 -1 952
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220596
transform 1 0 1856 0 -1 952
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220596
transform 1 0 3568 0 1 840
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220596
transform 1 0 1856 0 1 840
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220596
transform 1 0 3568 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220596
transform 1 0 1856 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220596
transform 1 0 3568 0 1 696
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220596
transform 1 0 1856 0 1 696
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220596
transform 1 0 3568 0 -1 660
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220596
transform 1 0 1856 0 -1 660
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220596
transform 1 0 3568 0 1 552
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220596
transform 1 0 1856 0 1 552
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220596
transform 1 0 3568 0 -1 512
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220596
transform 1 0 1856 0 -1 512
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220596
transform 1 0 3568 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220596
transform 1 0 1856 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220596
transform 1 0 3568 0 -1 368
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220596
transform 1 0 1856 0 -1 368
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220596
transform 1 0 3568 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220596
transform 1 0 1856 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220596
transform 1 0 3568 0 -1 232
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220596
transform 1 0 1856 0 -1 232
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220596
transform 1 0 3568 0 1 96
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220596
transform 1 0 1856 0 1 96
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220596
transform 1 0 1816 0 -1 3652
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220596
transform 1 0 104 0 -1 3652
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220596
transform 1 0 1816 0 1 3548
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220596
transform 1 0 104 0 1 3548
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220596
transform 1 0 1816 0 -1 3516
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220596
transform 1 0 104 0 -1 3516
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220596
transform 1 0 1816 0 1 3412
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220596
transform 1 0 104 0 1 3412
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220596
transform 1 0 1816 0 -1 3380
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220596
transform 1 0 104 0 -1 3380
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220596
transform 1 0 1816 0 1 3272
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220596
transform 1 0 104 0 1 3272
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220596
transform 1 0 1816 0 -1 3236
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220596
transform 1 0 104 0 -1 3236
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220596
transform 1 0 1816 0 1 3124
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220596
transform 1 0 104 0 1 3124
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220596
transform 1 0 1816 0 -1 3084
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220596
transform 1 0 104 0 -1 3084
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220596
transform 1 0 1816 0 1 2976
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220596
transform 1 0 104 0 1 2976
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220596
transform 1 0 1816 0 -1 2944
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220596
transform 1 0 104 0 -1 2944
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220596
transform 1 0 1816 0 1 2836
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220596
transform 1 0 104 0 1 2836
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220596
transform 1 0 1816 0 -1 2796
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220596
transform 1 0 104 0 -1 2796
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220596
transform 1 0 1816 0 1 2684
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220596
transform 1 0 104 0 1 2684
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220596
transform 1 0 1816 0 -1 2648
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220596
transform 1 0 104 0 -1 2648
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220596
transform 1 0 1816 0 1 2540
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220596
transform 1 0 104 0 1 2540
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220596
transform 1 0 1816 0 -1 2508
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220596
transform 1 0 104 0 -1 2508
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220596
transform 1 0 1816 0 1 2404
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220596
transform 1 0 104 0 1 2404
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220596
transform 1 0 1816 0 -1 2360
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220596
transform 1 0 104 0 -1 2360
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220596
transform 1 0 1816 0 1 2248
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220596
transform 1 0 104 0 1 2248
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220596
transform 1 0 1816 0 -1 2208
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220596
transform 1 0 104 0 -1 2208
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220596
transform 1 0 1816 0 1 2104
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220596
transform 1 0 104 0 1 2104
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220596
transform 1 0 1816 0 -1 2068
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220596
transform 1 0 104 0 -1 2068
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220596
transform 1 0 1816 0 1 1960
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220596
transform 1 0 104 0 1 1960
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220596
transform 1 0 1816 0 -1 1924
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220596
transform 1 0 104 0 -1 1924
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220596
transform 1 0 1816 0 1 1812
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220596
transform 1 0 104 0 1 1812
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220596
transform 1 0 1816 0 -1 1768
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220596
transform 1 0 104 0 -1 1768
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220596
transform 1 0 1816 0 1 1660
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220596
transform 1 0 104 0 1 1660
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220596
transform 1 0 1816 0 -1 1620
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220596
transform 1 0 104 0 -1 1620
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220596
transform 1 0 1816 0 1 1516
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220596
transform 1 0 104 0 1 1516
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220596
transform 1 0 1816 0 -1 1480
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220596
transform 1 0 104 0 -1 1480
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220596
transform 1 0 1816 0 1 1368
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220596
transform 1 0 104 0 1 1368
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220596
transform 1 0 1816 0 -1 1332
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220596
transform 1 0 104 0 -1 1332
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220596
transform 1 0 1816 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220596
transform 1 0 104 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220596
transform 1 0 1816 0 -1 1188
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220596
transform 1 0 104 0 -1 1188
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220596
transform 1 0 1816 0 1 1084
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220596
transform 1 0 104 0 1 1084
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220596
transform 1 0 1816 0 -1 1052
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220596
transform 1 0 104 0 -1 1052
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220596
transform 1 0 1816 0 1 944
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220596
transform 1 0 104 0 1 944
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220596
transform 1 0 1816 0 -1 904
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220596
transform 1 0 104 0 -1 904
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220596
transform 1 0 1816 0 1 800
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220596
transform 1 0 104 0 1 800
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220596
transform 1 0 1816 0 -1 764
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220596
transform 1 0 104 0 -1 764
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220596
transform 1 0 1816 0 1 656
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220596
transform 1 0 104 0 1 656
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220596
transform 1 0 1816 0 -1 616
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220596
transform 1 0 104 0 -1 616
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220596
transform 1 0 1816 0 1 508
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220596
transform 1 0 104 0 1 508
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220596
transform 1 0 1816 0 -1 468
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220596
transform 1 0 104 0 -1 468
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220596
transform 1 0 1816 0 1 364
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220596
transform 1 0 104 0 1 364
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220596
transform 1 0 1816 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220596
transform 1 0 104 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220596
transform 1 0 1816 0 1 208
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220596
transform 1 0 104 0 1 208
box 7 3 12 24
use _0_0std_0_0cells_0_0MUX2X1  tst_5999_6
timestamp 1731220596
transform 1 0 3384 0 1 80
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5998_6
timestamp 1731220596
transform 1 0 3472 0 1 80
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5997_6
timestamp 1731220596
transform 1 0 3472 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5996_6
timestamp 1731220596
transform 1 0 3456 0 1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5995_6
timestamp 1731220596
transform 1 0 3424 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5994_6
timestamp 1731220596
transform 1 0 3424 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5993_6
timestamp 1731220596
transform 1 0 3352 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5992_6
timestamp 1731220596
transform 1 0 3296 0 1 80
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5991_6
timestamp 1731220596
transform 1 0 3208 0 1 80
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5990_6
timestamp 1731220596
transform 1 0 3120 0 1 80
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5989_6
timestamp 1731220596
transform 1 0 3032 0 1 80
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5988_6
timestamp 1731220596
transform 1 0 2944 0 1 80
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5987_6
timestamp 1731220596
transform 1 0 2856 0 1 80
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5986_6
timestamp 1731220596
transform 1 0 2768 0 1 80
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5985_6
timestamp 1731220596
transform 1 0 3216 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5984_6
timestamp 1731220596
transform 1 0 3080 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5983_6
timestamp 1731220596
transform 1 0 2944 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5982_6
timestamp 1731220596
transform 1 0 2808 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5981_6
timestamp 1731220596
transform 1 0 3144 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5980_6
timestamp 1731220596
transform 1 0 3024 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5979_6
timestamp 1731220596
transform 1 0 2904 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5978_6
timestamp 1731220596
transform 1 0 2792 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5977_6
timestamp 1731220596
transform 1 0 2680 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5976_6
timestamp 1731220596
transform 1 0 3224 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5975_6
timestamp 1731220596
transform 1 0 3024 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5974_6
timestamp 1731220596
transform 1 0 2840 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5973_6
timestamp 1731220596
transform 1 0 2664 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5972_6
timestamp 1731220596
transform 1 0 3224 0 1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5971_6
timestamp 1731220596
transform 1 0 2992 0 1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5970_6
timestamp 1731220596
transform 1 0 2768 0 1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5969_6
timestamp 1731220596
transform 1 0 2560 0 1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5968_6
timestamp 1731220596
transform 1 0 2368 0 1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5967_6
timestamp 1731220596
transform 1 0 3208 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5966_6
timestamp 1731220596
transform 1 0 3000 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5965_6
timestamp 1731220596
transform 1 0 2800 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5964_6
timestamp 1731220596
transform 1 0 2624 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5963_6
timestamp 1731220596
transform 1 0 2480 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5962_6
timestamp 1731220596
transform 1 0 2376 0 1 536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5961_6
timestamp 1731220596
transform 1 0 2568 0 1 536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5960_6
timestamp 1731220596
transform 1 0 3240 0 1 536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5959_6
timestamp 1731220596
transform 1 0 3008 0 1 536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5958_6
timestamp 1731220596
transform 1 0 2784 0 1 536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5957_6
timestamp 1731220596
transform 1 0 2760 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5956_6
timestamp 1731220596
transform 1 0 2608 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5955_6
timestamp 1731220596
transform 1 0 3304 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5954_6
timestamp 1731220596
transform 1 0 3112 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5953_6
timestamp 1731220596
transform 1 0 2928 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5952_6
timestamp 1731220596
transform 1 0 2784 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5951_6
timestamp 1731220596
transform 1 0 2608 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5950_6
timestamp 1731220596
transform 1 0 2960 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5949_6
timestamp 1731220596
transform 1 0 3312 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5948_6
timestamp 1731220596
transform 1 0 3136 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5947_6
timestamp 1731220596
transform 1 0 3080 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5946_6
timestamp 1731220596
transform 1 0 2936 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5945_6
timestamp 1731220596
transform 1 0 2784 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5944_6
timestamp 1731220596
transform 1 0 2824 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5943_6
timestamp 1731220596
transform 1 0 2968 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5942_6
timestamp 1731220596
transform 1 0 3104 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5941_6
timestamp 1731220596
transform 1 0 3232 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5940_6
timestamp 1731220596
transform 1 0 3360 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5939_6
timestamp 1731220596
transform 1 0 3352 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5938_6
timestamp 1731220596
transform 1 0 3216 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5937_6
timestamp 1731220596
transform 1 0 3472 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5936_6
timestamp 1731220596
transform 1 0 3472 0 1 536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5935_6
timestamp 1731220596
transform 1 0 3472 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5934_6
timestamp 1731220596
transform 1 0 3472 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5933_6
timestamp 1731220596
transform 1 0 3472 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5932_6
timestamp 1731220596
transform 1 0 3472 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5931_6
timestamp 1731220596
transform 1 0 3472 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5930_6
timestamp 1731220596
transform 1 0 3472 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5929_6
timestamp 1731220596
transform 1 0 3472 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5928_6
timestamp 1731220596
transform 1 0 3424 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5927_6
timestamp 1731220596
transform 1 0 3472 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5926_6
timestamp 1731220596
transform 1 0 3472 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5925_6
timestamp 1731220596
transform 1 0 3472 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5924_6
timestamp 1731220596
transform 1 0 3472 0 1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5923_6
timestamp 1731220596
transform 1 0 3472 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5922_6
timestamp 1731220596
transform 1 0 3424 0 -1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5921_6
timestamp 1731220596
transform 1 0 3264 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5920_6
timestamp 1731220596
transform 1 0 3152 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5919_6
timestamp 1731220596
transform 1 0 3312 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5918_6
timestamp 1731220596
transform 1 0 3312 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5917_6
timestamp 1731220596
transform 1 0 3328 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5916_6
timestamp 1731220596
transform 1 0 3360 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5915_6
timestamp 1731220596
transform 1 0 3224 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5914_6
timestamp 1731220596
transform 1 0 3088 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5913_6
timestamp 1731220596
transform 1 0 2944 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5912_6
timestamp 1731220596
transform 1 0 2792 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5911_6
timestamp 1731220596
transform 1 0 3168 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5910_6
timestamp 1731220596
transform 1 0 3008 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5909_6
timestamp 1731220596
transform 1 0 2848 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5908_6
timestamp 1731220596
transform 1 0 2680 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5907_6
timestamp 1731220596
transform 1 0 3144 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5906_6
timestamp 1731220596
transform 1 0 2984 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5905_6
timestamp 1731220596
transform 1 0 2832 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5904_6
timestamp 1731220596
transform 1 0 2680 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5903_6
timestamp 1731220596
transform 1 0 2696 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5902_6
timestamp 1731220596
transform 1 0 2848 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5901_6
timestamp 1731220596
transform 1 0 3000 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5900_6
timestamp 1731220596
transform 1 0 3224 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5899_6
timestamp 1731220596
transform 1 0 3032 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5898_6
timestamp 1731220596
transform 1 0 2848 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5897_6
timestamp 1731220596
transform 1 0 2680 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5896_6
timestamp 1731220596
transform 1 0 2544 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5895_6
timestamp 1731220596
transform 1 0 3056 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5894_6
timestamp 1731220596
transform 1 0 2856 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5893_6
timestamp 1731220596
transform 1 0 2672 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5892_6
timestamp 1731220596
transform 1 0 2496 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5891_6
timestamp 1731220596
transform 1 0 2344 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5890_6
timestamp 1731220596
transform 1 0 2432 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5889_6
timestamp 1731220596
transform 1 0 2600 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5888_6
timestamp 1731220596
transform 1 0 3256 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5887_6
timestamp 1731220596
transform 1 0 3024 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5886_6
timestamp 1731220596
transform 1 0 2800 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5885_6
timestamp 1731220596
transform 1 0 2688 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5884_6
timestamp 1731220596
transform 1 0 2520 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5883_6
timestamp 1731220596
transform 1 0 2872 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5882_6
timestamp 1731220596
transform 1 0 3280 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5881_6
timestamp 1731220596
transform 1 0 3072 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5880_6
timestamp 1731220596
transform 1 0 2944 0 -1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5879_6
timestamp 1731220596
transform 1 0 2784 0 -1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5878_6
timestamp 1731220596
transform 1 0 2616 0 -1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5877_6
timestamp 1731220596
transform 1 0 3264 0 -1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5876_6
timestamp 1731220596
transform 1 0 3104 0 -1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5875_6
timestamp 1731220596
transform 1 0 3016 0 1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5874_6
timestamp 1731220596
transform 1 0 2856 0 1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5873_6
timestamp 1731220596
transform 1 0 3176 0 1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5872_6
timestamp 1731220596
transform 1 0 3336 0 1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5871_6
timestamp 1731220596
transform 1 0 3360 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5870_6
timestamp 1731220596
transform 1 0 3240 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5869_6
timestamp 1731220596
transform 1 0 3128 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5868_6
timestamp 1731220596
transform 1 0 3008 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5867_6
timestamp 1731220596
transform 1 0 2880 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5866_6
timestamp 1731220596
transform 1 0 3160 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5865_6
timestamp 1731220596
transform 1 0 3056 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5864_6
timestamp 1731220596
transform 1 0 2952 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5863_6
timestamp 1731220596
transform 1 0 2848 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5862_6
timestamp 1731220596
transform 1 0 2744 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5861_6
timestamp 1731220596
transform 1 0 2984 0 -1 1856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5860_6
timestamp 1731220596
transform 1 0 2856 0 -1 1856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5859_6
timestamp 1731220596
transform 1 0 2736 0 -1 1856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5858_6
timestamp 1731220596
transform 1 0 2616 0 -1 1856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5857_6
timestamp 1731220596
transform 1 0 2488 0 -1 1856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5856_6
timestamp 1731220596
transform 1 0 2496 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5855_6
timestamp 1731220596
transform 1 0 2616 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5854_6
timestamp 1731220596
transform 1 0 2736 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5853_6
timestamp 1731220596
transform 1 0 2864 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5852_6
timestamp 1731220596
transform 1 0 2992 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5851_6
timestamp 1731220596
transform 1 0 2864 0 -1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5850_6
timestamp 1731220596
transform 1 0 2704 0 -1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5849_6
timestamp 1731220596
transform 1 0 3200 0 -1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5848_6
timestamp 1731220596
transform 1 0 3032 0 -1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5847_6
timestamp 1731220596
transform 1 0 2896 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5846_6
timestamp 1731220596
transform 1 0 2760 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5845_6
timestamp 1731220596
transform 1 0 2888 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5844_6
timestamp 1731220596
transform 1 0 3016 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5843_6
timestamp 1731220596
transform 1 0 3136 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5842_6
timestamp 1731220596
transform 1 0 3256 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5841_6
timestamp 1731220596
transform 1 0 3144 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5840_6
timestamp 1731220596
transform 1 0 3024 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5839_6
timestamp 1731220596
transform 1 0 3264 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5838_6
timestamp 1731220596
transform 1 0 3376 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5837_6
timestamp 1731220596
transform 1 0 3472 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5836_6
timestamp 1731220596
transform 1 0 3376 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5835_6
timestamp 1731220596
transform 1 0 3472 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5834_6
timestamp 1731220596
transform 1 0 3472 0 1 2156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5833_6
timestamp 1731220596
transform 1 0 3472 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5832_6
timestamp 1731220596
transform 1 0 3472 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5831_6
timestamp 1731220596
transform 1 0 3384 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5830_6
timestamp 1731220596
transform 1 0 3272 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5829_6
timestamp 1731220596
transform 1 0 3264 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5828_6
timestamp 1731220596
transform 1 0 3376 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5827_6
timestamp 1731220596
transform 1 0 3288 0 1 2156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5826_6
timestamp 1731220596
transform 1 0 3088 0 1 2156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5825_6
timestamp 1731220596
transform 1 0 3152 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5824_6
timestamp 1731220596
transform 1 0 3032 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5823_6
timestamp 1731220596
transform 1 0 2912 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5822_6
timestamp 1731220596
transform 1 0 2776 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5821_6
timestamp 1731220596
transform 1 0 3168 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5820_6
timestamp 1731220596
transform 1 0 3056 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5819_6
timestamp 1731220596
transform 1 0 2936 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5818_6
timestamp 1731220596
transform 1 0 2816 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5817_6
timestamp 1731220596
transform 1 0 2688 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5816_6
timestamp 1731220596
transform 1 0 3104 0 -1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5815_6
timestamp 1731220596
transform 1 0 2944 0 -1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5814_6
timestamp 1731220596
transform 1 0 2792 0 -1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5813_6
timestamp 1731220596
transform 1 0 2640 0 -1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5812_6
timestamp 1731220596
transform 1 0 3000 0 1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5811_6
timestamp 1731220596
transform 1 0 2864 0 1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5810_6
timestamp 1731220596
transform 1 0 2736 0 1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5809_6
timestamp 1731220596
transform 1 0 2608 0 1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5808_6
timestamp 1731220596
transform 1 0 2472 0 1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5807_6
timestamp 1731220596
transform 1 0 2824 0 -1 2576
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5806_6
timestamp 1731220596
transform 1 0 2704 0 -1 2576
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5805_6
timestamp 1731220596
transform 1 0 2584 0 -1 2576
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5804_6
timestamp 1731220596
transform 1 0 2464 0 -1 2576
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5803_6
timestamp 1731220596
transform 1 0 2440 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5802_6
timestamp 1731220596
transform 1 0 2536 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5801_6
timestamp 1731220596
transform 1 0 2848 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5800_6
timestamp 1731220596
transform 1 0 2744 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5799_6
timestamp 1731220596
transform 1 0 2640 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5798_6
timestamp 1731220596
transform 1 0 2616 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5797_6
timestamp 1731220596
transform 1 0 2736 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5796_6
timestamp 1731220596
transform 1 0 2856 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5795_6
timestamp 1731220596
transform 1 0 3096 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5794_6
timestamp 1731220596
transform 1 0 2976 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5793_6
timestamp 1731220596
transform 1 0 2920 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5792_6
timestamp 1731220596
transform 1 0 2768 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5791_6
timestamp 1731220596
transform 1 0 3208 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5790_6
timestamp 1731220596
transform 1 0 3064 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5789_6
timestamp 1731220596
transform 1 0 2928 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5788_6
timestamp 1731220596
transform 1 0 2800 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5787_6
timestamp 1731220596
transform 1 0 2664 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5786_6
timestamp 1731220596
transform 1 0 3048 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5785_6
timestamp 1731220596
transform 1 0 3152 0 1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5784_6
timestamp 1731220596
transform 1 0 3160 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5783_6
timestamp 1731220596
transform 1 0 3272 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5782_6
timestamp 1731220596
transform 1 0 3384 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5781_6
timestamp 1731220596
transform 1 0 3352 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5780_6
timestamp 1731220596
transform 1 0 3472 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5779_6
timestamp 1731220596
transform 1 0 3472 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5778_6
timestamp 1731220596
transform 1 0 3472 0 1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5777_6
timestamp 1731220596
transform 1 0 3472 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5776_6
timestamp 1731220596
transform 1 0 3472 0 1 3012
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5775_6
timestamp 1731220596
transform 1 0 3472 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5774_6
timestamp 1731220596
transform 1 0 3472 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5773_6
timestamp 1731220596
transform 1 0 3472 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5772_6
timestamp 1731220596
transform 1 0 3304 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5771_6
timestamp 1731220596
transform 1 0 3472 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5770_6
timestamp 1731220596
transform 1 0 3328 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5769_6
timestamp 1731220596
transform 1 0 3176 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5768_6
timestamp 1731220596
transform 1 0 3024 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5767_6
timestamp 1731220596
transform 1 0 3352 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5766_6
timestamp 1731220596
transform 1 0 3184 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5765_6
timestamp 1731220596
transform 1 0 3024 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5764_6
timestamp 1731220596
transform 1 0 2864 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5763_6
timestamp 1731220596
transform 1 0 2920 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5762_6
timestamp 1731220596
transform 1 0 3064 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5761_6
timestamp 1731220596
transform 1 0 3208 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5760_6
timestamp 1731220596
transform 1 0 3216 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5759_6
timestamp 1731220596
transform 1 0 3112 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5758_6
timestamp 1731220596
transform 1 0 3008 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5757_6
timestamp 1731220596
transform 1 0 2912 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5756_6
timestamp 1731220596
transform 1 0 2816 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5755_6
timestamp 1731220596
transform 1 0 2720 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5754_6
timestamp 1731220596
transform 1 0 2624 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5753_6
timestamp 1731220596
transform 1 0 2640 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5752_6
timestamp 1731220596
transform 1 0 2776 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5751_6
timestamp 1731220596
transform 1 0 2704 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5750_6
timestamp 1731220596
transform 1 0 2704 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5749_6
timestamp 1731220596
transform 1 0 2864 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5748_6
timestamp 1731220596
transform 1 0 2792 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5747_6
timestamp 1731220596
transform 1 0 2960 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5746_6
timestamp 1731220596
transform 1 0 3128 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5745_6
timestamp 1731220596
transform 1 0 3312 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5744_6
timestamp 1731220596
transform 1 0 3152 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5743_6
timestamp 1731220596
transform 1 0 3000 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5742_6
timestamp 1731220596
transform 1 0 2856 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5741_6
timestamp 1731220596
transform 1 0 2720 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5740_6
timestamp 1731220596
transform 1 0 2864 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5739_6
timestamp 1731220596
transform 1 0 3064 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5738_6
timestamp 1731220596
transform 1 0 3280 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5737_6
timestamp 1731220596
transform 1 0 3224 0 1 3012
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5736_6
timestamp 1731220596
transform 1 0 3312 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5735_6
timestamp 1731220596
transform 1 0 3136 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5734_6
timestamp 1731220596
transform 1 0 2960 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5733_6
timestamp 1731220596
transform 1 0 2800 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5732_6
timestamp 1731220596
transform 1 0 2656 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5731_6
timestamp 1731220596
transform 1 0 2528 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5730_6
timestamp 1731220596
transform 1 0 2408 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5729_6
timestamp 1731220596
transform 1 0 2472 0 1 3012
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5728_6
timestamp 1731220596
transform 1 0 2960 0 1 3012
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5727_6
timestamp 1731220596
transform 1 0 2704 0 1 3012
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5726_6
timestamp 1731220596
transform 1 0 2672 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5725_6
timestamp 1731220596
transform 1 0 2504 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5724_6
timestamp 1731220596
transform 1 0 2344 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5723_6
timestamp 1731220596
transform 1 0 2192 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5722_6
timestamp 1731220596
transform 1 0 2584 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5721_6
timestamp 1731220596
transform 1 0 2448 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5720_6
timestamp 1731220596
transform 1 0 2312 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5719_6
timestamp 1731220596
transform 1 0 2160 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5718_6
timestamp 1731220596
transform 1 0 2624 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5717_6
timestamp 1731220596
transform 1 0 2456 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5716_6
timestamp 1731220596
transform 1 0 2296 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5715_6
timestamp 1731220596
transform 1 0 2144 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5714_6
timestamp 1731220596
transform 1 0 2536 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5713_6
timestamp 1731220596
transform 1 0 2360 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5712_6
timestamp 1731220596
transform 1 0 2184 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5711_6
timestamp 1731220596
transform 1 0 2016 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5710_6
timestamp 1731220596
transform 1 0 2184 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5709_6
timestamp 1731220596
transform 1 0 2360 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5708_6
timestamp 1731220596
transform 1 0 2536 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5707_6
timestamp 1731220596
transform 1 0 2496 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5706_6
timestamp 1731220596
transform 1 0 2352 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5705_6
timestamp 1731220596
transform 1 0 2216 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5704_6
timestamp 1731220596
transform 1 0 2088 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5703_6
timestamp 1731220596
transform 1 0 2528 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5702_6
timestamp 1731220596
transform 1 0 2424 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5701_6
timestamp 1731220596
transform 1 0 2320 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5700_6
timestamp 1731220596
transform 1 0 2232 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5699_6
timestamp 1731220596
transform 1 0 2144 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5698_6
timestamp 1731220596
transform 1 0 2056 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5697_6
timestamp 1731220596
transform 1 0 1968 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5696_6
timestamp 1731220596
transform 1 0 1880 0 -1 3592
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5695_6
timestamp 1731220596
transform 1 0 1880 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5694_6
timestamp 1731220596
transform 1 0 1968 0 1 3456
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5693_6
timestamp 1731220596
transform 1 0 2016 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5692_6
timestamp 1731220596
transform 1 0 1880 0 -1 3448
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5691_6
timestamp 1731220596
transform 1 0 1880 0 1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5690_6
timestamp 1731220596
transform 1 0 1880 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5689_6
timestamp 1731220596
transform 1 0 2000 0 -1 3304
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5688_6
timestamp 1731220596
transform 1 0 1880 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5687_6
timestamp 1731220596
transform 1 0 2008 0 1 3160
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5686_6
timestamp 1731220596
transform 1 0 2040 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5685_6
timestamp 1731220596
transform 1 0 1880 0 -1 3156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5684_6
timestamp 1731220596
transform 1 0 1904 0 1 3012
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5683_6
timestamp 1731220596
transform 1 0 2072 0 1 3012
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5682_6
timestamp 1731220596
transform 1 0 2264 0 1 3012
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5681_6
timestamp 1731220596
transform 1 0 2280 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5680_6
timestamp 1731220596
transform 1 0 2152 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5679_6
timestamp 1731220596
transform 1 0 2016 0 -1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5678_6
timestamp 1731220596
transform 1 0 2160 0 1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5677_6
timestamp 1731220596
transform 1 0 2480 0 1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5676_6
timestamp 1731220596
transform 1 0 2808 0 1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5675_6
timestamp 1731220596
transform 1 0 2512 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5674_6
timestamp 1731220596
transform 1 0 2352 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5673_6
timestamp 1731220596
transform 1 0 2184 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5672_6
timestamp 1731220596
transform 1 0 2240 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5671_6
timestamp 1731220596
transform 1 0 2424 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5670_6
timestamp 1731220596
transform 1 0 2600 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5669_6
timestamp 1731220596
transform 1 0 2488 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5668_6
timestamp 1731220596
transform 1 0 2352 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5667_6
timestamp 1731220596
transform 1 0 2200 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5666_6
timestamp 1731220596
transform 1 0 2336 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5665_6
timestamp 1731220596
transform 1 0 2224 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5664_6
timestamp 1731220596
transform 1 0 2104 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5663_6
timestamp 1731220596
transform 1 0 2104 0 -1 2576
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5662_6
timestamp 1731220596
transform 1 0 2224 0 -1 2576
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5661_6
timestamp 1731220596
transform 1 0 2344 0 -1 2576
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5660_6
timestamp 1731220596
transform 1 0 2328 0 1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5659_6
timestamp 1731220596
transform 1 0 2176 0 1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5658_6
timestamp 1731220596
transform 1 0 2168 0 -1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5657_6
timestamp 1731220596
transform 1 0 2328 0 -1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5656_6
timestamp 1731220596
transform 1 0 2488 0 -1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5655_6
timestamp 1731220596
transform 1 0 2392 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5654_6
timestamp 1731220596
transform 1 0 2232 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5653_6
timestamp 1731220596
transform 1 0 2544 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5652_6
timestamp 1731220596
transform 1 0 2632 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5651_6
timestamp 1731220596
transform 1 0 2472 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5650_6
timestamp 1731220596
transform 1 0 2304 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5649_6
timestamp 1731220596
transform 1 0 2504 0 1 2156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5648_6
timestamp 1731220596
transform 1 0 2696 0 1 2156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5647_6
timestamp 1731220596
transform 1 0 2888 0 1 2156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5646_6
timestamp 1731220596
transform 1 0 2752 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5645_6
timestamp 1731220596
transform 1 0 2608 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5644_6
timestamp 1731220596
transform 1 0 2464 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5643_6
timestamp 1731220596
transform 1 0 2312 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5642_6
timestamp 1731220596
transform 1 0 2296 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5641_6
timestamp 1731220596
transform 1 0 2456 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5640_6
timestamp 1731220596
transform 1 0 2616 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5639_6
timestamp 1731220596
transform 1 0 2536 0 -1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5638_6
timestamp 1731220596
transform 1 0 2368 0 -1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5637_6
timestamp 1731220596
transform 1 0 2240 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5636_6
timestamp 1731220596
transform 1 0 2368 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5635_6
timestamp 1731220596
transform 1 0 2352 0 -1 1856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5634_6
timestamp 1731220596
transform 1 0 2216 0 -1 1856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5633_6
timestamp 1731220596
transform 1 0 2256 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5632_6
timestamp 1731220596
transform 1 0 2344 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5631_6
timestamp 1731220596
transform 1 0 2440 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5630_6
timestamp 1731220596
transform 1 0 2544 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5629_6
timestamp 1731220596
transform 1 0 2648 0 1 1716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5628_6
timestamp 1731220596
transform 1 0 2752 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5627_6
timestamp 1731220596
transform 1 0 2616 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5626_6
timestamp 1731220596
transform 1 0 2488 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5625_6
timestamp 1731220596
transform 1 0 2360 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5624_6
timestamp 1731220596
transform 1 0 2240 0 -1 1712
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5623_6
timestamp 1731220596
transform 1 0 2688 0 1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5622_6
timestamp 1731220596
transform 1 0 2512 0 1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5621_6
timestamp 1731220596
transform 1 0 2328 0 1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5620_6
timestamp 1731220596
transform 1 0 2136 0 1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5619_6
timestamp 1731220596
transform 1 0 2080 0 -1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5618_6
timestamp 1731220596
transform 1 0 2448 0 -1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5617_6
timestamp 1731220596
transform 1 0 2272 0 -1 1572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5616_6
timestamp 1731220596
transform 1 0 2104 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5615_6
timestamp 1731220596
transform 1 0 2232 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5614_6
timestamp 1731220596
transform 1 0 2368 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5613_6
timestamp 1731220596
transform 1 0 2296 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5612_6
timestamp 1731220596
transform 1 0 2176 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5611_6
timestamp 1731220596
transform 1 0 2208 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5610_6
timestamp 1731220596
transform 1 0 2088 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5609_6
timestamp 1731220596
transform 1 0 1968 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5608_6
timestamp 1731220596
transform 1 0 1880 0 1 1284
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5607_6
timestamp 1731220596
transform 1 0 1880 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5606_6
timestamp 1731220596
transform 1 0 1968 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5605_6
timestamp 1731220596
transform 1 0 2064 0 -1 1424
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5604_6
timestamp 1731220596
transform 1 0 1976 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5603_6
timestamp 1731220596
transform 1 0 1880 0 1 1428
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5602_6
timestamp 1731220596
transform 1 0 1720 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5601_6
timestamp 1731220596
transform 1 0 1576 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5600_6
timestamp 1731220596
transform 1 0 1448 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5599_6
timestamp 1731220596
transform 1 0 1592 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5598_6
timestamp 1731220596
transform 1 0 1720 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5597_6
timestamp 1731220596
transform 1 0 1680 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5596_6
timestamp 1731220596
transform 1 0 1696 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5595_6
timestamp 1731220596
transform 1 0 1368 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5594_6
timestamp 1731220596
transform 1 0 1344 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5593_6
timestamp 1731220596
transform 1 0 1248 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5592_6
timestamp 1731220596
transform 1 0 1440 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5591_6
timestamp 1731220596
transform 1 0 1456 0 -1 1940
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5590_6
timestamp 1731220596
transform 1 0 1144 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5589_6
timestamp 1731220596
transform 1 0 1040 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5588_6
timestamp 1731220596
transform 1 0 1208 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5587_6
timestamp 1731220596
transform 1 0 1040 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5586_6
timestamp 1731220596
transform 1 0 1008 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5585_6
timestamp 1731220596
transform 1 0 984 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5584_6
timestamp 1731220596
transform 1 0 1088 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5583_6
timestamp 1731220596
transform 1 0 920 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5582_6
timestamp 1731220596
transform 1 0 864 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5581_6
timestamp 1731220596
transform 1 0 984 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5580_6
timestamp 1731220596
transform 1 0 1112 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5579_6
timestamp 1731220596
transform 1 0 1104 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5578_6
timestamp 1731220596
transform 1 0 1000 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5577_6
timestamp 1731220596
transform 1 0 904 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5576_6
timestamp 1731220596
transform 1 0 800 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5575_6
timestamp 1731220596
transform 1 0 696 0 -1 1348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5574_6
timestamp 1731220596
transform 1 0 568 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5573_6
timestamp 1731220596
transform 1 0 448 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5572_6
timestamp 1731220596
transform 1 0 688 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5571_6
timestamp 1731220596
transform 1 0 736 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5570_6
timestamp 1731220596
transform 1 0 600 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5569_6
timestamp 1731220596
transform 1 0 464 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5568_6
timestamp 1731220596
transform 1 0 320 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5567_6
timestamp 1731220596
transform 1 0 416 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5566_6
timestamp 1731220596
transform 1 0 584 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5565_6
timestamp 1731220596
transform 1 0 752 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5564_6
timestamp 1731220596
transform 1 0 808 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5563_6
timestamp 1731220596
transform 1 0 624 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5562_6
timestamp 1731220596
transform 1 0 440 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5561_6
timestamp 1731220596
transform 1 0 264 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5560_6
timestamp 1731220596
transform 1 0 272 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5559_6
timestamp 1731220596
transform 1 0 456 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5558_6
timestamp 1731220596
transform 1 0 640 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5557_6
timestamp 1731220596
transform 1 0 824 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5556_6
timestamp 1731220596
transform 1 0 864 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5555_6
timestamp 1731220596
transform 1 0 680 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5554_6
timestamp 1731220596
transform 1 0 488 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5553_6
timestamp 1731220596
transform 1 0 544 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5552_6
timestamp 1731220596
transform 1 0 680 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5551_6
timestamp 1731220596
transform 1 0 808 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5550_6
timestamp 1731220596
transform 1 0 928 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5549_6
timestamp 1731220596
transform 1 0 1240 0 -1 1940
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5548_6
timestamp 1731220596
transform 1 0 1032 0 -1 1940
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5547_6
timestamp 1731220596
transform 1 0 832 0 -1 1940
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5546_6
timestamp 1731220596
transform 1 0 760 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5545_6
timestamp 1731220596
transform 1 0 880 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5544_6
timestamp 1731220596
transform 1 0 1000 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5543_6
timestamp 1731220596
transform 1 0 1240 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5542_6
timestamp 1731220596
transform 1 0 1120 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5541_6
timestamp 1731220596
transform 1 0 1032 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5540_6
timestamp 1731220596
transform 1 0 912 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5539_6
timestamp 1731220596
transform 1 0 1152 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5538_6
timestamp 1731220596
transform 1 0 1272 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5537_6
timestamp 1731220596
transform 1 0 1400 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5536_6
timestamp 1731220596
transform 1 0 1312 0 1 2088
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5535_6
timestamp 1731220596
transform 1 0 1168 0 1 2088
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5534_6
timestamp 1731220596
transform 1 0 1456 0 1 2088
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5533_6
timestamp 1731220596
transform 1 0 1608 0 1 2088
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5532_6
timestamp 1731220596
transform 1 0 1720 0 -1 2224
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5531_6
timestamp 1731220596
transform 1 0 1568 0 -1 2224
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5530_6
timestamp 1731220596
transform 1 0 1400 0 -1 2224
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5529_6
timestamp 1731220596
transform 1 0 1232 0 -1 2224
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5528_6
timestamp 1731220596
transform 1 0 1720 0 1 2232
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5527_6
timestamp 1731220596
transform 1 0 1584 0 1 2232
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5526_6
timestamp 1731220596
transform 1 0 1448 0 1 2232
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5525_6
timestamp 1731220596
transform 1 0 1304 0 1 2232
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5524_6
timestamp 1731220596
transform 1 0 1160 0 1 2232
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5523_6
timestamp 1731220596
transform 1 0 1576 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5522_6
timestamp 1731220596
transform 1 0 1448 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5521_6
timestamp 1731220596
transform 1 0 1320 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5520_6
timestamp 1731220596
transform 1 0 1200 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5519_6
timestamp 1731220596
transform 1 0 1072 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5518_6
timestamp 1731220596
transform 1 0 1392 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5517_6
timestamp 1731220596
transform 1 0 1256 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5516_6
timestamp 1731220596
transform 1 0 1120 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5515_6
timestamp 1731220596
transform 1 0 984 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5514_6
timestamp 1731220596
transform 1 0 1272 0 -1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5513_6
timestamp 1731220596
transform 1 0 1136 0 -1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5512_6
timestamp 1731220596
transform 1 0 1000 0 -1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5511_6
timestamp 1731220596
transform 1 0 864 0 -1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5510_6
timestamp 1731220596
transform 1 0 912 0 1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5509_6
timestamp 1731220596
transform 1 0 1032 0 1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5508_6
timestamp 1731220596
transform 1 0 1160 0 1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5507_6
timestamp 1731220596
transform 1 0 1304 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5506_6
timestamp 1731220596
transform 1 0 1200 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5505_6
timestamp 1731220596
transform 1 0 1096 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5504_6
timestamp 1731220596
transform 1 0 992 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5503_6
timestamp 1731220596
transform 1 0 896 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5502_6
timestamp 1731220596
transform 1 0 792 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5501_6
timestamp 1731220596
transform 1 0 688 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5500_6
timestamp 1731220596
transform 1 0 792 0 1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5499_6
timestamp 1731220596
transform 1 0 728 0 -1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5498_6
timestamp 1731220596
transform 1 0 848 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5497_6
timestamp 1731220596
transform 1 0 944 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5496_6
timestamp 1731220596
transform 1 0 848 0 1 2232
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5495_6
timestamp 1731220596
transform 1 0 680 0 1 2232
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5494_6
timestamp 1731220596
transform 1 0 1008 0 1 2232
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5493_6
timestamp 1731220596
transform 1 0 1064 0 -1 2224
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5492_6
timestamp 1731220596
transform 1 0 888 0 -1 2224
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5491_6
timestamp 1731220596
transform 1 0 712 0 -1 2224
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5490_6
timestamp 1731220596
transform 1 0 528 0 -1 2224
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5489_6
timestamp 1731220596
transform 1 0 1024 0 1 2088
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5488_6
timestamp 1731220596
transform 1 0 880 0 1 2088
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5487_6
timestamp 1731220596
transform 1 0 744 0 1 2088
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5486_6
timestamp 1731220596
transform 1 0 608 0 1 2088
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5485_6
timestamp 1731220596
transform 1 0 480 0 1 2088
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5484_6
timestamp 1731220596
transform 1 0 792 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5483_6
timestamp 1731220596
transform 1 0 672 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5482_6
timestamp 1731220596
transform 1 0 544 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5481_6
timestamp 1731220596
transform 1 0 424 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5480_6
timestamp 1731220596
transform 1 0 312 0 -1 2084
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5479_6
timestamp 1731220596
transform 1 0 640 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5478_6
timestamp 1731220596
transform 1 0 520 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5477_6
timestamp 1731220596
transform 1 0 400 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5476_6
timestamp 1731220596
transform 1 0 280 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5475_6
timestamp 1731220596
transform 1 0 168 0 1 1944
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5474_6
timestamp 1731220596
transform 1 0 648 0 -1 1940
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5473_6
timestamp 1731220596
transform 1 0 488 0 -1 1940
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5472_6
timestamp 1731220596
transform 1 0 344 0 -1 1940
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5471_6
timestamp 1731220596
transform 1 0 216 0 -1 1940
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5470_6
timestamp 1731220596
transform 1 0 128 0 -1 1940
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5469_6
timestamp 1731220596
transform 1 0 128 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5468_6
timestamp 1731220596
transform 1 0 256 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5467_6
timestamp 1731220596
transform 1 0 400 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5466_6
timestamp 1731220596
transform 1 0 296 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5465_6
timestamp 1731220596
transform 1 0 128 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5464_6
timestamp 1731220596
transform 1 0 128 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5463_6
timestamp 1731220596
transform 1 0 128 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5462_6
timestamp 1731220596
transform 1 0 128 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5461_6
timestamp 1731220596
transform 1 0 256 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5460_6
timestamp 1731220596
transform 1 0 176 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5459_6
timestamp 1731220596
transform 1 0 184 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5458_6
timestamp 1731220596
transform 1 0 320 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5457_6
timestamp 1731220596
transform 1 0 224 0 -1 1348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5456_6
timestamp 1731220596
transform 1 0 376 0 -1 1348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5455_6
timestamp 1731220596
transform 1 0 536 0 -1 1348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5454_6
timestamp 1731220596
transform 1 0 864 0 -1 1348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5453_6
timestamp 1731220596
transform 1 0 824 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5452_6
timestamp 1731220596
transform 1 0 664 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5451_6
timestamp 1731220596
transform 1 0 504 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5450_6
timestamp 1731220596
transform 1 0 344 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5449_6
timestamp 1731220596
transform 1 0 200 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5448_6
timestamp 1731220596
transform 1 0 128 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5447_6
timestamp 1731220596
transform 1 0 264 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5446_6
timestamp 1731220596
transform 1 0 416 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5445_6
timestamp 1731220596
transform 1 0 280 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5444_6
timestamp 1731220596
transform 1 0 128 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5443_6
timestamp 1731220596
transform 1 0 128 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5442_6
timestamp 1731220596
transform 1 0 272 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5441_6
timestamp 1731220596
transform 1 0 128 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5440_6
timestamp 1731220596
transform 1 0 128 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5439_6
timestamp 1731220596
transform 1 0 264 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5438_6
timestamp 1731220596
transform 1 0 128 0 1 784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5437_6
timestamp 1731220596
transform 1 0 128 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5436_6
timestamp 1731220596
transform 1 0 264 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5435_6
timestamp 1731220596
transform 1 0 272 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5434_6
timestamp 1731220596
transform 1 0 128 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5433_6
timestamp 1731220596
transform 1 0 128 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5432_6
timestamp 1731220596
transform 1 0 280 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5431_6
timestamp 1731220596
transform 1 0 296 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5430_6
timestamp 1731220596
transform 1 0 136 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5429_6
timestamp 1731220596
transform 1 0 152 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5428_6
timestamp 1731220596
transform 1 0 304 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5427_6
timestamp 1731220596
transform 1 0 256 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5426_6
timestamp 1731220596
transform 1 0 136 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5425_6
timestamp 1731220596
transform 1 0 392 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5424_6
timestamp 1731220596
transform 1 0 392 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5423_6
timestamp 1731220596
transform 1 0 304 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5422_6
timestamp 1731220596
transform 1 0 216 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5421_6
timestamp 1731220596
transform 1 0 128 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5420_6
timestamp 1731220596
transform 1 0 128 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5419_6
timestamp 1731220596
transform 1 0 216 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5418_6
timestamp 1731220596
transform 1 0 304 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5417_6
timestamp 1731220596
transform 1 0 392 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5416_6
timestamp 1731220596
transform 1 0 480 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5415_6
timestamp 1731220596
transform 1 0 568 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5414_6
timestamp 1731220596
transform 1 0 656 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5413_6
timestamp 1731220596
transform 1 0 920 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5412_6
timestamp 1731220596
transform 1 0 832 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5411_6
timestamp 1731220596
transform 1 0 744 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5410_6
timestamp 1731220596
transform 1 0 656 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5409_6
timestamp 1731220596
transform 1 0 568 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5408_6
timestamp 1731220596
transform 1 0 480 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5407_6
timestamp 1731220596
transform 1 0 744 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5406_6
timestamp 1731220596
transform 1 0 832 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5405_6
timestamp 1731220596
transform 1 0 872 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5404_6
timestamp 1731220596
transform 1 0 696 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5403_6
timestamp 1731220596
transform 1 0 536 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5402_6
timestamp 1731220596
transform 1 0 456 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5401_6
timestamp 1731220596
transform 1 0 608 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5400_6
timestamp 1731220596
transform 1 0 752 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5399_6
timestamp 1731220596
transform 1 0 768 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5398_6
timestamp 1731220596
transform 1 0 616 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5397_6
timestamp 1731220596
transform 1 0 456 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5396_6
timestamp 1731220596
transform 1 0 448 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5395_6
timestamp 1731220596
transform 1 0 624 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5394_6
timestamp 1731220596
transform 1 0 792 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5393_6
timestamp 1731220596
transform 1 0 776 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5392_6
timestamp 1731220596
transform 1 0 608 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5391_6
timestamp 1731220596
transform 1 0 440 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5390_6
timestamp 1731220596
transform 1 0 432 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5389_6
timestamp 1731220596
transform 1 0 600 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5388_6
timestamp 1731220596
transform 1 0 768 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5387_6
timestamp 1731220596
transform 1 0 792 0 1 784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5386_6
timestamp 1731220596
transform 1 0 624 0 1 784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5385_6
timestamp 1731220596
transform 1 0 448 0 1 784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5384_6
timestamp 1731220596
transform 1 0 272 0 1 784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5383_6
timestamp 1731220596
transform 1 0 432 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5382_6
timestamp 1731220596
transform 1 0 768 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5381_6
timestamp 1731220596
transform 1 0 600 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5380_6
timestamp 1731220596
transform 1 0 448 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5379_6
timestamp 1731220596
transform 1 0 632 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5378_6
timestamp 1731220596
transform 1 0 808 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5377_6
timestamp 1731220596
transform 1 0 728 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5376_6
timestamp 1731220596
transform 1 0 576 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5375_6
timestamp 1731220596
transform 1 0 424 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5374_6
timestamp 1731220596
transform 1 0 264 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5373_6
timestamp 1731220596
transform 1 0 464 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5372_6
timestamp 1731220596
transform 1 0 832 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5371_6
timestamp 1731220596
transform 1 0 648 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5370_6
timestamp 1731220596
transform 1 0 568 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5369_6
timestamp 1731220596
transform 1 0 720 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5368_6
timestamp 1731220596
transform 1 0 880 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5367_6
timestamp 1731220596
transform 1 0 1048 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5366_6
timestamp 1731220596
transform 1 0 1224 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5365_6
timestamp 1731220596
transform 1 0 1192 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5364_6
timestamp 1731220596
transform 1 0 1016 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5363_6
timestamp 1731220596
transform 1 0 880 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5362_6
timestamp 1731220596
transform 1 0 1040 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5361_6
timestamp 1731220596
transform 1 0 1376 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5360_6
timestamp 1731220596
transform 1 0 1208 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5359_6
timestamp 1731220596
transform 1 0 1152 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5358_6
timestamp 1731220596
transform 1 0 984 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5357_6
timestamp 1731220596
transform 1 0 928 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5356_6
timestamp 1731220596
transform 1 0 1088 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5355_6
timestamp 1731220596
transform 1 0 968 0 1 784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5354_6
timestamp 1731220596
transform 1 0 1144 0 1 784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5353_6
timestamp 1731220596
transform 1 0 1080 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5352_6
timestamp 1731220596
transform 1 0 928 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5351_6
timestamp 1731220596
transform 1 0 944 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5350_6
timestamp 1731220596
transform 1 0 1104 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5349_6
timestamp 1731220596
transform 1 0 1112 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5348_6
timestamp 1731220596
transform 1 0 960 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5347_6
timestamp 1731220596
transform 1 0 912 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5346_6
timestamp 1731220596
transform 1 0 1048 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5345_6
timestamp 1731220596
transform 1 0 1000 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5344_6
timestamp 1731220596
transform 1 0 880 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5343_6
timestamp 1731220596
transform 1 0 1232 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5342_6
timestamp 1731220596
transform 1 0 1048 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5341_6
timestamp 1731220596
transform 1 0 1008 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5340_6
timestamp 1731220596
transform 1 0 920 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5339_6
timestamp 1731220596
transform 1 0 1096 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5338_6
timestamp 1731220596
transform 1 0 1184 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5337_6
timestamp 1731220596
transform 1 0 1184 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5336_6
timestamp 1731220596
transform 1 0 1096 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5335_6
timestamp 1731220596
transform 1 0 1008 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5334_6
timestamp 1731220596
transform 1 0 1272 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5333_6
timestamp 1731220596
transform 1 0 1360 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5332_6
timestamp 1731220596
transform 1 0 1448 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5331_6
timestamp 1731220596
transform 1 0 1712 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5330_6
timestamp 1731220596
transform 1 0 1624 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5329_6
timestamp 1731220596
transform 1 0 1536 0 1 192
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5328_6
timestamp 1731220596
transform 1 0 1472 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5327_6
timestamp 1731220596
transform 1 0 1376 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5326_6
timestamp 1731220596
transform 1 0 1280 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5325_6
timestamp 1731220596
transform 1 0 1568 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5324_6
timestamp 1731220596
transform 1 0 1664 0 -1 332
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5323_6
timestamp 1731220596
transform 1 0 1624 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5322_6
timestamp 1731220596
transform 1 0 1424 0 1 348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5321_6
timestamp 1731220596
transform 1 0 1336 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5320_6
timestamp 1731220596
transform 1 0 1232 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5319_6
timestamp 1731220596
transform 1 0 1120 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5318_6
timestamp 1731220596
transform 1 0 1520 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5317_6
timestamp 1731220596
transform 1 0 1632 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5316_6
timestamp 1731220596
transform 1 0 1720 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5315_6
timestamp 1731220596
transform 1 0 1880 0 1 536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5314_6
timestamp 1731220596
transform 1 0 1880 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5313_6
timestamp 1731220596
transform 1 0 1968 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5312_6
timestamp 1731220596
transform 1 0 2088 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5311_6
timestamp 1731220596
transform 1 0 2056 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5310_6
timestamp 1731220596
transform 1 0 1880 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5309_6
timestamp 1731220596
transform 1 0 2064 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5308_6
timestamp 1731220596
transform 1 0 1880 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5307_6
timestamp 1731220596
transform 1 0 1880 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5306_6
timestamp 1731220596
transform 1 0 2008 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5305_6
timestamp 1731220596
transform 1 0 2168 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5304_6
timestamp 1731220596
transform 1 0 2064 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5303_6
timestamp 1731220596
transform 1 0 1880 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5302_6
timestamp 1731220596
transform 1 0 1904 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5301_6
timestamp 1731220596
transform 1 0 2112 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5300_6
timestamp 1731220596
transform 1 0 2224 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5299_6
timestamp 1731220596
transform 1 0 2080 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5298_6
timestamp 1731220596
transform 1 0 1936 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5297_6
timestamp 1731220596
transform 1 0 2024 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5296_6
timestamp 1731220596
transform 1 0 2264 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5295_6
timestamp 1731220596
transform 1 0 2136 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5294_6
timestamp 1731220596
transform 1 0 2048 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5293_6
timestamp 1731220596
transform 1 0 2136 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5292_6
timestamp 1731220596
transform 1 0 2232 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5291_6
timestamp 1731220596
transform 1 0 2328 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5290_6
timestamp 1731220596
transform 1 0 2424 0 -1 1272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5289_6
timestamp 1731220596
transform 1 0 2400 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5288_6
timestamp 1731220596
transform 1 0 2544 0 1 1132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5287_6
timestamp 1731220596
transform 1 0 2528 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5286_6
timestamp 1731220596
transform 1 0 2376 0 -1 1120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5285_6
timestamp 1731220596
transform 1 0 2312 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5284_6
timestamp 1731220596
transform 1 0 2504 0 1 972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5283_6
timestamp 1731220596
transform 1 0 2624 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5282_6
timestamp 1731220596
transform 1 0 2448 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5281_6
timestamp 1731220596
transform 1 0 2256 0 -1 968
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5280_6
timestamp 1731220596
transform 1 0 2336 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5279_6
timestamp 1731220596
transform 1 0 2504 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5278_6
timestamp 1731220596
transform 1 0 2672 0 1 824
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5277_6
timestamp 1731220596
transform 1 0 2616 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5276_6
timestamp 1731220596
transform 1 0 2440 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5275_6
timestamp 1731220596
transform 1 0 2256 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5274_6
timestamp 1731220596
transform 1 0 2248 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5273_6
timestamp 1731220596
transform 1 0 2432 0 1 680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5272_6
timestamp 1731220596
transform 1 0 2472 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5271_6
timestamp 1731220596
transform 1 0 2344 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5270_6
timestamp 1731220596
transform 1 0 2216 0 -1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5269_6
timestamp 1731220596
transform 1 0 2200 0 1 536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5268_6
timestamp 1731220596
transform 1 0 2032 0 1 536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5267_6
timestamp 1731220596
transform 1 0 2368 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5266_6
timestamp 1731220596
transform 1 0 2272 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5265_6
timestamp 1731220596
transform 1 0 2184 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5264_6
timestamp 1731220596
transform 1 0 2024 0 1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5263_6
timestamp 1731220596
transform 1 0 2192 0 1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5262_6
timestamp 1731220596
transform 1 0 2256 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5261_6
timestamp 1731220596
transform 1 0 2376 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5260_6
timestamp 1731220596
transform 1 0 2512 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5259_6
timestamp 1731220596
transform 1 0 2456 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5258_6
timestamp 1731220596
transform 1 0 2344 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5257_6
timestamp 1731220596
transform 1 0 2568 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5256_6
timestamp 1731220596
transform 1 0 2672 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5255_6
timestamp 1731220596
transform 1 0 2528 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5254_6
timestamp 1731220596
transform 1 0 2392 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5253_6
timestamp 1731220596
transform 1 0 2256 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5252_6
timestamp 1731220596
transform 1 0 2144 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5251_6
timestamp 1731220596
transform 1 0 2056 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5250_6
timestamp 1731220596
transform 1 0 1968 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5249_6
timestamp 1731220596
transform 1 0 1880 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5248_6
timestamp 1731220596
transform 1 0 2232 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5247_6
timestamp 1731220596
transform 1 0 2144 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5246_6
timestamp 1731220596
transform 1 0 2056 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5245_6
timestamp 1731220596
transform 1 0 1968 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5244_6
timestamp 1731220596
transform 1 0 1880 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5243_6
timestamp 1731220596
transform 1 0 2144 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5242_6
timestamp 1731220596
transform 1 0 2056 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5241_6
timestamp 1731220596
transform 1 0 1968 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5240_6
timestamp 1731220596
transform 1 0 1880 0 -1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5239_6
timestamp 1731220596
transform 1 0 1880 0 1 384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5238_6
timestamp 1731220596
transform 1 0 1720 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5237_6
timestamp 1731220596
transform 1 0 1632 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5236_6
timestamp 1731220596
transform 1 0 1536 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5235_6
timestamp 1731220596
transform 1 0 1432 0 -1 484
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5234_6
timestamp 1731220596
transform 1 0 1408 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5233_6
timestamp 1731220596
transform 1 0 1296 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5232_6
timestamp 1731220596
transform 1 0 1176 0 1 492
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5231_6
timestamp 1731220596
transform 1 0 1704 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5230_6
timestamp 1731220596
transform 1 0 1552 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5229_6
timestamp 1731220596
transform 1 0 1408 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5228_6
timestamp 1731220596
transform 1 0 1264 0 -1 632
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5227_6
timestamp 1731220596
transform 1 0 1264 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5226_6
timestamp 1731220596
transform 1 0 1424 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5225_6
timestamp 1731220596
transform 1 0 1584 0 1 640
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5224_6
timestamp 1731220596
transform 1 0 1544 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5223_6
timestamp 1731220596
transform 1 0 1384 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5222_6
timestamp 1731220596
transform 1 0 1232 0 -1 780
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5221_6
timestamp 1731220596
transform 1 0 1320 0 1 784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5220_6
timestamp 1731220596
transform 1 0 1496 0 1 784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5219_6
timestamp 1731220596
transform 1 0 1392 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5218_6
timestamp 1731220596
transform 1 0 1240 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5217_6
timestamp 1731220596
transform 1 0 1544 0 -1 920
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5216_6
timestamp 1731220596
transform 1 0 1472 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5215_6
timestamp 1731220596
transform 1 0 1312 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5214_6
timestamp 1731220596
transform 1 0 1640 0 1 928
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5213_6
timestamp 1731220596
transform 1 0 1552 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5212_6
timestamp 1731220596
transform 1 0 1720 0 -1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5211_6
timestamp 1731220596
transform 1 0 1720 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5210_6
timestamp 1731220596
transform 1 0 1560 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5209_6
timestamp 1731220596
transform 1 0 1376 0 1 1068
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5208_6
timestamp 1731220596
transform 1 0 1408 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5207_6
timestamp 1731220596
transform 1 0 1592 0 -1 1204
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5206_6
timestamp 1731220596
transform 1 0 1576 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5205_6
timestamp 1731220596
transform 1 0 1424 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5204_6
timestamp 1731220596
transform 1 0 1280 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5203_6
timestamp 1731220596
transform 1 0 1136 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5202_6
timestamp 1731220596
transform 1 0 984 0 1 1212
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5201_6
timestamp 1731220596
transform 1 0 1032 0 -1 1348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5200_6
timestamp 1731220596
transform 1 0 1200 0 -1 1348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5199_6
timestamp 1731220596
transform 1 0 1368 0 -1 1348
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5198_6
timestamp 1731220596
transform 1 0 1312 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5197_6
timestamp 1731220596
transform 1 0 1208 0 1 1352
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5196_6
timestamp 1731220596
transform 1 0 1240 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5195_6
timestamp 1731220596
transform 1 0 1368 0 -1 1496
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5194_6
timestamp 1731220596
transform 1 0 1408 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5193_6
timestamp 1731220596
transform 1 0 1248 0 1 1500
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5192_6
timestamp 1731220596
transform 1 0 1296 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5191_6
timestamp 1731220596
transform 1 0 1144 0 -1 1636
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5190_6
timestamp 1731220596
transform 1 0 1176 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5189_6
timestamp 1731220596
transform 1 0 1344 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5188_6
timestamp 1731220596
transform 1 0 1512 0 1 1644
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5187_6
timestamp 1731220596
transform 1 0 1528 0 -1 1784
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5186_6
timestamp 1731220596
transform 1 0 1536 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5185_6
timestamp 1731220596
transform 1 0 1632 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5184_6
timestamp 1731220596
transform 1 0 1720 0 1 1796
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5183_6
timestamp 1731220596
transform 1 0 1880 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5182_6
timestamp 1731220596
transform 1 0 2104 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5181_6
timestamp 1731220596
transform 1 0 1976 0 1 1864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5180_6
timestamp 1731220596
transform 1 0 1880 0 -1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5179_6
timestamp 1731220596
transform 1 0 2024 0 -1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5178_6
timestamp 1731220596
transform 1 0 2192 0 -1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5177_6
timestamp 1731220596
transform 1 0 2128 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5176_6
timestamp 1731220596
transform 1 0 1968 0 1 2008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5175_6
timestamp 1731220596
transform 1 0 2016 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5174_6
timestamp 1731220596
transform 1 0 2160 0 -1 2148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5173_6
timestamp 1731220596
transform 1 0 2320 0 1 2156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5172_6
timestamp 1731220596
transform 1 0 2152 0 1 2156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5171_6
timestamp 1731220596
transform 1 0 1992 0 1 2156
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5170_6
timestamp 1731220596
transform 1 0 1968 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5169_6
timestamp 1731220596
transform 1 0 2136 0 -1 2292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5168_6
timestamp 1731220596
transform 1 0 2072 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5167_6
timestamp 1731220596
transform 1 0 1912 0 1 2296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5166_6
timestamp 1731220596
transform 1 0 1880 0 -1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5165_6
timestamp 1731220596
transform 1 0 2008 0 -1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5164_6
timestamp 1731220596
transform 1 0 2016 0 1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5163_6
timestamp 1731220596
transform 1 0 1880 0 1 2436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5162_6
timestamp 1731220596
transform 1 0 1880 0 -1 2576
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5161_6
timestamp 1731220596
transform 1 0 1984 0 -1 2576
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5160_6
timestamp 1731220596
transform 1 0 1984 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5159_6
timestamp 1731220596
transform 1 0 1880 0 1 2580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5158_6
timestamp 1731220596
transform 1 0 1880 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5157_6
timestamp 1731220596
transform 1 0 2040 0 -1 2724
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5156_6
timestamp 1731220596
transform 1 0 1880 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5155_6
timestamp 1731220596
transform 1 0 2048 0 1 2728
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5154_6
timestamp 1731220596
transform 1 0 2016 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5153_6
timestamp 1731220596
transform 1 0 1880 0 -1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5152_6
timestamp 1731220596
transform 1 0 1880 0 1 2864
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5151_6
timestamp 1731220596
transform 1 0 1720 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5150_6
timestamp 1731220596
transform 1 0 1632 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5149_6
timestamp 1731220596
transform 1 0 1720 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5148_6
timestamp 1731220596
transform 1 0 1688 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5147_6
timestamp 1731220596
transform 1 0 1552 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5146_6
timestamp 1731220596
transform 1 0 1448 0 1 3108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5145_6
timestamp 1731220596
transform 1 0 1624 0 1 3108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5144_6
timestamp 1731220596
transform 1 0 1568 0 -1 3252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5143_6
timestamp 1731220596
transform 1 0 1408 0 -1 3252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5142_6
timestamp 1731220596
transform 1 0 1336 0 1 3256
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5141_6
timestamp 1731220596
transform 1 0 1528 0 1 3256
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5140_6
timestamp 1731220596
transform 1 0 1520 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5139_6
timestamp 1731220596
transform 1 0 1360 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5138_6
timestamp 1731220596
transform 1 0 1200 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5137_6
timestamp 1731220596
transform 1 0 1168 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5136_6
timestamp 1731220596
transform 1 0 1312 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5135_6
timestamp 1731220596
transform 1 0 1464 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5134_6
timestamp 1731220596
transform 1 0 1568 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5133_6
timestamp 1731220596
transform 1 0 1464 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5132_6
timestamp 1731220596
transform 1 0 1360 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5131_6
timestamp 1731220596
transform 1 0 1264 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5130_6
timestamp 1731220596
transform 1 0 1168 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5129_6
timestamp 1731220596
transform 1 0 1072 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5128_6
timestamp 1731220596
transform 1 0 968 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5127_6
timestamp 1731220596
transform 1 0 856 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5126_6
timestamp 1731220596
transform 1 0 736 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5125_6
timestamp 1731220596
transform 1 0 880 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5124_6
timestamp 1731220596
transform 1 0 1024 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5123_6
timestamp 1731220596
transform 1 0 1040 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5122_6
timestamp 1731220596
transform 1 0 880 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5121_6
timestamp 1731220596
transform 1 0 968 0 1 3256
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5120_6
timestamp 1731220596
transform 1 0 1152 0 1 3256
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5119_6
timestamp 1731220596
transform 1 0 1088 0 -1 3252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5118_6
timestamp 1731220596
transform 1 0 928 0 -1 3252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5117_6
timestamp 1731220596
transform 1 0 1248 0 -1 3252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5116_6
timestamp 1731220596
transform 1 0 1120 0 1 3108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5115_6
timestamp 1731220596
transform 1 0 1280 0 1 3108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5114_6
timestamp 1731220596
transform 1 0 1416 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5113_6
timestamp 1731220596
transform 1 0 1280 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5112_6
timestamp 1731220596
transform 1 0 1152 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5111_6
timestamp 1731220596
transform 1 0 1224 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5110_6
timestamp 1731220596
transform 1 0 1352 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5109_6
timestamp 1731220596
transform 1 0 1480 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5108_6
timestamp 1731220596
transform 1 0 1608 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5107_6
timestamp 1731220596
transform 1 0 1520 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5106_6
timestamp 1731220596
transform 1 0 1408 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5105_6
timestamp 1731220596
transform 1 0 1296 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5104_6
timestamp 1731220596
transform 1 0 1176 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5103_6
timestamp 1731220596
transform 1 0 1048 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5102_6
timestamp 1731220596
transform 1 0 1536 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5101_6
timestamp 1731220596
transform 1 0 1400 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5100_6
timestamp 1731220596
transform 1 0 1264 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_599_6
timestamp 1731220596
transform 1 0 1128 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_598_6
timestamp 1731220596
transform 1 0 992 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_597_6
timestamp 1731220596
transform 1 0 1336 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_596_6
timestamp 1731220596
transform 1 0 1200 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_595_6
timestamp 1731220596
transform 1 0 1072 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_594_6
timestamp 1731220596
transform 1 0 944 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_593_6
timestamp 1731220596
transform 1 0 816 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_592_6
timestamp 1731220596
transform 1 0 1032 0 1 2668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_591_6
timestamp 1731220596
transform 1 0 888 0 1 2668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_590_6
timestamp 1731220596
transform 1 0 744 0 1 2668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_589_6
timestamp 1731220596
transform 1 0 576 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_588_6
timestamp 1731220596
transform 1 0 536 0 1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_587_6
timestamp 1731220596
transform 1 0 664 0 1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_586_6
timestamp 1731220596
transform 1 0 584 0 -1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_585_6
timestamp 1731220596
transform 1 0 576 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_584_6
timestamp 1731220596
transform 1 0 712 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_583_6
timestamp 1731220596
transform 1 0 808 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_582_6
timestamp 1731220596
transform 1 0 680 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_581_6
timestamp 1731220596
transform 1 0 552 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_580_6
timestamp 1731220596
transform 1 0 432 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_579_6
timestamp 1731220596
transform 1 0 328 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_578_6
timestamp 1731220596
transform 1 0 240 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_577_6
timestamp 1731220596
transform 1 0 152 0 -1 2376
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_576_6
timestamp 1731220596
transform 1 0 176 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_575_6
timestamp 1731220596
transform 1 0 304 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_574_6
timestamp 1731220596
transform 1 0 440 0 1 2388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_573_6
timestamp 1731220596
transform 1 0 432 0 -1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_572_6
timestamp 1731220596
transform 1 0 272 0 -1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_571_6
timestamp 1731220596
transform 1 0 128 0 -1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_570_6
timestamp 1731220596
transform 1 0 128 0 1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_569_6
timestamp 1731220596
transform 1 0 256 0 1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_568_6
timestamp 1731220596
transform 1 0 400 0 1 2524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_567_6
timestamp 1731220596
transform 1 0 464 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_566_6
timestamp 1731220596
transform 1 0 344 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_565_6
timestamp 1731220596
transform 1 0 224 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_564_6
timestamp 1731220596
transform 1 0 128 0 -1 2664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_563_6
timestamp 1731220596
transform 1 0 128 0 1 2668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_562_6
timestamp 1731220596
transform 1 0 216 0 1 2668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_561_6
timestamp 1731220596
transform 1 0 600 0 1 2668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_560_6
timestamp 1731220596
transform 1 0 464 0 1 2668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_559_6
timestamp 1731220596
transform 1 0 336 0 1 2668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_558_6
timestamp 1731220596
transform 1 0 288 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_557_6
timestamp 1731220596
transform 1 0 160 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_556_6
timestamp 1731220596
transform 1 0 688 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_555_6
timestamp 1731220596
transform 1 0 552 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_554_6
timestamp 1731220596
transform 1 0 416 0 -1 2812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_553_6
timestamp 1731220596
transform 1 0 312 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_552_6
timestamp 1731220596
transform 1 0 440 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_551_6
timestamp 1731220596
transform 1 0 576 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_550_6
timestamp 1731220596
transform 1 0 712 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_549_6
timestamp 1731220596
transform 1 0 856 0 1 2820
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_548_6
timestamp 1731220596
transform 1 0 912 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_547_6
timestamp 1731220596
transform 1 0 776 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_546_6
timestamp 1731220596
transform 1 0 632 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_545_6
timestamp 1731220596
transform 1 0 488 0 -1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_544_6
timestamp 1731220596
transform 1 0 560 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_543_6
timestamp 1731220596
transform 1 0 688 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_542_6
timestamp 1731220596
transform 1 0 816 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_541_6
timestamp 1731220596
transform 1 0 952 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_540_6
timestamp 1731220596
transform 1 0 1088 0 1 2960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_539_6
timestamp 1731220596
transform 1 0 1024 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_538_6
timestamp 1731220596
transform 1 0 896 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_537_6
timestamp 1731220596
transform 1 0 776 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_536_6
timestamp 1731220596
transform 1 0 656 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_535_6
timestamp 1731220596
transform 1 0 544 0 -1 3100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_534_6
timestamp 1731220596
transform 1 0 960 0 1 3108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_533_6
timestamp 1731220596
transform 1 0 808 0 1 3108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_532_6
timestamp 1731220596
transform 1 0 672 0 1 3108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_531_6
timestamp 1731220596
transform 1 0 544 0 1 3108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_530_6
timestamp 1731220596
transform 1 0 432 0 1 3108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_529_6
timestamp 1731220596
transform 1 0 776 0 -1 3252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_528_6
timestamp 1731220596
transform 1 0 632 0 -1 3252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_527_6
timestamp 1731220596
transform 1 0 496 0 -1 3252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_526_6
timestamp 1731220596
transform 1 0 360 0 -1 3252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_525_6
timestamp 1731220596
transform 1 0 792 0 1 3256
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_524_6
timestamp 1731220596
transform 1 0 624 0 1 3256
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_523_6
timestamp 1731220596
transform 1 0 464 0 1 3256
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_522_6
timestamp 1731220596
transform 1 0 320 0 1 3256
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_521_6
timestamp 1731220596
transform 1 0 192 0 1 3256
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_520_6
timestamp 1731220596
transform 1 0 720 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_519_6
timestamp 1731220596
transform 1 0 560 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_518_6
timestamp 1731220596
transform 1 0 400 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_517_6
timestamp 1731220596
transform 1 0 256 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_516_6
timestamp 1731220596
transform 1 0 128 0 -1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_515_6
timestamp 1731220596
transform 1 0 160 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_514_6
timestamp 1731220596
transform 1 0 288 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_513_6
timestamp 1731220596
transform 1 0 432 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_512_6
timestamp 1731220596
transform 1 0 576 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_511_6
timestamp 1731220596
transform 1 0 728 0 1 3396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_510_6
timestamp 1731220596
transform 1 0 616 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_59_6
timestamp 1731220596
transform 1 0 496 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_58_6
timestamp 1731220596
transform 1 0 368 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_57_6
timestamp 1731220596
transform 1 0 240 0 -1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_56_6
timestamp 1731220596
transform 1 0 480 0 1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_55_6
timestamp 1731220596
transform 1 0 392 0 1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_54_6
timestamp 1731220596
transform 1 0 304 0 1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_53_6
timestamp 1731220596
transform 1 0 216 0 1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_52_6
timestamp 1731220596
transform 1 0 128 0 1 3532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_51_6
timestamp 1731220596
transform 1 0 216 0 -1 3668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_50_6
timestamp 1731220596
transform 1 0 128 0 -1 3668
box 8 4 80 64
<< end >>
