magic
tech sky130l
timestamp 1731220305
<< checkpaint >>
rect 12 89 108 104
rect -18 88 108 89
rect -18 85 110 88
rect -18 83 111 85
rect -19 81 111 83
rect -24 73 111 81
rect -24 5 124 73
rect -24 4 119 5
rect -24 -2 111 4
rect -19 -4 106 -2
rect -12 -9 101 -4
rect 17 -11 101 -9
rect 21 -13 97 -11
rect 24 -21 96 -13
rect 25 -26 96 -21
rect 28 -27 96 -26
<< ndiffusion >>
rect 8 34 13 36
rect 8 31 9 34
rect 12 31 13 34
rect 8 30 13 31
rect 41 30 44 36
rect 46 35 53 36
rect 46 32 49 35
rect 52 32 53 35
rect 46 30 53 32
rect 49 21 53 30
rect 55 21 58 36
rect 60 21 63 36
rect 65 34 70 36
rect 65 31 66 34
rect 69 31 70 34
rect 65 30 70 31
rect 74 35 79 36
rect 74 32 75 35
rect 78 32 79 35
rect 74 30 79 32
rect 65 21 69 30
<< ndc >>
rect 9 31 12 34
rect 49 32 52 35
rect 66 31 69 34
rect 75 32 78 35
<< ntransistor >>
rect 13 30 41 36
rect 44 30 46 36
rect 53 21 55 36
rect 58 21 60 36
rect 63 21 65 36
rect 70 30 74 36
<< pdiffusion >>
rect 49 49 53 61
rect 8 48 13 49
rect 8 45 9 48
rect 12 45 13 48
rect 8 43 13 45
rect 27 43 44 49
rect 46 47 53 49
rect 46 44 49 47
rect 52 44 53 47
rect 46 43 53 44
rect 55 43 58 61
rect 60 43 63 61
rect 65 53 69 61
rect 65 48 70 53
rect 65 45 66 48
rect 69 45 70 48
rect 65 43 70 45
rect 74 47 79 53
rect 74 44 75 47
rect 78 44 79 47
rect 74 43 79 44
<< pdc >>
rect 9 45 12 48
rect 49 44 52 47
rect 66 45 69 48
rect 75 44 78 47
<< ptransistor >>
rect 13 43 27 49
rect 44 43 46 49
rect 53 43 55 61
rect 58 43 60 61
rect 63 43 65 61
rect 70 43 74 53
<< polysilicon >>
rect 50 68 55 69
rect 50 65 51 68
rect 54 65 55 68
rect 50 64 55 65
rect 53 61 55 64
rect 63 68 68 69
rect 63 65 64 68
rect 67 65 68 68
rect 63 64 68 65
rect 58 61 60 63
rect 63 61 65 64
rect 14 56 19 57
rect 14 53 15 56
rect 18 53 19 56
rect 14 51 19 53
rect 41 56 46 57
rect 41 53 42 56
rect 45 53 46 56
rect 41 52 46 53
rect 13 49 27 51
rect 44 49 46 52
rect 70 53 74 55
rect 13 41 27 43
rect 13 36 41 38
rect 44 36 46 43
rect 53 36 55 43
rect 58 36 60 43
rect 63 36 65 43
rect 70 41 74 43
rect 70 40 87 41
rect 70 39 83 40
rect 70 36 74 39
rect 82 37 83 39
rect 86 37 87 40
rect 82 36 87 37
rect 13 28 41 30
rect 44 28 46 30
rect 20 27 25 28
rect 20 24 21 27
rect 24 24 25 27
rect 20 23 25 24
rect 70 28 74 30
rect 53 19 55 21
rect 58 16 60 21
rect 63 19 65 21
rect 56 15 61 16
rect 56 12 57 15
rect 60 12 61 15
rect 56 11 61 12
<< pc >>
rect 51 65 54 68
rect 64 65 67 68
rect 15 53 18 56
rect 42 53 45 56
rect 83 37 86 40
rect 21 24 24 27
rect 57 12 60 15
<< m1 >>
rect 44 68 48 72
rect 72 68 76 72
rect 44 66 51 68
rect 45 65 51 66
rect 54 65 55 68
rect 63 65 64 68
rect 67 65 75 68
rect 15 56 18 57
rect 41 53 42 56
rect 45 53 78 56
rect 9 48 12 49
rect 9 44 12 45
rect 9 34 12 35
rect 9 30 12 31
rect 15 34 18 53
rect 15 30 18 31
rect 21 48 24 49
rect 66 48 69 49
rect 21 27 24 45
rect 49 47 52 48
rect 66 44 69 45
rect 75 47 78 53
rect 49 41 52 44
rect 49 35 52 38
rect 75 35 78 44
rect 88 40 92 41
rect 82 37 83 40
rect 86 37 92 40
rect 49 31 52 32
rect 66 34 69 35
rect 75 31 78 32
rect 66 30 69 31
rect 21 23 24 24
rect 57 15 60 16
rect 57 9 60 12
rect 57 6 64 9
rect 60 5 64 6
<< m2c >>
rect 9 45 12 48
rect 9 31 12 34
rect 15 31 18 34
rect 21 45 24 48
rect 66 45 69 48
rect 49 38 52 41
rect 83 37 86 40
rect 66 31 69 34
<< m2 >>
rect 8 48 70 49
rect 8 45 9 48
rect 12 45 21 48
rect 24 45 66 48
rect 69 45 70 48
rect 8 44 70 45
rect 48 41 53 42
rect 48 38 49 41
rect 52 40 53 41
rect 82 40 87 41
rect 52 38 83 40
rect 48 37 53 38
rect 82 37 83 38
rect 86 37 87 40
rect 82 36 87 37
rect 8 34 70 35
rect 8 31 9 34
rect 12 31 15 34
rect 18 31 66 34
rect 69 31 70 34
rect 8 30 70 31
<< labels >>
rlabel space 0 0 96 76 6 prboundary
rlabel pdiffusion 79 45 79 45 3 #10
rlabel ndiffusion 79 33 79 33 3 #10
rlabel polysilicon 71 37 71 37 3 out
rlabel polysilicon 71 40 71 40 3 out
rlabel polysilicon 71 41 71 41 3 out
rlabel polysilicon 71 42 71 42 3 out
rlabel pdiffusion 75 44 75 44 3 #10
rlabel pdiffusion 75 45 75 45 3 #10
rlabel pdiffusion 75 48 75 48 3 #10
rlabel polysilicon 71 54 71 54 3 out
rlabel polysilicon 64 62 64 62 3 in(0)
rlabel polysilicon 64 65 64 65 3 in(0)
rlabel polysilicon 64 69 64 69 3 in(0)
rlabel polysilicon 71 29 71 29 3 out
rlabel ndiffusion 75 31 75 31 3 #10
rlabel ndiffusion 75 33 75 33 3 #10
rlabel ndiffusion 75 36 75 36 3 #10
rlabel polysilicon 64 37 64 37 3 in(0)
rlabel ptransistor 71 44 71 44 3 out
rlabel ntransistor 71 31 71 31 3 out
rlabel pdiffusion 66 44 66 44 3 Vdd
rlabel pdiffusion 66 46 66 46 3 Vdd
rlabel pdiffusion 66 49 66 49 3 Vdd
rlabel pdiffusion 66 54 66 54 3 Vdd
rlabel polysilicon 59 62 59 62 3 in(1)
rlabel ndiffusion 66 22 66 22 3 GND
rlabel ndiffusion 66 31 66 31 3 GND
rlabel ndiffusion 66 32 66 32 3 GND
rlabel ndiffusion 66 35 66 35 3 GND
rlabel polysilicon 59 37 59 37 3 in(1)
rlabel ptransistor 64 44 64 44 3 in(0)
rlabel polysilicon 64 20 64 20 3 in(0)
rlabel ntransistor 64 22 64 22 3 in(0)
rlabel polysilicon 54 62 54 62 3 in(2)
rlabel polysilicon 61 13 61 13 3 in(1)
rlabel polysilicon 54 37 54 37 3 in(2)
rlabel ptransistor 59 44 59 44 3 in(1)
rlabel polysilicon 51 65 51 65 3 in(2)
rlabel polysilicon 51 66 51 66 3 in(2)
rlabel polysilicon 51 69 51 69 3 in(2)
rlabel polysilicon 59 17 59 17 3 in(1)
rlabel ntransistor 59 22 59 22 3 in(1)
rlabel ndiffusion 53 33 53 33 3 out
rlabel pdiffusion 53 45 53 45 3 out
rlabel pdiffusion 50 50 50 50 3 out
rlabel polysilicon 57 12 57 12 3 in(1)
rlabel polysilicon 57 13 57 13 3 in(1)
rlabel polysilicon 57 16 57 16 3 in(1)
rlabel ptransistor 54 44 54 44 3 in(2)
rlabel polysilicon 54 20 54 20 3 in(2)
rlabel ntransistor 54 22 54 22 3 in(2)
rlabel polysilicon 25 25 25 25 3 Vdd
rlabel ndiffusion 47 31 47 31 3 out
rlabel ndiffusion 47 33 47 33 3 out
rlabel ndiffusion 47 36 47 36 3 out
rlabel pdiffusion 47 44 47 44 3 out
rlabel pdiffusion 47 45 47 45 3 out
rlabel pdiffusion 47 48 47 48 3 out
rlabel polysilicon 45 50 45 50 3 #10
rlabel polysilicon 19 54 19 54 3 GND
rlabel ndiffusion 50 22 50 22 3 out
rlabel polysilicon 45 29 45 29 3 #10
rlabel ntransistor 45 31 45 31 3 #10
rlabel polysilicon 45 37 45 37 3 #10
rlabel ptransistor 45 44 45 44 3 #10
rlabel polysilicon 42 53 42 53 3 #10
rlabel polysilicon 42 57 42 57 3 #10
rlabel polysilicon 21 24 21 24 3 Vdd
rlabel polysilicon 21 25 21 25 3 Vdd
rlabel polysilicon 21 28 21 28 3 Vdd
rlabel polysilicon 15 52 15 52 3 GND
rlabel polysilicon 15 54 15 54 3 GND
rlabel polysilicon 15 57 15 57 3 GND
rlabel polysilicon 14 29 14 29 3 Vdd
rlabel ntransistor 14 31 14 31 3 Vdd
rlabel polysilicon 14 37 14 37 3 Vdd
rlabel polysilicon 14 42 14 42 3 GND
rlabel ptransistor 14 44 14 44 3 GND
rlabel polysilicon 14 50 14 50 3 GND
rlabel pdiffusion 9 44 9 44 3 Vdd
rlabel m1 73 69 73 69 3 in(0)
port 1 e
rlabel m1 89 41 89 41 3 out
port 2 e
rlabel m1 68 66 68 66 3 in(0)
port 1 e
rlabel pc 65 66 65 66 3 in(0)
port 1 e
rlabel m1 64 66 64 66 3 in(0)
port 1 e
rlabel m1 55 66 55 66 3 in(2)
port 3 e
rlabel ndc 76 33 76 33 3 #10
rlabel m1 76 36 76 36 3 #10
rlabel pdc 76 45 76 45 3 #10
rlabel m1 76 48 76 48 3 #10
rlabel pc 52 66 52 66 3 in(2)
port 3 e
rlabel m1 76 32 76 32 3 #10
rlabel m1 46 66 46 66 3 in(2)
port 3 e
rlabel m1 46 54 46 54 3 #10
rlabel m1 45 67 45 67 3 in(2)
port 3 e
rlabel m1 45 69 45 69 3 in(2)
port 3 e
rlabel m1 67 35 67 35 3 GND
rlabel m1 67 45 67 45 3 Vdd
rlabel m1 67 49 67 49 3 Vdd
rlabel pc 43 54 43 54 3 #10
rlabel m1 22 49 22 49 3 Vdd
rlabel m1 42 54 42 54 3 #10
rlabel m1 61 6 61 6 3 in(1)
port 4 e
rlabel m1 67 31 67 31 3 GND
rlabel m1 50 32 50 32 3 out
port 2 e
rlabel ndc 50 33 50 33 3 out
port 2 e
rlabel m1 50 36 50 36 3 out
port 2 e
rlabel m1 50 42 50 42 3 out
port 2 e
rlabel pdc 50 45 50 45 3 out
port 2 e
rlabel m1 50 48 50 48 3 out
port 2 e
rlabel m1 58 7 58 7 3 in(1)
port 4 e
rlabel m1 58 10 58 10 3 in(1)
port 4 e
rlabel pc 58 13 58 13 3 in(1)
port 4 e
rlabel m1 58 16 58 16 3 in(1)
port 4 e
rlabel m1 16 31 16 31 3 GND
rlabel m1 16 35 16 35 3 GND
rlabel pc 16 54 16 54 3 GND
rlabel m1 16 57 16 57 3 GND
rlabel m1 22 24 22 24 3 Vdd
rlabel pc 22 25 22 25 3 Vdd
rlabel m1 22 28 22 28 3 Vdd
rlabel m1 10 31 10 31 3 GND
rlabel m1 10 35 10 35 3 GND
rlabel m1 10 45 10 45 3 Vdd
rlabel m1 10 49 10 49 3 Vdd
rlabel m2 83 41 83 41 3 out
port 2 e
rlabel m2 53 39 53 39 3 out
port 2 e
rlabel m2 53 41 53 41 3 out
port 2 e
rlabel m2 70 32 70 32 3 GND
rlabel m2c 50 39 50 39 3 out
port 2 e
rlabel m2 70 46 70 46 3 Vdd
rlabel m2c 67 32 67 32 3 GND
rlabel m2 49 38 49 38 3 out
port 2 e
rlabel m2 49 39 49 39 3 out
port 2 e
rlabel m2 49 42 49 42 3 out
port 2 e
rlabel m2c 67 46 67 46 3 Vdd
rlabel m2 19 32 19 32 3 GND
rlabel m2 87 38 87 38 3 out
port 2 e
rlabel m2 25 46 25 46 3 Vdd
rlabel m2c 16 32 16 32 3 GND
rlabel m2c 84 38 84 38 3 out
port 2 e
rlabel m2c 22 46 22 46 3 Vdd
rlabel m2 13 32 13 32 3 GND
rlabel m2 83 37 83 37 3 out
port 2 e
rlabel m2 83 38 83 38 3 out
port 2 e
rlabel m2 13 46 13 46 3 Vdd
rlabel m2c 10 32 10 32 3 GND
rlabel m2c 10 46 10 46 3 Vdd
rlabel m2 9 31 9 31 3 GND
rlabel m2 9 32 9 32 3 GND
rlabel m2 9 35 9 35 3 GND
rlabel m2 9 45 9 45 3 Vdd
rlabel m2 9 46 9 46 3 Vdd
rlabel m2 9 49 9 49 3 Vdd
<< end >>
