magic
tech sky130l
timestamp 1730768468
<< m1 >>
rect 8 97 12 98
rect 8 94 9 97
rect 8 72 12 94
rect 30 97 33 98
rect 30 93 33 94
rect 44 97 47 98
rect 44 93 47 94
rect 69 97 72 98
rect 69 93 72 94
rect 22 89 25 90
rect 22 85 25 86
rect 36 89 39 90
rect 36 85 39 86
rect 50 89 53 90
rect 64 89 68 90
rect 50 85 53 86
rect 15 81 18 82
rect 15 77 18 78
rect 58 81 61 87
rect 58 77 61 78
rect 67 86 68 89
rect 64 72 68 86
rect 72 81 76 82
rect 75 78 76 81
rect 72 72 76 78
rect 81 81 84 98
rect 89 89 92 98
rect 97 97 100 98
rect 97 93 100 94
rect 81 77 84 78
rect 8 44 12 52
rect 15 46 36 49
rect 54 47 75 50
rect 8 41 9 44
rect 47 44 50 45
rect 97 44 100 45
rect 8 40 12 41
rect 9 19 12 28
rect 17 5 20 27
rect 24 5 29 43
rect 62 41 63 44
rect 66 41 67 44
rect 47 40 50 41
rect 32 30 35 31
rect 47 30 50 31
rect 32 16 35 27
rect 39 19 42 28
rect 62 27 63 30
rect 66 27 67 30
rect 47 26 50 27
rect 54 21 75 24
rect 80 19 83 44
rect 97 40 100 41
rect 97 30 100 31
rect 104 27 108 52
rect 112 37 118 52
rect 122 44 125 45
rect 122 40 125 41
rect 112 34 125 37
rect 115 30 118 31
rect 122 27 125 34
rect 97 26 100 27
rect 115 26 118 27
rect 116 20 121 23
rect 32 12 36 16
rect 75 6 80 9
rect 101 6 106 9
<< m2c >>
rect 9 94 12 97
rect 30 94 33 97
rect 44 94 47 97
rect 69 94 72 97
rect 22 86 25 89
rect 36 86 39 89
rect 50 86 53 89
rect 15 78 18 81
rect 58 78 61 81
rect 64 86 67 89
rect 72 78 75 81
rect 97 94 100 97
rect 89 86 92 89
rect 81 78 84 81
rect 9 41 12 44
rect 47 41 50 44
rect 63 41 66 44
rect 32 27 35 30
rect 47 27 50 30
rect 63 27 66 30
rect 97 41 100 44
rect 97 27 100 30
rect 122 41 125 44
rect 115 27 118 30
<< m2 >>
rect 8 97 101 98
rect 8 94 9 97
rect 12 94 30 97
rect 33 94 44 97
rect 47 94 69 97
rect 72 94 97 97
rect 100 94 101 97
rect 8 93 101 94
rect 21 89 93 90
rect 21 86 22 89
rect 25 86 36 89
rect 39 86 50 89
rect 53 86 64 89
rect 67 86 89 89
rect 92 86 93 89
rect 21 85 93 86
rect 14 81 85 82
rect 14 78 15 81
rect 18 78 58 81
rect 61 78 72 81
rect 75 78 81 81
rect 84 78 85 81
rect 14 77 85 78
rect 8 44 126 45
rect 8 41 9 44
rect 12 41 47 44
rect 50 41 63 44
rect 66 41 97 44
rect 100 41 122 44
rect 125 41 126 44
rect 8 40 126 41
rect 31 30 119 31
rect 31 27 32 30
rect 35 27 47 30
rect 50 27 63 30
rect 66 27 97 30
rect 100 27 115 30
rect 118 27 119 30
rect 31 26 119 27
rect 8 19 43 24
rect 79 19 121 24
rect 16 5 106 10
<< labels >>
rlabel m2 s 100 94 101 97 6 A
port 1 nsew signal input
rlabel m2 s 97 94 100 97 6 A
port 1 nsew signal input
rlabel m2 s 72 94 97 97 6 A
port 1 nsew signal input
rlabel m2 s 69 94 72 97 6 A
port 1 nsew signal input
rlabel m2 s 47 94 69 97 6 A
port 1 nsew signal input
rlabel m2 s 44 94 47 97 6 A
port 1 nsew signal input
rlabel m2 s 33 94 44 97 6 A
port 1 nsew signal input
rlabel m2 s 30 94 33 97 6 A
port 1 nsew signal input
rlabel m2 s 12 94 30 97 6 A
port 1 nsew signal input
rlabel m2 s 9 94 12 97 6 A
port 1 nsew signal input
rlabel m2 s 8 93 101 94 6 A
port 1 nsew signal input
rlabel m2 s 8 94 9 97 6 A
port 1 nsew signal input
rlabel m2 s 8 97 101 98 6 A
port 1 nsew signal input
rlabel m2c s 97 94 100 97 6 A
port 1 nsew signal input
rlabel m2c s 69 94 72 97 6 A
port 1 nsew signal input
rlabel m2c s 44 94 47 97 6 A
port 1 nsew signal input
rlabel m2c s 30 94 33 97 6 A
port 1 nsew signal input
rlabel m2c s 9 94 12 97 6 A
port 1 nsew signal input
rlabel m1 s 97 93 100 94 6 A
port 1 nsew signal input
rlabel m1 s 97 94 100 97 6 A
port 1 nsew signal input
rlabel m1 s 97 97 100 98 6 A
port 1 nsew signal input
rlabel m1 s 69 93 72 94 6 A
port 1 nsew signal input
rlabel m1 s 69 94 72 97 6 A
port 1 nsew signal input
rlabel m1 s 69 97 72 98 6 A
port 1 nsew signal input
rlabel m1 s 44 93 47 94 6 A
port 1 nsew signal input
rlabel m1 s 44 94 47 97 6 A
port 1 nsew signal input
rlabel m1 s 44 97 47 98 6 A
port 1 nsew signal input
rlabel m1 s 30 93 33 94 6 A
port 1 nsew signal input
rlabel m1 s 30 94 33 97 6 A
port 1 nsew signal input
rlabel m1 s 30 97 33 98 6 A
port 1 nsew signal input
rlabel m1 s 9 94 12 97 6 A
port 1 nsew signal input
rlabel m1 s 8 72 12 94 6 A
port 1 nsew signal input
rlabel m1 s 8 94 9 97 6 A
port 1 nsew signal input
rlabel m1 s 8 97 12 98 6 A
port 1 nsew signal input
rlabel m2 s 92 86 93 89 6 B
port 2 nsew signal input
rlabel m2 s 89 86 92 89 6 B
port 2 nsew signal input
rlabel m2 s 67 86 89 89 6 B
port 2 nsew signal input
rlabel m2 s 64 86 67 89 6 B
port 2 nsew signal input
rlabel m2 s 53 86 64 89 6 B
port 2 nsew signal input
rlabel m2 s 50 86 53 89 6 B
port 2 nsew signal input
rlabel m2 s 39 86 50 89 6 B
port 2 nsew signal input
rlabel m2 s 36 86 39 89 6 B
port 2 nsew signal input
rlabel m2 s 25 86 36 89 6 B
port 2 nsew signal input
rlabel m2 s 22 86 25 89 6 B
port 2 nsew signal input
rlabel m2 s 21 85 93 86 6 B
port 2 nsew signal input
rlabel m2 s 21 86 22 89 6 B
port 2 nsew signal input
rlabel m2 s 21 89 93 90 6 B
port 2 nsew signal input
rlabel m2c s 89 86 92 89 6 B
port 2 nsew signal input
rlabel m2c s 64 86 67 89 6 B
port 2 nsew signal input
rlabel m2c s 50 86 53 89 6 B
port 2 nsew signal input
rlabel m2c s 36 86 39 89 6 B
port 2 nsew signal input
rlabel m2c s 22 86 25 89 6 B
port 2 nsew signal input
rlabel m1 s 89 86 92 89 6 B
port 2 nsew signal input
rlabel m1 s 89 89 92 94 6 B
port 2 nsew signal input
rlabel m1 s 89 94 92 97 6 B
port 2 nsew signal input
rlabel m1 s 89 97 92 98 6 B
port 2 nsew signal input
rlabel m1 s 67 86 68 89 6 B
port 2 nsew signal input
rlabel m1 s 64 72 68 86 6 B
port 2 nsew signal input
rlabel m1 s 64 86 67 89 6 B
port 2 nsew signal input
rlabel m1 s 64 89 68 90 6 B
port 2 nsew signal input
rlabel m1 s 50 85 53 86 6 B
port 2 nsew signal input
rlabel m1 s 50 86 53 89 6 B
port 2 nsew signal input
rlabel m1 s 50 89 53 90 6 B
port 2 nsew signal input
rlabel m1 s 36 85 39 86 6 B
port 2 nsew signal input
rlabel m1 s 36 86 39 89 6 B
port 2 nsew signal input
rlabel m1 s 36 89 39 90 6 B
port 2 nsew signal input
rlabel m1 s 22 85 25 86 6 B
port 2 nsew signal input
rlabel m1 s 22 86 25 89 6 B
port 2 nsew signal input
rlabel m1 s 22 89 25 90 6 B
port 2 nsew signal input
rlabel m2 s 84 78 85 81 6 C
port 3 nsew signal input
rlabel m2 s 81 78 84 81 6 C
port 3 nsew signal input
rlabel m2 s 75 78 81 81 6 C
port 3 nsew signal input
rlabel m2 s 72 78 75 81 6 C
port 3 nsew signal input
rlabel m2 s 61 78 72 81 6 C
port 3 nsew signal input
rlabel m2 s 58 78 61 81 6 C
port 3 nsew signal input
rlabel m2 s 18 78 58 81 6 C
port 3 nsew signal input
rlabel m2 s 15 78 18 81 6 C
port 3 nsew signal input
rlabel m2 s 14 77 85 78 6 C
port 3 nsew signal input
rlabel m2 s 14 78 15 81 6 C
port 3 nsew signal input
rlabel m2 s 14 81 85 82 6 C
port 3 nsew signal input
rlabel m2c s 81 78 84 81 6 C
port 3 nsew signal input
rlabel m2c s 72 78 75 81 6 C
port 3 nsew signal input
rlabel m2c s 58 78 61 81 6 C
port 3 nsew signal input
rlabel m2c s 15 78 18 81 6 C
port 3 nsew signal input
rlabel m1 s 81 77 84 78 6 C
port 3 nsew signal input
rlabel m1 s 81 78 84 81 6 C
port 3 nsew signal input
rlabel m1 s 81 81 84 94 6 C
port 3 nsew signal input
rlabel m1 s 81 94 84 97 6 C
port 3 nsew signal input
rlabel m1 s 81 97 84 98 6 C
port 3 nsew signal input
rlabel m1 s 75 78 76 81 6 C
port 3 nsew signal input
rlabel m1 s 72 72 76 78 6 C
port 3 nsew signal input
rlabel m1 s 72 78 75 81 6 C
port 3 nsew signal input
rlabel m1 s 72 81 76 82 6 C
port 3 nsew signal input
rlabel m1 s 58 77 61 78 6 C
port 3 nsew signal input
rlabel m1 s 58 78 61 81 6 C
port 3 nsew signal input
rlabel m1 s 58 81 61 83 6 C
port 3 nsew signal input
rlabel m1 s 58 83 61 86 6 C
port 3 nsew signal input
rlabel m1 s 58 86 61 87 6 C
port 3 nsew signal input
rlabel m1 s 15 77 18 78 6 C
port 3 nsew signal input
rlabel m1 s 15 78 18 81 6 C
port 3 nsew signal input
rlabel m1 s 15 81 18 82 6 C
port 3 nsew signal input
rlabel m1 s 107 28 108 31 6 YC
port 4 nsew signal output
rlabel m1 s 107 43 108 46 6 YC
port 4 nsew signal output
rlabel m1 s 104 27 108 28 6 YC
port 4 nsew signal output
rlabel m1 s 104 28 107 31 6 YC
port 4 nsew signal output
rlabel m1 s 104 31 108 43 6 YC
port 4 nsew signal output
rlabel m1 s 104 43 107 46 6 YC
port 4 nsew signal output
rlabel m1 s 104 46 108 52 6 YC
port 4 nsew signal output
rlabel m1 s 122 27 125 28 6 YS
port 5 nsew signal output
rlabel m1 s 122 28 125 31 6 YS
port 5 nsew signal output
rlabel m1 s 122 31 125 34 6 YS
port 5 nsew signal output
rlabel m1 s 115 43 118 46 6 YS
port 5 nsew signal output
rlabel m1 s 112 34 125 37 6 YS
port 5 nsew signal output
rlabel m1 s 112 37 118 43 6 YS
port 5 nsew signal output
rlabel m1 s 112 43 115 46 6 YS
port 5 nsew signal output
rlabel m1 s 112 46 118 52 6 YS
port 5 nsew signal output
rlabel m2 s 125 41 126 44 6 Vdd
port 6 nsew power input
rlabel m2 s 122 41 125 44 6 Vdd
port 6 nsew power input
rlabel m2 s 100 41 122 44 6 Vdd
port 6 nsew power input
rlabel m2 s 97 41 100 44 6 Vdd
port 6 nsew power input
rlabel m2 s 66 41 97 44 6 Vdd
port 6 nsew power input
rlabel m2 s 63 41 66 44 6 Vdd
port 6 nsew power input
rlabel m2 s 50 41 63 44 6 Vdd
port 6 nsew power input
rlabel m2 s 47 41 50 44 6 Vdd
port 6 nsew power input
rlabel m2 s 12 41 47 44 6 Vdd
port 6 nsew power input
rlabel m2 s 9 41 12 44 6 Vdd
port 6 nsew power input
rlabel m2 s 8 40 126 41 6 Vdd
port 6 nsew power input
rlabel m2 s 8 41 9 44 6 Vdd
port 6 nsew power input
rlabel m2 s 8 44 126 45 6 Vdd
port 6 nsew power input
rlabel m2c s 122 41 125 44 6 Vdd
port 6 nsew power input
rlabel m2c s 97 41 100 44 6 Vdd
port 6 nsew power input
rlabel m2c s 63 41 66 44 6 Vdd
port 6 nsew power input
rlabel m2c s 47 41 50 44 6 Vdd
port 6 nsew power input
rlabel m2c s 9 41 12 44 6 Vdd
port 6 nsew power input
rlabel m1 s 122 40 125 41 6 Vdd
port 6 nsew power input
rlabel m1 s 122 41 125 44 6 Vdd
port 6 nsew power input
rlabel m1 s 122 44 125 45 6 Vdd
port 6 nsew power input
rlabel m1 s 97 40 100 41 6 Vdd
port 6 nsew power input
rlabel m1 s 97 41 100 44 6 Vdd
port 6 nsew power input
rlabel m1 s 97 44 100 45 6 Vdd
port 6 nsew power input
rlabel m1 s 66 41 67 44 6 Vdd
port 6 nsew power input
rlabel m1 s 63 41 66 44 6 Vdd
port 6 nsew power input
rlabel m1 s 62 41 63 44 6 Vdd
port 6 nsew power input
rlabel m1 s 47 40 50 41 6 Vdd
port 6 nsew power input
rlabel m1 s 47 41 50 44 6 Vdd
port 6 nsew power input
rlabel m1 s 47 44 50 45 6 Vdd
port 6 nsew power input
rlabel m1 s 9 41 12 44 6 Vdd
port 6 nsew power input
rlabel m1 s 8 40 12 41 6 Vdd
port 6 nsew power input
rlabel m1 s 8 41 9 44 6 Vdd
port 6 nsew power input
rlabel m1 s 8 44 12 52 6 Vdd
port 6 nsew power input
rlabel m2 s 118 27 119 30 6 GND
port 7 nsew ground input
rlabel m2 s 115 27 118 30 6 GND
port 7 nsew ground input
rlabel m2 s 100 27 115 30 6 GND
port 7 nsew ground input
rlabel m2 s 97 27 100 30 6 GND
port 7 nsew ground input
rlabel m2 s 66 27 97 30 6 GND
port 7 nsew ground input
rlabel m2 s 63 27 66 30 6 GND
port 7 nsew ground input
rlabel m2 s 50 27 63 30 6 GND
port 7 nsew ground input
rlabel m2 s 47 27 50 30 6 GND
port 7 nsew ground input
rlabel m2 s 35 27 47 30 6 GND
port 7 nsew ground input
rlabel m2 s 32 27 35 30 6 GND
port 7 nsew ground input
rlabel m2 s 31 26 119 27 6 GND
port 7 nsew ground input
rlabel m2 s 31 27 32 30 6 GND
port 7 nsew ground input
rlabel m2 s 31 30 119 31 6 GND
port 7 nsew ground input
rlabel m2c s 115 27 118 30 6 GND
port 7 nsew ground input
rlabel m2c s 97 27 100 30 6 GND
port 7 nsew ground input
rlabel m2c s 63 27 66 30 6 GND
port 7 nsew ground input
rlabel m2c s 47 27 50 30 6 GND
port 7 nsew ground input
rlabel m2c s 32 27 35 30 6 GND
port 7 nsew ground input
rlabel m1 s 115 26 118 27 6 GND
port 7 nsew ground input
rlabel m1 s 115 27 118 30 6 GND
port 7 nsew ground input
rlabel m1 s 115 30 118 31 6 GND
port 7 nsew ground input
rlabel m1 s 97 26 100 27 6 GND
port 7 nsew ground input
rlabel m1 s 97 27 100 30 6 GND
port 7 nsew ground input
rlabel m1 s 97 30 100 31 6 GND
port 7 nsew ground input
rlabel m1 s 66 27 67 30 6 GND
port 7 nsew ground input
rlabel m1 s 63 27 66 30 6 GND
port 7 nsew ground input
rlabel m1 s 62 27 63 30 6 GND
port 7 nsew ground input
rlabel m1 s 47 26 50 27 6 GND
port 7 nsew ground input
rlabel m1 s 47 27 50 30 6 GND
port 7 nsew ground input
rlabel m1 s 47 30 50 31 6 GND
port 7 nsew ground input
rlabel m1 s 32 12 36 16 6 GND
port 7 nsew ground input
rlabel m1 s 32 16 35 27 6 GND
port 7 nsew ground input
rlabel m1 s 32 27 35 30 6 GND
port 7 nsew ground input
rlabel m1 s 32 30 35 31 6 GND
port 7 nsew ground input
<< properties >>
string LEFsite CoreSite
string LEFclass CORE
string FIXED_BBOX 0 0 136 100
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
