magic
tech sky130l
timestamp 1731220378
<< m1 >>
rect 616 1555 620 1579
rect 280 1527 284 1547
rect 344 1511 348 1535
rect 1064 1523 1068 1539
rect 440 1479 444 1523
rect 600 1451 604 1467
rect 1424 1451 1428 1467
rect 1264 1379 1268 1395
rect 1088 1335 1092 1363
rect 696 1263 700 1291
rect 1032 1207 1036 1247
rect 1064 1179 1068 1203
rect 1568 1179 1572 1203
rect 288 1151 292 1175
rect 1568 1107 1572 1131
rect 472 1011 476 1035
rect 1568 943 1572 967
rect 848 879 852 911
rect 872 867 876 903
rect 1400 895 1404 939
rect 368 851 372 867
rect 416 819 420 863
rect 448 795 452 831
rect 1128 803 1132 851
rect 1240 839 1244 863
rect 224 747 228 791
rect 328 775 332 791
rect 760 775 764 791
rect 280 555 284 571
rect 448 527 452 571
rect 864 555 868 579
rect 1568 571 1572 595
rect 792 499 796 523
rect 952 511 956 551
rect 1192 511 1196 555
rect 1472 499 1476 523
rect 1568 439 1572 523
rect 456 379 460 419
rect 744 379 748 419
rect 1568 351 1572 375
rect 1144 259 1148 275
rect 1328 259 1332 275
rect 1384 263 1388 287
rect 752 207 756 227
rect 1568 199 1572 227
rect 240 183 244 199
rect 968 123 972 151
<< m2c >>
rect 152 1635 156 1639
rect 184 1635 188 1639
rect 216 1635 220 1639
rect 152 1619 156 1623
rect 184 1619 188 1623
rect 152 1607 156 1611
rect 192 1607 196 1611
rect 256 1607 260 1611
rect 312 1607 316 1611
rect 368 1607 372 1611
rect 424 1607 428 1611
rect 472 1607 476 1611
rect 520 1607 524 1611
rect 568 1607 572 1611
rect 616 1607 620 1611
rect 664 1607 668 1611
rect 712 1607 716 1611
rect 760 1607 764 1611
rect 808 1607 812 1611
rect 856 1607 860 1611
rect 904 1607 908 1611
rect 952 1607 956 1611
rect 1008 1607 1012 1611
rect 1064 1607 1068 1611
rect 1112 1607 1116 1611
rect 1160 1607 1164 1611
rect 1208 1607 1212 1611
rect 1256 1607 1260 1611
rect 1304 1607 1308 1611
rect 1344 1607 1348 1611
rect 1384 1607 1388 1611
rect 1424 1607 1428 1611
rect 1464 1607 1468 1611
rect 1496 1607 1500 1611
rect 1528 1607 1532 1611
rect 1560 1607 1564 1611
rect 152 1591 156 1595
rect 192 1591 196 1595
rect 256 1591 260 1595
rect 312 1591 316 1595
rect 368 1591 372 1595
rect 424 1591 428 1595
rect 472 1591 476 1595
rect 520 1591 524 1595
rect 568 1591 572 1595
rect 616 1591 620 1595
rect 664 1591 668 1595
rect 712 1591 716 1595
rect 760 1591 764 1595
rect 808 1591 812 1595
rect 856 1591 860 1595
rect 904 1591 908 1595
rect 952 1591 956 1595
rect 1008 1591 1012 1595
rect 1064 1591 1068 1595
rect 1112 1591 1116 1595
rect 1160 1591 1164 1595
rect 1208 1591 1212 1595
rect 1256 1591 1260 1595
rect 1304 1591 1308 1595
rect 1344 1591 1348 1595
rect 1384 1591 1388 1595
rect 1424 1591 1428 1595
rect 1464 1591 1468 1595
rect 1496 1591 1500 1595
rect 1528 1591 1532 1595
rect 1560 1591 1564 1595
rect 616 1579 620 1583
rect 192 1563 196 1567
rect 232 1563 236 1567
rect 272 1563 276 1567
rect 312 1563 316 1567
rect 360 1563 364 1567
rect 408 1563 412 1567
rect 456 1563 460 1567
rect 504 1563 508 1567
rect 552 1563 556 1567
rect 600 1563 604 1567
rect 656 1563 660 1567
rect 720 1563 724 1567
rect 792 1563 796 1567
rect 872 1563 876 1567
rect 952 1563 956 1567
rect 1032 1563 1036 1567
rect 1104 1563 1108 1567
rect 1176 1563 1180 1567
rect 1256 1563 1260 1567
rect 1336 1563 1340 1567
rect 1416 1563 1420 1567
rect 1496 1563 1500 1567
rect 1560 1563 1564 1567
rect 192 1547 196 1551
rect 232 1547 236 1551
rect 272 1547 276 1551
rect 280 1547 284 1551
rect 312 1547 316 1551
rect 360 1547 364 1551
rect 408 1547 412 1551
rect 456 1547 460 1551
rect 504 1547 508 1551
rect 552 1547 556 1551
rect 600 1549 604 1553
rect 616 1551 620 1555
rect 656 1547 660 1551
rect 720 1547 724 1551
rect 792 1547 796 1551
rect 872 1547 876 1551
rect 952 1547 956 1551
rect 1032 1547 1036 1551
rect 1104 1547 1108 1551
rect 1176 1547 1180 1551
rect 1256 1547 1260 1551
rect 1336 1547 1340 1551
rect 1416 1547 1420 1551
rect 1496 1549 1500 1553
rect 1560 1547 1564 1551
rect 176 1535 180 1539
rect 224 1535 228 1539
rect 272 1537 276 1541
rect 1064 1539 1068 1543
rect 328 1535 332 1539
rect 344 1535 348 1539
rect 376 1535 380 1539
rect 432 1535 436 1539
rect 488 1535 492 1539
rect 544 1535 548 1539
rect 600 1535 604 1539
rect 656 1535 660 1539
rect 712 1535 716 1539
rect 776 1535 780 1539
rect 840 1535 844 1539
rect 912 1535 916 1539
rect 984 1535 988 1539
rect 1056 1535 1060 1539
rect 176 1519 180 1523
rect 224 1519 228 1523
rect 272 1521 276 1525
rect 280 1523 284 1527
rect 328 1519 332 1523
rect 440 1523 444 1527
rect 1120 1535 1124 1539
rect 1184 1535 1188 1539
rect 1248 1535 1252 1539
rect 1312 1535 1316 1539
rect 1376 1535 1380 1539
rect 1440 1535 1444 1539
rect 1512 1535 1516 1539
rect 1560 1535 1564 1539
rect 376 1519 380 1523
rect 432 1519 436 1523
rect 344 1507 348 1511
rect 176 1491 180 1495
rect 224 1491 228 1495
rect 272 1491 276 1495
rect 320 1491 324 1495
rect 368 1491 372 1495
rect 424 1491 428 1495
rect 488 1519 492 1523
rect 544 1519 548 1523
rect 600 1519 604 1523
rect 656 1519 660 1523
rect 712 1519 716 1523
rect 776 1519 780 1523
rect 840 1519 844 1523
rect 912 1519 916 1523
rect 984 1519 988 1523
rect 1056 1519 1060 1523
rect 1064 1519 1068 1523
rect 1120 1519 1124 1523
rect 1184 1519 1188 1523
rect 1248 1519 1252 1523
rect 1312 1519 1316 1523
rect 1376 1519 1380 1523
rect 1440 1519 1444 1523
rect 1512 1519 1516 1523
rect 1560 1519 1564 1523
rect 480 1491 484 1495
rect 544 1491 548 1495
rect 608 1491 612 1495
rect 672 1491 676 1495
rect 736 1491 740 1495
rect 800 1491 804 1495
rect 872 1491 876 1495
rect 952 1491 956 1495
rect 1024 1491 1028 1495
rect 1096 1491 1100 1495
rect 1168 1491 1172 1495
rect 1232 1491 1236 1495
rect 1296 1491 1300 1495
rect 1368 1491 1372 1495
rect 1440 1491 1444 1495
rect 1512 1491 1516 1495
rect 1560 1491 1564 1495
rect 176 1475 180 1479
rect 224 1475 228 1479
rect 272 1475 276 1479
rect 320 1475 324 1479
rect 368 1475 372 1479
rect 424 1475 428 1479
rect 440 1475 444 1479
rect 480 1475 484 1479
rect 544 1475 548 1479
rect 608 1475 612 1479
rect 672 1475 676 1479
rect 736 1475 740 1479
rect 800 1475 804 1479
rect 872 1475 876 1479
rect 952 1475 956 1479
rect 1024 1475 1028 1479
rect 1096 1475 1100 1479
rect 1168 1475 1172 1479
rect 1232 1475 1236 1479
rect 1296 1475 1300 1479
rect 1368 1475 1372 1479
rect 1440 1475 1444 1479
rect 1512 1475 1516 1479
rect 1560 1475 1564 1479
rect 600 1467 604 1471
rect 1424 1467 1428 1471
rect 152 1463 156 1467
rect 200 1463 204 1467
rect 248 1463 252 1467
rect 304 1463 308 1467
rect 360 1463 364 1467
rect 416 1463 420 1467
rect 472 1463 476 1467
rect 528 1463 532 1467
rect 592 1463 596 1467
rect 648 1463 652 1467
rect 704 1463 708 1467
rect 768 1463 772 1467
rect 832 1463 836 1467
rect 896 1463 900 1467
rect 960 1463 964 1467
rect 1032 1463 1036 1467
rect 1104 1463 1108 1467
rect 1176 1463 1180 1467
rect 1256 1463 1260 1467
rect 1336 1463 1340 1467
rect 1416 1463 1420 1467
rect 1496 1463 1500 1467
rect 1560 1463 1564 1467
rect 152 1447 156 1451
rect 200 1447 204 1451
rect 248 1447 252 1451
rect 304 1447 308 1451
rect 360 1447 364 1451
rect 416 1447 420 1451
rect 472 1447 476 1451
rect 528 1447 532 1451
rect 592 1447 596 1451
rect 600 1447 604 1451
rect 648 1447 652 1451
rect 704 1447 708 1451
rect 768 1447 772 1451
rect 832 1447 836 1451
rect 896 1447 900 1451
rect 960 1447 964 1451
rect 1032 1447 1036 1451
rect 1104 1447 1108 1451
rect 1176 1447 1180 1451
rect 1256 1447 1260 1451
rect 1336 1447 1340 1451
rect 1416 1447 1420 1451
rect 1424 1447 1428 1451
rect 1496 1447 1500 1451
rect 1560 1447 1564 1451
rect 152 1419 156 1423
rect 200 1419 204 1423
rect 272 1419 276 1423
rect 344 1419 348 1423
rect 416 1419 420 1423
rect 488 1419 492 1423
rect 560 1419 564 1423
rect 632 1419 636 1423
rect 696 1419 700 1423
rect 760 1419 764 1423
rect 832 1419 836 1423
rect 896 1419 900 1423
rect 968 1419 972 1423
rect 1040 1419 1044 1423
rect 1112 1419 1116 1423
rect 1176 1419 1180 1423
rect 1240 1419 1244 1423
rect 1304 1419 1308 1423
rect 1360 1419 1364 1423
rect 1416 1419 1420 1423
rect 1472 1419 1476 1423
rect 1528 1419 1532 1423
rect 1560 1419 1564 1423
rect 152 1403 156 1407
rect 200 1403 204 1407
rect 272 1403 276 1407
rect 344 1403 348 1407
rect 416 1403 420 1407
rect 488 1403 492 1407
rect 560 1403 564 1407
rect 632 1403 636 1407
rect 696 1403 700 1407
rect 760 1403 764 1407
rect 832 1403 836 1407
rect 896 1403 900 1407
rect 968 1405 972 1409
rect 1040 1403 1044 1407
rect 1112 1403 1116 1407
rect 1176 1403 1180 1407
rect 1240 1403 1244 1407
rect 1304 1403 1308 1407
rect 1360 1403 1364 1407
rect 1416 1403 1420 1407
rect 1472 1403 1476 1407
rect 1528 1403 1532 1407
rect 1560 1403 1564 1407
rect 1264 1395 1268 1399
rect 152 1391 156 1395
rect 192 1391 196 1395
rect 264 1391 268 1395
rect 336 1391 340 1395
rect 408 1391 412 1395
rect 472 1391 476 1395
rect 536 1391 540 1395
rect 600 1391 604 1395
rect 664 1391 668 1395
rect 728 1391 732 1395
rect 792 1391 796 1395
rect 856 1391 860 1395
rect 912 1391 916 1395
rect 968 1391 972 1395
rect 1016 1391 1020 1395
rect 1072 1391 1076 1395
rect 1128 1391 1132 1395
rect 1192 1391 1196 1395
rect 1256 1391 1260 1395
rect 1312 1391 1316 1395
rect 1368 1391 1372 1395
rect 1432 1391 1436 1395
rect 1496 1391 1500 1395
rect 1560 1391 1564 1395
rect 152 1375 156 1379
rect 192 1375 196 1379
rect 264 1375 268 1379
rect 336 1375 340 1379
rect 408 1375 412 1379
rect 472 1375 476 1379
rect 536 1375 540 1379
rect 600 1375 604 1379
rect 664 1375 668 1379
rect 728 1375 732 1379
rect 792 1375 796 1379
rect 856 1375 860 1379
rect 912 1375 916 1379
rect 968 1375 972 1379
rect 1016 1375 1020 1379
rect 1072 1375 1076 1379
rect 1128 1375 1132 1379
rect 1192 1375 1196 1379
rect 1256 1375 1260 1379
rect 1264 1375 1268 1379
rect 1312 1375 1316 1379
rect 1368 1375 1372 1379
rect 1432 1375 1436 1379
rect 1496 1375 1500 1379
rect 1560 1375 1564 1379
rect 1088 1363 1092 1367
rect 152 1347 156 1351
rect 184 1347 188 1351
rect 232 1347 236 1351
rect 320 1347 324 1351
rect 432 1347 436 1351
rect 544 1347 548 1351
rect 656 1347 660 1351
rect 768 1347 772 1351
rect 880 1347 884 1351
rect 984 1347 988 1351
rect 1080 1347 1084 1351
rect 1168 1347 1172 1351
rect 1248 1347 1252 1351
rect 1328 1347 1332 1351
rect 1400 1347 1404 1351
rect 1472 1347 1476 1351
rect 1552 1347 1556 1351
rect 152 1331 156 1335
rect 184 1331 188 1335
rect 232 1331 236 1335
rect 320 1331 324 1335
rect 432 1331 436 1335
rect 544 1331 548 1335
rect 656 1331 660 1335
rect 768 1331 772 1335
rect 880 1331 884 1335
rect 984 1331 988 1335
rect 1080 1331 1084 1335
rect 1088 1331 1092 1335
rect 1168 1331 1172 1335
rect 1248 1331 1252 1335
rect 1328 1331 1332 1335
rect 1400 1331 1404 1335
rect 1472 1331 1476 1335
rect 1552 1331 1556 1335
rect 152 1319 156 1323
rect 200 1319 204 1323
rect 264 1319 268 1323
rect 328 1319 332 1323
rect 392 1319 396 1323
rect 456 1319 460 1323
rect 512 1319 516 1323
rect 560 1319 564 1323
rect 608 1319 612 1323
rect 656 1319 660 1323
rect 704 1319 708 1323
rect 760 1319 764 1323
rect 808 1319 812 1323
rect 856 1319 860 1323
rect 904 1319 908 1323
rect 952 1319 956 1323
rect 1008 1319 1012 1323
rect 1064 1319 1068 1323
rect 1120 1319 1124 1323
rect 1176 1319 1180 1323
rect 1232 1319 1236 1323
rect 1288 1319 1292 1323
rect 1344 1319 1348 1323
rect 1392 1319 1396 1323
rect 1440 1319 1444 1323
rect 1488 1319 1492 1323
rect 1544 1319 1548 1323
rect 152 1303 156 1307
rect 200 1303 204 1307
rect 264 1303 268 1307
rect 328 1303 332 1307
rect 392 1303 396 1307
rect 456 1303 460 1307
rect 512 1303 516 1307
rect 560 1303 564 1307
rect 608 1303 612 1307
rect 656 1303 660 1307
rect 704 1303 708 1307
rect 760 1303 764 1307
rect 808 1303 812 1307
rect 856 1303 860 1307
rect 904 1303 908 1307
rect 952 1303 956 1307
rect 1008 1303 1012 1307
rect 1064 1303 1068 1307
rect 1120 1303 1124 1307
rect 1176 1303 1180 1307
rect 1232 1303 1236 1307
rect 1288 1303 1292 1307
rect 1344 1303 1348 1307
rect 1392 1303 1396 1307
rect 1440 1303 1444 1307
rect 1488 1303 1492 1307
rect 1544 1303 1548 1307
rect 696 1291 700 1295
rect 152 1275 156 1279
rect 208 1275 212 1279
rect 272 1275 276 1279
rect 344 1275 348 1279
rect 408 1275 412 1279
rect 480 1275 484 1279
rect 552 1275 556 1279
rect 616 1275 620 1279
rect 680 1275 684 1279
rect 744 1275 748 1279
rect 808 1275 812 1279
rect 872 1275 876 1279
rect 944 1275 948 1279
rect 1016 1275 1020 1279
rect 1080 1275 1084 1279
rect 1144 1275 1148 1279
rect 1208 1275 1212 1279
rect 1264 1275 1268 1279
rect 1320 1275 1324 1279
rect 1384 1275 1388 1279
rect 1448 1275 1452 1279
rect 152 1259 156 1263
rect 208 1259 212 1263
rect 272 1259 276 1263
rect 344 1259 348 1263
rect 408 1259 412 1263
rect 480 1259 484 1263
rect 552 1259 556 1263
rect 616 1259 620 1263
rect 680 1259 684 1263
rect 696 1259 700 1263
rect 744 1259 748 1263
rect 808 1259 812 1263
rect 872 1259 876 1263
rect 944 1259 948 1263
rect 1016 1259 1020 1263
rect 1080 1259 1084 1263
rect 1144 1259 1148 1263
rect 1208 1259 1212 1263
rect 1264 1259 1268 1263
rect 1320 1259 1324 1263
rect 1384 1259 1388 1263
rect 1448 1259 1452 1263
rect 152 1247 156 1251
rect 192 1247 196 1251
rect 248 1247 252 1251
rect 304 1247 308 1251
rect 368 1247 372 1251
rect 432 1247 436 1251
rect 496 1247 500 1251
rect 560 1247 564 1251
rect 624 1247 628 1251
rect 688 1247 692 1251
rect 752 1247 756 1251
rect 816 1247 820 1251
rect 880 1247 884 1251
rect 944 1247 948 1251
rect 1008 1247 1012 1251
rect 1032 1247 1036 1251
rect 1072 1247 1076 1251
rect 1136 1247 1140 1251
rect 1200 1247 1204 1251
rect 1264 1247 1268 1251
rect 1328 1247 1332 1251
rect 1392 1247 1396 1251
rect 1456 1247 1460 1251
rect 1520 1247 1524 1251
rect 1560 1247 1564 1251
rect 152 1231 156 1235
rect 192 1231 196 1235
rect 248 1231 252 1235
rect 304 1231 308 1235
rect 368 1231 372 1235
rect 432 1231 436 1235
rect 496 1231 500 1235
rect 560 1231 564 1235
rect 624 1231 628 1235
rect 688 1231 692 1235
rect 752 1231 756 1235
rect 816 1231 820 1235
rect 880 1231 884 1235
rect 944 1231 948 1235
rect 1008 1231 1012 1235
rect 1072 1231 1076 1235
rect 1136 1231 1140 1235
rect 1200 1231 1204 1235
rect 1264 1231 1268 1235
rect 1328 1231 1332 1235
rect 1392 1231 1396 1235
rect 1456 1231 1460 1235
rect 1520 1231 1524 1235
rect 1560 1231 1564 1235
rect 160 1203 164 1207
rect 192 1203 196 1207
rect 232 1203 236 1207
rect 280 1203 284 1207
rect 328 1203 332 1207
rect 376 1203 380 1207
rect 432 1203 436 1207
rect 488 1203 492 1207
rect 544 1203 548 1207
rect 600 1203 604 1207
rect 656 1203 660 1207
rect 704 1203 708 1207
rect 752 1203 756 1207
rect 800 1203 804 1207
rect 848 1203 852 1207
rect 896 1203 900 1207
rect 952 1203 956 1207
rect 1000 1203 1004 1207
rect 1032 1203 1036 1207
rect 1056 1203 1060 1207
rect 1064 1203 1068 1207
rect 1112 1203 1116 1207
rect 1176 1203 1180 1207
rect 1248 1203 1252 1207
rect 1320 1203 1324 1207
rect 1400 1203 1404 1207
rect 1488 1203 1492 1207
rect 1560 1203 1564 1207
rect 1568 1203 1572 1207
rect 160 1187 164 1191
rect 192 1187 196 1191
rect 232 1187 236 1191
rect 280 1187 284 1191
rect 328 1187 332 1191
rect 376 1187 380 1191
rect 432 1187 436 1191
rect 488 1187 492 1191
rect 544 1187 548 1191
rect 600 1187 604 1191
rect 656 1187 660 1191
rect 704 1187 708 1191
rect 752 1187 756 1191
rect 800 1187 804 1191
rect 848 1187 852 1191
rect 896 1187 900 1191
rect 952 1187 956 1191
rect 1000 1187 1004 1191
rect 1056 1187 1060 1191
rect 1112 1187 1116 1191
rect 1176 1187 1180 1191
rect 1248 1187 1252 1191
rect 1320 1187 1324 1191
rect 1400 1187 1404 1191
rect 1488 1187 1492 1191
rect 1560 1187 1564 1191
rect 160 1175 164 1179
rect 192 1175 196 1179
rect 232 1175 236 1179
rect 272 1175 276 1179
rect 288 1175 292 1179
rect 320 1175 324 1179
rect 376 1175 380 1179
rect 432 1175 436 1179
rect 488 1175 492 1179
rect 544 1175 548 1179
rect 608 1175 612 1179
rect 672 1175 676 1179
rect 736 1175 740 1179
rect 808 1175 812 1179
rect 872 1175 876 1179
rect 936 1175 940 1179
rect 1000 1175 1004 1179
rect 1056 1175 1060 1179
rect 1064 1175 1068 1179
rect 1120 1175 1124 1179
rect 1184 1175 1188 1179
rect 1256 1175 1260 1179
rect 1328 1175 1332 1179
rect 1408 1175 1412 1179
rect 1496 1175 1500 1179
rect 1560 1175 1564 1179
rect 1568 1175 1572 1179
rect 160 1159 164 1163
rect 192 1159 196 1163
rect 232 1159 236 1163
rect 272 1159 276 1163
rect 320 1159 324 1163
rect 376 1159 380 1163
rect 432 1159 436 1163
rect 488 1159 492 1163
rect 544 1159 548 1163
rect 608 1159 612 1163
rect 672 1159 676 1163
rect 736 1159 740 1163
rect 808 1159 812 1163
rect 872 1159 876 1163
rect 936 1159 940 1163
rect 1000 1159 1004 1163
rect 1056 1159 1060 1163
rect 1120 1159 1124 1163
rect 1184 1159 1188 1163
rect 1256 1159 1260 1163
rect 1328 1159 1332 1163
rect 1408 1159 1412 1163
rect 1496 1159 1500 1163
rect 1560 1159 1564 1163
rect 288 1147 292 1151
rect 152 1131 156 1135
rect 184 1131 188 1135
rect 216 1131 220 1135
rect 248 1131 252 1135
rect 280 1131 284 1135
rect 312 1131 316 1135
rect 344 1131 348 1135
rect 376 1131 380 1135
rect 408 1131 412 1135
rect 464 1131 468 1135
rect 520 1131 524 1135
rect 576 1131 580 1135
rect 632 1131 636 1135
rect 688 1131 692 1135
rect 744 1131 748 1135
rect 800 1131 804 1135
rect 856 1131 860 1135
rect 912 1131 916 1135
rect 968 1131 972 1135
rect 1024 1131 1028 1135
rect 1080 1131 1084 1135
rect 1144 1131 1148 1135
rect 1208 1131 1212 1135
rect 1272 1131 1276 1135
rect 1344 1131 1348 1135
rect 1416 1131 1420 1135
rect 1496 1131 1500 1135
rect 1560 1131 1564 1135
rect 1568 1131 1572 1135
rect 152 1115 156 1119
rect 184 1115 188 1119
rect 216 1115 220 1119
rect 248 1115 252 1119
rect 280 1115 284 1119
rect 312 1115 316 1119
rect 344 1115 348 1119
rect 376 1115 380 1119
rect 408 1115 412 1119
rect 464 1115 468 1119
rect 520 1115 524 1119
rect 576 1115 580 1119
rect 632 1115 636 1119
rect 688 1115 692 1119
rect 744 1115 748 1119
rect 800 1115 804 1119
rect 856 1115 860 1119
rect 912 1115 916 1119
rect 968 1115 972 1119
rect 1024 1115 1028 1119
rect 1080 1115 1084 1119
rect 1144 1115 1148 1119
rect 1208 1115 1212 1119
rect 1272 1115 1276 1119
rect 1344 1115 1348 1119
rect 1416 1115 1420 1119
rect 1496 1115 1500 1119
rect 1560 1115 1564 1119
rect 168 1103 172 1107
rect 200 1103 204 1107
rect 240 1103 244 1107
rect 288 1103 292 1107
rect 344 1103 348 1107
rect 400 1103 404 1107
rect 456 1103 460 1107
rect 520 1103 524 1107
rect 584 1103 588 1107
rect 656 1103 660 1107
rect 728 1103 732 1107
rect 800 1103 804 1107
rect 872 1103 876 1107
rect 936 1103 940 1107
rect 1000 1103 1004 1107
rect 1056 1103 1060 1107
rect 1112 1103 1116 1107
rect 1168 1103 1172 1107
rect 1224 1103 1228 1107
rect 1280 1103 1284 1107
rect 1336 1103 1340 1107
rect 1392 1103 1396 1107
rect 1456 1103 1460 1107
rect 1520 1103 1524 1107
rect 1560 1103 1564 1107
rect 1568 1103 1572 1107
rect 168 1087 172 1091
rect 200 1087 204 1091
rect 240 1087 244 1091
rect 288 1087 292 1091
rect 344 1087 348 1091
rect 400 1087 404 1091
rect 456 1087 460 1091
rect 520 1087 524 1091
rect 584 1087 588 1091
rect 656 1087 660 1091
rect 728 1087 732 1091
rect 800 1087 804 1091
rect 872 1087 876 1091
rect 936 1087 940 1091
rect 1000 1087 1004 1091
rect 1056 1087 1060 1091
rect 1112 1087 1116 1091
rect 1168 1087 1172 1091
rect 1224 1087 1228 1091
rect 1280 1087 1284 1091
rect 1336 1087 1340 1091
rect 1392 1087 1396 1091
rect 1456 1087 1460 1091
rect 1520 1087 1524 1091
rect 1560 1087 1564 1091
rect 464 1051 468 1055
rect 504 1051 508 1055
rect 560 1051 564 1055
rect 616 1051 620 1055
rect 680 1051 684 1055
rect 744 1051 748 1055
rect 808 1051 812 1055
rect 880 1051 884 1055
rect 952 1051 956 1055
rect 1024 1051 1028 1055
rect 1096 1051 1100 1055
rect 1168 1051 1172 1055
rect 1232 1051 1236 1055
rect 1296 1051 1300 1055
rect 1352 1051 1356 1055
rect 1408 1051 1412 1055
rect 1464 1051 1468 1055
rect 1520 1051 1524 1055
rect 1560 1051 1564 1055
rect 464 1035 468 1039
rect 472 1035 476 1039
rect 504 1035 508 1039
rect 560 1035 564 1039
rect 616 1035 620 1039
rect 680 1035 684 1039
rect 744 1035 748 1039
rect 808 1035 812 1039
rect 880 1035 884 1039
rect 952 1035 956 1039
rect 1024 1035 1028 1039
rect 1096 1035 1100 1039
rect 1168 1035 1172 1039
rect 1232 1035 1236 1039
rect 1296 1035 1300 1039
rect 1352 1035 1356 1039
rect 1408 1035 1412 1039
rect 1464 1035 1468 1039
rect 1520 1035 1524 1039
rect 1560 1035 1564 1039
rect 528 1019 532 1023
rect 560 1019 564 1023
rect 592 1019 596 1023
rect 632 1019 636 1023
rect 680 1019 684 1023
rect 728 1019 732 1023
rect 792 1019 796 1023
rect 864 1019 868 1023
rect 944 1019 948 1023
rect 1024 1019 1028 1023
rect 1104 1019 1108 1023
rect 1184 1019 1188 1023
rect 1256 1019 1260 1023
rect 1320 1019 1324 1023
rect 1376 1019 1380 1023
rect 1424 1019 1428 1023
rect 1472 1019 1476 1023
rect 1528 1019 1532 1023
rect 1560 1019 1564 1023
rect 472 1007 476 1011
rect 528 1003 532 1007
rect 560 1003 564 1007
rect 592 1003 596 1007
rect 632 1003 636 1007
rect 680 1003 684 1007
rect 728 1003 732 1007
rect 792 1003 796 1007
rect 864 1003 868 1007
rect 944 1003 948 1007
rect 1024 1003 1028 1007
rect 1104 1003 1108 1007
rect 1184 1003 1188 1007
rect 1256 1003 1260 1007
rect 1320 1003 1324 1007
rect 1376 1003 1380 1007
rect 1424 1003 1428 1007
rect 1472 1003 1476 1007
rect 1528 1003 1532 1007
rect 1560 1003 1564 1007
rect 176 967 180 971
rect 216 967 220 971
rect 272 967 276 971
rect 328 967 332 971
rect 392 967 396 971
rect 456 967 460 971
rect 520 967 524 971
rect 576 967 580 971
rect 632 967 636 971
rect 680 967 684 971
rect 720 967 724 971
rect 752 967 756 971
rect 792 967 796 971
rect 848 967 852 971
rect 912 967 916 971
rect 984 967 988 971
rect 1064 967 1068 971
rect 1144 967 1148 971
rect 1216 967 1220 971
rect 1288 967 1292 971
rect 1360 967 1364 971
rect 1432 967 1436 971
rect 1504 967 1508 971
rect 1560 967 1564 971
rect 1568 967 1572 971
rect 176 951 180 955
rect 216 951 220 955
rect 272 951 276 955
rect 328 951 332 955
rect 392 951 396 955
rect 456 951 460 955
rect 520 951 524 955
rect 576 951 580 955
rect 632 951 636 955
rect 680 951 684 955
rect 720 951 724 955
rect 752 951 756 955
rect 792 951 796 955
rect 848 951 852 955
rect 912 951 916 955
rect 984 951 988 955
rect 1064 951 1068 955
rect 1144 951 1148 955
rect 1216 951 1220 955
rect 1288 951 1292 955
rect 1360 951 1364 955
rect 1432 951 1436 955
rect 1504 951 1508 955
rect 1560 951 1564 955
rect 168 939 172 943
rect 208 939 212 943
rect 264 939 268 943
rect 320 939 324 943
rect 384 939 388 943
rect 448 939 452 943
rect 512 939 516 943
rect 576 939 580 943
rect 632 939 636 943
rect 688 939 692 943
rect 736 939 740 943
rect 784 939 788 943
rect 832 939 836 943
rect 888 939 892 943
rect 952 939 956 943
rect 1024 939 1028 943
rect 1096 939 1100 943
rect 1160 939 1164 943
rect 1224 939 1228 943
rect 1288 939 1292 943
rect 1344 939 1348 943
rect 1392 939 1396 943
rect 1400 939 1404 943
rect 1440 939 1444 943
rect 1488 939 1492 943
rect 1528 939 1532 943
rect 1560 939 1564 943
rect 1568 939 1572 943
rect 168 923 172 927
rect 208 923 212 927
rect 264 923 268 927
rect 320 923 324 927
rect 384 923 388 927
rect 448 923 452 927
rect 512 923 516 927
rect 576 923 580 927
rect 632 923 636 927
rect 688 923 692 927
rect 736 923 740 927
rect 784 923 788 927
rect 832 923 836 927
rect 888 923 892 927
rect 952 923 956 927
rect 1024 923 1028 927
rect 1096 923 1100 927
rect 1160 923 1164 927
rect 1224 923 1228 927
rect 1288 923 1292 927
rect 1344 923 1348 927
rect 1392 923 1396 927
rect 848 911 852 915
rect 152 891 156 895
rect 184 891 188 895
rect 240 891 244 895
rect 296 891 300 895
rect 352 891 356 895
rect 408 891 412 895
rect 464 891 468 895
rect 520 891 524 895
rect 576 891 580 895
rect 640 891 644 895
rect 712 891 716 895
rect 776 891 780 895
rect 840 891 844 895
rect 152 875 156 879
rect 184 875 188 879
rect 240 875 244 879
rect 296 875 300 879
rect 352 875 356 879
rect 408 875 412 879
rect 464 875 468 879
rect 520 875 524 879
rect 576 875 580 879
rect 640 875 644 879
rect 712 875 716 879
rect 776 875 780 879
rect 840 875 844 879
rect 848 875 852 879
rect 872 903 876 907
rect 368 867 372 871
rect 1440 923 1444 927
rect 1488 923 1492 927
rect 1528 923 1532 927
rect 1560 923 1564 927
rect 904 891 908 895
rect 968 891 972 895
rect 1032 891 1036 895
rect 1096 891 1100 895
rect 1152 891 1156 895
rect 1208 891 1212 895
rect 1264 891 1268 895
rect 1320 891 1324 895
rect 1376 891 1380 895
rect 1400 891 1404 895
rect 1424 891 1428 895
rect 1472 891 1476 895
rect 1528 891 1532 895
rect 1560 891 1564 895
rect 904 875 908 879
rect 968 875 972 879
rect 1032 875 1036 879
rect 1096 875 1100 879
rect 1152 875 1156 879
rect 1208 875 1212 879
rect 1264 875 1268 879
rect 1320 875 1324 879
rect 1376 875 1380 879
rect 1424 875 1428 879
rect 1472 875 1476 879
rect 1528 875 1532 879
rect 1560 875 1564 879
rect 152 863 156 867
rect 184 863 188 867
rect 224 863 228 867
rect 272 863 276 867
rect 320 863 324 867
rect 360 863 364 867
rect 400 863 404 867
rect 416 863 420 867
rect 456 863 460 867
rect 528 863 532 867
rect 608 863 612 867
rect 696 863 700 867
rect 784 863 788 867
rect 864 863 868 867
rect 872 863 876 867
rect 936 863 940 867
rect 1000 863 1004 867
rect 1056 863 1060 867
rect 1112 863 1116 867
rect 1168 863 1172 867
rect 1224 863 1228 867
rect 1240 863 1244 867
rect 1280 863 1284 867
rect 1344 863 1348 867
rect 1416 863 1420 867
rect 1496 863 1500 867
rect 1560 863 1564 867
rect 152 847 156 851
rect 184 847 188 851
rect 224 847 228 851
rect 272 847 276 851
rect 320 847 324 851
rect 360 847 364 851
rect 368 847 372 851
rect 400 847 404 851
rect 1128 851 1132 855
rect 456 847 460 851
rect 528 847 532 851
rect 608 847 612 851
rect 696 847 700 851
rect 784 847 788 851
rect 864 847 868 851
rect 936 847 940 851
rect 1000 847 1004 851
rect 1056 847 1060 851
rect 1112 847 1116 851
rect 448 831 452 835
rect 152 815 156 819
rect 184 815 188 819
rect 240 815 244 819
rect 304 815 308 819
rect 368 815 372 819
rect 416 815 420 819
rect 440 815 444 819
rect 152 799 156 803
rect 184 799 188 803
rect 240 799 244 803
rect 304 799 308 803
rect 368 799 372 803
rect 440 799 444 803
rect 512 815 516 819
rect 584 815 588 819
rect 656 815 660 819
rect 736 815 740 819
rect 808 815 812 819
rect 880 815 884 819
rect 952 815 956 819
rect 1016 815 1020 819
rect 1072 815 1076 819
rect 1120 815 1124 819
rect 1168 847 1172 851
rect 1224 847 1228 851
rect 1280 847 1284 851
rect 1344 847 1348 851
rect 1416 847 1420 851
rect 1496 847 1500 851
rect 1560 847 1564 851
rect 1240 835 1244 839
rect 1160 815 1164 819
rect 1200 815 1204 819
rect 1248 815 1252 819
rect 1296 815 1300 819
rect 1344 815 1348 819
rect 512 799 516 803
rect 584 799 588 803
rect 656 799 660 803
rect 736 799 740 803
rect 808 799 812 803
rect 880 799 884 803
rect 952 799 956 803
rect 1016 799 1020 803
rect 1072 799 1076 803
rect 1120 799 1124 803
rect 1128 799 1132 803
rect 1160 799 1164 803
rect 1200 799 1204 803
rect 1248 799 1252 803
rect 1296 799 1300 803
rect 1344 799 1348 803
rect 224 791 228 795
rect 328 791 332 795
rect 152 787 156 791
rect 184 787 188 791
rect 216 787 220 791
rect 152 771 156 775
rect 184 771 188 775
rect 216 771 220 775
rect 264 787 268 791
rect 320 787 324 791
rect 376 787 380 791
rect 440 789 444 793
rect 448 791 452 795
rect 760 791 764 795
rect 504 787 508 791
rect 568 787 572 791
rect 624 787 628 791
rect 688 787 692 791
rect 752 787 756 791
rect 816 787 820 791
rect 888 787 892 791
rect 952 787 956 791
rect 1016 787 1020 791
rect 1080 787 1084 791
rect 1144 787 1148 791
rect 1208 787 1212 791
rect 1272 787 1276 791
rect 1336 787 1340 791
rect 1400 787 1404 791
rect 264 771 268 775
rect 320 771 324 775
rect 328 771 332 775
rect 376 771 380 775
rect 440 771 444 775
rect 504 771 508 775
rect 568 771 572 775
rect 624 771 628 775
rect 688 771 692 775
rect 752 771 756 775
rect 760 771 764 775
rect 816 771 820 775
rect 888 771 892 775
rect 952 771 956 775
rect 1016 771 1020 775
rect 1080 771 1084 775
rect 1144 771 1148 775
rect 1208 771 1212 775
rect 1272 771 1276 775
rect 1336 771 1340 775
rect 1400 771 1404 775
rect 152 743 156 747
rect 184 743 188 747
rect 216 743 220 747
rect 224 743 228 747
rect 272 743 276 747
rect 336 743 340 747
rect 408 743 412 747
rect 480 743 484 747
rect 560 743 564 747
rect 640 743 644 747
rect 720 743 724 747
rect 792 743 796 747
rect 864 743 868 747
rect 936 743 940 747
rect 1008 743 1012 747
rect 1080 743 1084 747
rect 1152 743 1156 747
rect 1224 743 1228 747
rect 1288 743 1292 747
rect 1344 743 1348 747
rect 1392 743 1396 747
rect 1440 743 1444 747
rect 1488 743 1492 747
rect 1528 743 1532 747
rect 1560 743 1564 747
rect 152 727 156 731
rect 184 727 188 731
rect 216 727 220 731
rect 272 727 276 731
rect 336 727 340 731
rect 408 727 412 731
rect 480 727 484 731
rect 560 727 564 731
rect 640 727 644 731
rect 720 727 724 731
rect 792 727 796 731
rect 864 727 868 731
rect 936 727 940 731
rect 1008 727 1012 731
rect 1080 727 1084 731
rect 1152 727 1156 731
rect 1224 727 1228 731
rect 1288 727 1292 731
rect 1344 727 1348 731
rect 1392 727 1396 731
rect 1440 727 1444 731
rect 1488 727 1492 731
rect 1528 727 1532 731
rect 1560 727 1564 731
rect 152 715 156 719
rect 184 715 188 719
rect 224 715 228 719
rect 272 715 276 719
rect 328 715 332 719
rect 384 715 388 719
rect 440 715 444 719
rect 496 715 500 719
rect 560 715 564 719
rect 632 715 636 719
rect 704 715 708 719
rect 776 715 780 719
rect 856 715 860 719
rect 936 715 940 719
rect 1024 715 1028 719
rect 1104 715 1108 719
rect 1184 715 1188 719
rect 1256 715 1260 719
rect 1320 715 1324 719
rect 1376 715 1380 719
rect 1424 715 1428 719
rect 1472 715 1476 719
rect 1528 715 1532 719
rect 1560 715 1564 719
rect 152 699 156 703
rect 184 699 188 703
rect 224 699 228 703
rect 272 699 276 703
rect 328 699 332 703
rect 384 699 388 703
rect 440 699 444 703
rect 496 699 500 703
rect 560 699 564 703
rect 632 699 636 703
rect 704 699 708 703
rect 776 699 780 703
rect 856 699 860 703
rect 936 699 940 703
rect 1024 699 1028 703
rect 1104 699 1108 703
rect 1184 699 1188 703
rect 1256 699 1260 703
rect 1320 699 1324 703
rect 1376 699 1380 703
rect 1424 699 1428 703
rect 1472 701 1476 705
rect 1528 699 1532 703
rect 1560 699 1564 703
rect 176 671 180 675
rect 224 671 228 675
rect 272 671 276 675
rect 320 671 324 675
rect 376 671 380 675
rect 432 671 436 675
rect 488 671 492 675
rect 544 671 548 675
rect 600 671 604 675
rect 656 671 660 675
rect 712 671 716 675
rect 776 671 780 675
rect 840 671 844 675
rect 904 671 908 675
rect 968 671 972 675
rect 1032 671 1036 675
rect 1096 671 1100 675
rect 1152 671 1156 675
rect 1208 671 1212 675
rect 1264 671 1268 675
rect 1320 671 1324 675
rect 1376 671 1380 675
rect 176 655 180 659
rect 224 655 228 659
rect 272 655 276 659
rect 320 655 324 659
rect 376 655 380 659
rect 432 655 436 659
rect 488 655 492 659
rect 544 655 548 659
rect 600 655 604 659
rect 656 655 660 659
rect 712 655 716 659
rect 776 655 780 659
rect 840 655 844 659
rect 904 655 908 659
rect 968 655 972 659
rect 1032 655 1036 659
rect 1096 655 1100 659
rect 1152 655 1156 659
rect 1208 655 1212 659
rect 1264 655 1268 659
rect 1320 655 1324 659
rect 1376 655 1380 659
rect 184 639 188 643
rect 232 639 236 643
rect 288 639 292 643
rect 344 639 348 643
rect 400 639 404 643
rect 448 639 452 643
rect 504 639 508 643
rect 552 639 556 643
rect 608 639 612 643
rect 664 639 668 643
rect 720 639 724 643
rect 776 639 780 643
rect 840 639 844 643
rect 904 639 908 643
rect 960 639 964 643
rect 1016 639 1020 643
rect 1072 639 1076 643
rect 1128 639 1132 643
rect 1184 639 1188 643
rect 1232 639 1236 643
rect 1288 639 1292 643
rect 1344 639 1348 643
rect 1400 639 1404 643
rect 1456 639 1460 643
rect 1520 639 1524 643
rect 1560 639 1564 643
rect 184 623 188 627
rect 232 623 236 627
rect 288 623 292 627
rect 344 623 348 627
rect 400 623 404 627
rect 448 623 452 627
rect 504 623 508 627
rect 552 623 556 627
rect 608 623 612 627
rect 664 623 668 627
rect 720 623 724 627
rect 776 623 780 627
rect 840 623 844 627
rect 904 623 908 627
rect 960 623 964 627
rect 1016 623 1020 627
rect 1072 623 1076 627
rect 1128 623 1132 627
rect 1184 623 1188 627
rect 1232 623 1236 627
rect 1288 623 1292 627
rect 1344 623 1348 627
rect 1400 623 1404 627
rect 1456 623 1460 627
rect 1520 623 1524 627
rect 1560 623 1564 627
rect 240 595 244 599
rect 272 595 276 599
rect 304 595 308 599
rect 336 597 340 601
rect 368 595 372 599
rect 400 595 404 599
rect 440 595 444 599
rect 480 595 484 599
rect 536 595 540 599
rect 600 595 604 599
rect 664 595 668 599
rect 736 595 740 599
rect 816 595 820 599
rect 904 595 908 599
rect 992 595 996 599
rect 1080 595 1084 599
rect 1160 595 1164 599
rect 1232 595 1236 599
rect 1304 595 1308 599
rect 1368 595 1372 599
rect 1424 595 1428 599
rect 1472 595 1476 599
rect 1528 595 1532 599
rect 1560 595 1564 599
rect 1568 595 1572 599
rect 240 579 244 583
rect 272 579 276 583
rect 304 579 308 583
rect 336 579 340 583
rect 368 579 372 583
rect 400 579 404 583
rect 440 579 444 583
rect 480 579 484 583
rect 536 579 540 583
rect 600 579 604 583
rect 664 579 668 583
rect 736 579 740 583
rect 816 579 820 583
rect 864 579 868 583
rect 904 579 908 583
rect 992 579 996 583
rect 1080 579 1084 583
rect 1160 579 1164 583
rect 1232 581 1236 585
rect 1304 579 1308 583
rect 1368 579 1372 583
rect 1424 579 1428 583
rect 1472 579 1476 583
rect 1528 579 1532 583
rect 1560 579 1564 583
rect 280 571 284 575
rect 448 571 452 575
rect 208 567 212 571
rect 272 567 276 571
rect 344 567 348 571
rect 416 567 420 571
rect 208 551 212 555
rect 272 551 276 555
rect 280 551 284 555
rect 344 551 348 555
rect 416 551 420 555
rect 488 567 492 571
rect 552 567 556 571
rect 616 567 620 571
rect 680 567 684 571
rect 744 567 748 571
rect 800 567 804 571
rect 856 567 860 571
rect 920 567 924 571
rect 984 567 988 571
rect 1056 567 1060 571
rect 1120 567 1124 571
rect 1184 567 1188 571
rect 1248 567 1252 571
rect 1304 567 1308 571
rect 1352 567 1356 571
rect 1400 567 1404 571
rect 1440 567 1444 571
rect 1488 567 1492 571
rect 1528 569 1532 573
rect 1560 567 1564 571
rect 1568 567 1572 571
rect 1192 555 1196 559
rect 488 551 492 555
rect 552 551 556 555
rect 616 551 620 555
rect 680 551 684 555
rect 744 551 748 555
rect 800 551 804 555
rect 856 551 860 555
rect 864 551 868 555
rect 920 551 924 555
rect 952 551 956 555
rect 984 551 988 555
rect 1056 551 1060 555
rect 1120 551 1124 555
rect 1184 551 1188 555
rect 152 523 156 527
rect 192 523 196 527
rect 248 523 252 527
rect 312 523 316 527
rect 376 523 380 527
rect 440 523 444 527
rect 448 523 452 527
rect 496 523 500 527
rect 560 523 564 527
rect 616 523 620 527
rect 672 523 676 527
rect 728 523 732 527
rect 784 523 788 527
rect 792 523 796 527
rect 848 523 852 527
rect 912 523 916 527
rect 152 507 156 511
rect 192 507 196 511
rect 248 507 252 511
rect 312 507 316 511
rect 376 507 380 511
rect 440 507 444 511
rect 496 507 500 511
rect 560 507 564 511
rect 616 507 620 511
rect 672 507 676 511
rect 728 507 732 511
rect 784 507 788 511
rect 984 523 988 527
rect 1048 523 1052 527
rect 1112 523 1116 527
rect 1184 523 1188 527
rect 1248 551 1252 555
rect 1304 551 1308 555
rect 1352 551 1356 555
rect 1400 551 1404 555
rect 1440 551 1444 555
rect 1488 551 1492 555
rect 1528 551 1532 555
rect 1560 551 1564 555
rect 1256 523 1260 527
rect 1328 523 1332 527
rect 1408 523 1412 527
rect 1472 523 1476 527
rect 1496 523 1500 527
rect 1560 523 1564 527
rect 1568 523 1572 527
rect 848 507 852 511
rect 912 507 916 511
rect 952 507 956 511
rect 984 507 988 511
rect 1048 507 1052 511
rect 1112 507 1116 511
rect 1184 507 1188 511
rect 1192 507 1196 511
rect 1256 507 1260 511
rect 1328 507 1332 511
rect 1408 507 1412 511
rect 1496 507 1500 511
rect 1560 507 1564 511
rect 152 495 156 499
rect 184 495 188 499
rect 216 495 220 499
rect 264 495 268 499
rect 312 495 316 499
rect 360 495 364 499
rect 416 495 420 499
rect 472 495 476 499
rect 528 495 532 499
rect 584 495 588 499
rect 640 495 644 499
rect 696 495 700 499
rect 760 495 764 499
rect 792 495 796 499
rect 832 495 836 499
rect 904 495 908 499
rect 976 495 980 499
rect 1056 495 1060 499
rect 1144 495 1148 499
rect 1240 495 1244 499
rect 1344 495 1348 499
rect 1456 495 1460 499
rect 1472 495 1476 499
rect 1560 495 1564 499
rect 152 479 156 483
rect 184 479 188 483
rect 216 479 220 483
rect 264 479 268 483
rect 312 479 316 483
rect 360 479 364 483
rect 416 479 420 483
rect 472 479 476 483
rect 528 479 532 483
rect 584 479 588 483
rect 640 479 644 483
rect 696 479 700 483
rect 760 479 764 483
rect 832 479 836 483
rect 904 479 908 483
rect 976 479 980 483
rect 1056 479 1060 483
rect 1144 479 1148 483
rect 1240 479 1244 483
rect 1344 479 1348 483
rect 1456 479 1460 483
rect 1560 479 1564 483
rect 152 451 156 455
rect 184 451 188 455
rect 216 451 220 455
rect 272 451 276 455
rect 328 451 332 455
rect 384 451 388 455
rect 440 451 444 455
rect 496 451 500 455
rect 552 451 556 455
rect 616 451 620 455
rect 680 451 684 455
rect 752 451 756 455
rect 824 451 828 455
rect 888 451 892 455
rect 952 451 956 455
rect 1008 451 1012 455
rect 1064 451 1068 455
rect 1112 451 1116 455
rect 1160 451 1164 455
rect 1216 451 1220 455
rect 1280 451 1284 455
rect 1344 451 1348 455
rect 1416 451 1420 455
rect 1496 451 1500 455
rect 1560 451 1564 455
rect 152 435 156 439
rect 184 435 188 439
rect 216 435 220 439
rect 272 435 276 439
rect 328 435 332 439
rect 384 435 388 439
rect 440 435 444 439
rect 496 435 500 439
rect 552 435 556 439
rect 616 435 620 439
rect 680 435 684 439
rect 752 435 756 439
rect 824 435 828 439
rect 888 435 892 439
rect 952 435 956 439
rect 1008 435 1012 439
rect 1064 435 1068 439
rect 1112 435 1116 439
rect 1160 435 1164 439
rect 1216 435 1220 439
rect 1280 435 1284 439
rect 1344 435 1348 439
rect 1416 435 1420 439
rect 1496 435 1500 439
rect 1560 435 1564 439
rect 1568 435 1572 439
rect 152 419 156 423
rect 184 419 188 423
rect 248 419 252 423
rect 312 419 316 423
rect 376 419 380 423
rect 440 419 444 423
rect 456 419 460 423
rect 504 419 508 423
rect 560 419 564 423
rect 608 419 612 423
rect 656 419 660 423
rect 696 419 700 423
rect 736 419 740 423
rect 744 419 748 423
rect 776 419 780 423
rect 824 419 828 423
rect 880 419 884 423
rect 936 419 940 423
rect 992 419 996 423
rect 1048 419 1052 423
rect 1104 419 1108 423
rect 1168 419 1172 423
rect 1240 419 1244 423
rect 1320 419 1324 423
rect 1400 419 1404 423
rect 1488 419 1492 423
rect 1560 419 1564 423
rect 152 403 156 407
rect 184 403 188 407
rect 248 403 252 407
rect 312 403 316 407
rect 376 403 380 407
rect 440 403 444 407
rect 504 403 508 407
rect 560 403 564 407
rect 608 403 612 407
rect 656 403 660 407
rect 696 403 700 407
rect 736 403 740 407
rect 776 403 780 407
rect 824 403 828 407
rect 880 403 884 407
rect 936 403 940 407
rect 992 403 996 407
rect 1048 403 1052 407
rect 1104 403 1108 407
rect 1168 403 1172 407
rect 1240 403 1244 407
rect 1320 403 1324 407
rect 1400 403 1404 407
rect 1488 403 1492 407
rect 1560 403 1564 407
rect 152 375 156 379
rect 224 375 228 379
rect 312 375 316 379
rect 400 375 404 379
rect 456 375 460 379
rect 480 375 484 379
rect 552 375 556 379
rect 616 375 620 379
rect 672 375 676 379
rect 720 375 724 379
rect 744 375 748 379
rect 768 375 772 379
rect 824 375 828 379
rect 880 375 884 379
rect 936 375 940 379
rect 1000 375 1004 379
rect 1072 375 1076 379
rect 1144 375 1148 379
rect 1216 375 1220 379
rect 1288 375 1292 379
rect 1360 375 1364 379
rect 1432 375 1436 379
rect 1504 375 1508 379
rect 1560 375 1564 379
rect 1568 375 1572 379
rect 152 359 156 363
rect 224 359 228 363
rect 312 359 316 363
rect 400 359 404 363
rect 480 359 484 363
rect 552 359 556 363
rect 616 359 620 363
rect 672 359 676 363
rect 720 359 724 363
rect 768 359 772 363
rect 824 359 828 363
rect 880 359 884 363
rect 936 359 940 363
rect 1000 359 1004 363
rect 1072 359 1076 363
rect 1144 359 1148 363
rect 1216 359 1220 363
rect 1288 359 1292 363
rect 1360 359 1364 363
rect 1432 359 1436 363
rect 1504 359 1508 363
rect 1560 359 1564 363
rect 152 347 156 351
rect 192 347 196 351
rect 240 347 244 351
rect 296 347 300 351
rect 352 347 356 351
rect 408 347 412 351
rect 464 347 468 351
rect 520 347 524 351
rect 584 347 588 351
rect 648 347 652 351
rect 704 347 708 351
rect 768 347 772 351
rect 832 347 836 351
rect 896 347 900 351
rect 968 347 972 351
rect 1048 347 1052 351
rect 1120 347 1124 351
rect 1192 347 1196 351
rect 1264 347 1268 351
rect 1344 347 1348 351
rect 1424 347 1428 351
rect 1504 347 1508 351
rect 1560 347 1564 351
rect 1568 347 1572 351
rect 152 331 156 335
rect 192 331 196 335
rect 240 331 244 335
rect 296 331 300 335
rect 352 331 356 335
rect 408 331 412 335
rect 464 331 468 335
rect 520 331 524 335
rect 584 331 588 335
rect 648 331 652 335
rect 704 331 708 335
rect 768 331 772 335
rect 832 331 836 335
rect 896 331 900 335
rect 968 331 972 335
rect 1048 331 1052 335
rect 1120 331 1124 335
rect 1192 331 1196 335
rect 1264 331 1268 335
rect 1344 331 1348 335
rect 1424 331 1428 335
rect 1504 331 1508 335
rect 1560 331 1564 335
rect 208 303 212 307
rect 240 303 244 307
rect 272 303 276 307
rect 312 303 316 307
rect 352 303 356 307
rect 384 303 388 307
rect 424 303 428 307
rect 472 303 476 307
rect 536 303 540 307
rect 608 303 612 307
rect 680 303 684 307
rect 752 303 756 307
rect 824 303 828 307
rect 896 303 900 307
rect 968 303 972 307
rect 1040 303 1044 307
rect 1112 303 1116 307
rect 1184 303 1188 307
rect 1248 303 1252 307
rect 1312 303 1316 307
rect 1368 303 1372 307
rect 1416 303 1420 307
rect 1472 303 1476 307
rect 1528 303 1532 307
rect 1560 303 1564 307
rect 208 287 212 291
rect 240 287 244 291
rect 272 287 276 291
rect 312 287 316 291
rect 352 287 356 291
rect 384 287 388 291
rect 424 287 428 291
rect 472 287 476 291
rect 536 287 540 291
rect 608 287 612 291
rect 680 287 684 291
rect 752 287 756 291
rect 824 287 828 291
rect 896 287 900 291
rect 968 287 972 291
rect 1040 287 1044 291
rect 1112 287 1116 291
rect 1184 287 1188 291
rect 1248 287 1252 291
rect 1312 287 1316 291
rect 1368 287 1372 291
rect 1384 287 1388 291
rect 1416 287 1420 291
rect 1472 287 1476 291
rect 1528 287 1532 291
rect 1560 287 1564 291
rect 1144 275 1148 279
rect 1328 275 1332 279
rect 168 271 172 275
rect 200 271 204 275
rect 232 271 236 275
rect 264 271 268 275
rect 296 271 300 275
rect 328 271 332 275
rect 368 271 372 275
rect 424 271 428 275
rect 496 271 500 275
rect 576 271 580 275
rect 664 271 668 275
rect 752 271 756 275
rect 840 271 844 275
rect 920 271 924 275
rect 1000 271 1004 275
rect 1072 271 1076 275
rect 1136 271 1140 275
rect 1192 271 1196 275
rect 1240 271 1244 275
rect 1280 271 1284 275
rect 1320 271 1324 275
rect 1368 271 1372 275
rect 1416 271 1420 275
rect 1464 271 1468 275
rect 1520 271 1524 275
rect 1560 271 1564 275
rect 1384 259 1388 263
rect 168 255 172 259
rect 200 255 204 259
rect 232 255 236 259
rect 264 255 268 259
rect 296 255 300 259
rect 328 255 332 259
rect 368 255 372 259
rect 424 255 428 259
rect 496 255 500 259
rect 576 255 580 259
rect 664 255 668 259
rect 752 255 756 259
rect 840 255 844 259
rect 920 255 924 259
rect 1000 255 1004 259
rect 1072 255 1076 259
rect 1136 255 1140 259
rect 1144 255 1148 259
rect 1192 255 1196 259
rect 1240 255 1244 259
rect 1280 255 1284 259
rect 1320 255 1324 259
rect 1328 255 1332 259
rect 1368 255 1372 259
rect 1416 255 1420 259
rect 1464 255 1468 259
rect 1520 255 1524 259
rect 1560 255 1564 259
rect 152 227 156 231
rect 184 227 188 231
rect 224 227 228 231
rect 272 227 276 231
rect 320 227 324 231
rect 360 227 364 231
rect 400 227 404 231
rect 456 227 460 231
rect 528 227 532 231
rect 608 227 612 231
rect 696 227 700 231
rect 752 227 756 231
rect 784 227 788 231
rect 864 227 868 231
rect 936 227 940 231
rect 1000 227 1004 231
rect 1064 227 1068 231
rect 1120 227 1124 231
rect 1176 227 1180 231
rect 1232 227 1236 231
rect 1288 227 1292 231
rect 1344 227 1348 231
rect 1400 227 1404 231
rect 1456 227 1460 231
rect 1520 227 1524 231
rect 1560 227 1564 231
rect 1568 227 1572 231
rect 152 211 156 215
rect 184 211 188 215
rect 224 211 228 215
rect 272 211 276 215
rect 320 211 324 215
rect 360 211 364 215
rect 400 211 404 215
rect 456 211 460 215
rect 528 211 532 215
rect 608 211 612 215
rect 696 211 700 215
rect 784 211 788 215
rect 864 211 868 215
rect 936 211 940 215
rect 1000 211 1004 215
rect 1064 211 1068 215
rect 1120 211 1124 215
rect 1176 211 1180 215
rect 1232 211 1236 215
rect 1288 211 1292 215
rect 1344 211 1348 215
rect 1400 211 1404 215
rect 1456 211 1460 215
rect 1520 211 1524 215
rect 1560 211 1564 215
rect 752 203 756 207
rect 240 199 244 203
rect 152 195 156 199
rect 184 195 188 199
rect 232 195 236 199
rect 280 195 284 199
rect 328 195 332 199
rect 376 195 380 199
rect 432 195 436 199
rect 488 195 492 199
rect 552 195 556 199
rect 624 195 628 199
rect 696 195 700 199
rect 768 195 772 199
rect 832 195 836 199
rect 896 195 900 199
rect 960 195 964 199
rect 1024 195 1028 199
rect 1080 195 1084 199
rect 1136 195 1140 199
rect 1192 195 1196 199
rect 1248 195 1252 199
rect 1304 195 1308 199
rect 1360 195 1364 199
rect 1416 195 1420 199
rect 1472 195 1476 199
rect 1528 195 1532 199
rect 1560 195 1564 199
rect 1568 195 1572 199
rect 152 179 156 183
rect 184 179 188 183
rect 232 179 236 183
rect 240 179 244 183
rect 280 179 284 183
rect 328 179 332 183
rect 376 179 380 183
rect 432 179 436 183
rect 488 179 492 183
rect 552 179 556 183
rect 624 179 628 183
rect 696 179 700 183
rect 768 179 772 183
rect 832 179 836 183
rect 896 179 900 183
rect 960 179 964 183
rect 1024 179 1028 183
rect 1080 179 1084 183
rect 1136 179 1140 183
rect 1192 179 1196 183
rect 1248 179 1252 183
rect 1304 179 1308 183
rect 1360 179 1364 183
rect 1416 179 1420 183
rect 1472 179 1476 183
rect 1528 179 1532 183
rect 1560 179 1564 183
rect 160 151 164 155
rect 208 151 212 155
rect 256 151 260 155
rect 312 151 316 155
rect 368 151 372 155
rect 424 151 428 155
rect 480 151 484 155
rect 536 151 540 155
rect 592 151 596 155
rect 648 151 652 155
rect 704 151 708 155
rect 760 151 764 155
rect 816 151 820 155
rect 872 151 876 155
rect 928 151 932 155
rect 968 151 972 155
rect 992 151 996 155
rect 1056 151 1060 155
rect 1112 151 1116 155
rect 1168 151 1172 155
rect 1224 151 1228 155
rect 1272 151 1276 155
rect 1320 151 1324 155
rect 1368 151 1372 155
rect 1416 151 1420 155
rect 1472 151 1476 155
rect 1528 151 1532 155
rect 1560 151 1564 155
rect 160 135 164 139
rect 208 135 212 139
rect 256 135 260 139
rect 312 135 316 139
rect 368 135 372 139
rect 424 135 428 139
rect 480 135 484 139
rect 536 135 540 139
rect 592 135 596 139
rect 648 135 652 139
rect 704 135 708 139
rect 760 135 764 139
rect 816 135 820 139
rect 872 135 876 139
rect 928 135 932 139
rect 992 135 996 139
rect 1056 135 1060 139
rect 1112 135 1116 139
rect 1168 135 1172 139
rect 1224 135 1228 139
rect 1272 135 1276 139
rect 1320 135 1324 139
rect 1368 135 1372 139
rect 1416 135 1420 139
rect 1472 135 1476 139
rect 1528 135 1532 139
rect 1560 135 1564 139
rect 968 119 972 123
rect 152 111 156 115
rect 184 111 188 115
rect 216 111 220 115
rect 248 111 252 115
rect 280 111 284 115
rect 312 111 316 115
rect 344 111 348 115
rect 376 111 380 115
rect 408 111 412 115
rect 440 111 444 115
rect 472 111 476 115
rect 504 111 508 115
rect 536 111 540 115
rect 568 111 572 115
rect 600 111 604 115
rect 632 111 636 115
rect 664 111 668 115
rect 696 111 700 115
rect 728 111 732 115
rect 760 111 764 115
rect 792 111 796 115
rect 824 111 828 115
rect 856 111 860 115
rect 888 111 892 115
rect 920 111 924 115
rect 960 111 964 115
rect 1000 111 1004 115
rect 1048 111 1052 115
rect 1096 111 1100 115
rect 1144 111 1148 115
rect 1192 111 1196 115
rect 1240 111 1244 115
rect 1280 111 1284 115
rect 1320 111 1324 115
rect 1360 111 1364 115
rect 1400 111 1404 115
rect 1440 111 1444 115
rect 1488 111 1492 115
rect 1528 111 1532 115
rect 1560 111 1564 115
rect 152 95 156 99
rect 184 95 188 99
rect 216 95 220 99
rect 248 95 252 99
rect 280 95 284 99
rect 312 95 316 99
rect 344 95 348 99
rect 376 95 380 99
rect 408 95 412 99
rect 440 95 444 99
rect 472 95 476 99
rect 504 95 508 99
rect 536 95 540 99
rect 568 95 572 99
rect 600 95 604 99
rect 632 97 636 101
rect 664 95 668 99
rect 696 95 700 99
rect 728 95 732 99
rect 760 95 764 99
rect 792 95 796 99
rect 824 95 828 99
rect 856 95 860 99
rect 888 95 892 99
rect 920 95 924 99
rect 960 95 964 99
rect 1000 95 1004 99
rect 1048 95 1052 99
rect 1096 95 1100 99
rect 1144 95 1148 99
rect 1192 95 1196 99
rect 1240 95 1244 99
rect 1280 95 1284 99
rect 1320 95 1324 99
rect 1360 95 1364 99
rect 1400 95 1404 99
rect 1440 95 1444 99
rect 1488 95 1492 99
rect 1560 95 1564 99
<< m2 >>
rect 134 1647 140 1648
rect 110 1645 116 1646
rect 110 1641 111 1645
rect 115 1641 116 1645
rect 134 1643 135 1647
rect 139 1643 140 1647
rect 134 1642 140 1643
rect 166 1647 172 1648
rect 166 1643 167 1647
rect 171 1643 172 1647
rect 166 1642 172 1643
rect 198 1647 204 1648
rect 198 1643 199 1647
rect 203 1643 204 1647
rect 198 1642 204 1643
rect 1582 1645 1588 1646
rect 110 1640 116 1641
rect 1582 1641 1583 1645
rect 1587 1641 1588 1645
rect 1582 1640 1588 1641
rect 150 1639 157 1640
rect 150 1635 151 1639
rect 156 1635 157 1639
rect 183 1639 189 1640
rect 183 1638 184 1639
rect 150 1634 157 1635
rect 176 1636 184 1638
rect 134 1629 140 1630
rect 110 1628 116 1629
rect 110 1624 111 1628
rect 115 1624 116 1628
rect 134 1625 135 1629
rect 139 1625 140 1629
rect 134 1624 140 1625
rect 166 1629 172 1630
rect 166 1625 167 1629
rect 171 1625 172 1629
rect 166 1624 172 1625
rect 110 1623 116 1624
rect 151 1623 157 1624
rect 151 1619 152 1623
rect 156 1622 157 1623
rect 176 1622 178 1636
rect 183 1635 184 1636
rect 188 1635 189 1639
rect 183 1634 189 1635
rect 215 1639 221 1640
rect 215 1635 216 1639
rect 220 1635 221 1639
rect 215 1634 221 1635
rect 198 1629 204 1630
rect 198 1625 199 1629
rect 203 1625 204 1629
rect 198 1624 204 1625
rect 156 1620 178 1622
rect 183 1623 189 1624
rect 156 1619 157 1620
rect 151 1618 157 1619
rect 183 1619 184 1623
rect 188 1622 189 1623
rect 217 1622 219 1634
rect 1582 1628 1588 1629
rect 1582 1624 1583 1628
rect 1587 1624 1588 1628
rect 1582 1623 1588 1624
rect 188 1620 219 1622
rect 188 1619 189 1620
rect 183 1618 189 1619
rect 150 1611 157 1612
rect 110 1608 116 1609
rect 110 1604 111 1608
rect 115 1604 116 1608
rect 110 1603 116 1604
rect 134 1607 140 1608
rect 134 1603 135 1607
rect 139 1603 140 1607
rect 150 1607 151 1611
rect 156 1607 157 1611
rect 191 1611 197 1612
rect 191 1610 192 1611
rect 184 1608 192 1610
rect 150 1606 157 1607
rect 174 1607 180 1608
rect 134 1602 140 1603
rect 174 1603 175 1607
rect 179 1603 180 1607
rect 174 1602 180 1603
rect 184 1598 186 1608
rect 191 1607 192 1608
rect 196 1607 197 1611
rect 255 1611 261 1612
rect 255 1610 256 1611
rect 248 1608 256 1610
rect 191 1606 197 1607
rect 238 1607 244 1608
rect 238 1603 239 1607
rect 243 1603 244 1607
rect 238 1602 244 1603
rect 248 1598 250 1608
rect 255 1607 256 1608
rect 260 1607 261 1611
rect 311 1611 317 1612
rect 311 1610 312 1611
rect 304 1608 312 1610
rect 255 1606 261 1607
rect 294 1607 300 1608
rect 294 1603 295 1607
rect 299 1603 300 1607
rect 294 1602 300 1603
rect 304 1598 306 1608
rect 311 1607 312 1608
rect 316 1607 317 1611
rect 367 1611 373 1612
rect 311 1606 317 1607
rect 350 1607 356 1608
rect 350 1603 351 1607
rect 355 1603 356 1607
rect 367 1607 368 1611
rect 372 1610 373 1611
rect 398 1611 404 1612
rect 398 1610 399 1611
rect 372 1608 399 1610
rect 372 1607 373 1608
rect 367 1606 373 1607
rect 398 1607 399 1608
rect 403 1607 404 1611
rect 423 1611 429 1612
rect 423 1610 424 1611
rect 416 1608 424 1610
rect 398 1606 404 1607
rect 406 1607 412 1608
rect 350 1602 356 1603
rect 406 1603 407 1607
rect 411 1603 412 1607
rect 406 1602 412 1603
rect 416 1598 418 1608
rect 423 1607 424 1608
rect 428 1607 429 1611
rect 471 1611 477 1612
rect 471 1610 472 1611
rect 464 1608 472 1610
rect 423 1606 429 1607
rect 454 1607 460 1608
rect 454 1603 455 1607
rect 459 1603 460 1607
rect 454 1602 460 1603
rect 464 1598 466 1608
rect 471 1607 472 1608
rect 476 1607 477 1611
rect 519 1611 525 1612
rect 519 1610 520 1611
rect 512 1608 520 1610
rect 471 1606 477 1607
rect 502 1607 508 1608
rect 502 1603 503 1607
rect 507 1603 508 1607
rect 502 1602 508 1603
rect 512 1598 514 1608
rect 519 1607 520 1608
rect 524 1607 525 1611
rect 567 1611 573 1612
rect 567 1610 568 1611
rect 560 1608 568 1610
rect 519 1606 525 1607
rect 550 1607 556 1608
rect 550 1603 551 1607
rect 555 1603 556 1607
rect 550 1602 556 1603
rect 560 1598 562 1608
rect 567 1607 568 1608
rect 572 1607 573 1611
rect 615 1611 621 1612
rect 615 1610 616 1611
rect 608 1608 616 1610
rect 567 1606 573 1607
rect 598 1607 604 1608
rect 598 1603 599 1607
rect 603 1603 604 1607
rect 598 1602 604 1603
rect 608 1598 610 1608
rect 615 1607 616 1608
rect 620 1607 621 1611
rect 663 1611 669 1612
rect 663 1610 664 1611
rect 656 1608 664 1610
rect 615 1606 621 1607
rect 646 1607 652 1608
rect 646 1603 647 1607
rect 651 1603 652 1607
rect 646 1602 652 1603
rect 656 1598 658 1608
rect 663 1607 664 1608
rect 668 1607 669 1611
rect 711 1611 717 1612
rect 711 1610 712 1611
rect 704 1608 712 1610
rect 663 1606 669 1607
rect 694 1607 700 1608
rect 694 1603 695 1607
rect 699 1603 700 1607
rect 694 1602 700 1603
rect 704 1598 706 1608
rect 711 1607 712 1608
rect 716 1607 717 1611
rect 759 1611 765 1612
rect 759 1610 760 1611
rect 752 1608 760 1610
rect 711 1606 717 1607
rect 742 1607 748 1608
rect 742 1603 743 1607
rect 747 1603 748 1607
rect 742 1602 748 1603
rect 752 1598 754 1608
rect 759 1607 760 1608
rect 764 1607 765 1611
rect 807 1611 813 1612
rect 759 1606 765 1607
rect 790 1607 796 1608
rect 790 1603 791 1607
rect 795 1603 796 1607
rect 807 1607 808 1611
rect 812 1610 813 1611
rect 830 1611 836 1612
rect 830 1610 831 1611
rect 812 1608 831 1610
rect 812 1607 813 1608
rect 807 1606 813 1607
rect 830 1607 831 1608
rect 835 1607 836 1611
rect 855 1611 861 1612
rect 855 1610 856 1611
rect 848 1608 856 1610
rect 830 1606 836 1607
rect 838 1607 844 1608
rect 790 1602 796 1603
rect 838 1603 839 1607
rect 843 1603 844 1607
rect 838 1602 844 1603
rect 848 1598 850 1608
rect 855 1607 856 1608
rect 860 1607 861 1611
rect 903 1611 909 1612
rect 903 1610 904 1611
rect 896 1608 904 1610
rect 855 1606 861 1607
rect 886 1607 892 1608
rect 886 1603 887 1607
rect 891 1603 892 1607
rect 886 1602 892 1603
rect 896 1598 898 1608
rect 903 1607 904 1608
rect 908 1607 909 1611
rect 951 1611 957 1612
rect 951 1610 952 1611
rect 944 1608 952 1610
rect 903 1606 909 1607
rect 934 1607 940 1608
rect 934 1603 935 1607
rect 939 1603 940 1607
rect 934 1602 940 1603
rect 944 1598 946 1608
rect 951 1607 952 1608
rect 956 1607 957 1611
rect 1007 1611 1013 1612
rect 1007 1610 1008 1611
rect 1000 1608 1008 1610
rect 951 1606 957 1607
rect 990 1607 996 1608
rect 990 1603 991 1607
rect 995 1603 996 1607
rect 990 1602 996 1603
rect 1000 1598 1002 1608
rect 1007 1607 1008 1608
rect 1012 1607 1013 1611
rect 1063 1611 1069 1612
rect 1063 1610 1064 1611
rect 1056 1608 1064 1610
rect 1007 1606 1013 1607
rect 1046 1607 1052 1608
rect 1046 1603 1047 1607
rect 1051 1603 1052 1607
rect 1046 1602 1052 1603
rect 1056 1598 1058 1608
rect 1063 1607 1064 1608
rect 1068 1607 1069 1611
rect 1111 1611 1117 1612
rect 1111 1610 1112 1611
rect 1104 1608 1112 1610
rect 1063 1606 1069 1607
rect 1094 1607 1100 1608
rect 1094 1603 1095 1607
rect 1099 1603 1100 1607
rect 1094 1602 1100 1603
rect 1104 1598 1106 1608
rect 1111 1607 1112 1608
rect 1116 1607 1117 1611
rect 1159 1611 1165 1612
rect 1159 1610 1160 1611
rect 1152 1608 1160 1610
rect 1111 1606 1117 1607
rect 1142 1607 1148 1608
rect 1142 1603 1143 1607
rect 1147 1603 1148 1607
rect 1142 1602 1148 1603
rect 1152 1598 1154 1608
rect 1159 1607 1160 1608
rect 1164 1607 1165 1611
rect 1202 1611 1213 1612
rect 1159 1606 1165 1607
rect 1190 1607 1196 1608
rect 1190 1603 1191 1607
rect 1195 1603 1196 1607
rect 1202 1607 1203 1611
rect 1207 1607 1208 1611
rect 1212 1607 1213 1611
rect 1255 1611 1261 1612
rect 1255 1610 1256 1611
rect 1248 1608 1256 1610
rect 1202 1606 1213 1607
rect 1238 1607 1244 1608
rect 1190 1602 1196 1603
rect 1238 1603 1239 1607
rect 1243 1603 1244 1607
rect 1238 1602 1244 1603
rect 1248 1598 1250 1608
rect 1255 1607 1256 1608
rect 1260 1607 1261 1611
rect 1303 1611 1309 1612
rect 1303 1610 1304 1611
rect 1296 1608 1304 1610
rect 1255 1606 1261 1607
rect 1286 1607 1292 1608
rect 1286 1603 1287 1607
rect 1291 1603 1292 1607
rect 1286 1602 1292 1603
rect 1296 1598 1298 1608
rect 1303 1607 1304 1608
rect 1308 1607 1309 1611
rect 1343 1611 1349 1612
rect 1343 1610 1344 1611
rect 1336 1608 1344 1610
rect 1303 1606 1309 1607
rect 1326 1607 1332 1608
rect 1326 1603 1327 1607
rect 1331 1603 1332 1607
rect 1326 1602 1332 1603
rect 1336 1598 1338 1608
rect 1343 1607 1344 1608
rect 1348 1607 1349 1611
rect 1383 1611 1389 1612
rect 1383 1610 1384 1611
rect 1376 1608 1384 1610
rect 1343 1606 1349 1607
rect 1366 1607 1372 1608
rect 1366 1603 1367 1607
rect 1371 1603 1372 1607
rect 1366 1602 1372 1603
rect 1376 1598 1378 1608
rect 1383 1607 1384 1608
rect 1388 1607 1389 1611
rect 1423 1611 1429 1612
rect 1423 1610 1424 1611
rect 1416 1608 1424 1610
rect 1383 1606 1389 1607
rect 1406 1607 1412 1608
rect 1406 1603 1407 1607
rect 1411 1603 1412 1607
rect 1406 1602 1412 1603
rect 1416 1598 1418 1608
rect 1423 1607 1424 1608
rect 1428 1607 1429 1611
rect 1463 1611 1469 1612
rect 1463 1610 1464 1611
rect 1456 1608 1464 1610
rect 1423 1606 1429 1607
rect 1446 1607 1452 1608
rect 1446 1603 1447 1607
rect 1451 1603 1452 1607
rect 1446 1602 1452 1603
rect 1456 1598 1458 1608
rect 1463 1607 1464 1608
rect 1468 1607 1469 1611
rect 1495 1611 1501 1612
rect 1495 1610 1496 1611
rect 1488 1608 1496 1610
rect 1463 1606 1469 1607
rect 1478 1607 1484 1608
rect 1478 1603 1479 1607
rect 1483 1603 1484 1607
rect 1478 1602 1484 1603
rect 1488 1598 1490 1608
rect 1495 1607 1496 1608
rect 1500 1607 1501 1611
rect 1527 1611 1533 1612
rect 1527 1610 1528 1611
rect 1520 1608 1528 1610
rect 1495 1606 1501 1607
rect 1510 1607 1516 1608
rect 1510 1603 1511 1607
rect 1515 1603 1516 1607
rect 1510 1602 1516 1603
rect 1520 1598 1522 1608
rect 1527 1607 1528 1608
rect 1532 1607 1533 1611
rect 1559 1611 1565 1612
rect 1559 1610 1560 1611
rect 1552 1608 1560 1610
rect 1527 1606 1533 1607
rect 1542 1607 1548 1608
rect 1542 1603 1543 1607
rect 1547 1603 1548 1607
rect 1542 1602 1548 1603
rect 1552 1598 1554 1608
rect 1559 1607 1560 1608
rect 1564 1607 1565 1611
rect 1559 1606 1565 1607
rect 1582 1608 1588 1609
rect 1582 1604 1583 1608
rect 1587 1604 1588 1608
rect 1582 1603 1588 1604
rect 153 1596 186 1598
rect 224 1596 250 1598
rect 259 1596 306 1598
rect 396 1596 418 1598
rect 448 1596 466 1598
rect 496 1596 514 1598
rect 521 1596 562 1598
rect 592 1596 610 1598
rect 640 1596 658 1598
rect 689 1596 706 1598
rect 736 1596 754 1598
rect 832 1596 850 1598
rect 857 1596 898 1598
rect 928 1596 946 1598
rect 980 1596 1002 1598
rect 1036 1596 1058 1598
rect 1081 1596 1106 1598
rect 1136 1596 1154 1598
rect 1209 1596 1250 1598
rect 1280 1596 1298 1598
rect 1324 1596 1338 1598
rect 1345 1596 1378 1598
rect 1404 1596 1418 1598
rect 1444 1596 1458 1598
rect 1476 1596 1490 1598
rect 1497 1596 1522 1598
rect 1540 1596 1554 1598
rect 151 1595 157 1596
rect 110 1591 116 1592
rect 110 1587 111 1591
rect 115 1587 116 1591
rect 151 1591 152 1595
rect 156 1591 157 1595
rect 151 1590 157 1591
rect 191 1595 197 1596
rect 191 1591 192 1595
rect 196 1594 197 1595
rect 224 1594 226 1596
rect 196 1592 226 1594
rect 255 1595 261 1596
rect 196 1591 197 1592
rect 191 1590 197 1591
rect 255 1591 256 1595
rect 260 1591 261 1595
rect 255 1590 261 1591
rect 311 1595 317 1596
rect 311 1591 312 1595
rect 316 1591 317 1595
rect 311 1590 317 1591
rect 367 1595 373 1596
rect 367 1591 368 1595
rect 372 1594 373 1595
rect 396 1594 398 1596
rect 372 1592 398 1594
rect 423 1595 429 1596
rect 372 1591 373 1592
rect 367 1590 373 1591
rect 423 1591 424 1595
rect 428 1594 429 1595
rect 448 1594 450 1596
rect 428 1592 450 1594
rect 471 1595 477 1596
rect 428 1591 429 1592
rect 423 1590 429 1591
rect 471 1591 472 1595
rect 476 1594 477 1595
rect 496 1594 498 1596
rect 476 1592 498 1594
rect 519 1595 525 1596
rect 476 1591 477 1592
rect 471 1590 477 1591
rect 519 1591 520 1595
rect 524 1591 525 1595
rect 519 1590 525 1591
rect 567 1595 573 1596
rect 567 1591 568 1595
rect 572 1594 573 1595
rect 592 1594 594 1596
rect 572 1592 594 1594
rect 615 1595 621 1596
rect 572 1591 573 1592
rect 567 1590 573 1591
rect 615 1591 616 1595
rect 620 1594 621 1595
rect 640 1594 642 1596
rect 620 1592 642 1594
rect 663 1595 669 1596
rect 620 1591 621 1592
rect 615 1590 621 1591
rect 663 1591 664 1595
rect 668 1594 669 1595
rect 689 1594 691 1596
rect 668 1592 691 1594
rect 711 1595 717 1596
rect 668 1591 669 1592
rect 663 1590 669 1591
rect 711 1591 712 1595
rect 716 1594 717 1595
rect 736 1594 738 1596
rect 716 1592 738 1594
rect 759 1595 765 1596
rect 716 1591 717 1592
rect 711 1590 717 1591
rect 759 1591 760 1595
rect 764 1591 765 1595
rect 759 1590 765 1591
rect 807 1595 813 1596
rect 807 1591 808 1595
rect 812 1594 813 1595
rect 832 1594 834 1596
rect 812 1592 834 1594
rect 855 1595 861 1596
rect 812 1591 813 1592
rect 807 1590 813 1591
rect 855 1591 856 1595
rect 860 1591 861 1595
rect 855 1590 861 1591
rect 903 1595 909 1596
rect 903 1591 904 1595
rect 908 1594 909 1595
rect 928 1594 930 1596
rect 908 1592 930 1594
rect 951 1595 957 1596
rect 908 1591 909 1592
rect 903 1590 909 1591
rect 951 1591 952 1595
rect 956 1594 957 1595
rect 980 1594 982 1596
rect 956 1592 982 1594
rect 1007 1595 1013 1596
rect 956 1591 957 1592
rect 951 1590 957 1591
rect 1007 1591 1008 1595
rect 1012 1594 1013 1595
rect 1036 1594 1038 1596
rect 1012 1592 1038 1594
rect 1063 1595 1069 1596
rect 1012 1591 1013 1592
rect 1007 1590 1013 1591
rect 1063 1591 1064 1595
rect 1068 1594 1069 1595
rect 1081 1594 1083 1596
rect 1068 1592 1083 1594
rect 1111 1595 1117 1596
rect 1068 1591 1069 1592
rect 1063 1590 1069 1591
rect 1111 1591 1112 1595
rect 1116 1594 1117 1595
rect 1136 1594 1138 1596
rect 1116 1592 1138 1594
rect 1158 1595 1165 1596
rect 1116 1591 1117 1592
rect 1111 1590 1117 1591
rect 1158 1591 1159 1595
rect 1164 1591 1165 1595
rect 1158 1590 1165 1591
rect 1207 1595 1213 1596
rect 1207 1591 1208 1595
rect 1212 1591 1213 1595
rect 1207 1590 1213 1591
rect 1255 1595 1261 1596
rect 1255 1591 1256 1595
rect 1260 1594 1261 1595
rect 1280 1594 1282 1596
rect 1260 1592 1282 1594
rect 1303 1595 1309 1596
rect 1260 1591 1261 1592
rect 1255 1590 1261 1591
rect 1303 1591 1304 1595
rect 1308 1594 1309 1595
rect 1324 1594 1326 1596
rect 1308 1592 1326 1594
rect 1343 1595 1349 1596
rect 1308 1591 1309 1592
rect 1303 1590 1309 1591
rect 1343 1591 1344 1595
rect 1348 1591 1349 1595
rect 1343 1590 1349 1591
rect 1383 1595 1389 1596
rect 1383 1591 1384 1595
rect 1388 1594 1389 1595
rect 1404 1594 1406 1596
rect 1388 1592 1406 1594
rect 1423 1595 1429 1596
rect 1388 1591 1389 1592
rect 1383 1590 1389 1591
rect 1423 1591 1424 1595
rect 1428 1594 1429 1595
rect 1444 1594 1446 1596
rect 1428 1592 1446 1594
rect 1463 1595 1469 1596
rect 1428 1591 1429 1592
rect 1423 1590 1429 1591
rect 1463 1591 1464 1595
rect 1468 1594 1469 1595
rect 1476 1594 1478 1596
rect 1468 1592 1478 1594
rect 1495 1595 1501 1596
rect 1468 1591 1469 1592
rect 1463 1590 1469 1591
rect 1495 1591 1496 1595
rect 1500 1591 1501 1595
rect 1495 1590 1501 1591
rect 1527 1595 1533 1596
rect 1527 1591 1528 1595
rect 1532 1594 1533 1595
rect 1540 1594 1542 1596
rect 1532 1592 1542 1594
rect 1559 1595 1565 1596
rect 1532 1591 1533 1592
rect 1527 1590 1533 1591
rect 1559 1591 1560 1595
rect 1564 1591 1565 1595
rect 1559 1590 1565 1591
rect 1582 1591 1588 1592
rect 110 1586 116 1587
rect 134 1589 140 1590
rect 134 1585 135 1589
rect 139 1585 140 1589
rect 134 1584 140 1585
rect 174 1589 180 1590
rect 174 1585 175 1589
rect 179 1585 180 1589
rect 174 1584 180 1585
rect 238 1589 244 1590
rect 238 1585 239 1589
rect 243 1585 244 1589
rect 238 1584 244 1585
rect 294 1589 300 1590
rect 294 1585 295 1589
rect 299 1585 300 1589
rect 294 1584 300 1585
rect 194 1583 200 1584
rect 194 1579 195 1583
rect 199 1582 200 1583
rect 313 1582 315 1590
rect 350 1589 356 1590
rect 350 1585 351 1589
rect 355 1585 356 1589
rect 350 1584 356 1585
rect 406 1589 412 1590
rect 406 1585 407 1589
rect 411 1585 412 1589
rect 406 1584 412 1585
rect 454 1589 460 1590
rect 454 1585 455 1589
rect 459 1585 460 1589
rect 454 1584 460 1585
rect 502 1589 508 1590
rect 502 1585 503 1589
rect 507 1585 508 1589
rect 502 1584 508 1585
rect 550 1589 556 1590
rect 550 1585 551 1589
rect 555 1585 556 1589
rect 550 1584 556 1585
rect 598 1589 604 1590
rect 598 1585 599 1589
rect 603 1585 604 1589
rect 598 1584 604 1585
rect 646 1589 652 1590
rect 646 1585 647 1589
rect 651 1585 652 1589
rect 646 1584 652 1585
rect 694 1589 700 1590
rect 694 1585 695 1589
rect 699 1585 700 1589
rect 694 1584 700 1585
rect 742 1589 748 1590
rect 742 1585 743 1589
rect 747 1585 748 1589
rect 742 1584 748 1585
rect 199 1580 315 1582
rect 398 1583 404 1584
rect 199 1579 200 1580
rect 194 1578 200 1579
rect 398 1579 399 1583
rect 403 1582 404 1583
rect 615 1583 621 1584
rect 403 1580 546 1582
rect 403 1579 404 1580
rect 398 1578 404 1579
rect 174 1575 180 1576
rect 110 1573 116 1574
rect 110 1569 111 1573
rect 115 1569 116 1573
rect 174 1571 175 1575
rect 179 1571 180 1575
rect 174 1570 180 1571
rect 214 1575 220 1576
rect 214 1571 215 1575
rect 219 1571 220 1575
rect 214 1570 220 1571
rect 254 1575 260 1576
rect 254 1571 255 1575
rect 259 1571 260 1575
rect 254 1570 260 1571
rect 294 1575 300 1576
rect 294 1571 295 1575
rect 299 1571 300 1575
rect 294 1570 300 1571
rect 342 1575 348 1576
rect 342 1571 343 1575
rect 347 1571 348 1575
rect 342 1570 348 1571
rect 390 1575 396 1576
rect 390 1571 391 1575
rect 395 1571 396 1575
rect 390 1570 396 1571
rect 438 1575 444 1576
rect 438 1571 439 1575
rect 443 1571 444 1575
rect 438 1570 444 1571
rect 486 1575 492 1576
rect 486 1571 487 1575
rect 491 1571 492 1575
rect 486 1570 492 1571
rect 534 1575 540 1576
rect 534 1571 535 1575
rect 539 1571 540 1575
rect 534 1570 540 1571
rect 110 1568 116 1569
rect 191 1567 197 1568
rect 191 1563 192 1567
rect 196 1566 197 1567
rect 231 1567 237 1568
rect 196 1564 210 1566
rect 196 1563 197 1564
rect 191 1562 197 1563
rect 174 1557 180 1558
rect 110 1556 116 1557
rect 110 1552 111 1556
rect 115 1552 116 1556
rect 174 1553 175 1557
rect 179 1553 180 1557
rect 174 1552 180 1553
rect 110 1551 116 1552
rect 191 1551 200 1552
rect 191 1547 192 1551
rect 199 1547 200 1551
rect 208 1550 210 1564
rect 231 1563 232 1567
rect 236 1566 237 1567
rect 246 1567 252 1568
rect 246 1566 247 1567
rect 236 1564 247 1566
rect 236 1563 237 1564
rect 231 1562 237 1563
rect 246 1563 247 1564
rect 251 1563 252 1567
rect 246 1562 252 1563
rect 271 1567 277 1568
rect 271 1563 272 1567
rect 276 1566 277 1567
rect 311 1567 317 1568
rect 276 1564 291 1566
rect 276 1563 277 1564
rect 271 1562 277 1563
rect 214 1557 220 1558
rect 214 1553 215 1557
rect 219 1553 220 1557
rect 214 1552 220 1553
rect 254 1557 260 1558
rect 254 1553 255 1557
rect 259 1553 260 1557
rect 254 1552 260 1553
rect 231 1551 237 1552
rect 231 1550 232 1551
rect 208 1548 232 1550
rect 191 1546 200 1547
rect 231 1547 232 1548
rect 236 1547 237 1551
rect 231 1546 237 1547
rect 271 1551 277 1552
rect 271 1547 272 1551
rect 276 1550 277 1551
rect 279 1551 285 1552
rect 279 1550 280 1551
rect 276 1548 280 1550
rect 276 1547 277 1548
rect 271 1546 277 1547
rect 279 1547 280 1548
rect 284 1547 285 1551
rect 289 1550 291 1564
rect 311 1563 312 1567
rect 316 1566 317 1567
rect 359 1567 365 1568
rect 316 1564 354 1566
rect 316 1563 317 1564
rect 311 1562 317 1563
rect 294 1557 300 1558
rect 294 1553 295 1557
rect 299 1553 300 1557
rect 294 1552 300 1553
rect 342 1557 348 1558
rect 342 1553 343 1557
rect 347 1553 348 1557
rect 342 1552 348 1553
rect 311 1551 317 1552
rect 311 1550 312 1551
rect 289 1548 312 1550
rect 279 1546 285 1547
rect 311 1547 312 1548
rect 316 1547 317 1551
rect 352 1550 354 1564
rect 359 1563 360 1567
rect 364 1566 365 1567
rect 407 1567 413 1568
rect 364 1564 386 1566
rect 364 1563 365 1564
rect 359 1562 365 1563
rect 359 1551 365 1552
rect 359 1550 360 1551
rect 352 1548 360 1550
rect 311 1546 317 1547
rect 359 1547 360 1548
rect 364 1547 365 1551
rect 384 1550 386 1564
rect 407 1563 408 1567
rect 412 1566 413 1567
rect 455 1567 461 1568
rect 412 1564 450 1566
rect 412 1563 413 1564
rect 407 1562 413 1563
rect 390 1557 396 1558
rect 390 1553 391 1557
rect 395 1553 396 1557
rect 390 1552 396 1553
rect 438 1557 444 1558
rect 438 1553 439 1557
rect 443 1553 444 1557
rect 438 1552 444 1553
rect 407 1551 413 1552
rect 407 1550 408 1551
rect 384 1548 408 1550
rect 359 1546 365 1547
rect 407 1547 408 1548
rect 412 1547 413 1551
rect 448 1550 450 1564
rect 455 1563 456 1567
rect 460 1566 461 1567
rect 503 1567 509 1568
rect 460 1564 482 1566
rect 460 1563 461 1564
rect 455 1562 461 1563
rect 455 1551 461 1552
rect 455 1550 456 1551
rect 448 1548 456 1550
rect 407 1546 413 1547
rect 455 1547 456 1548
rect 460 1547 461 1551
rect 480 1550 482 1564
rect 503 1563 504 1567
rect 508 1566 509 1567
rect 544 1566 546 1580
rect 615 1579 616 1583
rect 620 1582 621 1583
rect 761 1582 763 1590
rect 790 1589 796 1590
rect 790 1585 791 1589
rect 795 1585 796 1589
rect 790 1584 796 1585
rect 838 1589 844 1590
rect 838 1585 839 1589
rect 843 1585 844 1589
rect 838 1584 844 1585
rect 886 1589 892 1590
rect 886 1585 887 1589
rect 891 1585 892 1589
rect 886 1584 892 1585
rect 934 1589 940 1590
rect 934 1585 935 1589
rect 939 1585 940 1589
rect 934 1584 940 1585
rect 990 1589 996 1590
rect 990 1585 991 1589
rect 995 1585 996 1589
rect 990 1584 996 1585
rect 1046 1589 1052 1590
rect 1046 1585 1047 1589
rect 1051 1585 1052 1589
rect 1046 1584 1052 1585
rect 1094 1589 1100 1590
rect 1094 1585 1095 1589
rect 1099 1585 1100 1589
rect 1094 1584 1100 1585
rect 1142 1589 1148 1590
rect 1142 1585 1143 1589
rect 1147 1585 1148 1589
rect 1142 1584 1148 1585
rect 1190 1589 1196 1590
rect 1190 1585 1191 1589
rect 1195 1585 1196 1589
rect 1190 1584 1196 1585
rect 1238 1589 1244 1590
rect 1238 1585 1239 1589
rect 1243 1585 1244 1589
rect 1238 1584 1244 1585
rect 1286 1589 1292 1590
rect 1286 1585 1287 1589
rect 1291 1585 1292 1589
rect 1286 1584 1292 1585
rect 1326 1589 1332 1590
rect 1326 1585 1327 1589
rect 1331 1585 1332 1589
rect 1326 1584 1332 1585
rect 1366 1589 1372 1590
rect 1366 1585 1367 1589
rect 1371 1585 1372 1589
rect 1366 1584 1372 1585
rect 1406 1589 1412 1590
rect 1406 1585 1407 1589
rect 1411 1585 1412 1589
rect 1406 1584 1412 1585
rect 1446 1589 1452 1590
rect 1446 1585 1447 1589
rect 1451 1585 1452 1589
rect 1446 1584 1452 1585
rect 1478 1589 1484 1590
rect 1478 1585 1479 1589
rect 1483 1585 1484 1589
rect 1478 1584 1484 1585
rect 1510 1589 1516 1590
rect 1510 1585 1511 1589
rect 1515 1585 1516 1589
rect 1510 1584 1516 1585
rect 1542 1589 1548 1590
rect 1542 1585 1543 1589
rect 1547 1585 1548 1589
rect 1542 1584 1548 1585
rect 620 1580 763 1582
rect 1498 1583 1504 1584
rect 620 1579 621 1580
rect 615 1578 621 1579
rect 1498 1579 1499 1583
rect 1503 1582 1504 1583
rect 1561 1582 1563 1590
rect 1582 1587 1583 1591
rect 1587 1587 1588 1591
rect 1582 1586 1588 1587
rect 1503 1580 1563 1582
rect 1503 1579 1504 1580
rect 1498 1578 1504 1579
rect 582 1575 588 1576
rect 582 1571 583 1575
rect 587 1571 588 1575
rect 582 1570 588 1571
rect 638 1575 644 1576
rect 638 1571 639 1575
rect 643 1571 644 1575
rect 638 1570 644 1571
rect 702 1575 708 1576
rect 702 1571 703 1575
rect 707 1571 708 1575
rect 702 1570 708 1571
rect 774 1575 780 1576
rect 774 1571 775 1575
rect 779 1571 780 1575
rect 774 1570 780 1571
rect 854 1575 860 1576
rect 854 1571 855 1575
rect 859 1571 860 1575
rect 854 1570 860 1571
rect 934 1575 940 1576
rect 934 1571 935 1575
rect 939 1571 940 1575
rect 934 1570 940 1571
rect 1014 1575 1020 1576
rect 1014 1571 1015 1575
rect 1019 1571 1020 1575
rect 1014 1570 1020 1571
rect 1086 1575 1092 1576
rect 1086 1571 1087 1575
rect 1091 1571 1092 1575
rect 1086 1570 1092 1571
rect 1158 1575 1164 1576
rect 1158 1571 1159 1575
rect 1163 1571 1164 1575
rect 1158 1570 1164 1571
rect 1238 1575 1244 1576
rect 1238 1571 1239 1575
rect 1243 1571 1244 1575
rect 1238 1570 1244 1571
rect 1318 1575 1324 1576
rect 1318 1571 1319 1575
rect 1323 1571 1324 1575
rect 1398 1575 1404 1576
rect 1318 1570 1324 1571
rect 1328 1572 1382 1574
rect 551 1567 557 1568
rect 551 1566 552 1567
rect 508 1564 530 1566
rect 544 1564 552 1566
rect 508 1563 509 1564
rect 503 1562 509 1563
rect 486 1557 492 1558
rect 486 1553 487 1557
rect 491 1553 492 1557
rect 486 1552 492 1553
rect 503 1551 509 1552
rect 503 1550 504 1551
rect 480 1548 504 1550
rect 455 1546 461 1547
rect 503 1547 504 1548
rect 508 1547 509 1551
rect 528 1550 530 1564
rect 551 1563 552 1564
rect 556 1563 557 1567
rect 551 1562 557 1563
rect 599 1567 605 1568
rect 599 1563 600 1567
rect 604 1566 605 1567
rect 655 1567 661 1568
rect 604 1564 630 1566
rect 604 1563 605 1564
rect 599 1562 605 1563
rect 534 1557 540 1558
rect 534 1553 535 1557
rect 539 1553 540 1557
rect 534 1552 540 1553
rect 582 1557 588 1558
rect 582 1553 583 1557
rect 587 1553 588 1557
rect 615 1555 621 1556
rect 615 1554 616 1555
rect 582 1552 588 1553
rect 599 1553 616 1554
rect 551 1551 557 1552
rect 551 1550 552 1551
rect 528 1548 552 1550
rect 503 1546 509 1547
rect 551 1547 552 1548
rect 556 1547 557 1551
rect 599 1549 600 1553
rect 604 1552 616 1553
rect 604 1549 605 1552
rect 615 1551 616 1552
rect 620 1551 621 1555
rect 615 1550 621 1551
rect 628 1550 630 1564
rect 655 1563 656 1567
rect 660 1566 661 1567
rect 719 1567 725 1568
rect 660 1564 690 1566
rect 660 1563 661 1564
rect 655 1562 661 1563
rect 638 1557 644 1558
rect 638 1553 639 1557
rect 643 1553 644 1557
rect 638 1552 644 1553
rect 655 1551 661 1552
rect 655 1550 656 1551
rect 599 1548 605 1549
rect 628 1548 656 1550
rect 551 1546 557 1547
rect 655 1547 656 1548
rect 660 1547 661 1551
rect 688 1550 690 1564
rect 719 1563 720 1567
rect 724 1566 725 1567
rect 766 1567 772 1568
rect 724 1564 758 1566
rect 724 1563 725 1564
rect 719 1562 725 1563
rect 702 1557 708 1558
rect 702 1553 703 1557
rect 707 1553 708 1557
rect 702 1552 708 1553
rect 719 1551 725 1552
rect 719 1550 720 1551
rect 688 1548 720 1550
rect 655 1546 661 1547
rect 719 1547 720 1548
rect 724 1547 725 1551
rect 756 1550 758 1564
rect 766 1563 767 1567
rect 771 1566 772 1567
rect 791 1567 797 1568
rect 791 1566 792 1567
rect 771 1564 792 1566
rect 771 1563 772 1564
rect 766 1562 772 1563
rect 791 1563 792 1564
rect 796 1563 797 1567
rect 791 1562 797 1563
rect 830 1567 836 1568
rect 830 1563 831 1567
rect 835 1566 836 1567
rect 871 1567 877 1568
rect 871 1566 872 1567
rect 835 1564 872 1566
rect 835 1563 836 1564
rect 830 1562 836 1563
rect 871 1563 872 1564
rect 876 1563 877 1567
rect 951 1567 957 1568
rect 951 1566 952 1567
rect 871 1562 877 1563
rect 896 1564 952 1566
rect 774 1557 780 1558
rect 774 1553 775 1557
rect 779 1553 780 1557
rect 774 1552 780 1553
rect 854 1557 860 1558
rect 854 1553 855 1557
rect 859 1553 860 1557
rect 854 1552 860 1553
rect 791 1551 797 1552
rect 791 1550 792 1551
rect 756 1548 792 1550
rect 719 1546 725 1547
rect 791 1547 792 1548
rect 796 1547 797 1551
rect 791 1546 797 1547
rect 871 1551 877 1552
rect 871 1547 872 1551
rect 876 1550 877 1551
rect 896 1550 898 1564
rect 951 1563 952 1564
rect 956 1563 957 1567
rect 951 1562 957 1563
rect 986 1567 992 1568
rect 986 1563 987 1567
rect 991 1566 992 1567
rect 1031 1567 1037 1568
rect 1031 1566 1032 1567
rect 991 1564 1032 1566
rect 991 1563 992 1564
rect 986 1562 992 1563
rect 1031 1563 1032 1564
rect 1036 1563 1037 1567
rect 1103 1567 1109 1568
rect 1103 1566 1104 1567
rect 1031 1562 1037 1563
rect 1099 1564 1104 1566
rect 934 1557 940 1558
rect 934 1553 935 1557
rect 939 1553 940 1557
rect 934 1552 940 1553
rect 1014 1557 1020 1558
rect 1014 1553 1015 1557
rect 1019 1553 1020 1557
rect 1014 1552 1020 1553
rect 1086 1557 1092 1558
rect 1086 1553 1087 1557
rect 1091 1553 1092 1557
rect 1086 1552 1092 1553
rect 876 1548 898 1550
rect 914 1551 920 1552
rect 876 1547 877 1548
rect 871 1546 877 1547
rect 914 1547 915 1551
rect 919 1550 920 1551
rect 951 1551 957 1552
rect 951 1550 952 1551
rect 919 1548 952 1550
rect 919 1547 920 1548
rect 914 1546 920 1547
rect 951 1547 952 1548
rect 956 1547 957 1551
rect 951 1546 957 1547
rect 1031 1551 1037 1552
rect 1031 1547 1032 1551
rect 1036 1550 1037 1551
rect 1099 1550 1101 1564
rect 1103 1563 1104 1564
rect 1108 1563 1109 1567
rect 1103 1562 1109 1563
rect 1175 1567 1181 1568
rect 1175 1563 1176 1567
rect 1180 1566 1181 1567
rect 1202 1567 1208 1568
rect 1202 1566 1203 1567
rect 1180 1564 1203 1566
rect 1180 1563 1181 1564
rect 1175 1562 1181 1563
rect 1202 1563 1203 1564
rect 1207 1563 1208 1567
rect 1255 1567 1261 1568
rect 1255 1566 1256 1567
rect 1202 1562 1208 1563
rect 1220 1564 1256 1566
rect 1158 1557 1164 1558
rect 1158 1553 1159 1557
rect 1163 1553 1164 1557
rect 1158 1552 1164 1553
rect 1036 1548 1101 1550
rect 1103 1551 1109 1552
rect 1036 1547 1037 1548
rect 1031 1546 1037 1547
rect 1103 1547 1104 1551
rect 1108 1550 1109 1551
rect 1150 1551 1156 1552
rect 1150 1550 1151 1551
rect 1108 1548 1151 1550
rect 1108 1547 1109 1548
rect 1103 1546 1109 1547
rect 1150 1547 1151 1548
rect 1155 1547 1156 1551
rect 1150 1546 1156 1547
rect 1175 1551 1181 1552
rect 1175 1547 1176 1551
rect 1180 1550 1181 1551
rect 1220 1550 1222 1564
rect 1255 1563 1256 1564
rect 1260 1563 1261 1567
rect 1328 1566 1330 1572
rect 1255 1562 1261 1563
rect 1312 1564 1330 1566
rect 1335 1567 1341 1568
rect 1238 1557 1244 1558
rect 1238 1553 1239 1557
rect 1243 1553 1244 1557
rect 1238 1552 1244 1553
rect 1180 1548 1222 1550
rect 1255 1551 1261 1552
rect 1180 1547 1181 1548
rect 1175 1546 1181 1547
rect 1255 1547 1256 1551
rect 1260 1550 1261 1551
rect 1312 1550 1314 1564
rect 1335 1563 1336 1567
rect 1340 1566 1341 1567
rect 1380 1566 1382 1572
rect 1398 1571 1399 1575
rect 1403 1571 1404 1575
rect 1398 1570 1404 1571
rect 1478 1575 1484 1576
rect 1478 1571 1479 1575
rect 1483 1571 1484 1575
rect 1478 1570 1484 1571
rect 1542 1575 1548 1576
rect 1542 1571 1543 1575
rect 1547 1571 1548 1575
rect 1542 1570 1548 1571
rect 1582 1573 1588 1574
rect 1582 1569 1583 1573
rect 1587 1569 1588 1573
rect 1582 1568 1588 1569
rect 1415 1567 1421 1568
rect 1415 1566 1416 1567
rect 1340 1564 1378 1566
rect 1380 1564 1416 1566
rect 1340 1563 1341 1564
rect 1335 1562 1341 1563
rect 1318 1557 1324 1558
rect 1318 1553 1319 1557
rect 1323 1553 1324 1557
rect 1318 1552 1324 1553
rect 1260 1548 1314 1550
rect 1326 1551 1332 1552
rect 1260 1547 1261 1548
rect 1255 1546 1261 1547
rect 1326 1547 1327 1551
rect 1331 1550 1332 1551
rect 1335 1551 1341 1552
rect 1335 1550 1336 1551
rect 1331 1548 1336 1550
rect 1331 1547 1332 1548
rect 1326 1546 1332 1547
rect 1335 1547 1336 1548
rect 1340 1547 1341 1551
rect 1376 1550 1378 1564
rect 1415 1563 1416 1564
rect 1420 1563 1421 1567
rect 1415 1562 1421 1563
rect 1495 1567 1501 1568
rect 1495 1563 1496 1567
rect 1500 1566 1501 1567
rect 1558 1567 1565 1568
rect 1500 1564 1554 1566
rect 1500 1563 1501 1564
rect 1495 1562 1501 1563
rect 1398 1557 1404 1558
rect 1398 1553 1399 1557
rect 1403 1553 1404 1557
rect 1398 1552 1404 1553
rect 1478 1557 1484 1558
rect 1478 1553 1479 1557
rect 1483 1553 1484 1557
rect 1542 1557 1548 1558
rect 1498 1555 1504 1556
rect 1498 1554 1499 1555
rect 1478 1552 1484 1553
rect 1495 1553 1499 1554
rect 1415 1551 1421 1552
rect 1415 1550 1416 1551
rect 1376 1548 1416 1550
rect 1335 1546 1341 1547
rect 1415 1547 1416 1548
rect 1420 1547 1421 1551
rect 1495 1549 1496 1553
rect 1503 1551 1504 1555
rect 1542 1553 1543 1557
rect 1547 1553 1548 1557
rect 1542 1552 1548 1553
rect 1500 1550 1504 1551
rect 1552 1550 1554 1564
rect 1558 1563 1559 1567
rect 1564 1563 1565 1567
rect 1558 1562 1565 1563
rect 1582 1556 1588 1557
rect 1582 1552 1583 1556
rect 1587 1552 1588 1556
rect 1559 1551 1565 1552
rect 1582 1551 1588 1552
rect 1559 1550 1560 1551
rect 1500 1549 1501 1550
rect 1495 1548 1501 1549
rect 1552 1548 1560 1550
rect 1415 1546 1421 1547
rect 1559 1547 1560 1548
rect 1564 1547 1565 1551
rect 1559 1546 1565 1547
rect 246 1543 252 1544
rect 175 1539 181 1540
rect 110 1536 116 1537
rect 110 1532 111 1536
rect 115 1532 116 1536
rect 110 1531 116 1532
rect 158 1535 164 1536
rect 158 1531 159 1535
rect 163 1531 164 1535
rect 175 1535 176 1539
rect 180 1538 181 1539
rect 223 1539 229 1540
rect 180 1536 202 1538
rect 180 1535 181 1536
rect 175 1534 181 1535
rect 158 1530 164 1531
rect 200 1526 202 1536
rect 206 1535 212 1536
rect 206 1531 207 1535
rect 211 1531 212 1535
rect 223 1535 224 1539
rect 228 1538 229 1539
rect 246 1539 247 1543
rect 251 1542 252 1543
rect 766 1543 772 1544
rect 766 1542 767 1543
rect 251 1541 277 1542
rect 251 1540 272 1541
rect 251 1539 252 1540
rect 246 1538 252 1539
rect 228 1536 242 1538
rect 271 1537 272 1540
rect 276 1537 277 1541
rect 752 1540 767 1542
rect 271 1536 277 1537
rect 327 1539 333 1540
rect 228 1535 229 1536
rect 223 1534 229 1535
rect 206 1530 212 1531
rect 240 1526 242 1536
rect 254 1535 260 1536
rect 254 1531 255 1535
rect 259 1531 260 1535
rect 254 1530 260 1531
rect 310 1535 316 1536
rect 310 1531 311 1535
rect 315 1531 316 1535
rect 327 1535 328 1539
rect 332 1538 333 1539
rect 343 1539 349 1540
rect 343 1538 344 1539
rect 332 1536 344 1538
rect 332 1535 333 1536
rect 327 1534 333 1535
rect 343 1535 344 1536
rect 348 1535 349 1539
rect 370 1539 381 1540
rect 343 1534 349 1535
rect 358 1535 364 1536
rect 310 1530 316 1531
rect 358 1531 359 1535
rect 363 1531 364 1535
rect 370 1535 371 1539
rect 375 1535 376 1539
rect 380 1535 381 1539
rect 431 1539 437 1540
rect 431 1538 432 1539
rect 424 1536 432 1538
rect 370 1534 381 1535
rect 414 1535 420 1536
rect 358 1530 364 1531
rect 414 1531 415 1535
rect 419 1531 420 1535
rect 414 1530 420 1531
rect 264 1528 274 1530
rect 264 1526 266 1528
rect 272 1526 274 1528
rect 279 1527 285 1528
rect 200 1524 218 1526
rect 240 1524 266 1526
rect 271 1525 277 1526
rect 174 1523 181 1524
rect 110 1519 116 1520
rect 110 1515 111 1519
rect 115 1515 116 1519
rect 174 1519 175 1523
rect 180 1519 181 1523
rect 216 1522 218 1524
rect 223 1523 229 1524
rect 223 1522 224 1523
rect 216 1520 224 1522
rect 174 1518 181 1519
rect 223 1519 224 1520
rect 228 1519 229 1523
rect 271 1521 272 1525
rect 276 1521 277 1525
rect 279 1523 280 1527
rect 284 1526 285 1527
rect 424 1526 426 1536
rect 431 1535 432 1536
rect 436 1535 437 1539
rect 487 1539 493 1540
rect 431 1534 437 1535
rect 470 1535 476 1536
rect 470 1531 471 1535
rect 475 1531 476 1535
rect 487 1535 488 1539
rect 492 1538 493 1539
rect 543 1539 549 1540
rect 492 1536 522 1538
rect 492 1535 493 1536
rect 487 1534 493 1535
rect 470 1530 476 1531
rect 284 1524 322 1526
rect 377 1524 426 1526
rect 439 1527 445 1528
rect 284 1523 285 1524
rect 279 1522 285 1523
rect 320 1522 322 1524
rect 327 1523 333 1524
rect 327 1522 328 1523
rect 271 1520 277 1521
rect 320 1520 328 1522
rect 223 1518 229 1519
rect 327 1519 328 1520
rect 332 1519 333 1523
rect 327 1518 333 1519
rect 375 1523 381 1524
rect 375 1519 376 1523
rect 380 1519 381 1523
rect 431 1523 437 1524
rect 431 1522 432 1523
rect 375 1518 381 1519
rect 424 1520 432 1522
rect 110 1514 116 1515
rect 158 1517 164 1518
rect 158 1513 159 1517
rect 163 1513 164 1517
rect 158 1512 164 1513
rect 206 1517 212 1518
rect 206 1513 207 1517
rect 211 1513 212 1517
rect 206 1512 212 1513
rect 254 1517 260 1518
rect 254 1513 255 1517
rect 259 1513 260 1517
rect 254 1512 260 1513
rect 310 1517 316 1518
rect 310 1513 311 1517
rect 315 1513 316 1517
rect 310 1512 316 1513
rect 358 1517 364 1518
rect 358 1513 359 1517
rect 363 1513 364 1517
rect 358 1512 364 1513
rect 414 1517 420 1518
rect 414 1513 415 1517
rect 419 1513 420 1517
rect 414 1512 420 1513
rect 343 1511 349 1512
rect 343 1507 344 1511
rect 348 1510 349 1511
rect 424 1510 426 1520
rect 431 1519 432 1520
rect 436 1519 437 1523
rect 439 1523 440 1527
rect 444 1526 445 1527
rect 520 1526 522 1536
rect 526 1535 532 1536
rect 526 1531 527 1535
rect 531 1531 532 1535
rect 543 1535 544 1539
rect 548 1538 549 1539
rect 599 1539 605 1540
rect 548 1536 578 1538
rect 548 1535 549 1536
rect 543 1534 549 1535
rect 526 1530 532 1531
rect 576 1526 578 1536
rect 582 1535 588 1536
rect 582 1531 583 1535
rect 587 1531 588 1535
rect 599 1535 600 1539
rect 604 1538 605 1539
rect 655 1539 661 1540
rect 604 1536 634 1538
rect 604 1535 605 1536
rect 599 1534 605 1535
rect 582 1530 588 1531
rect 632 1526 634 1536
rect 638 1535 644 1536
rect 638 1531 639 1535
rect 643 1531 644 1535
rect 655 1535 656 1539
rect 660 1538 661 1539
rect 711 1539 717 1540
rect 660 1536 690 1538
rect 660 1535 661 1536
rect 655 1534 661 1535
rect 638 1530 644 1531
rect 688 1526 690 1536
rect 694 1535 700 1536
rect 694 1531 695 1535
rect 699 1531 700 1535
rect 711 1535 712 1539
rect 716 1538 717 1539
rect 752 1538 754 1540
rect 766 1539 767 1540
rect 771 1539 772 1543
rect 1063 1543 1069 1544
rect 766 1538 772 1539
rect 775 1539 781 1540
rect 716 1536 754 1538
rect 775 1536 776 1539
rect 716 1535 717 1536
rect 711 1534 717 1535
rect 758 1535 764 1536
rect 694 1530 700 1531
rect 758 1531 759 1535
rect 763 1531 764 1535
rect 758 1530 764 1531
rect 774 1535 776 1536
rect 780 1535 781 1539
rect 839 1539 845 1540
rect 839 1538 840 1539
rect 832 1536 840 1538
rect 774 1531 775 1535
rect 779 1534 781 1535
rect 822 1535 828 1536
rect 779 1531 780 1534
rect 774 1530 780 1531
rect 822 1531 823 1535
rect 827 1531 828 1535
rect 822 1530 828 1531
rect 832 1526 834 1536
rect 839 1535 840 1536
rect 844 1535 845 1539
rect 911 1539 917 1540
rect 911 1538 912 1539
rect 904 1536 912 1538
rect 839 1534 845 1535
rect 894 1535 900 1536
rect 894 1531 895 1535
rect 899 1531 900 1535
rect 894 1530 900 1531
rect 904 1526 906 1536
rect 911 1535 912 1536
rect 916 1535 917 1539
rect 983 1539 992 1540
rect 911 1534 917 1535
rect 966 1535 972 1536
rect 966 1531 967 1535
rect 971 1531 972 1535
rect 983 1535 984 1539
rect 991 1535 992 1539
rect 1055 1539 1061 1540
rect 1055 1538 1056 1539
rect 1048 1536 1056 1538
rect 983 1534 992 1535
rect 1038 1535 1044 1536
rect 966 1530 972 1531
rect 1038 1531 1039 1535
rect 1043 1531 1044 1535
rect 1038 1530 1044 1531
rect 1048 1526 1050 1536
rect 1055 1535 1056 1536
rect 1060 1535 1061 1539
rect 1063 1539 1064 1543
rect 1068 1542 1069 1543
rect 1068 1540 1114 1542
rect 1068 1539 1069 1540
rect 1063 1538 1069 1539
rect 1112 1538 1114 1540
rect 1119 1539 1125 1540
rect 1119 1538 1120 1539
rect 1112 1536 1120 1538
rect 1055 1534 1061 1535
rect 1102 1535 1108 1536
rect 1102 1531 1103 1535
rect 1107 1531 1108 1535
rect 1119 1535 1120 1536
rect 1124 1535 1125 1539
rect 1183 1539 1189 1540
rect 1119 1534 1125 1535
rect 1166 1535 1172 1536
rect 1102 1530 1108 1531
rect 1166 1531 1167 1535
rect 1171 1531 1172 1535
rect 1183 1535 1184 1539
rect 1188 1538 1189 1539
rect 1222 1539 1228 1540
rect 1222 1538 1223 1539
rect 1188 1536 1223 1538
rect 1188 1535 1189 1536
rect 1183 1534 1189 1535
rect 1222 1535 1223 1536
rect 1227 1535 1228 1539
rect 1247 1539 1253 1540
rect 1247 1538 1248 1539
rect 1240 1536 1248 1538
rect 1222 1534 1228 1535
rect 1230 1535 1236 1536
rect 1166 1530 1172 1531
rect 1230 1531 1231 1535
rect 1235 1531 1236 1535
rect 1230 1530 1236 1531
rect 1240 1526 1242 1536
rect 1247 1535 1248 1536
rect 1252 1535 1253 1539
rect 1311 1539 1317 1540
rect 1311 1538 1312 1539
rect 1304 1536 1312 1538
rect 1247 1534 1253 1535
rect 1294 1535 1300 1536
rect 1294 1531 1295 1535
rect 1299 1531 1300 1535
rect 1294 1530 1300 1531
rect 1304 1526 1306 1536
rect 1311 1535 1312 1536
rect 1316 1535 1317 1539
rect 1375 1539 1381 1540
rect 1311 1534 1317 1535
rect 1358 1535 1364 1536
rect 1358 1531 1359 1535
rect 1363 1531 1364 1535
rect 1375 1535 1376 1539
rect 1380 1538 1381 1539
rect 1438 1539 1445 1540
rect 1380 1536 1418 1538
rect 1380 1535 1381 1536
rect 1375 1534 1381 1535
rect 1358 1530 1364 1531
rect 444 1524 482 1526
rect 520 1524 538 1526
rect 576 1524 594 1526
rect 632 1524 650 1526
rect 688 1524 706 1526
rect 808 1524 834 1526
rect 876 1524 906 1526
rect 1020 1524 1050 1526
rect 1216 1524 1242 1526
rect 1280 1524 1306 1526
rect 1416 1526 1418 1536
rect 1422 1535 1428 1536
rect 1422 1531 1423 1535
rect 1427 1531 1428 1535
rect 1438 1535 1439 1539
rect 1444 1535 1445 1539
rect 1511 1539 1517 1540
rect 1438 1534 1445 1535
rect 1494 1535 1500 1536
rect 1422 1530 1428 1531
rect 1494 1531 1495 1535
rect 1499 1531 1500 1535
rect 1511 1535 1512 1539
rect 1516 1538 1517 1539
rect 1558 1539 1565 1540
rect 1516 1536 1538 1538
rect 1516 1535 1517 1536
rect 1511 1534 1517 1535
rect 1494 1530 1500 1531
rect 1536 1526 1538 1536
rect 1542 1535 1548 1536
rect 1542 1531 1543 1535
rect 1547 1531 1548 1535
rect 1558 1535 1559 1539
rect 1564 1535 1565 1539
rect 1558 1534 1565 1535
rect 1582 1536 1588 1537
rect 1582 1532 1583 1536
rect 1587 1532 1588 1536
rect 1582 1531 1588 1532
rect 1542 1530 1548 1531
rect 1416 1524 1434 1526
rect 1536 1524 1563 1526
rect 444 1523 445 1524
rect 439 1522 445 1523
rect 480 1522 482 1524
rect 487 1523 493 1524
rect 487 1522 488 1523
rect 480 1520 488 1522
rect 431 1518 437 1519
rect 487 1519 488 1520
rect 492 1519 493 1523
rect 536 1522 538 1524
rect 543 1523 549 1524
rect 543 1522 544 1523
rect 536 1520 544 1522
rect 487 1518 493 1519
rect 543 1519 544 1520
rect 548 1519 549 1523
rect 592 1522 594 1524
rect 599 1523 605 1524
rect 599 1522 600 1523
rect 592 1520 600 1522
rect 543 1518 549 1519
rect 599 1519 600 1520
rect 604 1519 605 1523
rect 648 1522 650 1524
rect 655 1523 661 1524
rect 655 1522 656 1523
rect 648 1520 656 1522
rect 599 1518 605 1519
rect 655 1519 656 1520
rect 660 1519 661 1523
rect 704 1522 706 1524
rect 711 1523 717 1524
rect 711 1522 712 1523
rect 704 1520 712 1522
rect 655 1518 661 1519
rect 711 1519 712 1520
rect 716 1519 717 1523
rect 711 1518 717 1519
rect 775 1523 781 1524
rect 775 1519 776 1523
rect 780 1522 781 1523
rect 808 1522 810 1524
rect 780 1520 810 1522
rect 839 1523 845 1524
rect 780 1519 781 1520
rect 775 1518 781 1519
rect 839 1519 840 1523
rect 844 1522 845 1523
rect 876 1522 878 1524
rect 844 1520 878 1522
rect 911 1523 920 1524
rect 844 1519 845 1520
rect 839 1518 845 1519
rect 911 1519 912 1523
rect 919 1519 920 1523
rect 911 1518 920 1519
rect 983 1523 989 1524
rect 983 1519 984 1523
rect 988 1522 989 1523
rect 1020 1522 1022 1524
rect 988 1520 1022 1522
rect 1055 1523 1061 1524
rect 988 1519 989 1520
rect 983 1518 989 1519
rect 1055 1519 1056 1523
rect 1060 1522 1061 1523
rect 1063 1523 1069 1524
rect 1063 1522 1064 1523
rect 1060 1520 1064 1522
rect 1060 1519 1061 1520
rect 1055 1518 1061 1519
rect 1063 1519 1064 1520
rect 1068 1519 1069 1523
rect 1063 1518 1069 1519
rect 1114 1523 1125 1524
rect 1114 1519 1115 1523
rect 1119 1519 1120 1523
rect 1124 1519 1125 1523
rect 1114 1518 1125 1519
rect 1183 1523 1189 1524
rect 1183 1519 1184 1523
rect 1188 1522 1189 1523
rect 1216 1522 1218 1524
rect 1188 1520 1218 1522
rect 1247 1523 1253 1524
rect 1188 1519 1189 1520
rect 1183 1518 1189 1519
rect 1247 1519 1248 1523
rect 1252 1522 1253 1523
rect 1280 1522 1282 1524
rect 1252 1520 1282 1522
rect 1311 1523 1317 1524
rect 1252 1519 1253 1520
rect 1247 1518 1253 1519
rect 1311 1519 1312 1523
rect 1316 1522 1317 1523
rect 1326 1523 1332 1524
rect 1326 1522 1327 1523
rect 1316 1520 1327 1522
rect 1316 1519 1317 1520
rect 1311 1518 1317 1519
rect 1326 1519 1327 1520
rect 1331 1519 1332 1523
rect 1375 1523 1381 1524
rect 1375 1522 1376 1523
rect 1326 1518 1332 1519
rect 1368 1520 1376 1522
rect 470 1517 476 1518
rect 470 1513 471 1517
rect 475 1513 476 1517
rect 470 1512 476 1513
rect 526 1517 532 1518
rect 526 1513 527 1517
rect 531 1513 532 1517
rect 526 1512 532 1513
rect 582 1517 588 1518
rect 582 1513 583 1517
rect 587 1513 588 1517
rect 582 1512 588 1513
rect 638 1517 644 1518
rect 638 1513 639 1517
rect 643 1513 644 1517
rect 638 1512 644 1513
rect 694 1517 700 1518
rect 694 1513 695 1517
rect 699 1513 700 1517
rect 694 1512 700 1513
rect 758 1517 764 1518
rect 758 1513 759 1517
rect 763 1513 764 1517
rect 758 1512 764 1513
rect 822 1517 828 1518
rect 822 1513 823 1517
rect 827 1513 828 1517
rect 822 1512 828 1513
rect 894 1517 900 1518
rect 894 1513 895 1517
rect 899 1513 900 1517
rect 894 1512 900 1513
rect 966 1517 972 1518
rect 966 1513 967 1517
rect 971 1513 972 1517
rect 966 1512 972 1513
rect 1038 1517 1044 1518
rect 1038 1513 1039 1517
rect 1043 1513 1044 1517
rect 1038 1512 1044 1513
rect 1102 1517 1108 1518
rect 1102 1513 1103 1517
rect 1107 1513 1108 1517
rect 1102 1512 1108 1513
rect 1166 1517 1172 1518
rect 1166 1513 1167 1517
rect 1171 1513 1172 1517
rect 1166 1512 1172 1513
rect 1230 1517 1236 1518
rect 1230 1513 1231 1517
rect 1235 1513 1236 1517
rect 1230 1512 1236 1513
rect 1294 1517 1300 1518
rect 1294 1513 1295 1517
rect 1299 1513 1300 1517
rect 1294 1512 1300 1513
rect 1358 1517 1364 1518
rect 1358 1513 1359 1517
rect 1363 1513 1364 1517
rect 1358 1512 1364 1513
rect 348 1508 426 1510
rect 482 1511 488 1512
rect 348 1507 349 1508
rect 343 1506 349 1507
rect 482 1507 483 1511
rect 487 1510 488 1511
rect 1222 1511 1228 1512
rect 487 1508 646 1510
rect 487 1507 488 1508
rect 482 1506 488 1507
rect 158 1503 164 1504
rect 110 1501 116 1502
rect 110 1497 111 1501
rect 115 1497 116 1501
rect 158 1499 159 1503
rect 163 1499 164 1503
rect 158 1498 164 1499
rect 206 1503 212 1504
rect 206 1499 207 1503
rect 211 1499 212 1503
rect 206 1498 212 1499
rect 254 1503 260 1504
rect 254 1499 255 1503
rect 259 1499 260 1503
rect 254 1498 260 1499
rect 302 1503 308 1504
rect 302 1499 303 1503
rect 307 1499 308 1503
rect 302 1498 308 1499
rect 350 1503 356 1504
rect 350 1499 351 1503
rect 355 1499 356 1503
rect 350 1498 356 1499
rect 406 1503 412 1504
rect 406 1499 407 1503
rect 411 1499 412 1503
rect 406 1498 412 1499
rect 462 1503 468 1504
rect 462 1499 463 1503
rect 467 1499 468 1503
rect 462 1498 468 1499
rect 526 1503 532 1504
rect 526 1499 527 1503
rect 531 1499 532 1503
rect 526 1498 532 1499
rect 590 1503 596 1504
rect 590 1499 591 1503
rect 595 1499 596 1503
rect 590 1498 596 1499
rect 110 1496 116 1497
rect 175 1495 181 1496
rect 175 1491 176 1495
rect 180 1494 181 1495
rect 218 1495 229 1496
rect 180 1492 202 1494
rect 180 1491 181 1492
rect 175 1490 181 1491
rect 158 1485 164 1486
rect 110 1484 116 1485
rect 110 1480 111 1484
rect 115 1480 116 1484
rect 158 1481 159 1485
rect 163 1481 164 1485
rect 158 1480 164 1481
rect 110 1479 116 1480
rect 174 1479 181 1480
rect 174 1475 175 1479
rect 180 1475 181 1479
rect 200 1478 202 1492
rect 218 1491 219 1495
rect 223 1491 224 1495
rect 228 1491 229 1495
rect 218 1490 229 1491
rect 271 1495 277 1496
rect 271 1491 272 1495
rect 276 1494 277 1495
rect 319 1495 325 1496
rect 276 1492 298 1494
rect 276 1491 277 1492
rect 271 1490 277 1491
rect 206 1485 212 1486
rect 206 1481 207 1485
rect 211 1481 212 1485
rect 206 1480 212 1481
rect 254 1485 260 1486
rect 254 1481 255 1485
rect 259 1481 260 1485
rect 254 1480 260 1481
rect 223 1479 229 1480
rect 223 1478 224 1479
rect 200 1476 224 1478
rect 174 1474 181 1475
rect 223 1475 224 1476
rect 228 1475 229 1479
rect 223 1474 229 1475
rect 271 1479 280 1480
rect 271 1475 272 1479
rect 279 1475 280 1479
rect 296 1478 298 1492
rect 319 1491 320 1495
rect 324 1494 325 1495
rect 367 1495 376 1496
rect 324 1492 346 1494
rect 324 1491 325 1492
rect 319 1490 325 1491
rect 302 1485 308 1486
rect 302 1481 303 1485
rect 307 1481 308 1485
rect 302 1480 308 1481
rect 319 1479 325 1480
rect 319 1478 320 1479
rect 296 1476 320 1478
rect 271 1474 280 1475
rect 319 1475 320 1476
rect 324 1475 325 1479
rect 344 1478 346 1492
rect 367 1491 368 1495
rect 375 1491 376 1495
rect 367 1490 376 1491
rect 423 1495 429 1496
rect 423 1491 424 1495
rect 428 1494 429 1495
rect 479 1495 485 1496
rect 428 1492 454 1494
rect 428 1491 429 1492
rect 423 1490 429 1491
rect 350 1485 356 1486
rect 350 1481 351 1485
rect 355 1481 356 1485
rect 350 1480 356 1481
rect 406 1485 412 1486
rect 406 1481 407 1485
rect 411 1481 412 1485
rect 406 1480 412 1481
rect 367 1479 373 1480
rect 367 1478 368 1479
rect 344 1476 368 1478
rect 319 1474 325 1475
rect 367 1475 368 1476
rect 372 1475 373 1479
rect 367 1474 373 1475
rect 423 1479 429 1480
rect 423 1475 424 1479
rect 428 1478 429 1479
rect 439 1479 445 1480
rect 439 1478 440 1479
rect 428 1476 440 1478
rect 428 1475 429 1476
rect 423 1474 429 1475
rect 439 1475 440 1476
rect 444 1475 445 1479
rect 452 1478 454 1492
rect 479 1491 480 1495
rect 484 1494 485 1495
rect 543 1495 549 1496
rect 484 1492 514 1494
rect 484 1491 485 1492
rect 479 1490 485 1491
rect 462 1485 468 1486
rect 462 1481 463 1485
rect 467 1481 468 1485
rect 462 1480 468 1481
rect 479 1479 485 1480
rect 479 1478 480 1479
rect 452 1476 480 1478
rect 439 1474 445 1475
rect 479 1475 480 1476
rect 484 1475 485 1479
rect 512 1478 514 1492
rect 543 1491 544 1495
rect 548 1494 549 1495
rect 607 1495 613 1496
rect 548 1492 578 1494
rect 548 1491 549 1492
rect 543 1490 549 1491
rect 526 1485 532 1486
rect 526 1481 527 1485
rect 531 1481 532 1485
rect 526 1480 532 1481
rect 543 1479 549 1480
rect 543 1478 544 1479
rect 512 1476 544 1478
rect 479 1474 485 1475
rect 543 1475 544 1476
rect 548 1475 549 1479
rect 576 1478 578 1492
rect 607 1491 608 1495
rect 612 1494 613 1495
rect 644 1494 646 1508
rect 1222 1507 1223 1511
rect 1227 1510 1228 1511
rect 1368 1510 1370 1520
rect 1375 1519 1376 1520
rect 1380 1519 1381 1523
rect 1432 1522 1434 1524
rect 1439 1523 1445 1524
rect 1439 1522 1440 1523
rect 1432 1520 1440 1522
rect 1375 1518 1381 1519
rect 1439 1519 1440 1520
rect 1444 1519 1445 1523
rect 1439 1518 1445 1519
rect 1510 1523 1517 1524
rect 1510 1519 1511 1523
rect 1516 1519 1517 1523
rect 1510 1518 1517 1519
rect 1559 1523 1565 1524
rect 1559 1519 1560 1523
rect 1564 1519 1565 1523
rect 1559 1518 1565 1519
rect 1582 1519 1588 1520
rect 1422 1517 1428 1518
rect 1422 1513 1423 1517
rect 1427 1513 1428 1517
rect 1422 1512 1428 1513
rect 1494 1517 1500 1518
rect 1494 1513 1495 1517
rect 1499 1513 1500 1517
rect 1494 1512 1500 1513
rect 1542 1517 1548 1518
rect 1542 1513 1543 1517
rect 1547 1513 1548 1517
rect 1582 1515 1583 1519
rect 1587 1515 1588 1519
rect 1582 1514 1588 1515
rect 1542 1512 1548 1513
rect 1227 1508 1370 1510
rect 1227 1507 1228 1508
rect 1222 1506 1228 1507
rect 654 1503 660 1504
rect 654 1499 655 1503
rect 659 1499 660 1503
rect 654 1498 660 1499
rect 718 1503 724 1504
rect 718 1499 719 1503
rect 723 1499 724 1503
rect 718 1498 724 1499
rect 782 1503 788 1504
rect 782 1499 783 1503
rect 787 1499 788 1503
rect 782 1498 788 1499
rect 854 1503 860 1504
rect 854 1499 855 1503
rect 859 1499 860 1503
rect 854 1498 860 1499
rect 934 1503 940 1504
rect 934 1499 935 1503
rect 939 1499 940 1503
rect 934 1498 940 1499
rect 1006 1503 1012 1504
rect 1006 1499 1007 1503
rect 1011 1499 1012 1503
rect 1006 1498 1012 1499
rect 1078 1503 1084 1504
rect 1078 1499 1079 1503
rect 1083 1499 1084 1503
rect 1078 1498 1084 1499
rect 1150 1503 1156 1504
rect 1150 1499 1151 1503
rect 1155 1499 1156 1503
rect 1150 1498 1156 1499
rect 1214 1503 1220 1504
rect 1214 1499 1215 1503
rect 1219 1499 1220 1503
rect 1214 1498 1220 1499
rect 1278 1503 1284 1504
rect 1278 1499 1279 1503
rect 1283 1499 1284 1503
rect 1278 1498 1284 1499
rect 1350 1503 1356 1504
rect 1350 1499 1351 1503
rect 1355 1499 1356 1503
rect 1350 1498 1356 1499
rect 1422 1503 1428 1504
rect 1422 1499 1423 1503
rect 1427 1499 1428 1503
rect 1422 1498 1428 1499
rect 1494 1503 1500 1504
rect 1494 1499 1495 1503
rect 1499 1499 1500 1503
rect 1494 1498 1500 1499
rect 1542 1503 1548 1504
rect 1542 1499 1543 1503
rect 1547 1499 1548 1503
rect 1542 1498 1548 1499
rect 1582 1501 1588 1502
rect 1582 1497 1583 1501
rect 1587 1497 1588 1501
rect 1582 1496 1588 1497
rect 671 1495 677 1496
rect 671 1494 672 1495
rect 612 1492 642 1494
rect 644 1492 672 1494
rect 612 1491 613 1492
rect 607 1490 613 1491
rect 590 1485 596 1486
rect 590 1481 591 1485
rect 595 1481 596 1485
rect 590 1480 596 1481
rect 607 1479 613 1480
rect 607 1478 608 1479
rect 576 1476 608 1478
rect 543 1474 549 1475
rect 607 1475 608 1476
rect 612 1475 613 1479
rect 640 1478 642 1492
rect 671 1491 672 1492
rect 676 1491 677 1495
rect 671 1490 677 1491
rect 735 1495 741 1496
rect 735 1491 736 1495
rect 740 1494 741 1495
rect 774 1495 780 1496
rect 774 1494 775 1495
rect 740 1492 775 1494
rect 740 1491 741 1492
rect 735 1490 741 1491
rect 774 1491 775 1492
rect 779 1491 780 1495
rect 799 1495 805 1496
rect 799 1494 800 1495
rect 774 1490 780 1491
rect 792 1492 800 1494
rect 654 1485 660 1486
rect 654 1481 655 1485
rect 659 1481 660 1485
rect 654 1480 660 1481
rect 718 1485 724 1486
rect 718 1481 719 1485
rect 723 1481 724 1485
rect 718 1480 724 1481
rect 782 1485 788 1486
rect 782 1481 783 1485
rect 787 1481 788 1485
rect 782 1480 788 1481
rect 671 1479 677 1480
rect 671 1478 672 1479
rect 640 1476 672 1478
rect 607 1474 613 1475
rect 671 1475 672 1476
rect 676 1475 677 1479
rect 671 1474 677 1475
rect 735 1479 741 1480
rect 735 1475 736 1479
rect 740 1478 741 1479
rect 792 1478 794 1492
rect 799 1491 800 1492
rect 804 1491 805 1495
rect 871 1495 877 1496
rect 871 1494 872 1495
rect 799 1490 805 1491
rect 836 1492 872 1494
rect 836 1486 838 1492
rect 871 1491 872 1492
rect 876 1491 877 1495
rect 871 1490 877 1491
rect 898 1495 904 1496
rect 898 1491 899 1495
rect 903 1494 904 1495
rect 951 1495 957 1496
rect 951 1494 952 1495
rect 903 1492 952 1494
rect 903 1491 904 1492
rect 898 1490 904 1491
rect 951 1491 952 1492
rect 956 1491 957 1495
rect 1023 1495 1029 1496
rect 1023 1494 1024 1495
rect 951 1490 957 1491
rect 988 1492 1024 1494
rect 801 1484 838 1486
rect 854 1485 860 1486
rect 801 1480 803 1484
rect 854 1481 855 1485
rect 859 1481 860 1485
rect 854 1480 860 1481
rect 934 1485 940 1486
rect 934 1481 935 1485
rect 939 1481 940 1485
rect 934 1480 940 1481
rect 740 1476 794 1478
rect 799 1479 805 1480
rect 740 1475 741 1476
rect 735 1474 741 1475
rect 799 1475 800 1479
rect 804 1475 805 1479
rect 799 1474 805 1475
rect 834 1479 840 1480
rect 834 1475 835 1479
rect 839 1478 840 1479
rect 871 1479 877 1480
rect 871 1478 872 1479
rect 839 1476 872 1478
rect 839 1475 840 1476
rect 834 1474 840 1475
rect 871 1475 872 1476
rect 876 1475 877 1479
rect 871 1474 877 1475
rect 951 1479 957 1480
rect 951 1475 952 1479
rect 956 1478 957 1479
rect 988 1478 990 1492
rect 1023 1491 1024 1492
rect 1028 1491 1029 1495
rect 1095 1495 1101 1496
rect 1095 1494 1096 1495
rect 1023 1490 1029 1491
rect 1060 1492 1096 1494
rect 1006 1485 1012 1486
rect 1006 1481 1007 1485
rect 1011 1481 1012 1485
rect 1006 1480 1012 1481
rect 956 1476 990 1478
rect 1023 1479 1029 1480
rect 956 1475 957 1476
rect 951 1474 957 1475
rect 1023 1475 1024 1479
rect 1028 1478 1029 1479
rect 1060 1478 1062 1492
rect 1095 1491 1096 1492
rect 1100 1491 1101 1495
rect 1095 1490 1101 1491
rect 1167 1495 1173 1496
rect 1167 1491 1168 1495
rect 1172 1494 1173 1495
rect 1231 1495 1237 1496
rect 1172 1492 1202 1494
rect 1172 1491 1173 1492
rect 1167 1490 1173 1491
rect 1078 1485 1084 1486
rect 1078 1481 1079 1485
rect 1083 1481 1084 1485
rect 1078 1480 1084 1481
rect 1150 1485 1156 1486
rect 1150 1481 1151 1485
rect 1155 1481 1156 1485
rect 1150 1480 1156 1481
rect 1028 1476 1062 1478
rect 1095 1479 1101 1480
rect 1028 1475 1029 1476
rect 1023 1474 1029 1475
rect 1095 1475 1096 1479
rect 1100 1478 1101 1479
rect 1114 1479 1120 1480
rect 1114 1478 1115 1479
rect 1100 1476 1115 1478
rect 1100 1475 1101 1476
rect 1095 1474 1101 1475
rect 1114 1475 1115 1476
rect 1119 1475 1120 1479
rect 1114 1474 1120 1475
rect 1167 1479 1173 1480
rect 1167 1475 1168 1479
rect 1172 1478 1173 1479
rect 1200 1478 1202 1492
rect 1231 1491 1232 1495
rect 1236 1494 1237 1495
rect 1295 1495 1301 1496
rect 1236 1492 1266 1494
rect 1236 1491 1237 1492
rect 1231 1490 1237 1491
rect 1214 1485 1220 1486
rect 1214 1481 1215 1485
rect 1219 1481 1220 1485
rect 1214 1480 1220 1481
rect 1231 1479 1237 1480
rect 1231 1478 1232 1479
rect 1172 1476 1198 1478
rect 1200 1476 1232 1478
rect 1172 1475 1173 1476
rect 1167 1474 1173 1475
rect 599 1471 605 1472
rect 151 1467 157 1468
rect 110 1464 116 1465
rect 110 1460 111 1464
rect 115 1460 116 1464
rect 110 1459 116 1460
rect 134 1463 140 1464
rect 134 1459 135 1463
rect 139 1459 140 1463
rect 151 1463 152 1467
rect 156 1463 157 1467
rect 199 1467 205 1468
rect 151 1462 157 1463
rect 182 1463 188 1464
rect 134 1458 140 1459
rect 153 1458 155 1462
rect 182 1459 183 1463
rect 187 1459 188 1463
rect 199 1463 200 1467
rect 204 1466 205 1467
rect 218 1467 224 1468
rect 218 1466 219 1467
rect 204 1464 219 1466
rect 204 1463 205 1464
rect 199 1462 205 1463
rect 218 1463 219 1464
rect 223 1463 224 1467
rect 247 1467 253 1468
rect 218 1462 224 1463
rect 230 1463 236 1464
rect 182 1458 188 1459
rect 230 1459 231 1463
rect 235 1459 236 1463
rect 247 1463 248 1467
rect 252 1466 253 1467
rect 303 1467 309 1468
rect 303 1466 304 1467
rect 252 1464 261 1466
rect 296 1464 304 1466
rect 252 1463 253 1464
rect 247 1462 253 1463
rect 258 1463 264 1464
rect 230 1458 236 1459
rect 258 1459 259 1463
rect 263 1459 264 1463
rect 258 1458 264 1459
rect 286 1463 292 1464
rect 286 1459 287 1463
rect 291 1459 292 1463
rect 286 1458 292 1459
rect 153 1456 178 1458
rect 176 1454 178 1456
rect 296 1454 298 1464
rect 303 1463 304 1464
rect 308 1463 309 1467
rect 359 1467 365 1468
rect 359 1466 360 1467
rect 352 1464 360 1466
rect 303 1462 309 1463
rect 342 1463 348 1464
rect 342 1459 343 1463
rect 347 1459 348 1463
rect 342 1458 348 1459
rect 352 1454 354 1464
rect 359 1463 360 1464
rect 364 1463 365 1467
rect 415 1467 421 1468
rect 415 1466 416 1467
rect 408 1464 416 1466
rect 359 1462 365 1463
rect 398 1463 404 1464
rect 398 1459 399 1463
rect 403 1459 404 1463
rect 398 1458 404 1459
rect 408 1454 410 1464
rect 415 1463 416 1464
rect 420 1463 421 1467
rect 471 1467 477 1468
rect 415 1462 421 1463
rect 454 1463 460 1464
rect 454 1459 455 1463
rect 459 1459 460 1463
rect 471 1463 472 1467
rect 476 1466 477 1467
rect 482 1467 488 1468
rect 482 1466 483 1467
rect 476 1464 483 1466
rect 476 1463 477 1464
rect 471 1462 477 1463
rect 482 1463 483 1464
rect 487 1463 488 1467
rect 527 1467 533 1468
rect 527 1466 528 1467
rect 520 1464 528 1466
rect 482 1462 488 1463
rect 510 1463 516 1464
rect 454 1458 460 1459
rect 510 1459 511 1463
rect 515 1459 516 1463
rect 510 1458 516 1459
rect 520 1454 522 1464
rect 527 1463 528 1464
rect 532 1463 533 1467
rect 591 1467 597 1468
rect 591 1466 592 1467
rect 584 1464 592 1466
rect 527 1462 533 1463
rect 574 1463 580 1464
rect 574 1459 575 1463
rect 579 1459 580 1463
rect 574 1458 580 1459
rect 584 1454 586 1464
rect 591 1463 592 1464
rect 596 1463 597 1467
rect 599 1467 600 1471
rect 604 1470 605 1471
rect 1196 1470 1198 1476
rect 1231 1475 1232 1476
rect 1236 1475 1237 1479
rect 1264 1478 1266 1492
rect 1295 1491 1296 1495
rect 1300 1494 1301 1495
rect 1367 1495 1373 1496
rect 1300 1492 1334 1494
rect 1300 1491 1301 1492
rect 1295 1490 1301 1491
rect 1278 1485 1284 1486
rect 1278 1481 1279 1485
rect 1283 1481 1284 1485
rect 1278 1480 1284 1481
rect 1295 1479 1301 1480
rect 1295 1478 1296 1479
rect 1264 1476 1296 1478
rect 1231 1474 1237 1475
rect 1295 1475 1296 1476
rect 1300 1475 1301 1479
rect 1332 1478 1334 1492
rect 1367 1491 1368 1495
rect 1372 1494 1373 1495
rect 1438 1495 1445 1496
rect 1372 1492 1406 1494
rect 1372 1491 1373 1492
rect 1367 1490 1373 1491
rect 1350 1485 1356 1486
rect 1350 1481 1351 1485
rect 1355 1481 1356 1485
rect 1350 1480 1356 1481
rect 1367 1479 1373 1480
rect 1367 1478 1368 1479
rect 1332 1476 1368 1478
rect 1295 1474 1301 1475
rect 1367 1475 1368 1476
rect 1372 1475 1373 1479
rect 1404 1478 1406 1492
rect 1438 1491 1439 1495
rect 1444 1491 1445 1495
rect 1438 1490 1445 1491
rect 1511 1495 1517 1496
rect 1511 1491 1512 1495
rect 1516 1494 1517 1495
rect 1558 1495 1565 1496
rect 1516 1492 1538 1494
rect 1516 1491 1517 1492
rect 1511 1490 1517 1491
rect 1422 1485 1428 1486
rect 1422 1481 1423 1485
rect 1427 1481 1428 1485
rect 1422 1480 1428 1481
rect 1494 1485 1500 1486
rect 1494 1481 1495 1485
rect 1499 1481 1500 1485
rect 1494 1480 1500 1481
rect 1439 1479 1445 1480
rect 1439 1478 1440 1479
rect 1404 1476 1440 1478
rect 1367 1474 1373 1475
rect 1439 1475 1440 1476
rect 1444 1475 1445 1479
rect 1439 1474 1445 1475
rect 1510 1479 1517 1480
rect 1510 1475 1511 1479
rect 1516 1475 1517 1479
rect 1536 1478 1538 1492
rect 1558 1491 1559 1495
rect 1564 1491 1565 1495
rect 1558 1490 1565 1491
rect 1542 1485 1548 1486
rect 1542 1481 1543 1485
rect 1547 1481 1548 1485
rect 1542 1480 1548 1481
rect 1582 1484 1588 1485
rect 1582 1480 1583 1484
rect 1587 1480 1588 1484
rect 1559 1479 1565 1480
rect 1582 1479 1588 1480
rect 1559 1478 1560 1479
rect 1536 1476 1560 1478
rect 1510 1474 1517 1475
rect 1559 1475 1560 1476
rect 1564 1475 1565 1479
rect 1559 1474 1565 1475
rect 1248 1472 1290 1474
rect 1248 1470 1250 1472
rect 604 1468 642 1470
rect 1196 1468 1250 1470
rect 1288 1470 1290 1472
rect 1328 1472 1362 1474
rect 1328 1470 1330 1472
rect 1288 1468 1330 1470
rect 1360 1470 1362 1472
rect 1408 1472 1426 1474
rect 1408 1470 1410 1472
rect 1360 1468 1410 1470
rect 1423 1471 1429 1472
rect 604 1467 605 1468
rect 599 1466 605 1467
rect 640 1466 642 1468
rect 647 1467 653 1468
rect 647 1466 648 1467
rect 640 1464 648 1466
rect 591 1462 597 1463
rect 630 1463 636 1464
rect 630 1459 631 1463
rect 635 1459 636 1463
rect 647 1463 648 1464
rect 652 1463 653 1467
rect 698 1467 709 1468
rect 647 1462 653 1463
rect 686 1463 692 1464
rect 630 1458 636 1459
rect 686 1459 687 1463
rect 691 1459 692 1463
rect 698 1463 699 1467
rect 703 1463 704 1467
rect 708 1463 709 1467
rect 767 1467 773 1468
rect 767 1466 768 1467
rect 760 1464 768 1466
rect 698 1462 709 1463
rect 750 1463 756 1464
rect 686 1458 692 1459
rect 750 1459 751 1463
rect 755 1459 756 1463
rect 750 1458 756 1459
rect 760 1454 762 1464
rect 767 1463 768 1464
rect 772 1463 773 1467
rect 831 1467 837 1468
rect 831 1466 832 1467
rect 824 1464 832 1466
rect 767 1462 773 1463
rect 814 1463 820 1464
rect 814 1459 815 1463
rect 819 1459 820 1463
rect 814 1458 820 1459
rect 824 1454 826 1464
rect 831 1463 832 1464
rect 836 1463 837 1467
rect 895 1467 904 1468
rect 831 1462 837 1463
rect 878 1463 884 1464
rect 878 1459 879 1463
rect 883 1459 884 1463
rect 895 1463 896 1467
rect 903 1463 904 1467
rect 959 1467 965 1468
rect 959 1466 960 1467
rect 952 1464 960 1466
rect 895 1462 904 1463
rect 942 1463 948 1464
rect 878 1458 884 1459
rect 942 1459 943 1463
rect 947 1459 948 1463
rect 942 1458 948 1459
rect 952 1454 954 1464
rect 959 1463 960 1464
rect 964 1463 965 1467
rect 1031 1467 1037 1468
rect 1031 1466 1032 1467
rect 1024 1464 1032 1466
rect 959 1462 965 1463
rect 1014 1463 1020 1464
rect 1014 1459 1015 1463
rect 1019 1459 1020 1463
rect 1014 1458 1020 1459
rect 1024 1454 1026 1464
rect 1031 1463 1032 1464
rect 1036 1463 1037 1467
rect 1103 1467 1109 1468
rect 1103 1466 1104 1467
rect 1096 1464 1104 1466
rect 1031 1462 1037 1463
rect 1086 1463 1092 1464
rect 1086 1459 1087 1463
rect 1091 1459 1092 1463
rect 1086 1458 1092 1459
rect 1096 1454 1098 1464
rect 1103 1463 1104 1464
rect 1108 1463 1109 1467
rect 1174 1467 1181 1468
rect 1103 1462 1109 1463
rect 1158 1463 1164 1464
rect 1158 1459 1159 1463
rect 1163 1459 1164 1463
rect 1174 1463 1175 1467
rect 1180 1463 1181 1467
rect 1255 1467 1261 1468
rect 1255 1466 1256 1467
rect 1248 1464 1256 1466
rect 1174 1462 1181 1463
rect 1238 1463 1244 1464
rect 1158 1458 1164 1459
rect 1238 1459 1239 1463
rect 1243 1459 1244 1463
rect 1238 1458 1244 1459
rect 1248 1454 1250 1464
rect 1255 1463 1256 1464
rect 1260 1463 1261 1467
rect 1335 1467 1341 1468
rect 1335 1466 1336 1467
rect 1328 1464 1336 1466
rect 1255 1462 1261 1463
rect 1318 1463 1324 1464
rect 1318 1459 1319 1463
rect 1323 1459 1324 1463
rect 1318 1458 1324 1459
rect 1328 1454 1330 1464
rect 1335 1463 1336 1464
rect 1340 1463 1341 1467
rect 1415 1467 1421 1468
rect 1415 1466 1416 1467
rect 1408 1464 1416 1466
rect 1335 1462 1341 1463
rect 1398 1463 1404 1464
rect 1398 1459 1399 1463
rect 1403 1459 1404 1463
rect 1398 1458 1404 1459
rect 1408 1454 1410 1464
rect 1415 1463 1416 1464
rect 1420 1463 1421 1467
rect 1423 1467 1424 1471
rect 1428 1467 1429 1471
rect 1423 1466 1429 1467
rect 1495 1467 1501 1468
rect 1415 1462 1421 1463
rect 1478 1463 1484 1464
rect 1478 1459 1479 1463
rect 1483 1459 1484 1463
rect 1495 1463 1496 1467
rect 1500 1463 1501 1467
rect 1558 1467 1565 1468
rect 1495 1462 1501 1463
rect 1542 1463 1548 1464
rect 1478 1458 1484 1459
rect 1497 1458 1499 1462
rect 1542 1459 1543 1463
rect 1547 1459 1548 1463
rect 1558 1463 1559 1467
rect 1564 1463 1565 1467
rect 1558 1462 1565 1463
rect 1582 1464 1588 1465
rect 1582 1460 1583 1464
rect 1587 1460 1588 1464
rect 1582 1459 1588 1460
rect 1542 1458 1548 1459
rect 1497 1456 1538 1458
rect 176 1452 194 1454
rect 259 1452 298 1454
rect 332 1452 354 1454
rect 388 1452 410 1454
rect 500 1452 522 1454
rect 560 1452 586 1454
rect 736 1452 762 1454
rect 801 1452 826 1454
rect 928 1452 954 1454
rect 996 1452 1026 1454
rect 1064 1452 1098 1454
rect 1216 1452 1250 1454
rect 1296 1452 1330 1454
rect 1376 1452 1410 1454
rect 1536 1454 1538 1456
rect 1536 1452 1563 1454
rect 150 1451 157 1452
rect 110 1447 116 1448
rect 110 1443 111 1447
rect 115 1443 116 1447
rect 150 1447 151 1451
rect 156 1447 157 1451
rect 192 1450 194 1452
rect 199 1451 205 1452
rect 199 1450 200 1451
rect 192 1448 200 1450
rect 150 1446 157 1447
rect 199 1447 200 1448
rect 204 1447 205 1451
rect 199 1446 205 1447
rect 247 1451 253 1452
rect 247 1447 248 1451
rect 252 1450 253 1451
rect 259 1450 261 1452
rect 252 1448 261 1450
rect 303 1451 309 1452
rect 252 1447 253 1448
rect 247 1446 253 1447
rect 303 1447 304 1451
rect 308 1450 309 1451
rect 332 1450 334 1452
rect 308 1448 334 1450
rect 359 1451 365 1452
rect 308 1447 309 1448
rect 303 1446 309 1447
rect 359 1447 360 1451
rect 364 1450 365 1451
rect 388 1450 390 1452
rect 415 1451 421 1452
rect 415 1450 416 1451
rect 364 1448 390 1450
rect 408 1448 416 1450
rect 364 1447 365 1448
rect 359 1446 365 1447
rect 110 1442 116 1443
rect 134 1445 140 1446
rect 134 1441 135 1445
rect 139 1441 140 1445
rect 134 1440 140 1441
rect 182 1445 188 1446
rect 182 1441 183 1445
rect 187 1441 188 1445
rect 182 1440 188 1441
rect 230 1445 236 1446
rect 230 1441 231 1445
rect 235 1441 236 1445
rect 230 1440 236 1441
rect 286 1445 292 1446
rect 286 1441 287 1445
rect 291 1441 292 1445
rect 286 1440 292 1441
rect 342 1445 348 1446
rect 342 1441 343 1445
rect 347 1441 348 1445
rect 342 1440 348 1441
rect 398 1445 404 1446
rect 398 1441 399 1445
rect 403 1441 404 1445
rect 398 1440 404 1441
rect 274 1439 280 1440
rect 274 1435 275 1439
rect 279 1438 280 1439
rect 408 1438 410 1448
rect 415 1447 416 1448
rect 420 1447 421 1451
rect 415 1446 421 1447
rect 471 1451 477 1452
rect 471 1447 472 1451
rect 476 1450 477 1451
rect 500 1450 502 1452
rect 476 1448 502 1450
rect 527 1451 533 1452
rect 476 1447 477 1448
rect 471 1446 477 1447
rect 527 1447 528 1451
rect 532 1450 533 1451
rect 560 1450 562 1452
rect 532 1448 562 1450
rect 591 1451 597 1452
rect 532 1447 533 1448
rect 527 1446 533 1447
rect 591 1447 592 1451
rect 596 1450 597 1451
rect 599 1451 605 1452
rect 599 1450 600 1451
rect 596 1448 600 1450
rect 596 1447 597 1448
rect 591 1446 597 1447
rect 599 1447 600 1448
rect 604 1447 605 1451
rect 599 1446 605 1447
rect 642 1451 653 1452
rect 642 1447 643 1451
rect 647 1447 648 1451
rect 652 1447 653 1451
rect 642 1446 653 1447
rect 703 1451 709 1452
rect 703 1447 704 1451
rect 708 1450 709 1451
rect 736 1450 738 1452
rect 708 1448 738 1450
rect 767 1451 773 1452
rect 708 1447 709 1448
rect 703 1446 709 1447
rect 767 1447 768 1451
rect 772 1450 773 1451
rect 801 1450 803 1452
rect 772 1448 803 1450
rect 831 1451 840 1452
rect 772 1447 773 1448
rect 767 1446 773 1447
rect 831 1447 832 1451
rect 839 1447 840 1451
rect 831 1446 840 1447
rect 895 1451 901 1452
rect 895 1447 896 1451
rect 900 1450 901 1451
rect 928 1450 930 1452
rect 900 1448 930 1450
rect 959 1451 965 1452
rect 900 1447 901 1448
rect 895 1446 901 1447
rect 959 1447 960 1451
rect 964 1450 965 1451
rect 996 1450 998 1452
rect 964 1448 998 1450
rect 1031 1451 1037 1452
rect 964 1447 965 1448
rect 959 1446 965 1447
rect 1031 1447 1032 1451
rect 1036 1450 1037 1451
rect 1064 1450 1066 1452
rect 1036 1448 1066 1450
rect 1102 1451 1109 1452
rect 1036 1447 1037 1448
rect 1031 1446 1037 1447
rect 1102 1447 1103 1451
rect 1108 1447 1109 1451
rect 1102 1446 1109 1447
rect 1175 1451 1181 1452
rect 1175 1447 1176 1451
rect 1180 1450 1181 1451
rect 1216 1450 1218 1452
rect 1180 1448 1218 1450
rect 1255 1451 1261 1452
rect 1180 1447 1181 1448
rect 1175 1446 1181 1447
rect 1255 1447 1256 1451
rect 1260 1450 1261 1451
rect 1296 1450 1298 1452
rect 1260 1448 1298 1450
rect 1335 1451 1341 1452
rect 1260 1447 1261 1448
rect 1255 1446 1261 1447
rect 1335 1447 1336 1451
rect 1340 1450 1341 1451
rect 1376 1450 1378 1452
rect 1340 1448 1378 1450
rect 1415 1451 1421 1452
rect 1340 1447 1341 1448
rect 1335 1446 1341 1447
rect 1415 1447 1416 1451
rect 1420 1450 1421 1451
rect 1423 1451 1429 1452
rect 1423 1450 1424 1451
rect 1420 1448 1424 1450
rect 1420 1447 1421 1448
rect 1415 1446 1421 1447
rect 1423 1447 1424 1448
rect 1428 1447 1429 1451
rect 1423 1446 1429 1447
rect 1495 1451 1501 1452
rect 1495 1447 1496 1451
rect 1500 1450 1501 1451
rect 1526 1451 1532 1452
rect 1526 1450 1527 1451
rect 1500 1448 1527 1450
rect 1500 1447 1501 1448
rect 1495 1446 1501 1447
rect 1526 1447 1527 1448
rect 1531 1447 1532 1451
rect 1526 1446 1532 1447
rect 1559 1451 1565 1452
rect 1559 1447 1560 1451
rect 1564 1447 1565 1451
rect 1559 1446 1565 1447
rect 1582 1447 1588 1448
rect 454 1445 460 1446
rect 454 1441 455 1445
rect 459 1441 460 1445
rect 454 1440 460 1441
rect 510 1445 516 1446
rect 510 1441 511 1445
rect 515 1441 516 1445
rect 510 1440 516 1441
rect 574 1445 580 1446
rect 574 1441 575 1445
rect 579 1441 580 1445
rect 574 1440 580 1441
rect 630 1445 636 1446
rect 630 1441 631 1445
rect 635 1441 636 1445
rect 630 1440 636 1441
rect 686 1445 692 1446
rect 686 1441 687 1445
rect 691 1441 692 1445
rect 686 1440 692 1441
rect 750 1445 756 1446
rect 750 1441 751 1445
rect 755 1441 756 1445
rect 750 1440 756 1441
rect 814 1445 820 1446
rect 814 1441 815 1445
rect 819 1441 820 1445
rect 814 1440 820 1441
rect 878 1445 884 1446
rect 878 1441 879 1445
rect 883 1441 884 1445
rect 878 1440 884 1441
rect 942 1445 948 1446
rect 942 1441 943 1445
rect 947 1441 948 1445
rect 942 1440 948 1441
rect 1014 1445 1020 1446
rect 1014 1441 1015 1445
rect 1019 1441 1020 1445
rect 1014 1440 1020 1441
rect 1086 1445 1092 1446
rect 1086 1441 1087 1445
rect 1091 1441 1092 1445
rect 1086 1440 1092 1441
rect 1158 1445 1164 1446
rect 1158 1441 1159 1445
rect 1163 1441 1164 1445
rect 1158 1440 1164 1441
rect 1238 1445 1244 1446
rect 1238 1441 1239 1445
rect 1243 1441 1244 1445
rect 1238 1440 1244 1441
rect 1318 1445 1324 1446
rect 1318 1441 1319 1445
rect 1323 1441 1324 1445
rect 1318 1440 1324 1441
rect 1398 1445 1404 1446
rect 1398 1441 1399 1445
rect 1403 1441 1404 1445
rect 1398 1440 1404 1441
rect 1478 1445 1484 1446
rect 1478 1441 1479 1445
rect 1483 1441 1484 1445
rect 1478 1440 1484 1441
rect 1542 1445 1548 1446
rect 1542 1441 1543 1445
rect 1547 1441 1548 1445
rect 1582 1443 1583 1447
rect 1587 1443 1588 1447
rect 1582 1442 1588 1443
rect 1542 1440 1548 1441
rect 279 1436 410 1438
rect 910 1439 916 1440
rect 279 1435 280 1436
rect 274 1434 280 1435
rect 910 1435 911 1439
rect 915 1438 916 1439
rect 1362 1439 1368 1440
rect 915 1436 1078 1438
rect 915 1435 916 1436
rect 910 1434 916 1435
rect 134 1431 140 1432
rect 110 1429 116 1430
rect 110 1425 111 1429
rect 115 1425 116 1429
rect 134 1427 135 1431
rect 139 1427 140 1431
rect 134 1426 140 1427
rect 182 1431 188 1432
rect 182 1427 183 1431
rect 187 1427 188 1431
rect 182 1426 188 1427
rect 254 1431 260 1432
rect 254 1427 255 1431
rect 259 1427 260 1431
rect 254 1426 260 1427
rect 326 1431 332 1432
rect 326 1427 327 1431
rect 331 1427 332 1431
rect 326 1426 332 1427
rect 398 1431 404 1432
rect 398 1427 399 1431
rect 403 1427 404 1431
rect 398 1426 404 1427
rect 470 1431 476 1432
rect 470 1427 471 1431
rect 475 1427 476 1431
rect 470 1426 476 1427
rect 542 1431 548 1432
rect 542 1427 543 1431
rect 547 1427 548 1431
rect 542 1426 548 1427
rect 614 1431 620 1432
rect 614 1427 615 1431
rect 619 1427 620 1431
rect 614 1426 620 1427
rect 678 1431 684 1432
rect 678 1427 679 1431
rect 683 1427 684 1431
rect 678 1426 684 1427
rect 742 1431 748 1432
rect 742 1427 743 1431
rect 747 1427 748 1431
rect 742 1426 748 1427
rect 814 1431 820 1432
rect 814 1427 815 1431
rect 819 1427 820 1431
rect 814 1426 820 1427
rect 878 1431 884 1432
rect 878 1427 879 1431
rect 883 1427 884 1431
rect 878 1426 884 1427
rect 950 1431 956 1432
rect 950 1427 951 1431
rect 955 1427 956 1431
rect 950 1426 956 1427
rect 1022 1431 1028 1432
rect 1022 1427 1023 1431
rect 1027 1427 1028 1431
rect 1022 1426 1028 1427
rect 110 1424 116 1425
rect 151 1423 157 1424
rect 151 1419 152 1423
rect 156 1419 157 1423
rect 151 1418 157 1419
rect 194 1423 205 1424
rect 194 1419 195 1423
rect 199 1419 200 1423
rect 204 1419 205 1423
rect 194 1418 205 1419
rect 271 1423 277 1424
rect 271 1419 272 1423
rect 276 1422 277 1423
rect 343 1423 349 1424
rect 276 1420 310 1422
rect 276 1419 277 1420
rect 271 1418 277 1419
rect 153 1414 155 1418
rect 134 1413 140 1414
rect 110 1412 116 1413
rect 110 1408 111 1412
rect 115 1408 116 1412
rect 134 1409 135 1413
rect 139 1409 140 1413
rect 153 1412 178 1414
rect 134 1408 140 1409
rect 110 1407 116 1408
rect 150 1407 157 1408
rect 150 1403 151 1407
rect 156 1403 157 1407
rect 176 1406 178 1412
rect 182 1413 188 1414
rect 182 1409 183 1413
rect 187 1409 188 1413
rect 182 1408 188 1409
rect 254 1413 260 1414
rect 254 1409 255 1413
rect 259 1409 260 1413
rect 254 1408 260 1409
rect 199 1407 205 1408
rect 199 1406 200 1407
rect 176 1404 200 1406
rect 150 1402 157 1403
rect 199 1403 200 1404
rect 204 1403 205 1407
rect 199 1402 205 1403
rect 262 1407 268 1408
rect 262 1403 263 1407
rect 267 1406 268 1407
rect 271 1407 277 1408
rect 271 1406 272 1407
rect 267 1404 272 1406
rect 267 1403 268 1404
rect 262 1402 268 1403
rect 271 1403 272 1404
rect 276 1403 277 1407
rect 308 1406 310 1420
rect 343 1419 344 1423
rect 348 1422 349 1423
rect 414 1423 421 1424
rect 348 1420 410 1422
rect 348 1419 349 1420
rect 343 1418 349 1419
rect 326 1413 332 1414
rect 326 1409 327 1413
rect 331 1409 332 1413
rect 326 1408 332 1409
rect 398 1413 404 1414
rect 398 1409 399 1413
rect 403 1409 404 1413
rect 398 1408 404 1409
rect 343 1407 349 1408
rect 343 1406 344 1407
rect 308 1404 344 1406
rect 271 1402 277 1403
rect 343 1403 344 1404
rect 348 1403 349 1407
rect 408 1406 410 1420
rect 414 1419 415 1423
rect 420 1419 421 1423
rect 414 1418 421 1419
rect 482 1423 493 1424
rect 482 1419 483 1423
rect 487 1419 488 1423
rect 492 1419 493 1423
rect 559 1423 565 1424
rect 559 1422 560 1423
rect 482 1418 493 1419
rect 524 1420 560 1422
rect 470 1413 476 1414
rect 470 1409 471 1413
rect 475 1409 476 1413
rect 470 1408 476 1409
rect 415 1407 421 1408
rect 415 1406 416 1407
rect 408 1404 416 1406
rect 343 1402 349 1403
rect 415 1403 416 1404
rect 420 1403 421 1407
rect 415 1402 421 1403
rect 487 1407 493 1408
rect 487 1403 488 1407
rect 492 1406 493 1407
rect 524 1406 526 1420
rect 559 1419 560 1420
rect 564 1419 565 1423
rect 631 1423 637 1424
rect 631 1422 632 1423
rect 559 1418 565 1419
rect 596 1420 632 1422
rect 542 1413 548 1414
rect 542 1409 543 1413
rect 547 1409 548 1413
rect 542 1408 548 1409
rect 492 1404 526 1406
rect 559 1407 565 1408
rect 492 1403 493 1404
rect 487 1402 493 1403
rect 559 1403 560 1407
rect 564 1406 565 1407
rect 596 1406 598 1420
rect 631 1419 632 1420
rect 636 1419 637 1423
rect 631 1418 637 1419
rect 695 1423 704 1424
rect 695 1419 696 1423
rect 703 1419 704 1423
rect 759 1423 765 1424
rect 759 1422 760 1423
rect 695 1418 704 1419
rect 732 1420 760 1422
rect 614 1413 620 1414
rect 614 1409 615 1413
rect 619 1409 620 1413
rect 678 1413 684 1414
rect 642 1411 648 1412
rect 642 1410 643 1411
rect 614 1408 620 1409
rect 633 1408 643 1410
rect 564 1404 598 1406
rect 631 1407 637 1408
rect 564 1403 565 1404
rect 559 1402 565 1403
rect 631 1403 632 1407
rect 636 1403 637 1407
rect 642 1407 643 1408
rect 647 1407 648 1411
rect 678 1409 679 1413
rect 683 1409 684 1413
rect 678 1408 684 1409
rect 642 1406 648 1407
rect 695 1407 701 1408
rect 631 1402 637 1403
rect 695 1403 696 1407
rect 700 1406 701 1407
rect 732 1406 734 1420
rect 759 1419 760 1420
rect 764 1419 765 1423
rect 831 1423 837 1424
rect 831 1422 832 1423
rect 759 1418 765 1419
rect 800 1420 832 1422
rect 742 1413 748 1414
rect 742 1409 743 1413
rect 747 1409 748 1413
rect 742 1408 748 1409
rect 700 1404 734 1406
rect 759 1407 765 1408
rect 700 1403 701 1404
rect 695 1402 701 1403
rect 759 1403 760 1407
rect 764 1406 765 1407
rect 800 1406 802 1420
rect 831 1419 832 1420
rect 836 1419 837 1423
rect 831 1418 837 1419
rect 895 1423 901 1424
rect 895 1419 896 1423
rect 900 1422 901 1423
rect 967 1423 973 1424
rect 900 1420 962 1422
rect 900 1419 901 1420
rect 895 1418 901 1419
rect 960 1414 962 1420
rect 967 1419 968 1423
rect 972 1422 973 1423
rect 1039 1423 1045 1424
rect 972 1420 1034 1422
rect 972 1419 973 1420
rect 967 1418 973 1419
rect 814 1413 820 1414
rect 814 1409 815 1413
rect 819 1409 820 1413
rect 814 1408 820 1409
rect 878 1413 884 1414
rect 878 1409 879 1413
rect 883 1409 884 1413
rect 878 1408 884 1409
rect 950 1413 956 1414
rect 950 1409 951 1413
rect 955 1409 956 1413
rect 960 1412 971 1414
rect 969 1410 971 1412
rect 1022 1413 1028 1414
rect 950 1408 956 1409
rect 967 1409 973 1410
rect 764 1404 802 1406
rect 831 1407 837 1408
rect 764 1403 765 1404
rect 759 1402 765 1403
rect 831 1403 832 1407
rect 836 1406 837 1407
rect 854 1407 860 1408
rect 854 1406 855 1407
rect 836 1404 855 1406
rect 836 1403 837 1404
rect 831 1402 837 1403
rect 854 1403 855 1404
rect 859 1403 860 1407
rect 854 1402 860 1403
rect 895 1407 901 1408
rect 895 1403 896 1407
rect 900 1406 901 1407
rect 900 1404 930 1406
rect 967 1405 968 1409
rect 972 1405 973 1409
rect 1022 1409 1023 1413
rect 1027 1409 1028 1413
rect 1022 1408 1028 1409
rect 967 1404 973 1405
rect 1032 1406 1034 1420
rect 1039 1419 1040 1423
rect 1044 1422 1045 1423
rect 1076 1422 1078 1436
rect 1362 1435 1363 1439
rect 1367 1438 1368 1439
rect 1367 1436 1563 1438
rect 1367 1435 1368 1436
rect 1362 1434 1368 1435
rect 1094 1431 1100 1432
rect 1094 1427 1095 1431
rect 1099 1427 1100 1431
rect 1094 1426 1100 1427
rect 1158 1431 1164 1432
rect 1158 1427 1159 1431
rect 1163 1427 1164 1431
rect 1158 1426 1164 1427
rect 1222 1431 1228 1432
rect 1222 1427 1223 1431
rect 1227 1427 1228 1431
rect 1222 1426 1228 1427
rect 1286 1431 1292 1432
rect 1286 1427 1287 1431
rect 1291 1427 1292 1431
rect 1286 1426 1292 1427
rect 1342 1431 1348 1432
rect 1342 1427 1343 1431
rect 1347 1427 1348 1431
rect 1342 1426 1348 1427
rect 1398 1431 1404 1432
rect 1398 1427 1399 1431
rect 1403 1427 1404 1431
rect 1398 1426 1404 1427
rect 1454 1431 1460 1432
rect 1454 1427 1455 1431
rect 1459 1427 1460 1431
rect 1454 1426 1460 1427
rect 1510 1431 1516 1432
rect 1510 1427 1511 1431
rect 1515 1427 1516 1431
rect 1510 1426 1516 1427
rect 1542 1431 1548 1432
rect 1542 1427 1543 1431
rect 1547 1427 1548 1431
rect 1542 1426 1548 1427
rect 1561 1424 1563 1436
rect 1582 1429 1588 1430
rect 1582 1425 1583 1429
rect 1587 1425 1588 1429
rect 1582 1424 1588 1425
rect 1111 1423 1117 1424
rect 1111 1422 1112 1423
rect 1044 1420 1074 1422
rect 1076 1420 1112 1422
rect 1044 1419 1045 1420
rect 1039 1418 1045 1419
rect 1039 1407 1045 1408
rect 1039 1406 1040 1407
rect 1032 1404 1040 1406
rect 900 1403 901 1404
rect 895 1402 901 1403
rect 928 1402 930 1404
rect 1039 1403 1040 1404
rect 1044 1403 1045 1407
rect 1072 1406 1074 1420
rect 1111 1419 1112 1420
rect 1116 1419 1117 1423
rect 1111 1418 1117 1419
rect 1174 1423 1181 1424
rect 1174 1419 1175 1423
rect 1180 1419 1181 1423
rect 1239 1423 1245 1424
rect 1239 1422 1240 1423
rect 1174 1418 1181 1419
rect 1209 1420 1240 1422
rect 1094 1413 1100 1414
rect 1094 1409 1095 1413
rect 1099 1409 1100 1413
rect 1094 1408 1100 1409
rect 1158 1413 1164 1414
rect 1158 1409 1159 1413
rect 1163 1409 1164 1413
rect 1158 1408 1164 1409
rect 1111 1407 1117 1408
rect 1111 1406 1112 1407
rect 1072 1404 1112 1406
rect 1039 1402 1045 1403
rect 1111 1403 1112 1404
rect 1116 1403 1117 1407
rect 1111 1402 1117 1403
rect 1175 1407 1181 1408
rect 1175 1403 1176 1407
rect 1180 1406 1181 1407
rect 1209 1406 1211 1420
rect 1239 1419 1240 1420
rect 1244 1419 1245 1423
rect 1303 1423 1309 1424
rect 1303 1422 1304 1423
rect 1239 1418 1245 1419
rect 1273 1420 1304 1422
rect 1222 1413 1228 1414
rect 1222 1409 1223 1413
rect 1227 1409 1228 1413
rect 1222 1408 1228 1409
rect 1180 1404 1211 1406
rect 1239 1407 1245 1408
rect 1180 1403 1181 1404
rect 1175 1402 1181 1403
rect 1239 1403 1240 1407
rect 1244 1406 1245 1407
rect 1273 1406 1275 1420
rect 1303 1419 1304 1420
rect 1308 1419 1309 1423
rect 1303 1418 1309 1419
rect 1359 1423 1365 1424
rect 1359 1419 1360 1423
rect 1364 1422 1365 1423
rect 1415 1423 1421 1424
rect 1364 1420 1390 1422
rect 1364 1419 1365 1420
rect 1359 1418 1365 1419
rect 1286 1413 1292 1414
rect 1286 1409 1287 1413
rect 1291 1409 1292 1413
rect 1286 1408 1292 1409
rect 1342 1413 1348 1414
rect 1342 1409 1343 1413
rect 1347 1409 1348 1413
rect 1342 1408 1348 1409
rect 1244 1404 1275 1406
rect 1303 1407 1312 1408
rect 1244 1403 1245 1404
rect 1239 1402 1245 1403
rect 1303 1403 1304 1407
rect 1311 1403 1312 1407
rect 1303 1402 1312 1403
rect 1359 1407 1368 1408
rect 1359 1403 1360 1407
rect 1367 1403 1368 1407
rect 1388 1406 1390 1420
rect 1415 1419 1416 1423
rect 1420 1422 1421 1423
rect 1471 1423 1477 1424
rect 1420 1420 1466 1422
rect 1420 1419 1421 1420
rect 1415 1418 1421 1419
rect 1398 1413 1404 1414
rect 1398 1409 1399 1413
rect 1403 1409 1404 1413
rect 1398 1408 1404 1409
rect 1454 1413 1460 1414
rect 1454 1409 1455 1413
rect 1459 1409 1460 1413
rect 1454 1408 1460 1409
rect 1415 1407 1421 1408
rect 1415 1406 1416 1407
rect 1388 1404 1416 1406
rect 1359 1402 1368 1403
rect 1415 1403 1416 1404
rect 1420 1403 1421 1407
rect 1464 1406 1466 1420
rect 1471 1419 1472 1423
rect 1476 1422 1477 1423
rect 1494 1423 1500 1424
rect 1494 1422 1495 1423
rect 1476 1420 1495 1422
rect 1476 1419 1477 1420
rect 1471 1418 1477 1419
rect 1494 1419 1495 1420
rect 1499 1419 1500 1423
rect 1494 1418 1500 1419
rect 1527 1423 1533 1424
rect 1527 1419 1528 1423
rect 1532 1422 1533 1423
rect 1559 1423 1565 1424
rect 1532 1420 1554 1422
rect 1532 1419 1533 1420
rect 1527 1418 1533 1419
rect 1510 1413 1516 1414
rect 1510 1409 1511 1413
rect 1515 1409 1516 1413
rect 1510 1408 1516 1409
rect 1542 1413 1548 1414
rect 1542 1409 1543 1413
rect 1547 1409 1548 1413
rect 1542 1408 1548 1409
rect 1471 1407 1477 1408
rect 1471 1406 1472 1407
rect 1464 1404 1472 1406
rect 1415 1402 1421 1403
rect 1471 1403 1472 1404
rect 1476 1403 1477 1407
rect 1471 1402 1477 1403
rect 1526 1407 1533 1408
rect 1526 1403 1527 1407
rect 1532 1403 1533 1407
rect 1552 1406 1554 1420
rect 1559 1419 1560 1423
rect 1564 1419 1565 1423
rect 1559 1418 1565 1419
rect 1582 1412 1588 1413
rect 1582 1408 1583 1412
rect 1587 1408 1588 1412
rect 1559 1407 1565 1408
rect 1582 1407 1588 1408
rect 1559 1406 1560 1407
rect 1552 1404 1560 1406
rect 1526 1402 1533 1403
rect 1559 1403 1560 1404
rect 1564 1403 1565 1407
rect 1559 1402 1565 1403
rect 928 1400 1027 1402
rect 1025 1398 1027 1400
rect 1048 1400 1106 1402
rect 1048 1398 1050 1400
rect 1025 1396 1050 1398
rect 1102 1399 1108 1400
rect 151 1395 157 1396
rect 110 1392 116 1393
rect 110 1388 111 1392
rect 115 1388 116 1392
rect 110 1387 116 1388
rect 134 1391 140 1392
rect 134 1387 135 1391
rect 139 1387 140 1391
rect 151 1391 152 1395
rect 156 1391 157 1395
rect 191 1395 200 1396
rect 151 1390 157 1391
rect 174 1391 180 1392
rect 134 1386 140 1387
rect 153 1386 155 1390
rect 174 1387 175 1391
rect 179 1387 180 1391
rect 191 1391 192 1395
rect 199 1391 200 1395
rect 263 1395 269 1396
rect 191 1390 200 1391
rect 246 1391 252 1392
rect 174 1386 180 1387
rect 246 1387 247 1391
rect 251 1387 252 1391
rect 263 1391 264 1395
rect 268 1394 269 1395
rect 335 1395 341 1396
rect 268 1392 315 1394
rect 268 1391 269 1392
rect 263 1390 269 1391
rect 246 1386 252 1387
rect 153 1384 170 1386
rect 168 1382 170 1384
rect 313 1382 315 1392
rect 318 1391 324 1392
rect 318 1387 319 1391
rect 323 1387 324 1391
rect 335 1391 336 1395
rect 340 1394 341 1395
rect 407 1395 413 1396
rect 340 1392 378 1394
rect 340 1391 341 1392
rect 335 1390 341 1391
rect 318 1386 324 1387
rect 376 1382 378 1392
rect 390 1391 396 1392
rect 390 1387 391 1391
rect 395 1387 396 1391
rect 407 1391 408 1395
rect 412 1394 413 1395
rect 446 1395 452 1396
rect 446 1394 447 1395
rect 412 1392 447 1394
rect 412 1391 413 1392
rect 407 1390 413 1391
rect 446 1391 447 1392
rect 451 1391 452 1395
rect 471 1395 477 1396
rect 446 1390 452 1391
rect 454 1391 460 1392
rect 390 1386 396 1387
rect 454 1387 455 1391
rect 459 1387 460 1391
rect 471 1391 472 1395
rect 476 1394 477 1395
rect 482 1395 488 1396
rect 482 1394 483 1395
rect 476 1392 483 1394
rect 476 1391 477 1392
rect 471 1390 477 1391
rect 482 1391 483 1392
rect 487 1391 488 1395
rect 535 1395 541 1396
rect 535 1394 536 1395
rect 528 1392 536 1394
rect 482 1390 488 1391
rect 518 1391 524 1392
rect 454 1386 460 1387
rect 518 1387 519 1391
rect 523 1387 524 1391
rect 518 1386 524 1387
rect 528 1382 530 1392
rect 535 1391 536 1392
rect 540 1391 541 1395
rect 599 1395 605 1396
rect 599 1394 600 1395
rect 592 1392 600 1394
rect 535 1390 541 1391
rect 582 1391 588 1392
rect 582 1387 583 1391
rect 587 1387 588 1391
rect 582 1386 588 1387
rect 592 1382 594 1392
rect 599 1391 600 1392
rect 604 1391 605 1395
rect 663 1395 669 1396
rect 663 1394 664 1395
rect 656 1392 664 1394
rect 599 1390 605 1391
rect 646 1391 652 1392
rect 646 1387 647 1391
rect 651 1387 652 1391
rect 646 1386 652 1387
rect 656 1382 658 1392
rect 663 1391 664 1392
rect 668 1391 669 1395
rect 727 1395 733 1396
rect 727 1394 728 1395
rect 720 1392 728 1394
rect 663 1390 669 1391
rect 710 1391 716 1392
rect 710 1387 711 1391
rect 715 1387 716 1391
rect 710 1386 716 1387
rect 720 1382 722 1392
rect 727 1391 728 1392
rect 732 1391 733 1395
rect 791 1395 797 1396
rect 791 1394 792 1395
rect 784 1392 792 1394
rect 727 1390 733 1391
rect 774 1391 780 1392
rect 774 1387 775 1391
rect 779 1387 780 1391
rect 774 1386 780 1387
rect 784 1382 786 1392
rect 791 1391 792 1392
rect 796 1391 797 1395
rect 855 1395 861 1396
rect 855 1394 856 1395
rect 848 1392 856 1394
rect 791 1390 797 1391
rect 838 1391 844 1392
rect 838 1387 839 1391
rect 843 1387 844 1391
rect 838 1386 844 1387
rect 848 1382 850 1392
rect 855 1391 856 1392
rect 860 1391 861 1395
rect 910 1395 917 1396
rect 855 1390 861 1391
rect 894 1391 900 1392
rect 894 1387 895 1391
rect 899 1387 900 1391
rect 910 1391 911 1395
rect 916 1391 917 1395
rect 967 1395 973 1396
rect 967 1394 968 1395
rect 960 1392 968 1394
rect 910 1390 917 1391
rect 950 1391 956 1392
rect 894 1386 900 1387
rect 950 1387 951 1391
rect 955 1387 956 1391
rect 950 1386 956 1387
rect 960 1382 962 1392
rect 967 1391 968 1392
rect 972 1391 973 1395
rect 1015 1395 1021 1396
rect 1015 1394 1016 1395
rect 1008 1392 1016 1394
rect 967 1390 973 1391
rect 998 1391 1004 1392
rect 998 1387 999 1391
rect 1003 1387 1004 1391
rect 998 1386 1004 1387
rect 1008 1382 1010 1392
rect 1015 1391 1016 1392
rect 1020 1391 1021 1395
rect 1071 1395 1077 1396
rect 1071 1394 1072 1395
rect 1064 1392 1072 1394
rect 1015 1390 1021 1391
rect 1054 1391 1060 1392
rect 1054 1387 1055 1391
rect 1059 1387 1060 1391
rect 1054 1386 1060 1387
rect 1064 1382 1066 1392
rect 1071 1391 1072 1392
rect 1076 1391 1077 1395
rect 1102 1395 1103 1399
rect 1107 1395 1108 1399
rect 1263 1399 1269 1400
rect 1102 1394 1108 1395
rect 1127 1395 1133 1396
rect 1127 1394 1128 1395
rect 1120 1392 1128 1394
rect 1071 1390 1077 1391
rect 1110 1391 1116 1392
rect 1110 1387 1111 1391
rect 1115 1387 1116 1391
rect 1110 1386 1116 1387
rect 1120 1382 1122 1392
rect 1127 1391 1128 1392
rect 1132 1391 1133 1395
rect 1186 1395 1197 1396
rect 1127 1390 1133 1391
rect 1174 1391 1180 1392
rect 1174 1387 1175 1391
rect 1179 1387 1180 1391
rect 1186 1391 1187 1395
rect 1191 1391 1192 1395
rect 1196 1391 1197 1395
rect 1255 1395 1261 1396
rect 1255 1394 1256 1395
rect 1248 1392 1256 1394
rect 1186 1390 1197 1391
rect 1238 1391 1244 1392
rect 1174 1386 1180 1387
rect 1238 1387 1239 1391
rect 1243 1387 1244 1391
rect 1238 1386 1244 1387
rect 1248 1382 1250 1392
rect 1255 1391 1256 1392
rect 1260 1391 1261 1395
rect 1263 1395 1264 1399
rect 1268 1398 1269 1399
rect 1268 1396 1306 1398
rect 1268 1395 1269 1396
rect 1263 1394 1269 1395
rect 1304 1394 1306 1396
rect 1311 1395 1317 1396
rect 1311 1394 1312 1395
rect 1304 1392 1312 1394
rect 1255 1390 1261 1391
rect 1294 1391 1300 1392
rect 1294 1387 1295 1391
rect 1299 1387 1300 1391
rect 1311 1391 1312 1392
rect 1316 1391 1317 1395
rect 1367 1395 1373 1396
rect 1311 1390 1317 1391
rect 1350 1391 1356 1392
rect 1294 1386 1300 1387
rect 1350 1387 1351 1391
rect 1355 1387 1356 1391
rect 1367 1391 1368 1395
rect 1372 1394 1373 1395
rect 1406 1395 1412 1396
rect 1406 1394 1407 1395
rect 1372 1392 1407 1394
rect 1372 1391 1373 1392
rect 1367 1390 1373 1391
rect 1406 1391 1407 1392
rect 1411 1391 1412 1395
rect 1431 1395 1437 1396
rect 1431 1394 1432 1395
rect 1424 1392 1432 1394
rect 1406 1390 1412 1391
rect 1414 1391 1420 1392
rect 1350 1386 1356 1387
rect 1414 1387 1415 1391
rect 1419 1387 1420 1391
rect 1414 1386 1420 1387
rect 1424 1382 1426 1392
rect 1431 1391 1432 1392
rect 1436 1391 1437 1395
rect 1494 1395 1501 1396
rect 1431 1390 1437 1391
rect 1478 1391 1484 1392
rect 1478 1387 1479 1391
rect 1483 1387 1484 1391
rect 1494 1391 1495 1395
rect 1500 1391 1501 1395
rect 1559 1395 1565 1396
rect 1559 1394 1560 1395
rect 1552 1392 1560 1394
rect 1494 1390 1501 1391
rect 1542 1391 1548 1392
rect 1478 1386 1484 1387
rect 1542 1387 1543 1391
rect 1547 1387 1548 1391
rect 1542 1386 1548 1387
rect 1552 1382 1554 1392
rect 1559 1391 1560 1392
rect 1564 1391 1565 1395
rect 1559 1390 1565 1391
rect 1582 1392 1588 1393
rect 1582 1388 1583 1392
rect 1587 1388 1588 1392
rect 1582 1387 1588 1388
rect 168 1380 186 1382
rect 313 1380 330 1382
rect 376 1380 411 1382
rect 504 1380 530 1382
rect 568 1380 594 1382
rect 633 1380 658 1382
rect 696 1380 722 1382
rect 760 1380 786 1382
rect 824 1380 850 1382
rect 913 1380 962 1382
rect 969 1380 1010 1382
rect 1044 1380 1066 1382
rect 1099 1380 1122 1382
rect 1224 1380 1250 1382
rect 1400 1380 1426 1382
rect 1497 1380 1554 1382
rect 150 1379 157 1380
rect 110 1375 116 1376
rect 110 1371 111 1375
rect 115 1371 116 1375
rect 150 1375 151 1379
rect 156 1375 157 1379
rect 184 1378 186 1380
rect 191 1379 197 1380
rect 191 1378 192 1379
rect 184 1376 192 1378
rect 150 1374 157 1375
rect 191 1375 192 1376
rect 196 1375 197 1379
rect 191 1374 197 1375
rect 262 1379 269 1380
rect 262 1375 263 1379
rect 268 1375 269 1379
rect 328 1378 330 1380
rect 335 1379 341 1380
rect 335 1378 336 1379
rect 328 1376 336 1378
rect 262 1374 269 1375
rect 335 1375 336 1376
rect 340 1375 341 1379
rect 335 1374 341 1375
rect 407 1379 413 1380
rect 407 1375 408 1379
rect 412 1375 413 1379
rect 407 1374 413 1375
rect 471 1379 477 1380
rect 471 1375 472 1379
rect 476 1378 477 1379
rect 504 1378 506 1380
rect 476 1376 506 1378
rect 535 1379 541 1380
rect 476 1375 477 1376
rect 471 1374 477 1375
rect 535 1375 536 1379
rect 540 1378 541 1379
rect 568 1378 570 1380
rect 540 1376 570 1378
rect 599 1379 605 1380
rect 540 1375 541 1376
rect 535 1374 541 1375
rect 599 1375 600 1379
rect 604 1378 605 1379
rect 633 1378 635 1380
rect 604 1376 635 1378
rect 663 1379 669 1380
rect 604 1375 605 1376
rect 599 1374 605 1375
rect 663 1375 664 1379
rect 668 1378 669 1379
rect 696 1378 698 1380
rect 668 1376 698 1378
rect 727 1379 733 1380
rect 668 1375 669 1376
rect 663 1374 669 1375
rect 727 1375 728 1379
rect 732 1378 733 1379
rect 760 1378 762 1380
rect 732 1376 762 1378
rect 791 1379 797 1380
rect 732 1375 733 1376
rect 727 1374 733 1375
rect 791 1375 792 1379
rect 796 1378 797 1379
rect 824 1378 826 1380
rect 796 1376 826 1378
rect 854 1379 861 1380
rect 796 1375 797 1376
rect 791 1374 797 1375
rect 854 1375 855 1379
rect 860 1375 861 1379
rect 854 1374 861 1375
rect 911 1379 917 1380
rect 911 1375 912 1379
rect 916 1375 917 1379
rect 911 1374 917 1375
rect 967 1379 973 1380
rect 967 1375 968 1379
rect 972 1375 973 1379
rect 967 1374 973 1375
rect 1015 1379 1021 1380
rect 1015 1375 1016 1379
rect 1020 1378 1021 1379
rect 1044 1378 1046 1380
rect 1020 1376 1046 1378
rect 1071 1379 1077 1380
rect 1020 1375 1021 1376
rect 1015 1374 1021 1375
rect 1071 1375 1072 1379
rect 1076 1378 1077 1379
rect 1099 1378 1101 1380
rect 1076 1376 1101 1378
rect 1126 1379 1133 1380
rect 1076 1375 1077 1376
rect 1071 1374 1077 1375
rect 1126 1375 1127 1379
rect 1132 1375 1133 1379
rect 1126 1374 1133 1375
rect 1191 1379 1197 1380
rect 1191 1375 1192 1379
rect 1196 1378 1197 1379
rect 1224 1378 1226 1380
rect 1196 1376 1226 1378
rect 1255 1379 1261 1380
rect 1196 1375 1197 1376
rect 1191 1374 1197 1375
rect 1255 1375 1256 1379
rect 1260 1378 1261 1379
rect 1263 1379 1269 1380
rect 1263 1378 1264 1379
rect 1260 1376 1264 1378
rect 1260 1375 1261 1376
rect 1255 1374 1261 1375
rect 1263 1375 1264 1376
rect 1268 1375 1269 1379
rect 1263 1374 1269 1375
rect 1306 1379 1317 1380
rect 1306 1375 1307 1379
rect 1311 1375 1312 1379
rect 1316 1375 1317 1379
rect 1306 1374 1317 1375
rect 1367 1379 1373 1380
rect 1367 1375 1368 1379
rect 1372 1378 1373 1379
rect 1400 1378 1402 1380
rect 1372 1376 1402 1378
rect 1431 1379 1437 1380
rect 1372 1375 1373 1376
rect 1367 1374 1373 1375
rect 1431 1375 1432 1379
rect 1436 1378 1437 1379
rect 1462 1379 1468 1380
rect 1462 1378 1463 1379
rect 1436 1376 1463 1378
rect 1436 1375 1437 1376
rect 1431 1374 1437 1375
rect 1462 1375 1463 1376
rect 1467 1375 1468 1379
rect 1462 1374 1468 1375
rect 1495 1379 1501 1380
rect 1495 1375 1496 1379
rect 1500 1375 1501 1379
rect 1495 1374 1501 1375
rect 1559 1379 1565 1380
rect 1559 1375 1560 1379
rect 1564 1375 1565 1379
rect 1559 1374 1565 1375
rect 1582 1375 1588 1376
rect 110 1370 116 1371
rect 134 1373 140 1374
rect 134 1369 135 1373
rect 139 1369 140 1373
rect 134 1368 140 1369
rect 174 1373 180 1374
rect 174 1369 175 1373
rect 179 1369 180 1373
rect 174 1368 180 1369
rect 246 1373 252 1374
rect 246 1369 247 1373
rect 251 1369 252 1373
rect 246 1368 252 1369
rect 318 1373 324 1374
rect 318 1369 319 1373
rect 323 1369 324 1373
rect 318 1368 324 1369
rect 390 1373 396 1374
rect 390 1369 391 1373
rect 395 1369 396 1373
rect 390 1368 396 1369
rect 454 1373 460 1374
rect 454 1369 455 1373
rect 459 1369 460 1373
rect 454 1368 460 1369
rect 518 1373 524 1374
rect 518 1369 519 1373
rect 523 1369 524 1373
rect 518 1368 524 1369
rect 582 1373 588 1374
rect 582 1369 583 1373
rect 587 1369 588 1373
rect 582 1368 588 1369
rect 646 1373 652 1374
rect 646 1369 647 1373
rect 651 1369 652 1373
rect 646 1368 652 1369
rect 710 1373 716 1374
rect 710 1369 711 1373
rect 715 1369 716 1373
rect 710 1368 716 1369
rect 774 1373 780 1374
rect 774 1369 775 1373
rect 779 1369 780 1373
rect 774 1368 780 1369
rect 838 1373 844 1374
rect 838 1369 839 1373
rect 843 1369 844 1373
rect 838 1368 844 1369
rect 894 1373 900 1374
rect 894 1369 895 1373
rect 899 1369 900 1373
rect 894 1368 900 1369
rect 950 1373 956 1374
rect 950 1369 951 1373
rect 955 1369 956 1373
rect 950 1368 956 1369
rect 998 1373 1004 1374
rect 998 1369 999 1373
rect 1003 1369 1004 1373
rect 998 1368 1004 1369
rect 1054 1373 1060 1374
rect 1054 1369 1055 1373
rect 1059 1369 1060 1373
rect 1054 1368 1060 1369
rect 1110 1373 1116 1374
rect 1110 1369 1111 1373
rect 1115 1369 1116 1373
rect 1110 1368 1116 1369
rect 1174 1373 1180 1374
rect 1174 1369 1175 1373
rect 1179 1369 1180 1373
rect 1174 1368 1180 1369
rect 1238 1373 1244 1374
rect 1238 1369 1239 1373
rect 1243 1369 1244 1373
rect 1238 1368 1244 1369
rect 1294 1373 1300 1374
rect 1294 1369 1295 1373
rect 1299 1369 1300 1373
rect 1294 1368 1300 1369
rect 1350 1373 1356 1374
rect 1350 1369 1351 1373
rect 1355 1369 1356 1373
rect 1350 1368 1356 1369
rect 1414 1373 1420 1374
rect 1414 1369 1415 1373
rect 1419 1369 1420 1373
rect 1414 1368 1420 1369
rect 1478 1373 1484 1374
rect 1478 1369 1479 1373
rect 1483 1369 1484 1373
rect 1478 1368 1484 1369
rect 1542 1373 1548 1374
rect 1542 1369 1543 1373
rect 1547 1369 1548 1373
rect 1542 1368 1548 1369
rect 446 1367 452 1368
rect 446 1363 447 1367
rect 451 1366 452 1367
rect 1087 1367 1093 1368
rect 451 1364 606 1366
rect 451 1363 452 1364
rect 446 1362 452 1363
rect 134 1359 140 1360
rect 110 1357 116 1358
rect 110 1353 111 1357
rect 115 1353 116 1357
rect 134 1355 135 1359
rect 139 1355 140 1359
rect 134 1354 140 1355
rect 166 1359 172 1360
rect 166 1355 167 1359
rect 171 1355 172 1359
rect 166 1354 172 1355
rect 214 1359 220 1360
rect 214 1355 215 1359
rect 219 1355 220 1359
rect 214 1354 220 1355
rect 302 1359 308 1360
rect 302 1355 303 1359
rect 307 1355 308 1359
rect 302 1354 308 1355
rect 414 1359 420 1360
rect 414 1355 415 1359
rect 419 1355 420 1359
rect 414 1354 420 1355
rect 526 1359 532 1360
rect 526 1355 527 1359
rect 531 1355 532 1359
rect 526 1354 532 1355
rect 110 1352 116 1353
rect 151 1351 157 1352
rect 151 1347 152 1351
rect 156 1350 157 1351
rect 183 1351 189 1352
rect 156 1348 178 1350
rect 156 1347 157 1348
rect 151 1346 157 1347
rect 134 1341 140 1342
rect 110 1340 116 1341
rect 110 1336 111 1340
rect 115 1336 116 1340
rect 134 1337 135 1341
rect 139 1337 140 1341
rect 134 1336 140 1337
rect 166 1341 172 1342
rect 166 1337 167 1341
rect 171 1337 172 1341
rect 166 1336 172 1337
rect 110 1335 116 1336
rect 150 1335 157 1336
rect 150 1331 151 1335
rect 156 1331 157 1335
rect 176 1334 178 1348
rect 183 1347 184 1351
rect 188 1347 189 1351
rect 183 1346 189 1347
rect 202 1351 208 1352
rect 202 1347 203 1351
rect 207 1350 208 1351
rect 231 1351 237 1352
rect 231 1350 232 1351
rect 207 1348 232 1350
rect 207 1347 208 1348
rect 202 1346 208 1347
rect 231 1347 232 1348
rect 236 1347 237 1351
rect 231 1346 237 1347
rect 319 1351 325 1352
rect 319 1347 320 1351
rect 324 1350 325 1351
rect 431 1351 437 1352
rect 324 1348 378 1350
rect 324 1347 325 1348
rect 319 1346 325 1347
rect 185 1342 187 1346
rect 185 1340 210 1342
rect 183 1335 189 1336
rect 183 1334 184 1335
rect 176 1332 184 1334
rect 150 1330 157 1331
rect 183 1331 184 1332
rect 188 1331 189 1335
rect 208 1334 210 1340
rect 214 1341 220 1342
rect 214 1337 215 1341
rect 219 1337 220 1341
rect 214 1336 220 1337
rect 302 1341 308 1342
rect 302 1337 303 1341
rect 307 1337 308 1341
rect 302 1336 308 1337
rect 231 1335 237 1336
rect 231 1334 232 1335
rect 208 1332 232 1334
rect 183 1330 189 1331
rect 231 1331 232 1332
rect 236 1331 237 1335
rect 231 1330 237 1331
rect 266 1335 272 1336
rect 266 1331 267 1335
rect 271 1334 272 1335
rect 319 1335 325 1336
rect 319 1334 320 1335
rect 271 1332 320 1334
rect 271 1331 272 1332
rect 266 1330 272 1331
rect 319 1331 320 1332
rect 324 1331 325 1335
rect 376 1334 378 1348
rect 431 1347 432 1351
rect 436 1350 437 1351
rect 543 1351 549 1352
rect 436 1348 490 1350
rect 436 1347 437 1348
rect 431 1346 437 1347
rect 414 1341 420 1342
rect 414 1337 415 1341
rect 419 1337 420 1341
rect 414 1336 420 1337
rect 431 1335 437 1336
rect 431 1334 432 1335
rect 376 1332 432 1334
rect 319 1330 325 1331
rect 431 1331 432 1332
rect 436 1331 437 1335
rect 488 1334 490 1348
rect 543 1347 544 1351
rect 548 1350 549 1351
rect 604 1350 606 1364
rect 1087 1363 1088 1367
rect 1092 1366 1093 1367
rect 1406 1367 1412 1368
rect 1092 1364 1242 1366
rect 1092 1363 1093 1364
rect 1087 1362 1093 1363
rect 638 1359 644 1360
rect 638 1355 639 1359
rect 643 1355 644 1359
rect 638 1354 644 1355
rect 750 1359 756 1360
rect 750 1355 751 1359
rect 755 1355 756 1359
rect 750 1354 756 1355
rect 862 1359 868 1360
rect 862 1355 863 1359
rect 867 1355 868 1359
rect 862 1354 868 1355
rect 966 1359 972 1360
rect 966 1355 967 1359
rect 971 1355 972 1359
rect 966 1354 972 1355
rect 1062 1359 1068 1360
rect 1062 1355 1063 1359
rect 1067 1355 1068 1359
rect 1126 1359 1132 1360
rect 1126 1358 1127 1359
rect 1062 1354 1068 1355
rect 1072 1356 1127 1358
rect 655 1351 661 1352
rect 655 1350 656 1351
rect 548 1348 602 1350
rect 604 1348 656 1350
rect 548 1347 549 1348
rect 543 1346 549 1347
rect 526 1341 532 1342
rect 526 1337 527 1341
rect 531 1337 532 1341
rect 526 1336 532 1337
rect 543 1335 549 1336
rect 543 1334 544 1335
rect 488 1332 544 1334
rect 431 1330 437 1331
rect 543 1331 544 1332
rect 548 1331 549 1335
rect 600 1334 602 1348
rect 655 1347 656 1348
rect 660 1347 661 1351
rect 655 1346 661 1347
rect 767 1351 773 1352
rect 767 1347 768 1351
rect 772 1350 773 1351
rect 879 1351 885 1352
rect 772 1348 826 1350
rect 772 1347 773 1348
rect 767 1346 773 1347
rect 638 1341 644 1342
rect 638 1337 639 1341
rect 643 1337 644 1341
rect 638 1336 644 1337
rect 750 1341 756 1342
rect 750 1337 751 1341
rect 755 1337 756 1341
rect 750 1336 756 1337
rect 655 1335 661 1336
rect 655 1334 656 1335
rect 600 1332 656 1334
rect 543 1330 549 1331
rect 655 1331 656 1332
rect 660 1331 661 1335
rect 655 1330 661 1331
rect 767 1335 773 1336
rect 767 1331 768 1335
rect 772 1334 773 1335
rect 824 1334 826 1348
rect 879 1347 880 1351
rect 884 1350 885 1351
rect 902 1351 908 1352
rect 902 1350 903 1351
rect 884 1348 903 1350
rect 884 1347 885 1348
rect 879 1346 885 1347
rect 902 1347 903 1348
rect 907 1347 908 1351
rect 902 1346 908 1347
rect 910 1351 916 1352
rect 910 1347 911 1351
rect 915 1350 916 1351
rect 983 1351 989 1352
rect 983 1350 984 1351
rect 915 1348 984 1350
rect 915 1347 916 1348
rect 910 1346 916 1347
rect 983 1347 984 1348
rect 988 1347 989 1351
rect 983 1346 989 1347
rect 862 1341 868 1342
rect 862 1337 863 1341
rect 867 1337 868 1341
rect 862 1336 868 1337
rect 966 1341 972 1342
rect 966 1337 967 1341
rect 971 1337 972 1341
rect 966 1336 972 1337
rect 1062 1341 1068 1342
rect 1062 1337 1063 1341
rect 1067 1337 1068 1341
rect 1062 1336 1068 1337
rect 879 1335 885 1336
rect 879 1334 880 1335
rect 772 1332 822 1334
rect 824 1332 880 1334
rect 772 1331 773 1332
rect 767 1330 773 1331
rect 820 1330 822 1332
rect 879 1331 880 1332
rect 884 1331 885 1335
rect 983 1335 989 1336
rect 879 1330 885 1331
rect 910 1331 916 1332
rect 910 1330 911 1331
rect 820 1328 866 1330
rect 864 1326 866 1328
rect 888 1328 911 1330
rect 888 1326 890 1328
rect 910 1327 911 1328
rect 915 1327 916 1331
rect 983 1331 984 1335
rect 988 1334 989 1335
rect 1072 1334 1074 1356
rect 1126 1355 1127 1356
rect 1131 1355 1132 1359
rect 1126 1354 1132 1355
rect 1150 1359 1156 1360
rect 1150 1355 1151 1359
rect 1155 1355 1156 1359
rect 1150 1354 1156 1355
rect 1230 1359 1236 1360
rect 1230 1355 1231 1359
rect 1235 1355 1236 1359
rect 1230 1354 1236 1355
rect 1079 1351 1085 1352
rect 1079 1347 1080 1351
rect 1084 1350 1085 1351
rect 1167 1351 1173 1352
rect 1084 1348 1101 1350
rect 1084 1347 1085 1348
rect 1079 1346 1085 1347
rect 988 1332 1074 1334
rect 1079 1335 1085 1336
rect 988 1331 989 1332
rect 983 1330 989 1331
rect 1079 1331 1080 1335
rect 1084 1334 1085 1335
rect 1087 1335 1093 1336
rect 1087 1334 1088 1335
rect 1084 1332 1088 1334
rect 1084 1331 1085 1332
rect 1079 1330 1085 1331
rect 1087 1331 1088 1332
rect 1092 1331 1093 1335
rect 1099 1334 1101 1348
rect 1167 1347 1168 1351
rect 1172 1350 1173 1351
rect 1186 1351 1192 1352
rect 1186 1350 1187 1351
rect 1172 1348 1187 1350
rect 1172 1347 1173 1348
rect 1167 1346 1173 1347
rect 1186 1347 1187 1348
rect 1191 1347 1192 1351
rect 1240 1350 1242 1364
rect 1406 1363 1407 1367
rect 1411 1366 1412 1367
rect 1561 1366 1563 1374
rect 1582 1371 1583 1375
rect 1587 1371 1588 1375
rect 1582 1370 1588 1371
rect 1411 1364 1563 1366
rect 1411 1363 1412 1364
rect 1406 1362 1412 1363
rect 1310 1359 1316 1360
rect 1310 1355 1311 1359
rect 1315 1355 1316 1359
rect 1310 1354 1316 1355
rect 1382 1359 1388 1360
rect 1382 1355 1383 1359
rect 1387 1355 1388 1359
rect 1382 1354 1388 1355
rect 1454 1359 1460 1360
rect 1454 1355 1455 1359
rect 1459 1355 1460 1359
rect 1534 1359 1540 1360
rect 1454 1354 1460 1355
rect 1464 1356 1518 1358
rect 1247 1351 1253 1352
rect 1247 1350 1248 1351
rect 1240 1348 1248 1350
rect 1186 1346 1192 1347
rect 1247 1347 1248 1348
rect 1252 1347 1253 1351
rect 1247 1346 1253 1347
rect 1327 1351 1333 1352
rect 1327 1347 1328 1351
rect 1332 1350 1333 1351
rect 1399 1351 1405 1352
rect 1332 1348 1366 1350
rect 1332 1347 1333 1348
rect 1327 1346 1333 1347
rect 1150 1341 1156 1342
rect 1150 1337 1151 1341
rect 1155 1337 1156 1341
rect 1150 1336 1156 1337
rect 1230 1341 1236 1342
rect 1230 1337 1231 1341
rect 1235 1337 1236 1341
rect 1230 1336 1236 1337
rect 1310 1341 1316 1342
rect 1310 1337 1311 1341
rect 1315 1337 1316 1341
rect 1310 1336 1316 1337
rect 1354 1339 1360 1340
rect 1167 1335 1173 1336
rect 1167 1334 1168 1335
rect 1099 1332 1168 1334
rect 1087 1330 1093 1331
rect 1167 1331 1168 1332
rect 1172 1331 1173 1335
rect 1167 1330 1173 1331
rect 1238 1335 1244 1336
rect 1238 1331 1239 1335
rect 1243 1334 1244 1335
rect 1247 1335 1253 1336
rect 1247 1334 1248 1335
rect 1243 1332 1248 1334
rect 1243 1331 1244 1332
rect 1238 1330 1244 1331
rect 1247 1331 1248 1332
rect 1252 1331 1253 1335
rect 1247 1330 1253 1331
rect 1327 1335 1333 1336
rect 1327 1331 1328 1335
rect 1332 1334 1333 1335
rect 1354 1335 1355 1339
rect 1359 1335 1360 1339
rect 1354 1334 1360 1335
rect 1364 1334 1366 1348
rect 1399 1347 1400 1351
rect 1404 1350 1405 1351
rect 1438 1351 1444 1352
rect 1438 1350 1439 1351
rect 1404 1348 1439 1350
rect 1404 1347 1405 1348
rect 1399 1346 1405 1347
rect 1438 1347 1439 1348
rect 1443 1347 1444 1351
rect 1438 1346 1444 1347
rect 1446 1351 1452 1352
rect 1446 1347 1447 1351
rect 1451 1350 1452 1351
rect 1464 1350 1466 1356
rect 1451 1348 1466 1350
rect 1471 1351 1477 1352
rect 1451 1347 1452 1348
rect 1446 1346 1452 1347
rect 1471 1347 1472 1351
rect 1476 1350 1477 1351
rect 1516 1350 1518 1356
rect 1534 1355 1535 1359
rect 1539 1355 1540 1359
rect 1534 1354 1540 1355
rect 1582 1357 1588 1358
rect 1582 1353 1583 1357
rect 1587 1353 1588 1357
rect 1582 1352 1588 1353
rect 1551 1351 1557 1352
rect 1551 1350 1552 1351
rect 1476 1348 1514 1350
rect 1516 1348 1552 1350
rect 1476 1347 1477 1348
rect 1471 1346 1477 1347
rect 1382 1341 1388 1342
rect 1382 1337 1383 1341
rect 1387 1337 1388 1341
rect 1382 1336 1388 1337
rect 1454 1341 1460 1342
rect 1454 1337 1455 1341
rect 1459 1337 1460 1341
rect 1454 1336 1460 1337
rect 1399 1335 1405 1336
rect 1399 1334 1400 1335
rect 1332 1332 1358 1334
rect 1364 1332 1400 1334
rect 1332 1331 1333 1332
rect 1327 1330 1333 1331
rect 1399 1331 1400 1332
rect 1404 1331 1405 1335
rect 1399 1330 1405 1331
rect 1462 1335 1468 1336
rect 1462 1331 1463 1335
rect 1467 1334 1468 1335
rect 1471 1335 1477 1336
rect 1471 1334 1472 1335
rect 1467 1332 1472 1334
rect 1467 1331 1468 1332
rect 1462 1330 1468 1331
rect 1471 1331 1472 1332
rect 1476 1331 1477 1335
rect 1512 1334 1514 1348
rect 1551 1347 1552 1348
rect 1556 1347 1557 1351
rect 1551 1346 1557 1347
rect 1534 1341 1540 1342
rect 1534 1337 1535 1341
rect 1539 1337 1540 1341
rect 1534 1336 1540 1337
rect 1582 1340 1588 1341
rect 1582 1336 1583 1340
rect 1587 1336 1588 1340
rect 1551 1335 1557 1336
rect 1582 1335 1588 1336
rect 1551 1334 1552 1335
rect 1512 1332 1552 1334
rect 1471 1330 1477 1331
rect 1551 1331 1552 1332
rect 1556 1331 1557 1335
rect 1551 1330 1557 1331
rect 1336 1328 1386 1330
rect 910 1326 916 1327
rect 1054 1327 1060 1328
rect 864 1324 890 1326
rect 151 1323 157 1324
rect 110 1320 116 1321
rect 110 1316 111 1320
rect 115 1316 116 1320
rect 110 1315 116 1316
rect 134 1319 140 1320
rect 134 1315 135 1319
rect 139 1315 140 1319
rect 151 1319 152 1323
rect 156 1319 157 1323
rect 199 1323 208 1324
rect 151 1318 157 1319
rect 182 1319 188 1320
rect 134 1314 140 1315
rect 153 1314 155 1318
rect 182 1315 183 1319
rect 187 1315 188 1319
rect 199 1319 200 1323
rect 207 1319 208 1323
rect 263 1323 269 1324
rect 199 1318 208 1319
rect 246 1319 252 1320
rect 182 1314 188 1315
rect 246 1315 247 1319
rect 251 1315 252 1319
rect 263 1319 264 1323
rect 268 1322 269 1323
rect 327 1323 333 1324
rect 268 1320 306 1322
rect 268 1319 269 1320
rect 263 1318 269 1319
rect 246 1314 252 1315
rect 153 1312 178 1314
rect 176 1310 178 1312
rect 304 1310 306 1320
rect 310 1319 316 1320
rect 310 1315 311 1319
rect 315 1315 316 1319
rect 327 1319 328 1323
rect 332 1322 333 1323
rect 391 1323 397 1324
rect 332 1320 370 1322
rect 332 1319 333 1320
rect 327 1318 333 1319
rect 310 1314 316 1315
rect 368 1310 370 1320
rect 374 1319 380 1320
rect 374 1315 375 1319
rect 379 1315 380 1319
rect 391 1319 392 1323
rect 396 1322 397 1323
rect 406 1323 412 1324
rect 406 1322 407 1323
rect 396 1320 407 1322
rect 396 1319 397 1320
rect 391 1318 397 1319
rect 406 1319 407 1320
rect 411 1319 412 1323
rect 455 1323 461 1324
rect 406 1318 412 1319
rect 438 1319 444 1320
rect 374 1314 380 1315
rect 438 1315 439 1319
rect 443 1315 444 1319
rect 455 1319 456 1323
rect 460 1322 461 1323
rect 478 1323 484 1324
rect 478 1322 479 1323
rect 460 1320 479 1322
rect 460 1319 461 1320
rect 455 1318 461 1319
rect 478 1319 479 1320
rect 483 1319 484 1323
rect 511 1323 517 1324
rect 511 1322 512 1323
rect 504 1320 512 1322
rect 478 1318 484 1319
rect 494 1319 500 1320
rect 438 1314 444 1315
rect 494 1315 495 1319
rect 499 1315 500 1319
rect 494 1314 500 1315
rect 504 1310 506 1320
rect 511 1319 512 1320
rect 516 1319 517 1323
rect 559 1323 565 1324
rect 559 1322 560 1323
rect 552 1320 560 1322
rect 511 1318 517 1319
rect 542 1319 548 1320
rect 542 1315 543 1319
rect 547 1315 548 1319
rect 542 1314 548 1315
rect 552 1310 554 1320
rect 559 1319 560 1320
rect 564 1319 565 1323
rect 607 1323 613 1324
rect 607 1322 608 1323
rect 600 1320 608 1322
rect 559 1318 565 1319
rect 590 1319 596 1320
rect 590 1315 591 1319
rect 595 1315 596 1319
rect 590 1314 596 1315
rect 600 1310 602 1320
rect 607 1319 608 1320
rect 612 1319 613 1323
rect 655 1323 661 1324
rect 655 1322 656 1323
rect 648 1320 656 1322
rect 607 1318 613 1319
rect 638 1319 644 1320
rect 638 1315 639 1319
rect 643 1315 644 1319
rect 638 1314 644 1315
rect 648 1310 650 1320
rect 655 1319 656 1320
rect 660 1319 661 1323
rect 703 1323 709 1324
rect 703 1322 704 1323
rect 696 1320 704 1322
rect 655 1318 661 1319
rect 686 1319 692 1320
rect 686 1315 687 1319
rect 691 1315 692 1319
rect 686 1314 692 1315
rect 696 1310 698 1320
rect 703 1319 704 1320
rect 708 1319 709 1323
rect 759 1323 765 1324
rect 759 1322 760 1323
rect 752 1320 760 1322
rect 703 1318 709 1319
rect 742 1319 748 1320
rect 742 1315 743 1319
rect 747 1315 748 1319
rect 742 1314 748 1315
rect 752 1310 754 1320
rect 759 1319 760 1320
rect 764 1319 765 1323
rect 807 1323 813 1324
rect 807 1322 808 1323
rect 800 1320 808 1322
rect 759 1318 765 1319
rect 790 1319 796 1320
rect 790 1315 791 1319
rect 795 1315 796 1319
rect 790 1314 796 1315
rect 800 1310 802 1320
rect 807 1319 808 1320
rect 812 1319 813 1323
rect 855 1323 861 1324
rect 855 1322 856 1323
rect 848 1320 856 1322
rect 807 1318 813 1319
rect 838 1319 844 1320
rect 838 1315 839 1319
rect 843 1315 844 1319
rect 838 1314 844 1315
rect 848 1310 850 1320
rect 855 1319 856 1320
rect 860 1319 861 1323
rect 902 1323 909 1324
rect 855 1318 861 1319
rect 886 1319 892 1320
rect 886 1315 887 1319
rect 891 1315 892 1319
rect 902 1319 903 1323
rect 908 1319 909 1323
rect 951 1323 957 1324
rect 951 1322 952 1323
rect 944 1320 952 1322
rect 902 1318 909 1319
rect 934 1319 940 1320
rect 886 1314 892 1315
rect 934 1315 935 1319
rect 939 1315 940 1319
rect 934 1314 940 1315
rect 944 1310 946 1320
rect 951 1319 952 1320
rect 956 1319 957 1323
rect 1007 1323 1013 1324
rect 1007 1322 1008 1323
rect 1000 1320 1008 1322
rect 951 1318 957 1319
rect 990 1319 996 1320
rect 990 1315 991 1319
rect 995 1315 996 1319
rect 990 1314 996 1315
rect 1000 1310 1002 1320
rect 1007 1319 1008 1320
rect 1012 1319 1013 1323
rect 1054 1323 1055 1327
rect 1059 1323 1060 1327
rect 1336 1326 1338 1328
rect 1320 1324 1338 1326
rect 1054 1322 1060 1323
rect 1063 1323 1069 1324
rect 1063 1322 1064 1323
rect 1056 1320 1064 1322
rect 1007 1318 1013 1319
rect 1046 1319 1052 1320
rect 1046 1315 1047 1319
rect 1051 1315 1052 1319
rect 1063 1319 1064 1320
rect 1068 1319 1069 1323
rect 1119 1323 1125 1324
rect 1119 1322 1120 1323
rect 1112 1320 1120 1322
rect 1063 1318 1069 1319
rect 1102 1319 1108 1320
rect 1046 1314 1052 1315
rect 1102 1315 1103 1319
rect 1107 1315 1108 1319
rect 1102 1314 1108 1315
rect 1112 1310 1114 1320
rect 1119 1319 1120 1320
rect 1124 1319 1125 1323
rect 1175 1323 1181 1324
rect 1175 1322 1176 1323
rect 1168 1320 1176 1322
rect 1119 1318 1125 1319
rect 1158 1319 1164 1320
rect 1158 1315 1159 1319
rect 1163 1315 1164 1319
rect 1158 1314 1164 1315
rect 1168 1310 1170 1320
rect 1175 1319 1176 1320
rect 1180 1319 1181 1323
rect 1231 1323 1237 1324
rect 1231 1322 1232 1323
rect 1224 1320 1232 1322
rect 1175 1318 1181 1319
rect 1214 1319 1220 1320
rect 1214 1315 1215 1319
rect 1219 1315 1220 1319
rect 1214 1314 1220 1315
rect 1224 1310 1226 1320
rect 1231 1319 1232 1320
rect 1236 1319 1237 1323
rect 1287 1323 1293 1324
rect 1231 1318 1237 1319
rect 1270 1319 1276 1320
rect 1270 1315 1271 1319
rect 1275 1315 1276 1319
rect 1287 1319 1288 1323
rect 1292 1322 1293 1323
rect 1320 1322 1322 1324
rect 1343 1323 1349 1324
rect 1343 1322 1344 1323
rect 1292 1320 1322 1322
rect 1336 1320 1344 1322
rect 1292 1319 1293 1320
rect 1287 1318 1293 1319
rect 1326 1319 1332 1320
rect 1270 1314 1276 1315
rect 1326 1315 1327 1319
rect 1331 1315 1332 1319
rect 1326 1314 1332 1315
rect 1336 1310 1338 1320
rect 1343 1319 1344 1320
rect 1348 1319 1349 1323
rect 1343 1318 1349 1319
rect 1374 1319 1380 1320
rect 1374 1315 1375 1319
rect 1379 1315 1380 1319
rect 1374 1314 1380 1315
rect 176 1308 194 1310
rect 304 1308 322 1310
rect 368 1308 386 1310
rect 484 1308 506 1310
rect 536 1308 554 1310
rect 584 1308 602 1310
rect 633 1308 650 1310
rect 680 1308 698 1310
rect 732 1308 754 1310
rect 784 1308 802 1310
rect 832 1308 850 1310
rect 928 1308 946 1310
rect 980 1308 1002 1310
rect 1099 1308 1114 1310
rect 1148 1308 1170 1310
rect 1204 1308 1226 1310
rect 1316 1308 1338 1310
rect 150 1307 157 1308
rect 110 1303 116 1304
rect 110 1299 111 1303
rect 115 1299 116 1303
rect 150 1303 151 1307
rect 156 1303 157 1307
rect 192 1306 194 1308
rect 199 1307 205 1308
rect 199 1306 200 1307
rect 192 1304 200 1306
rect 150 1302 157 1303
rect 199 1303 200 1304
rect 204 1303 205 1307
rect 199 1302 205 1303
rect 263 1307 272 1308
rect 263 1303 264 1307
rect 271 1303 272 1307
rect 320 1306 322 1308
rect 327 1307 333 1308
rect 327 1306 328 1307
rect 320 1304 328 1306
rect 263 1302 272 1303
rect 327 1303 328 1304
rect 332 1303 333 1307
rect 384 1306 386 1308
rect 391 1307 397 1308
rect 391 1306 392 1307
rect 384 1304 392 1306
rect 327 1302 333 1303
rect 391 1303 392 1304
rect 396 1303 397 1307
rect 391 1302 397 1303
rect 455 1307 461 1308
rect 455 1303 456 1307
rect 460 1306 461 1307
rect 484 1306 486 1308
rect 460 1304 486 1306
rect 511 1307 517 1308
rect 460 1303 461 1304
rect 455 1302 461 1303
rect 511 1303 512 1307
rect 516 1306 517 1307
rect 536 1306 538 1308
rect 516 1304 538 1306
rect 559 1307 565 1308
rect 516 1303 517 1304
rect 511 1302 517 1303
rect 559 1303 560 1307
rect 564 1306 565 1307
rect 584 1306 586 1308
rect 564 1304 586 1306
rect 607 1307 613 1308
rect 564 1303 565 1304
rect 559 1302 565 1303
rect 607 1303 608 1307
rect 612 1306 613 1307
rect 633 1306 635 1308
rect 612 1304 635 1306
rect 655 1307 661 1308
rect 612 1303 613 1304
rect 607 1302 613 1303
rect 655 1303 656 1307
rect 660 1306 661 1307
rect 680 1306 682 1308
rect 660 1304 682 1306
rect 703 1307 709 1308
rect 660 1303 661 1304
rect 655 1302 661 1303
rect 703 1303 704 1307
rect 708 1306 709 1307
rect 732 1306 734 1308
rect 708 1304 734 1306
rect 759 1307 765 1308
rect 708 1303 709 1304
rect 703 1302 709 1303
rect 759 1303 760 1307
rect 764 1306 765 1307
rect 784 1306 786 1308
rect 764 1304 786 1306
rect 807 1307 813 1308
rect 764 1303 765 1304
rect 759 1302 765 1303
rect 807 1303 808 1307
rect 812 1306 813 1307
rect 832 1306 834 1308
rect 812 1304 834 1306
rect 854 1307 861 1308
rect 812 1303 813 1304
rect 807 1302 813 1303
rect 854 1303 855 1307
rect 860 1303 861 1307
rect 854 1302 861 1303
rect 903 1307 909 1308
rect 903 1303 904 1307
rect 908 1306 909 1307
rect 928 1306 930 1308
rect 908 1304 930 1306
rect 951 1307 957 1308
rect 908 1303 909 1304
rect 903 1302 909 1303
rect 951 1303 952 1307
rect 956 1306 957 1307
rect 980 1306 982 1308
rect 956 1304 982 1306
rect 1006 1307 1013 1308
rect 956 1303 957 1304
rect 951 1302 957 1303
rect 1006 1303 1007 1307
rect 1012 1303 1013 1307
rect 1006 1302 1013 1303
rect 1063 1307 1069 1308
rect 1063 1303 1064 1307
rect 1068 1306 1069 1307
rect 1099 1306 1101 1308
rect 1068 1304 1101 1306
rect 1119 1307 1125 1308
rect 1068 1303 1069 1304
rect 1063 1302 1069 1303
rect 1119 1303 1120 1307
rect 1124 1306 1125 1307
rect 1148 1306 1150 1308
rect 1124 1304 1150 1306
rect 1175 1307 1181 1308
rect 1124 1303 1125 1304
rect 1119 1302 1125 1303
rect 1175 1303 1176 1307
rect 1180 1306 1181 1307
rect 1204 1306 1206 1308
rect 1180 1304 1206 1306
rect 1231 1307 1237 1308
rect 1180 1303 1181 1304
rect 1175 1302 1181 1303
rect 1231 1303 1232 1307
rect 1236 1303 1237 1307
rect 1231 1302 1237 1303
rect 1287 1307 1293 1308
rect 1287 1303 1288 1307
rect 1292 1306 1293 1307
rect 1316 1306 1318 1308
rect 1292 1304 1318 1306
rect 1343 1307 1349 1308
rect 1292 1303 1293 1304
rect 1287 1302 1293 1303
rect 1343 1303 1344 1307
rect 1348 1306 1349 1307
rect 1358 1307 1364 1308
rect 1358 1306 1359 1307
rect 1348 1304 1359 1306
rect 1348 1303 1349 1304
rect 1343 1302 1349 1303
rect 1358 1303 1359 1304
rect 1363 1303 1364 1307
rect 1384 1306 1386 1328
rect 1391 1323 1397 1324
rect 1391 1319 1392 1323
rect 1396 1322 1397 1323
rect 1414 1323 1420 1324
rect 1414 1322 1415 1323
rect 1396 1320 1415 1322
rect 1396 1319 1397 1320
rect 1391 1318 1397 1319
rect 1414 1319 1415 1320
rect 1419 1319 1420 1323
rect 1438 1323 1445 1324
rect 1414 1318 1420 1319
rect 1422 1319 1428 1320
rect 1422 1315 1423 1319
rect 1427 1315 1428 1319
rect 1438 1319 1439 1323
rect 1444 1319 1445 1323
rect 1487 1323 1493 1324
rect 1487 1322 1488 1323
rect 1480 1320 1488 1322
rect 1438 1318 1445 1319
rect 1470 1319 1476 1320
rect 1422 1314 1428 1315
rect 1470 1315 1471 1319
rect 1475 1315 1476 1319
rect 1470 1314 1476 1315
rect 1480 1310 1482 1320
rect 1487 1319 1488 1320
rect 1492 1319 1493 1323
rect 1543 1323 1549 1324
rect 1543 1322 1544 1323
rect 1536 1320 1544 1322
rect 1487 1318 1493 1319
rect 1526 1319 1532 1320
rect 1526 1315 1527 1319
rect 1531 1315 1532 1319
rect 1526 1314 1532 1315
rect 1536 1310 1538 1320
rect 1543 1319 1544 1320
rect 1548 1319 1549 1323
rect 1543 1318 1549 1319
rect 1582 1320 1588 1321
rect 1582 1316 1583 1320
rect 1587 1316 1588 1320
rect 1582 1315 1588 1316
rect 1464 1308 1482 1310
rect 1516 1308 1538 1310
rect 1391 1307 1397 1308
rect 1391 1306 1392 1307
rect 1384 1304 1392 1306
rect 1358 1302 1364 1303
rect 1391 1303 1392 1304
rect 1396 1303 1397 1307
rect 1391 1302 1397 1303
rect 1439 1307 1445 1308
rect 1439 1303 1440 1307
rect 1444 1306 1445 1307
rect 1464 1306 1466 1308
rect 1444 1304 1466 1306
rect 1487 1307 1493 1308
rect 1444 1303 1445 1304
rect 1439 1302 1445 1303
rect 1487 1303 1488 1307
rect 1492 1306 1493 1307
rect 1516 1306 1518 1308
rect 1543 1307 1549 1308
rect 1543 1306 1544 1307
rect 1492 1304 1518 1306
rect 1536 1304 1544 1306
rect 1492 1303 1493 1304
rect 1487 1302 1493 1303
rect 110 1298 116 1299
rect 134 1301 140 1302
rect 134 1297 135 1301
rect 139 1297 140 1301
rect 134 1296 140 1297
rect 182 1301 188 1302
rect 182 1297 183 1301
rect 187 1297 188 1301
rect 182 1296 188 1297
rect 246 1301 252 1302
rect 246 1297 247 1301
rect 251 1297 252 1301
rect 246 1296 252 1297
rect 310 1301 316 1302
rect 310 1297 311 1301
rect 315 1297 316 1301
rect 310 1296 316 1297
rect 374 1301 380 1302
rect 374 1297 375 1301
rect 379 1297 380 1301
rect 374 1296 380 1297
rect 438 1301 444 1302
rect 438 1297 439 1301
rect 443 1297 444 1301
rect 438 1296 444 1297
rect 494 1301 500 1302
rect 494 1297 495 1301
rect 499 1297 500 1301
rect 494 1296 500 1297
rect 542 1301 548 1302
rect 542 1297 543 1301
rect 547 1297 548 1301
rect 542 1296 548 1297
rect 590 1301 596 1302
rect 590 1297 591 1301
rect 595 1297 596 1301
rect 590 1296 596 1297
rect 638 1301 644 1302
rect 638 1297 639 1301
rect 643 1297 644 1301
rect 638 1296 644 1297
rect 686 1301 692 1302
rect 686 1297 687 1301
rect 691 1297 692 1301
rect 686 1296 692 1297
rect 742 1301 748 1302
rect 742 1297 743 1301
rect 747 1297 748 1301
rect 742 1296 748 1297
rect 790 1301 796 1302
rect 790 1297 791 1301
rect 795 1297 796 1301
rect 790 1296 796 1297
rect 838 1301 844 1302
rect 838 1297 839 1301
rect 843 1297 844 1301
rect 838 1296 844 1297
rect 886 1301 892 1302
rect 886 1297 887 1301
rect 891 1297 892 1301
rect 886 1296 892 1297
rect 934 1301 940 1302
rect 934 1297 935 1301
rect 939 1297 940 1301
rect 934 1296 940 1297
rect 990 1301 996 1302
rect 990 1297 991 1301
rect 995 1297 996 1301
rect 990 1296 996 1297
rect 1046 1301 1052 1302
rect 1046 1297 1047 1301
rect 1051 1297 1052 1301
rect 1046 1296 1052 1297
rect 1102 1301 1108 1302
rect 1102 1297 1103 1301
rect 1107 1297 1108 1301
rect 1102 1296 1108 1297
rect 1158 1301 1164 1302
rect 1158 1297 1159 1301
rect 1163 1297 1164 1301
rect 1158 1296 1164 1297
rect 1214 1301 1220 1302
rect 1214 1297 1215 1301
rect 1219 1297 1220 1301
rect 1214 1296 1220 1297
rect 1270 1301 1276 1302
rect 1270 1297 1271 1301
rect 1275 1297 1276 1301
rect 1270 1296 1276 1297
rect 1326 1301 1332 1302
rect 1326 1297 1327 1301
rect 1331 1297 1332 1301
rect 1326 1296 1332 1297
rect 1374 1301 1380 1302
rect 1374 1297 1375 1301
rect 1379 1297 1380 1301
rect 1374 1296 1380 1297
rect 1422 1301 1428 1302
rect 1422 1297 1423 1301
rect 1427 1297 1428 1301
rect 1422 1296 1428 1297
rect 1470 1301 1476 1302
rect 1470 1297 1471 1301
rect 1475 1297 1476 1301
rect 1470 1296 1476 1297
rect 1526 1301 1532 1302
rect 1526 1297 1527 1301
rect 1531 1297 1532 1301
rect 1526 1296 1532 1297
rect 695 1295 701 1296
rect 695 1291 696 1295
rect 700 1294 701 1295
rect 1018 1295 1024 1296
rect 700 1292 810 1294
rect 700 1291 701 1292
rect 695 1290 701 1291
rect 134 1287 140 1288
rect 110 1285 116 1286
rect 110 1281 111 1285
rect 115 1281 116 1285
rect 134 1283 135 1287
rect 139 1283 140 1287
rect 134 1282 140 1283
rect 190 1287 196 1288
rect 190 1283 191 1287
rect 195 1283 196 1287
rect 190 1282 196 1283
rect 254 1287 260 1288
rect 254 1283 255 1287
rect 259 1283 260 1287
rect 254 1282 260 1283
rect 326 1287 332 1288
rect 326 1283 327 1287
rect 331 1283 332 1287
rect 326 1282 332 1283
rect 390 1287 396 1288
rect 390 1283 391 1287
rect 395 1283 396 1287
rect 390 1282 396 1283
rect 462 1287 468 1288
rect 462 1283 463 1287
rect 467 1283 468 1287
rect 462 1282 468 1283
rect 534 1287 540 1288
rect 534 1283 535 1287
rect 539 1283 540 1287
rect 534 1282 540 1283
rect 598 1287 604 1288
rect 598 1283 599 1287
rect 603 1283 604 1287
rect 598 1282 604 1283
rect 662 1287 668 1288
rect 662 1283 663 1287
rect 667 1283 668 1287
rect 662 1282 668 1283
rect 726 1287 732 1288
rect 726 1283 727 1287
rect 731 1283 732 1287
rect 726 1282 732 1283
rect 790 1287 796 1288
rect 790 1283 791 1287
rect 795 1283 796 1287
rect 790 1282 796 1283
rect 110 1280 116 1281
rect 808 1280 810 1292
rect 1018 1291 1019 1295
rect 1023 1294 1024 1295
rect 1222 1295 1228 1296
rect 1023 1292 1101 1294
rect 1023 1291 1024 1292
rect 1018 1290 1024 1291
rect 854 1287 860 1288
rect 854 1283 855 1287
rect 859 1283 860 1287
rect 854 1282 860 1283
rect 926 1287 932 1288
rect 926 1283 927 1287
rect 931 1283 932 1287
rect 926 1282 932 1283
rect 998 1287 1004 1288
rect 998 1283 999 1287
rect 1003 1283 1004 1287
rect 998 1282 1004 1283
rect 1062 1287 1068 1288
rect 1062 1283 1063 1287
rect 1067 1283 1068 1287
rect 1062 1282 1068 1283
rect 1099 1282 1101 1292
rect 1222 1291 1223 1295
rect 1227 1294 1228 1295
rect 1414 1295 1420 1296
rect 1227 1292 1274 1294
rect 1227 1291 1228 1292
rect 1222 1290 1228 1291
rect 1126 1287 1132 1288
rect 1126 1283 1127 1287
rect 1131 1283 1132 1287
rect 1126 1282 1132 1283
rect 1190 1287 1196 1288
rect 1190 1283 1191 1287
rect 1195 1283 1196 1287
rect 1190 1282 1196 1283
rect 1246 1287 1252 1288
rect 1246 1283 1247 1287
rect 1251 1283 1252 1287
rect 1246 1282 1252 1283
rect 1099 1280 1122 1282
rect 151 1279 157 1280
rect 151 1275 152 1279
rect 156 1278 157 1279
rect 207 1279 213 1280
rect 156 1276 202 1278
rect 156 1275 157 1276
rect 151 1274 157 1275
rect 134 1269 140 1270
rect 110 1268 116 1269
rect 110 1264 111 1268
rect 115 1264 116 1268
rect 134 1265 135 1269
rect 139 1265 140 1269
rect 134 1264 140 1265
rect 190 1269 196 1270
rect 190 1265 191 1269
rect 195 1265 196 1269
rect 190 1264 196 1265
rect 110 1263 116 1264
rect 150 1263 157 1264
rect 150 1259 151 1263
rect 156 1259 157 1263
rect 200 1262 202 1276
rect 207 1275 208 1279
rect 212 1278 213 1279
rect 246 1279 252 1280
rect 246 1278 247 1279
rect 212 1276 247 1278
rect 212 1275 213 1276
rect 207 1274 213 1275
rect 246 1275 247 1276
rect 251 1275 252 1279
rect 246 1274 252 1275
rect 271 1279 277 1280
rect 271 1275 272 1279
rect 276 1278 277 1279
rect 343 1279 349 1280
rect 276 1276 314 1278
rect 276 1275 277 1276
rect 271 1274 277 1275
rect 254 1269 260 1270
rect 254 1265 255 1269
rect 259 1265 260 1269
rect 254 1264 260 1265
rect 207 1263 213 1264
rect 207 1262 208 1263
rect 200 1260 208 1262
rect 150 1258 157 1259
rect 207 1259 208 1260
rect 212 1259 213 1263
rect 207 1258 213 1259
rect 271 1263 277 1264
rect 271 1259 272 1263
rect 276 1262 277 1263
rect 302 1263 308 1264
rect 302 1262 303 1263
rect 276 1260 303 1262
rect 276 1259 277 1260
rect 271 1258 277 1259
rect 302 1259 303 1260
rect 307 1259 308 1263
rect 312 1262 314 1276
rect 343 1275 344 1279
rect 348 1278 349 1279
rect 406 1279 413 1280
rect 348 1276 402 1278
rect 348 1275 349 1276
rect 343 1274 349 1275
rect 326 1269 332 1270
rect 326 1265 327 1269
rect 331 1265 332 1269
rect 326 1264 332 1265
rect 390 1269 396 1270
rect 390 1265 391 1269
rect 395 1265 396 1269
rect 390 1264 396 1265
rect 343 1263 349 1264
rect 343 1262 344 1263
rect 312 1260 344 1262
rect 302 1258 308 1259
rect 343 1259 344 1260
rect 348 1259 349 1263
rect 400 1262 402 1276
rect 406 1275 407 1279
rect 412 1275 413 1279
rect 406 1274 413 1275
rect 478 1279 485 1280
rect 478 1275 479 1279
rect 484 1275 485 1279
rect 551 1279 557 1280
rect 551 1278 552 1279
rect 478 1274 485 1275
rect 520 1276 552 1278
rect 462 1269 468 1270
rect 462 1265 463 1269
rect 467 1265 468 1269
rect 462 1264 468 1265
rect 407 1263 413 1264
rect 407 1262 408 1263
rect 400 1260 408 1262
rect 343 1258 349 1259
rect 407 1259 408 1260
rect 412 1259 413 1263
rect 407 1258 413 1259
rect 479 1263 485 1264
rect 479 1259 480 1263
rect 484 1262 485 1263
rect 520 1262 522 1276
rect 551 1275 552 1276
rect 556 1275 557 1279
rect 615 1279 621 1280
rect 615 1278 616 1279
rect 551 1274 557 1275
rect 588 1276 616 1278
rect 534 1269 540 1270
rect 534 1265 535 1269
rect 539 1265 540 1269
rect 534 1264 540 1265
rect 484 1260 522 1262
rect 551 1263 557 1264
rect 484 1259 485 1260
rect 479 1258 485 1259
rect 551 1259 552 1263
rect 556 1262 557 1263
rect 588 1262 590 1276
rect 615 1275 616 1276
rect 620 1275 621 1279
rect 615 1274 621 1275
rect 679 1279 685 1280
rect 679 1275 680 1279
rect 684 1278 685 1279
rect 743 1279 749 1280
rect 684 1276 714 1278
rect 684 1275 685 1276
rect 679 1274 685 1275
rect 598 1269 604 1270
rect 598 1265 599 1269
rect 603 1265 604 1269
rect 598 1264 604 1265
rect 662 1269 668 1270
rect 662 1265 663 1269
rect 667 1265 668 1269
rect 662 1264 668 1265
rect 556 1260 590 1262
rect 615 1263 624 1264
rect 556 1259 557 1260
rect 551 1258 557 1259
rect 615 1259 616 1263
rect 623 1259 624 1263
rect 615 1258 624 1259
rect 679 1263 685 1264
rect 679 1259 680 1263
rect 684 1262 685 1263
rect 695 1263 701 1264
rect 695 1262 696 1263
rect 684 1260 696 1262
rect 684 1259 685 1260
rect 679 1258 685 1259
rect 695 1259 696 1260
rect 700 1259 701 1263
rect 712 1262 714 1276
rect 743 1275 744 1279
rect 748 1278 749 1279
rect 807 1279 813 1280
rect 748 1276 802 1278
rect 748 1275 749 1276
rect 743 1274 749 1275
rect 800 1270 802 1276
rect 807 1275 808 1279
rect 812 1275 813 1279
rect 807 1274 813 1275
rect 871 1279 880 1280
rect 871 1275 872 1279
rect 879 1275 880 1279
rect 943 1279 949 1280
rect 943 1278 944 1279
rect 871 1274 880 1275
rect 912 1276 944 1278
rect 814 1271 820 1272
rect 814 1270 815 1271
rect 726 1269 732 1270
rect 726 1265 727 1269
rect 731 1265 732 1269
rect 726 1264 732 1265
rect 790 1269 796 1270
rect 790 1265 791 1269
rect 795 1265 796 1269
rect 800 1268 815 1270
rect 814 1267 815 1268
rect 819 1267 820 1271
rect 814 1266 820 1267
rect 854 1269 860 1270
rect 790 1264 796 1265
rect 854 1265 855 1269
rect 859 1265 860 1269
rect 854 1264 860 1265
rect 743 1263 749 1264
rect 743 1262 744 1263
rect 712 1260 744 1262
rect 695 1258 701 1259
rect 743 1259 744 1260
rect 748 1259 749 1263
rect 743 1258 749 1259
rect 807 1263 813 1264
rect 807 1259 808 1263
rect 812 1262 813 1263
rect 846 1263 852 1264
rect 846 1262 847 1263
rect 812 1260 847 1262
rect 812 1259 813 1260
rect 807 1258 813 1259
rect 846 1259 847 1260
rect 851 1259 852 1263
rect 846 1258 852 1259
rect 871 1263 877 1264
rect 871 1259 872 1263
rect 876 1262 877 1263
rect 912 1262 914 1276
rect 943 1275 944 1276
rect 948 1275 949 1279
rect 943 1274 949 1275
rect 1015 1279 1021 1280
rect 1015 1275 1016 1279
rect 1020 1278 1021 1279
rect 1054 1279 1060 1280
rect 1054 1278 1055 1279
rect 1020 1276 1055 1278
rect 1020 1275 1021 1276
rect 1015 1274 1021 1275
rect 1054 1275 1055 1276
rect 1059 1275 1060 1279
rect 1054 1274 1060 1275
rect 1079 1279 1085 1280
rect 1079 1275 1080 1279
rect 1084 1278 1085 1279
rect 1120 1278 1122 1280
rect 1143 1279 1149 1280
rect 1143 1278 1144 1279
rect 1084 1276 1101 1278
rect 1120 1276 1144 1278
rect 1084 1275 1085 1276
rect 1079 1274 1085 1275
rect 926 1269 932 1270
rect 926 1265 927 1269
rect 931 1265 932 1269
rect 926 1264 932 1265
rect 998 1269 1004 1270
rect 998 1265 999 1269
rect 1003 1265 1004 1269
rect 998 1264 1004 1265
rect 1062 1269 1068 1270
rect 1062 1265 1063 1269
rect 1067 1265 1068 1269
rect 1062 1264 1068 1265
rect 876 1260 914 1262
rect 943 1263 949 1264
rect 876 1259 877 1260
rect 871 1258 877 1259
rect 943 1259 944 1263
rect 948 1262 949 1263
rect 1006 1263 1012 1264
rect 1006 1262 1007 1263
rect 948 1260 1007 1262
rect 948 1259 949 1260
rect 943 1258 949 1259
rect 1006 1259 1007 1260
rect 1011 1259 1012 1263
rect 1006 1258 1012 1259
rect 1015 1263 1024 1264
rect 1015 1259 1016 1263
rect 1023 1259 1024 1263
rect 1015 1258 1024 1259
rect 1074 1263 1085 1264
rect 1074 1259 1075 1263
rect 1079 1259 1080 1263
rect 1084 1259 1085 1263
rect 1099 1262 1101 1276
rect 1143 1275 1144 1276
rect 1148 1275 1149 1279
rect 1143 1274 1149 1275
rect 1207 1279 1213 1280
rect 1207 1275 1208 1279
rect 1212 1278 1213 1279
rect 1263 1279 1269 1280
rect 1212 1276 1258 1278
rect 1212 1275 1213 1276
rect 1207 1274 1213 1275
rect 1126 1269 1132 1270
rect 1126 1265 1127 1269
rect 1131 1265 1132 1269
rect 1126 1264 1132 1265
rect 1190 1269 1196 1270
rect 1190 1265 1191 1269
rect 1195 1265 1196 1269
rect 1190 1264 1196 1265
rect 1246 1269 1252 1270
rect 1246 1265 1247 1269
rect 1251 1265 1252 1269
rect 1246 1264 1252 1265
rect 1143 1263 1149 1264
rect 1143 1262 1144 1263
rect 1099 1260 1144 1262
rect 1074 1258 1085 1259
rect 1143 1259 1144 1260
rect 1148 1259 1149 1263
rect 1143 1258 1149 1259
rect 1207 1263 1213 1264
rect 1207 1259 1208 1263
rect 1212 1262 1213 1263
rect 1222 1263 1228 1264
rect 1222 1262 1223 1263
rect 1212 1260 1223 1262
rect 1212 1259 1213 1260
rect 1207 1258 1213 1259
rect 1222 1259 1223 1260
rect 1227 1259 1228 1263
rect 1256 1262 1258 1276
rect 1263 1275 1264 1279
rect 1268 1278 1269 1279
rect 1272 1278 1274 1292
rect 1414 1291 1415 1295
rect 1419 1294 1420 1295
rect 1536 1294 1538 1304
rect 1543 1303 1544 1304
rect 1548 1303 1549 1307
rect 1543 1302 1549 1303
rect 1582 1303 1588 1304
rect 1582 1299 1583 1303
rect 1587 1299 1588 1303
rect 1582 1298 1588 1299
rect 1419 1292 1538 1294
rect 1419 1291 1420 1292
rect 1414 1290 1420 1291
rect 1302 1287 1308 1288
rect 1302 1283 1303 1287
rect 1307 1283 1308 1287
rect 1302 1282 1308 1283
rect 1366 1287 1372 1288
rect 1366 1283 1367 1287
rect 1371 1283 1372 1287
rect 1430 1287 1436 1288
rect 1366 1282 1372 1283
rect 1376 1284 1422 1286
rect 1319 1279 1325 1280
rect 1319 1278 1320 1279
rect 1268 1275 1270 1278
rect 1272 1276 1320 1278
rect 1263 1274 1270 1275
rect 1319 1275 1320 1276
rect 1324 1275 1325 1279
rect 1376 1278 1378 1284
rect 1319 1274 1325 1275
rect 1352 1276 1378 1278
rect 1383 1279 1389 1280
rect 1268 1270 1270 1274
rect 1268 1268 1298 1270
rect 1263 1263 1269 1264
rect 1263 1262 1264 1263
rect 1256 1260 1264 1262
rect 1222 1258 1228 1259
rect 1263 1259 1264 1260
rect 1268 1259 1269 1263
rect 1263 1258 1269 1259
rect 334 1255 340 1256
rect 151 1251 157 1252
rect 110 1248 116 1249
rect 110 1244 111 1248
rect 115 1244 116 1248
rect 110 1243 116 1244
rect 134 1247 140 1248
rect 134 1243 135 1247
rect 139 1243 140 1247
rect 151 1247 152 1251
rect 156 1247 157 1251
rect 191 1251 197 1252
rect 151 1246 157 1247
rect 174 1247 180 1248
rect 134 1242 140 1243
rect 153 1242 155 1246
rect 174 1243 175 1247
rect 179 1243 180 1247
rect 191 1247 192 1251
rect 196 1250 197 1251
rect 246 1251 253 1252
rect 196 1248 222 1250
rect 196 1247 197 1248
rect 191 1246 197 1247
rect 174 1242 180 1243
rect 153 1240 170 1242
rect 168 1238 170 1240
rect 220 1238 222 1248
rect 230 1247 236 1248
rect 230 1243 231 1247
rect 235 1243 236 1247
rect 246 1247 247 1251
rect 252 1247 253 1251
rect 303 1251 309 1252
rect 246 1246 253 1247
rect 286 1247 292 1248
rect 230 1242 236 1243
rect 286 1243 287 1247
rect 291 1243 292 1247
rect 303 1247 304 1251
rect 308 1250 309 1251
rect 334 1251 335 1255
rect 339 1254 340 1255
rect 570 1255 576 1256
rect 339 1252 371 1254
rect 339 1251 340 1252
rect 334 1250 340 1251
rect 367 1251 373 1252
rect 308 1248 330 1250
rect 308 1247 309 1248
rect 303 1246 309 1247
rect 286 1242 292 1243
rect 328 1238 330 1248
rect 350 1247 356 1248
rect 350 1243 351 1247
rect 355 1243 356 1247
rect 367 1247 368 1251
rect 372 1247 373 1251
rect 430 1251 437 1252
rect 367 1246 373 1247
rect 414 1247 420 1248
rect 350 1242 356 1243
rect 414 1243 415 1247
rect 419 1243 420 1247
rect 430 1247 431 1251
rect 436 1247 437 1251
rect 495 1251 501 1252
rect 495 1250 496 1251
rect 488 1248 496 1250
rect 430 1246 437 1247
rect 478 1247 484 1248
rect 414 1242 420 1243
rect 478 1243 479 1247
rect 483 1243 484 1247
rect 478 1242 484 1243
rect 488 1238 490 1248
rect 495 1247 496 1248
rect 500 1247 501 1251
rect 559 1251 565 1252
rect 559 1250 560 1251
rect 552 1248 560 1250
rect 495 1246 501 1247
rect 542 1247 548 1248
rect 542 1243 543 1247
rect 547 1243 548 1247
rect 542 1242 548 1243
rect 552 1238 554 1248
rect 559 1247 560 1248
rect 564 1247 565 1251
rect 570 1251 571 1255
rect 575 1254 576 1255
rect 1296 1254 1298 1268
rect 1302 1269 1308 1270
rect 1302 1265 1303 1269
rect 1307 1265 1308 1269
rect 1302 1264 1308 1265
rect 1319 1263 1325 1264
rect 1319 1259 1320 1263
rect 1324 1262 1325 1263
rect 1352 1262 1354 1276
rect 1383 1275 1384 1279
rect 1388 1278 1389 1279
rect 1420 1278 1422 1284
rect 1430 1283 1431 1287
rect 1435 1283 1436 1287
rect 1430 1282 1436 1283
rect 1582 1285 1588 1286
rect 1582 1281 1583 1285
rect 1587 1281 1588 1285
rect 1582 1280 1588 1281
rect 1447 1279 1453 1280
rect 1447 1278 1448 1279
rect 1388 1276 1418 1278
rect 1420 1276 1448 1278
rect 1388 1275 1389 1276
rect 1383 1274 1389 1275
rect 1366 1269 1372 1270
rect 1366 1265 1367 1269
rect 1371 1265 1372 1269
rect 1366 1264 1372 1265
rect 1324 1260 1354 1262
rect 1358 1263 1364 1264
rect 1324 1259 1325 1260
rect 1319 1258 1325 1259
rect 1358 1259 1359 1263
rect 1363 1262 1364 1263
rect 1383 1263 1389 1264
rect 1383 1262 1384 1263
rect 1363 1260 1384 1262
rect 1363 1259 1364 1260
rect 1358 1258 1364 1259
rect 1383 1259 1384 1260
rect 1388 1259 1389 1263
rect 1416 1262 1418 1276
rect 1447 1275 1448 1276
rect 1452 1275 1453 1279
rect 1447 1274 1453 1275
rect 1430 1269 1436 1270
rect 1430 1265 1431 1269
rect 1435 1265 1436 1269
rect 1430 1264 1436 1265
rect 1582 1268 1588 1269
rect 1582 1264 1583 1268
rect 1587 1264 1588 1268
rect 1447 1263 1453 1264
rect 1582 1263 1588 1264
rect 1447 1262 1448 1263
rect 1416 1260 1448 1262
rect 1383 1258 1389 1259
rect 1447 1259 1448 1260
rect 1452 1259 1453 1263
rect 1447 1258 1453 1259
rect 575 1252 618 1254
rect 1296 1252 1322 1254
rect 575 1251 576 1252
rect 570 1250 576 1251
rect 616 1250 618 1252
rect 623 1251 629 1252
rect 623 1250 624 1251
rect 616 1248 624 1250
rect 559 1246 565 1247
rect 606 1247 612 1248
rect 606 1243 607 1247
rect 611 1243 612 1247
rect 623 1247 624 1248
rect 628 1247 629 1251
rect 687 1251 693 1252
rect 623 1246 629 1247
rect 670 1247 676 1248
rect 606 1242 612 1243
rect 670 1243 671 1247
rect 675 1243 676 1247
rect 687 1247 688 1251
rect 692 1247 693 1251
rect 751 1251 757 1252
rect 687 1246 693 1247
rect 734 1247 740 1248
rect 670 1242 676 1243
rect 689 1242 691 1246
rect 734 1243 735 1247
rect 739 1243 740 1247
rect 751 1247 752 1251
rect 756 1250 757 1251
rect 814 1251 821 1252
rect 756 1248 794 1250
rect 756 1247 757 1248
rect 751 1246 757 1247
rect 734 1242 740 1243
rect 689 1240 730 1242
rect 168 1236 186 1238
rect 220 1236 251 1238
rect 328 1236 362 1238
rect 465 1236 490 1238
rect 528 1236 554 1238
rect 728 1238 730 1240
rect 792 1238 794 1248
rect 798 1247 804 1248
rect 798 1243 799 1247
rect 803 1243 804 1247
rect 814 1247 815 1251
rect 820 1247 821 1251
rect 874 1251 885 1252
rect 814 1246 821 1247
rect 862 1247 868 1248
rect 798 1242 804 1243
rect 862 1243 863 1247
rect 867 1243 868 1247
rect 874 1247 875 1251
rect 879 1247 880 1251
rect 884 1247 885 1251
rect 943 1251 949 1252
rect 943 1250 944 1251
rect 936 1248 944 1250
rect 874 1246 885 1247
rect 926 1247 932 1248
rect 862 1242 868 1243
rect 926 1243 927 1247
rect 931 1243 932 1247
rect 926 1242 932 1243
rect 936 1238 938 1248
rect 943 1247 944 1248
rect 948 1247 949 1251
rect 1007 1251 1013 1252
rect 943 1246 949 1247
rect 990 1247 996 1248
rect 990 1243 991 1247
rect 995 1243 996 1247
rect 1007 1247 1008 1251
rect 1012 1250 1013 1251
rect 1031 1251 1037 1252
rect 1031 1250 1032 1251
rect 1012 1248 1032 1250
rect 1012 1247 1013 1248
rect 1007 1246 1013 1247
rect 1031 1247 1032 1248
rect 1036 1247 1037 1251
rect 1071 1251 1077 1252
rect 1071 1250 1072 1251
rect 1064 1248 1072 1250
rect 1031 1246 1037 1247
rect 1054 1247 1060 1248
rect 990 1242 996 1243
rect 1054 1243 1055 1247
rect 1059 1243 1060 1247
rect 1054 1242 1060 1243
rect 1064 1238 1066 1248
rect 1071 1247 1072 1248
rect 1076 1247 1077 1251
rect 1135 1251 1141 1252
rect 1071 1246 1077 1247
rect 1118 1247 1124 1248
rect 1118 1243 1119 1247
rect 1123 1243 1124 1247
rect 1135 1247 1136 1251
rect 1140 1250 1141 1251
rect 1174 1251 1180 1252
rect 1174 1250 1175 1251
rect 1140 1248 1175 1250
rect 1140 1247 1141 1248
rect 1135 1246 1141 1247
rect 1174 1247 1175 1248
rect 1179 1247 1180 1251
rect 1199 1251 1205 1252
rect 1199 1250 1200 1251
rect 1192 1248 1200 1250
rect 1174 1246 1180 1247
rect 1182 1247 1188 1248
rect 1118 1242 1124 1243
rect 1182 1243 1183 1247
rect 1187 1243 1188 1247
rect 1182 1242 1188 1243
rect 1192 1238 1194 1248
rect 1199 1247 1200 1248
rect 1204 1247 1205 1251
rect 1263 1251 1269 1252
rect 1263 1250 1264 1251
rect 1256 1248 1264 1250
rect 1199 1246 1205 1247
rect 1246 1247 1252 1248
rect 1246 1243 1247 1247
rect 1251 1243 1252 1247
rect 1246 1242 1252 1243
rect 1256 1238 1258 1248
rect 1263 1247 1264 1248
rect 1268 1247 1269 1251
rect 1320 1250 1322 1252
rect 1327 1251 1333 1252
rect 1327 1250 1328 1251
rect 1320 1248 1328 1250
rect 1263 1246 1269 1247
rect 1310 1247 1316 1248
rect 1310 1243 1311 1247
rect 1315 1243 1316 1247
rect 1327 1247 1328 1248
rect 1332 1247 1333 1251
rect 1391 1251 1397 1252
rect 1391 1250 1392 1251
rect 1384 1248 1392 1250
rect 1327 1246 1333 1247
rect 1374 1247 1380 1248
rect 1310 1242 1316 1243
rect 1374 1243 1375 1247
rect 1379 1243 1380 1247
rect 1374 1242 1380 1243
rect 1384 1238 1386 1248
rect 1391 1247 1392 1248
rect 1396 1247 1397 1251
rect 1455 1251 1461 1252
rect 1391 1246 1397 1247
rect 1438 1247 1444 1248
rect 1438 1243 1439 1247
rect 1443 1243 1444 1247
rect 1455 1247 1456 1251
rect 1460 1250 1461 1251
rect 1486 1251 1492 1252
rect 1486 1250 1487 1251
rect 1460 1248 1487 1250
rect 1460 1247 1461 1248
rect 1455 1246 1461 1247
rect 1486 1247 1487 1248
rect 1491 1247 1492 1251
rect 1519 1251 1525 1252
rect 1519 1250 1520 1251
rect 1512 1248 1520 1250
rect 1486 1246 1492 1247
rect 1502 1247 1508 1248
rect 1438 1242 1444 1243
rect 1502 1243 1503 1247
rect 1507 1243 1508 1247
rect 1502 1242 1508 1243
rect 1512 1238 1514 1248
rect 1519 1247 1520 1248
rect 1524 1247 1525 1251
rect 1559 1251 1565 1252
rect 1559 1250 1560 1251
rect 1552 1248 1560 1250
rect 1519 1246 1525 1247
rect 1542 1247 1548 1248
rect 1542 1243 1543 1247
rect 1547 1243 1548 1247
rect 1542 1242 1548 1243
rect 1552 1238 1554 1248
rect 1559 1247 1560 1248
rect 1564 1247 1565 1251
rect 1559 1246 1565 1247
rect 1582 1248 1588 1249
rect 1582 1244 1583 1248
rect 1587 1244 1588 1248
rect 1582 1243 1588 1244
rect 728 1236 746 1238
rect 792 1236 810 1238
rect 913 1236 938 1238
rect 1040 1236 1066 1238
rect 1168 1236 1194 1238
rect 1232 1236 1258 1238
rect 1360 1236 1386 1238
rect 1484 1236 1514 1238
rect 1540 1236 1554 1238
rect 151 1235 160 1236
rect 110 1231 116 1232
rect 110 1227 111 1231
rect 115 1227 116 1231
rect 151 1231 152 1235
rect 159 1231 160 1235
rect 184 1234 186 1236
rect 191 1235 197 1236
rect 191 1234 192 1235
rect 184 1232 192 1234
rect 151 1230 160 1231
rect 191 1231 192 1232
rect 196 1231 197 1235
rect 191 1230 197 1231
rect 247 1235 253 1236
rect 247 1231 248 1235
rect 252 1231 253 1235
rect 247 1230 253 1231
rect 302 1235 309 1236
rect 302 1231 303 1235
rect 308 1231 309 1235
rect 360 1234 362 1236
rect 367 1235 373 1236
rect 367 1234 368 1235
rect 360 1232 368 1234
rect 302 1230 309 1231
rect 367 1231 368 1232
rect 372 1231 373 1235
rect 367 1230 373 1231
rect 431 1235 437 1236
rect 431 1231 432 1235
rect 436 1234 437 1235
rect 465 1234 467 1236
rect 436 1232 467 1234
rect 495 1235 501 1236
rect 436 1231 437 1232
rect 431 1230 437 1231
rect 495 1231 496 1235
rect 500 1234 501 1235
rect 528 1234 530 1236
rect 500 1232 530 1234
rect 559 1235 565 1236
rect 500 1231 501 1232
rect 495 1230 501 1231
rect 559 1231 560 1235
rect 564 1234 565 1235
rect 570 1235 576 1236
rect 570 1234 571 1235
rect 564 1232 571 1234
rect 564 1231 565 1232
rect 559 1230 565 1231
rect 570 1231 571 1232
rect 575 1231 576 1235
rect 570 1230 576 1231
rect 618 1235 629 1236
rect 618 1231 619 1235
rect 623 1231 624 1235
rect 628 1231 629 1235
rect 618 1230 629 1231
rect 687 1235 693 1236
rect 687 1231 688 1235
rect 692 1234 693 1235
rect 702 1235 708 1236
rect 702 1234 703 1235
rect 692 1232 703 1234
rect 692 1231 693 1232
rect 687 1230 693 1231
rect 702 1231 703 1232
rect 707 1231 708 1235
rect 744 1234 746 1236
rect 751 1235 757 1236
rect 751 1234 752 1235
rect 744 1232 752 1234
rect 702 1230 708 1231
rect 751 1231 752 1232
rect 756 1231 757 1235
rect 808 1234 810 1236
rect 815 1235 821 1236
rect 815 1234 816 1235
rect 808 1232 816 1234
rect 751 1230 757 1231
rect 815 1231 816 1232
rect 820 1231 821 1235
rect 815 1230 821 1231
rect 879 1235 885 1236
rect 879 1231 880 1235
rect 884 1234 885 1235
rect 913 1234 915 1236
rect 884 1232 915 1234
rect 943 1235 952 1236
rect 884 1231 885 1232
rect 879 1230 885 1231
rect 943 1231 944 1235
rect 951 1231 952 1235
rect 943 1230 952 1231
rect 1007 1235 1013 1236
rect 1007 1231 1008 1235
rect 1012 1234 1013 1235
rect 1040 1234 1042 1236
rect 1012 1232 1042 1234
rect 1071 1235 1080 1236
rect 1012 1231 1013 1232
rect 1007 1230 1013 1231
rect 1071 1231 1072 1235
rect 1079 1231 1080 1235
rect 1071 1230 1080 1231
rect 1135 1235 1141 1236
rect 1135 1231 1136 1235
rect 1140 1234 1141 1235
rect 1168 1234 1170 1236
rect 1140 1232 1170 1234
rect 1199 1235 1205 1236
rect 1140 1231 1141 1232
rect 1135 1230 1141 1231
rect 1199 1231 1200 1235
rect 1204 1234 1205 1235
rect 1232 1234 1234 1236
rect 1204 1232 1234 1234
rect 1263 1235 1269 1236
rect 1204 1231 1205 1232
rect 1199 1230 1205 1231
rect 1263 1231 1264 1235
rect 1268 1234 1269 1235
rect 1294 1235 1300 1236
rect 1294 1234 1295 1235
rect 1268 1232 1295 1234
rect 1268 1231 1269 1232
rect 1263 1230 1269 1231
rect 1294 1231 1295 1232
rect 1299 1231 1300 1235
rect 1294 1230 1300 1231
rect 1327 1235 1333 1236
rect 1327 1231 1328 1235
rect 1332 1234 1333 1235
rect 1360 1234 1362 1236
rect 1391 1235 1397 1236
rect 1391 1234 1392 1235
rect 1332 1232 1362 1234
rect 1384 1232 1392 1234
rect 1332 1231 1333 1232
rect 1327 1230 1333 1231
rect 110 1226 116 1227
rect 134 1229 140 1230
rect 134 1225 135 1229
rect 139 1225 140 1229
rect 134 1224 140 1225
rect 174 1229 180 1230
rect 174 1225 175 1229
rect 179 1225 180 1229
rect 174 1224 180 1225
rect 230 1229 236 1230
rect 230 1225 231 1229
rect 235 1225 236 1229
rect 230 1224 236 1225
rect 286 1229 292 1230
rect 286 1225 287 1229
rect 291 1225 292 1229
rect 286 1224 292 1225
rect 350 1229 356 1230
rect 350 1225 351 1229
rect 355 1225 356 1229
rect 350 1224 356 1225
rect 414 1229 420 1230
rect 414 1225 415 1229
rect 419 1225 420 1229
rect 414 1224 420 1225
rect 478 1229 484 1230
rect 478 1225 479 1229
rect 483 1225 484 1229
rect 478 1224 484 1225
rect 542 1229 548 1230
rect 542 1225 543 1229
rect 547 1225 548 1229
rect 542 1224 548 1225
rect 606 1229 612 1230
rect 606 1225 607 1229
rect 611 1225 612 1229
rect 606 1224 612 1225
rect 670 1229 676 1230
rect 670 1225 671 1229
rect 675 1225 676 1229
rect 670 1224 676 1225
rect 734 1229 740 1230
rect 734 1225 735 1229
rect 739 1225 740 1229
rect 734 1224 740 1225
rect 798 1229 804 1230
rect 798 1225 799 1229
rect 803 1225 804 1229
rect 798 1224 804 1225
rect 862 1229 868 1230
rect 862 1225 863 1229
rect 867 1225 868 1229
rect 862 1224 868 1225
rect 926 1229 932 1230
rect 926 1225 927 1229
rect 931 1225 932 1229
rect 926 1224 932 1225
rect 990 1229 996 1230
rect 990 1225 991 1229
rect 995 1225 996 1229
rect 990 1224 996 1225
rect 1054 1229 1060 1230
rect 1054 1225 1055 1229
rect 1059 1225 1060 1229
rect 1054 1224 1060 1225
rect 1118 1229 1124 1230
rect 1118 1225 1119 1229
rect 1123 1225 1124 1229
rect 1118 1224 1124 1225
rect 1182 1229 1188 1230
rect 1182 1225 1183 1229
rect 1187 1225 1188 1229
rect 1182 1224 1188 1225
rect 1246 1229 1252 1230
rect 1246 1225 1247 1229
rect 1251 1225 1252 1229
rect 1246 1224 1252 1225
rect 1310 1229 1316 1230
rect 1310 1225 1311 1229
rect 1315 1225 1316 1229
rect 1310 1224 1316 1225
rect 1374 1229 1380 1230
rect 1374 1225 1375 1229
rect 1379 1225 1380 1229
rect 1374 1224 1380 1225
rect 294 1223 300 1224
rect 294 1219 295 1223
rect 299 1222 300 1223
rect 1046 1223 1052 1224
rect 1046 1222 1047 1223
rect 299 1220 379 1222
rect 299 1219 300 1220
rect 294 1218 300 1219
rect 142 1215 148 1216
rect 110 1213 116 1214
rect 110 1209 111 1213
rect 115 1209 116 1213
rect 142 1211 143 1215
rect 147 1211 148 1215
rect 142 1210 148 1211
rect 174 1215 180 1216
rect 174 1211 175 1215
rect 179 1211 180 1215
rect 174 1210 180 1211
rect 214 1215 220 1216
rect 214 1211 215 1215
rect 219 1211 220 1215
rect 214 1210 220 1211
rect 262 1215 268 1216
rect 262 1211 263 1215
rect 267 1211 268 1215
rect 262 1210 268 1211
rect 310 1215 316 1216
rect 310 1211 311 1215
rect 315 1211 316 1215
rect 310 1210 316 1211
rect 358 1215 364 1216
rect 358 1211 359 1215
rect 363 1211 364 1215
rect 358 1210 364 1211
rect 110 1208 116 1209
rect 377 1208 379 1220
rect 944 1220 1047 1222
rect 414 1215 420 1216
rect 414 1211 415 1215
rect 419 1211 420 1215
rect 414 1210 420 1211
rect 470 1215 476 1216
rect 470 1211 471 1215
rect 475 1211 476 1215
rect 470 1210 476 1211
rect 526 1215 532 1216
rect 526 1211 527 1215
rect 531 1211 532 1215
rect 526 1210 532 1211
rect 582 1215 588 1216
rect 582 1211 583 1215
rect 587 1211 588 1215
rect 582 1210 588 1211
rect 638 1215 644 1216
rect 638 1211 639 1215
rect 643 1211 644 1215
rect 638 1210 644 1211
rect 686 1215 692 1216
rect 686 1211 687 1215
rect 691 1211 692 1215
rect 686 1210 692 1211
rect 734 1215 740 1216
rect 734 1211 735 1215
rect 739 1211 740 1215
rect 734 1210 740 1211
rect 782 1215 788 1216
rect 782 1211 783 1215
rect 787 1211 788 1215
rect 782 1210 788 1211
rect 830 1215 836 1216
rect 830 1211 831 1215
rect 835 1211 836 1215
rect 830 1210 836 1211
rect 878 1215 884 1216
rect 878 1211 879 1215
rect 883 1211 884 1215
rect 878 1210 884 1211
rect 934 1215 940 1216
rect 934 1211 935 1215
rect 939 1211 940 1215
rect 934 1210 940 1211
rect 159 1207 165 1208
rect 159 1203 160 1207
rect 164 1206 165 1207
rect 191 1207 197 1208
rect 164 1204 186 1206
rect 164 1203 165 1204
rect 159 1202 165 1203
rect 142 1197 148 1198
rect 110 1196 116 1197
rect 110 1192 111 1196
rect 115 1192 116 1196
rect 142 1193 143 1197
rect 147 1193 148 1197
rect 142 1192 148 1193
rect 174 1197 180 1198
rect 174 1193 175 1197
rect 179 1193 180 1197
rect 174 1192 180 1193
rect 110 1191 116 1192
rect 154 1191 165 1192
rect 154 1187 155 1191
rect 159 1187 160 1191
rect 164 1187 165 1191
rect 184 1190 186 1204
rect 191 1203 192 1207
rect 196 1206 197 1207
rect 230 1207 237 1208
rect 196 1204 210 1206
rect 196 1203 197 1204
rect 191 1202 197 1203
rect 191 1191 197 1192
rect 191 1190 192 1191
rect 184 1188 192 1190
rect 154 1186 165 1187
rect 191 1187 192 1188
rect 196 1187 197 1191
rect 208 1190 210 1204
rect 230 1203 231 1207
rect 236 1203 237 1207
rect 230 1202 237 1203
rect 279 1207 285 1208
rect 279 1203 280 1207
rect 284 1206 285 1207
rect 327 1207 333 1208
rect 284 1204 322 1206
rect 284 1203 285 1204
rect 279 1202 285 1203
rect 214 1197 220 1198
rect 214 1193 215 1197
rect 219 1193 220 1197
rect 214 1192 220 1193
rect 262 1197 268 1198
rect 262 1193 263 1197
rect 267 1193 268 1197
rect 262 1192 268 1193
rect 310 1197 316 1198
rect 310 1193 311 1197
rect 315 1193 316 1197
rect 310 1192 316 1193
rect 231 1191 237 1192
rect 231 1190 232 1191
rect 208 1188 232 1190
rect 191 1186 197 1187
rect 231 1187 232 1188
rect 236 1187 237 1191
rect 231 1186 237 1187
rect 279 1191 285 1192
rect 279 1187 280 1191
rect 284 1190 285 1191
rect 294 1191 300 1192
rect 294 1190 295 1191
rect 284 1188 295 1190
rect 284 1187 285 1188
rect 279 1186 285 1187
rect 294 1187 295 1188
rect 299 1187 300 1191
rect 320 1190 322 1204
rect 327 1203 328 1207
rect 332 1203 333 1207
rect 327 1202 333 1203
rect 375 1207 381 1208
rect 375 1203 376 1207
rect 380 1203 381 1207
rect 375 1202 381 1203
rect 430 1207 437 1208
rect 430 1203 431 1207
rect 436 1203 437 1207
rect 487 1207 493 1208
rect 487 1206 488 1207
rect 430 1202 437 1203
rect 464 1204 488 1206
rect 358 1197 364 1198
rect 358 1193 359 1197
rect 363 1193 364 1197
rect 358 1192 364 1193
rect 414 1197 420 1198
rect 414 1193 415 1197
rect 419 1193 420 1197
rect 414 1192 420 1193
rect 327 1191 333 1192
rect 327 1190 328 1191
rect 320 1188 328 1190
rect 294 1186 300 1187
rect 327 1187 328 1188
rect 332 1187 333 1191
rect 327 1186 333 1187
rect 375 1191 381 1192
rect 375 1187 376 1191
rect 380 1190 381 1191
rect 422 1191 428 1192
rect 422 1190 423 1191
rect 380 1188 423 1190
rect 380 1187 381 1188
rect 375 1186 381 1187
rect 422 1187 423 1188
rect 427 1187 428 1191
rect 422 1186 428 1187
rect 431 1191 437 1192
rect 431 1187 432 1191
rect 436 1190 437 1191
rect 464 1190 466 1204
rect 487 1203 488 1204
rect 492 1203 493 1207
rect 543 1207 549 1208
rect 543 1206 544 1207
rect 487 1202 493 1203
rect 520 1204 544 1206
rect 470 1197 476 1198
rect 470 1193 471 1197
rect 475 1193 476 1197
rect 470 1192 476 1193
rect 436 1188 466 1190
rect 487 1191 493 1192
rect 436 1187 437 1188
rect 431 1186 437 1187
rect 487 1187 488 1191
rect 492 1190 493 1191
rect 520 1190 522 1204
rect 543 1203 544 1204
rect 548 1203 549 1207
rect 599 1207 605 1208
rect 599 1206 600 1207
rect 543 1202 549 1203
rect 576 1204 600 1206
rect 526 1197 532 1198
rect 526 1193 527 1197
rect 531 1193 532 1197
rect 526 1192 532 1193
rect 492 1188 522 1190
rect 543 1191 549 1192
rect 492 1187 493 1188
rect 487 1186 493 1187
rect 543 1187 544 1191
rect 548 1190 549 1191
rect 576 1190 578 1204
rect 599 1203 600 1204
rect 604 1203 605 1207
rect 655 1207 661 1208
rect 655 1206 656 1207
rect 599 1202 605 1203
rect 624 1204 656 1206
rect 624 1198 626 1204
rect 655 1203 656 1204
rect 660 1203 661 1207
rect 655 1202 661 1203
rect 703 1207 709 1208
rect 703 1203 704 1207
rect 708 1206 709 1207
rect 751 1207 757 1208
rect 708 1204 730 1206
rect 708 1203 709 1204
rect 703 1202 709 1203
rect 582 1197 588 1198
rect 582 1193 583 1197
rect 587 1193 588 1197
rect 582 1192 588 1193
rect 604 1196 626 1198
rect 638 1197 644 1198
rect 604 1192 606 1196
rect 638 1193 639 1197
rect 643 1193 644 1197
rect 638 1192 644 1193
rect 686 1197 692 1198
rect 686 1193 687 1197
rect 691 1193 692 1197
rect 686 1192 692 1193
rect 548 1188 578 1190
rect 599 1191 606 1192
rect 548 1187 549 1188
rect 543 1186 549 1187
rect 599 1187 600 1191
rect 604 1188 606 1191
rect 610 1191 616 1192
rect 604 1187 605 1188
rect 599 1186 605 1187
rect 610 1187 611 1191
rect 615 1190 616 1191
rect 655 1191 661 1192
rect 655 1190 656 1191
rect 615 1188 656 1190
rect 615 1187 616 1188
rect 610 1186 616 1187
rect 655 1187 656 1188
rect 660 1187 661 1191
rect 655 1186 661 1187
rect 702 1191 709 1192
rect 702 1187 703 1191
rect 708 1187 709 1191
rect 728 1190 730 1204
rect 751 1203 752 1207
rect 756 1206 757 1207
rect 799 1207 805 1208
rect 756 1204 778 1206
rect 756 1203 757 1204
rect 751 1202 757 1203
rect 734 1197 740 1198
rect 734 1193 735 1197
rect 739 1193 740 1197
rect 734 1192 740 1193
rect 751 1191 757 1192
rect 751 1190 752 1191
rect 728 1188 752 1190
rect 702 1186 709 1187
rect 751 1187 752 1188
rect 756 1187 757 1191
rect 776 1190 778 1204
rect 799 1203 800 1207
rect 804 1206 805 1207
rect 847 1207 853 1208
rect 804 1204 842 1206
rect 804 1203 805 1204
rect 799 1202 805 1203
rect 782 1197 788 1198
rect 782 1193 783 1197
rect 787 1193 788 1197
rect 782 1192 788 1193
rect 830 1197 836 1198
rect 830 1193 831 1197
rect 835 1193 836 1197
rect 830 1192 836 1193
rect 799 1191 805 1192
rect 799 1190 800 1191
rect 776 1188 800 1190
rect 751 1186 757 1187
rect 799 1187 800 1188
rect 804 1187 805 1191
rect 840 1190 842 1204
rect 847 1203 848 1207
rect 852 1206 853 1207
rect 895 1207 901 1208
rect 852 1204 874 1206
rect 852 1203 853 1204
rect 847 1202 853 1203
rect 847 1191 853 1192
rect 847 1190 848 1191
rect 840 1188 848 1190
rect 799 1186 805 1187
rect 847 1187 848 1188
rect 852 1187 853 1191
rect 872 1190 874 1204
rect 895 1203 896 1207
rect 900 1206 901 1207
rect 944 1206 946 1220
rect 1046 1219 1047 1220
rect 1051 1219 1052 1223
rect 1046 1218 1052 1219
rect 1174 1223 1180 1224
rect 1174 1219 1175 1223
rect 1179 1222 1180 1223
rect 1384 1222 1386 1232
rect 1391 1231 1392 1232
rect 1396 1231 1397 1235
rect 1391 1230 1397 1231
rect 1455 1235 1461 1236
rect 1455 1231 1456 1235
rect 1460 1234 1461 1235
rect 1484 1234 1486 1236
rect 1460 1232 1486 1234
rect 1519 1235 1525 1236
rect 1460 1231 1461 1232
rect 1455 1230 1461 1231
rect 1519 1231 1520 1235
rect 1524 1234 1525 1235
rect 1540 1234 1542 1236
rect 1524 1232 1542 1234
rect 1558 1235 1565 1236
rect 1524 1231 1525 1232
rect 1519 1230 1525 1231
rect 1558 1231 1559 1235
rect 1564 1231 1565 1235
rect 1558 1230 1565 1231
rect 1582 1231 1588 1232
rect 1438 1229 1444 1230
rect 1438 1225 1439 1229
rect 1443 1225 1444 1229
rect 1438 1224 1444 1225
rect 1502 1229 1508 1230
rect 1502 1225 1503 1229
rect 1507 1225 1508 1229
rect 1502 1224 1508 1225
rect 1542 1229 1548 1230
rect 1542 1225 1543 1229
rect 1547 1225 1548 1229
rect 1582 1227 1583 1231
rect 1587 1227 1588 1231
rect 1582 1226 1588 1227
rect 1542 1224 1548 1225
rect 1179 1220 1386 1222
rect 1179 1219 1180 1220
rect 1174 1218 1180 1219
rect 982 1215 988 1216
rect 982 1211 983 1215
rect 987 1211 988 1215
rect 982 1210 988 1211
rect 1038 1215 1044 1216
rect 1038 1211 1039 1215
rect 1043 1211 1044 1215
rect 1038 1210 1044 1211
rect 1094 1215 1100 1216
rect 1094 1211 1095 1215
rect 1099 1211 1100 1215
rect 1094 1210 1100 1211
rect 1158 1215 1164 1216
rect 1158 1211 1159 1215
rect 1163 1211 1164 1215
rect 1158 1210 1164 1211
rect 1230 1215 1236 1216
rect 1230 1211 1231 1215
rect 1235 1211 1236 1215
rect 1230 1210 1236 1211
rect 1302 1215 1308 1216
rect 1302 1211 1303 1215
rect 1307 1211 1308 1215
rect 1382 1215 1388 1216
rect 1302 1210 1308 1211
rect 1312 1212 1366 1214
rect 900 1204 946 1206
rect 951 1207 957 1208
rect 900 1203 901 1204
rect 895 1202 901 1203
rect 951 1203 952 1207
rect 956 1206 957 1207
rect 998 1207 1005 1208
rect 956 1204 978 1206
rect 956 1203 957 1204
rect 951 1202 957 1203
rect 878 1197 884 1198
rect 878 1193 879 1197
rect 883 1193 884 1197
rect 878 1192 884 1193
rect 934 1197 940 1198
rect 934 1193 935 1197
rect 939 1193 940 1197
rect 934 1192 940 1193
rect 895 1191 901 1192
rect 895 1190 896 1191
rect 872 1188 896 1190
rect 847 1186 853 1187
rect 895 1187 896 1188
rect 900 1187 901 1191
rect 895 1186 901 1187
rect 946 1191 957 1192
rect 946 1187 947 1191
rect 951 1187 952 1191
rect 956 1187 957 1191
rect 976 1190 978 1204
rect 998 1203 999 1207
rect 1004 1203 1005 1207
rect 998 1202 1005 1203
rect 1031 1207 1037 1208
rect 1031 1203 1032 1207
rect 1036 1206 1037 1207
rect 1055 1207 1061 1208
rect 1055 1206 1056 1207
rect 1036 1204 1056 1206
rect 1036 1203 1037 1204
rect 1031 1202 1037 1203
rect 1055 1203 1056 1204
rect 1060 1203 1061 1207
rect 1055 1202 1061 1203
rect 1063 1207 1069 1208
rect 1063 1203 1064 1207
rect 1068 1206 1069 1207
rect 1111 1207 1117 1208
rect 1111 1206 1112 1207
rect 1068 1204 1112 1206
rect 1068 1203 1069 1204
rect 1063 1202 1069 1203
rect 1111 1203 1112 1204
rect 1116 1203 1117 1207
rect 1175 1207 1181 1208
rect 1175 1206 1176 1207
rect 1111 1202 1117 1203
rect 1145 1204 1176 1206
rect 982 1197 988 1198
rect 982 1193 983 1197
rect 987 1193 988 1197
rect 982 1192 988 1193
rect 1038 1197 1044 1198
rect 1038 1193 1039 1197
rect 1043 1193 1044 1197
rect 1038 1192 1044 1193
rect 1094 1197 1100 1198
rect 1094 1193 1095 1197
rect 1099 1193 1100 1197
rect 1094 1192 1100 1193
rect 999 1191 1005 1192
rect 999 1190 1000 1191
rect 976 1188 1000 1190
rect 946 1186 957 1187
rect 999 1187 1000 1188
rect 1004 1187 1005 1191
rect 999 1186 1005 1187
rect 1046 1191 1052 1192
rect 1046 1187 1047 1191
rect 1051 1190 1052 1191
rect 1055 1191 1061 1192
rect 1055 1190 1056 1191
rect 1051 1188 1056 1190
rect 1051 1187 1052 1188
rect 1046 1186 1052 1187
rect 1055 1187 1056 1188
rect 1060 1187 1061 1191
rect 1055 1186 1061 1187
rect 1111 1191 1117 1192
rect 1111 1187 1112 1191
rect 1116 1190 1117 1191
rect 1145 1190 1147 1204
rect 1175 1203 1176 1204
rect 1180 1203 1181 1207
rect 1247 1207 1253 1208
rect 1247 1206 1248 1207
rect 1175 1202 1181 1203
rect 1212 1204 1248 1206
rect 1158 1197 1164 1198
rect 1158 1193 1159 1197
rect 1163 1193 1164 1197
rect 1158 1192 1164 1193
rect 1116 1188 1147 1190
rect 1175 1191 1181 1192
rect 1116 1187 1117 1188
rect 1111 1186 1117 1187
rect 1175 1187 1176 1191
rect 1180 1190 1181 1191
rect 1212 1190 1214 1204
rect 1247 1203 1248 1204
rect 1252 1203 1253 1207
rect 1312 1206 1314 1212
rect 1247 1202 1253 1203
rect 1288 1204 1314 1206
rect 1319 1207 1325 1208
rect 1230 1197 1236 1198
rect 1230 1193 1231 1197
rect 1235 1193 1236 1197
rect 1230 1192 1236 1193
rect 1180 1188 1214 1190
rect 1247 1191 1253 1192
rect 1180 1187 1181 1188
rect 1175 1186 1181 1187
rect 1247 1187 1248 1191
rect 1252 1190 1253 1191
rect 1288 1190 1290 1204
rect 1319 1203 1320 1207
rect 1324 1206 1325 1207
rect 1364 1206 1366 1212
rect 1382 1211 1383 1215
rect 1387 1211 1388 1215
rect 1382 1210 1388 1211
rect 1470 1215 1476 1216
rect 1470 1211 1471 1215
rect 1475 1211 1476 1215
rect 1470 1210 1476 1211
rect 1542 1215 1548 1216
rect 1542 1211 1543 1215
rect 1547 1211 1548 1215
rect 1542 1210 1548 1211
rect 1582 1213 1588 1214
rect 1582 1209 1583 1213
rect 1587 1209 1588 1213
rect 1582 1208 1588 1209
rect 1399 1207 1405 1208
rect 1399 1206 1400 1207
rect 1324 1204 1362 1206
rect 1364 1204 1400 1206
rect 1324 1203 1325 1204
rect 1319 1202 1325 1203
rect 1302 1197 1308 1198
rect 1302 1193 1303 1197
rect 1307 1193 1308 1197
rect 1302 1192 1308 1193
rect 1252 1188 1290 1190
rect 1294 1191 1300 1192
rect 1252 1187 1253 1188
rect 1247 1186 1253 1187
rect 1294 1187 1295 1191
rect 1299 1190 1300 1191
rect 1319 1191 1325 1192
rect 1319 1190 1320 1191
rect 1299 1188 1320 1190
rect 1299 1187 1300 1188
rect 1294 1186 1300 1187
rect 1319 1187 1320 1188
rect 1324 1187 1325 1191
rect 1360 1190 1362 1204
rect 1399 1203 1400 1204
rect 1404 1203 1405 1207
rect 1399 1202 1405 1203
rect 1486 1207 1493 1208
rect 1486 1203 1487 1207
rect 1492 1203 1493 1207
rect 1486 1202 1493 1203
rect 1559 1207 1565 1208
rect 1559 1203 1560 1207
rect 1564 1206 1565 1207
rect 1567 1207 1573 1208
rect 1567 1206 1568 1207
rect 1564 1204 1568 1206
rect 1564 1203 1565 1204
rect 1559 1202 1565 1203
rect 1567 1203 1568 1204
rect 1572 1203 1573 1207
rect 1567 1202 1573 1203
rect 1382 1197 1388 1198
rect 1382 1193 1383 1197
rect 1387 1193 1388 1197
rect 1382 1192 1388 1193
rect 1470 1197 1476 1198
rect 1470 1193 1471 1197
rect 1475 1193 1476 1197
rect 1470 1192 1476 1193
rect 1542 1197 1548 1198
rect 1542 1193 1543 1197
rect 1547 1193 1548 1197
rect 1542 1192 1548 1193
rect 1582 1196 1588 1197
rect 1582 1192 1583 1196
rect 1587 1192 1588 1196
rect 1399 1191 1405 1192
rect 1399 1190 1400 1191
rect 1360 1188 1400 1190
rect 1319 1186 1325 1187
rect 1399 1187 1400 1188
rect 1404 1187 1405 1191
rect 1399 1186 1405 1187
rect 1487 1191 1493 1192
rect 1487 1187 1488 1191
rect 1492 1187 1493 1191
rect 1487 1186 1493 1187
rect 1558 1191 1565 1192
rect 1582 1191 1588 1192
rect 1558 1187 1559 1191
rect 1564 1187 1565 1191
rect 1558 1186 1565 1187
rect 159 1179 165 1180
rect 110 1176 116 1177
rect 110 1172 111 1176
rect 115 1172 116 1176
rect 110 1171 116 1172
rect 142 1175 148 1176
rect 142 1171 143 1175
rect 147 1171 148 1175
rect 159 1175 160 1179
rect 164 1178 165 1179
rect 191 1179 197 1180
rect 164 1176 170 1178
rect 164 1175 165 1176
rect 159 1174 165 1175
rect 142 1170 148 1171
rect 168 1166 170 1176
rect 174 1175 180 1176
rect 174 1171 175 1175
rect 179 1171 180 1175
rect 191 1175 192 1179
rect 196 1178 197 1179
rect 230 1179 237 1180
rect 196 1176 210 1178
rect 196 1175 197 1176
rect 191 1174 197 1175
rect 174 1170 180 1171
rect 208 1166 210 1176
rect 214 1175 220 1176
rect 214 1171 215 1175
rect 219 1171 220 1175
rect 230 1175 231 1179
rect 236 1175 237 1179
rect 271 1179 277 1180
rect 230 1174 237 1175
rect 254 1175 260 1176
rect 214 1170 220 1171
rect 254 1171 255 1175
rect 259 1171 260 1175
rect 271 1175 272 1179
rect 276 1178 277 1179
rect 287 1179 293 1180
rect 287 1178 288 1179
rect 276 1176 288 1178
rect 276 1175 277 1176
rect 271 1174 277 1175
rect 287 1175 288 1176
rect 292 1175 293 1179
rect 319 1179 325 1180
rect 319 1178 320 1179
rect 312 1176 320 1178
rect 287 1174 293 1175
rect 302 1175 308 1176
rect 254 1170 260 1171
rect 302 1171 303 1175
rect 307 1171 308 1175
rect 302 1170 308 1171
rect 312 1166 314 1176
rect 319 1175 320 1176
rect 324 1175 325 1179
rect 375 1179 381 1180
rect 375 1178 376 1179
rect 368 1176 376 1178
rect 319 1174 325 1175
rect 358 1175 364 1176
rect 358 1171 359 1175
rect 363 1171 364 1175
rect 358 1170 364 1171
rect 368 1166 370 1176
rect 375 1175 376 1176
rect 380 1175 381 1179
rect 431 1179 437 1180
rect 431 1178 432 1179
rect 424 1176 432 1178
rect 375 1174 381 1175
rect 414 1175 420 1176
rect 414 1171 415 1175
rect 419 1171 420 1175
rect 414 1170 420 1171
rect 424 1166 426 1176
rect 431 1175 432 1176
rect 436 1175 437 1179
rect 487 1179 493 1180
rect 431 1174 437 1175
rect 470 1175 476 1176
rect 470 1171 471 1175
rect 475 1171 476 1175
rect 487 1175 488 1179
rect 492 1178 493 1179
rect 518 1179 524 1180
rect 518 1178 519 1179
rect 492 1176 519 1178
rect 492 1175 493 1176
rect 487 1174 493 1175
rect 518 1175 519 1176
rect 523 1175 524 1179
rect 543 1179 549 1180
rect 543 1178 544 1179
rect 536 1176 544 1178
rect 518 1174 524 1175
rect 526 1175 532 1176
rect 470 1170 476 1171
rect 526 1171 527 1175
rect 531 1171 532 1175
rect 526 1170 532 1171
rect 536 1166 538 1176
rect 543 1175 544 1176
rect 548 1175 549 1179
rect 607 1179 613 1180
rect 607 1178 608 1179
rect 600 1176 608 1178
rect 543 1174 549 1175
rect 590 1175 596 1176
rect 590 1171 591 1175
rect 595 1171 596 1175
rect 590 1170 596 1171
rect 600 1166 602 1176
rect 607 1175 608 1176
rect 612 1175 613 1179
rect 671 1179 677 1180
rect 607 1174 613 1175
rect 654 1175 660 1176
rect 654 1171 655 1175
rect 659 1171 660 1175
rect 671 1175 672 1179
rect 676 1178 677 1179
rect 735 1179 741 1180
rect 676 1176 714 1178
rect 676 1175 677 1176
rect 671 1174 677 1175
rect 654 1170 660 1171
rect 168 1164 186 1166
rect 208 1164 226 1166
rect 296 1164 314 1166
rect 348 1164 370 1166
rect 377 1164 426 1166
rect 516 1164 538 1166
rect 577 1164 602 1166
rect 712 1166 714 1176
rect 718 1175 724 1176
rect 718 1171 719 1175
rect 723 1171 724 1175
rect 735 1175 736 1179
rect 740 1178 741 1179
rect 802 1179 813 1180
rect 740 1176 778 1178
rect 740 1175 741 1176
rect 735 1174 741 1175
rect 718 1170 724 1171
rect 776 1166 778 1176
rect 790 1175 796 1176
rect 790 1171 791 1175
rect 795 1171 796 1175
rect 802 1175 803 1179
rect 807 1175 808 1179
rect 812 1175 813 1179
rect 871 1179 877 1180
rect 802 1174 813 1175
rect 854 1175 860 1176
rect 790 1170 796 1171
rect 854 1171 855 1175
rect 859 1171 860 1175
rect 871 1175 872 1179
rect 876 1178 877 1179
rect 935 1179 941 1180
rect 876 1176 914 1178
rect 876 1175 877 1176
rect 871 1174 877 1175
rect 854 1170 860 1171
rect 912 1166 914 1176
rect 918 1175 924 1176
rect 918 1171 919 1175
rect 923 1171 924 1175
rect 935 1175 936 1179
rect 940 1178 941 1179
rect 998 1179 1005 1180
rect 940 1176 978 1178
rect 940 1175 941 1176
rect 935 1174 941 1175
rect 918 1170 924 1171
rect 976 1166 978 1176
rect 982 1175 988 1176
rect 982 1171 983 1175
rect 987 1171 988 1175
rect 998 1175 999 1179
rect 1004 1175 1005 1179
rect 1055 1179 1061 1180
rect 998 1174 1005 1175
rect 1038 1175 1044 1176
rect 982 1170 988 1171
rect 1038 1171 1039 1175
rect 1043 1171 1044 1175
rect 1055 1175 1056 1179
rect 1060 1178 1061 1179
rect 1063 1179 1069 1180
rect 1063 1178 1064 1179
rect 1060 1176 1064 1178
rect 1060 1175 1061 1176
rect 1055 1174 1061 1175
rect 1063 1175 1064 1176
rect 1068 1175 1069 1179
rect 1119 1179 1125 1180
rect 1119 1178 1120 1179
rect 1112 1176 1120 1178
rect 1063 1174 1069 1175
rect 1102 1175 1108 1176
rect 1038 1170 1044 1171
rect 1102 1171 1103 1175
rect 1107 1171 1108 1175
rect 1102 1170 1108 1171
rect 1112 1166 1114 1176
rect 1119 1175 1120 1176
rect 1124 1175 1125 1179
rect 1183 1179 1189 1180
rect 1183 1178 1184 1179
rect 1176 1176 1184 1178
rect 1119 1174 1125 1175
rect 1166 1175 1172 1176
rect 1166 1171 1167 1175
rect 1171 1171 1172 1175
rect 1166 1170 1172 1171
rect 1176 1166 1178 1176
rect 1183 1175 1184 1176
rect 1188 1175 1189 1179
rect 1255 1179 1261 1180
rect 1255 1178 1256 1179
rect 1248 1176 1256 1178
rect 1183 1174 1189 1175
rect 1238 1175 1244 1176
rect 1238 1171 1239 1175
rect 1243 1171 1244 1175
rect 1238 1170 1244 1171
rect 1248 1166 1250 1176
rect 1255 1175 1256 1176
rect 1260 1175 1261 1179
rect 1327 1179 1333 1180
rect 1327 1178 1328 1179
rect 1320 1176 1328 1178
rect 1255 1174 1261 1175
rect 1310 1175 1316 1176
rect 1310 1171 1311 1175
rect 1315 1171 1316 1175
rect 1310 1170 1316 1171
rect 1320 1166 1322 1176
rect 1327 1175 1328 1176
rect 1332 1175 1333 1179
rect 1407 1179 1413 1180
rect 1407 1178 1408 1179
rect 1400 1176 1408 1178
rect 1327 1174 1333 1175
rect 1390 1175 1396 1176
rect 1390 1171 1391 1175
rect 1395 1171 1396 1175
rect 1390 1170 1396 1171
rect 1400 1166 1402 1176
rect 1407 1175 1408 1176
rect 1412 1175 1413 1179
rect 1407 1174 1413 1175
rect 1478 1175 1484 1176
rect 1478 1171 1479 1175
rect 1483 1171 1484 1175
rect 1478 1170 1484 1171
rect 712 1164 730 1166
rect 776 1164 802 1166
rect 912 1164 930 1166
rect 976 1164 994 1166
rect 1099 1164 1114 1166
rect 1152 1164 1178 1166
rect 1220 1164 1250 1166
rect 1292 1164 1322 1166
rect 1368 1164 1402 1166
rect 154 1163 165 1164
rect 110 1159 116 1160
rect 110 1155 111 1159
rect 115 1155 116 1159
rect 154 1159 155 1163
rect 159 1159 160 1163
rect 164 1159 165 1163
rect 184 1162 186 1164
rect 191 1163 197 1164
rect 191 1162 192 1163
rect 184 1160 192 1162
rect 154 1158 165 1159
rect 191 1159 192 1160
rect 196 1159 197 1163
rect 224 1162 226 1164
rect 231 1163 237 1164
rect 231 1162 232 1163
rect 224 1160 232 1162
rect 191 1158 197 1159
rect 231 1159 232 1160
rect 236 1159 237 1163
rect 231 1158 237 1159
rect 271 1163 277 1164
rect 271 1159 272 1163
rect 276 1162 277 1163
rect 296 1162 298 1164
rect 276 1160 298 1162
rect 319 1163 325 1164
rect 276 1159 277 1160
rect 271 1158 277 1159
rect 319 1159 320 1163
rect 324 1162 325 1163
rect 348 1162 350 1164
rect 324 1160 350 1162
rect 375 1163 381 1164
rect 324 1159 325 1160
rect 319 1158 325 1159
rect 375 1159 376 1163
rect 380 1159 381 1163
rect 375 1158 381 1159
rect 430 1163 437 1164
rect 430 1159 431 1163
rect 436 1159 437 1163
rect 430 1158 437 1159
rect 487 1163 493 1164
rect 487 1159 488 1163
rect 492 1162 493 1163
rect 516 1162 518 1164
rect 492 1160 518 1162
rect 543 1163 549 1164
rect 492 1159 493 1160
rect 487 1158 493 1159
rect 543 1159 544 1163
rect 548 1162 549 1163
rect 577 1162 579 1164
rect 548 1160 579 1162
rect 607 1163 616 1164
rect 548 1159 549 1160
rect 543 1158 549 1159
rect 607 1159 608 1163
rect 615 1159 616 1163
rect 671 1163 677 1164
rect 671 1162 672 1163
rect 607 1158 616 1159
rect 664 1160 672 1162
rect 110 1154 116 1155
rect 142 1157 148 1158
rect 142 1153 143 1157
rect 147 1153 148 1157
rect 142 1152 148 1153
rect 174 1157 180 1158
rect 174 1153 175 1157
rect 179 1153 180 1157
rect 174 1152 180 1153
rect 214 1157 220 1158
rect 214 1153 215 1157
rect 219 1153 220 1157
rect 214 1152 220 1153
rect 254 1157 260 1158
rect 254 1153 255 1157
rect 259 1153 260 1157
rect 254 1152 260 1153
rect 302 1157 308 1158
rect 302 1153 303 1157
rect 307 1153 308 1157
rect 302 1152 308 1153
rect 358 1157 364 1158
rect 358 1153 359 1157
rect 363 1153 364 1157
rect 358 1152 364 1153
rect 414 1157 420 1158
rect 414 1153 415 1157
rect 419 1153 420 1157
rect 414 1152 420 1153
rect 470 1157 476 1158
rect 470 1153 471 1157
rect 475 1153 476 1157
rect 470 1152 476 1153
rect 526 1157 532 1158
rect 526 1153 527 1157
rect 531 1153 532 1157
rect 526 1152 532 1153
rect 590 1157 596 1158
rect 590 1153 591 1157
rect 595 1153 596 1157
rect 590 1152 596 1153
rect 654 1157 660 1158
rect 654 1153 655 1157
rect 659 1153 660 1157
rect 654 1152 660 1153
rect 287 1151 293 1152
rect 287 1147 288 1151
rect 292 1150 293 1151
rect 518 1151 524 1152
rect 292 1148 498 1150
rect 292 1147 293 1148
rect 287 1146 293 1147
rect 134 1143 140 1144
rect 110 1141 116 1142
rect 110 1137 111 1141
rect 115 1137 116 1141
rect 134 1139 135 1143
rect 139 1139 140 1143
rect 134 1138 140 1139
rect 166 1143 172 1144
rect 166 1139 167 1143
rect 171 1139 172 1143
rect 166 1138 172 1139
rect 198 1143 204 1144
rect 198 1139 199 1143
rect 203 1139 204 1143
rect 198 1138 204 1139
rect 230 1143 236 1144
rect 230 1139 231 1143
rect 235 1139 236 1143
rect 230 1138 236 1139
rect 262 1143 268 1144
rect 262 1139 263 1143
rect 267 1139 268 1143
rect 262 1138 268 1139
rect 294 1143 300 1144
rect 294 1139 295 1143
rect 299 1139 300 1143
rect 294 1138 300 1139
rect 326 1143 332 1144
rect 326 1139 327 1143
rect 331 1139 332 1143
rect 326 1138 332 1139
rect 358 1143 364 1144
rect 358 1139 359 1143
rect 363 1139 364 1143
rect 358 1138 364 1139
rect 390 1143 396 1144
rect 390 1139 391 1143
rect 395 1139 396 1143
rect 390 1138 396 1139
rect 446 1143 452 1144
rect 446 1139 447 1143
rect 451 1139 452 1143
rect 446 1138 452 1139
rect 110 1136 116 1137
rect 151 1135 157 1136
rect 151 1131 152 1135
rect 156 1134 157 1135
rect 183 1135 189 1136
rect 156 1132 178 1134
rect 156 1131 157 1132
rect 151 1130 157 1131
rect 134 1125 140 1126
rect 110 1124 116 1125
rect 110 1120 111 1124
rect 115 1120 116 1124
rect 134 1121 135 1125
rect 139 1121 140 1125
rect 166 1125 172 1126
rect 134 1120 140 1121
rect 154 1123 160 1124
rect 154 1120 155 1123
rect 110 1119 116 1120
rect 151 1119 155 1120
rect 159 1119 160 1123
rect 166 1121 167 1125
rect 171 1121 172 1125
rect 166 1120 172 1121
rect 151 1115 152 1119
rect 156 1118 160 1119
rect 176 1118 178 1132
rect 183 1131 184 1135
rect 188 1134 189 1135
rect 215 1135 221 1136
rect 188 1132 210 1134
rect 188 1131 189 1132
rect 183 1130 189 1131
rect 198 1125 204 1126
rect 198 1121 199 1125
rect 203 1121 204 1125
rect 198 1120 204 1121
rect 183 1119 189 1120
rect 183 1118 184 1119
rect 156 1116 158 1118
rect 176 1116 184 1118
rect 156 1115 157 1116
rect 151 1114 157 1115
rect 183 1115 184 1116
rect 188 1115 189 1119
rect 208 1118 210 1132
rect 215 1131 216 1135
rect 220 1134 221 1135
rect 247 1135 253 1136
rect 220 1132 242 1134
rect 220 1131 221 1132
rect 215 1130 221 1131
rect 230 1125 236 1126
rect 230 1121 231 1125
rect 235 1121 236 1125
rect 230 1120 236 1121
rect 215 1119 221 1120
rect 215 1118 216 1119
rect 208 1116 216 1118
rect 183 1114 189 1115
rect 215 1115 216 1116
rect 220 1115 221 1119
rect 240 1118 242 1132
rect 247 1131 248 1135
rect 252 1134 253 1135
rect 279 1135 285 1136
rect 252 1132 274 1134
rect 252 1131 253 1132
rect 247 1130 253 1131
rect 262 1125 268 1126
rect 262 1121 263 1125
rect 267 1121 268 1125
rect 262 1120 268 1121
rect 247 1119 253 1120
rect 247 1118 248 1119
rect 240 1116 248 1118
rect 215 1114 221 1115
rect 247 1115 248 1116
rect 252 1115 253 1119
rect 272 1118 274 1132
rect 279 1131 280 1135
rect 284 1134 285 1135
rect 310 1135 317 1136
rect 284 1132 306 1134
rect 284 1131 285 1132
rect 279 1130 285 1131
rect 294 1125 300 1126
rect 294 1121 295 1125
rect 299 1121 300 1125
rect 294 1120 300 1121
rect 279 1119 285 1120
rect 279 1118 280 1119
rect 272 1116 280 1118
rect 247 1114 253 1115
rect 279 1115 280 1116
rect 284 1115 285 1119
rect 304 1118 306 1132
rect 310 1131 311 1135
rect 316 1131 317 1135
rect 310 1130 317 1131
rect 343 1135 349 1136
rect 343 1131 344 1135
rect 348 1134 349 1135
rect 375 1135 381 1136
rect 348 1132 370 1134
rect 348 1131 349 1132
rect 343 1130 349 1131
rect 326 1125 332 1126
rect 326 1121 327 1125
rect 331 1121 332 1125
rect 326 1120 332 1121
rect 358 1125 364 1126
rect 358 1121 359 1125
rect 363 1121 364 1125
rect 358 1120 364 1121
rect 311 1119 317 1120
rect 311 1118 312 1119
rect 304 1116 312 1118
rect 279 1114 285 1115
rect 311 1115 312 1116
rect 316 1115 317 1119
rect 311 1114 317 1115
rect 343 1119 352 1120
rect 343 1115 344 1119
rect 351 1115 352 1119
rect 368 1118 370 1132
rect 375 1131 376 1135
rect 380 1134 381 1135
rect 407 1135 413 1136
rect 380 1132 402 1134
rect 380 1131 381 1132
rect 375 1130 381 1131
rect 390 1125 396 1126
rect 390 1121 391 1125
rect 395 1121 396 1125
rect 390 1120 396 1121
rect 375 1119 381 1120
rect 375 1118 376 1119
rect 368 1116 376 1118
rect 343 1114 352 1115
rect 375 1115 376 1116
rect 380 1115 381 1119
rect 400 1118 402 1132
rect 407 1131 408 1135
rect 412 1134 413 1135
rect 463 1135 469 1136
rect 412 1132 438 1134
rect 412 1131 413 1132
rect 407 1130 413 1131
rect 407 1119 413 1120
rect 407 1118 408 1119
rect 400 1116 408 1118
rect 375 1114 381 1115
rect 407 1115 408 1116
rect 412 1115 413 1119
rect 436 1118 438 1132
rect 463 1131 464 1135
rect 468 1134 469 1135
rect 496 1134 498 1148
rect 518 1147 519 1151
rect 523 1150 524 1151
rect 664 1150 666 1160
rect 671 1159 672 1160
rect 676 1159 677 1163
rect 728 1162 730 1164
rect 735 1163 741 1164
rect 735 1162 736 1163
rect 728 1160 736 1162
rect 671 1158 677 1159
rect 735 1159 736 1160
rect 740 1159 741 1163
rect 800 1162 802 1164
rect 807 1163 813 1164
rect 807 1162 808 1163
rect 800 1160 808 1162
rect 735 1158 741 1159
rect 807 1159 808 1160
rect 812 1159 813 1163
rect 807 1158 813 1159
rect 866 1163 877 1164
rect 866 1159 867 1163
rect 871 1159 872 1163
rect 876 1159 877 1163
rect 928 1162 930 1164
rect 935 1163 941 1164
rect 935 1162 936 1163
rect 928 1160 936 1162
rect 866 1158 877 1159
rect 935 1159 936 1160
rect 940 1159 941 1163
rect 992 1162 994 1164
rect 999 1163 1005 1164
rect 999 1162 1000 1163
rect 992 1160 1000 1162
rect 935 1158 941 1159
rect 999 1159 1000 1160
rect 1004 1159 1005 1163
rect 999 1158 1005 1159
rect 1055 1163 1061 1164
rect 1055 1159 1056 1163
rect 1060 1162 1061 1163
rect 1099 1162 1101 1164
rect 1060 1160 1101 1162
rect 1119 1163 1125 1164
rect 1060 1159 1061 1160
rect 1055 1158 1061 1159
rect 1119 1159 1120 1163
rect 1124 1162 1125 1163
rect 1152 1162 1154 1164
rect 1124 1160 1154 1162
rect 1183 1163 1189 1164
rect 1124 1159 1125 1160
rect 1119 1158 1125 1159
rect 1183 1159 1184 1163
rect 1188 1162 1189 1163
rect 1220 1162 1222 1164
rect 1188 1160 1222 1162
rect 1255 1163 1261 1164
rect 1188 1159 1189 1160
rect 1183 1158 1189 1159
rect 1255 1159 1256 1163
rect 1260 1162 1261 1163
rect 1292 1162 1294 1164
rect 1260 1160 1294 1162
rect 1327 1163 1333 1164
rect 1260 1159 1261 1160
rect 1255 1158 1261 1159
rect 1327 1159 1328 1163
rect 1332 1162 1333 1163
rect 1368 1162 1370 1164
rect 1332 1160 1370 1162
rect 1407 1163 1413 1164
rect 1332 1159 1333 1160
rect 1327 1158 1333 1159
rect 1407 1159 1408 1163
rect 1412 1162 1413 1163
rect 1418 1163 1424 1164
rect 1418 1162 1419 1163
rect 1412 1160 1419 1162
rect 1412 1159 1413 1160
rect 1407 1158 1413 1159
rect 1418 1159 1419 1160
rect 1423 1159 1424 1163
rect 1489 1162 1491 1186
rect 1494 1179 1501 1180
rect 1494 1175 1495 1179
rect 1500 1175 1501 1179
rect 1559 1179 1565 1180
rect 1494 1174 1501 1175
rect 1542 1175 1548 1176
rect 1542 1171 1543 1175
rect 1547 1171 1548 1175
rect 1559 1175 1560 1179
rect 1564 1178 1565 1179
rect 1567 1179 1573 1180
rect 1567 1178 1568 1179
rect 1564 1176 1568 1178
rect 1564 1175 1565 1176
rect 1559 1174 1565 1175
rect 1567 1175 1568 1176
rect 1572 1175 1573 1179
rect 1567 1174 1573 1175
rect 1582 1176 1588 1177
rect 1582 1172 1583 1176
rect 1587 1172 1588 1176
rect 1582 1171 1588 1172
rect 1542 1170 1548 1171
rect 1495 1163 1501 1164
rect 1495 1162 1496 1163
rect 1489 1160 1496 1162
rect 1418 1158 1424 1159
rect 1495 1159 1496 1160
rect 1500 1159 1501 1163
rect 1495 1158 1501 1159
rect 1558 1163 1565 1164
rect 1558 1159 1559 1163
rect 1564 1159 1565 1163
rect 1558 1158 1565 1159
rect 1582 1159 1588 1160
rect 718 1157 724 1158
rect 718 1153 719 1157
rect 723 1153 724 1157
rect 718 1152 724 1153
rect 790 1157 796 1158
rect 790 1153 791 1157
rect 795 1153 796 1157
rect 790 1152 796 1153
rect 854 1157 860 1158
rect 854 1153 855 1157
rect 859 1153 860 1157
rect 854 1152 860 1153
rect 918 1157 924 1158
rect 918 1153 919 1157
rect 923 1153 924 1157
rect 918 1152 924 1153
rect 982 1157 988 1158
rect 982 1153 983 1157
rect 987 1153 988 1157
rect 982 1152 988 1153
rect 1038 1157 1044 1158
rect 1038 1153 1039 1157
rect 1043 1153 1044 1157
rect 1038 1152 1044 1153
rect 1102 1157 1108 1158
rect 1102 1153 1103 1157
rect 1107 1153 1108 1157
rect 1102 1152 1108 1153
rect 1166 1157 1172 1158
rect 1166 1153 1167 1157
rect 1171 1153 1172 1157
rect 1166 1152 1172 1153
rect 1238 1157 1244 1158
rect 1238 1153 1239 1157
rect 1243 1153 1244 1157
rect 1238 1152 1244 1153
rect 1310 1157 1316 1158
rect 1310 1153 1311 1157
rect 1315 1153 1316 1157
rect 1310 1152 1316 1153
rect 1390 1157 1396 1158
rect 1390 1153 1391 1157
rect 1395 1153 1396 1157
rect 1390 1152 1396 1153
rect 1478 1157 1484 1158
rect 1478 1153 1479 1157
rect 1483 1153 1484 1157
rect 1478 1152 1484 1153
rect 1542 1157 1548 1158
rect 1542 1153 1543 1157
rect 1547 1153 1548 1157
rect 1582 1155 1583 1159
rect 1587 1155 1588 1159
rect 1582 1154 1588 1155
rect 1542 1152 1548 1153
rect 523 1148 666 1150
rect 874 1151 880 1152
rect 523 1147 524 1148
rect 518 1146 524 1147
rect 874 1147 875 1151
rect 879 1150 880 1151
rect 1226 1151 1232 1152
rect 879 1148 1058 1150
rect 879 1147 880 1148
rect 874 1146 880 1147
rect 502 1143 508 1144
rect 502 1139 503 1143
rect 507 1139 508 1143
rect 502 1138 508 1139
rect 558 1143 564 1144
rect 558 1139 559 1143
rect 563 1139 564 1143
rect 558 1138 564 1139
rect 614 1143 620 1144
rect 614 1139 615 1143
rect 619 1139 620 1143
rect 614 1138 620 1139
rect 670 1143 676 1144
rect 670 1139 671 1143
rect 675 1139 676 1143
rect 670 1138 676 1139
rect 726 1143 732 1144
rect 726 1139 727 1143
rect 731 1139 732 1143
rect 726 1138 732 1139
rect 782 1143 788 1144
rect 782 1139 783 1143
rect 787 1139 788 1143
rect 782 1138 788 1139
rect 838 1143 844 1144
rect 838 1139 839 1143
rect 843 1139 844 1143
rect 838 1138 844 1139
rect 894 1143 900 1144
rect 894 1139 895 1143
rect 899 1139 900 1143
rect 894 1138 900 1139
rect 950 1143 956 1144
rect 950 1139 951 1143
rect 955 1139 956 1143
rect 950 1138 956 1139
rect 1006 1143 1012 1144
rect 1006 1139 1007 1143
rect 1011 1139 1012 1143
rect 1006 1138 1012 1139
rect 519 1135 525 1136
rect 519 1134 520 1135
rect 468 1132 494 1134
rect 496 1132 520 1134
rect 468 1131 469 1132
rect 463 1130 469 1131
rect 446 1125 452 1126
rect 446 1121 447 1125
rect 451 1121 452 1125
rect 446 1120 452 1121
rect 463 1119 469 1120
rect 463 1118 464 1119
rect 436 1116 464 1118
rect 407 1114 413 1115
rect 463 1115 464 1116
rect 468 1115 469 1119
rect 492 1118 494 1132
rect 519 1131 520 1132
rect 524 1131 525 1135
rect 519 1130 525 1131
rect 575 1135 581 1136
rect 575 1131 576 1135
rect 580 1134 581 1135
rect 631 1135 637 1136
rect 580 1132 626 1134
rect 580 1131 581 1132
rect 575 1130 581 1131
rect 502 1125 508 1126
rect 502 1121 503 1125
rect 507 1121 508 1125
rect 502 1120 508 1121
rect 558 1125 564 1126
rect 558 1121 559 1125
rect 563 1121 564 1125
rect 558 1120 564 1121
rect 614 1125 620 1126
rect 614 1121 615 1125
rect 619 1121 620 1125
rect 614 1120 620 1121
rect 519 1119 525 1120
rect 519 1118 520 1119
rect 492 1116 520 1118
rect 463 1114 469 1115
rect 519 1115 520 1116
rect 524 1115 525 1119
rect 519 1114 525 1115
rect 575 1119 581 1120
rect 575 1115 576 1119
rect 580 1118 581 1119
rect 606 1119 612 1120
rect 606 1118 607 1119
rect 580 1116 607 1118
rect 580 1115 581 1116
rect 575 1114 581 1115
rect 606 1115 607 1116
rect 611 1115 612 1119
rect 624 1118 626 1132
rect 631 1131 632 1135
rect 636 1134 637 1135
rect 687 1135 693 1136
rect 636 1132 662 1134
rect 636 1131 637 1132
rect 631 1130 637 1131
rect 631 1119 637 1120
rect 631 1118 632 1119
rect 624 1116 632 1118
rect 606 1114 612 1115
rect 631 1115 632 1116
rect 636 1115 637 1119
rect 660 1118 662 1132
rect 687 1131 688 1135
rect 692 1134 693 1135
rect 743 1135 749 1136
rect 692 1132 718 1134
rect 692 1131 693 1132
rect 687 1130 693 1131
rect 670 1125 676 1126
rect 670 1121 671 1125
rect 675 1121 676 1125
rect 670 1120 676 1121
rect 687 1119 693 1120
rect 687 1118 688 1119
rect 660 1116 688 1118
rect 631 1114 637 1115
rect 687 1115 688 1116
rect 692 1115 693 1119
rect 716 1118 718 1132
rect 743 1131 744 1135
rect 748 1134 749 1135
rect 799 1135 808 1136
rect 748 1132 774 1134
rect 748 1131 749 1132
rect 743 1130 749 1131
rect 726 1125 732 1126
rect 726 1121 727 1125
rect 731 1121 732 1125
rect 726 1120 732 1121
rect 743 1119 749 1120
rect 743 1118 744 1119
rect 716 1116 744 1118
rect 687 1114 693 1115
rect 743 1115 744 1116
rect 748 1115 749 1119
rect 772 1118 774 1132
rect 799 1131 800 1135
rect 807 1131 808 1135
rect 799 1130 808 1131
rect 855 1135 861 1136
rect 855 1131 856 1135
rect 860 1134 861 1135
rect 911 1135 917 1136
rect 860 1132 886 1134
rect 860 1131 861 1132
rect 855 1130 861 1131
rect 782 1125 788 1126
rect 782 1121 783 1125
rect 787 1121 788 1125
rect 782 1120 788 1121
rect 838 1125 844 1126
rect 838 1121 839 1125
rect 843 1121 844 1125
rect 838 1120 844 1121
rect 799 1119 805 1120
rect 799 1118 800 1119
rect 772 1116 800 1118
rect 743 1114 749 1115
rect 799 1115 800 1116
rect 804 1115 805 1119
rect 799 1114 805 1115
rect 855 1119 861 1120
rect 855 1115 856 1119
rect 860 1118 861 1119
rect 866 1119 872 1120
rect 866 1118 867 1119
rect 860 1116 867 1118
rect 860 1115 861 1116
rect 855 1114 861 1115
rect 866 1115 867 1116
rect 871 1115 872 1119
rect 884 1118 886 1132
rect 911 1131 912 1135
rect 916 1134 917 1135
rect 967 1135 973 1136
rect 916 1132 942 1134
rect 916 1131 917 1132
rect 911 1130 917 1131
rect 894 1125 900 1126
rect 894 1121 895 1125
rect 899 1121 900 1125
rect 894 1120 900 1121
rect 911 1119 917 1120
rect 911 1118 912 1119
rect 884 1116 912 1118
rect 866 1114 872 1115
rect 911 1115 912 1116
rect 916 1115 917 1119
rect 940 1118 942 1132
rect 967 1131 968 1135
rect 972 1134 973 1135
rect 1023 1135 1029 1136
rect 972 1132 1018 1134
rect 972 1131 973 1132
rect 967 1130 973 1131
rect 950 1125 956 1126
rect 950 1121 951 1125
rect 955 1121 956 1125
rect 950 1120 956 1121
rect 1006 1125 1012 1126
rect 1006 1121 1007 1125
rect 1011 1121 1012 1125
rect 1006 1120 1012 1121
rect 967 1119 973 1120
rect 967 1118 968 1119
rect 940 1116 968 1118
rect 911 1114 917 1115
rect 967 1115 968 1116
rect 972 1115 973 1119
rect 1016 1118 1018 1132
rect 1023 1131 1024 1135
rect 1028 1134 1029 1135
rect 1056 1134 1058 1148
rect 1226 1147 1227 1151
rect 1231 1150 1232 1151
rect 1231 1148 1386 1150
rect 1231 1147 1232 1148
rect 1226 1146 1232 1147
rect 1062 1143 1068 1144
rect 1062 1139 1063 1143
rect 1067 1139 1068 1143
rect 1062 1138 1068 1139
rect 1126 1143 1132 1144
rect 1126 1139 1127 1143
rect 1131 1139 1132 1143
rect 1126 1138 1132 1139
rect 1190 1143 1196 1144
rect 1190 1139 1191 1143
rect 1195 1139 1196 1143
rect 1190 1138 1196 1139
rect 1254 1143 1260 1144
rect 1254 1139 1255 1143
rect 1259 1139 1260 1143
rect 1254 1138 1260 1139
rect 1326 1143 1332 1144
rect 1326 1139 1327 1143
rect 1331 1139 1332 1143
rect 1326 1138 1332 1139
rect 1079 1135 1085 1136
rect 1079 1134 1080 1135
rect 1028 1132 1054 1134
rect 1056 1132 1080 1134
rect 1028 1131 1029 1132
rect 1023 1130 1029 1131
rect 1023 1119 1029 1120
rect 1023 1118 1024 1119
rect 1016 1116 1024 1118
rect 967 1114 973 1115
rect 1023 1115 1024 1116
rect 1028 1115 1029 1119
rect 1052 1118 1054 1132
rect 1079 1131 1080 1132
rect 1084 1131 1085 1135
rect 1079 1130 1085 1131
rect 1143 1135 1149 1136
rect 1143 1131 1144 1135
rect 1148 1134 1149 1135
rect 1207 1135 1213 1136
rect 1148 1132 1178 1134
rect 1148 1131 1149 1132
rect 1143 1130 1149 1131
rect 1062 1125 1068 1126
rect 1062 1121 1063 1125
rect 1067 1121 1068 1125
rect 1062 1120 1068 1121
rect 1126 1125 1132 1126
rect 1126 1121 1127 1125
rect 1131 1121 1132 1125
rect 1126 1120 1132 1121
rect 1079 1119 1085 1120
rect 1079 1118 1080 1119
rect 1052 1116 1080 1118
rect 1023 1114 1029 1115
rect 1079 1115 1080 1116
rect 1084 1115 1085 1119
rect 1079 1114 1085 1115
rect 1143 1119 1149 1120
rect 1143 1115 1144 1119
rect 1148 1118 1149 1119
rect 1158 1119 1164 1120
rect 1158 1118 1159 1119
rect 1148 1116 1159 1118
rect 1148 1115 1149 1116
rect 1143 1114 1149 1115
rect 1158 1115 1159 1116
rect 1163 1115 1164 1119
rect 1176 1118 1178 1132
rect 1207 1131 1208 1135
rect 1212 1134 1213 1135
rect 1271 1135 1277 1136
rect 1212 1132 1266 1134
rect 1212 1131 1213 1132
rect 1207 1130 1213 1131
rect 1190 1125 1196 1126
rect 1190 1121 1191 1125
rect 1195 1121 1196 1125
rect 1190 1120 1196 1121
rect 1254 1125 1260 1126
rect 1254 1121 1255 1125
rect 1259 1121 1260 1125
rect 1254 1120 1260 1121
rect 1207 1119 1213 1120
rect 1207 1118 1208 1119
rect 1176 1116 1208 1118
rect 1158 1114 1164 1115
rect 1207 1115 1208 1116
rect 1212 1115 1213 1119
rect 1264 1118 1266 1132
rect 1271 1131 1272 1135
rect 1276 1134 1277 1135
rect 1343 1135 1349 1136
rect 1276 1132 1310 1134
rect 1276 1131 1277 1132
rect 1271 1130 1277 1131
rect 1271 1119 1277 1120
rect 1271 1118 1272 1119
rect 1264 1116 1272 1118
rect 1207 1114 1213 1115
rect 1271 1115 1272 1116
rect 1276 1115 1277 1119
rect 1308 1118 1310 1132
rect 1343 1131 1344 1135
rect 1348 1134 1349 1135
rect 1384 1134 1386 1148
rect 1398 1143 1404 1144
rect 1398 1139 1399 1143
rect 1403 1139 1404 1143
rect 1398 1138 1404 1139
rect 1478 1143 1484 1144
rect 1478 1139 1479 1143
rect 1483 1139 1484 1143
rect 1478 1138 1484 1139
rect 1542 1143 1548 1144
rect 1542 1139 1543 1143
rect 1547 1139 1548 1143
rect 1542 1138 1548 1139
rect 1582 1141 1588 1142
rect 1582 1137 1583 1141
rect 1587 1137 1588 1141
rect 1582 1136 1588 1137
rect 1415 1135 1421 1136
rect 1415 1134 1416 1135
rect 1348 1132 1382 1134
rect 1384 1132 1416 1134
rect 1348 1131 1349 1132
rect 1343 1130 1349 1131
rect 1326 1125 1332 1126
rect 1326 1121 1327 1125
rect 1331 1121 1332 1125
rect 1326 1120 1332 1121
rect 1343 1119 1349 1120
rect 1343 1118 1344 1119
rect 1308 1116 1344 1118
rect 1271 1114 1277 1115
rect 1343 1115 1344 1116
rect 1348 1115 1349 1119
rect 1380 1118 1382 1132
rect 1415 1131 1416 1132
rect 1420 1131 1421 1135
rect 1415 1130 1421 1131
rect 1494 1135 1501 1136
rect 1494 1131 1495 1135
rect 1500 1131 1501 1135
rect 1494 1130 1501 1131
rect 1559 1135 1565 1136
rect 1559 1131 1560 1135
rect 1564 1134 1565 1135
rect 1567 1135 1573 1136
rect 1567 1134 1568 1135
rect 1564 1132 1568 1134
rect 1564 1131 1565 1132
rect 1559 1130 1565 1131
rect 1567 1131 1568 1132
rect 1572 1131 1573 1135
rect 1567 1130 1573 1131
rect 1398 1125 1404 1126
rect 1398 1121 1399 1125
rect 1403 1121 1404 1125
rect 1398 1120 1404 1121
rect 1478 1125 1484 1126
rect 1478 1121 1479 1125
rect 1483 1121 1484 1125
rect 1478 1120 1484 1121
rect 1542 1125 1548 1126
rect 1542 1121 1543 1125
rect 1547 1121 1548 1125
rect 1542 1120 1548 1121
rect 1582 1124 1588 1125
rect 1582 1120 1583 1124
rect 1587 1120 1588 1124
rect 1415 1119 1421 1120
rect 1415 1118 1416 1119
rect 1380 1116 1416 1118
rect 1343 1114 1349 1115
rect 1415 1115 1416 1116
rect 1420 1115 1421 1119
rect 1415 1114 1421 1115
rect 1495 1119 1501 1120
rect 1495 1115 1496 1119
rect 1500 1118 1501 1119
rect 1518 1119 1524 1120
rect 1518 1118 1519 1119
rect 1500 1116 1519 1118
rect 1500 1115 1501 1116
rect 1495 1114 1501 1115
rect 1518 1115 1519 1116
rect 1523 1115 1524 1119
rect 1518 1114 1524 1115
rect 1558 1119 1565 1120
rect 1582 1119 1588 1120
rect 1558 1115 1559 1119
rect 1564 1115 1565 1119
rect 1558 1114 1565 1115
rect 1410 1111 1416 1112
rect 167 1107 173 1108
rect 110 1104 116 1105
rect 167 1104 168 1107
rect 110 1100 111 1104
rect 115 1100 116 1104
rect 110 1099 116 1100
rect 150 1103 156 1104
rect 150 1099 151 1103
rect 155 1099 156 1103
rect 150 1098 156 1099
rect 166 1103 168 1104
rect 172 1103 173 1107
rect 199 1107 205 1108
rect 199 1106 200 1107
rect 192 1104 200 1106
rect 166 1099 167 1103
rect 171 1102 173 1103
rect 182 1103 188 1104
rect 171 1099 172 1102
rect 166 1098 172 1099
rect 182 1099 183 1103
rect 187 1099 188 1103
rect 182 1098 188 1099
rect 192 1094 194 1104
rect 199 1103 200 1104
rect 204 1103 205 1107
rect 239 1107 245 1108
rect 239 1106 240 1107
rect 232 1104 240 1106
rect 199 1102 205 1103
rect 222 1103 228 1104
rect 222 1099 223 1103
rect 227 1099 228 1103
rect 222 1098 228 1099
rect 232 1094 234 1104
rect 239 1103 240 1104
rect 244 1103 245 1107
rect 287 1107 293 1108
rect 287 1106 288 1107
rect 280 1104 288 1106
rect 239 1102 245 1103
rect 270 1103 276 1104
rect 270 1099 271 1103
rect 275 1099 276 1103
rect 270 1098 276 1099
rect 280 1094 282 1104
rect 287 1103 288 1104
rect 292 1103 293 1107
rect 343 1107 349 1108
rect 343 1106 344 1107
rect 336 1104 344 1106
rect 287 1102 293 1103
rect 326 1103 332 1104
rect 326 1099 327 1103
rect 331 1099 332 1103
rect 326 1098 332 1099
rect 336 1094 338 1104
rect 343 1103 344 1104
rect 348 1103 349 1107
rect 399 1107 405 1108
rect 399 1106 400 1107
rect 392 1104 400 1106
rect 343 1102 349 1103
rect 382 1103 388 1104
rect 382 1099 383 1103
rect 387 1099 388 1103
rect 382 1098 388 1099
rect 392 1094 394 1104
rect 399 1103 400 1104
rect 404 1103 405 1107
rect 455 1107 461 1108
rect 399 1102 405 1103
rect 438 1103 444 1104
rect 438 1099 439 1103
rect 443 1099 444 1103
rect 455 1103 456 1107
rect 460 1106 461 1107
rect 494 1107 500 1108
rect 494 1106 495 1107
rect 460 1104 495 1106
rect 460 1103 461 1104
rect 455 1102 461 1103
rect 494 1103 495 1104
rect 499 1103 500 1107
rect 519 1107 525 1108
rect 519 1106 520 1107
rect 512 1104 520 1106
rect 494 1102 500 1103
rect 502 1103 508 1104
rect 438 1098 444 1099
rect 502 1099 503 1103
rect 507 1099 508 1103
rect 502 1098 508 1099
rect 512 1094 514 1104
rect 519 1103 520 1104
rect 524 1103 525 1107
rect 583 1107 589 1108
rect 583 1106 584 1107
rect 576 1104 584 1106
rect 519 1102 525 1103
rect 566 1103 572 1104
rect 566 1099 567 1103
rect 571 1099 572 1103
rect 566 1098 572 1099
rect 576 1094 578 1104
rect 583 1103 584 1104
rect 588 1103 589 1107
rect 655 1107 661 1108
rect 655 1106 656 1107
rect 648 1104 656 1106
rect 583 1102 589 1103
rect 638 1103 644 1104
rect 638 1099 639 1103
rect 643 1099 644 1103
rect 638 1098 644 1099
rect 648 1094 650 1104
rect 655 1103 656 1104
rect 660 1103 661 1107
rect 727 1107 733 1108
rect 727 1106 728 1107
rect 720 1104 728 1106
rect 655 1102 661 1103
rect 710 1103 716 1104
rect 710 1099 711 1103
rect 715 1099 716 1103
rect 710 1098 716 1099
rect 720 1094 722 1104
rect 727 1103 728 1104
rect 732 1103 733 1107
rect 799 1107 805 1108
rect 799 1106 800 1107
rect 792 1104 800 1106
rect 727 1102 733 1103
rect 782 1103 788 1104
rect 782 1099 783 1103
rect 787 1099 788 1103
rect 782 1098 788 1099
rect 792 1094 794 1104
rect 799 1103 800 1104
rect 804 1103 805 1107
rect 871 1107 880 1108
rect 799 1102 805 1103
rect 854 1103 860 1104
rect 854 1099 855 1103
rect 859 1099 860 1103
rect 871 1103 872 1107
rect 879 1103 880 1107
rect 935 1107 941 1108
rect 935 1106 936 1107
rect 928 1104 936 1106
rect 871 1102 880 1103
rect 918 1103 924 1104
rect 854 1098 860 1099
rect 918 1099 919 1103
rect 923 1099 924 1103
rect 918 1098 924 1099
rect 928 1094 930 1104
rect 935 1103 936 1104
rect 940 1103 941 1107
rect 999 1107 1005 1108
rect 999 1106 1000 1107
rect 992 1104 1000 1106
rect 935 1102 941 1103
rect 982 1103 988 1104
rect 982 1099 983 1103
rect 987 1099 988 1103
rect 982 1098 988 1099
rect 992 1094 994 1104
rect 999 1103 1000 1104
rect 1004 1103 1005 1107
rect 1055 1107 1061 1108
rect 1055 1106 1056 1107
rect 1048 1104 1056 1106
rect 999 1102 1005 1103
rect 1038 1103 1044 1104
rect 1038 1099 1039 1103
rect 1043 1099 1044 1103
rect 1038 1098 1044 1099
rect 1048 1094 1050 1104
rect 1055 1103 1056 1104
rect 1060 1103 1061 1107
rect 1111 1107 1117 1108
rect 1111 1106 1112 1107
rect 1104 1104 1112 1106
rect 1055 1102 1061 1103
rect 1094 1103 1100 1104
rect 1094 1099 1095 1103
rect 1099 1099 1100 1103
rect 1094 1098 1100 1099
rect 1104 1094 1106 1104
rect 1111 1103 1112 1104
rect 1116 1103 1117 1107
rect 1167 1107 1173 1108
rect 1167 1106 1168 1107
rect 1160 1104 1168 1106
rect 1111 1102 1117 1103
rect 1150 1103 1156 1104
rect 1150 1099 1151 1103
rect 1155 1099 1156 1103
rect 1150 1098 1156 1099
rect 1160 1094 1162 1104
rect 1167 1103 1168 1104
rect 1172 1103 1173 1107
rect 1223 1107 1232 1108
rect 1167 1102 1173 1103
rect 1206 1103 1212 1104
rect 1206 1099 1207 1103
rect 1211 1099 1212 1103
rect 1223 1103 1224 1107
rect 1231 1103 1232 1107
rect 1279 1107 1285 1108
rect 1279 1106 1280 1107
rect 1272 1104 1280 1106
rect 1223 1102 1232 1103
rect 1262 1103 1268 1104
rect 1206 1098 1212 1099
rect 1262 1099 1263 1103
rect 1267 1099 1268 1103
rect 1262 1098 1268 1099
rect 1272 1094 1274 1104
rect 1279 1103 1280 1104
rect 1284 1103 1285 1107
rect 1335 1107 1341 1108
rect 1335 1106 1336 1107
rect 1328 1104 1336 1106
rect 1279 1102 1285 1103
rect 1318 1103 1324 1104
rect 1318 1099 1319 1103
rect 1323 1099 1324 1103
rect 1318 1098 1324 1099
rect 1328 1094 1330 1104
rect 1335 1103 1336 1104
rect 1340 1103 1341 1107
rect 1391 1107 1397 1108
rect 1391 1106 1392 1107
rect 1384 1104 1392 1106
rect 1335 1102 1341 1103
rect 1374 1103 1380 1104
rect 1374 1099 1375 1103
rect 1379 1099 1380 1103
rect 1374 1098 1380 1099
rect 1384 1094 1386 1104
rect 1391 1103 1392 1104
rect 1396 1103 1397 1107
rect 1410 1107 1411 1111
rect 1415 1110 1416 1111
rect 1415 1108 1450 1110
rect 1415 1107 1416 1108
rect 1410 1106 1416 1107
rect 1448 1106 1450 1108
rect 1455 1107 1461 1108
rect 1455 1106 1456 1107
rect 1448 1104 1456 1106
rect 1391 1102 1397 1103
rect 1438 1103 1444 1104
rect 1438 1099 1439 1103
rect 1443 1099 1444 1103
rect 1455 1103 1456 1104
rect 1460 1103 1461 1107
rect 1519 1107 1525 1108
rect 1519 1106 1520 1107
rect 1512 1104 1520 1106
rect 1455 1102 1461 1103
rect 1502 1103 1508 1104
rect 1438 1098 1444 1099
rect 1502 1099 1503 1103
rect 1507 1099 1508 1103
rect 1502 1098 1508 1099
rect 1512 1094 1514 1104
rect 1519 1103 1520 1104
rect 1524 1103 1525 1107
rect 1559 1107 1565 1108
rect 1519 1102 1525 1103
rect 1542 1103 1548 1104
rect 1542 1099 1543 1103
rect 1547 1099 1548 1103
rect 1559 1103 1560 1107
rect 1564 1106 1565 1107
rect 1567 1107 1573 1108
rect 1567 1106 1568 1107
rect 1564 1104 1568 1106
rect 1564 1103 1565 1104
rect 1559 1102 1565 1103
rect 1567 1103 1568 1104
rect 1572 1103 1573 1107
rect 1567 1102 1573 1103
rect 1582 1104 1588 1105
rect 1582 1100 1583 1104
rect 1587 1100 1588 1104
rect 1582 1099 1588 1100
rect 1542 1098 1548 1099
rect 180 1092 194 1094
rect 220 1092 234 1094
rect 259 1092 282 1094
rect 289 1092 338 1094
rect 372 1092 394 1094
rect 489 1092 514 1094
rect 552 1092 578 1094
rect 620 1092 650 1094
rect 692 1092 722 1094
rect 764 1092 794 1094
rect 873 1092 930 1094
rect 937 1092 994 1094
rect 1001 1092 1050 1094
rect 1057 1092 1106 1094
rect 1140 1092 1162 1094
rect 1252 1092 1274 1094
rect 1308 1092 1330 1094
rect 1364 1092 1386 1094
rect 1459 1092 1514 1094
rect 167 1091 173 1092
rect 110 1087 116 1088
rect 110 1083 111 1087
rect 115 1083 116 1087
rect 167 1087 168 1091
rect 172 1090 173 1091
rect 180 1090 182 1092
rect 172 1088 182 1090
rect 199 1091 205 1092
rect 172 1087 173 1088
rect 167 1086 173 1087
rect 199 1087 200 1091
rect 204 1090 205 1091
rect 220 1090 222 1092
rect 204 1088 222 1090
rect 239 1091 245 1092
rect 204 1087 205 1088
rect 199 1086 205 1087
rect 239 1087 240 1091
rect 244 1090 245 1091
rect 259 1090 261 1092
rect 244 1088 261 1090
rect 287 1091 293 1092
rect 244 1087 245 1088
rect 239 1086 245 1087
rect 287 1087 288 1091
rect 292 1087 293 1091
rect 287 1086 293 1087
rect 343 1091 349 1092
rect 343 1087 344 1091
rect 348 1090 349 1091
rect 372 1090 374 1092
rect 399 1091 405 1092
rect 399 1090 400 1091
rect 348 1088 374 1090
rect 392 1088 400 1090
rect 348 1087 349 1088
rect 343 1086 349 1087
rect 110 1082 116 1083
rect 150 1085 156 1086
rect 150 1081 151 1085
rect 155 1081 156 1085
rect 150 1080 156 1081
rect 182 1085 188 1086
rect 182 1081 183 1085
rect 187 1081 188 1085
rect 182 1080 188 1081
rect 222 1085 228 1086
rect 222 1081 223 1085
rect 227 1081 228 1085
rect 222 1080 228 1081
rect 270 1085 276 1086
rect 270 1081 271 1085
rect 275 1081 276 1085
rect 270 1080 276 1081
rect 326 1085 332 1086
rect 326 1081 327 1085
rect 331 1081 332 1085
rect 326 1080 332 1081
rect 382 1085 388 1086
rect 382 1081 383 1085
rect 387 1081 388 1085
rect 382 1080 388 1081
rect 346 1079 352 1080
rect 346 1075 347 1079
rect 351 1078 352 1079
rect 392 1078 394 1088
rect 399 1087 400 1088
rect 404 1087 405 1091
rect 399 1086 405 1087
rect 455 1091 461 1092
rect 455 1087 456 1091
rect 460 1090 461 1091
rect 489 1090 491 1092
rect 460 1088 491 1090
rect 519 1091 525 1092
rect 460 1087 461 1088
rect 455 1086 461 1087
rect 519 1087 520 1091
rect 524 1090 525 1091
rect 552 1090 554 1092
rect 524 1088 554 1090
rect 583 1091 589 1092
rect 524 1087 525 1088
rect 519 1086 525 1087
rect 583 1087 584 1091
rect 588 1090 589 1091
rect 620 1090 622 1092
rect 588 1088 622 1090
rect 655 1091 661 1092
rect 588 1087 589 1088
rect 583 1086 589 1087
rect 655 1087 656 1091
rect 660 1090 661 1091
rect 692 1090 694 1092
rect 660 1088 694 1090
rect 727 1091 733 1092
rect 660 1087 661 1088
rect 655 1086 661 1087
rect 727 1087 728 1091
rect 732 1090 733 1091
rect 764 1090 766 1092
rect 799 1091 805 1092
rect 799 1090 800 1091
rect 732 1088 766 1090
rect 792 1088 800 1090
rect 732 1087 733 1088
rect 727 1086 733 1087
rect 438 1085 444 1086
rect 438 1081 439 1085
rect 443 1081 444 1085
rect 438 1080 444 1081
rect 502 1085 508 1086
rect 502 1081 503 1085
rect 507 1081 508 1085
rect 502 1080 508 1081
rect 566 1085 572 1086
rect 566 1081 567 1085
rect 571 1081 572 1085
rect 566 1080 572 1081
rect 638 1085 644 1086
rect 638 1081 639 1085
rect 643 1081 644 1085
rect 638 1080 644 1081
rect 710 1085 716 1086
rect 710 1081 711 1085
rect 715 1081 716 1085
rect 710 1080 716 1081
rect 782 1085 788 1086
rect 782 1081 783 1085
rect 787 1081 788 1085
rect 782 1080 788 1081
rect 351 1076 394 1078
rect 606 1079 612 1080
rect 351 1075 352 1076
rect 346 1074 352 1075
rect 606 1075 607 1079
rect 611 1078 612 1079
rect 792 1078 794 1088
rect 799 1087 800 1088
rect 804 1087 805 1091
rect 799 1086 805 1087
rect 871 1091 877 1092
rect 871 1087 872 1091
rect 876 1087 877 1091
rect 871 1086 877 1087
rect 935 1091 941 1092
rect 935 1087 936 1091
rect 940 1087 941 1091
rect 935 1086 941 1087
rect 999 1091 1005 1092
rect 999 1087 1000 1091
rect 1004 1087 1005 1091
rect 999 1086 1005 1087
rect 1055 1091 1061 1092
rect 1055 1087 1056 1091
rect 1060 1087 1061 1091
rect 1055 1086 1061 1087
rect 1111 1091 1117 1092
rect 1111 1087 1112 1091
rect 1116 1090 1117 1091
rect 1140 1090 1142 1092
rect 1116 1088 1142 1090
rect 1166 1091 1173 1092
rect 1116 1087 1117 1088
rect 1111 1086 1117 1087
rect 1166 1087 1167 1091
rect 1172 1087 1173 1091
rect 1166 1086 1173 1087
rect 1223 1091 1229 1092
rect 1223 1087 1224 1091
rect 1228 1090 1229 1091
rect 1252 1090 1254 1092
rect 1228 1088 1254 1090
rect 1279 1091 1285 1092
rect 1228 1087 1229 1088
rect 1223 1086 1229 1087
rect 1279 1087 1280 1091
rect 1284 1090 1285 1091
rect 1308 1090 1310 1092
rect 1284 1088 1310 1090
rect 1335 1091 1341 1092
rect 1284 1087 1285 1088
rect 1279 1086 1285 1087
rect 1335 1087 1336 1091
rect 1340 1090 1341 1091
rect 1364 1090 1366 1092
rect 1340 1088 1366 1090
rect 1390 1091 1397 1092
rect 1340 1087 1341 1088
rect 1335 1086 1341 1087
rect 1390 1087 1391 1091
rect 1396 1087 1397 1091
rect 1390 1086 1397 1087
rect 1455 1091 1461 1092
rect 1455 1087 1456 1091
rect 1460 1087 1461 1091
rect 1455 1086 1461 1087
rect 1518 1091 1525 1092
rect 1518 1087 1519 1091
rect 1524 1087 1525 1091
rect 1518 1086 1525 1087
rect 1558 1091 1565 1092
rect 1558 1087 1559 1091
rect 1564 1087 1565 1091
rect 1558 1086 1565 1087
rect 1582 1087 1588 1088
rect 854 1085 860 1086
rect 854 1081 855 1085
rect 859 1081 860 1085
rect 854 1080 860 1081
rect 918 1085 924 1086
rect 918 1081 919 1085
rect 923 1081 924 1085
rect 918 1080 924 1081
rect 982 1085 988 1086
rect 982 1081 983 1085
rect 987 1081 988 1085
rect 982 1080 988 1081
rect 1038 1085 1044 1086
rect 1038 1081 1039 1085
rect 1043 1081 1044 1085
rect 1038 1080 1044 1081
rect 1094 1085 1100 1086
rect 1094 1081 1095 1085
rect 1099 1081 1100 1085
rect 1094 1080 1100 1081
rect 1150 1085 1156 1086
rect 1150 1081 1151 1085
rect 1155 1081 1156 1085
rect 1150 1080 1156 1081
rect 1206 1085 1212 1086
rect 1206 1081 1207 1085
rect 1211 1081 1212 1085
rect 1206 1080 1212 1081
rect 1262 1085 1268 1086
rect 1262 1081 1263 1085
rect 1267 1081 1268 1085
rect 1262 1080 1268 1081
rect 1318 1085 1324 1086
rect 1318 1081 1319 1085
rect 1323 1081 1324 1085
rect 1318 1080 1324 1081
rect 1374 1085 1380 1086
rect 1374 1081 1375 1085
rect 1379 1081 1380 1085
rect 1374 1080 1380 1081
rect 1438 1085 1444 1086
rect 1438 1081 1439 1085
rect 1443 1081 1444 1085
rect 1438 1080 1444 1081
rect 1502 1085 1508 1086
rect 1502 1081 1503 1085
rect 1507 1081 1508 1085
rect 1502 1080 1508 1081
rect 1542 1085 1548 1086
rect 1542 1081 1543 1085
rect 1547 1081 1548 1085
rect 1582 1083 1583 1087
rect 1587 1083 1588 1087
rect 1582 1082 1588 1083
rect 1542 1080 1548 1081
rect 611 1076 794 1078
rect 1158 1079 1164 1080
rect 611 1075 612 1076
rect 606 1074 612 1075
rect 1158 1075 1159 1079
rect 1163 1078 1164 1079
rect 1418 1079 1424 1080
rect 1418 1078 1419 1079
rect 1163 1076 1419 1078
rect 1163 1075 1164 1076
rect 1158 1074 1164 1075
rect 1418 1075 1419 1076
rect 1423 1075 1424 1079
rect 1418 1074 1424 1075
rect 494 1071 500 1072
rect 494 1067 495 1071
rect 499 1070 500 1071
rect 499 1068 746 1070
rect 499 1067 500 1068
rect 494 1066 500 1067
rect 446 1063 452 1064
rect 110 1061 116 1062
rect 110 1057 111 1061
rect 115 1057 116 1061
rect 446 1059 447 1063
rect 451 1059 452 1063
rect 446 1058 452 1059
rect 486 1063 492 1064
rect 486 1059 487 1063
rect 491 1059 492 1063
rect 486 1058 492 1059
rect 542 1063 548 1064
rect 542 1059 543 1063
rect 547 1059 548 1063
rect 542 1058 548 1059
rect 598 1063 604 1064
rect 598 1059 599 1063
rect 603 1059 604 1063
rect 598 1058 604 1059
rect 662 1063 668 1064
rect 662 1059 663 1063
rect 667 1059 668 1063
rect 662 1058 668 1059
rect 726 1063 732 1064
rect 726 1059 727 1063
rect 731 1059 732 1063
rect 726 1058 732 1059
rect 110 1056 116 1057
rect 744 1056 746 1068
rect 790 1063 796 1064
rect 790 1059 791 1063
rect 795 1059 796 1063
rect 790 1058 796 1059
rect 862 1063 868 1064
rect 862 1059 863 1063
rect 867 1059 868 1063
rect 862 1058 868 1059
rect 934 1063 940 1064
rect 934 1059 935 1063
rect 939 1059 940 1063
rect 934 1058 940 1059
rect 1006 1063 1012 1064
rect 1006 1059 1007 1063
rect 1011 1059 1012 1063
rect 1006 1058 1012 1059
rect 1078 1063 1084 1064
rect 1078 1059 1079 1063
rect 1083 1059 1084 1063
rect 1078 1058 1084 1059
rect 1150 1063 1156 1064
rect 1150 1059 1151 1063
rect 1155 1059 1156 1063
rect 1150 1058 1156 1059
rect 1214 1063 1220 1064
rect 1214 1059 1215 1063
rect 1219 1059 1220 1063
rect 1214 1058 1220 1059
rect 1278 1063 1284 1064
rect 1278 1059 1279 1063
rect 1283 1059 1284 1063
rect 1278 1058 1284 1059
rect 1334 1063 1340 1064
rect 1334 1059 1335 1063
rect 1339 1059 1340 1063
rect 1334 1058 1340 1059
rect 1390 1063 1396 1064
rect 1390 1059 1391 1063
rect 1395 1059 1396 1063
rect 1390 1058 1396 1059
rect 1446 1063 1452 1064
rect 1446 1059 1447 1063
rect 1451 1059 1452 1063
rect 1446 1058 1452 1059
rect 1502 1063 1508 1064
rect 1502 1059 1503 1063
rect 1507 1059 1508 1063
rect 1502 1058 1508 1059
rect 1542 1063 1548 1064
rect 1542 1059 1543 1063
rect 1547 1059 1548 1063
rect 1542 1058 1548 1059
rect 1582 1061 1588 1062
rect 1582 1057 1583 1061
rect 1587 1057 1588 1061
rect 1582 1056 1588 1057
rect 463 1055 469 1056
rect 463 1051 464 1055
rect 468 1054 469 1055
rect 503 1055 509 1056
rect 468 1052 482 1054
rect 468 1051 469 1052
rect 463 1050 469 1051
rect 446 1045 452 1046
rect 110 1044 116 1045
rect 110 1040 111 1044
rect 115 1040 116 1044
rect 446 1041 447 1045
rect 451 1041 452 1045
rect 446 1040 452 1041
rect 110 1039 116 1040
rect 463 1039 469 1040
rect 463 1035 464 1039
rect 468 1038 469 1039
rect 471 1039 477 1040
rect 471 1038 472 1039
rect 468 1036 472 1038
rect 468 1035 469 1036
rect 463 1034 469 1035
rect 471 1035 472 1036
rect 476 1035 477 1039
rect 480 1038 482 1052
rect 503 1051 504 1055
rect 508 1054 509 1055
rect 559 1055 565 1056
rect 508 1052 534 1054
rect 508 1051 509 1052
rect 503 1050 509 1051
rect 486 1045 492 1046
rect 486 1041 487 1045
rect 491 1041 492 1045
rect 486 1040 492 1041
rect 503 1039 509 1040
rect 503 1038 504 1039
rect 480 1036 504 1038
rect 471 1034 477 1035
rect 503 1035 504 1036
rect 508 1035 509 1039
rect 532 1038 534 1052
rect 559 1051 560 1055
rect 564 1054 565 1055
rect 615 1055 621 1056
rect 564 1052 590 1054
rect 564 1051 565 1052
rect 559 1050 565 1051
rect 542 1045 548 1046
rect 542 1041 543 1045
rect 547 1041 548 1045
rect 542 1040 548 1041
rect 559 1039 565 1040
rect 559 1038 560 1039
rect 532 1036 560 1038
rect 503 1034 509 1035
rect 559 1035 560 1036
rect 564 1035 565 1039
rect 588 1038 590 1052
rect 615 1051 616 1055
rect 620 1054 621 1055
rect 679 1055 685 1056
rect 620 1052 650 1054
rect 620 1051 621 1052
rect 615 1050 621 1051
rect 598 1045 604 1046
rect 598 1041 599 1045
rect 603 1041 604 1045
rect 598 1040 604 1041
rect 615 1039 621 1040
rect 615 1038 616 1039
rect 588 1036 616 1038
rect 559 1034 565 1035
rect 615 1035 616 1036
rect 620 1035 621 1039
rect 648 1038 650 1052
rect 679 1051 680 1055
rect 684 1054 685 1055
rect 743 1055 749 1056
rect 684 1052 738 1054
rect 684 1051 685 1052
rect 679 1050 685 1051
rect 662 1045 668 1046
rect 662 1041 663 1045
rect 667 1041 668 1045
rect 662 1040 668 1041
rect 726 1045 732 1046
rect 726 1041 727 1045
rect 731 1041 732 1045
rect 726 1040 732 1041
rect 679 1039 685 1040
rect 679 1038 680 1039
rect 648 1036 680 1038
rect 615 1034 621 1035
rect 679 1035 680 1036
rect 684 1035 685 1039
rect 736 1038 738 1052
rect 743 1051 744 1055
rect 748 1051 749 1055
rect 743 1050 749 1051
rect 807 1055 813 1056
rect 807 1051 808 1055
rect 812 1054 813 1055
rect 879 1055 885 1056
rect 812 1052 874 1054
rect 812 1051 813 1052
rect 807 1050 813 1051
rect 790 1045 796 1046
rect 790 1041 791 1045
rect 795 1041 796 1045
rect 790 1040 796 1041
rect 862 1045 868 1046
rect 862 1041 863 1045
rect 867 1041 868 1045
rect 862 1040 868 1041
rect 743 1039 749 1040
rect 743 1038 744 1039
rect 736 1036 744 1038
rect 679 1034 685 1035
rect 743 1035 744 1036
rect 748 1035 749 1039
rect 743 1034 749 1035
rect 807 1039 813 1040
rect 807 1035 808 1039
rect 812 1035 813 1039
rect 872 1038 874 1052
rect 879 1051 880 1055
rect 884 1054 885 1055
rect 951 1055 957 1056
rect 884 1052 918 1054
rect 884 1051 885 1052
rect 879 1050 885 1051
rect 879 1039 885 1040
rect 879 1038 880 1039
rect 872 1036 880 1038
rect 807 1034 813 1035
rect 879 1035 880 1036
rect 884 1035 885 1039
rect 916 1038 918 1052
rect 951 1051 952 1055
rect 956 1054 957 1055
rect 986 1055 992 1056
rect 986 1054 987 1055
rect 956 1052 987 1054
rect 956 1051 957 1052
rect 951 1050 957 1051
rect 986 1051 987 1052
rect 991 1051 992 1055
rect 986 1050 992 1051
rect 994 1055 1000 1056
rect 994 1051 995 1055
rect 999 1054 1000 1055
rect 1023 1055 1029 1056
rect 1023 1054 1024 1055
rect 999 1052 1024 1054
rect 999 1051 1000 1052
rect 994 1050 1000 1051
rect 1023 1051 1024 1052
rect 1028 1051 1029 1055
rect 1095 1055 1101 1056
rect 1095 1054 1096 1055
rect 1023 1050 1029 1051
rect 1064 1052 1096 1054
rect 934 1045 940 1046
rect 934 1041 935 1045
rect 939 1041 940 1045
rect 934 1040 940 1041
rect 1006 1045 1012 1046
rect 1006 1041 1007 1045
rect 1011 1041 1012 1045
rect 1006 1040 1012 1041
rect 951 1039 957 1040
rect 951 1038 952 1039
rect 916 1036 952 1038
rect 879 1034 885 1035
rect 951 1035 952 1036
rect 956 1035 957 1039
rect 1023 1039 1029 1040
rect 951 1034 957 1035
rect 994 1035 1000 1036
rect 994 1034 995 1035
rect 718 1031 724 1032
rect 718 1030 719 1031
rect 593 1028 719 1030
rect 593 1024 595 1028
rect 718 1027 719 1028
rect 723 1027 724 1031
rect 809 1030 811 1034
rect 960 1032 995 1034
rect 960 1030 962 1032
rect 994 1031 995 1032
rect 999 1031 1000 1035
rect 1023 1035 1024 1039
rect 1028 1038 1029 1039
rect 1064 1038 1066 1052
rect 1095 1051 1096 1052
rect 1100 1051 1101 1055
rect 1167 1055 1173 1056
rect 1167 1054 1168 1055
rect 1095 1050 1101 1051
rect 1132 1052 1168 1054
rect 1078 1045 1084 1046
rect 1078 1041 1079 1045
rect 1083 1041 1084 1045
rect 1078 1040 1084 1041
rect 1028 1036 1066 1038
rect 1095 1039 1101 1040
rect 1028 1035 1029 1036
rect 1023 1034 1029 1035
rect 1095 1035 1096 1039
rect 1100 1038 1101 1039
rect 1132 1038 1134 1052
rect 1167 1051 1168 1052
rect 1172 1051 1173 1055
rect 1167 1050 1173 1051
rect 1186 1055 1192 1056
rect 1186 1051 1187 1055
rect 1191 1054 1192 1055
rect 1231 1055 1237 1056
rect 1231 1054 1232 1055
rect 1191 1052 1232 1054
rect 1191 1051 1192 1052
rect 1186 1050 1192 1051
rect 1231 1051 1232 1052
rect 1236 1051 1237 1055
rect 1295 1055 1301 1056
rect 1295 1054 1296 1055
rect 1231 1050 1237 1051
rect 1265 1052 1296 1054
rect 1150 1045 1156 1046
rect 1150 1041 1151 1045
rect 1155 1041 1156 1045
rect 1150 1040 1156 1041
rect 1214 1045 1220 1046
rect 1214 1041 1215 1045
rect 1219 1041 1220 1045
rect 1214 1040 1220 1041
rect 1100 1036 1134 1038
rect 1166 1039 1173 1040
rect 1100 1035 1101 1036
rect 1095 1034 1101 1035
rect 1166 1035 1167 1039
rect 1172 1035 1173 1039
rect 1166 1034 1173 1035
rect 1231 1039 1237 1040
rect 1231 1035 1232 1039
rect 1236 1038 1237 1039
rect 1265 1038 1267 1052
rect 1295 1051 1296 1052
rect 1300 1051 1301 1055
rect 1351 1055 1357 1056
rect 1351 1054 1352 1055
rect 1295 1050 1301 1051
rect 1324 1052 1352 1054
rect 1278 1045 1284 1046
rect 1278 1041 1279 1045
rect 1283 1041 1284 1045
rect 1278 1040 1284 1041
rect 1236 1036 1267 1038
rect 1295 1039 1301 1040
rect 1236 1035 1237 1036
rect 1231 1034 1237 1035
rect 1295 1035 1296 1039
rect 1300 1038 1301 1039
rect 1324 1038 1326 1052
rect 1351 1051 1352 1052
rect 1356 1051 1357 1055
rect 1351 1050 1357 1051
rect 1407 1055 1416 1056
rect 1407 1051 1408 1055
rect 1415 1051 1416 1055
rect 1463 1055 1469 1056
rect 1463 1054 1464 1055
rect 1407 1050 1416 1051
rect 1459 1052 1464 1054
rect 1334 1045 1340 1046
rect 1334 1041 1335 1045
rect 1339 1041 1340 1045
rect 1334 1040 1340 1041
rect 1390 1045 1396 1046
rect 1390 1041 1391 1045
rect 1395 1041 1396 1045
rect 1390 1040 1396 1041
rect 1446 1045 1452 1046
rect 1446 1041 1447 1045
rect 1451 1041 1452 1045
rect 1446 1040 1452 1041
rect 1300 1036 1326 1038
rect 1351 1039 1357 1040
rect 1300 1035 1301 1036
rect 1295 1034 1301 1035
rect 1351 1035 1352 1039
rect 1356 1038 1357 1039
rect 1382 1039 1388 1040
rect 1382 1038 1383 1039
rect 1356 1036 1383 1038
rect 1356 1035 1357 1036
rect 1351 1034 1357 1035
rect 1382 1035 1383 1036
rect 1387 1035 1388 1039
rect 1382 1034 1388 1035
rect 1407 1039 1413 1040
rect 1407 1035 1408 1039
rect 1412 1038 1413 1039
rect 1459 1038 1461 1052
rect 1463 1051 1464 1052
rect 1468 1051 1469 1055
rect 1519 1055 1525 1056
rect 1519 1054 1520 1055
rect 1463 1050 1469 1051
rect 1488 1052 1520 1054
rect 1488 1046 1490 1052
rect 1519 1051 1520 1052
rect 1524 1051 1525 1055
rect 1519 1050 1525 1051
rect 1530 1055 1536 1056
rect 1530 1051 1531 1055
rect 1535 1054 1536 1055
rect 1559 1055 1565 1056
rect 1559 1054 1560 1055
rect 1535 1052 1560 1054
rect 1535 1051 1536 1052
rect 1530 1050 1536 1051
rect 1559 1051 1560 1052
rect 1564 1051 1565 1055
rect 1559 1050 1565 1051
rect 1468 1044 1490 1046
rect 1502 1045 1508 1046
rect 1468 1040 1470 1044
rect 1502 1041 1503 1045
rect 1507 1041 1508 1045
rect 1502 1040 1508 1041
rect 1542 1045 1548 1046
rect 1542 1041 1543 1045
rect 1547 1041 1548 1045
rect 1542 1040 1548 1041
rect 1582 1044 1588 1045
rect 1582 1040 1583 1044
rect 1587 1040 1588 1044
rect 1412 1036 1461 1038
rect 1463 1039 1470 1040
rect 1412 1035 1413 1036
rect 1407 1034 1413 1035
rect 1463 1035 1464 1039
rect 1468 1036 1470 1039
rect 1474 1039 1480 1040
rect 1468 1035 1469 1036
rect 1463 1034 1469 1035
rect 1474 1035 1475 1039
rect 1479 1038 1480 1039
rect 1519 1039 1525 1040
rect 1519 1038 1520 1039
rect 1479 1036 1520 1038
rect 1479 1035 1480 1036
rect 1474 1034 1480 1035
rect 1519 1035 1520 1036
rect 1524 1035 1525 1039
rect 1519 1034 1525 1035
rect 1558 1039 1565 1040
rect 1582 1039 1588 1040
rect 1558 1035 1559 1039
rect 1564 1035 1565 1039
rect 1558 1034 1565 1035
rect 994 1030 1000 1031
rect 809 1028 962 1030
rect 718 1026 724 1027
rect 986 1027 992 1028
rect 527 1023 533 1024
rect 110 1020 116 1021
rect 110 1016 111 1020
rect 115 1016 116 1020
rect 110 1015 116 1016
rect 510 1019 516 1020
rect 510 1015 511 1019
rect 515 1015 516 1019
rect 527 1019 528 1023
rect 532 1022 533 1023
rect 559 1023 565 1024
rect 532 1020 539 1022
rect 532 1019 533 1020
rect 527 1018 533 1019
rect 510 1014 516 1015
rect 471 1011 477 1012
rect 471 1007 472 1011
rect 476 1010 477 1011
rect 537 1010 539 1020
rect 542 1019 548 1020
rect 542 1015 543 1019
rect 547 1015 548 1019
rect 559 1019 560 1023
rect 564 1022 565 1023
rect 591 1023 597 1024
rect 564 1020 570 1022
rect 564 1019 565 1020
rect 559 1018 565 1019
rect 542 1014 548 1015
rect 568 1010 570 1020
rect 574 1019 580 1020
rect 574 1015 575 1019
rect 579 1015 580 1019
rect 591 1019 592 1023
rect 596 1019 597 1023
rect 626 1023 637 1024
rect 591 1018 597 1019
rect 614 1019 620 1020
rect 574 1014 580 1015
rect 614 1015 615 1019
rect 619 1015 620 1019
rect 626 1019 627 1023
rect 631 1019 632 1023
rect 636 1019 637 1023
rect 679 1023 685 1024
rect 679 1022 680 1023
rect 672 1020 680 1022
rect 626 1018 637 1019
rect 662 1019 668 1020
rect 614 1014 620 1015
rect 662 1015 663 1019
rect 667 1015 668 1019
rect 662 1014 668 1015
rect 672 1010 674 1020
rect 679 1019 680 1020
rect 684 1019 685 1023
rect 727 1023 733 1024
rect 727 1022 728 1023
rect 720 1020 728 1022
rect 679 1018 685 1019
rect 710 1019 716 1020
rect 710 1015 711 1019
rect 715 1015 716 1019
rect 710 1014 716 1015
rect 720 1010 722 1020
rect 727 1019 728 1020
rect 732 1019 733 1023
rect 791 1023 797 1024
rect 727 1018 733 1019
rect 774 1019 780 1020
rect 774 1015 775 1019
rect 779 1015 780 1019
rect 791 1019 792 1023
rect 796 1022 797 1023
rect 863 1023 869 1024
rect 796 1020 830 1022
rect 796 1019 797 1020
rect 791 1018 797 1019
rect 774 1014 780 1015
rect 476 1008 522 1010
rect 537 1008 554 1010
rect 568 1008 586 1010
rect 656 1008 674 1010
rect 681 1008 722 1010
rect 828 1010 830 1020
rect 846 1019 852 1020
rect 846 1015 847 1019
rect 851 1015 852 1019
rect 863 1019 864 1023
rect 868 1022 869 1023
rect 943 1023 949 1024
rect 868 1020 906 1022
rect 868 1019 869 1020
rect 863 1018 869 1019
rect 846 1014 852 1015
rect 904 1010 906 1020
rect 926 1019 932 1020
rect 926 1015 927 1019
rect 931 1015 932 1019
rect 943 1019 944 1023
rect 948 1022 949 1023
rect 978 1023 984 1024
rect 978 1022 979 1023
rect 948 1020 979 1022
rect 948 1019 949 1020
rect 943 1018 949 1019
rect 978 1019 979 1020
rect 983 1019 984 1023
rect 986 1023 987 1027
rect 991 1026 992 1027
rect 991 1024 1018 1026
rect 991 1023 992 1024
rect 986 1022 992 1023
rect 1016 1022 1018 1024
rect 1023 1023 1029 1024
rect 1023 1022 1024 1023
rect 1016 1020 1024 1022
rect 978 1018 984 1019
rect 1006 1019 1012 1020
rect 926 1014 932 1015
rect 1006 1015 1007 1019
rect 1011 1015 1012 1019
rect 1023 1019 1024 1020
rect 1028 1019 1029 1023
rect 1103 1023 1109 1024
rect 1103 1022 1104 1023
rect 1099 1020 1104 1022
rect 1023 1018 1029 1019
rect 1086 1019 1092 1020
rect 1006 1014 1012 1015
rect 1086 1015 1087 1019
rect 1091 1015 1092 1019
rect 1086 1014 1092 1015
rect 1099 1010 1101 1020
rect 1103 1019 1104 1020
rect 1108 1019 1109 1023
rect 1183 1023 1192 1024
rect 1103 1018 1109 1019
rect 1166 1019 1172 1020
rect 1166 1015 1167 1019
rect 1171 1015 1172 1019
rect 1183 1019 1184 1023
rect 1191 1019 1192 1023
rect 1255 1023 1261 1024
rect 1255 1022 1256 1023
rect 1248 1020 1256 1022
rect 1183 1018 1192 1019
rect 1238 1019 1244 1020
rect 1166 1014 1172 1015
rect 1238 1015 1239 1019
rect 1243 1015 1244 1019
rect 1238 1014 1244 1015
rect 1248 1010 1250 1020
rect 1255 1019 1256 1020
rect 1260 1019 1261 1023
rect 1319 1023 1325 1024
rect 1319 1022 1320 1023
rect 1312 1020 1320 1022
rect 1255 1018 1261 1019
rect 1302 1019 1308 1020
rect 1302 1015 1303 1019
rect 1307 1015 1308 1019
rect 1302 1014 1308 1015
rect 1312 1010 1314 1020
rect 1319 1019 1320 1020
rect 1324 1019 1325 1023
rect 1375 1023 1381 1024
rect 1375 1022 1376 1023
rect 1368 1020 1376 1022
rect 1319 1018 1325 1019
rect 1358 1019 1364 1020
rect 1358 1015 1359 1019
rect 1363 1015 1364 1019
rect 1358 1014 1364 1015
rect 1368 1010 1370 1020
rect 1375 1019 1376 1020
rect 1380 1019 1381 1023
rect 1423 1023 1429 1024
rect 1423 1022 1424 1023
rect 1416 1020 1424 1022
rect 1375 1018 1381 1019
rect 1406 1019 1412 1020
rect 1406 1015 1407 1019
rect 1411 1015 1412 1019
rect 1406 1014 1412 1015
rect 1416 1010 1418 1020
rect 1423 1019 1424 1020
rect 1428 1019 1429 1023
rect 1471 1023 1477 1024
rect 1471 1022 1472 1023
rect 1464 1020 1472 1022
rect 1423 1018 1429 1019
rect 1454 1019 1460 1020
rect 1454 1015 1455 1019
rect 1459 1015 1460 1019
rect 1454 1014 1460 1015
rect 1464 1010 1466 1020
rect 1471 1019 1472 1020
rect 1476 1019 1477 1023
rect 1527 1023 1536 1024
rect 1471 1018 1477 1019
rect 1510 1019 1516 1020
rect 1510 1015 1511 1019
rect 1515 1015 1516 1019
rect 1527 1019 1528 1023
rect 1535 1019 1536 1023
rect 1559 1023 1565 1024
rect 1559 1022 1560 1023
rect 1552 1020 1560 1022
rect 1527 1018 1536 1019
rect 1542 1019 1548 1020
rect 1510 1014 1516 1015
rect 1542 1015 1543 1019
rect 1547 1015 1548 1019
rect 1542 1014 1548 1015
rect 1552 1010 1554 1020
rect 1559 1019 1560 1020
rect 1564 1019 1565 1023
rect 1559 1018 1565 1019
rect 1582 1020 1588 1021
rect 1582 1016 1583 1020
rect 1587 1016 1588 1020
rect 1582 1015 1588 1016
rect 828 1008 858 1010
rect 904 1008 938 1010
rect 1060 1008 1101 1010
rect 1185 1008 1250 1010
rect 1288 1008 1314 1010
rect 1321 1008 1370 1010
rect 1377 1008 1418 1010
rect 1441 1008 1466 1010
rect 1540 1008 1554 1010
rect 476 1007 477 1008
rect 471 1006 477 1007
rect 520 1006 522 1008
rect 527 1007 533 1008
rect 527 1006 528 1007
rect 520 1004 528 1006
rect 110 1003 116 1004
rect 110 999 111 1003
rect 115 999 116 1003
rect 527 1003 528 1004
rect 532 1003 533 1007
rect 552 1006 554 1008
rect 559 1007 565 1008
rect 559 1006 560 1007
rect 552 1004 560 1006
rect 527 1002 533 1003
rect 559 1003 560 1004
rect 564 1003 565 1007
rect 584 1006 586 1008
rect 591 1007 597 1008
rect 591 1006 592 1007
rect 584 1004 592 1006
rect 559 1002 565 1003
rect 591 1003 592 1004
rect 596 1003 597 1007
rect 591 1002 597 1003
rect 631 1007 637 1008
rect 631 1003 632 1007
rect 636 1006 637 1007
rect 656 1006 658 1008
rect 636 1004 658 1006
rect 679 1007 685 1008
rect 636 1003 637 1004
rect 631 1002 637 1003
rect 679 1003 680 1007
rect 684 1003 685 1007
rect 679 1002 685 1003
rect 726 1007 733 1008
rect 726 1003 727 1007
rect 732 1003 733 1007
rect 726 1002 733 1003
rect 790 1007 797 1008
rect 790 1003 791 1007
rect 796 1003 797 1007
rect 856 1006 858 1008
rect 863 1007 869 1008
rect 863 1006 864 1007
rect 856 1004 864 1006
rect 790 1002 797 1003
rect 863 1003 864 1004
rect 868 1003 869 1007
rect 936 1006 938 1008
rect 943 1007 949 1008
rect 943 1006 944 1007
rect 936 1004 944 1006
rect 863 1002 869 1003
rect 943 1003 944 1004
rect 948 1003 949 1007
rect 943 1002 949 1003
rect 1023 1007 1029 1008
rect 1023 1003 1024 1007
rect 1028 1006 1029 1007
rect 1060 1006 1062 1008
rect 1103 1007 1109 1008
rect 1103 1006 1104 1007
rect 1028 1004 1062 1006
rect 1099 1004 1104 1006
rect 1028 1003 1029 1004
rect 1023 1002 1029 1003
rect 110 998 116 999
rect 510 1001 516 1002
rect 510 997 511 1001
rect 515 997 516 1001
rect 510 996 516 997
rect 542 1001 548 1002
rect 542 997 543 1001
rect 547 997 548 1001
rect 542 996 548 997
rect 574 1001 580 1002
rect 574 997 575 1001
rect 579 997 580 1001
rect 574 996 580 997
rect 614 1001 620 1002
rect 614 997 615 1001
rect 619 997 620 1001
rect 614 996 620 997
rect 662 1001 668 1002
rect 662 997 663 1001
rect 667 997 668 1001
rect 662 996 668 997
rect 710 1001 716 1002
rect 710 997 711 1001
rect 715 997 716 1001
rect 710 996 716 997
rect 774 1001 780 1002
rect 774 997 775 1001
rect 779 997 780 1001
rect 774 996 780 997
rect 846 1001 852 1002
rect 846 997 847 1001
rect 851 997 852 1001
rect 846 996 852 997
rect 926 1001 932 1002
rect 926 997 927 1001
rect 931 997 932 1001
rect 926 996 932 997
rect 1006 1001 1012 1002
rect 1006 997 1007 1001
rect 1011 997 1012 1001
rect 1006 996 1012 997
rect 1086 1001 1092 1002
rect 1086 997 1087 1001
rect 1091 997 1092 1001
rect 1086 996 1092 997
rect 978 995 984 996
rect 978 991 979 995
rect 983 994 984 995
rect 1099 994 1101 1004
rect 1103 1003 1104 1004
rect 1108 1003 1109 1007
rect 1103 1002 1109 1003
rect 1183 1007 1189 1008
rect 1183 1003 1184 1007
rect 1188 1003 1189 1007
rect 1183 1002 1189 1003
rect 1255 1007 1261 1008
rect 1255 1003 1256 1007
rect 1260 1006 1261 1007
rect 1288 1006 1290 1008
rect 1260 1004 1290 1006
rect 1319 1007 1325 1008
rect 1260 1003 1261 1004
rect 1255 1002 1261 1003
rect 1319 1003 1320 1007
rect 1324 1003 1325 1007
rect 1319 1002 1325 1003
rect 1375 1007 1381 1008
rect 1375 1003 1376 1007
rect 1380 1003 1381 1007
rect 1375 1002 1381 1003
rect 1423 1007 1429 1008
rect 1423 1003 1424 1007
rect 1428 1006 1429 1007
rect 1441 1006 1443 1008
rect 1428 1004 1443 1006
rect 1471 1007 1480 1008
rect 1428 1003 1429 1004
rect 1423 1002 1429 1003
rect 1471 1003 1472 1007
rect 1479 1003 1480 1007
rect 1471 1002 1480 1003
rect 1527 1007 1533 1008
rect 1527 1003 1528 1007
rect 1532 1006 1533 1007
rect 1540 1006 1542 1008
rect 1532 1004 1542 1006
rect 1558 1007 1565 1008
rect 1532 1003 1533 1004
rect 1527 1002 1533 1003
rect 1558 1003 1559 1007
rect 1564 1003 1565 1007
rect 1558 1002 1565 1003
rect 1582 1003 1588 1004
rect 1166 1001 1172 1002
rect 1166 997 1167 1001
rect 1171 997 1172 1001
rect 1166 996 1172 997
rect 1238 1001 1244 1002
rect 1238 997 1239 1001
rect 1243 997 1244 1001
rect 1238 996 1244 997
rect 1302 1001 1308 1002
rect 1302 997 1303 1001
rect 1307 997 1308 1001
rect 1302 996 1308 997
rect 1358 1001 1364 1002
rect 1358 997 1359 1001
rect 1363 997 1364 1001
rect 1358 996 1364 997
rect 1406 1001 1412 1002
rect 1406 997 1407 1001
rect 1411 997 1412 1001
rect 1406 996 1412 997
rect 1454 1001 1460 1002
rect 1454 997 1455 1001
rect 1459 997 1460 1001
rect 1454 996 1460 997
rect 1510 1001 1516 1002
rect 1510 997 1511 1001
rect 1515 997 1516 1001
rect 1510 996 1516 997
rect 1542 1001 1548 1002
rect 1542 997 1543 1001
rect 1547 997 1548 1001
rect 1582 999 1583 1003
rect 1587 999 1588 1003
rect 1582 998 1588 999
rect 1542 996 1548 997
rect 983 992 1101 994
rect 983 991 984 992
rect 978 990 984 991
rect 626 987 632 988
rect 626 986 627 987
rect 577 984 627 986
rect 158 979 164 980
rect 110 977 116 978
rect 110 973 111 977
rect 115 973 116 977
rect 158 975 159 979
rect 163 975 164 979
rect 158 974 164 975
rect 198 979 204 980
rect 198 975 199 979
rect 203 975 204 979
rect 198 974 204 975
rect 254 979 260 980
rect 254 975 255 979
rect 259 975 260 979
rect 254 974 260 975
rect 310 979 316 980
rect 310 975 311 979
rect 315 975 316 979
rect 310 974 316 975
rect 374 979 380 980
rect 374 975 375 979
rect 379 975 380 979
rect 374 974 380 975
rect 438 979 444 980
rect 438 975 439 979
rect 443 975 444 979
rect 438 974 444 975
rect 502 979 508 980
rect 502 975 503 979
rect 507 975 508 979
rect 502 974 508 975
rect 558 979 564 980
rect 558 975 559 979
rect 563 975 564 979
rect 558 974 564 975
rect 110 972 116 973
rect 577 972 579 984
rect 626 983 627 984
rect 631 983 632 987
rect 626 982 632 983
rect 822 987 828 988
rect 822 983 823 987
rect 827 986 828 987
rect 827 984 1147 986
rect 827 983 828 984
rect 822 982 828 983
rect 614 979 620 980
rect 614 975 615 979
rect 619 975 620 979
rect 614 974 620 975
rect 662 979 668 980
rect 662 975 663 979
rect 667 975 668 979
rect 662 974 668 975
rect 702 979 708 980
rect 702 975 703 979
rect 707 975 708 979
rect 702 974 708 975
rect 734 979 740 980
rect 734 975 735 979
rect 739 975 740 979
rect 734 974 740 975
rect 774 979 780 980
rect 774 975 775 979
rect 779 975 780 979
rect 774 974 780 975
rect 830 979 836 980
rect 830 975 831 979
rect 835 975 836 979
rect 830 974 836 975
rect 894 979 900 980
rect 894 975 895 979
rect 899 975 900 979
rect 894 974 900 975
rect 966 979 972 980
rect 966 975 967 979
rect 971 975 972 979
rect 966 974 972 975
rect 1046 979 1052 980
rect 1046 975 1047 979
rect 1051 975 1052 979
rect 1046 974 1052 975
rect 1126 979 1132 980
rect 1126 975 1127 979
rect 1131 975 1132 979
rect 1126 974 1132 975
rect 1145 972 1147 984
rect 1198 979 1204 980
rect 1198 975 1199 979
rect 1203 975 1204 979
rect 1198 974 1204 975
rect 1270 979 1276 980
rect 1270 975 1271 979
rect 1275 975 1276 979
rect 1270 974 1276 975
rect 1342 979 1348 980
rect 1342 975 1343 979
rect 1347 975 1348 979
rect 1342 974 1348 975
rect 1414 979 1420 980
rect 1414 975 1415 979
rect 1419 975 1420 979
rect 1414 974 1420 975
rect 1486 979 1492 980
rect 1486 975 1487 979
rect 1491 975 1492 979
rect 1486 974 1492 975
rect 1542 979 1548 980
rect 1542 975 1543 979
rect 1547 975 1548 979
rect 1542 974 1548 975
rect 1582 977 1588 978
rect 1582 973 1583 977
rect 1587 973 1588 977
rect 1582 972 1588 973
rect 170 971 181 972
rect 170 967 171 971
rect 175 967 176 971
rect 180 967 181 971
rect 215 971 221 972
rect 215 970 216 971
rect 170 966 181 967
rect 193 968 216 970
rect 158 961 164 962
rect 110 960 116 961
rect 110 956 111 960
rect 115 956 116 960
rect 158 957 159 961
rect 163 957 164 961
rect 158 956 164 957
rect 110 955 116 956
rect 175 955 181 956
rect 175 951 176 955
rect 180 954 181 955
rect 193 954 195 968
rect 215 967 216 968
rect 220 967 221 971
rect 271 971 277 972
rect 271 970 272 971
rect 215 966 221 967
rect 240 968 272 970
rect 198 961 204 962
rect 198 957 199 961
rect 203 957 204 961
rect 198 956 204 957
rect 180 952 195 954
rect 215 955 221 956
rect 180 951 181 952
rect 175 950 181 951
rect 215 951 216 955
rect 220 954 221 955
rect 240 954 242 968
rect 271 967 272 968
rect 276 967 277 971
rect 327 971 333 972
rect 327 970 328 971
rect 271 966 277 967
rect 300 968 328 970
rect 254 961 260 962
rect 254 957 255 961
rect 259 957 260 961
rect 254 956 260 957
rect 220 952 242 954
rect 271 955 277 956
rect 220 951 221 952
rect 215 950 221 951
rect 271 951 272 955
rect 276 954 277 955
rect 300 954 302 968
rect 327 967 328 968
rect 332 967 333 971
rect 391 971 397 972
rect 391 970 392 971
rect 327 966 333 967
rect 364 968 392 970
rect 310 961 316 962
rect 310 957 311 961
rect 315 957 316 961
rect 310 956 316 957
rect 276 952 302 954
rect 327 955 333 956
rect 276 951 277 952
rect 271 950 277 951
rect 327 951 328 955
rect 332 954 333 955
rect 364 954 366 968
rect 391 967 392 968
rect 396 967 397 971
rect 455 971 461 972
rect 455 970 456 971
rect 391 966 397 967
rect 425 968 456 970
rect 374 961 380 962
rect 374 957 375 961
rect 379 957 380 961
rect 374 956 380 957
rect 332 952 366 954
rect 391 955 397 956
rect 332 951 333 952
rect 327 950 333 951
rect 391 951 392 955
rect 396 954 397 955
rect 425 954 427 968
rect 455 967 456 968
rect 460 967 461 971
rect 455 966 461 967
rect 519 971 525 972
rect 519 967 520 971
rect 524 970 525 971
rect 575 971 581 972
rect 524 968 570 970
rect 524 967 525 968
rect 519 966 525 967
rect 438 961 444 962
rect 438 957 439 961
rect 443 957 444 961
rect 438 956 444 957
rect 502 961 508 962
rect 502 957 503 961
rect 507 957 508 961
rect 502 956 508 957
rect 558 961 564 962
rect 558 957 559 961
rect 563 957 564 961
rect 558 956 564 957
rect 568 958 570 968
rect 575 967 576 971
rect 580 967 581 971
rect 575 966 581 967
rect 586 971 592 972
rect 586 967 587 971
rect 591 970 592 971
rect 631 971 637 972
rect 631 970 632 971
rect 591 968 632 970
rect 591 967 592 968
rect 586 966 592 967
rect 631 967 632 968
rect 636 967 637 971
rect 679 971 685 972
rect 679 970 680 971
rect 631 966 637 967
rect 656 968 680 970
rect 614 961 620 962
rect 568 956 579 958
rect 614 957 615 961
rect 619 957 620 961
rect 614 956 620 957
rect 396 952 427 954
rect 450 955 461 956
rect 396 951 397 952
rect 391 950 397 951
rect 450 951 451 955
rect 455 951 456 955
rect 460 951 461 955
rect 450 950 461 951
rect 519 955 528 956
rect 519 951 520 955
rect 527 951 528 955
rect 519 950 528 951
rect 575 955 581 956
rect 575 951 576 955
rect 580 951 581 955
rect 575 950 581 951
rect 631 955 637 956
rect 631 951 632 955
rect 636 954 637 955
rect 656 954 658 968
rect 679 967 680 968
rect 684 967 685 971
rect 719 971 725 972
rect 719 970 720 971
rect 679 966 685 967
rect 696 968 720 970
rect 662 961 668 962
rect 662 957 663 961
rect 667 957 668 961
rect 662 956 668 957
rect 636 952 658 954
rect 679 955 685 956
rect 636 951 637 952
rect 631 950 637 951
rect 679 951 680 955
rect 684 954 685 955
rect 696 954 698 968
rect 719 967 720 968
rect 724 967 725 971
rect 751 971 757 972
rect 751 970 752 971
rect 719 966 725 967
rect 744 968 752 970
rect 702 961 708 962
rect 702 957 703 961
rect 707 957 708 961
rect 702 956 708 957
rect 734 961 740 962
rect 734 957 735 961
rect 739 957 740 961
rect 734 956 740 957
rect 684 952 698 954
rect 719 955 725 956
rect 684 951 685 952
rect 679 950 685 951
rect 719 951 720 955
rect 724 954 725 955
rect 744 954 746 968
rect 751 967 752 968
rect 756 967 757 971
rect 751 966 757 967
rect 791 971 797 972
rect 791 967 792 971
rect 796 970 797 971
rect 847 971 853 972
rect 796 968 822 970
rect 796 967 797 968
rect 791 966 797 967
rect 774 961 780 962
rect 774 957 775 961
rect 779 957 780 961
rect 774 956 780 957
rect 724 952 746 954
rect 751 955 757 956
rect 724 951 725 952
rect 719 950 725 951
rect 751 951 752 955
rect 756 954 757 955
rect 782 955 788 956
rect 782 954 783 955
rect 756 952 783 954
rect 756 951 757 952
rect 751 950 757 951
rect 782 951 783 952
rect 787 951 788 955
rect 782 950 788 951
rect 790 955 797 956
rect 790 951 791 955
rect 796 951 797 955
rect 820 954 822 968
rect 847 967 848 971
rect 852 970 853 971
rect 911 971 917 972
rect 852 968 882 970
rect 852 967 853 968
rect 847 966 853 967
rect 830 961 836 962
rect 830 957 831 961
rect 835 957 836 961
rect 830 956 836 957
rect 847 955 853 956
rect 847 954 848 955
rect 820 952 848 954
rect 790 950 797 951
rect 847 951 848 952
rect 852 951 853 955
rect 880 954 882 968
rect 911 967 912 971
rect 916 970 917 971
rect 983 971 989 972
rect 916 968 950 970
rect 916 967 917 968
rect 911 966 917 967
rect 894 961 900 962
rect 894 957 895 961
rect 899 957 900 961
rect 894 956 900 957
rect 911 955 917 956
rect 911 954 912 955
rect 880 952 912 954
rect 847 950 853 951
rect 911 951 912 952
rect 916 951 917 955
rect 948 954 950 968
rect 983 967 984 971
rect 988 970 989 971
rect 1063 971 1069 972
rect 988 968 1026 970
rect 988 967 989 968
rect 983 966 989 967
rect 966 961 972 962
rect 966 957 967 961
rect 971 957 972 961
rect 966 956 972 957
rect 983 955 989 956
rect 983 954 984 955
rect 948 952 984 954
rect 911 950 917 951
rect 983 951 984 952
rect 988 951 989 955
rect 1024 954 1026 968
rect 1063 967 1064 971
rect 1068 970 1069 971
rect 1143 971 1149 972
rect 1068 968 1138 970
rect 1068 967 1069 968
rect 1063 966 1069 967
rect 1046 961 1052 962
rect 1046 957 1047 961
rect 1051 957 1052 961
rect 1046 956 1052 957
rect 1126 961 1132 962
rect 1126 957 1127 961
rect 1131 957 1132 961
rect 1126 956 1132 957
rect 1063 955 1069 956
rect 1063 954 1064 955
rect 1024 952 1064 954
rect 983 950 989 951
rect 1063 951 1064 952
rect 1068 951 1069 955
rect 1136 954 1138 968
rect 1143 967 1144 971
rect 1148 967 1149 971
rect 1143 966 1149 967
rect 1215 971 1224 972
rect 1215 967 1216 971
rect 1223 967 1224 971
rect 1287 971 1293 972
rect 1287 970 1288 971
rect 1215 966 1224 967
rect 1252 968 1288 970
rect 1198 961 1204 962
rect 1198 957 1199 961
rect 1203 957 1204 961
rect 1198 956 1204 957
rect 1143 955 1149 956
rect 1143 954 1144 955
rect 1136 952 1144 954
rect 1063 950 1069 951
rect 1143 951 1144 952
rect 1148 951 1149 955
rect 1143 950 1149 951
rect 1215 955 1221 956
rect 1215 951 1216 955
rect 1220 954 1221 955
rect 1252 954 1254 968
rect 1287 967 1288 968
rect 1292 967 1293 971
rect 1359 971 1365 972
rect 1359 970 1360 971
rect 1287 966 1293 967
rect 1324 968 1360 970
rect 1270 961 1276 962
rect 1270 957 1271 961
rect 1275 957 1276 961
rect 1270 956 1276 957
rect 1220 952 1254 954
rect 1287 955 1293 956
rect 1220 951 1221 952
rect 1215 950 1221 951
rect 1287 951 1288 955
rect 1292 954 1293 955
rect 1324 954 1326 968
rect 1359 967 1360 968
rect 1364 967 1365 971
rect 1431 971 1437 972
rect 1431 970 1432 971
rect 1359 966 1365 967
rect 1396 968 1432 970
rect 1342 961 1348 962
rect 1342 957 1343 961
rect 1347 957 1348 961
rect 1342 956 1348 957
rect 1292 952 1326 954
rect 1359 955 1365 956
rect 1292 951 1293 952
rect 1287 950 1293 951
rect 1359 951 1360 955
rect 1364 954 1365 955
rect 1396 954 1398 968
rect 1431 967 1432 968
rect 1436 967 1437 971
rect 1503 971 1509 972
rect 1503 970 1504 971
rect 1431 966 1437 967
rect 1459 968 1504 970
rect 1414 961 1420 962
rect 1414 957 1415 961
rect 1419 957 1420 961
rect 1414 956 1420 957
rect 1364 952 1398 954
rect 1431 955 1437 956
rect 1364 951 1365 952
rect 1359 950 1365 951
rect 1431 951 1432 955
rect 1436 954 1437 955
rect 1459 954 1461 968
rect 1503 967 1504 968
rect 1508 967 1509 971
rect 1503 966 1509 967
rect 1559 971 1565 972
rect 1559 967 1560 971
rect 1564 970 1565 971
rect 1567 971 1573 972
rect 1567 970 1568 971
rect 1564 968 1568 970
rect 1564 967 1565 968
rect 1559 966 1565 967
rect 1567 967 1568 968
rect 1572 967 1573 971
rect 1567 966 1573 967
rect 1486 961 1492 962
rect 1486 957 1487 961
rect 1491 957 1492 961
rect 1486 956 1492 957
rect 1542 961 1548 962
rect 1542 957 1543 961
rect 1547 957 1548 961
rect 1542 956 1548 957
rect 1582 960 1588 961
rect 1582 956 1583 960
rect 1587 956 1588 960
rect 1436 952 1461 954
rect 1498 955 1509 956
rect 1436 951 1437 952
rect 1431 950 1437 951
rect 1498 951 1499 955
rect 1503 951 1504 955
rect 1508 951 1509 955
rect 1498 950 1509 951
rect 1558 955 1565 956
rect 1582 955 1588 956
rect 1558 951 1559 955
rect 1564 951 1565 955
rect 1558 950 1565 951
rect 822 947 828 948
rect 167 943 176 944
rect 110 940 116 941
rect 110 936 111 940
rect 115 936 116 940
rect 110 935 116 936
rect 150 939 156 940
rect 150 935 151 939
rect 155 935 156 939
rect 167 939 168 943
rect 175 939 176 943
rect 207 943 213 944
rect 207 942 208 943
rect 200 940 208 942
rect 167 938 176 939
rect 190 939 196 940
rect 150 934 156 935
rect 190 935 191 939
rect 195 935 196 939
rect 190 934 196 935
rect 200 930 202 940
rect 207 939 208 940
rect 212 939 213 943
rect 263 943 269 944
rect 263 942 264 943
rect 256 940 264 942
rect 207 938 213 939
rect 246 939 252 940
rect 246 935 247 939
rect 251 935 252 939
rect 246 934 252 935
rect 256 930 258 940
rect 263 939 264 940
rect 268 939 269 943
rect 318 943 325 944
rect 263 938 269 939
rect 302 939 308 940
rect 302 935 303 939
rect 307 935 308 939
rect 318 939 319 943
rect 324 939 325 943
rect 383 943 389 944
rect 383 942 384 943
rect 376 940 384 942
rect 318 938 325 939
rect 366 939 372 940
rect 302 934 308 935
rect 366 935 367 939
rect 371 935 372 939
rect 366 934 372 935
rect 376 930 378 940
rect 383 939 384 940
rect 388 939 389 943
rect 447 943 453 944
rect 447 942 448 943
rect 440 940 448 942
rect 383 938 389 939
rect 430 939 436 940
rect 430 935 431 939
rect 435 935 436 939
rect 430 934 436 935
rect 440 930 442 940
rect 447 939 448 940
rect 452 939 453 943
rect 511 943 517 944
rect 447 938 453 939
rect 494 939 500 940
rect 494 935 495 939
rect 499 935 500 939
rect 511 939 512 943
rect 516 942 517 943
rect 550 943 556 944
rect 550 942 551 943
rect 516 940 551 942
rect 516 939 517 940
rect 511 938 517 939
rect 550 939 551 940
rect 555 939 556 943
rect 575 943 581 944
rect 575 942 576 943
rect 568 940 576 942
rect 550 938 556 939
rect 558 939 564 940
rect 494 934 500 935
rect 558 935 559 939
rect 563 935 564 939
rect 558 934 564 935
rect 568 930 570 940
rect 575 939 576 940
rect 580 939 581 943
rect 631 943 637 944
rect 631 942 632 943
rect 624 940 632 942
rect 575 938 581 939
rect 614 939 620 940
rect 614 935 615 939
rect 619 935 620 939
rect 614 934 620 935
rect 624 930 626 940
rect 631 939 632 940
rect 636 939 637 943
rect 687 943 693 944
rect 687 942 688 943
rect 680 940 688 942
rect 631 938 637 939
rect 670 939 676 940
rect 670 935 671 939
rect 675 935 676 939
rect 670 934 676 935
rect 680 930 682 940
rect 687 939 688 940
rect 692 939 693 943
rect 735 943 741 944
rect 735 942 736 943
rect 728 940 736 942
rect 687 938 693 939
rect 718 939 724 940
rect 718 935 719 939
rect 723 935 724 939
rect 718 934 724 935
rect 728 930 730 940
rect 735 939 736 940
rect 740 939 741 943
rect 783 943 789 944
rect 783 942 784 943
rect 776 940 784 942
rect 735 938 741 939
rect 766 939 772 940
rect 766 935 767 939
rect 771 935 772 939
rect 766 934 772 935
rect 776 930 778 940
rect 783 939 784 940
rect 788 939 789 943
rect 822 943 823 947
rect 827 943 828 947
rect 822 942 828 943
rect 831 943 837 944
rect 831 942 832 943
rect 824 940 832 942
rect 783 938 789 939
rect 814 939 820 940
rect 814 935 815 939
rect 819 935 820 939
rect 831 939 832 940
rect 836 939 837 943
rect 887 943 893 944
rect 887 942 888 943
rect 880 940 888 942
rect 831 938 837 939
rect 870 939 876 940
rect 814 934 820 935
rect 870 935 871 939
rect 875 935 876 939
rect 870 934 876 935
rect 880 930 882 940
rect 887 939 888 940
rect 892 939 893 943
rect 951 943 957 944
rect 951 942 952 943
rect 944 940 952 942
rect 887 938 893 939
rect 934 939 940 940
rect 934 935 935 939
rect 939 935 940 939
rect 934 934 940 935
rect 944 930 946 940
rect 951 939 952 940
rect 956 939 957 943
rect 1023 943 1029 944
rect 1023 942 1024 943
rect 1016 940 1024 942
rect 951 938 957 939
rect 1006 939 1012 940
rect 1006 935 1007 939
rect 1011 935 1012 939
rect 1006 934 1012 935
rect 1016 930 1018 940
rect 1023 939 1024 940
rect 1028 939 1029 943
rect 1095 943 1101 944
rect 1095 942 1096 943
rect 1088 940 1096 942
rect 1023 938 1029 939
rect 1078 939 1084 940
rect 1078 935 1079 939
rect 1083 935 1084 939
rect 1078 934 1084 935
rect 1088 930 1090 940
rect 1095 939 1096 940
rect 1100 939 1101 943
rect 1159 943 1165 944
rect 1159 942 1160 943
rect 1152 940 1160 942
rect 1095 938 1101 939
rect 1142 939 1148 940
rect 1142 935 1143 939
rect 1147 935 1148 939
rect 1142 934 1148 935
rect 1152 930 1154 940
rect 1159 939 1160 940
rect 1164 939 1165 943
rect 1218 943 1229 944
rect 1159 938 1165 939
rect 1206 939 1212 940
rect 1206 935 1207 939
rect 1211 935 1212 939
rect 1218 939 1219 943
rect 1223 939 1224 943
rect 1228 939 1229 943
rect 1287 943 1293 944
rect 1287 942 1288 943
rect 1280 940 1288 942
rect 1218 938 1229 939
rect 1270 939 1276 940
rect 1206 934 1212 935
rect 1270 935 1271 939
rect 1275 935 1276 939
rect 1270 934 1276 935
rect 1280 930 1282 940
rect 1287 939 1288 940
rect 1292 939 1293 943
rect 1343 943 1349 944
rect 1343 942 1344 943
rect 1336 940 1344 942
rect 1287 938 1293 939
rect 1326 939 1332 940
rect 1326 935 1327 939
rect 1331 935 1332 939
rect 1326 934 1332 935
rect 1336 930 1338 940
rect 1343 939 1344 940
rect 1348 939 1349 943
rect 1391 943 1397 944
rect 1343 938 1349 939
rect 1374 939 1380 940
rect 1374 935 1375 939
rect 1379 935 1380 939
rect 1391 939 1392 943
rect 1396 942 1397 943
rect 1399 943 1405 944
rect 1399 942 1400 943
rect 1396 940 1400 942
rect 1396 939 1397 940
rect 1391 938 1397 939
rect 1399 939 1400 940
rect 1404 939 1405 943
rect 1439 943 1445 944
rect 1439 942 1440 943
rect 1432 940 1440 942
rect 1399 938 1405 939
rect 1422 939 1428 940
rect 1374 934 1380 935
rect 1422 935 1423 939
rect 1427 935 1428 939
rect 1422 934 1428 935
rect 1432 930 1434 940
rect 1439 939 1440 940
rect 1444 939 1445 943
rect 1487 943 1493 944
rect 1487 942 1488 943
rect 1480 940 1488 942
rect 1439 938 1445 939
rect 1470 939 1476 940
rect 1470 935 1471 939
rect 1475 935 1476 939
rect 1470 934 1476 935
rect 1480 930 1482 940
rect 1487 939 1488 940
rect 1492 939 1493 943
rect 1527 943 1533 944
rect 1487 938 1493 939
rect 1510 939 1516 940
rect 1510 935 1511 939
rect 1515 935 1516 939
rect 1527 939 1528 943
rect 1532 942 1533 943
rect 1559 943 1565 944
rect 1532 940 1538 942
rect 1532 939 1533 940
rect 1527 938 1533 939
rect 1510 934 1516 935
rect 188 928 202 930
rect 209 928 258 930
rect 321 928 378 930
rect 385 928 442 930
rect 545 928 570 930
rect 577 928 626 930
rect 660 928 682 930
rect 712 928 730 930
rect 737 928 778 930
rect 860 928 882 930
rect 920 928 946 930
rect 988 928 1018 930
rect 1048 928 1090 930
rect 1099 928 1154 930
rect 1256 928 1282 930
rect 1316 928 1338 930
rect 1416 928 1434 930
rect 1441 928 1482 930
rect 1536 930 1538 940
rect 1542 939 1548 940
rect 1542 935 1543 939
rect 1547 935 1548 939
rect 1559 939 1560 943
rect 1564 942 1565 943
rect 1567 943 1573 944
rect 1567 942 1568 943
rect 1564 940 1568 942
rect 1564 939 1565 940
rect 1559 938 1565 939
rect 1567 939 1568 940
rect 1572 939 1573 943
rect 1567 938 1573 939
rect 1582 940 1588 941
rect 1582 936 1583 940
rect 1587 936 1588 940
rect 1582 935 1588 936
rect 1542 934 1548 935
rect 1536 928 1563 930
rect 167 927 173 928
rect 110 923 116 924
rect 110 919 111 923
rect 115 919 116 923
rect 167 923 168 927
rect 172 926 173 927
rect 188 926 190 928
rect 172 924 190 926
rect 207 927 213 928
rect 172 923 173 924
rect 167 922 173 923
rect 207 923 208 927
rect 212 923 213 927
rect 207 922 213 923
rect 262 927 269 928
rect 262 923 263 927
rect 268 923 269 927
rect 262 922 269 923
rect 319 927 325 928
rect 319 923 320 927
rect 324 923 325 927
rect 319 922 325 923
rect 383 927 389 928
rect 383 923 384 927
rect 388 923 389 927
rect 383 922 389 923
rect 447 927 456 928
rect 447 923 448 927
rect 455 923 456 927
rect 447 922 456 923
rect 511 927 517 928
rect 511 923 512 927
rect 516 926 517 927
rect 545 926 547 928
rect 516 924 547 926
rect 575 927 581 928
rect 516 923 517 924
rect 511 922 517 923
rect 575 923 576 927
rect 580 923 581 927
rect 575 922 581 923
rect 631 927 637 928
rect 631 923 632 927
rect 636 926 637 927
rect 660 926 662 928
rect 636 924 662 926
rect 687 927 693 928
rect 636 923 637 924
rect 631 922 637 923
rect 687 923 688 927
rect 692 926 693 927
rect 712 926 714 928
rect 692 924 714 926
rect 735 927 741 928
rect 692 923 693 924
rect 687 922 693 923
rect 735 923 736 927
rect 740 923 741 927
rect 735 922 741 923
rect 782 927 789 928
rect 782 923 783 927
rect 788 923 789 927
rect 782 922 789 923
rect 831 927 837 928
rect 831 923 832 927
rect 836 926 837 927
rect 860 926 862 928
rect 836 924 862 926
rect 887 927 893 928
rect 836 923 837 924
rect 831 922 837 923
rect 887 923 888 927
rect 892 926 893 927
rect 920 926 922 928
rect 892 924 922 926
rect 951 927 957 928
rect 892 923 893 924
rect 887 922 893 923
rect 951 923 952 927
rect 956 926 957 927
rect 988 926 990 928
rect 956 924 990 926
rect 1023 927 1029 928
rect 956 923 957 924
rect 951 922 957 923
rect 1023 923 1024 927
rect 1028 926 1029 927
rect 1048 926 1050 928
rect 1028 924 1050 926
rect 1095 927 1101 928
rect 1028 923 1029 924
rect 1023 922 1029 923
rect 1095 923 1096 927
rect 1100 923 1101 927
rect 1159 927 1165 928
rect 1159 926 1160 927
rect 1095 922 1101 923
rect 1152 924 1160 926
rect 110 918 116 919
rect 150 921 156 922
rect 150 917 151 921
rect 155 917 156 921
rect 150 916 156 917
rect 190 921 196 922
rect 190 917 191 921
rect 195 917 196 921
rect 190 916 196 917
rect 246 921 252 922
rect 246 917 247 921
rect 251 917 252 921
rect 246 916 252 917
rect 302 921 308 922
rect 302 917 303 921
rect 307 917 308 921
rect 302 916 308 917
rect 366 921 372 922
rect 366 917 367 921
rect 371 917 372 921
rect 366 916 372 917
rect 430 921 436 922
rect 430 917 431 921
rect 435 917 436 921
rect 430 916 436 917
rect 494 921 500 922
rect 494 917 495 921
rect 499 917 500 921
rect 494 916 500 917
rect 558 921 564 922
rect 558 917 559 921
rect 563 917 564 921
rect 558 916 564 917
rect 614 921 620 922
rect 614 917 615 921
rect 619 917 620 921
rect 614 916 620 917
rect 670 921 676 922
rect 670 917 671 921
rect 675 917 676 921
rect 670 916 676 917
rect 718 921 724 922
rect 718 917 719 921
rect 723 917 724 921
rect 718 916 724 917
rect 766 921 772 922
rect 766 917 767 921
rect 771 917 772 921
rect 766 916 772 917
rect 814 921 820 922
rect 814 917 815 921
rect 819 917 820 921
rect 814 916 820 917
rect 870 921 876 922
rect 870 917 871 921
rect 875 917 876 921
rect 870 916 876 917
rect 934 921 940 922
rect 934 917 935 921
rect 939 917 940 921
rect 934 916 940 917
rect 1006 921 1012 922
rect 1006 917 1007 921
rect 1011 917 1012 921
rect 1006 916 1012 917
rect 1078 921 1084 922
rect 1078 917 1079 921
rect 1083 917 1084 921
rect 1078 916 1084 917
rect 1142 921 1148 922
rect 1142 917 1143 921
rect 1147 917 1148 921
rect 1142 916 1148 917
rect 847 915 853 916
rect 550 911 556 912
rect 550 907 551 911
rect 555 910 556 911
rect 847 911 848 915
rect 852 914 853 915
rect 1152 914 1154 924
rect 1159 923 1160 924
rect 1164 923 1165 927
rect 1159 922 1165 923
rect 1223 927 1229 928
rect 1223 923 1224 927
rect 1228 926 1229 927
rect 1256 926 1258 928
rect 1228 924 1258 926
rect 1287 927 1293 928
rect 1228 923 1229 924
rect 1223 922 1229 923
rect 1287 923 1288 927
rect 1292 926 1293 927
rect 1316 926 1318 928
rect 1292 924 1318 926
rect 1343 927 1349 928
rect 1292 923 1293 924
rect 1287 922 1293 923
rect 1343 923 1344 927
rect 1348 926 1349 927
rect 1366 927 1372 928
rect 1366 926 1367 927
rect 1348 924 1367 926
rect 1348 923 1349 924
rect 1343 922 1349 923
rect 1366 923 1367 924
rect 1371 923 1372 927
rect 1366 922 1372 923
rect 1391 927 1397 928
rect 1391 923 1392 927
rect 1396 926 1397 927
rect 1416 926 1418 928
rect 1396 924 1418 926
rect 1439 927 1445 928
rect 1396 923 1397 924
rect 1391 922 1397 923
rect 1439 923 1440 927
rect 1444 923 1445 927
rect 1439 922 1445 923
rect 1487 927 1493 928
rect 1487 923 1488 927
rect 1492 926 1493 927
rect 1498 927 1504 928
rect 1498 926 1499 927
rect 1492 924 1499 926
rect 1492 923 1493 924
rect 1487 922 1493 923
rect 1498 923 1499 924
rect 1503 923 1504 927
rect 1527 927 1533 928
rect 1527 926 1528 927
rect 1498 922 1504 923
rect 1520 924 1528 926
rect 1206 921 1212 922
rect 1206 917 1207 921
rect 1211 917 1212 921
rect 1206 916 1212 917
rect 1270 921 1276 922
rect 1270 917 1271 921
rect 1275 917 1276 921
rect 1270 916 1276 917
rect 1326 921 1332 922
rect 1326 917 1327 921
rect 1331 917 1332 921
rect 1326 916 1332 917
rect 1374 921 1380 922
rect 1374 917 1375 921
rect 1379 917 1380 921
rect 1374 916 1380 917
rect 1422 921 1428 922
rect 1422 917 1423 921
rect 1427 917 1428 921
rect 1422 916 1428 917
rect 1470 921 1476 922
rect 1470 917 1471 921
rect 1475 917 1476 921
rect 1470 916 1476 917
rect 1510 921 1516 922
rect 1510 917 1511 921
rect 1515 917 1516 921
rect 1510 916 1516 917
rect 1520 914 1522 924
rect 1527 923 1528 924
rect 1532 923 1533 927
rect 1527 922 1533 923
rect 1559 927 1565 928
rect 1559 923 1560 927
rect 1564 923 1565 927
rect 1559 922 1565 923
rect 1582 923 1588 924
rect 1542 921 1548 922
rect 1542 917 1543 921
rect 1547 917 1548 921
rect 1582 919 1583 923
rect 1587 919 1588 923
rect 1582 918 1588 919
rect 1542 916 1548 917
rect 852 912 1154 914
rect 1459 912 1522 914
rect 852 911 853 912
rect 847 910 853 911
rect 1459 910 1461 912
rect 1526 911 1532 912
rect 1526 910 1527 911
rect 555 908 750 910
rect 873 908 1155 910
rect 1459 908 1527 910
rect 555 907 556 908
rect 550 906 556 907
rect 134 903 140 904
rect 110 901 116 902
rect 110 897 111 901
rect 115 897 116 901
rect 134 899 135 903
rect 139 899 140 903
rect 134 898 140 899
rect 166 903 172 904
rect 166 899 167 903
rect 171 899 172 903
rect 166 898 172 899
rect 222 903 228 904
rect 222 899 223 903
rect 227 899 228 903
rect 222 898 228 899
rect 278 903 284 904
rect 278 899 279 903
rect 283 899 284 903
rect 278 898 284 899
rect 334 903 340 904
rect 334 899 335 903
rect 339 899 340 903
rect 334 898 340 899
rect 390 903 396 904
rect 390 899 391 903
rect 395 899 396 903
rect 390 898 396 899
rect 446 903 452 904
rect 446 899 447 903
rect 451 899 452 903
rect 446 898 452 899
rect 502 903 508 904
rect 502 899 503 903
rect 507 899 508 903
rect 502 898 508 899
rect 558 903 564 904
rect 558 899 559 903
rect 563 899 564 903
rect 558 898 564 899
rect 622 903 628 904
rect 622 899 623 903
rect 627 899 628 903
rect 622 898 628 899
rect 694 903 700 904
rect 694 899 695 903
rect 699 899 700 903
rect 694 898 700 899
rect 110 896 116 897
rect 150 895 157 896
rect 150 891 151 895
rect 156 891 157 895
rect 183 895 189 896
rect 183 894 184 895
rect 150 890 157 891
rect 176 892 184 894
rect 134 885 140 886
rect 110 884 116 885
rect 110 880 111 884
rect 115 880 116 884
rect 134 881 135 885
rect 139 881 140 885
rect 134 880 140 881
rect 166 885 172 886
rect 166 881 167 885
rect 171 881 172 885
rect 166 880 172 881
rect 110 879 116 880
rect 151 879 157 880
rect 151 875 152 879
rect 156 878 157 879
rect 176 878 178 892
rect 183 891 184 892
rect 188 891 189 895
rect 239 895 245 896
rect 239 894 240 895
rect 183 890 189 891
rect 212 892 240 894
rect 156 876 178 878
rect 183 879 189 880
rect 156 875 157 876
rect 151 874 157 875
rect 183 875 184 879
rect 188 878 189 879
rect 212 878 214 892
rect 239 891 240 892
rect 244 891 245 895
rect 239 890 245 891
rect 295 895 301 896
rect 295 891 296 895
rect 300 894 301 895
rect 318 895 324 896
rect 318 894 319 895
rect 300 892 319 894
rect 300 891 301 892
rect 295 890 301 891
rect 318 891 319 892
rect 323 891 324 895
rect 351 895 357 896
rect 351 894 352 895
rect 318 890 324 891
rect 328 892 352 894
rect 222 885 228 886
rect 222 881 223 885
rect 227 881 228 885
rect 222 880 228 881
rect 278 885 284 886
rect 278 881 279 885
rect 283 881 284 885
rect 278 880 284 881
rect 188 876 214 878
rect 239 879 245 880
rect 188 875 189 876
rect 183 874 189 875
rect 239 875 240 879
rect 244 878 245 879
rect 262 879 268 880
rect 262 878 263 879
rect 244 876 263 878
rect 244 875 245 876
rect 239 874 245 875
rect 262 875 263 876
rect 267 875 268 879
rect 262 874 268 875
rect 295 879 301 880
rect 295 875 296 879
rect 300 878 301 879
rect 328 878 330 892
rect 351 891 352 892
rect 356 891 357 895
rect 407 895 413 896
rect 407 894 408 895
rect 351 890 357 891
rect 384 892 408 894
rect 334 885 340 886
rect 334 881 335 885
rect 339 881 340 885
rect 334 880 340 881
rect 300 876 330 878
rect 351 879 357 880
rect 300 875 301 876
rect 295 874 301 875
rect 351 875 352 879
rect 356 878 357 879
rect 384 878 386 892
rect 407 891 408 892
rect 412 891 413 895
rect 407 890 413 891
rect 463 895 469 896
rect 463 891 464 895
rect 468 894 469 895
rect 519 895 525 896
rect 468 892 494 894
rect 468 891 469 892
rect 463 890 469 891
rect 390 885 396 886
rect 390 881 391 885
rect 395 881 396 885
rect 390 880 396 881
rect 446 885 452 886
rect 446 881 447 885
rect 451 881 452 885
rect 446 880 452 881
rect 407 879 413 880
rect 407 878 408 879
rect 356 876 386 878
rect 388 876 408 878
rect 356 875 357 876
rect 351 874 357 875
rect 367 871 373 872
rect 150 867 157 868
rect 110 864 116 865
rect 110 860 111 864
rect 115 860 116 864
rect 110 859 116 860
rect 134 863 140 864
rect 134 859 135 863
rect 139 859 140 863
rect 150 863 151 867
rect 156 863 157 867
rect 183 867 189 868
rect 183 866 184 867
rect 176 864 184 866
rect 150 862 157 863
rect 166 863 172 864
rect 134 858 140 859
rect 166 859 167 863
rect 171 859 172 863
rect 166 858 172 859
rect 176 854 178 864
rect 183 863 184 864
rect 188 863 189 867
rect 223 867 229 868
rect 223 866 224 867
rect 216 864 224 866
rect 183 862 189 863
rect 206 863 212 864
rect 206 859 207 863
rect 211 859 212 863
rect 206 858 212 859
rect 216 854 218 864
rect 223 863 224 864
rect 228 863 229 867
rect 266 867 277 868
rect 223 862 229 863
rect 254 863 260 864
rect 254 859 255 863
rect 259 859 260 863
rect 266 863 267 867
rect 271 863 272 867
rect 276 863 277 867
rect 319 867 325 868
rect 319 866 320 867
rect 312 864 320 866
rect 266 862 277 863
rect 302 863 308 864
rect 254 858 260 859
rect 302 859 303 863
rect 307 859 308 863
rect 302 858 308 859
rect 312 854 314 864
rect 319 863 320 864
rect 324 863 325 867
rect 359 867 365 868
rect 359 866 360 867
rect 352 864 360 866
rect 319 862 325 863
rect 342 863 348 864
rect 342 859 343 863
rect 347 859 348 863
rect 342 858 348 859
rect 352 854 354 864
rect 359 863 360 864
rect 364 863 365 867
rect 367 867 368 871
rect 372 870 373 871
rect 388 870 390 876
rect 407 875 408 876
rect 412 875 413 879
rect 407 874 413 875
rect 463 879 469 880
rect 463 875 464 879
rect 468 878 469 879
rect 482 879 488 880
rect 482 878 483 879
rect 468 876 483 878
rect 468 875 469 876
rect 463 874 469 875
rect 482 875 483 876
rect 487 875 488 879
rect 492 878 494 892
rect 519 891 520 895
rect 524 894 525 895
rect 575 895 581 896
rect 524 892 550 894
rect 524 891 525 892
rect 519 890 525 891
rect 502 885 508 886
rect 502 881 503 885
rect 507 881 508 885
rect 502 880 508 881
rect 519 879 525 880
rect 519 878 520 879
rect 492 876 520 878
rect 482 874 488 875
rect 519 875 520 876
rect 524 875 525 879
rect 548 878 550 892
rect 575 891 576 895
rect 580 894 581 895
rect 639 895 645 896
rect 580 892 634 894
rect 580 891 581 892
rect 575 890 581 891
rect 558 885 564 886
rect 558 881 559 885
rect 563 881 564 885
rect 558 880 564 881
rect 622 885 628 886
rect 622 881 623 885
rect 627 881 628 885
rect 622 880 628 881
rect 575 879 581 880
rect 575 878 576 879
rect 548 876 576 878
rect 519 874 525 875
rect 575 875 576 876
rect 580 875 581 879
rect 632 878 634 892
rect 639 891 640 895
rect 644 894 645 895
rect 711 895 717 896
rect 644 892 678 894
rect 644 891 645 892
rect 639 890 645 891
rect 639 879 645 880
rect 639 878 640 879
rect 632 876 640 878
rect 575 874 581 875
rect 639 875 640 876
rect 644 875 645 879
rect 676 878 678 892
rect 711 891 712 895
rect 716 894 717 895
rect 748 894 750 908
rect 871 907 877 908
rect 758 903 764 904
rect 758 899 759 903
rect 763 899 764 903
rect 758 898 764 899
rect 822 903 828 904
rect 822 899 823 903
rect 827 899 828 903
rect 871 903 872 907
rect 876 903 877 907
rect 871 902 877 903
rect 886 903 892 904
rect 822 898 828 899
rect 886 899 887 903
rect 891 899 892 903
rect 886 898 892 899
rect 950 903 956 904
rect 950 899 951 903
rect 955 899 956 903
rect 950 898 956 899
rect 1014 903 1020 904
rect 1014 899 1015 903
rect 1019 899 1020 903
rect 1014 898 1020 899
rect 1078 903 1084 904
rect 1078 899 1079 903
rect 1083 899 1084 903
rect 1078 898 1084 899
rect 1134 903 1140 904
rect 1134 899 1135 903
rect 1139 899 1140 903
rect 1134 898 1140 899
rect 1153 896 1155 908
rect 1526 907 1527 908
rect 1531 907 1532 911
rect 1526 906 1532 907
rect 1190 903 1196 904
rect 1190 899 1191 903
rect 1195 899 1196 903
rect 1190 898 1196 899
rect 1246 903 1252 904
rect 1246 899 1247 903
rect 1251 899 1252 903
rect 1246 898 1252 899
rect 1302 903 1308 904
rect 1302 899 1303 903
rect 1307 899 1308 903
rect 1302 898 1308 899
rect 1358 903 1364 904
rect 1358 899 1359 903
rect 1363 899 1364 903
rect 1358 898 1364 899
rect 1406 903 1412 904
rect 1406 899 1407 903
rect 1411 899 1412 903
rect 1406 898 1412 899
rect 1454 903 1460 904
rect 1454 899 1455 903
rect 1459 899 1460 903
rect 1454 898 1460 899
rect 1510 903 1516 904
rect 1510 899 1511 903
rect 1515 899 1516 903
rect 1510 898 1516 899
rect 1542 903 1548 904
rect 1542 899 1543 903
rect 1547 899 1548 903
rect 1542 898 1548 899
rect 1582 901 1588 902
rect 1582 897 1583 901
rect 1587 897 1588 901
rect 1582 896 1588 897
rect 775 895 781 896
rect 775 894 776 895
rect 716 892 746 894
rect 748 892 776 894
rect 716 891 717 892
rect 711 890 717 891
rect 694 885 700 886
rect 694 881 695 885
rect 699 881 700 885
rect 694 880 700 881
rect 711 879 717 880
rect 711 878 712 879
rect 676 876 712 878
rect 639 874 645 875
rect 711 875 712 876
rect 716 875 717 879
rect 744 878 746 892
rect 775 891 776 892
rect 780 891 781 895
rect 775 890 781 891
rect 839 895 845 896
rect 839 891 840 895
rect 844 894 845 895
rect 903 895 909 896
rect 844 892 874 894
rect 844 891 845 892
rect 839 890 845 891
rect 758 885 764 886
rect 758 881 759 885
rect 763 881 764 885
rect 758 880 764 881
rect 822 885 828 886
rect 822 881 823 885
rect 827 881 828 885
rect 822 880 828 881
rect 775 879 781 880
rect 775 878 776 879
rect 744 876 776 878
rect 711 874 717 875
rect 775 875 776 876
rect 780 875 781 879
rect 775 874 781 875
rect 839 879 845 880
rect 839 875 840 879
rect 844 878 845 879
rect 847 879 853 880
rect 847 878 848 879
rect 844 876 848 878
rect 844 875 845 876
rect 839 874 845 875
rect 847 875 848 876
rect 852 875 853 879
rect 872 878 874 892
rect 903 891 904 895
rect 908 894 909 895
rect 967 895 973 896
rect 908 892 938 894
rect 908 891 909 892
rect 903 890 909 891
rect 886 885 892 886
rect 886 881 887 885
rect 891 881 892 885
rect 886 880 892 881
rect 903 879 909 880
rect 903 878 904 879
rect 872 876 904 878
rect 847 874 853 875
rect 903 875 904 876
rect 908 875 909 879
rect 936 878 938 892
rect 967 891 968 895
rect 972 894 973 895
rect 1031 895 1037 896
rect 972 892 1026 894
rect 972 891 973 892
rect 967 890 973 891
rect 950 885 956 886
rect 950 881 951 885
rect 955 881 956 885
rect 950 880 956 881
rect 1014 885 1020 886
rect 1014 881 1015 885
rect 1019 881 1020 885
rect 1014 880 1020 881
rect 967 879 973 880
rect 967 878 968 879
rect 936 876 968 878
rect 903 874 909 875
rect 967 875 968 876
rect 972 875 973 879
rect 1024 878 1026 892
rect 1031 891 1032 895
rect 1036 894 1037 895
rect 1095 895 1101 896
rect 1036 892 1066 894
rect 1036 891 1037 892
rect 1031 890 1037 891
rect 1031 879 1037 880
rect 1031 878 1032 879
rect 1024 876 1032 878
rect 967 874 973 875
rect 1031 875 1032 876
rect 1036 875 1037 879
rect 1064 878 1066 892
rect 1095 891 1096 895
rect 1100 894 1101 895
rect 1151 895 1157 896
rect 1100 892 1146 894
rect 1100 891 1101 892
rect 1095 890 1101 891
rect 1078 885 1084 886
rect 1078 881 1079 885
rect 1083 881 1084 885
rect 1078 880 1084 881
rect 1134 885 1140 886
rect 1134 881 1135 885
rect 1139 881 1140 885
rect 1134 880 1140 881
rect 1095 879 1101 880
rect 1095 878 1096 879
rect 1064 876 1096 878
rect 1031 874 1037 875
rect 1095 875 1096 876
rect 1100 875 1101 879
rect 1144 878 1146 892
rect 1151 891 1152 895
rect 1156 891 1157 895
rect 1151 890 1157 891
rect 1207 895 1213 896
rect 1207 891 1208 895
rect 1212 894 1213 895
rect 1263 895 1269 896
rect 1212 892 1258 894
rect 1212 891 1213 892
rect 1207 890 1213 891
rect 1190 885 1196 886
rect 1190 881 1191 885
rect 1195 881 1196 885
rect 1190 880 1196 881
rect 1246 885 1252 886
rect 1246 881 1247 885
rect 1251 881 1252 885
rect 1246 880 1252 881
rect 1151 879 1157 880
rect 1151 878 1152 879
rect 1144 876 1152 878
rect 1095 874 1101 875
rect 1151 875 1152 876
rect 1156 875 1157 879
rect 1151 874 1157 875
rect 1207 879 1213 880
rect 1207 875 1208 879
rect 1212 878 1213 879
rect 1256 878 1258 892
rect 1263 891 1264 895
rect 1268 894 1269 895
rect 1278 895 1284 896
rect 1278 894 1279 895
rect 1268 892 1279 894
rect 1268 891 1269 892
rect 1263 890 1269 891
rect 1278 891 1279 892
rect 1283 891 1284 895
rect 1278 890 1284 891
rect 1286 895 1292 896
rect 1286 891 1287 895
rect 1291 894 1292 895
rect 1319 895 1325 896
rect 1319 894 1320 895
rect 1291 892 1320 894
rect 1291 891 1292 892
rect 1286 890 1292 891
rect 1319 891 1320 892
rect 1324 891 1325 895
rect 1375 895 1381 896
rect 1375 894 1376 895
rect 1319 890 1325 891
rect 1348 892 1376 894
rect 1302 885 1308 886
rect 1302 881 1303 885
rect 1307 881 1308 885
rect 1302 880 1308 881
rect 1263 879 1269 880
rect 1263 878 1264 879
rect 1212 876 1254 878
rect 1256 876 1264 878
rect 1212 875 1213 876
rect 1207 874 1213 875
rect 372 868 390 870
rect 1252 870 1254 876
rect 1263 875 1264 876
rect 1268 875 1269 879
rect 1319 879 1325 880
rect 1263 874 1269 875
rect 1286 875 1292 876
rect 1286 874 1287 875
rect 1272 872 1287 874
rect 1272 870 1274 872
rect 1286 871 1287 872
rect 1291 871 1292 875
rect 1319 875 1320 879
rect 1324 878 1325 879
rect 1348 878 1350 892
rect 1375 891 1376 892
rect 1380 891 1381 895
rect 1375 890 1381 891
rect 1399 895 1405 896
rect 1399 891 1400 895
rect 1404 894 1405 895
rect 1423 895 1429 896
rect 1423 894 1424 895
rect 1404 892 1424 894
rect 1404 891 1405 892
rect 1399 890 1405 891
rect 1423 891 1424 892
rect 1428 891 1429 895
rect 1471 895 1477 896
rect 1471 894 1472 895
rect 1423 890 1429 891
rect 1441 892 1472 894
rect 1358 885 1364 886
rect 1358 881 1359 885
rect 1363 881 1364 885
rect 1358 880 1364 881
rect 1406 885 1412 886
rect 1406 881 1407 885
rect 1411 881 1412 885
rect 1406 880 1412 881
rect 1324 876 1350 878
rect 1366 879 1372 880
rect 1324 875 1325 876
rect 1319 874 1325 875
rect 1366 875 1367 879
rect 1371 878 1372 879
rect 1375 879 1381 880
rect 1375 878 1376 879
rect 1371 876 1376 878
rect 1371 875 1372 876
rect 1366 874 1372 875
rect 1375 875 1376 876
rect 1380 875 1381 879
rect 1375 874 1381 875
rect 1423 879 1429 880
rect 1423 875 1424 879
rect 1428 878 1429 879
rect 1441 878 1443 892
rect 1471 891 1472 892
rect 1476 891 1477 895
rect 1471 890 1477 891
rect 1527 895 1533 896
rect 1527 891 1528 895
rect 1532 894 1533 895
rect 1558 895 1565 896
rect 1532 892 1554 894
rect 1532 891 1533 892
rect 1527 890 1533 891
rect 1454 885 1460 886
rect 1454 881 1455 885
rect 1459 881 1460 885
rect 1454 880 1460 881
rect 1510 885 1516 886
rect 1510 881 1511 885
rect 1515 881 1516 885
rect 1510 880 1516 881
rect 1542 885 1548 886
rect 1542 881 1543 885
rect 1547 881 1548 885
rect 1542 880 1548 881
rect 1428 876 1443 878
rect 1471 879 1477 880
rect 1428 875 1429 876
rect 1423 874 1429 875
rect 1471 875 1472 879
rect 1476 878 1477 879
rect 1494 879 1500 880
rect 1494 878 1495 879
rect 1476 876 1495 878
rect 1476 875 1477 876
rect 1471 874 1477 875
rect 1494 875 1495 876
rect 1499 875 1500 879
rect 1494 874 1500 875
rect 1526 879 1533 880
rect 1526 875 1527 879
rect 1532 875 1533 879
rect 1552 878 1554 892
rect 1558 891 1559 895
rect 1564 891 1565 895
rect 1558 890 1565 891
rect 1582 884 1588 885
rect 1582 880 1583 884
rect 1587 880 1588 884
rect 1559 879 1565 880
rect 1582 879 1588 880
rect 1559 878 1560 879
rect 1552 876 1560 878
rect 1526 874 1533 875
rect 1559 875 1560 876
rect 1564 875 1565 879
rect 1559 874 1565 875
rect 1286 870 1292 871
rect 1252 868 1274 870
rect 372 867 373 868
rect 367 866 373 867
rect 399 867 405 868
rect 359 862 365 863
rect 382 863 388 864
rect 382 859 383 863
rect 387 859 388 863
rect 399 863 400 867
rect 404 866 405 867
rect 415 867 421 868
rect 415 866 416 867
rect 404 864 416 866
rect 404 863 405 864
rect 399 862 405 863
rect 415 863 416 864
rect 420 863 421 867
rect 455 867 461 868
rect 455 866 456 867
rect 448 864 456 866
rect 415 862 421 863
rect 438 863 444 864
rect 382 858 388 859
rect 438 859 439 863
rect 443 859 444 863
rect 438 858 444 859
rect 448 854 450 864
rect 455 863 456 864
rect 460 863 461 867
rect 527 867 533 868
rect 527 866 528 867
rect 520 864 528 866
rect 455 862 461 863
rect 510 863 516 864
rect 510 859 511 863
rect 515 859 516 863
rect 510 858 516 859
rect 520 854 522 864
rect 527 863 528 864
rect 532 863 533 867
rect 607 867 613 868
rect 607 866 608 867
rect 600 864 608 866
rect 527 862 533 863
rect 590 863 596 864
rect 590 859 591 863
rect 595 859 596 863
rect 590 858 596 859
rect 600 854 602 864
rect 607 863 608 864
rect 612 863 613 867
rect 695 867 701 868
rect 695 866 696 867
rect 688 864 696 866
rect 607 862 613 863
rect 678 863 684 864
rect 678 859 679 863
rect 683 859 684 863
rect 678 858 684 859
rect 688 854 690 864
rect 695 863 696 864
rect 700 863 701 867
rect 783 867 789 868
rect 783 866 784 867
rect 776 864 784 866
rect 695 862 701 863
rect 766 863 772 864
rect 766 859 767 863
rect 771 859 772 863
rect 766 858 772 859
rect 776 854 778 864
rect 783 863 784 864
rect 788 863 789 867
rect 863 867 869 868
rect 783 862 789 863
rect 846 863 852 864
rect 846 859 847 863
rect 851 859 852 863
rect 863 863 864 867
rect 868 866 869 867
rect 871 867 877 868
rect 871 866 872 867
rect 868 864 872 866
rect 868 863 869 864
rect 863 862 869 863
rect 871 863 872 864
rect 876 863 877 867
rect 935 867 941 868
rect 935 866 936 867
rect 928 864 936 866
rect 871 862 877 863
rect 918 863 924 864
rect 846 858 852 859
rect 918 859 919 863
rect 923 859 924 863
rect 918 858 924 859
rect 928 854 930 864
rect 935 863 936 864
rect 940 863 941 867
rect 999 867 1005 868
rect 999 866 1000 867
rect 992 864 1000 866
rect 935 862 941 863
rect 982 863 988 864
rect 982 859 983 863
rect 987 859 988 863
rect 982 858 988 859
rect 992 854 994 864
rect 999 863 1000 864
rect 1004 863 1005 867
rect 1055 867 1061 868
rect 1055 866 1056 867
rect 1048 864 1056 866
rect 999 862 1005 863
rect 1038 863 1044 864
rect 1038 859 1039 863
rect 1043 859 1044 863
rect 1038 858 1044 859
rect 1048 854 1050 864
rect 1055 863 1056 864
rect 1060 863 1061 867
rect 1111 867 1117 868
rect 1111 866 1112 867
rect 1104 864 1112 866
rect 1055 862 1061 863
rect 1094 863 1100 864
rect 1094 859 1095 863
rect 1099 859 1100 863
rect 1094 858 1100 859
rect 1104 854 1106 864
rect 1111 863 1112 864
rect 1116 863 1117 867
rect 1167 867 1173 868
rect 1111 862 1117 863
rect 1150 863 1156 864
rect 1150 859 1151 863
rect 1155 859 1156 863
rect 1167 863 1168 867
rect 1172 866 1173 867
rect 1223 867 1229 868
rect 1172 864 1202 866
rect 1172 863 1173 864
rect 1167 862 1173 863
rect 1150 858 1156 859
rect 164 852 178 854
rect 204 852 218 854
rect 273 852 314 854
rect 321 852 354 854
rect 428 852 450 854
rect 492 852 522 854
rect 568 852 602 854
rect 609 852 690 854
rect 740 852 778 854
rect 876 852 930 854
rect 937 852 994 854
rect 1001 852 1050 854
rect 1057 852 1106 854
rect 1127 855 1133 856
rect 151 851 157 852
rect 110 847 116 848
rect 110 843 111 847
rect 115 843 116 847
rect 151 847 152 851
rect 156 850 157 851
rect 164 850 166 852
rect 156 848 166 850
rect 183 851 189 852
rect 156 847 157 848
rect 151 846 157 847
rect 183 847 184 851
rect 188 850 189 851
rect 204 850 206 852
rect 188 848 206 850
rect 222 851 229 852
rect 188 847 189 848
rect 183 846 189 847
rect 222 847 223 851
rect 228 847 229 851
rect 222 846 229 847
rect 271 851 277 852
rect 271 847 272 851
rect 276 847 277 851
rect 271 846 277 847
rect 319 851 325 852
rect 319 847 320 851
rect 324 847 325 851
rect 319 846 325 847
rect 359 851 365 852
rect 359 847 360 851
rect 364 850 365 851
rect 367 851 373 852
rect 367 850 368 851
rect 364 848 368 850
rect 364 847 365 848
rect 359 846 365 847
rect 367 847 368 848
rect 372 847 373 851
rect 367 846 373 847
rect 399 851 405 852
rect 399 847 400 851
rect 404 850 405 851
rect 428 850 430 852
rect 404 848 430 850
rect 455 851 461 852
rect 404 847 405 848
rect 399 846 405 847
rect 455 847 456 851
rect 460 850 461 851
rect 492 850 494 852
rect 460 848 494 850
rect 527 851 533 852
rect 460 847 461 848
rect 455 846 461 847
rect 527 847 528 851
rect 532 850 533 851
rect 568 850 570 852
rect 532 848 570 850
rect 607 851 613 852
rect 532 847 533 848
rect 527 846 533 847
rect 607 847 608 851
rect 612 847 613 851
rect 607 846 613 847
rect 695 851 701 852
rect 695 847 696 851
rect 700 850 701 851
rect 740 850 742 852
rect 783 851 789 852
rect 783 850 784 851
rect 700 848 742 850
rect 776 848 784 850
rect 700 847 701 848
rect 695 846 701 847
rect 110 842 116 843
rect 134 845 140 846
rect 134 841 135 845
rect 139 841 140 845
rect 134 840 140 841
rect 166 845 172 846
rect 166 841 167 845
rect 171 841 172 845
rect 166 840 172 841
rect 206 845 212 846
rect 206 841 207 845
rect 211 841 212 845
rect 206 840 212 841
rect 254 845 260 846
rect 254 841 255 845
rect 259 841 260 845
rect 254 840 260 841
rect 302 845 308 846
rect 302 841 303 845
rect 307 841 308 845
rect 302 840 308 841
rect 342 845 348 846
rect 342 841 343 845
rect 347 841 348 845
rect 342 840 348 841
rect 382 845 388 846
rect 382 841 383 845
rect 387 841 388 845
rect 382 840 388 841
rect 438 845 444 846
rect 438 841 439 845
rect 443 841 444 845
rect 510 845 516 846
rect 438 840 444 841
rect 482 843 488 844
rect 482 839 483 843
rect 487 839 488 843
rect 510 841 511 845
rect 515 841 516 845
rect 510 840 516 841
rect 590 845 596 846
rect 590 841 591 845
rect 595 841 596 845
rect 590 840 596 841
rect 678 845 684 846
rect 678 841 679 845
rect 683 841 684 845
rect 678 840 684 841
rect 766 845 772 846
rect 766 841 767 845
rect 771 841 772 845
rect 766 840 772 841
rect 482 838 488 839
rect 776 838 778 848
rect 783 847 784 848
rect 788 847 789 851
rect 783 846 789 847
rect 863 851 869 852
rect 863 847 864 851
rect 868 850 869 851
rect 876 850 878 852
rect 868 848 878 850
rect 935 851 941 852
rect 868 847 869 848
rect 863 846 869 847
rect 935 847 936 851
rect 940 847 941 851
rect 935 846 941 847
rect 999 851 1005 852
rect 999 847 1000 851
rect 1004 847 1005 851
rect 999 846 1005 847
rect 1055 851 1061 852
rect 1055 847 1056 851
rect 1060 847 1061 851
rect 1111 851 1117 852
rect 1111 850 1112 851
rect 1055 846 1061 847
rect 1104 848 1112 850
rect 846 845 852 846
rect 846 841 847 845
rect 851 841 852 845
rect 846 840 852 841
rect 918 845 924 846
rect 918 841 919 845
rect 923 841 924 845
rect 918 840 924 841
rect 982 845 988 846
rect 982 841 983 845
rect 987 841 988 845
rect 982 840 988 841
rect 1038 845 1044 846
rect 1038 841 1039 845
rect 1043 841 1044 845
rect 1038 840 1044 841
rect 1094 845 1100 846
rect 1094 841 1095 845
rect 1099 841 1100 845
rect 1094 840 1100 841
rect 484 836 778 838
rect 1018 839 1024 840
rect 447 835 453 836
rect 447 831 448 835
rect 452 834 453 835
rect 1018 835 1019 839
rect 1023 838 1024 839
rect 1104 838 1106 848
rect 1111 847 1112 848
rect 1116 847 1117 851
rect 1127 851 1128 855
rect 1132 854 1133 855
rect 1200 854 1202 864
rect 1206 863 1212 864
rect 1206 859 1207 863
rect 1211 859 1212 863
rect 1223 863 1224 867
rect 1228 866 1229 867
rect 1239 867 1245 868
rect 1239 866 1240 867
rect 1228 864 1240 866
rect 1228 863 1229 864
rect 1223 862 1229 863
rect 1239 863 1240 864
rect 1244 863 1245 867
rect 1278 867 1285 868
rect 1239 862 1245 863
rect 1262 863 1268 864
rect 1206 858 1212 859
rect 1262 859 1263 863
rect 1267 859 1268 863
rect 1278 863 1279 867
rect 1284 863 1285 867
rect 1343 867 1349 868
rect 1343 866 1344 867
rect 1336 864 1344 866
rect 1278 862 1285 863
rect 1326 863 1332 864
rect 1262 858 1268 859
rect 1326 859 1327 863
rect 1331 859 1332 863
rect 1326 858 1332 859
rect 1336 854 1338 864
rect 1343 863 1344 864
rect 1348 863 1349 867
rect 1415 867 1421 868
rect 1415 866 1416 867
rect 1408 864 1416 866
rect 1343 862 1349 863
rect 1398 863 1404 864
rect 1398 859 1399 863
rect 1403 859 1404 863
rect 1398 858 1404 859
rect 1408 854 1410 864
rect 1415 863 1416 864
rect 1420 863 1421 867
rect 1495 867 1501 868
rect 1415 862 1421 863
rect 1478 863 1484 864
rect 1478 859 1479 863
rect 1483 859 1484 863
rect 1495 863 1496 867
rect 1500 866 1501 867
rect 1558 867 1565 868
rect 1500 864 1538 866
rect 1500 863 1501 864
rect 1495 862 1501 863
rect 1478 858 1484 859
rect 1132 852 1162 854
rect 1200 852 1218 854
rect 1313 852 1338 854
rect 1376 852 1410 854
rect 1536 854 1538 864
rect 1542 863 1548 864
rect 1542 859 1543 863
rect 1547 859 1548 863
rect 1558 863 1559 867
rect 1564 863 1565 867
rect 1558 862 1565 863
rect 1582 864 1588 865
rect 1582 860 1583 864
rect 1587 860 1588 864
rect 1582 859 1588 860
rect 1542 858 1548 859
rect 1536 852 1563 854
rect 1132 851 1133 852
rect 1127 850 1133 851
rect 1160 850 1162 852
rect 1167 851 1173 852
rect 1167 850 1168 851
rect 1160 848 1168 850
rect 1111 846 1117 847
rect 1167 847 1168 848
rect 1172 847 1173 851
rect 1216 850 1218 852
rect 1223 851 1229 852
rect 1223 850 1224 851
rect 1216 848 1224 850
rect 1167 846 1173 847
rect 1223 847 1224 848
rect 1228 847 1229 851
rect 1223 846 1229 847
rect 1279 851 1285 852
rect 1279 847 1280 851
rect 1284 850 1285 851
rect 1313 850 1315 852
rect 1284 848 1315 850
rect 1343 851 1349 852
rect 1284 847 1285 848
rect 1279 846 1285 847
rect 1343 847 1344 851
rect 1348 850 1349 851
rect 1376 850 1378 852
rect 1415 851 1421 852
rect 1415 850 1416 851
rect 1348 848 1378 850
rect 1408 848 1416 850
rect 1348 847 1349 848
rect 1343 846 1349 847
rect 1150 845 1156 846
rect 1150 841 1151 845
rect 1155 841 1156 845
rect 1150 840 1156 841
rect 1206 845 1212 846
rect 1206 841 1207 845
rect 1211 841 1212 845
rect 1206 840 1212 841
rect 1262 845 1268 846
rect 1262 841 1263 845
rect 1267 841 1268 845
rect 1262 840 1268 841
rect 1326 845 1332 846
rect 1326 841 1327 845
rect 1331 841 1332 845
rect 1326 840 1332 841
rect 1398 845 1404 846
rect 1398 841 1399 845
rect 1403 841 1404 845
rect 1398 840 1404 841
rect 1023 836 1106 838
rect 1239 839 1245 840
rect 1023 835 1024 836
rect 1018 834 1024 835
rect 1239 835 1240 839
rect 1244 838 1245 839
rect 1408 838 1410 848
rect 1415 847 1416 848
rect 1420 847 1421 851
rect 1415 846 1421 847
rect 1494 851 1501 852
rect 1494 847 1495 851
rect 1500 847 1501 851
rect 1494 846 1501 847
rect 1559 851 1565 852
rect 1559 847 1560 851
rect 1564 847 1565 851
rect 1559 846 1565 847
rect 1582 847 1588 848
rect 1478 845 1484 846
rect 1478 841 1479 845
rect 1483 841 1484 845
rect 1478 840 1484 841
rect 1542 845 1548 846
rect 1542 841 1543 845
rect 1547 841 1548 845
rect 1582 843 1583 847
rect 1587 843 1588 847
rect 1582 842 1588 843
rect 1542 840 1548 841
rect 1244 836 1410 838
rect 1244 835 1245 836
rect 1239 834 1245 835
rect 452 832 522 834
rect 1248 832 1338 834
rect 452 831 453 832
rect 447 830 453 831
rect 134 827 140 828
rect 110 825 116 826
rect 110 821 111 825
rect 115 821 116 825
rect 134 823 135 827
rect 139 823 140 827
rect 134 822 140 823
rect 166 827 172 828
rect 166 823 167 827
rect 171 823 172 827
rect 166 822 172 823
rect 222 827 228 828
rect 222 823 223 827
rect 227 823 228 827
rect 222 822 228 823
rect 286 827 292 828
rect 286 823 287 827
rect 291 823 292 827
rect 286 822 292 823
rect 350 827 356 828
rect 350 823 351 827
rect 355 823 356 827
rect 350 822 356 823
rect 422 827 428 828
rect 422 823 423 827
rect 427 823 428 827
rect 422 822 428 823
rect 494 827 500 828
rect 494 823 495 827
rect 499 823 500 827
rect 494 822 500 823
rect 110 820 116 821
rect 150 819 157 820
rect 150 815 151 819
rect 156 815 157 819
rect 183 819 189 820
rect 183 818 184 819
rect 150 814 157 815
rect 176 816 184 818
rect 134 809 140 810
rect 110 808 116 809
rect 110 804 111 808
rect 115 804 116 808
rect 134 805 135 809
rect 139 805 140 809
rect 134 804 140 805
rect 166 809 172 810
rect 166 805 167 809
rect 171 805 172 809
rect 166 804 172 805
rect 110 803 116 804
rect 151 803 157 804
rect 151 799 152 803
rect 156 802 157 803
rect 176 802 178 816
rect 183 815 184 816
rect 188 815 189 819
rect 183 814 189 815
rect 239 819 245 820
rect 239 815 240 819
rect 244 818 245 819
rect 266 819 272 820
rect 266 818 267 819
rect 244 816 267 818
rect 244 815 245 816
rect 239 814 245 815
rect 266 815 267 816
rect 271 815 272 819
rect 303 819 309 820
rect 303 818 304 819
rect 266 814 272 815
rect 280 816 304 818
rect 222 809 228 810
rect 222 805 223 809
rect 227 805 228 809
rect 222 804 228 805
rect 156 800 178 802
rect 183 803 189 804
rect 156 799 157 800
rect 151 798 157 799
rect 183 799 184 803
rect 188 802 189 803
rect 214 803 220 804
rect 214 802 215 803
rect 188 800 215 802
rect 188 799 189 800
rect 183 798 189 799
rect 214 799 215 800
rect 219 799 220 803
rect 214 798 220 799
rect 239 803 245 804
rect 239 799 240 803
rect 244 802 245 803
rect 280 802 282 816
rect 303 815 304 816
rect 308 815 309 819
rect 367 819 373 820
rect 367 818 368 819
rect 303 814 309 815
rect 340 816 368 818
rect 286 809 292 810
rect 286 805 287 809
rect 291 805 292 809
rect 286 804 292 805
rect 244 800 282 802
rect 303 803 309 804
rect 244 799 245 800
rect 239 798 245 799
rect 303 799 304 803
rect 308 802 309 803
rect 340 802 342 816
rect 367 815 368 816
rect 372 815 373 819
rect 367 814 373 815
rect 415 819 421 820
rect 415 815 416 819
rect 420 818 421 819
rect 439 819 445 820
rect 439 818 440 819
rect 420 816 440 818
rect 420 815 421 816
rect 415 814 421 815
rect 439 815 440 816
rect 444 815 445 819
rect 511 819 517 820
rect 511 818 512 819
rect 439 814 445 815
rect 476 816 512 818
rect 350 809 356 810
rect 350 805 351 809
rect 355 805 356 809
rect 350 804 356 805
rect 422 809 428 810
rect 422 805 423 809
rect 427 805 428 809
rect 422 804 428 805
rect 308 800 342 802
rect 367 803 376 804
rect 308 799 309 800
rect 303 798 309 799
rect 367 799 368 803
rect 375 799 376 803
rect 367 798 376 799
rect 439 803 445 804
rect 439 799 440 803
rect 444 802 445 803
rect 476 802 478 816
rect 511 815 512 816
rect 516 815 517 819
rect 520 818 522 832
rect 1246 831 1252 832
rect 566 827 572 828
rect 566 823 567 827
rect 571 823 572 827
rect 566 822 572 823
rect 638 827 644 828
rect 638 823 639 827
rect 643 823 644 827
rect 638 822 644 823
rect 718 827 724 828
rect 718 823 719 827
rect 723 823 724 827
rect 718 822 724 823
rect 790 827 796 828
rect 790 823 791 827
rect 795 823 796 827
rect 790 822 796 823
rect 862 827 868 828
rect 862 823 863 827
rect 867 823 868 827
rect 862 822 868 823
rect 934 827 940 828
rect 934 823 935 827
rect 939 823 940 827
rect 934 822 940 823
rect 998 827 1004 828
rect 998 823 999 827
rect 1003 823 1004 827
rect 998 822 1004 823
rect 1054 827 1060 828
rect 1054 823 1055 827
rect 1059 823 1060 827
rect 1054 822 1060 823
rect 1102 827 1108 828
rect 1102 823 1103 827
rect 1107 823 1108 827
rect 1102 822 1108 823
rect 1142 827 1148 828
rect 1142 823 1143 827
rect 1147 823 1148 827
rect 1142 822 1148 823
rect 1182 827 1188 828
rect 1182 823 1183 827
rect 1187 823 1188 827
rect 1182 822 1188 823
rect 1230 827 1236 828
rect 1230 823 1231 827
rect 1235 823 1236 827
rect 1246 827 1247 831
rect 1251 827 1252 831
rect 1246 826 1252 827
rect 1278 827 1284 828
rect 1230 822 1236 823
rect 1278 823 1279 827
rect 1283 823 1284 827
rect 1278 822 1284 823
rect 1326 827 1332 828
rect 1326 823 1327 827
rect 1331 823 1332 827
rect 1326 822 1332 823
rect 583 819 589 820
rect 583 818 584 819
rect 520 816 584 818
rect 511 814 517 815
rect 583 815 584 816
rect 588 815 589 819
rect 655 819 661 820
rect 655 818 656 819
rect 583 814 589 815
rect 620 816 656 818
rect 494 809 500 810
rect 494 805 495 809
rect 499 805 500 809
rect 494 804 500 805
rect 566 809 572 810
rect 566 805 567 809
rect 571 805 572 809
rect 566 804 572 805
rect 444 800 478 802
rect 502 803 508 804
rect 444 799 445 800
rect 439 798 445 799
rect 502 799 503 803
rect 507 802 508 803
rect 511 803 517 804
rect 511 802 512 803
rect 507 800 512 802
rect 507 799 508 800
rect 502 798 508 799
rect 511 799 512 800
rect 516 799 517 803
rect 511 798 517 799
rect 583 803 589 804
rect 583 799 584 803
rect 588 802 589 803
rect 620 802 622 816
rect 655 815 656 816
rect 660 815 661 819
rect 655 814 661 815
rect 735 819 741 820
rect 735 815 736 819
rect 740 818 741 819
rect 750 819 756 820
rect 750 818 751 819
rect 740 816 751 818
rect 740 815 741 816
rect 735 814 741 815
rect 750 815 751 816
rect 755 815 756 819
rect 807 819 813 820
rect 807 818 808 819
rect 750 814 756 815
rect 772 816 808 818
rect 638 809 644 810
rect 638 805 639 809
rect 643 805 644 809
rect 638 804 644 805
rect 718 809 724 810
rect 718 805 719 809
rect 723 805 724 809
rect 718 804 724 805
rect 588 800 622 802
rect 655 803 661 804
rect 588 799 589 800
rect 583 798 589 799
rect 655 799 656 803
rect 660 802 661 803
rect 686 803 692 804
rect 686 802 687 803
rect 660 800 687 802
rect 660 799 661 800
rect 655 798 661 799
rect 686 799 687 800
rect 691 799 692 803
rect 686 798 692 799
rect 735 803 741 804
rect 735 799 736 803
rect 740 802 741 803
rect 772 802 774 816
rect 807 815 808 816
rect 812 815 813 819
rect 879 819 885 820
rect 879 818 880 819
rect 807 814 813 815
rect 844 816 880 818
rect 790 809 796 810
rect 790 805 791 809
rect 795 805 796 809
rect 790 804 796 805
rect 740 800 774 802
rect 807 803 813 804
rect 740 799 741 800
rect 735 798 741 799
rect 807 799 808 803
rect 812 802 813 803
rect 844 802 846 816
rect 879 815 880 816
rect 884 815 885 819
rect 951 819 957 820
rect 951 818 952 819
rect 879 814 885 815
rect 916 816 952 818
rect 862 809 868 810
rect 862 805 863 809
rect 867 805 868 809
rect 862 804 868 805
rect 812 800 846 802
rect 879 803 885 804
rect 812 799 813 800
rect 807 798 813 799
rect 879 799 880 803
rect 884 802 885 803
rect 916 802 918 816
rect 951 815 952 816
rect 956 815 957 819
rect 951 814 957 815
rect 1015 819 1021 820
rect 1015 815 1016 819
rect 1020 818 1021 819
rect 1071 819 1077 820
rect 1020 816 1046 818
rect 1020 815 1021 816
rect 1015 814 1021 815
rect 934 809 940 810
rect 934 805 935 809
rect 939 805 940 809
rect 934 804 940 805
rect 998 809 1004 810
rect 998 805 999 809
rect 1003 805 1004 809
rect 998 804 1004 805
rect 884 800 918 802
rect 951 803 957 804
rect 884 799 885 800
rect 879 798 885 799
rect 951 799 952 803
rect 956 802 957 803
rect 1006 803 1012 804
rect 1006 802 1007 803
rect 956 800 1007 802
rect 956 799 957 800
rect 951 798 957 799
rect 1006 799 1007 800
rect 1011 799 1012 803
rect 1006 798 1012 799
rect 1015 803 1024 804
rect 1015 799 1016 803
rect 1023 799 1024 803
rect 1044 802 1046 816
rect 1071 815 1072 819
rect 1076 818 1077 819
rect 1086 819 1092 820
rect 1086 818 1087 819
rect 1076 816 1087 818
rect 1076 815 1077 816
rect 1071 814 1077 815
rect 1086 815 1087 816
rect 1091 815 1092 819
rect 1086 814 1092 815
rect 1119 819 1125 820
rect 1119 815 1120 819
rect 1124 818 1125 819
rect 1159 819 1165 820
rect 1124 816 1154 818
rect 1124 815 1125 816
rect 1119 814 1125 815
rect 1054 809 1060 810
rect 1054 805 1055 809
rect 1059 805 1060 809
rect 1054 804 1060 805
rect 1102 809 1108 810
rect 1102 805 1103 809
rect 1107 805 1108 809
rect 1102 804 1108 805
rect 1142 809 1148 810
rect 1142 805 1143 809
rect 1147 805 1148 809
rect 1142 804 1148 805
rect 1071 803 1077 804
rect 1071 802 1072 803
rect 1044 800 1072 802
rect 1015 798 1024 799
rect 1071 799 1072 800
rect 1076 799 1077 803
rect 1119 803 1125 804
rect 1071 798 1077 799
rect 1086 799 1092 800
rect 223 795 229 796
rect 150 791 157 792
rect 110 788 116 789
rect 110 784 111 788
rect 115 784 116 788
rect 110 783 116 784
rect 134 787 140 788
rect 134 783 135 787
rect 139 783 140 787
rect 150 787 151 791
rect 156 787 157 791
rect 183 791 189 792
rect 183 790 184 791
rect 176 788 184 790
rect 150 786 157 787
rect 166 787 172 788
rect 134 782 140 783
rect 166 783 167 787
rect 171 783 172 787
rect 166 782 172 783
rect 176 778 178 788
rect 183 787 184 788
rect 188 787 189 791
rect 215 791 221 792
rect 215 790 216 791
rect 208 788 216 790
rect 183 786 189 787
rect 198 787 204 788
rect 198 783 199 787
rect 203 783 204 787
rect 198 782 204 783
rect 208 778 210 788
rect 215 787 216 788
rect 220 787 221 791
rect 223 791 224 795
rect 228 794 229 795
rect 327 795 333 796
rect 228 792 261 794
rect 228 791 229 792
rect 223 790 229 791
rect 259 790 261 792
rect 263 791 269 792
rect 263 790 264 791
rect 259 788 264 790
rect 215 786 221 787
rect 246 787 252 788
rect 246 783 247 787
rect 251 783 252 787
rect 263 787 264 788
rect 268 787 269 791
rect 319 791 325 792
rect 319 790 320 791
rect 312 788 320 790
rect 263 786 269 787
rect 302 787 308 788
rect 246 782 252 783
rect 302 783 303 787
rect 307 783 308 787
rect 302 782 308 783
rect 312 778 314 788
rect 319 787 320 788
rect 324 787 325 791
rect 327 791 328 795
rect 332 794 333 795
rect 447 795 453 796
rect 447 794 448 795
rect 332 792 379 794
rect 439 793 448 794
rect 332 791 333 792
rect 327 790 333 791
rect 375 791 381 792
rect 319 786 325 787
rect 358 787 364 788
rect 358 783 359 787
rect 363 783 364 787
rect 375 787 376 791
rect 380 787 381 791
rect 439 789 440 793
rect 444 792 448 793
rect 444 789 445 792
rect 447 791 448 792
rect 452 791 453 795
rect 759 795 765 796
rect 447 790 453 791
rect 503 791 509 792
rect 503 790 504 791
rect 439 788 445 789
rect 496 788 504 790
rect 375 786 381 787
rect 422 787 428 788
rect 358 782 364 783
rect 422 783 423 787
rect 427 783 428 787
rect 422 782 428 783
rect 486 787 492 788
rect 486 783 487 787
rect 491 783 492 787
rect 486 782 492 783
rect 496 778 498 788
rect 503 787 504 788
rect 508 787 509 791
rect 567 791 573 792
rect 503 786 509 787
rect 550 787 556 788
rect 550 783 551 787
rect 555 783 556 787
rect 567 787 568 791
rect 572 790 573 791
rect 598 791 604 792
rect 598 790 599 791
rect 572 788 599 790
rect 572 787 573 788
rect 567 786 573 787
rect 598 787 599 788
rect 603 787 604 791
rect 623 791 629 792
rect 623 790 624 791
rect 616 788 624 790
rect 598 786 604 787
rect 606 787 612 788
rect 550 782 556 783
rect 606 783 607 787
rect 611 783 612 787
rect 606 782 612 783
rect 616 778 618 788
rect 623 787 624 788
rect 628 787 629 791
rect 687 791 693 792
rect 687 790 688 791
rect 680 788 688 790
rect 623 786 629 787
rect 670 787 676 788
rect 670 783 671 787
rect 675 783 676 787
rect 670 782 676 783
rect 680 778 682 788
rect 687 787 688 788
rect 692 787 693 791
rect 750 791 757 792
rect 687 786 693 787
rect 734 787 740 788
rect 734 783 735 787
rect 739 783 740 787
rect 750 787 751 791
rect 756 787 757 791
rect 759 791 760 795
rect 764 794 765 795
rect 1086 795 1087 799
rect 1091 798 1092 799
rect 1119 799 1120 803
rect 1124 802 1125 803
rect 1127 803 1133 804
rect 1127 802 1128 803
rect 1124 800 1128 802
rect 1124 799 1125 800
rect 1119 798 1125 799
rect 1127 799 1128 800
rect 1132 799 1133 803
rect 1152 802 1154 816
rect 1159 815 1160 819
rect 1164 818 1165 819
rect 1199 819 1205 820
rect 1164 816 1178 818
rect 1164 815 1165 816
rect 1159 814 1165 815
rect 1159 803 1165 804
rect 1159 802 1160 803
rect 1152 800 1160 802
rect 1127 798 1133 799
rect 1159 799 1160 800
rect 1164 799 1165 803
rect 1176 802 1178 816
rect 1199 815 1200 819
rect 1204 818 1205 819
rect 1247 819 1253 820
rect 1204 816 1226 818
rect 1204 815 1205 816
rect 1199 814 1205 815
rect 1182 809 1188 810
rect 1182 805 1183 809
rect 1187 805 1188 809
rect 1182 804 1188 805
rect 1199 803 1205 804
rect 1199 802 1200 803
rect 1176 800 1200 802
rect 1159 798 1165 799
rect 1199 799 1200 800
rect 1204 799 1205 803
rect 1224 802 1226 816
rect 1247 815 1248 819
rect 1252 818 1253 819
rect 1295 819 1301 820
rect 1252 816 1290 818
rect 1252 815 1253 816
rect 1247 814 1253 815
rect 1230 809 1236 810
rect 1230 805 1231 809
rect 1235 805 1236 809
rect 1230 804 1236 805
rect 1278 809 1284 810
rect 1278 805 1279 809
rect 1283 805 1284 809
rect 1278 804 1284 805
rect 1247 803 1253 804
rect 1247 802 1248 803
rect 1224 800 1248 802
rect 1199 798 1205 799
rect 1247 799 1248 800
rect 1252 799 1253 803
rect 1288 802 1290 816
rect 1295 815 1296 819
rect 1300 818 1301 819
rect 1336 818 1338 832
rect 1582 825 1588 826
rect 1582 821 1583 825
rect 1587 821 1588 825
rect 1582 820 1588 821
rect 1343 819 1349 820
rect 1343 818 1344 819
rect 1300 816 1322 818
rect 1336 816 1344 818
rect 1300 815 1301 816
rect 1295 814 1301 815
rect 1295 803 1301 804
rect 1295 802 1296 803
rect 1288 800 1296 802
rect 1247 798 1253 799
rect 1295 799 1296 800
rect 1300 799 1301 803
rect 1320 802 1322 816
rect 1343 815 1344 816
rect 1348 815 1349 819
rect 1343 814 1349 815
rect 1326 809 1332 810
rect 1326 805 1327 809
rect 1331 805 1332 809
rect 1326 804 1332 805
rect 1582 808 1588 809
rect 1582 804 1583 808
rect 1587 804 1588 808
rect 1343 803 1349 804
rect 1582 803 1588 804
rect 1343 802 1344 803
rect 1320 800 1344 802
rect 1295 798 1301 799
rect 1343 799 1344 800
rect 1348 799 1349 803
rect 1343 798 1349 799
rect 1091 796 1101 798
rect 1091 795 1092 796
rect 1086 794 1092 795
rect 1099 794 1101 796
rect 764 792 810 794
rect 1099 792 1138 794
rect 764 791 765 792
rect 759 790 765 791
rect 808 790 810 792
rect 815 791 821 792
rect 815 790 816 791
rect 808 788 816 790
rect 750 786 757 787
rect 798 787 804 788
rect 734 782 740 783
rect 798 783 799 787
rect 803 783 804 787
rect 815 787 816 788
rect 820 787 821 791
rect 882 791 893 792
rect 815 786 821 787
rect 870 787 876 788
rect 798 782 804 783
rect 870 783 871 787
rect 875 783 876 787
rect 882 787 883 791
rect 887 787 888 791
rect 892 787 893 791
rect 951 791 957 792
rect 951 790 952 791
rect 944 788 952 790
rect 882 786 893 787
rect 934 787 940 788
rect 870 782 876 783
rect 934 783 935 787
rect 939 783 940 787
rect 934 782 940 783
rect 944 778 946 788
rect 951 787 952 788
rect 956 787 957 791
rect 1015 791 1021 792
rect 1015 790 1016 791
rect 1008 788 1016 790
rect 951 786 957 787
rect 998 787 1004 788
rect 998 783 999 787
rect 1003 783 1004 787
rect 998 782 1004 783
rect 1008 778 1010 788
rect 1015 787 1016 788
rect 1020 787 1021 791
rect 1079 791 1085 792
rect 1015 786 1021 787
rect 1062 787 1068 788
rect 1062 783 1063 787
rect 1067 783 1068 787
rect 1079 787 1080 791
rect 1084 790 1085 791
rect 1136 790 1138 792
rect 1143 791 1149 792
rect 1143 790 1144 791
rect 1084 788 1122 790
rect 1136 788 1144 790
rect 1084 787 1085 788
rect 1079 786 1085 787
rect 1062 782 1068 783
rect 164 776 178 778
rect 196 776 210 778
rect 292 776 314 778
rect 473 776 498 778
rect 596 776 618 778
rect 656 776 682 778
rect 920 776 946 778
rect 984 776 1010 778
rect 1120 778 1122 788
rect 1126 787 1132 788
rect 1126 783 1127 787
rect 1131 783 1132 787
rect 1143 787 1144 788
rect 1148 787 1149 791
rect 1207 791 1213 792
rect 1143 786 1149 787
rect 1190 787 1196 788
rect 1126 782 1132 783
rect 1190 783 1191 787
rect 1195 783 1196 787
rect 1207 787 1208 791
rect 1212 790 1213 791
rect 1246 791 1252 792
rect 1246 790 1247 791
rect 1212 788 1247 790
rect 1212 787 1213 788
rect 1207 786 1213 787
rect 1246 787 1247 788
rect 1251 787 1252 791
rect 1271 791 1277 792
rect 1271 790 1272 791
rect 1264 788 1272 790
rect 1246 786 1252 787
rect 1254 787 1260 788
rect 1190 782 1196 783
rect 1254 783 1255 787
rect 1259 783 1260 787
rect 1254 782 1260 783
rect 1264 778 1266 788
rect 1271 787 1272 788
rect 1276 787 1277 791
rect 1335 791 1341 792
rect 1335 790 1336 791
rect 1328 788 1336 790
rect 1271 786 1277 787
rect 1318 787 1324 788
rect 1318 783 1319 787
rect 1323 783 1324 787
rect 1318 782 1324 783
rect 1328 778 1330 788
rect 1335 787 1336 788
rect 1340 787 1341 791
rect 1399 791 1405 792
rect 1399 790 1400 791
rect 1392 788 1400 790
rect 1335 786 1341 787
rect 1382 787 1388 788
rect 1382 783 1383 787
rect 1387 783 1388 787
rect 1382 782 1388 783
rect 1392 778 1394 788
rect 1399 787 1400 788
rect 1404 787 1405 791
rect 1399 786 1405 787
rect 1582 788 1588 789
rect 1582 784 1583 788
rect 1587 784 1588 788
rect 1582 783 1588 784
rect 1120 776 1138 778
rect 1209 776 1266 778
rect 1304 776 1330 778
rect 1368 776 1394 778
rect 151 775 157 776
rect 110 771 116 772
rect 110 767 111 771
rect 115 767 116 771
rect 151 771 152 775
rect 156 774 157 775
rect 164 774 166 776
rect 156 772 166 774
rect 183 775 189 776
rect 156 771 157 772
rect 151 770 157 771
rect 183 771 184 775
rect 188 774 189 775
rect 196 774 198 776
rect 188 772 198 774
rect 214 775 221 776
rect 188 771 189 772
rect 183 770 189 771
rect 214 771 215 775
rect 220 771 221 775
rect 214 770 221 771
rect 263 775 269 776
rect 263 771 264 775
rect 268 774 269 775
rect 292 774 294 776
rect 268 772 294 774
rect 319 775 325 776
rect 268 771 269 772
rect 263 770 269 771
rect 319 771 320 775
rect 324 774 325 775
rect 327 775 333 776
rect 327 774 328 775
rect 324 772 328 774
rect 324 771 325 772
rect 319 770 325 771
rect 327 771 328 772
rect 332 771 333 775
rect 327 770 333 771
rect 370 775 381 776
rect 370 771 371 775
rect 375 771 376 775
rect 380 771 381 775
rect 370 770 381 771
rect 439 775 445 776
rect 439 771 440 775
rect 444 774 445 775
rect 473 774 475 776
rect 444 772 475 774
rect 503 775 509 776
rect 444 771 445 772
rect 439 770 445 771
rect 503 771 504 775
rect 508 774 509 775
rect 534 775 540 776
rect 534 774 535 775
rect 508 772 535 774
rect 508 771 509 772
rect 503 770 509 771
rect 534 771 535 772
rect 539 771 540 775
rect 534 770 540 771
rect 567 775 573 776
rect 567 771 568 775
rect 572 774 573 775
rect 596 774 598 776
rect 572 772 598 774
rect 623 775 629 776
rect 572 771 573 772
rect 567 770 573 771
rect 623 771 624 775
rect 628 774 629 775
rect 656 774 658 776
rect 628 772 658 774
rect 686 775 693 776
rect 628 771 629 772
rect 623 770 629 771
rect 686 771 687 775
rect 692 771 693 775
rect 686 770 693 771
rect 751 775 757 776
rect 751 771 752 775
rect 756 774 757 775
rect 759 775 765 776
rect 759 774 760 775
rect 756 772 760 774
rect 756 771 757 772
rect 751 770 757 771
rect 759 771 760 772
rect 764 771 765 775
rect 759 770 765 771
rect 810 775 821 776
rect 810 771 811 775
rect 815 771 816 775
rect 820 771 821 775
rect 810 770 821 771
rect 887 775 893 776
rect 887 771 888 775
rect 892 774 893 775
rect 920 774 922 776
rect 892 772 922 774
rect 951 775 957 776
rect 892 771 893 772
rect 887 770 893 771
rect 951 771 952 775
rect 956 774 957 775
rect 984 774 986 776
rect 1015 775 1021 776
rect 1015 774 1016 775
rect 956 772 986 774
rect 1012 772 1016 774
rect 956 771 957 772
rect 951 770 957 771
rect 1010 771 1016 772
rect 1020 771 1021 775
rect 110 766 116 767
rect 134 769 140 770
rect 134 765 135 769
rect 139 765 140 769
rect 134 764 140 765
rect 166 769 172 770
rect 166 765 167 769
rect 171 765 172 769
rect 166 764 172 765
rect 198 769 204 770
rect 198 765 199 769
rect 203 765 204 769
rect 198 764 204 765
rect 246 769 252 770
rect 246 765 247 769
rect 251 765 252 769
rect 246 764 252 765
rect 302 769 308 770
rect 302 765 303 769
rect 307 765 308 769
rect 302 764 308 765
rect 358 769 364 770
rect 358 765 359 769
rect 363 765 364 769
rect 358 764 364 765
rect 422 769 428 770
rect 422 765 423 769
rect 427 765 428 769
rect 422 764 428 765
rect 486 769 492 770
rect 486 765 487 769
rect 491 765 492 769
rect 486 764 492 765
rect 550 769 556 770
rect 550 765 551 769
rect 555 765 556 769
rect 550 764 556 765
rect 606 769 612 770
rect 606 765 607 769
rect 611 765 612 769
rect 606 764 612 765
rect 670 769 676 770
rect 670 765 671 769
rect 675 765 676 769
rect 670 764 676 765
rect 734 769 740 770
rect 734 765 735 769
rect 739 765 740 769
rect 734 764 740 765
rect 798 769 804 770
rect 798 765 799 769
rect 803 765 804 769
rect 798 764 804 765
rect 870 769 876 770
rect 870 765 871 769
rect 875 765 876 769
rect 870 764 876 765
rect 934 769 940 770
rect 934 765 935 769
rect 939 765 940 769
rect 934 764 940 765
rect 998 769 1004 770
rect 998 765 999 769
rect 1003 765 1004 769
rect 1010 767 1011 771
rect 1015 770 1021 771
rect 1078 775 1085 776
rect 1078 771 1079 775
rect 1084 771 1085 775
rect 1136 774 1138 776
rect 1143 775 1149 776
rect 1143 774 1144 775
rect 1136 772 1144 774
rect 1078 770 1085 771
rect 1143 771 1144 772
rect 1148 771 1149 775
rect 1143 770 1149 771
rect 1207 775 1213 776
rect 1207 771 1208 775
rect 1212 771 1213 775
rect 1207 770 1213 771
rect 1271 775 1277 776
rect 1271 771 1272 775
rect 1276 774 1277 775
rect 1304 774 1306 776
rect 1276 772 1306 774
rect 1335 775 1341 776
rect 1276 771 1277 772
rect 1271 770 1277 771
rect 1335 771 1336 775
rect 1340 774 1341 775
rect 1368 774 1370 776
rect 1399 775 1405 776
rect 1399 774 1400 775
rect 1340 772 1370 774
rect 1392 772 1400 774
rect 1340 771 1341 772
rect 1335 770 1341 771
rect 1015 767 1016 770
rect 1010 766 1016 767
rect 1062 769 1068 770
rect 998 764 1004 765
rect 1062 765 1063 769
rect 1067 765 1068 769
rect 1062 764 1068 765
rect 1126 769 1132 770
rect 1126 765 1127 769
rect 1131 765 1132 769
rect 1126 764 1132 765
rect 1190 769 1196 770
rect 1190 765 1191 769
rect 1195 765 1196 769
rect 1190 764 1196 765
rect 1254 769 1260 770
rect 1254 765 1255 769
rect 1259 765 1260 769
rect 1254 764 1260 765
rect 1318 769 1324 770
rect 1318 765 1319 769
rect 1323 765 1324 769
rect 1318 764 1324 765
rect 1382 769 1388 770
rect 1382 765 1383 769
rect 1387 765 1388 769
rect 1382 764 1388 765
rect 1290 763 1296 764
rect 1290 759 1291 763
rect 1295 762 1296 763
rect 1392 762 1394 772
rect 1399 771 1400 772
rect 1404 771 1405 775
rect 1399 770 1405 771
rect 1582 771 1588 772
rect 1582 767 1583 771
rect 1587 767 1588 771
rect 1582 766 1588 767
rect 1295 760 1394 762
rect 1295 759 1296 760
rect 1290 758 1296 759
rect 134 755 140 756
rect 110 753 116 754
rect 110 749 111 753
rect 115 749 116 753
rect 134 751 135 755
rect 139 751 140 755
rect 134 750 140 751
rect 166 755 172 756
rect 166 751 167 755
rect 171 751 172 755
rect 166 750 172 751
rect 198 755 204 756
rect 198 751 199 755
rect 203 751 204 755
rect 198 750 204 751
rect 254 755 260 756
rect 254 751 255 755
rect 259 751 260 755
rect 254 750 260 751
rect 318 755 324 756
rect 318 751 319 755
rect 323 751 324 755
rect 318 750 324 751
rect 390 755 396 756
rect 390 751 391 755
rect 395 751 396 755
rect 390 750 396 751
rect 462 755 468 756
rect 462 751 463 755
rect 467 751 468 755
rect 462 750 468 751
rect 542 755 548 756
rect 542 751 543 755
rect 547 751 548 755
rect 542 750 548 751
rect 622 755 628 756
rect 622 751 623 755
rect 627 751 628 755
rect 622 750 628 751
rect 702 755 708 756
rect 702 751 703 755
rect 707 751 708 755
rect 702 750 708 751
rect 774 755 780 756
rect 774 751 775 755
rect 779 751 780 755
rect 774 750 780 751
rect 846 755 852 756
rect 846 751 847 755
rect 851 751 852 755
rect 846 750 852 751
rect 918 755 924 756
rect 918 751 919 755
rect 923 751 924 755
rect 918 750 924 751
rect 990 755 996 756
rect 990 751 991 755
rect 995 751 996 755
rect 990 750 996 751
rect 1062 755 1068 756
rect 1062 751 1063 755
rect 1067 751 1068 755
rect 1062 750 1068 751
rect 1134 755 1140 756
rect 1134 751 1135 755
rect 1139 751 1140 755
rect 1134 750 1140 751
rect 1206 755 1212 756
rect 1206 751 1207 755
rect 1211 751 1212 755
rect 1206 750 1212 751
rect 1270 755 1276 756
rect 1270 751 1271 755
rect 1275 751 1276 755
rect 1270 750 1276 751
rect 1326 755 1332 756
rect 1326 751 1327 755
rect 1331 751 1332 755
rect 1326 750 1332 751
rect 1374 755 1380 756
rect 1374 751 1375 755
rect 1379 751 1380 755
rect 1374 750 1380 751
rect 1422 755 1428 756
rect 1422 751 1423 755
rect 1427 751 1428 755
rect 1422 750 1428 751
rect 1470 755 1476 756
rect 1470 751 1471 755
rect 1475 751 1476 755
rect 1470 750 1476 751
rect 1510 755 1516 756
rect 1510 751 1511 755
rect 1515 751 1516 755
rect 1510 750 1516 751
rect 1542 755 1548 756
rect 1542 751 1543 755
rect 1547 751 1548 755
rect 1542 750 1548 751
rect 1582 753 1588 754
rect 110 748 116 749
rect 1582 749 1583 753
rect 1587 749 1588 753
rect 1582 748 1588 749
rect 150 747 157 748
rect 150 743 151 747
rect 156 743 157 747
rect 183 747 189 748
rect 183 746 184 747
rect 150 742 157 743
rect 176 744 184 746
rect 134 737 140 738
rect 110 736 116 737
rect 110 732 111 736
rect 115 732 116 736
rect 134 733 135 737
rect 139 733 140 737
rect 134 732 140 733
rect 166 737 172 738
rect 166 733 167 737
rect 171 733 172 737
rect 166 732 172 733
rect 110 731 116 732
rect 151 731 157 732
rect 151 727 152 731
rect 156 730 157 731
rect 176 730 178 744
rect 183 743 184 744
rect 188 743 189 747
rect 183 742 189 743
rect 215 747 221 748
rect 215 743 216 747
rect 220 746 221 747
rect 223 747 229 748
rect 223 746 224 747
rect 220 744 224 746
rect 220 743 221 744
rect 215 742 221 743
rect 223 743 224 744
rect 228 743 229 747
rect 271 747 277 748
rect 271 746 272 747
rect 223 742 229 743
rect 240 744 272 746
rect 214 739 220 740
rect 214 738 215 739
rect 198 737 204 738
rect 198 733 199 737
rect 203 733 204 737
rect 198 732 204 733
rect 208 736 215 738
rect 156 728 178 730
rect 183 731 189 732
rect 156 727 157 728
rect 151 726 157 727
rect 183 727 184 731
rect 188 730 189 731
rect 208 730 210 736
rect 214 735 215 736
rect 219 735 220 739
rect 214 734 220 735
rect 188 728 210 730
rect 215 731 221 732
rect 188 727 189 728
rect 183 726 189 727
rect 215 727 216 731
rect 220 730 221 731
rect 240 730 242 744
rect 271 743 272 744
rect 276 743 277 747
rect 335 747 341 748
rect 335 746 336 747
rect 271 742 277 743
rect 308 744 336 746
rect 254 737 260 738
rect 254 733 255 737
rect 259 733 260 737
rect 254 732 260 733
rect 220 728 242 730
rect 271 731 277 732
rect 220 727 221 728
rect 215 726 221 727
rect 271 727 272 731
rect 276 730 277 731
rect 308 730 310 744
rect 335 743 336 744
rect 340 743 341 747
rect 407 747 413 748
rect 407 746 408 747
rect 335 742 341 743
rect 376 744 408 746
rect 318 737 324 738
rect 318 733 319 737
rect 323 733 324 737
rect 318 732 324 733
rect 276 728 310 730
rect 335 731 341 732
rect 276 727 277 728
rect 271 726 277 727
rect 335 727 336 731
rect 340 730 341 731
rect 376 730 378 744
rect 407 743 408 744
rect 412 743 413 747
rect 407 742 413 743
rect 479 747 485 748
rect 479 743 480 747
rect 484 746 485 747
rect 502 747 508 748
rect 502 746 503 747
rect 484 744 503 746
rect 484 743 485 744
rect 479 742 485 743
rect 502 743 503 744
rect 507 743 508 747
rect 502 742 508 743
rect 558 747 565 748
rect 558 743 559 747
rect 564 743 565 747
rect 558 742 565 743
rect 598 747 604 748
rect 598 743 599 747
rect 603 746 604 747
rect 639 747 645 748
rect 639 746 640 747
rect 603 744 640 746
rect 603 743 604 744
rect 598 742 604 743
rect 639 743 640 744
rect 644 743 645 747
rect 639 742 645 743
rect 719 747 725 748
rect 719 743 720 747
rect 724 746 725 747
rect 766 747 772 748
rect 766 746 767 747
rect 724 744 767 746
rect 724 743 725 744
rect 719 742 725 743
rect 766 743 767 744
rect 771 743 772 747
rect 791 747 797 748
rect 791 746 792 747
rect 766 742 772 743
rect 784 744 792 746
rect 390 737 396 738
rect 390 733 391 737
rect 395 733 396 737
rect 390 732 396 733
rect 462 737 468 738
rect 462 733 463 737
rect 467 733 468 737
rect 462 732 468 733
rect 542 737 548 738
rect 542 733 543 737
rect 547 733 548 737
rect 542 732 548 733
rect 622 737 628 738
rect 622 733 623 737
rect 627 733 628 737
rect 622 732 628 733
rect 702 737 708 738
rect 702 733 703 737
rect 707 733 708 737
rect 702 732 708 733
rect 774 737 780 738
rect 774 733 775 737
rect 779 733 780 737
rect 774 732 780 733
rect 340 728 378 730
rect 398 731 404 732
rect 340 727 341 728
rect 335 726 341 727
rect 398 727 399 731
rect 403 730 404 731
rect 407 731 413 732
rect 407 730 408 731
rect 403 728 408 730
rect 403 727 404 728
rect 398 726 404 727
rect 407 727 408 728
rect 412 727 413 731
rect 407 726 413 727
rect 442 731 448 732
rect 442 727 443 731
rect 447 730 448 731
rect 479 731 485 732
rect 479 730 480 731
rect 447 728 480 730
rect 447 727 448 728
rect 442 726 448 727
rect 479 727 480 728
rect 484 727 485 731
rect 479 726 485 727
rect 534 731 540 732
rect 534 727 535 731
rect 539 730 540 731
rect 559 731 565 732
rect 559 730 560 731
rect 539 728 560 730
rect 539 727 540 728
rect 534 726 540 727
rect 559 727 560 728
rect 564 727 565 731
rect 559 726 565 727
rect 634 731 645 732
rect 634 727 635 731
rect 639 727 640 731
rect 644 727 645 731
rect 634 726 645 727
rect 719 731 725 732
rect 719 727 720 731
rect 724 730 725 731
rect 784 730 786 744
rect 791 743 792 744
rect 796 743 797 747
rect 791 742 797 743
rect 863 747 869 748
rect 863 743 864 747
rect 868 746 869 747
rect 882 747 888 748
rect 882 746 883 747
rect 868 744 883 746
rect 868 743 869 744
rect 863 742 869 743
rect 882 743 883 744
rect 887 743 888 747
rect 935 747 941 748
rect 935 746 936 747
rect 882 742 888 743
rect 900 744 936 746
rect 846 737 852 738
rect 846 733 847 737
rect 851 733 852 737
rect 846 732 852 733
rect 724 728 786 730
rect 791 731 797 732
rect 724 727 725 728
rect 719 726 725 727
rect 791 727 792 731
rect 796 730 797 731
rect 810 731 816 732
rect 810 730 811 731
rect 796 728 811 730
rect 796 727 797 728
rect 791 726 797 727
rect 810 727 811 728
rect 815 727 816 731
rect 810 726 816 727
rect 863 731 869 732
rect 863 727 864 731
rect 868 730 869 731
rect 900 730 902 744
rect 935 743 936 744
rect 940 743 941 747
rect 1007 747 1013 748
rect 1007 746 1008 747
rect 935 742 941 743
rect 972 744 1008 746
rect 918 737 924 738
rect 918 733 919 737
rect 923 733 924 737
rect 918 732 924 733
rect 868 728 902 730
rect 935 731 941 732
rect 868 727 869 728
rect 863 726 869 727
rect 935 727 936 731
rect 940 730 941 731
rect 972 730 974 744
rect 1007 743 1008 744
rect 1012 743 1013 747
rect 1007 742 1013 743
rect 1079 747 1085 748
rect 1079 743 1080 747
rect 1084 746 1085 747
rect 1151 747 1157 748
rect 1084 744 1118 746
rect 1084 743 1085 744
rect 1079 742 1085 743
rect 990 737 996 738
rect 990 733 991 737
rect 995 733 996 737
rect 990 732 996 733
rect 1062 737 1068 738
rect 1062 733 1063 737
rect 1067 733 1068 737
rect 1062 732 1068 733
rect 940 728 974 730
rect 1007 731 1013 732
rect 940 727 941 728
rect 935 726 941 727
rect 1007 727 1008 731
rect 1012 730 1013 731
rect 1022 731 1028 732
rect 1022 730 1023 731
rect 1012 728 1023 730
rect 1012 727 1013 728
rect 1007 726 1013 727
rect 1022 727 1023 728
rect 1027 727 1028 731
rect 1022 726 1028 727
rect 1078 731 1085 732
rect 1078 727 1079 731
rect 1084 727 1085 731
rect 1116 730 1118 744
rect 1151 743 1152 747
rect 1156 743 1157 747
rect 1151 742 1157 743
rect 1186 747 1192 748
rect 1186 743 1187 747
rect 1191 746 1192 747
rect 1223 747 1229 748
rect 1223 746 1224 747
rect 1191 744 1224 746
rect 1191 743 1192 744
rect 1186 742 1192 743
rect 1223 743 1224 744
rect 1228 743 1229 747
rect 1223 742 1229 743
rect 1287 747 1293 748
rect 1287 743 1288 747
rect 1292 746 1293 747
rect 1343 747 1349 748
rect 1292 744 1318 746
rect 1292 743 1293 744
rect 1287 742 1293 743
rect 1153 738 1155 742
rect 1134 737 1140 738
rect 1134 733 1135 737
rect 1139 733 1140 737
rect 1153 736 1190 738
rect 1134 732 1140 733
rect 1151 731 1157 732
rect 1151 730 1152 731
rect 1116 728 1152 730
rect 1078 726 1085 727
rect 1151 727 1152 728
rect 1156 727 1157 731
rect 1188 730 1190 736
rect 1206 737 1212 738
rect 1206 733 1207 737
rect 1211 733 1212 737
rect 1206 732 1212 733
rect 1270 737 1276 738
rect 1270 733 1271 737
rect 1275 733 1276 737
rect 1270 732 1276 733
rect 1223 731 1229 732
rect 1223 730 1224 731
rect 1188 728 1224 730
rect 1151 726 1157 727
rect 1223 727 1224 728
rect 1228 727 1229 731
rect 1223 726 1229 727
rect 1287 731 1296 732
rect 1287 727 1288 731
rect 1295 727 1296 731
rect 1316 730 1318 744
rect 1343 743 1344 747
rect 1348 746 1349 747
rect 1391 747 1397 748
rect 1348 744 1370 746
rect 1348 743 1349 744
rect 1343 742 1349 743
rect 1326 737 1332 738
rect 1326 733 1327 737
rect 1331 733 1332 737
rect 1326 732 1332 733
rect 1343 731 1349 732
rect 1343 730 1344 731
rect 1316 728 1344 730
rect 1287 726 1296 727
rect 1343 727 1344 728
rect 1348 727 1349 731
rect 1368 730 1370 744
rect 1391 743 1392 747
rect 1396 746 1397 747
rect 1439 747 1445 748
rect 1396 744 1418 746
rect 1396 743 1397 744
rect 1391 742 1397 743
rect 1374 737 1380 738
rect 1374 733 1375 737
rect 1379 733 1380 737
rect 1374 732 1380 733
rect 1391 731 1397 732
rect 1391 730 1392 731
rect 1368 728 1392 730
rect 1343 726 1349 727
rect 1391 727 1392 728
rect 1396 727 1397 731
rect 1416 730 1418 744
rect 1439 743 1440 747
rect 1444 746 1445 747
rect 1487 747 1493 748
rect 1444 744 1461 746
rect 1444 743 1445 744
rect 1439 742 1445 743
rect 1422 737 1428 738
rect 1422 733 1423 737
rect 1427 733 1428 737
rect 1422 732 1428 733
rect 1439 731 1445 732
rect 1439 730 1440 731
rect 1416 728 1440 730
rect 1391 726 1397 727
rect 1439 727 1440 728
rect 1444 727 1445 731
rect 1459 730 1461 744
rect 1487 743 1488 747
rect 1492 746 1493 747
rect 1527 747 1533 748
rect 1492 744 1506 746
rect 1492 743 1493 744
rect 1487 742 1493 743
rect 1470 737 1476 738
rect 1470 733 1471 737
rect 1475 733 1476 737
rect 1470 732 1476 733
rect 1487 731 1493 732
rect 1487 730 1488 731
rect 1459 728 1488 730
rect 1439 726 1445 727
rect 1487 727 1488 728
rect 1492 727 1493 731
rect 1504 730 1506 744
rect 1527 743 1528 747
rect 1532 746 1533 747
rect 1558 747 1565 748
rect 1532 744 1554 746
rect 1532 743 1533 744
rect 1527 742 1533 743
rect 1510 737 1516 738
rect 1510 733 1511 737
rect 1515 733 1516 737
rect 1510 732 1516 733
rect 1542 737 1548 738
rect 1542 733 1543 737
rect 1547 733 1548 737
rect 1542 732 1548 733
rect 1527 731 1533 732
rect 1527 730 1528 731
rect 1504 728 1528 730
rect 1487 726 1493 727
rect 1527 727 1528 728
rect 1532 727 1533 731
rect 1552 730 1554 744
rect 1558 743 1559 747
rect 1564 743 1565 747
rect 1558 742 1565 743
rect 1582 736 1588 737
rect 1582 732 1583 736
rect 1587 732 1588 736
rect 1559 731 1565 732
rect 1582 731 1588 732
rect 1559 730 1560 731
rect 1552 728 1560 730
rect 1527 726 1533 727
rect 1559 727 1560 728
rect 1564 727 1565 731
rect 1559 726 1565 727
rect 658 723 664 724
rect 537 720 554 722
rect 150 719 157 720
rect 110 716 116 717
rect 110 712 111 716
rect 115 712 116 716
rect 110 711 116 712
rect 134 715 140 716
rect 134 711 135 715
rect 139 711 140 715
rect 150 715 151 719
rect 156 715 157 719
rect 183 719 189 720
rect 183 718 184 719
rect 176 716 184 718
rect 150 714 157 715
rect 166 715 172 716
rect 134 710 140 711
rect 166 711 167 715
rect 171 711 172 715
rect 166 710 172 711
rect 176 706 178 716
rect 183 715 184 716
rect 188 715 189 719
rect 223 719 229 720
rect 223 718 224 719
rect 216 716 224 718
rect 183 714 189 715
rect 206 715 212 716
rect 206 711 207 715
rect 211 711 212 715
rect 206 710 212 711
rect 216 706 218 716
rect 223 715 224 716
rect 228 715 229 719
rect 270 719 277 720
rect 223 714 229 715
rect 254 715 260 716
rect 254 711 255 715
rect 259 711 260 715
rect 270 715 271 719
rect 276 715 277 719
rect 327 719 333 720
rect 327 718 328 719
rect 320 716 328 718
rect 270 714 277 715
rect 310 715 316 716
rect 254 710 260 711
rect 310 711 311 715
rect 315 711 316 715
rect 310 710 316 711
rect 320 706 322 716
rect 327 715 328 716
rect 332 715 333 719
rect 383 719 389 720
rect 383 718 384 719
rect 376 716 384 718
rect 327 714 333 715
rect 366 715 372 716
rect 366 711 367 715
rect 371 711 372 715
rect 366 710 372 711
rect 376 706 378 716
rect 383 715 384 716
rect 388 715 389 719
rect 434 719 445 720
rect 383 714 389 715
rect 422 715 428 716
rect 422 711 423 715
rect 427 711 428 715
rect 434 715 435 719
rect 439 715 440 719
rect 444 715 445 719
rect 495 719 501 720
rect 434 714 445 715
rect 478 715 484 716
rect 422 710 428 711
rect 478 711 479 715
rect 483 711 484 715
rect 495 715 496 719
rect 500 718 501 719
rect 537 718 539 720
rect 500 716 539 718
rect 500 715 501 716
rect 495 714 501 715
rect 542 715 548 716
rect 478 710 484 711
rect 542 711 543 715
rect 547 711 548 715
rect 542 710 548 711
rect 164 704 178 706
rect 204 704 218 706
rect 273 704 322 706
rect 356 704 378 706
rect 151 703 157 704
rect 110 699 116 700
rect 110 695 111 699
rect 115 695 116 699
rect 151 699 152 703
rect 156 702 157 703
rect 164 702 166 704
rect 156 700 166 702
rect 183 703 189 704
rect 156 699 157 700
rect 151 698 157 699
rect 183 699 184 703
rect 188 702 189 703
rect 204 702 206 704
rect 188 700 206 702
rect 222 703 229 704
rect 188 699 189 700
rect 183 698 189 699
rect 222 699 223 703
rect 228 699 229 703
rect 222 698 229 699
rect 271 703 277 704
rect 271 699 272 703
rect 276 699 277 703
rect 271 698 277 699
rect 327 703 333 704
rect 327 699 328 703
rect 332 702 333 703
rect 356 702 358 704
rect 332 700 358 702
rect 383 703 389 704
rect 332 699 333 700
rect 327 698 333 699
rect 383 699 384 703
rect 388 702 389 703
rect 398 703 404 704
rect 398 702 399 703
rect 388 700 399 702
rect 388 699 389 700
rect 383 698 389 699
rect 398 699 399 700
rect 403 699 404 703
rect 398 698 404 699
rect 439 703 448 704
rect 439 699 440 703
rect 447 699 448 703
rect 439 698 448 699
rect 495 703 501 704
rect 495 699 496 703
rect 500 702 501 703
rect 534 703 540 704
rect 534 702 535 703
rect 500 700 535 702
rect 500 699 501 700
rect 495 698 501 699
rect 534 699 535 700
rect 539 699 540 703
rect 552 702 554 720
rect 558 719 565 720
rect 558 715 559 719
rect 564 715 565 719
rect 631 719 637 720
rect 558 714 565 715
rect 614 715 620 716
rect 614 711 615 715
rect 619 711 620 715
rect 631 715 632 719
rect 636 718 637 719
rect 658 719 659 723
rect 663 722 664 723
rect 766 723 772 724
rect 663 720 698 722
rect 663 719 664 720
rect 658 718 664 719
rect 696 718 698 720
rect 703 719 709 720
rect 703 718 704 719
rect 636 716 654 718
rect 696 716 704 718
rect 636 715 637 716
rect 631 714 637 715
rect 614 710 620 711
rect 652 706 654 716
rect 686 715 692 716
rect 686 711 687 715
rect 691 711 692 715
rect 703 715 704 716
rect 708 715 709 719
rect 766 719 767 723
rect 771 719 772 723
rect 766 718 772 719
rect 775 719 781 720
rect 775 718 776 719
rect 768 716 776 718
rect 703 714 709 715
rect 758 715 764 716
rect 686 710 692 711
rect 758 711 759 715
rect 763 711 764 715
rect 775 715 776 716
rect 780 715 781 719
rect 854 719 861 720
rect 775 714 781 715
rect 838 715 844 716
rect 758 710 764 711
rect 838 711 839 715
rect 843 711 844 715
rect 854 715 855 719
rect 860 715 861 719
rect 935 719 941 720
rect 935 718 936 719
rect 928 716 936 718
rect 854 714 861 715
rect 918 715 924 716
rect 838 710 844 711
rect 918 711 919 715
rect 923 711 924 715
rect 918 710 924 711
rect 714 707 720 708
rect 652 704 698 706
rect 559 703 565 704
rect 559 702 560 703
rect 552 700 560 702
rect 534 698 540 699
rect 559 699 560 700
rect 564 699 565 703
rect 559 698 565 699
rect 631 703 640 704
rect 631 699 632 703
rect 639 699 640 703
rect 696 702 698 704
rect 703 703 709 704
rect 703 702 704 703
rect 696 700 704 702
rect 631 698 640 699
rect 703 699 704 700
rect 708 699 709 703
rect 714 703 715 707
rect 719 706 720 707
rect 928 706 930 716
rect 935 715 936 716
rect 940 715 941 719
rect 1023 719 1029 720
rect 1023 718 1024 719
rect 1016 716 1024 718
rect 935 714 941 715
rect 1006 715 1012 716
rect 1006 711 1007 715
rect 1011 711 1012 715
rect 1006 710 1012 711
rect 1016 706 1018 716
rect 1023 715 1024 716
rect 1028 715 1029 719
rect 1103 719 1109 720
rect 1023 714 1029 715
rect 1086 715 1092 716
rect 1086 711 1087 715
rect 1091 711 1092 715
rect 1103 715 1104 719
rect 1108 718 1109 719
rect 1183 719 1192 720
rect 1108 716 1150 718
rect 1108 715 1109 716
rect 1103 714 1109 715
rect 1086 710 1092 711
rect 719 704 770 706
rect 897 704 930 706
rect 937 704 1018 706
rect 1034 707 1040 708
rect 719 703 720 704
rect 714 702 720 703
rect 768 702 770 704
rect 775 703 781 704
rect 775 702 776 703
rect 768 700 776 702
rect 703 698 709 699
rect 775 699 776 700
rect 780 699 781 703
rect 775 698 781 699
rect 855 703 861 704
rect 855 699 856 703
rect 860 702 861 703
rect 897 702 899 704
rect 860 700 899 702
rect 935 703 941 704
rect 860 699 861 700
rect 855 698 861 699
rect 935 699 936 703
rect 940 699 941 703
rect 935 698 941 699
rect 1022 703 1029 704
rect 1022 699 1023 703
rect 1028 699 1029 703
rect 1034 703 1035 707
rect 1039 706 1040 707
rect 1148 706 1150 716
rect 1166 715 1172 716
rect 1166 711 1167 715
rect 1171 711 1172 715
rect 1183 715 1184 719
rect 1191 715 1192 719
rect 1255 719 1261 720
rect 1183 714 1192 715
rect 1238 715 1244 716
rect 1166 710 1172 711
rect 1238 711 1239 715
rect 1243 711 1244 715
rect 1255 715 1256 719
rect 1260 718 1261 719
rect 1294 719 1300 720
rect 1294 718 1295 719
rect 1260 716 1295 718
rect 1260 715 1261 716
rect 1255 714 1261 715
rect 1294 715 1295 716
rect 1299 715 1300 719
rect 1319 719 1325 720
rect 1319 718 1320 719
rect 1312 716 1320 718
rect 1294 714 1300 715
rect 1302 715 1308 716
rect 1238 710 1244 711
rect 1302 711 1303 715
rect 1307 711 1308 715
rect 1302 710 1308 711
rect 1312 706 1314 716
rect 1319 715 1320 716
rect 1324 715 1325 719
rect 1375 719 1381 720
rect 1319 714 1325 715
rect 1358 715 1364 716
rect 1358 711 1359 715
rect 1363 711 1364 715
rect 1375 715 1376 719
rect 1380 715 1381 719
rect 1423 719 1429 720
rect 1375 714 1381 715
rect 1406 715 1412 716
rect 1358 710 1364 711
rect 1377 710 1379 714
rect 1406 711 1407 715
rect 1411 711 1412 715
rect 1423 715 1424 719
rect 1428 718 1429 719
rect 1471 719 1477 720
rect 1428 716 1443 718
rect 1428 715 1429 716
rect 1423 714 1429 715
rect 1406 710 1412 711
rect 1377 708 1402 710
rect 1039 704 1101 706
rect 1148 704 1187 706
rect 1288 704 1314 706
rect 1400 706 1402 708
rect 1441 706 1443 716
rect 1454 715 1460 716
rect 1454 711 1455 715
rect 1459 711 1460 715
rect 1471 715 1472 719
rect 1476 718 1477 719
rect 1527 719 1533 720
rect 1476 716 1506 718
rect 1476 715 1477 716
rect 1471 714 1477 715
rect 1454 710 1460 711
rect 1464 708 1474 710
rect 1464 706 1466 708
rect 1472 706 1474 708
rect 1504 706 1506 716
rect 1510 715 1516 716
rect 1510 711 1511 715
rect 1515 711 1516 715
rect 1527 715 1528 719
rect 1532 718 1533 719
rect 1558 719 1565 720
rect 1532 716 1538 718
rect 1532 715 1533 716
rect 1527 714 1533 715
rect 1510 710 1516 711
rect 1536 706 1538 716
rect 1542 715 1548 716
rect 1542 711 1543 715
rect 1547 711 1548 715
rect 1558 715 1559 719
rect 1564 715 1565 719
rect 1558 714 1565 715
rect 1582 716 1588 717
rect 1582 712 1583 716
rect 1587 712 1588 716
rect 1582 711 1588 712
rect 1542 710 1548 711
rect 1400 704 1418 706
rect 1441 704 1466 706
rect 1471 705 1477 706
rect 1039 703 1040 704
rect 1034 702 1040 703
rect 1099 702 1101 704
rect 1103 703 1109 704
rect 1103 702 1104 703
rect 1099 700 1104 702
rect 1022 698 1029 699
rect 1103 699 1104 700
rect 1108 699 1109 703
rect 1103 698 1109 699
rect 1183 703 1189 704
rect 1183 699 1184 703
rect 1188 699 1189 703
rect 1183 698 1189 699
rect 1255 703 1261 704
rect 1255 699 1256 703
rect 1260 702 1261 703
rect 1288 702 1290 704
rect 1260 700 1290 702
rect 1319 703 1325 704
rect 1260 699 1261 700
rect 1255 698 1261 699
rect 1319 699 1320 703
rect 1324 702 1325 703
rect 1350 703 1356 704
rect 1350 702 1351 703
rect 1324 700 1351 702
rect 1324 699 1325 700
rect 1319 698 1325 699
rect 1350 699 1351 700
rect 1355 699 1356 703
rect 1350 698 1356 699
rect 1375 703 1381 704
rect 1375 699 1376 703
rect 1380 699 1381 703
rect 1416 702 1418 704
rect 1423 703 1429 704
rect 1423 702 1424 703
rect 1416 700 1424 702
rect 1375 698 1381 699
rect 1423 699 1424 700
rect 1428 699 1429 703
rect 1471 701 1472 705
rect 1476 701 1477 705
rect 1504 704 1522 706
rect 1536 704 1563 706
rect 1471 700 1477 701
rect 1520 702 1522 704
rect 1527 703 1533 704
rect 1527 702 1528 703
rect 1520 700 1528 702
rect 1423 698 1429 699
rect 1527 699 1528 700
rect 1532 699 1533 703
rect 1527 698 1533 699
rect 1559 703 1565 704
rect 1559 699 1560 703
rect 1564 699 1565 703
rect 1559 698 1565 699
rect 1582 699 1588 700
rect 110 694 116 695
rect 134 697 140 698
rect 134 693 135 697
rect 139 693 140 697
rect 134 692 140 693
rect 166 697 172 698
rect 166 693 167 697
rect 171 693 172 697
rect 166 692 172 693
rect 206 697 212 698
rect 206 693 207 697
rect 211 693 212 697
rect 206 692 212 693
rect 254 697 260 698
rect 254 693 255 697
rect 259 693 260 697
rect 254 692 260 693
rect 310 697 316 698
rect 310 693 311 697
rect 315 693 316 697
rect 310 692 316 693
rect 366 697 372 698
rect 366 693 367 697
rect 371 693 372 697
rect 366 692 372 693
rect 422 697 428 698
rect 422 693 423 697
rect 427 693 428 697
rect 422 692 428 693
rect 478 697 484 698
rect 478 693 479 697
rect 483 693 484 697
rect 478 692 484 693
rect 542 697 548 698
rect 542 693 543 697
rect 547 693 548 697
rect 542 692 548 693
rect 614 697 620 698
rect 614 693 615 697
rect 619 693 620 697
rect 614 692 620 693
rect 686 697 692 698
rect 686 693 687 697
rect 691 693 692 697
rect 686 692 692 693
rect 758 697 764 698
rect 758 693 759 697
rect 763 693 764 697
rect 758 692 764 693
rect 838 697 844 698
rect 838 693 839 697
rect 843 693 844 697
rect 838 692 844 693
rect 918 697 924 698
rect 918 693 919 697
rect 923 693 924 697
rect 918 692 924 693
rect 1006 697 1012 698
rect 1006 693 1007 697
rect 1011 693 1012 697
rect 1006 692 1012 693
rect 1086 697 1092 698
rect 1086 693 1087 697
rect 1091 693 1092 697
rect 1086 692 1092 693
rect 1166 697 1172 698
rect 1166 693 1167 697
rect 1171 693 1172 697
rect 1166 692 1172 693
rect 1238 697 1244 698
rect 1238 693 1239 697
rect 1243 693 1244 697
rect 1238 692 1244 693
rect 1302 697 1308 698
rect 1302 693 1303 697
rect 1307 693 1308 697
rect 1302 692 1308 693
rect 1358 697 1364 698
rect 1358 693 1359 697
rect 1363 693 1364 697
rect 1358 692 1364 693
rect 1294 691 1300 692
rect 1294 687 1295 691
rect 1299 690 1300 691
rect 1377 690 1379 698
rect 1406 697 1412 698
rect 1406 693 1407 697
rect 1411 693 1412 697
rect 1406 692 1412 693
rect 1454 697 1460 698
rect 1454 693 1455 697
rect 1459 693 1460 697
rect 1454 692 1460 693
rect 1510 697 1516 698
rect 1510 693 1511 697
rect 1515 693 1516 697
rect 1510 692 1516 693
rect 1542 697 1548 698
rect 1542 693 1543 697
rect 1547 693 1548 697
rect 1582 695 1583 699
rect 1587 695 1588 699
rect 1582 694 1588 695
rect 1542 692 1548 693
rect 1299 688 1379 690
rect 1299 687 1300 688
rect 1294 686 1300 687
rect 158 683 164 684
rect 110 681 116 682
rect 110 677 111 681
rect 115 677 116 681
rect 158 679 159 683
rect 163 679 164 683
rect 158 678 164 679
rect 206 683 212 684
rect 206 679 207 683
rect 211 679 212 683
rect 206 678 212 679
rect 254 683 260 684
rect 254 679 255 683
rect 259 679 260 683
rect 254 678 260 679
rect 302 683 308 684
rect 302 679 303 683
rect 307 679 308 683
rect 302 678 308 679
rect 358 683 364 684
rect 358 679 359 683
rect 363 679 364 683
rect 358 678 364 679
rect 414 683 420 684
rect 414 679 415 683
rect 419 679 420 683
rect 414 678 420 679
rect 470 683 476 684
rect 470 679 471 683
rect 475 679 476 683
rect 470 678 476 679
rect 526 683 532 684
rect 526 679 527 683
rect 531 679 532 683
rect 526 678 532 679
rect 582 683 588 684
rect 582 679 583 683
rect 587 679 588 683
rect 582 678 588 679
rect 638 683 644 684
rect 638 679 639 683
rect 643 679 644 683
rect 638 678 644 679
rect 694 683 700 684
rect 694 679 695 683
rect 699 679 700 683
rect 694 678 700 679
rect 758 683 764 684
rect 758 679 759 683
rect 763 679 764 683
rect 758 678 764 679
rect 822 683 828 684
rect 822 679 823 683
rect 827 679 828 683
rect 822 678 828 679
rect 886 683 892 684
rect 886 679 887 683
rect 891 679 892 683
rect 886 678 892 679
rect 950 683 956 684
rect 950 679 951 683
rect 955 679 956 683
rect 950 678 956 679
rect 1014 683 1020 684
rect 1014 679 1015 683
rect 1019 679 1020 683
rect 1014 678 1020 679
rect 1078 683 1084 684
rect 1078 679 1079 683
rect 1083 679 1084 683
rect 1078 678 1084 679
rect 1134 683 1140 684
rect 1134 679 1135 683
rect 1139 679 1140 683
rect 1134 678 1140 679
rect 1190 683 1196 684
rect 1190 679 1191 683
rect 1195 679 1196 683
rect 1190 678 1196 679
rect 1246 683 1252 684
rect 1246 679 1247 683
rect 1251 679 1252 683
rect 1246 678 1252 679
rect 1302 683 1308 684
rect 1302 679 1303 683
rect 1307 679 1308 683
rect 1302 678 1308 679
rect 1358 683 1364 684
rect 1358 679 1359 683
rect 1363 679 1364 683
rect 1358 678 1364 679
rect 1582 681 1588 682
rect 110 676 116 677
rect 1582 677 1583 681
rect 1587 677 1588 681
rect 1582 676 1588 677
rect 175 675 184 676
rect 175 671 176 675
rect 183 671 184 675
rect 223 675 229 676
rect 223 674 224 675
rect 175 670 184 671
rect 200 672 224 674
rect 158 665 164 666
rect 110 664 116 665
rect 110 660 111 664
rect 115 660 116 664
rect 158 661 159 665
rect 163 661 164 665
rect 158 660 164 661
rect 110 659 116 660
rect 175 659 181 660
rect 175 655 176 659
rect 180 658 181 659
rect 200 658 202 672
rect 223 671 224 672
rect 228 671 229 675
rect 223 670 229 671
rect 270 675 277 676
rect 270 671 271 675
rect 276 671 277 675
rect 319 675 325 676
rect 319 674 320 675
rect 270 670 277 671
rect 296 672 320 674
rect 206 665 212 666
rect 206 661 207 665
rect 211 661 212 665
rect 206 660 212 661
rect 254 665 260 666
rect 254 661 255 665
rect 259 661 260 665
rect 254 660 260 661
rect 180 656 202 658
rect 222 659 229 660
rect 180 655 181 656
rect 175 654 181 655
rect 222 655 223 659
rect 228 655 229 659
rect 222 654 229 655
rect 271 659 277 660
rect 271 655 272 659
rect 276 658 277 659
rect 296 658 298 672
rect 319 671 320 672
rect 324 671 325 675
rect 375 675 381 676
rect 375 674 376 675
rect 319 670 325 671
rect 352 672 376 674
rect 302 665 308 666
rect 302 661 303 665
rect 307 661 308 665
rect 302 660 308 661
rect 276 656 298 658
rect 319 659 325 660
rect 276 655 277 656
rect 271 654 277 655
rect 319 655 320 659
rect 324 658 325 659
rect 352 658 354 672
rect 375 671 376 672
rect 380 671 381 675
rect 375 670 381 671
rect 431 675 440 676
rect 431 671 432 675
rect 439 671 440 675
rect 431 670 440 671
rect 442 675 448 676
rect 442 671 443 675
rect 447 674 448 675
rect 487 675 493 676
rect 487 674 488 675
rect 447 672 488 674
rect 447 671 448 672
rect 442 670 448 671
rect 487 671 488 672
rect 492 671 493 675
rect 487 670 493 671
rect 506 675 512 676
rect 506 671 507 675
rect 511 674 512 675
rect 543 675 549 676
rect 543 674 544 675
rect 511 672 544 674
rect 511 671 512 672
rect 506 670 512 671
rect 543 671 544 672
rect 548 671 549 675
rect 543 670 549 671
rect 599 675 605 676
rect 599 671 600 675
rect 604 674 605 675
rect 655 675 664 676
rect 604 672 630 674
rect 604 671 605 672
rect 599 670 605 671
rect 358 665 364 666
rect 358 661 359 665
rect 363 661 364 665
rect 358 660 364 661
rect 414 665 420 666
rect 414 661 415 665
rect 419 661 420 665
rect 414 660 420 661
rect 470 665 476 666
rect 470 661 471 665
rect 475 661 476 665
rect 470 660 476 661
rect 526 665 532 666
rect 526 661 527 665
rect 531 661 532 665
rect 526 660 532 661
rect 582 665 588 666
rect 582 661 583 665
rect 587 661 588 665
rect 582 660 588 661
rect 324 656 354 658
rect 375 659 381 660
rect 324 655 325 656
rect 319 654 325 655
rect 375 655 376 659
rect 380 655 381 659
rect 375 654 381 655
rect 402 659 408 660
rect 402 655 403 659
rect 407 658 408 659
rect 431 659 437 660
rect 431 658 432 659
rect 407 656 432 658
rect 407 655 408 656
rect 402 654 408 655
rect 431 655 432 656
rect 436 655 437 659
rect 431 654 437 655
rect 450 659 456 660
rect 450 655 451 659
rect 455 658 456 659
rect 487 659 493 660
rect 487 658 488 659
rect 455 656 488 658
rect 455 655 456 656
rect 450 654 456 655
rect 487 655 488 656
rect 492 655 493 659
rect 487 654 493 655
rect 534 659 540 660
rect 534 655 535 659
rect 539 658 540 659
rect 543 659 549 660
rect 543 658 544 659
rect 539 656 544 658
rect 539 655 540 656
rect 534 654 540 655
rect 543 655 544 656
rect 548 655 549 659
rect 543 654 549 655
rect 599 659 608 660
rect 599 655 600 659
rect 607 655 608 659
rect 628 658 630 672
rect 655 671 656 675
rect 663 671 664 675
rect 655 670 664 671
rect 711 675 717 676
rect 711 671 712 675
rect 716 674 717 675
rect 774 675 781 676
rect 716 672 746 674
rect 716 671 717 672
rect 711 670 717 671
rect 638 665 644 666
rect 638 661 639 665
rect 643 661 644 665
rect 638 660 644 661
rect 694 665 700 666
rect 694 661 695 665
rect 699 661 700 665
rect 694 660 700 661
rect 655 659 661 660
rect 655 658 656 659
rect 628 656 656 658
rect 599 654 608 655
rect 655 655 656 656
rect 660 655 661 659
rect 655 654 661 655
rect 711 659 720 660
rect 711 655 712 659
rect 719 655 720 659
rect 744 658 746 672
rect 774 671 775 675
rect 780 671 781 675
rect 774 670 781 671
rect 839 675 845 676
rect 839 671 840 675
rect 844 674 845 675
rect 854 675 860 676
rect 854 674 855 675
rect 844 672 855 674
rect 844 671 845 672
rect 839 670 845 671
rect 854 671 855 672
rect 859 671 860 675
rect 903 675 909 676
rect 903 674 904 675
rect 854 670 860 671
rect 873 672 904 674
rect 758 665 764 666
rect 758 661 759 665
rect 763 661 764 665
rect 758 660 764 661
rect 822 665 828 666
rect 822 661 823 665
rect 827 661 828 665
rect 822 660 828 661
rect 775 659 781 660
rect 775 658 776 659
rect 744 656 776 658
rect 711 654 720 655
rect 775 655 776 656
rect 780 655 781 659
rect 775 654 781 655
rect 839 659 845 660
rect 839 655 840 659
rect 844 658 845 659
rect 873 658 875 672
rect 903 671 904 672
rect 908 671 909 675
rect 967 675 973 676
rect 967 674 968 675
rect 903 670 909 671
rect 937 672 968 674
rect 886 665 892 666
rect 886 661 887 665
rect 891 661 892 665
rect 886 660 892 661
rect 844 656 875 658
rect 903 659 909 660
rect 844 655 845 656
rect 839 654 845 655
rect 903 655 904 659
rect 908 658 909 659
rect 937 658 939 672
rect 967 671 968 672
rect 972 671 973 675
rect 967 670 973 671
rect 1031 675 1037 676
rect 1031 671 1032 675
rect 1036 674 1037 675
rect 1095 675 1101 676
rect 1036 672 1066 674
rect 1036 671 1037 672
rect 1031 670 1037 671
rect 950 665 956 666
rect 950 661 951 665
rect 955 661 956 665
rect 950 660 956 661
rect 1014 665 1020 666
rect 1014 661 1015 665
rect 1019 661 1020 665
rect 1014 660 1020 661
rect 908 656 939 658
rect 967 659 973 660
rect 908 655 909 656
rect 903 654 909 655
rect 967 655 968 659
rect 972 655 973 659
rect 967 654 973 655
rect 1031 659 1040 660
rect 1031 655 1032 659
rect 1039 655 1040 659
rect 1064 658 1066 672
rect 1095 671 1096 675
rect 1100 674 1101 675
rect 1126 675 1132 676
rect 1126 674 1127 675
rect 1100 672 1127 674
rect 1100 671 1101 672
rect 1095 670 1101 671
rect 1126 671 1127 672
rect 1131 671 1132 675
rect 1126 670 1132 671
rect 1151 675 1157 676
rect 1151 671 1152 675
rect 1156 674 1157 675
rect 1182 675 1188 676
rect 1182 674 1183 675
rect 1156 672 1183 674
rect 1156 671 1157 672
rect 1151 670 1157 671
rect 1182 671 1183 672
rect 1187 671 1188 675
rect 1207 675 1213 676
rect 1207 674 1208 675
rect 1182 670 1188 671
rect 1200 672 1208 674
rect 1078 665 1084 666
rect 1078 661 1079 665
rect 1083 661 1084 665
rect 1078 660 1084 661
rect 1134 665 1140 666
rect 1134 661 1135 665
rect 1139 661 1140 665
rect 1134 660 1140 661
rect 1190 665 1196 666
rect 1190 661 1191 665
rect 1195 661 1196 665
rect 1190 660 1196 661
rect 1095 659 1101 660
rect 1095 658 1096 659
rect 1064 656 1096 658
rect 1031 654 1040 655
rect 1095 655 1096 656
rect 1100 655 1101 659
rect 1095 654 1101 655
rect 1151 659 1157 660
rect 1151 655 1152 659
rect 1156 658 1157 659
rect 1200 658 1202 672
rect 1207 671 1208 672
rect 1212 671 1213 675
rect 1263 675 1269 676
rect 1263 674 1264 675
rect 1207 670 1213 671
rect 1236 672 1264 674
rect 1156 656 1202 658
rect 1207 659 1213 660
rect 1156 655 1157 656
rect 1151 654 1157 655
rect 1207 655 1208 659
rect 1212 658 1213 659
rect 1236 658 1238 672
rect 1263 671 1264 672
rect 1268 671 1269 675
rect 1319 675 1325 676
rect 1319 674 1320 675
rect 1263 670 1269 671
rect 1292 672 1320 674
rect 1246 665 1252 666
rect 1246 661 1247 665
rect 1251 661 1252 665
rect 1246 660 1252 661
rect 1212 656 1238 658
rect 1263 659 1269 660
rect 1212 655 1213 656
rect 1207 654 1213 655
rect 1263 655 1264 659
rect 1268 658 1269 659
rect 1292 658 1294 672
rect 1319 671 1320 672
rect 1324 671 1325 675
rect 1375 675 1381 676
rect 1375 674 1376 675
rect 1319 670 1325 671
rect 1348 672 1376 674
rect 1348 666 1350 672
rect 1375 671 1376 672
rect 1380 671 1381 675
rect 1375 670 1381 671
rect 1302 665 1308 666
rect 1302 661 1303 665
rect 1307 661 1308 665
rect 1302 660 1308 661
rect 1321 664 1350 666
rect 1358 665 1364 666
rect 1321 660 1323 664
rect 1358 661 1359 665
rect 1363 661 1364 665
rect 1358 660 1364 661
rect 1582 664 1588 665
rect 1582 660 1583 664
rect 1587 660 1588 664
rect 1268 656 1294 658
rect 1319 659 1325 660
rect 1268 655 1269 656
rect 1263 654 1269 655
rect 1319 655 1320 659
rect 1324 655 1325 659
rect 1319 654 1325 655
rect 1350 659 1356 660
rect 1350 655 1351 659
rect 1355 658 1356 659
rect 1375 659 1381 660
rect 1582 659 1588 660
rect 1375 658 1376 659
rect 1355 656 1376 658
rect 1355 655 1356 656
rect 1350 654 1356 655
rect 1375 655 1376 656
rect 1380 655 1381 659
rect 1375 654 1381 655
rect 377 650 379 654
rect 442 651 448 652
rect 442 650 443 651
rect 377 648 443 650
rect 442 647 443 648
rect 447 647 448 651
rect 442 646 448 647
rect 906 651 912 652
rect 906 647 907 651
rect 911 650 912 651
rect 969 650 971 654
rect 911 648 971 650
rect 911 647 912 648
rect 906 646 912 647
rect 992 644 1010 646
rect 178 643 189 644
rect 110 640 116 641
rect 110 636 111 640
rect 115 636 116 640
rect 110 635 116 636
rect 166 639 172 640
rect 166 635 167 639
rect 171 635 172 639
rect 178 639 179 643
rect 183 639 184 643
rect 188 639 189 643
rect 231 643 237 644
rect 231 642 232 643
rect 224 640 232 642
rect 178 638 189 639
rect 214 639 220 640
rect 166 634 172 635
rect 214 635 215 639
rect 219 635 220 639
rect 214 634 220 635
rect 224 630 226 640
rect 231 639 232 640
rect 236 639 237 643
rect 287 643 293 644
rect 287 642 288 643
rect 280 640 288 642
rect 231 638 237 639
rect 270 639 276 640
rect 270 635 271 639
rect 275 635 276 639
rect 270 634 276 635
rect 280 630 282 640
rect 287 639 288 640
rect 292 639 293 643
rect 338 643 349 644
rect 287 638 293 639
rect 326 639 332 640
rect 326 635 327 639
rect 331 635 332 639
rect 338 639 339 643
rect 343 639 344 643
rect 348 639 349 643
rect 399 643 405 644
rect 399 642 400 643
rect 392 640 400 642
rect 338 638 349 639
rect 382 639 388 640
rect 326 634 332 635
rect 382 635 383 639
rect 387 635 388 639
rect 382 634 388 635
rect 392 630 394 640
rect 399 639 400 640
rect 404 639 405 643
rect 442 643 453 644
rect 399 638 405 639
rect 430 639 436 640
rect 430 635 431 639
rect 435 635 436 639
rect 442 639 443 643
rect 447 639 448 643
rect 452 639 453 643
rect 503 643 512 644
rect 442 638 453 639
rect 486 639 492 640
rect 430 634 436 635
rect 486 635 487 639
rect 491 635 492 639
rect 503 639 504 643
rect 511 639 512 643
rect 551 643 557 644
rect 551 642 552 643
rect 544 640 552 642
rect 503 638 512 639
rect 534 639 540 640
rect 486 634 492 635
rect 534 635 535 639
rect 539 635 540 639
rect 534 634 540 635
rect 544 630 546 640
rect 551 639 552 640
rect 556 639 557 643
rect 607 643 613 644
rect 551 638 557 639
rect 590 639 596 640
rect 590 635 591 639
rect 595 635 596 639
rect 607 639 608 643
rect 612 639 613 643
rect 663 643 669 644
rect 607 638 613 639
rect 646 639 652 640
rect 590 634 596 635
rect 609 634 611 638
rect 646 635 647 639
rect 651 635 652 639
rect 663 639 664 643
rect 668 642 669 643
rect 719 643 725 644
rect 668 640 698 642
rect 668 639 669 640
rect 663 638 669 639
rect 646 634 652 635
rect 609 632 642 634
rect 209 628 226 630
rect 259 628 282 630
rect 372 628 394 630
rect 528 628 546 630
rect 640 630 642 632
rect 696 630 698 640
rect 702 639 708 640
rect 702 635 703 639
rect 707 635 708 639
rect 719 639 720 643
rect 724 642 725 643
rect 774 643 781 644
rect 724 640 754 642
rect 724 639 725 640
rect 719 638 725 639
rect 702 634 708 635
rect 752 630 754 640
rect 758 639 764 640
rect 758 635 759 639
rect 763 635 764 639
rect 774 639 775 643
rect 780 639 781 643
rect 834 643 845 644
rect 774 638 781 639
rect 822 639 828 640
rect 758 634 764 635
rect 822 635 823 639
rect 827 635 828 639
rect 834 639 835 643
rect 839 639 840 643
rect 844 639 845 643
rect 903 643 909 644
rect 903 642 904 643
rect 896 640 904 642
rect 834 638 845 639
rect 886 639 892 640
rect 822 634 828 635
rect 886 635 887 639
rect 891 635 892 639
rect 886 634 892 635
rect 896 630 898 640
rect 903 639 904 640
rect 908 639 909 643
rect 959 643 965 644
rect 903 638 909 639
rect 942 639 948 640
rect 942 635 943 639
rect 947 635 948 639
rect 959 639 960 643
rect 964 642 965 643
rect 992 642 994 644
rect 964 640 994 642
rect 964 639 965 640
rect 959 638 965 639
rect 998 639 1004 640
rect 942 634 948 635
rect 998 635 999 639
rect 1003 635 1004 639
rect 998 634 1004 635
rect 640 628 658 630
rect 696 628 714 630
rect 752 628 770 630
rect 873 628 898 630
rect 183 627 189 628
rect 110 623 116 624
rect 110 619 111 623
rect 115 619 116 623
rect 183 623 184 627
rect 188 626 189 627
rect 209 626 211 628
rect 188 624 211 626
rect 231 627 237 628
rect 188 623 189 624
rect 183 622 189 623
rect 231 623 232 627
rect 236 626 237 627
rect 259 626 261 628
rect 236 624 261 626
rect 287 627 293 628
rect 236 623 237 624
rect 231 622 237 623
rect 287 623 288 627
rect 292 626 293 627
rect 302 627 308 628
rect 302 626 303 627
rect 292 624 303 626
rect 292 623 293 624
rect 287 622 293 623
rect 302 623 303 624
rect 307 623 308 627
rect 302 622 308 623
rect 343 627 349 628
rect 343 623 344 627
rect 348 626 349 627
rect 372 626 374 628
rect 348 624 374 626
rect 399 627 408 628
rect 348 623 349 624
rect 343 622 349 623
rect 399 623 400 627
rect 407 623 408 627
rect 399 622 408 623
rect 447 627 456 628
rect 447 623 448 627
rect 455 623 456 627
rect 447 622 456 623
rect 503 627 509 628
rect 503 623 504 627
rect 508 626 509 627
rect 528 626 530 628
rect 508 624 530 626
rect 551 627 557 628
rect 508 623 509 624
rect 503 622 509 623
rect 551 623 552 627
rect 556 626 557 627
rect 574 627 580 628
rect 574 626 575 627
rect 556 624 575 626
rect 556 623 557 624
rect 551 622 557 623
rect 574 623 575 624
rect 579 623 580 627
rect 574 622 580 623
rect 602 627 613 628
rect 602 623 603 627
rect 607 623 608 627
rect 612 623 613 627
rect 656 626 658 628
rect 663 627 669 628
rect 663 626 664 627
rect 656 624 664 626
rect 602 622 613 623
rect 663 623 664 624
rect 668 623 669 627
rect 712 626 714 628
rect 719 627 725 628
rect 719 626 720 627
rect 712 624 720 626
rect 663 622 669 623
rect 719 623 720 624
rect 724 623 725 627
rect 768 626 770 628
rect 775 627 781 628
rect 775 626 776 627
rect 768 624 776 626
rect 719 622 725 623
rect 775 623 776 624
rect 780 623 781 627
rect 775 622 781 623
rect 839 627 845 628
rect 839 623 840 627
rect 844 626 845 627
rect 873 626 875 628
rect 844 624 875 626
rect 903 627 912 628
rect 844 623 845 624
rect 839 622 845 623
rect 903 623 904 627
rect 911 623 912 627
rect 903 622 912 623
rect 959 627 965 628
rect 959 623 960 627
rect 964 626 965 627
rect 990 627 996 628
rect 990 626 991 627
rect 964 624 991 626
rect 964 623 965 624
rect 959 622 965 623
rect 990 623 991 624
rect 995 623 996 627
rect 1008 626 1010 644
rect 1015 643 1021 644
rect 1015 639 1016 643
rect 1020 642 1021 643
rect 1071 643 1077 644
rect 1020 640 1046 642
rect 1020 639 1021 640
rect 1015 638 1021 639
rect 1044 630 1046 640
rect 1054 639 1060 640
rect 1054 635 1055 639
rect 1059 635 1060 639
rect 1071 639 1072 643
rect 1076 642 1077 643
rect 1126 643 1133 644
rect 1076 640 1102 642
rect 1076 639 1077 640
rect 1071 638 1077 639
rect 1054 634 1060 635
rect 1100 630 1102 640
rect 1110 639 1116 640
rect 1110 635 1111 639
rect 1115 635 1116 639
rect 1126 639 1127 643
rect 1132 639 1133 643
rect 1182 643 1189 644
rect 1126 638 1133 639
rect 1166 639 1172 640
rect 1110 634 1116 635
rect 1166 635 1167 639
rect 1171 635 1172 639
rect 1182 639 1183 643
rect 1188 639 1189 643
rect 1231 643 1237 644
rect 1231 642 1232 643
rect 1224 640 1232 642
rect 1182 638 1189 639
rect 1214 639 1220 640
rect 1166 634 1172 635
rect 1214 635 1215 639
rect 1219 635 1220 639
rect 1214 634 1220 635
rect 1224 630 1226 640
rect 1231 639 1232 640
rect 1236 639 1237 643
rect 1287 643 1293 644
rect 1287 642 1288 643
rect 1280 640 1288 642
rect 1231 638 1237 639
rect 1270 639 1276 640
rect 1270 635 1271 639
rect 1275 635 1276 639
rect 1270 634 1276 635
rect 1280 630 1282 640
rect 1287 639 1288 640
rect 1292 639 1293 643
rect 1343 643 1349 644
rect 1343 642 1344 643
rect 1336 640 1344 642
rect 1287 638 1293 639
rect 1326 639 1332 640
rect 1326 635 1327 639
rect 1331 635 1332 639
rect 1326 634 1332 635
rect 1336 630 1338 640
rect 1343 639 1344 640
rect 1348 639 1349 643
rect 1399 643 1405 644
rect 1399 642 1400 643
rect 1392 640 1400 642
rect 1343 638 1349 639
rect 1382 639 1388 640
rect 1382 635 1383 639
rect 1387 635 1388 639
rect 1382 634 1388 635
rect 1392 630 1394 640
rect 1399 639 1400 640
rect 1404 639 1405 643
rect 1455 643 1461 644
rect 1455 642 1456 643
rect 1448 640 1456 642
rect 1399 638 1405 639
rect 1438 639 1444 640
rect 1438 635 1439 639
rect 1443 635 1444 639
rect 1438 634 1444 635
rect 1448 630 1450 640
rect 1455 639 1456 640
rect 1460 639 1461 643
rect 1519 643 1528 644
rect 1455 638 1461 639
rect 1502 639 1508 640
rect 1502 635 1503 639
rect 1507 635 1508 639
rect 1519 639 1520 643
rect 1527 639 1528 643
rect 1559 643 1565 644
rect 1559 642 1560 643
rect 1552 640 1560 642
rect 1519 638 1528 639
rect 1542 639 1548 640
rect 1502 634 1508 635
rect 1542 635 1543 639
rect 1547 635 1548 639
rect 1542 634 1548 635
rect 1552 630 1554 640
rect 1559 639 1560 640
rect 1564 639 1565 643
rect 1559 638 1565 639
rect 1582 640 1588 641
rect 1582 636 1583 640
rect 1587 636 1588 640
rect 1582 635 1588 636
rect 1044 628 1066 630
rect 1100 628 1122 630
rect 1209 628 1226 630
rect 1260 628 1282 630
rect 1316 628 1338 630
rect 1372 628 1394 630
rect 1428 628 1450 630
rect 1540 628 1554 630
rect 1015 627 1021 628
rect 1015 626 1016 627
rect 1008 624 1016 626
rect 990 622 996 623
rect 1015 623 1016 624
rect 1020 623 1021 627
rect 1064 626 1066 628
rect 1071 627 1077 628
rect 1071 626 1072 627
rect 1064 624 1072 626
rect 1015 622 1021 623
rect 1071 623 1072 624
rect 1076 623 1077 627
rect 1120 626 1122 628
rect 1127 627 1133 628
rect 1127 626 1128 627
rect 1120 624 1128 626
rect 1071 622 1077 623
rect 1127 623 1128 624
rect 1132 623 1133 627
rect 1127 622 1133 623
rect 1183 627 1189 628
rect 1183 623 1184 627
rect 1188 626 1189 627
rect 1209 626 1211 628
rect 1188 624 1211 626
rect 1231 627 1237 628
rect 1188 623 1189 624
rect 1183 622 1189 623
rect 1231 623 1232 627
rect 1236 626 1237 627
rect 1260 626 1262 628
rect 1236 624 1262 626
rect 1287 627 1293 628
rect 1236 623 1237 624
rect 1231 622 1237 623
rect 1287 623 1288 627
rect 1292 626 1293 627
rect 1316 626 1318 628
rect 1292 624 1318 626
rect 1343 627 1349 628
rect 1292 623 1293 624
rect 1287 622 1293 623
rect 1343 623 1344 627
rect 1348 626 1349 627
rect 1372 626 1374 628
rect 1348 624 1374 626
rect 1399 627 1405 628
rect 1348 623 1349 624
rect 1343 622 1349 623
rect 1399 623 1400 627
rect 1404 626 1405 627
rect 1428 626 1430 628
rect 1455 627 1461 628
rect 1455 626 1456 627
rect 1404 624 1430 626
rect 1448 624 1456 626
rect 1404 623 1405 624
rect 1399 622 1405 623
rect 110 618 116 619
rect 166 621 172 622
rect 166 617 167 621
rect 171 617 172 621
rect 166 616 172 617
rect 214 621 220 622
rect 214 617 215 621
rect 219 617 220 621
rect 214 616 220 617
rect 270 621 276 622
rect 270 617 271 621
rect 275 617 276 621
rect 270 616 276 617
rect 326 621 332 622
rect 326 617 327 621
rect 331 617 332 621
rect 326 616 332 617
rect 382 621 388 622
rect 382 617 383 621
rect 387 617 388 621
rect 382 616 388 617
rect 430 621 436 622
rect 430 617 431 621
rect 435 617 436 621
rect 430 616 436 617
rect 486 621 492 622
rect 486 617 487 621
rect 491 617 492 621
rect 486 616 492 617
rect 534 621 540 622
rect 534 617 535 621
rect 539 617 540 621
rect 534 616 540 617
rect 590 621 596 622
rect 590 617 591 621
rect 595 617 596 621
rect 590 616 596 617
rect 646 621 652 622
rect 646 617 647 621
rect 651 617 652 621
rect 646 616 652 617
rect 702 621 708 622
rect 702 617 703 621
rect 707 617 708 621
rect 702 616 708 617
rect 758 621 764 622
rect 758 617 759 621
rect 763 617 764 621
rect 758 616 764 617
rect 822 621 828 622
rect 822 617 823 621
rect 827 617 828 621
rect 822 616 828 617
rect 886 621 892 622
rect 886 617 887 621
rect 891 617 892 621
rect 886 616 892 617
rect 942 621 948 622
rect 942 617 943 621
rect 947 617 948 621
rect 942 616 948 617
rect 998 621 1004 622
rect 998 617 999 621
rect 1003 617 1004 621
rect 998 616 1004 617
rect 1054 621 1060 622
rect 1054 617 1055 621
rect 1059 617 1060 621
rect 1054 616 1060 617
rect 1110 621 1116 622
rect 1110 617 1111 621
rect 1115 617 1116 621
rect 1110 616 1116 617
rect 1166 621 1172 622
rect 1166 617 1167 621
rect 1171 617 1172 621
rect 1166 616 1172 617
rect 1214 621 1220 622
rect 1214 617 1215 621
rect 1219 617 1220 621
rect 1214 616 1220 617
rect 1270 621 1276 622
rect 1270 617 1271 621
rect 1275 617 1276 621
rect 1270 616 1276 617
rect 1326 621 1332 622
rect 1326 617 1327 621
rect 1331 617 1332 621
rect 1326 616 1332 617
rect 1382 621 1388 622
rect 1382 617 1383 621
rect 1387 617 1388 621
rect 1382 616 1388 617
rect 1438 621 1444 622
rect 1438 617 1439 621
rect 1443 617 1444 621
rect 1438 616 1444 617
rect 1230 615 1236 616
rect 1230 611 1231 615
rect 1235 614 1236 615
rect 1448 614 1450 624
rect 1455 623 1456 624
rect 1460 623 1461 627
rect 1455 622 1461 623
rect 1519 627 1525 628
rect 1519 623 1520 627
rect 1524 626 1525 627
rect 1540 626 1542 628
rect 1524 624 1542 626
rect 1558 627 1565 628
rect 1524 623 1525 624
rect 1519 622 1525 623
rect 1558 623 1559 627
rect 1564 623 1565 627
rect 1558 622 1565 623
rect 1582 623 1588 624
rect 1502 621 1508 622
rect 1502 617 1503 621
rect 1507 617 1508 621
rect 1502 616 1508 617
rect 1542 621 1548 622
rect 1542 617 1543 621
rect 1547 617 1548 621
rect 1582 619 1583 623
rect 1587 619 1588 623
rect 1582 618 1588 619
rect 1542 616 1548 617
rect 1235 612 1450 614
rect 1235 611 1236 612
rect 1230 610 1236 611
rect 222 607 228 608
rect 110 605 116 606
rect 110 601 111 605
rect 115 601 116 605
rect 222 603 223 607
rect 227 603 228 607
rect 222 602 228 603
rect 254 607 260 608
rect 254 603 255 607
rect 259 603 260 607
rect 254 602 260 603
rect 286 607 292 608
rect 286 603 287 607
rect 291 603 292 607
rect 286 602 292 603
rect 318 607 324 608
rect 318 603 319 607
rect 323 603 324 607
rect 350 607 356 608
rect 318 602 324 603
rect 338 603 344 604
rect 338 602 339 603
rect 110 600 116 601
rect 335 601 339 602
rect 210 599 216 600
rect 210 595 211 599
rect 215 598 216 599
rect 239 599 245 600
rect 239 598 240 599
rect 215 596 240 598
rect 215 595 216 596
rect 210 594 216 595
rect 239 595 240 596
rect 244 595 245 599
rect 271 599 277 600
rect 271 598 272 599
rect 239 594 245 595
rect 264 596 272 598
rect 222 589 228 590
rect 110 588 116 589
rect 110 584 111 588
rect 115 584 116 588
rect 222 585 223 589
rect 227 585 228 589
rect 222 584 228 585
rect 254 589 260 590
rect 254 585 255 589
rect 259 585 260 589
rect 254 584 260 585
rect 110 583 116 584
rect 239 583 245 584
rect 239 579 240 583
rect 244 582 245 583
rect 264 582 266 596
rect 271 595 272 596
rect 276 595 277 599
rect 303 599 309 600
rect 303 598 304 599
rect 271 594 277 595
rect 296 596 304 598
rect 286 589 292 590
rect 286 585 287 589
rect 291 585 292 589
rect 286 584 292 585
rect 244 580 266 582
rect 271 583 277 584
rect 244 579 245 580
rect 239 578 245 579
rect 271 579 272 583
rect 276 582 277 583
rect 296 582 298 596
rect 303 595 304 596
rect 308 595 309 599
rect 335 597 336 601
rect 343 599 344 603
rect 350 603 351 607
rect 355 603 356 607
rect 350 602 356 603
rect 382 607 388 608
rect 382 603 383 607
rect 387 603 388 607
rect 382 602 388 603
rect 422 607 428 608
rect 422 603 423 607
rect 427 603 428 607
rect 422 602 428 603
rect 462 607 468 608
rect 462 603 463 607
rect 467 603 468 607
rect 462 602 468 603
rect 518 607 524 608
rect 518 603 519 607
rect 523 603 524 607
rect 518 602 524 603
rect 582 607 588 608
rect 582 603 583 607
rect 587 603 588 607
rect 646 607 652 608
rect 582 602 588 603
rect 592 604 638 606
rect 340 598 344 599
rect 367 599 373 600
rect 367 598 368 599
rect 340 597 341 598
rect 335 596 341 597
rect 360 596 368 598
rect 303 594 309 595
rect 318 589 324 590
rect 318 585 319 589
rect 323 585 324 589
rect 318 584 324 585
rect 350 589 356 590
rect 350 585 351 589
rect 355 585 356 589
rect 350 584 356 585
rect 276 580 298 582
rect 302 583 309 584
rect 276 579 277 580
rect 271 578 277 579
rect 302 579 303 583
rect 308 579 309 583
rect 302 578 309 579
rect 335 583 341 584
rect 335 579 336 583
rect 340 582 341 583
rect 360 582 362 596
rect 367 595 368 596
rect 372 595 373 599
rect 399 599 405 600
rect 399 598 400 599
rect 367 594 373 595
rect 392 596 400 598
rect 382 589 388 590
rect 382 585 383 589
rect 387 585 388 589
rect 382 584 388 585
rect 340 580 362 582
rect 367 583 373 584
rect 340 579 341 580
rect 335 578 341 579
rect 367 579 368 583
rect 372 582 373 583
rect 392 582 394 596
rect 399 595 400 596
rect 404 595 405 599
rect 399 594 405 595
rect 439 599 448 600
rect 439 595 440 599
rect 447 595 448 599
rect 479 599 485 600
rect 479 598 480 599
rect 439 594 448 595
rect 456 596 480 598
rect 422 589 428 590
rect 422 585 423 589
rect 427 585 428 589
rect 422 584 428 585
rect 372 580 394 582
rect 399 583 405 584
rect 372 579 373 580
rect 367 578 373 579
rect 399 579 400 583
rect 404 582 405 583
rect 414 583 420 584
rect 414 582 415 583
rect 404 580 415 582
rect 404 579 405 580
rect 399 578 405 579
rect 414 579 415 580
rect 419 579 420 583
rect 414 578 420 579
rect 439 583 445 584
rect 439 579 440 583
rect 444 582 445 583
rect 456 582 458 596
rect 479 595 480 596
rect 484 595 485 599
rect 535 599 541 600
rect 535 598 536 599
rect 479 594 485 595
rect 508 596 536 598
rect 462 589 468 590
rect 462 585 463 589
rect 467 585 468 589
rect 462 584 468 585
rect 444 580 458 582
rect 479 583 485 584
rect 444 579 445 580
rect 439 578 445 579
rect 479 579 480 583
rect 484 582 485 583
rect 508 582 510 596
rect 535 595 536 596
rect 540 595 541 599
rect 592 598 594 604
rect 535 594 541 595
rect 568 596 594 598
rect 599 599 605 600
rect 518 589 524 590
rect 518 585 519 589
rect 523 585 524 589
rect 518 584 524 585
rect 484 580 510 582
rect 535 583 541 584
rect 484 579 485 580
rect 479 578 485 579
rect 535 579 536 583
rect 540 582 541 583
rect 568 582 570 596
rect 599 595 600 599
rect 604 598 605 599
rect 636 598 638 604
rect 646 603 647 607
rect 651 603 652 607
rect 646 602 652 603
rect 718 607 724 608
rect 718 603 719 607
rect 723 603 724 607
rect 718 602 724 603
rect 798 607 804 608
rect 798 603 799 607
rect 803 603 804 607
rect 798 602 804 603
rect 886 607 892 608
rect 886 603 887 607
rect 891 603 892 607
rect 886 602 892 603
rect 974 607 980 608
rect 974 603 975 607
rect 979 603 980 607
rect 974 602 980 603
rect 1062 607 1068 608
rect 1062 603 1063 607
rect 1067 603 1068 607
rect 1062 602 1068 603
rect 1142 607 1148 608
rect 1142 603 1143 607
rect 1147 603 1148 607
rect 1142 602 1148 603
rect 1214 607 1220 608
rect 1214 603 1215 607
rect 1219 603 1220 607
rect 1214 602 1220 603
rect 1286 607 1292 608
rect 1286 603 1287 607
rect 1291 603 1292 607
rect 1286 602 1292 603
rect 1350 607 1356 608
rect 1350 603 1351 607
rect 1355 603 1356 607
rect 1350 602 1356 603
rect 1406 607 1412 608
rect 1406 603 1407 607
rect 1411 603 1412 607
rect 1406 602 1412 603
rect 1454 607 1460 608
rect 1454 603 1455 607
rect 1459 603 1460 607
rect 1454 602 1460 603
rect 1510 607 1516 608
rect 1510 603 1511 607
rect 1515 603 1516 607
rect 1510 602 1516 603
rect 1542 607 1548 608
rect 1542 603 1543 607
rect 1547 603 1548 607
rect 1542 602 1548 603
rect 1582 605 1588 606
rect 1582 601 1583 605
rect 1587 601 1588 605
rect 1582 600 1588 601
rect 663 599 669 600
rect 663 598 664 599
rect 604 596 634 598
rect 636 596 664 598
rect 604 595 605 596
rect 599 594 605 595
rect 582 589 588 590
rect 582 585 583 589
rect 587 585 588 589
rect 582 584 588 585
rect 540 580 570 582
rect 574 583 580 584
rect 540 579 541 580
rect 535 578 541 579
rect 574 579 575 583
rect 579 582 580 583
rect 599 583 605 584
rect 599 582 600 583
rect 579 580 600 582
rect 579 579 580 580
rect 574 578 580 579
rect 599 579 600 580
rect 604 579 605 583
rect 632 582 634 596
rect 663 595 664 596
rect 668 595 669 599
rect 663 594 669 595
rect 735 599 741 600
rect 735 595 736 599
rect 740 598 741 599
rect 815 599 821 600
rect 740 596 810 598
rect 740 595 741 596
rect 735 594 741 595
rect 646 589 652 590
rect 646 585 647 589
rect 651 585 652 589
rect 646 584 652 585
rect 718 589 724 590
rect 718 585 719 589
rect 723 585 724 589
rect 718 584 724 585
rect 798 589 804 590
rect 798 585 799 589
rect 803 585 804 589
rect 798 584 804 585
rect 663 583 669 584
rect 663 582 664 583
rect 632 580 664 582
rect 599 578 605 579
rect 663 579 664 580
rect 668 579 669 583
rect 663 578 669 579
rect 735 583 741 584
rect 735 579 736 583
rect 740 579 741 583
rect 808 582 810 596
rect 815 595 816 599
rect 820 598 821 599
rect 834 599 840 600
rect 834 598 835 599
rect 820 596 835 598
rect 820 595 821 596
rect 815 594 821 595
rect 834 595 835 596
rect 839 595 840 599
rect 834 594 840 595
rect 846 599 852 600
rect 846 595 847 599
rect 851 598 852 599
rect 903 599 909 600
rect 903 598 904 599
rect 851 596 904 598
rect 851 595 852 596
rect 846 594 852 595
rect 903 595 904 596
rect 908 595 909 599
rect 903 594 909 595
rect 991 599 997 600
rect 991 595 992 599
rect 996 598 997 599
rect 1079 599 1085 600
rect 996 596 1038 598
rect 996 595 997 596
rect 991 594 997 595
rect 886 589 892 590
rect 886 585 887 589
rect 891 585 892 589
rect 886 584 892 585
rect 974 589 980 590
rect 974 585 975 589
rect 979 585 980 589
rect 974 584 980 585
rect 815 583 821 584
rect 815 582 816 583
rect 808 580 816 582
rect 735 578 741 579
rect 815 579 816 580
rect 820 579 821 583
rect 863 583 869 584
rect 815 578 821 579
rect 846 579 852 580
rect 737 576 810 578
rect 279 575 285 576
rect 207 571 216 572
rect 110 568 116 569
rect 110 564 111 568
rect 115 564 116 568
rect 110 563 116 564
rect 190 567 196 568
rect 190 563 191 567
rect 195 563 196 567
rect 207 567 208 571
rect 215 567 216 571
rect 271 571 277 572
rect 271 570 272 571
rect 264 568 272 570
rect 207 566 216 567
rect 254 567 260 568
rect 190 562 196 563
rect 254 563 255 567
rect 259 563 260 567
rect 254 562 260 563
rect 264 558 266 568
rect 271 567 272 568
rect 276 567 277 571
rect 279 571 280 575
rect 284 574 285 575
rect 447 575 453 576
rect 284 572 338 574
rect 284 571 285 572
rect 279 570 285 571
rect 336 570 338 572
rect 343 571 349 572
rect 343 570 344 571
rect 336 568 344 570
rect 271 566 277 567
rect 326 567 332 568
rect 326 563 327 567
rect 331 563 332 567
rect 343 567 344 568
rect 348 567 349 571
rect 415 571 421 572
rect 343 566 349 567
rect 398 567 404 568
rect 326 562 332 563
rect 398 563 399 567
rect 403 563 404 567
rect 415 567 416 571
rect 420 570 421 571
rect 447 571 448 575
rect 452 574 453 575
rect 808 574 810 576
rect 846 575 847 579
rect 851 575 852 579
rect 863 579 864 583
rect 868 582 869 583
rect 903 583 909 584
rect 903 582 904 583
rect 868 580 904 582
rect 868 579 869 580
rect 863 578 869 579
rect 903 579 904 580
rect 908 579 909 583
rect 903 578 909 579
rect 990 583 997 584
rect 990 579 991 583
rect 996 579 997 583
rect 1036 582 1038 596
rect 1079 595 1080 599
rect 1084 598 1085 599
rect 1159 599 1165 600
rect 1084 596 1122 598
rect 1084 595 1085 596
rect 1079 594 1085 595
rect 1062 589 1068 590
rect 1062 585 1063 589
rect 1067 585 1068 589
rect 1062 584 1068 585
rect 1079 583 1085 584
rect 1079 582 1080 583
rect 1036 580 1080 582
rect 990 578 997 579
rect 1079 579 1080 580
rect 1084 579 1085 583
rect 1120 582 1122 596
rect 1159 595 1160 599
rect 1164 598 1165 599
rect 1182 599 1188 600
rect 1182 598 1183 599
rect 1164 596 1183 598
rect 1164 595 1165 596
rect 1159 594 1165 595
rect 1182 595 1183 596
rect 1187 595 1188 599
rect 1182 594 1188 595
rect 1231 599 1237 600
rect 1231 595 1232 599
rect 1236 598 1237 599
rect 1303 599 1309 600
rect 1236 596 1270 598
rect 1236 595 1237 596
rect 1231 594 1237 595
rect 1142 589 1148 590
rect 1142 585 1143 589
rect 1147 585 1148 589
rect 1142 584 1148 585
rect 1214 589 1220 590
rect 1214 585 1215 589
rect 1219 585 1220 589
rect 1214 584 1220 585
rect 1230 587 1236 588
rect 1159 583 1165 584
rect 1159 582 1160 583
rect 1120 580 1160 582
rect 1079 578 1085 579
rect 1159 579 1160 580
rect 1164 579 1165 583
rect 1230 583 1231 587
rect 1235 586 1236 587
rect 1235 585 1237 586
rect 1230 582 1232 583
rect 1231 581 1232 582
rect 1236 581 1237 585
rect 1231 580 1237 581
rect 1268 582 1270 596
rect 1303 595 1304 599
rect 1308 598 1309 599
rect 1367 599 1373 600
rect 1308 596 1338 598
rect 1308 595 1309 596
rect 1303 594 1309 595
rect 1286 589 1292 590
rect 1286 585 1287 589
rect 1291 585 1292 589
rect 1286 584 1292 585
rect 1303 583 1309 584
rect 1303 582 1304 583
rect 1268 580 1304 582
rect 1159 578 1165 579
rect 1303 579 1304 580
rect 1308 579 1309 583
rect 1336 582 1338 596
rect 1367 595 1368 599
rect 1372 598 1373 599
rect 1423 599 1429 600
rect 1372 596 1398 598
rect 1372 595 1373 596
rect 1367 594 1373 595
rect 1350 589 1356 590
rect 1350 585 1351 589
rect 1355 585 1356 589
rect 1350 584 1356 585
rect 1367 583 1373 584
rect 1367 582 1368 583
rect 1336 580 1368 582
rect 1303 578 1309 579
rect 1367 579 1368 580
rect 1372 579 1373 583
rect 1396 582 1398 596
rect 1423 595 1424 599
rect 1428 598 1429 599
rect 1471 599 1477 600
rect 1428 596 1442 598
rect 1428 595 1429 596
rect 1423 594 1429 595
rect 1406 589 1412 590
rect 1406 585 1407 589
rect 1411 585 1412 589
rect 1406 584 1412 585
rect 1423 583 1429 584
rect 1423 582 1424 583
rect 1396 580 1424 582
rect 1367 578 1373 579
rect 1423 579 1424 580
rect 1428 579 1429 583
rect 1440 582 1442 596
rect 1471 595 1472 599
rect 1476 598 1477 599
rect 1486 599 1492 600
rect 1486 598 1487 599
rect 1476 596 1487 598
rect 1476 595 1477 596
rect 1471 594 1477 595
rect 1486 595 1487 596
rect 1491 595 1492 599
rect 1486 594 1492 595
rect 1522 599 1533 600
rect 1522 595 1523 599
rect 1527 595 1528 599
rect 1532 595 1533 599
rect 1522 594 1533 595
rect 1559 599 1565 600
rect 1559 595 1560 599
rect 1564 598 1565 599
rect 1567 599 1573 600
rect 1567 598 1568 599
rect 1564 596 1568 598
rect 1564 595 1565 596
rect 1559 594 1565 595
rect 1567 595 1568 596
rect 1572 595 1573 599
rect 1567 594 1573 595
rect 1454 589 1460 590
rect 1454 585 1455 589
rect 1459 585 1460 589
rect 1454 584 1460 585
rect 1510 589 1516 590
rect 1510 585 1511 589
rect 1515 585 1516 589
rect 1510 584 1516 585
rect 1542 589 1548 590
rect 1542 585 1543 589
rect 1547 585 1548 589
rect 1542 584 1548 585
rect 1582 588 1588 589
rect 1582 584 1583 588
rect 1587 584 1588 588
rect 1471 583 1477 584
rect 1471 582 1472 583
rect 1440 580 1472 582
rect 1423 578 1429 579
rect 1471 579 1472 580
rect 1476 579 1477 583
rect 1471 578 1477 579
rect 1526 583 1533 584
rect 1526 579 1527 583
rect 1532 579 1533 583
rect 1526 578 1533 579
rect 1558 583 1565 584
rect 1582 583 1588 584
rect 1558 579 1559 583
rect 1564 579 1565 583
rect 1558 578 1565 579
rect 846 574 852 575
rect 1550 575 1556 576
rect 1550 574 1551 575
rect 452 572 491 574
rect 808 572 850 574
rect 1527 573 1551 574
rect 452 571 453 572
rect 447 570 453 571
rect 487 571 493 572
rect 420 568 442 570
rect 420 567 421 568
rect 415 566 421 567
rect 398 562 404 563
rect 209 556 266 558
rect 440 558 442 568
rect 470 567 476 568
rect 470 563 471 567
rect 475 563 476 567
rect 487 567 488 571
rect 492 567 493 571
rect 551 571 557 572
rect 487 566 493 567
rect 534 567 540 568
rect 470 562 476 563
rect 534 563 535 567
rect 539 563 540 567
rect 551 567 552 571
rect 556 570 557 571
rect 590 571 596 572
rect 590 570 591 571
rect 556 568 591 570
rect 556 567 557 568
rect 551 566 557 567
rect 590 567 591 568
rect 595 567 596 571
rect 615 571 621 572
rect 615 570 616 571
rect 608 568 616 570
rect 590 566 596 567
rect 598 567 604 568
rect 534 562 540 563
rect 598 563 599 567
rect 603 563 604 567
rect 598 562 604 563
rect 608 558 610 568
rect 615 567 616 568
rect 620 567 621 571
rect 679 571 685 572
rect 679 570 680 571
rect 672 568 680 570
rect 615 566 621 567
rect 662 567 668 568
rect 662 563 663 567
rect 667 563 668 567
rect 662 562 668 563
rect 672 558 674 568
rect 679 567 680 568
rect 684 567 685 571
rect 743 571 749 572
rect 743 570 744 571
rect 736 568 744 570
rect 679 566 685 567
rect 726 567 732 568
rect 726 563 727 567
rect 731 563 732 567
rect 726 562 732 563
rect 736 558 738 568
rect 743 567 744 568
rect 748 567 749 571
rect 799 571 805 572
rect 799 570 800 571
rect 792 568 800 570
rect 743 566 749 567
rect 782 567 788 568
rect 782 563 783 567
rect 787 563 788 567
rect 782 562 788 563
rect 792 558 794 568
rect 799 567 800 568
rect 804 567 805 571
rect 855 571 861 572
rect 855 570 856 571
rect 848 568 856 570
rect 799 566 805 567
rect 838 567 844 568
rect 838 563 839 567
rect 843 563 844 567
rect 838 562 844 563
rect 848 558 850 568
rect 855 567 856 568
rect 860 567 861 571
rect 919 571 925 572
rect 855 566 861 567
rect 902 567 908 568
rect 902 563 903 567
rect 907 563 908 567
rect 919 567 920 571
rect 924 570 925 571
rect 983 571 989 572
rect 924 568 962 570
rect 924 567 925 568
rect 919 566 925 567
rect 902 562 908 563
rect 440 556 491 558
rect 584 556 610 558
rect 648 556 674 558
rect 681 556 738 558
rect 772 556 794 558
rect 828 556 850 558
rect 960 558 962 568
rect 966 567 972 568
rect 966 563 967 567
rect 971 563 972 567
rect 983 567 984 571
rect 988 570 989 571
rect 1055 571 1061 572
rect 988 568 1030 570
rect 988 567 989 568
rect 983 566 989 567
rect 966 562 972 563
rect 1028 558 1030 568
rect 1038 567 1044 568
rect 1038 563 1039 567
rect 1043 563 1044 567
rect 1055 567 1056 571
rect 1060 567 1061 571
rect 1119 571 1125 572
rect 1055 566 1061 567
rect 1102 567 1108 568
rect 1038 562 1044 563
rect 1057 562 1059 566
rect 1102 563 1103 567
rect 1107 563 1108 567
rect 1119 567 1120 571
rect 1124 570 1125 571
rect 1182 571 1189 572
rect 1124 568 1162 570
rect 1124 567 1125 568
rect 1119 566 1125 567
rect 1102 562 1108 563
rect 1057 560 1082 562
rect 1080 558 1082 560
rect 1160 558 1162 568
rect 1166 567 1172 568
rect 1166 563 1167 567
rect 1171 563 1172 567
rect 1182 567 1183 571
rect 1188 567 1189 571
rect 1247 571 1253 572
rect 1182 566 1189 567
rect 1230 567 1236 568
rect 1166 562 1172 563
rect 1230 563 1231 567
rect 1235 563 1236 567
rect 1247 567 1248 571
rect 1252 570 1253 571
rect 1303 571 1309 572
rect 1252 568 1282 570
rect 1252 567 1253 568
rect 1247 566 1253 567
rect 1230 562 1236 563
rect 1191 559 1197 560
rect 960 556 978 558
rect 1028 556 1059 558
rect 1080 556 1114 558
rect 1160 556 1178 558
rect 207 555 213 556
rect 110 551 116 552
rect 110 547 111 551
rect 115 547 116 551
rect 207 551 208 555
rect 212 551 213 555
rect 207 550 213 551
rect 271 555 277 556
rect 271 551 272 555
rect 276 554 277 555
rect 279 555 285 556
rect 279 554 280 555
rect 276 552 280 554
rect 276 551 277 552
rect 271 550 277 551
rect 279 551 280 552
rect 284 551 285 555
rect 279 550 285 551
rect 338 555 349 556
rect 338 551 339 555
rect 343 551 344 555
rect 348 551 349 555
rect 338 550 349 551
rect 414 555 421 556
rect 414 551 415 555
rect 420 551 421 555
rect 414 550 421 551
rect 487 555 493 556
rect 487 551 488 555
rect 492 551 493 555
rect 487 550 493 551
rect 551 555 557 556
rect 551 551 552 555
rect 556 554 557 555
rect 584 554 586 556
rect 556 552 586 554
rect 615 555 621 556
rect 556 551 557 552
rect 551 550 557 551
rect 615 551 616 555
rect 620 554 621 555
rect 648 554 650 556
rect 620 552 650 554
rect 679 555 685 556
rect 620 551 621 552
rect 615 550 621 551
rect 679 551 680 555
rect 684 551 685 555
rect 679 550 685 551
rect 743 555 749 556
rect 743 551 744 555
rect 748 554 749 555
rect 772 554 774 556
rect 748 552 774 554
rect 799 555 805 556
rect 748 551 749 552
rect 743 550 749 551
rect 799 551 800 555
rect 804 554 805 555
rect 828 554 830 556
rect 804 552 830 554
rect 855 555 861 556
rect 804 551 805 552
rect 799 550 805 551
rect 855 551 856 555
rect 860 554 861 555
rect 863 555 869 556
rect 863 554 864 555
rect 860 552 864 554
rect 860 551 861 552
rect 855 550 861 551
rect 863 551 864 552
rect 868 551 869 555
rect 863 550 869 551
rect 919 555 925 556
rect 919 551 920 555
rect 924 554 925 555
rect 951 555 957 556
rect 951 554 952 555
rect 924 552 952 554
rect 924 551 925 552
rect 919 550 925 551
rect 951 551 952 552
rect 956 551 957 555
rect 976 554 978 556
rect 983 555 989 556
rect 983 554 984 555
rect 976 552 984 554
rect 951 550 957 551
rect 983 551 984 552
rect 988 551 989 555
rect 983 550 989 551
rect 1055 555 1061 556
rect 1055 551 1056 555
rect 1060 551 1061 555
rect 1112 554 1114 556
rect 1119 555 1125 556
rect 1119 554 1120 555
rect 1112 552 1120 554
rect 1055 550 1061 551
rect 1119 551 1120 552
rect 1124 551 1125 555
rect 1176 554 1178 556
rect 1183 555 1189 556
rect 1183 554 1184 555
rect 1176 552 1184 554
rect 1119 550 1125 551
rect 1183 551 1184 552
rect 1188 551 1189 555
rect 1191 555 1192 559
rect 1196 558 1197 559
rect 1280 558 1282 568
rect 1286 567 1292 568
rect 1286 563 1287 567
rect 1291 563 1292 567
rect 1303 567 1304 571
rect 1308 570 1309 571
rect 1351 571 1357 572
rect 1308 568 1330 570
rect 1308 567 1309 568
rect 1303 566 1309 567
rect 1286 562 1292 563
rect 1328 558 1330 568
rect 1334 567 1340 568
rect 1334 563 1335 567
rect 1339 563 1340 567
rect 1351 567 1352 571
rect 1356 570 1357 571
rect 1399 571 1405 572
rect 1356 568 1379 570
rect 1356 567 1357 568
rect 1351 566 1357 567
rect 1334 562 1340 563
rect 1377 558 1379 568
rect 1382 567 1388 568
rect 1382 563 1383 567
rect 1387 563 1388 567
rect 1399 567 1400 571
rect 1404 570 1405 571
rect 1439 571 1445 572
rect 1404 568 1418 570
rect 1404 567 1405 568
rect 1399 566 1405 567
rect 1382 562 1388 563
rect 1416 558 1418 568
rect 1422 567 1428 568
rect 1422 563 1423 567
rect 1427 563 1428 567
rect 1439 567 1440 571
rect 1444 570 1445 571
rect 1486 571 1493 572
rect 1444 568 1461 570
rect 1444 567 1445 568
rect 1439 566 1445 567
rect 1422 562 1428 563
rect 1459 558 1461 568
rect 1470 567 1476 568
rect 1470 563 1471 567
rect 1475 563 1476 567
rect 1486 567 1487 571
rect 1492 567 1493 571
rect 1527 569 1528 573
rect 1532 572 1551 573
rect 1532 569 1533 572
rect 1550 571 1551 572
rect 1555 571 1556 575
rect 1550 570 1556 571
rect 1559 571 1565 572
rect 1527 568 1533 569
rect 1486 566 1493 567
rect 1510 567 1516 568
rect 1470 562 1476 563
rect 1510 563 1511 567
rect 1515 563 1516 567
rect 1510 562 1516 563
rect 1542 567 1548 568
rect 1542 563 1543 567
rect 1547 563 1548 567
rect 1559 567 1560 571
rect 1564 570 1565 571
rect 1567 571 1573 572
rect 1567 570 1568 571
rect 1564 568 1568 570
rect 1564 567 1565 568
rect 1559 566 1565 567
rect 1567 567 1568 568
rect 1572 567 1573 571
rect 1567 566 1573 567
rect 1582 568 1588 569
rect 1582 564 1583 568
rect 1587 564 1588 568
rect 1582 563 1588 564
rect 1542 562 1548 563
rect 1196 556 1242 558
rect 1280 556 1298 558
rect 1328 556 1346 558
rect 1377 556 1394 558
rect 1416 556 1434 558
rect 1459 556 1482 558
rect 1196 555 1197 556
rect 1191 554 1197 555
rect 1240 554 1242 556
rect 1247 555 1253 556
rect 1247 554 1248 555
rect 1240 552 1248 554
rect 1183 550 1189 551
rect 1247 551 1248 552
rect 1252 551 1253 555
rect 1296 554 1298 556
rect 1303 555 1309 556
rect 1303 554 1304 555
rect 1296 552 1304 554
rect 1247 550 1253 551
rect 1303 551 1304 552
rect 1308 551 1309 555
rect 1344 554 1346 556
rect 1351 555 1357 556
rect 1351 554 1352 555
rect 1344 552 1352 554
rect 1303 550 1309 551
rect 1351 551 1352 552
rect 1356 551 1357 555
rect 1392 554 1394 556
rect 1399 555 1405 556
rect 1399 554 1400 555
rect 1392 552 1400 554
rect 1351 550 1357 551
rect 1399 551 1400 552
rect 1404 551 1405 555
rect 1432 554 1434 556
rect 1439 555 1445 556
rect 1439 554 1440 555
rect 1432 552 1440 554
rect 1399 550 1405 551
rect 1439 551 1440 552
rect 1444 551 1445 555
rect 1480 554 1482 556
rect 1487 555 1493 556
rect 1487 554 1488 555
rect 1480 552 1488 554
rect 1439 550 1445 551
rect 1487 551 1488 552
rect 1492 551 1493 555
rect 1487 550 1493 551
rect 1526 555 1533 556
rect 1526 551 1527 555
rect 1532 551 1533 555
rect 1526 550 1533 551
rect 1558 555 1565 556
rect 1558 551 1559 555
rect 1564 551 1565 555
rect 1558 550 1565 551
rect 1582 551 1588 552
rect 110 546 116 547
rect 190 549 196 550
rect 190 545 191 549
rect 195 545 196 549
rect 190 544 196 545
rect 254 549 260 550
rect 254 545 255 549
rect 259 545 260 549
rect 254 544 260 545
rect 326 549 332 550
rect 326 545 327 549
rect 331 545 332 549
rect 326 544 332 545
rect 398 549 404 550
rect 398 545 399 549
rect 403 545 404 549
rect 398 544 404 545
rect 470 549 476 550
rect 470 545 471 549
rect 475 545 476 549
rect 470 544 476 545
rect 534 549 540 550
rect 534 545 535 549
rect 539 545 540 549
rect 534 544 540 545
rect 598 549 604 550
rect 598 545 599 549
rect 603 545 604 549
rect 598 544 604 545
rect 662 549 668 550
rect 662 545 663 549
rect 667 545 668 549
rect 662 544 668 545
rect 726 549 732 550
rect 726 545 727 549
rect 731 545 732 549
rect 726 544 732 545
rect 782 549 788 550
rect 782 545 783 549
rect 787 545 788 549
rect 782 544 788 545
rect 838 549 844 550
rect 838 545 839 549
rect 843 545 844 549
rect 838 544 844 545
rect 902 549 908 550
rect 902 545 903 549
rect 907 545 908 549
rect 902 544 908 545
rect 966 549 972 550
rect 966 545 967 549
rect 971 545 972 549
rect 966 544 972 545
rect 1038 549 1044 550
rect 1038 545 1039 549
rect 1043 545 1044 549
rect 1038 544 1044 545
rect 1102 549 1108 550
rect 1102 545 1103 549
rect 1107 545 1108 549
rect 1102 544 1108 545
rect 1166 549 1172 550
rect 1166 545 1167 549
rect 1171 545 1172 549
rect 1166 544 1172 545
rect 1230 549 1236 550
rect 1230 545 1231 549
rect 1235 545 1236 549
rect 1230 544 1236 545
rect 1286 549 1292 550
rect 1286 545 1287 549
rect 1291 545 1292 549
rect 1286 544 1292 545
rect 1334 549 1340 550
rect 1334 545 1335 549
rect 1339 545 1340 549
rect 1334 544 1340 545
rect 1382 549 1388 550
rect 1382 545 1383 549
rect 1387 545 1388 549
rect 1382 544 1388 545
rect 1422 549 1428 550
rect 1422 545 1423 549
rect 1427 545 1428 549
rect 1422 544 1428 545
rect 1470 549 1476 550
rect 1470 545 1471 549
rect 1475 545 1476 549
rect 1470 544 1476 545
rect 1510 549 1516 550
rect 1510 545 1511 549
rect 1515 545 1516 549
rect 1510 544 1516 545
rect 1542 549 1548 550
rect 1542 545 1543 549
rect 1547 545 1548 549
rect 1582 547 1583 551
rect 1587 547 1588 551
rect 1582 546 1588 547
rect 1542 544 1548 545
rect 590 543 596 544
rect 590 539 591 543
rect 595 542 596 543
rect 910 543 916 544
rect 595 540 762 542
rect 595 539 596 540
rect 590 538 596 539
rect 134 535 140 536
rect 110 533 116 534
rect 110 529 111 533
rect 115 529 116 533
rect 134 531 135 535
rect 139 531 140 535
rect 134 530 140 531
rect 174 535 180 536
rect 174 531 175 535
rect 179 531 180 535
rect 174 530 180 531
rect 230 535 236 536
rect 230 531 231 535
rect 235 531 236 535
rect 230 530 236 531
rect 294 535 300 536
rect 294 531 295 535
rect 299 531 300 535
rect 294 530 300 531
rect 358 535 364 536
rect 358 531 359 535
rect 363 531 364 535
rect 358 530 364 531
rect 422 535 428 536
rect 422 531 423 535
rect 427 531 428 535
rect 422 530 428 531
rect 478 535 484 536
rect 478 531 479 535
rect 483 531 484 535
rect 478 530 484 531
rect 542 535 548 536
rect 542 531 543 535
rect 547 531 548 535
rect 542 530 548 531
rect 598 535 604 536
rect 598 531 599 535
rect 603 531 604 535
rect 598 530 604 531
rect 654 535 660 536
rect 654 531 655 535
rect 659 531 660 535
rect 654 530 660 531
rect 710 535 716 536
rect 710 531 711 535
rect 715 531 716 535
rect 710 530 716 531
rect 110 528 116 529
rect 150 527 157 528
rect 150 523 151 527
rect 156 523 157 527
rect 191 527 197 528
rect 191 526 192 527
rect 150 522 157 523
rect 168 524 192 526
rect 134 517 140 518
rect 110 516 116 517
rect 110 512 111 516
rect 115 512 116 516
rect 134 513 135 517
rect 139 513 140 517
rect 134 512 140 513
rect 110 511 116 512
rect 151 511 157 512
rect 151 507 152 511
rect 156 510 157 511
rect 168 510 170 524
rect 191 523 192 524
rect 196 523 197 527
rect 247 527 253 528
rect 247 526 248 527
rect 191 522 197 523
rect 220 524 248 526
rect 174 517 180 518
rect 174 513 175 517
rect 179 513 180 517
rect 174 512 180 513
rect 156 508 170 510
rect 191 511 197 512
rect 156 507 157 508
rect 151 506 157 507
rect 191 507 192 511
rect 196 510 197 511
rect 220 510 222 524
rect 247 523 248 524
rect 252 523 253 527
rect 311 527 317 528
rect 311 526 312 527
rect 247 522 253 523
rect 259 524 312 526
rect 230 517 236 518
rect 230 513 231 517
rect 235 513 236 517
rect 230 512 236 513
rect 196 508 222 510
rect 247 511 253 512
rect 196 507 197 508
rect 191 506 197 507
rect 247 507 248 511
rect 252 510 253 511
rect 259 510 261 524
rect 311 523 312 524
rect 316 523 317 527
rect 311 522 317 523
rect 375 527 381 528
rect 375 523 376 527
rect 380 526 381 527
rect 439 527 445 528
rect 380 524 434 526
rect 380 523 381 524
rect 375 522 381 523
rect 294 517 300 518
rect 294 513 295 517
rect 299 513 300 517
rect 358 517 364 518
rect 294 512 300 513
rect 338 515 344 516
rect 252 508 261 510
rect 311 511 317 512
rect 252 507 253 508
rect 247 506 253 507
rect 311 507 312 511
rect 316 510 317 511
rect 338 511 339 515
rect 343 511 344 515
rect 358 513 359 517
rect 363 513 364 517
rect 358 512 364 513
rect 422 517 428 518
rect 422 513 423 517
rect 427 513 428 517
rect 422 512 428 513
rect 338 510 344 511
rect 366 511 372 512
rect 316 508 342 510
rect 316 507 317 508
rect 311 506 317 507
rect 366 507 367 511
rect 371 510 372 511
rect 375 511 381 512
rect 375 510 376 511
rect 371 508 376 510
rect 371 507 372 508
rect 366 506 372 507
rect 375 507 376 508
rect 380 507 381 511
rect 432 510 434 524
rect 439 523 440 527
rect 444 526 445 527
rect 447 527 453 528
rect 447 526 448 527
rect 444 524 448 526
rect 444 523 445 524
rect 439 522 445 523
rect 447 523 448 524
rect 452 523 453 527
rect 447 522 453 523
rect 495 527 501 528
rect 495 523 496 527
rect 500 526 501 527
rect 559 527 565 528
rect 500 524 530 526
rect 500 523 501 524
rect 495 522 501 523
rect 478 517 484 518
rect 478 513 479 517
rect 483 513 484 517
rect 478 512 484 513
rect 439 511 445 512
rect 439 510 440 511
rect 432 508 440 510
rect 375 506 381 507
rect 439 507 440 508
rect 444 507 445 511
rect 439 506 445 507
rect 495 511 501 512
rect 495 507 496 511
rect 500 510 501 511
rect 528 510 530 524
rect 559 523 560 527
rect 564 526 565 527
rect 615 527 621 528
rect 564 524 590 526
rect 564 523 565 524
rect 559 522 565 523
rect 542 517 548 518
rect 542 513 543 517
rect 547 513 548 517
rect 542 512 548 513
rect 559 511 565 512
rect 559 510 560 511
rect 500 508 526 510
rect 528 508 560 510
rect 500 507 501 508
rect 495 506 501 507
rect 524 506 526 508
rect 559 507 560 508
rect 564 507 565 511
rect 588 510 590 524
rect 615 523 616 527
rect 620 526 621 527
rect 671 527 677 528
rect 620 524 646 526
rect 620 523 621 524
rect 615 522 621 523
rect 598 517 604 518
rect 598 513 599 517
rect 603 513 604 517
rect 598 512 604 513
rect 615 511 621 512
rect 615 510 616 511
rect 588 508 616 510
rect 559 506 565 507
rect 615 507 616 508
rect 620 507 621 511
rect 644 510 646 524
rect 671 523 672 527
rect 676 526 677 527
rect 727 527 733 528
rect 676 524 722 526
rect 676 523 677 524
rect 671 522 677 523
rect 654 517 660 518
rect 654 513 655 517
rect 659 513 660 517
rect 654 512 660 513
rect 710 517 716 518
rect 710 513 711 517
rect 715 513 716 517
rect 710 512 716 513
rect 671 511 677 512
rect 671 510 672 511
rect 644 508 672 510
rect 615 506 621 507
rect 671 507 672 508
rect 676 507 677 511
rect 720 510 722 524
rect 727 523 728 527
rect 732 526 733 527
rect 760 526 762 540
rect 910 539 911 543
rect 915 542 916 543
rect 915 540 1082 542
rect 915 539 916 540
rect 910 538 916 539
rect 766 535 772 536
rect 766 531 767 535
rect 771 531 772 535
rect 766 530 772 531
rect 830 535 836 536
rect 830 531 831 535
rect 835 531 836 535
rect 830 530 836 531
rect 894 535 900 536
rect 894 531 895 535
rect 899 531 900 535
rect 894 530 900 531
rect 966 535 972 536
rect 966 531 967 535
rect 971 531 972 535
rect 966 530 972 531
rect 1030 535 1036 536
rect 1030 531 1031 535
rect 1035 531 1036 535
rect 1030 530 1036 531
rect 783 527 789 528
rect 783 526 784 527
rect 732 524 758 526
rect 760 524 784 526
rect 732 523 733 524
rect 727 522 733 523
rect 727 511 733 512
rect 727 510 728 511
rect 720 508 728 510
rect 671 506 677 507
rect 694 507 700 508
rect 694 506 695 507
rect 524 504 554 506
rect 552 502 554 504
rect 577 504 611 506
rect 577 502 579 504
rect 552 500 579 502
rect 609 502 611 504
rect 632 504 666 506
rect 632 502 634 504
rect 609 500 634 502
rect 664 502 666 504
rect 688 504 695 506
rect 688 502 690 504
rect 694 503 695 504
rect 699 503 700 507
rect 727 507 728 508
rect 732 507 733 511
rect 756 510 758 524
rect 783 523 784 524
rect 788 523 789 527
rect 783 522 789 523
rect 791 527 797 528
rect 791 523 792 527
rect 796 526 797 527
rect 847 527 853 528
rect 847 526 848 527
rect 796 524 848 526
rect 796 523 797 524
rect 791 522 797 523
rect 847 523 848 524
rect 852 523 853 527
rect 911 527 917 528
rect 911 526 912 527
rect 847 522 853 523
rect 884 524 912 526
rect 766 517 772 518
rect 766 513 767 517
rect 771 513 772 517
rect 766 512 772 513
rect 830 517 836 518
rect 830 513 831 517
rect 835 513 836 517
rect 830 512 836 513
rect 783 511 789 512
rect 783 510 784 511
rect 756 508 784 510
rect 727 506 733 507
rect 783 507 784 508
rect 788 507 789 511
rect 783 506 789 507
rect 847 511 853 512
rect 847 507 848 511
rect 852 510 853 511
rect 884 510 886 524
rect 911 523 912 524
rect 916 523 917 527
rect 911 522 917 523
rect 983 527 989 528
rect 983 523 984 527
rect 988 526 989 527
rect 1047 527 1053 528
rect 988 524 1018 526
rect 988 523 989 524
rect 983 522 989 523
rect 894 517 900 518
rect 894 513 895 517
rect 899 513 900 517
rect 894 512 900 513
rect 966 517 972 518
rect 966 513 967 517
rect 971 513 972 517
rect 966 512 972 513
rect 852 508 886 510
rect 910 511 917 512
rect 852 507 853 508
rect 847 506 853 507
rect 910 507 911 511
rect 916 507 917 511
rect 910 506 917 507
rect 951 511 957 512
rect 951 507 952 511
rect 956 510 957 511
rect 983 511 989 512
rect 983 510 984 511
rect 956 508 984 510
rect 956 507 957 508
rect 951 506 957 507
rect 983 507 984 508
rect 988 507 989 511
rect 1016 510 1018 524
rect 1047 523 1048 527
rect 1052 526 1053 527
rect 1080 526 1082 540
rect 1094 535 1100 536
rect 1094 531 1095 535
rect 1099 531 1100 535
rect 1094 530 1100 531
rect 1166 535 1172 536
rect 1166 531 1167 535
rect 1171 531 1172 535
rect 1166 530 1172 531
rect 1238 535 1244 536
rect 1238 531 1239 535
rect 1243 531 1244 535
rect 1238 530 1244 531
rect 1310 535 1316 536
rect 1310 531 1311 535
rect 1315 531 1316 535
rect 1310 530 1316 531
rect 1390 535 1396 536
rect 1390 531 1391 535
rect 1395 531 1396 535
rect 1390 530 1396 531
rect 1478 535 1484 536
rect 1478 531 1479 535
rect 1483 531 1484 535
rect 1478 530 1484 531
rect 1542 535 1548 536
rect 1542 531 1543 535
rect 1547 531 1548 535
rect 1542 530 1548 531
rect 1582 533 1588 534
rect 1582 529 1583 533
rect 1587 529 1588 533
rect 1582 528 1588 529
rect 1111 527 1117 528
rect 1111 526 1112 527
rect 1052 524 1078 526
rect 1080 524 1112 526
rect 1052 523 1053 524
rect 1047 522 1053 523
rect 1030 517 1036 518
rect 1030 513 1031 517
rect 1035 513 1036 517
rect 1030 512 1036 513
rect 1047 511 1053 512
rect 1047 510 1048 511
rect 1016 508 1048 510
rect 983 506 989 507
rect 1047 507 1048 508
rect 1052 507 1053 511
rect 1076 510 1078 524
rect 1111 523 1112 524
rect 1116 523 1117 527
rect 1111 522 1117 523
rect 1183 527 1189 528
rect 1183 523 1184 527
rect 1188 526 1189 527
rect 1255 527 1261 528
rect 1188 524 1222 526
rect 1188 523 1189 524
rect 1183 522 1189 523
rect 1094 517 1100 518
rect 1094 513 1095 517
rect 1099 513 1100 517
rect 1094 512 1100 513
rect 1166 517 1172 518
rect 1166 513 1167 517
rect 1171 513 1172 517
rect 1166 512 1172 513
rect 1111 511 1117 512
rect 1111 510 1112 511
rect 1076 508 1112 510
rect 1047 506 1053 507
rect 1111 507 1112 508
rect 1116 507 1117 511
rect 1111 506 1117 507
rect 1183 511 1189 512
rect 1183 507 1184 511
rect 1188 510 1189 511
rect 1191 511 1197 512
rect 1191 510 1192 511
rect 1188 508 1192 510
rect 1188 507 1189 508
rect 1183 506 1189 507
rect 1191 507 1192 508
rect 1196 507 1197 511
rect 1220 510 1222 524
rect 1255 523 1256 527
rect 1260 526 1261 527
rect 1327 527 1333 528
rect 1260 524 1294 526
rect 1260 523 1261 524
rect 1255 522 1261 523
rect 1238 517 1244 518
rect 1238 513 1239 517
rect 1243 513 1244 517
rect 1238 512 1244 513
rect 1255 511 1261 512
rect 1255 510 1256 511
rect 1220 508 1256 510
rect 1191 506 1197 507
rect 1255 507 1256 508
rect 1260 507 1261 511
rect 1292 510 1294 524
rect 1327 523 1328 527
rect 1332 526 1333 527
rect 1407 527 1413 528
rect 1332 524 1370 526
rect 1332 523 1333 524
rect 1327 522 1333 523
rect 1310 517 1316 518
rect 1310 513 1311 517
rect 1315 513 1316 517
rect 1310 512 1316 513
rect 1327 511 1333 512
rect 1327 510 1328 511
rect 1292 508 1328 510
rect 1255 506 1261 507
rect 1327 507 1328 508
rect 1332 507 1333 511
rect 1368 510 1370 524
rect 1407 523 1408 527
rect 1412 526 1413 527
rect 1471 527 1477 528
rect 1412 524 1461 526
rect 1412 523 1413 524
rect 1407 522 1413 523
rect 1390 517 1396 518
rect 1390 513 1391 517
rect 1395 513 1396 517
rect 1390 512 1396 513
rect 1407 511 1413 512
rect 1407 510 1408 511
rect 1368 508 1408 510
rect 1327 506 1333 507
rect 1407 507 1408 508
rect 1412 507 1413 511
rect 1459 510 1461 524
rect 1471 523 1472 527
rect 1476 526 1477 527
rect 1495 527 1501 528
rect 1495 526 1496 527
rect 1476 524 1496 526
rect 1476 523 1477 524
rect 1471 522 1477 523
rect 1495 523 1496 524
rect 1500 523 1501 527
rect 1495 522 1501 523
rect 1559 527 1565 528
rect 1559 523 1560 527
rect 1564 526 1565 527
rect 1567 527 1573 528
rect 1567 526 1568 527
rect 1564 524 1568 526
rect 1564 523 1565 524
rect 1559 522 1565 523
rect 1567 523 1568 524
rect 1572 523 1573 527
rect 1567 522 1573 523
rect 1478 517 1484 518
rect 1478 513 1479 517
rect 1483 513 1484 517
rect 1478 512 1484 513
rect 1542 517 1548 518
rect 1542 513 1543 517
rect 1547 513 1548 517
rect 1542 512 1548 513
rect 1582 516 1588 517
rect 1582 512 1583 516
rect 1587 512 1588 516
rect 1495 511 1501 512
rect 1495 510 1496 511
rect 1459 508 1496 510
rect 1407 506 1413 507
rect 1495 507 1496 508
rect 1500 507 1501 511
rect 1495 506 1501 507
rect 1558 511 1565 512
rect 1582 511 1588 512
rect 1558 507 1559 511
rect 1564 507 1565 511
rect 1558 506 1565 507
rect 694 502 700 503
rect 1498 503 1504 504
rect 664 500 690 502
rect 150 499 157 500
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 110 491 116 492
rect 134 495 140 496
rect 134 491 135 495
rect 139 491 140 495
rect 150 495 151 499
rect 156 495 157 499
rect 183 499 189 500
rect 183 498 184 499
rect 176 496 184 498
rect 150 494 157 495
rect 166 495 172 496
rect 134 490 140 491
rect 166 491 167 495
rect 171 491 172 495
rect 166 490 172 491
rect 176 486 178 496
rect 183 495 184 496
rect 188 495 189 499
rect 215 499 221 500
rect 215 498 216 499
rect 208 496 216 498
rect 183 494 189 495
rect 198 495 204 496
rect 198 491 199 495
rect 203 491 204 495
rect 198 490 204 491
rect 208 486 210 496
rect 215 495 216 496
rect 220 495 221 499
rect 263 499 269 500
rect 263 498 264 499
rect 259 496 264 498
rect 215 494 221 495
rect 246 495 252 496
rect 246 491 247 495
rect 251 491 252 495
rect 246 490 252 491
rect 259 486 261 496
rect 263 495 264 496
rect 268 495 269 499
rect 311 499 317 500
rect 263 494 269 495
rect 294 495 300 496
rect 294 491 295 495
rect 299 491 300 495
rect 311 495 312 499
rect 316 498 317 499
rect 326 499 332 500
rect 326 498 327 499
rect 316 496 327 498
rect 316 495 317 496
rect 311 494 317 495
rect 326 495 327 496
rect 331 495 332 499
rect 359 499 365 500
rect 359 498 360 499
rect 352 496 360 498
rect 326 494 332 495
rect 342 495 348 496
rect 294 490 300 491
rect 342 491 343 495
rect 347 491 348 495
rect 342 490 348 491
rect 352 486 354 496
rect 359 495 360 496
rect 364 495 365 499
rect 415 499 421 500
rect 359 494 365 495
rect 398 495 404 496
rect 398 491 399 495
rect 403 491 404 495
rect 415 495 416 499
rect 420 498 421 499
rect 438 499 444 500
rect 438 498 439 499
rect 420 496 439 498
rect 420 495 421 496
rect 415 494 421 495
rect 438 495 439 496
rect 443 495 444 499
rect 471 499 477 500
rect 471 498 472 499
rect 464 496 472 498
rect 438 494 444 495
rect 454 495 460 496
rect 398 490 404 491
rect 454 491 455 495
rect 459 491 460 495
rect 454 490 460 491
rect 464 486 466 496
rect 471 495 472 496
rect 476 495 477 499
rect 527 499 533 500
rect 527 498 528 499
rect 520 496 528 498
rect 471 494 477 495
rect 510 495 516 496
rect 510 491 511 495
rect 515 491 516 495
rect 510 490 516 491
rect 520 486 522 496
rect 527 495 528 496
rect 532 495 533 499
rect 583 499 589 500
rect 583 498 584 499
rect 576 496 584 498
rect 527 494 533 495
rect 566 495 572 496
rect 566 491 567 495
rect 571 491 572 495
rect 566 490 572 491
rect 576 486 578 496
rect 583 495 584 496
rect 588 495 589 499
rect 639 499 645 500
rect 639 498 640 499
rect 632 496 640 498
rect 583 494 589 495
rect 622 495 628 496
rect 622 491 623 495
rect 627 491 628 495
rect 622 490 628 491
rect 632 486 634 496
rect 639 495 640 496
rect 644 495 645 499
rect 695 499 701 500
rect 695 498 696 499
rect 688 496 696 498
rect 639 494 645 495
rect 678 495 684 496
rect 678 491 679 495
rect 683 491 684 495
rect 678 490 684 491
rect 688 486 690 496
rect 695 495 696 496
rect 700 495 701 499
rect 759 499 765 500
rect 695 494 701 495
rect 742 495 748 496
rect 742 491 743 495
rect 747 491 748 495
rect 759 495 760 499
rect 764 498 765 499
rect 791 499 797 500
rect 791 498 792 499
rect 764 496 792 498
rect 764 495 765 496
rect 759 494 765 495
rect 791 495 792 496
rect 796 495 797 499
rect 831 499 837 500
rect 831 498 832 499
rect 824 496 832 498
rect 791 494 797 495
rect 814 495 820 496
rect 742 490 748 491
rect 814 491 815 495
rect 819 491 820 495
rect 814 490 820 491
rect 824 486 826 496
rect 831 495 832 496
rect 836 495 837 499
rect 903 499 909 500
rect 903 498 904 499
rect 896 496 904 498
rect 831 494 837 495
rect 886 495 892 496
rect 886 491 887 495
rect 891 491 892 495
rect 886 490 892 491
rect 896 486 898 496
rect 903 495 904 496
rect 908 495 909 499
rect 975 499 981 500
rect 975 498 976 499
rect 968 496 976 498
rect 903 494 909 495
rect 958 495 964 496
rect 958 491 959 495
rect 963 491 964 495
rect 958 490 964 491
rect 968 486 970 496
rect 975 495 976 496
rect 980 495 981 499
rect 1055 499 1061 500
rect 1055 498 1056 499
rect 1048 496 1056 498
rect 975 494 981 495
rect 1038 495 1044 496
rect 1038 491 1039 495
rect 1043 491 1044 495
rect 1038 490 1044 491
rect 1048 486 1050 496
rect 1055 495 1056 496
rect 1060 495 1061 499
rect 1143 499 1149 500
rect 1055 494 1061 495
rect 1126 495 1132 496
rect 1126 491 1127 495
rect 1131 491 1132 495
rect 1143 495 1144 499
rect 1148 498 1149 499
rect 1214 499 1220 500
rect 1214 498 1215 499
rect 1148 496 1215 498
rect 1148 495 1149 496
rect 1143 494 1149 495
rect 1214 495 1215 496
rect 1219 495 1220 499
rect 1239 499 1245 500
rect 1239 498 1240 499
rect 1232 496 1240 498
rect 1214 494 1220 495
rect 1222 495 1228 496
rect 1126 490 1132 491
rect 1222 491 1223 495
rect 1227 491 1228 495
rect 1222 490 1228 491
rect 1232 486 1234 496
rect 1239 495 1240 496
rect 1244 495 1245 499
rect 1343 499 1349 500
rect 1239 494 1245 495
rect 1326 495 1332 496
rect 1326 491 1327 495
rect 1331 491 1332 495
rect 1343 495 1344 499
rect 1348 498 1349 499
rect 1455 499 1461 500
rect 1348 496 1410 498
rect 1348 495 1349 496
rect 1343 494 1349 495
rect 1326 490 1332 491
rect 164 484 178 486
rect 196 484 210 486
rect 236 484 261 486
rect 313 484 354 486
rect 444 484 466 486
rect 473 484 522 486
rect 556 484 578 486
rect 612 484 634 486
rect 668 484 690 486
rect 796 484 826 486
rect 868 484 898 486
rect 940 484 970 486
rect 1016 484 1050 486
rect 1192 484 1234 486
rect 1408 486 1410 496
rect 1438 495 1444 496
rect 1438 491 1439 495
rect 1443 491 1444 495
rect 1455 495 1456 499
rect 1460 498 1461 499
rect 1471 499 1477 500
rect 1471 498 1472 499
rect 1460 496 1472 498
rect 1460 495 1461 496
rect 1455 494 1461 495
rect 1471 495 1472 496
rect 1476 495 1477 499
rect 1498 499 1499 503
rect 1503 502 1504 503
rect 1503 500 1554 502
rect 1503 499 1504 500
rect 1498 498 1504 499
rect 1552 498 1554 500
rect 1559 499 1565 500
rect 1559 498 1560 499
rect 1552 496 1560 498
rect 1471 494 1477 495
rect 1542 495 1548 496
rect 1438 490 1444 491
rect 1542 491 1543 495
rect 1547 491 1548 495
rect 1559 495 1560 496
rect 1564 495 1565 499
rect 1559 494 1565 495
rect 1582 496 1588 497
rect 1582 492 1583 496
rect 1587 492 1588 496
rect 1582 491 1588 492
rect 1542 490 1548 491
rect 1408 484 1450 486
rect 151 483 157 484
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 151 479 152 483
rect 156 482 157 483
rect 164 482 166 484
rect 156 480 166 482
rect 183 483 189 484
rect 156 479 157 480
rect 151 478 157 479
rect 183 479 184 483
rect 188 482 189 483
rect 196 482 198 484
rect 188 480 198 482
rect 215 483 221 484
rect 188 479 189 480
rect 183 478 189 479
rect 215 479 216 483
rect 220 482 221 483
rect 236 482 238 484
rect 220 480 238 482
rect 263 483 272 484
rect 220 479 221 480
rect 215 478 221 479
rect 263 479 264 483
rect 271 479 272 483
rect 263 478 272 479
rect 311 483 317 484
rect 311 479 312 483
rect 316 479 317 483
rect 311 478 317 479
rect 359 483 365 484
rect 359 479 360 483
rect 364 479 365 483
rect 359 478 365 479
rect 415 483 421 484
rect 415 479 416 483
rect 420 482 421 483
rect 444 482 446 484
rect 420 480 446 482
rect 471 483 477 484
rect 420 479 421 480
rect 415 478 421 479
rect 471 479 472 483
rect 476 479 477 483
rect 471 478 477 479
rect 527 483 533 484
rect 527 479 528 483
rect 532 482 533 483
rect 556 482 558 484
rect 532 480 558 482
rect 583 483 589 484
rect 532 479 533 480
rect 527 478 533 479
rect 583 479 584 483
rect 588 482 589 483
rect 612 482 614 484
rect 588 480 614 482
rect 639 483 645 484
rect 588 479 589 480
rect 583 478 589 479
rect 639 479 640 483
rect 644 482 645 483
rect 668 482 670 484
rect 644 480 670 482
rect 694 483 701 484
rect 644 479 645 480
rect 639 478 645 479
rect 694 479 695 483
rect 700 479 701 483
rect 694 478 701 479
rect 759 483 765 484
rect 759 479 760 483
rect 764 482 765 483
rect 796 482 798 484
rect 764 480 798 482
rect 831 483 837 484
rect 764 479 765 480
rect 759 478 765 479
rect 831 479 832 483
rect 836 482 837 483
rect 868 482 870 484
rect 836 480 870 482
rect 903 483 909 484
rect 836 479 837 480
rect 831 478 837 479
rect 903 479 904 483
rect 908 482 909 483
rect 940 482 942 484
rect 908 480 942 482
rect 975 483 981 484
rect 908 479 909 480
rect 903 478 909 479
rect 975 479 976 483
rect 980 482 981 483
rect 1016 482 1018 484
rect 980 480 1018 482
rect 1055 483 1061 484
rect 980 479 981 480
rect 975 478 981 479
rect 1055 479 1056 483
rect 1060 479 1061 483
rect 1055 478 1061 479
rect 1143 483 1149 484
rect 1143 479 1144 483
rect 1148 482 1149 483
rect 1192 482 1194 484
rect 1148 480 1194 482
rect 1239 483 1245 484
rect 1148 479 1149 480
rect 1143 478 1149 479
rect 1239 479 1240 483
rect 1244 482 1245 483
rect 1278 483 1284 484
rect 1278 482 1279 483
rect 1244 480 1279 482
rect 1244 479 1245 480
rect 1239 478 1245 479
rect 1278 479 1279 480
rect 1283 479 1284 483
rect 1343 483 1349 484
rect 1343 482 1344 483
rect 1278 478 1284 479
rect 1336 480 1344 482
rect 110 474 116 475
rect 134 477 140 478
rect 134 473 135 477
rect 139 473 140 477
rect 134 472 140 473
rect 166 477 172 478
rect 166 473 167 477
rect 171 473 172 477
rect 166 472 172 473
rect 198 477 204 478
rect 198 473 199 477
rect 203 473 204 477
rect 198 472 204 473
rect 246 477 252 478
rect 246 473 247 477
rect 251 473 252 477
rect 246 472 252 473
rect 294 477 300 478
rect 294 473 295 477
rect 299 473 300 477
rect 294 472 300 473
rect 342 477 348 478
rect 342 473 343 477
rect 347 473 348 477
rect 342 472 348 473
rect 398 477 404 478
rect 398 473 399 477
rect 403 473 404 477
rect 398 472 404 473
rect 454 477 460 478
rect 454 473 455 477
rect 459 473 460 477
rect 454 472 460 473
rect 510 477 516 478
rect 510 473 511 477
rect 515 473 516 477
rect 510 472 516 473
rect 566 477 572 478
rect 566 473 567 477
rect 571 473 572 477
rect 566 472 572 473
rect 622 477 628 478
rect 622 473 623 477
rect 627 473 628 477
rect 622 472 628 473
rect 678 477 684 478
rect 678 473 679 477
rect 683 473 684 477
rect 678 472 684 473
rect 742 477 748 478
rect 742 473 743 477
rect 747 473 748 477
rect 742 472 748 473
rect 814 477 820 478
rect 814 473 815 477
rect 819 473 820 477
rect 814 472 820 473
rect 886 477 892 478
rect 886 473 887 477
rect 891 473 892 477
rect 886 472 892 473
rect 958 477 964 478
rect 958 473 959 477
rect 963 473 964 477
rect 958 472 964 473
rect 1038 477 1044 478
rect 1038 473 1039 477
rect 1043 473 1044 477
rect 1038 472 1044 473
rect 554 471 560 472
rect 554 467 555 471
rect 559 470 560 471
rect 894 471 900 472
rect 559 468 755 470
rect 559 467 560 468
rect 554 466 560 467
rect 134 463 140 464
rect 110 461 116 462
rect 110 457 111 461
rect 115 457 116 461
rect 134 459 135 463
rect 139 459 140 463
rect 134 458 140 459
rect 166 463 172 464
rect 166 459 167 463
rect 171 459 172 463
rect 166 458 172 459
rect 198 463 204 464
rect 198 459 199 463
rect 203 459 204 463
rect 198 458 204 459
rect 254 463 260 464
rect 254 459 255 463
rect 259 459 260 463
rect 254 458 260 459
rect 310 463 316 464
rect 310 459 311 463
rect 315 459 316 463
rect 310 458 316 459
rect 366 463 372 464
rect 366 459 367 463
rect 371 459 372 463
rect 366 458 372 459
rect 422 463 428 464
rect 422 459 423 463
rect 427 459 428 463
rect 422 458 428 459
rect 478 463 484 464
rect 478 459 479 463
rect 483 459 484 463
rect 478 458 484 459
rect 534 463 540 464
rect 534 459 535 463
rect 539 459 540 463
rect 534 458 540 459
rect 598 463 604 464
rect 598 459 599 463
rect 603 459 604 463
rect 598 458 604 459
rect 662 463 668 464
rect 662 459 663 463
rect 667 459 668 463
rect 662 458 668 459
rect 734 463 740 464
rect 734 459 735 463
rect 739 459 740 463
rect 734 458 740 459
rect 110 456 116 457
rect 753 456 755 468
rect 894 467 895 471
rect 899 470 900 471
rect 1057 470 1059 478
rect 1126 477 1132 478
rect 1126 473 1127 477
rect 1131 473 1132 477
rect 1126 472 1132 473
rect 1222 477 1228 478
rect 1222 473 1223 477
rect 1227 473 1228 477
rect 1222 472 1228 473
rect 1326 477 1332 478
rect 1326 473 1327 477
rect 1331 473 1332 477
rect 1326 472 1332 473
rect 899 468 1059 470
rect 1214 471 1220 472
rect 899 467 900 468
rect 894 466 900 467
rect 1214 467 1215 471
rect 1219 470 1220 471
rect 1336 470 1338 480
rect 1343 479 1344 480
rect 1348 479 1349 483
rect 1448 482 1450 484
rect 1455 483 1461 484
rect 1455 482 1456 483
rect 1448 480 1456 482
rect 1343 478 1349 479
rect 1455 479 1456 480
rect 1460 479 1461 483
rect 1455 478 1461 479
rect 1554 483 1565 484
rect 1554 479 1555 483
rect 1559 479 1560 483
rect 1564 479 1565 483
rect 1554 478 1565 479
rect 1582 479 1588 480
rect 1438 477 1444 478
rect 1438 473 1439 477
rect 1443 473 1444 477
rect 1438 472 1444 473
rect 1542 477 1548 478
rect 1542 473 1543 477
rect 1547 473 1548 477
rect 1582 475 1583 479
rect 1587 475 1588 479
rect 1582 474 1588 475
rect 1542 472 1548 473
rect 1219 468 1338 470
rect 1219 467 1220 468
rect 1214 466 1220 467
rect 806 463 812 464
rect 806 459 807 463
rect 811 459 812 463
rect 806 458 812 459
rect 870 463 876 464
rect 870 459 871 463
rect 875 459 876 463
rect 870 458 876 459
rect 934 463 940 464
rect 934 459 935 463
rect 939 459 940 463
rect 934 458 940 459
rect 990 463 996 464
rect 990 459 991 463
rect 995 459 996 463
rect 990 458 996 459
rect 1046 463 1052 464
rect 1046 459 1047 463
rect 1051 459 1052 463
rect 1046 458 1052 459
rect 1094 463 1100 464
rect 1094 459 1095 463
rect 1099 459 1100 463
rect 1094 458 1100 459
rect 1142 463 1148 464
rect 1142 459 1143 463
rect 1147 459 1148 463
rect 1142 458 1148 459
rect 1198 463 1204 464
rect 1198 459 1199 463
rect 1203 459 1204 463
rect 1198 458 1204 459
rect 1262 463 1268 464
rect 1262 459 1263 463
rect 1267 459 1268 463
rect 1262 458 1268 459
rect 1326 463 1332 464
rect 1326 459 1327 463
rect 1331 459 1332 463
rect 1326 458 1332 459
rect 1398 463 1404 464
rect 1398 459 1399 463
rect 1403 459 1404 463
rect 1398 458 1404 459
rect 1478 463 1484 464
rect 1478 459 1479 463
rect 1483 459 1484 463
rect 1478 458 1484 459
rect 1542 463 1548 464
rect 1542 459 1543 463
rect 1547 459 1548 463
rect 1542 458 1548 459
rect 1582 461 1588 462
rect 1582 457 1583 461
rect 1587 457 1588 461
rect 1582 456 1588 457
rect 150 455 157 456
rect 150 451 151 455
rect 156 451 157 455
rect 183 455 189 456
rect 183 454 184 455
rect 150 450 157 451
rect 176 452 184 454
rect 134 445 140 446
rect 110 444 116 445
rect 110 440 111 444
rect 115 440 116 444
rect 134 441 135 445
rect 139 441 140 445
rect 134 440 140 441
rect 166 445 172 446
rect 166 441 167 445
rect 171 441 172 445
rect 166 440 172 441
rect 110 439 116 440
rect 151 439 157 440
rect 151 435 152 439
rect 156 438 157 439
rect 176 438 178 452
rect 183 451 184 452
rect 188 451 189 455
rect 215 455 221 456
rect 215 454 216 455
rect 183 450 189 451
rect 208 452 216 454
rect 198 445 204 446
rect 198 441 199 445
rect 203 441 204 445
rect 198 440 204 441
rect 156 436 178 438
rect 183 439 189 440
rect 156 435 157 436
rect 151 434 157 435
rect 183 435 184 439
rect 188 438 189 439
rect 208 438 210 452
rect 215 451 216 452
rect 220 451 221 455
rect 271 455 277 456
rect 271 454 272 455
rect 215 450 221 451
rect 240 452 272 454
rect 188 436 210 438
rect 215 439 221 440
rect 188 435 189 436
rect 183 434 189 435
rect 215 435 216 439
rect 220 438 221 439
rect 240 438 242 452
rect 271 451 272 452
rect 276 451 277 455
rect 271 450 277 451
rect 326 455 333 456
rect 326 451 327 455
rect 332 451 333 455
rect 383 455 389 456
rect 383 454 384 455
rect 326 450 333 451
rect 356 452 384 454
rect 254 445 260 446
rect 254 441 255 445
rect 259 441 260 445
rect 254 440 260 441
rect 310 445 316 446
rect 310 441 311 445
rect 315 441 316 445
rect 310 440 316 441
rect 220 436 242 438
rect 266 439 277 440
rect 220 435 221 436
rect 215 434 221 435
rect 266 435 267 439
rect 271 435 272 439
rect 276 435 277 439
rect 266 434 277 435
rect 327 439 333 440
rect 327 435 328 439
rect 332 438 333 439
rect 356 438 358 452
rect 383 451 384 452
rect 388 451 389 455
rect 383 450 389 451
rect 438 455 445 456
rect 438 451 439 455
rect 444 451 445 455
rect 495 455 501 456
rect 495 454 496 455
rect 438 450 445 451
rect 472 452 496 454
rect 366 445 372 446
rect 366 441 367 445
rect 371 441 372 445
rect 366 440 372 441
rect 422 445 428 446
rect 422 441 423 445
rect 427 441 428 445
rect 422 440 428 441
rect 332 436 358 438
rect 378 439 389 440
rect 332 435 333 436
rect 327 434 333 435
rect 378 435 379 439
rect 383 435 384 439
rect 388 435 389 439
rect 378 434 389 435
rect 439 439 445 440
rect 439 435 440 439
rect 444 438 445 439
rect 472 438 474 452
rect 495 451 496 452
rect 500 451 501 455
rect 551 455 557 456
rect 551 454 552 455
rect 495 450 501 451
rect 524 452 552 454
rect 478 445 484 446
rect 478 441 479 445
rect 483 441 484 445
rect 478 440 484 441
rect 444 436 474 438
rect 495 439 501 440
rect 444 435 445 436
rect 439 434 445 435
rect 495 435 496 439
rect 500 438 501 439
rect 524 438 526 452
rect 551 451 552 452
rect 556 451 557 455
rect 551 450 557 451
rect 615 455 621 456
rect 615 451 616 455
rect 620 454 621 455
rect 679 455 685 456
rect 620 452 650 454
rect 620 451 621 452
rect 615 450 621 451
rect 534 445 540 446
rect 534 441 535 445
rect 539 441 540 445
rect 534 440 540 441
rect 598 445 604 446
rect 598 441 599 445
rect 603 441 604 445
rect 598 440 604 441
rect 500 436 526 438
rect 551 439 560 440
rect 500 435 501 436
rect 495 434 501 435
rect 551 435 552 439
rect 559 435 560 439
rect 551 434 560 435
rect 562 439 568 440
rect 562 435 563 439
rect 567 438 568 439
rect 615 439 621 440
rect 615 438 616 439
rect 567 436 616 438
rect 567 435 568 436
rect 562 434 568 435
rect 615 435 616 436
rect 620 435 621 439
rect 648 438 650 452
rect 679 451 680 455
rect 684 454 685 455
rect 751 455 757 456
rect 684 452 746 454
rect 684 451 685 452
rect 679 450 685 451
rect 662 445 668 446
rect 662 441 663 445
rect 667 441 668 445
rect 662 440 668 441
rect 734 445 740 446
rect 734 441 735 445
rect 739 441 740 445
rect 734 440 740 441
rect 679 439 685 440
rect 679 438 680 439
rect 648 436 680 438
rect 615 434 621 435
rect 679 435 680 436
rect 684 435 685 439
rect 744 438 746 452
rect 751 451 752 455
rect 756 451 757 455
rect 751 450 757 451
rect 778 455 784 456
rect 778 451 779 455
rect 783 454 784 455
rect 823 455 829 456
rect 823 454 824 455
rect 783 452 824 454
rect 783 451 784 452
rect 778 450 784 451
rect 823 451 824 452
rect 828 451 829 455
rect 887 455 893 456
rect 887 454 888 455
rect 823 450 829 451
rect 860 452 888 454
rect 806 445 812 446
rect 806 441 807 445
rect 811 441 812 445
rect 806 440 812 441
rect 751 439 757 440
rect 751 438 752 439
rect 744 436 752 438
rect 679 434 685 435
rect 751 435 752 436
rect 756 435 757 439
rect 751 434 757 435
rect 823 439 829 440
rect 823 435 824 439
rect 828 438 829 439
rect 860 438 862 452
rect 887 451 888 452
rect 892 451 893 455
rect 887 450 893 451
rect 951 455 957 456
rect 951 451 952 455
rect 956 454 957 455
rect 1007 455 1013 456
rect 956 452 982 454
rect 956 451 957 452
rect 951 450 957 451
rect 870 445 876 446
rect 870 441 871 445
rect 875 441 876 445
rect 870 440 876 441
rect 934 445 940 446
rect 934 441 935 445
rect 939 441 940 445
rect 934 440 940 441
rect 828 436 862 438
rect 887 439 893 440
rect 828 435 829 436
rect 823 434 829 435
rect 887 435 888 439
rect 892 435 893 439
rect 887 434 893 435
rect 951 439 957 440
rect 951 435 952 439
rect 956 438 957 439
rect 980 438 982 452
rect 1007 451 1008 455
rect 1012 454 1013 455
rect 1038 455 1044 456
rect 1038 454 1039 455
rect 1012 452 1039 454
rect 1012 451 1013 452
rect 1007 450 1013 451
rect 1038 451 1039 452
rect 1043 451 1044 455
rect 1063 455 1069 456
rect 1063 454 1064 455
rect 1038 450 1044 451
rect 1056 452 1064 454
rect 990 445 996 446
rect 990 441 991 445
rect 995 441 996 445
rect 990 440 996 441
rect 1046 445 1052 446
rect 1046 441 1047 445
rect 1051 441 1052 445
rect 1046 440 1052 441
rect 1007 439 1013 440
rect 1007 438 1008 439
rect 956 436 978 438
rect 980 436 1008 438
rect 956 435 957 436
rect 951 434 957 435
rect 606 431 612 432
rect 606 430 607 431
rect 537 428 607 430
rect 150 423 157 424
rect 110 420 116 421
rect 110 416 111 420
rect 115 416 116 420
rect 110 415 116 416
rect 134 419 140 420
rect 134 415 135 419
rect 139 415 140 419
rect 150 419 151 423
rect 156 419 157 423
rect 183 423 189 424
rect 183 422 184 423
rect 176 420 184 422
rect 150 418 157 419
rect 166 419 172 420
rect 134 414 140 415
rect 166 415 167 419
rect 171 415 172 419
rect 166 414 172 415
rect 176 410 178 420
rect 183 419 184 420
rect 188 419 189 423
rect 247 423 253 424
rect 247 422 248 423
rect 240 420 248 422
rect 183 418 189 419
rect 230 419 236 420
rect 230 415 231 419
rect 235 415 236 419
rect 230 414 236 415
rect 240 410 242 420
rect 247 419 248 420
rect 252 419 253 423
rect 311 423 317 424
rect 311 422 312 423
rect 304 420 312 422
rect 247 418 253 419
rect 294 419 300 420
rect 294 415 295 419
rect 299 415 300 419
rect 294 414 300 415
rect 304 410 306 420
rect 311 419 312 420
rect 316 419 317 423
rect 375 423 381 424
rect 311 418 317 419
rect 358 419 364 420
rect 358 415 359 419
rect 363 415 364 419
rect 375 419 376 423
rect 380 419 381 423
rect 439 423 445 424
rect 375 418 381 419
rect 422 419 428 420
rect 358 414 364 415
rect 377 414 379 418
rect 422 415 423 419
rect 427 415 428 419
rect 439 419 440 423
rect 444 422 445 423
rect 455 423 461 424
rect 455 422 456 423
rect 444 420 456 422
rect 444 419 445 420
rect 439 418 445 419
rect 455 419 456 420
rect 460 419 461 423
rect 503 423 509 424
rect 455 418 461 419
rect 486 419 492 420
rect 422 414 428 415
rect 486 415 487 419
rect 491 415 492 419
rect 503 419 504 423
rect 508 422 509 423
rect 537 422 539 428
rect 606 427 607 428
rect 611 427 612 431
rect 976 430 978 436
rect 1007 435 1008 436
rect 1012 435 1013 439
rect 1056 438 1058 452
rect 1063 451 1064 452
rect 1068 451 1069 455
rect 1111 455 1117 456
rect 1111 454 1112 455
rect 1063 450 1069 451
rect 1084 452 1112 454
rect 1007 434 1013 435
rect 1016 436 1058 438
rect 1063 439 1069 440
rect 1016 430 1018 436
rect 1063 435 1064 439
rect 1068 438 1069 439
rect 1084 438 1086 452
rect 1111 451 1112 452
rect 1116 451 1117 455
rect 1159 455 1165 456
rect 1159 454 1160 455
rect 1111 450 1117 451
rect 1136 452 1160 454
rect 1094 445 1100 446
rect 1094 441 1095 445
rect 1099 441 1100 445
rect 1094 440 1100 441
rect 1068 436 1086 438
rect 1111 439 1117 440
rect 1068 435 1069 436
rect 1063 434 1069 435
rect 1111 435 1112 439
rect 1116 438 1117 439
rect 1136 438 1138 452
rect 1159 451 1160 452
rect 1164 451 1165 455
rect 1215 455 1221 456
rect 1215 454 1216 455
rect 1159 450 1165 451
rect 1188 452 1216 454
rect 1142 445 1148 446
rect 1142 441 1143 445
rect 1147 441 1148 445
rect 1142 440 1148 441
rect 1116 436 1138 438
rect 1159 439 1165 440
rect 1116 435 1117 436
rect 1111 434 1117 435
rect 1159 435 1160 439
rect 1164 438 1165 439
rect 1188 438 1190 452
rect 1215 451 1216 452
rect 1220 451 1221 455
rect 1215 450 1221 451
rect 1279 455 1285 456
rect 1279 451 1280 455
rect 1284 454 1285 455
rect 1343 455 1349 456
rect 1284 452 1314 454
rect 1284 451 1285 452
rect 1279 450 1285 451
rect 1198 445 1204 446
rect 1198 441 1199 445
rect 1203 441 1204 445
rect 1198 440 1204 441
rect 1262 445 1268 446
rect 1262 441 1263 445
rect 1267 441 1268 445
rect 1262 440 1268 441
rect 1164 436 1190 438
rect 1215 439 1221 440
rect 1164 435 1165 436
rect 1159 434 1165 435
rect 1215 435 1216 439
rect 1220 438 1221 439
rect 1278 439 1285 440
rect 1220 436 1274 438
rect 1220 435 1221 436
rect 1215 434 1221 435
rect 976 428 1018 430
rect 1272 430 1274 436
rect 1278 435 1279 439
rect 1284 435 1285 439
rect 1312 438 1314 452
rect 1343 451 1344 455
rect 1348 454 1349 455
rect 1390 455 1396 456
rect 1348 452 1382 454
rect 1348 451 1349 452
rect 1343 450 1349 451
rect 1326 445 1332 446
rect 1326 441 1327 445
rect 1331 441 1332 445
rect 1326 440 1332 441
rect 1343 439 1349 440
rect 1343 438 1344 439
rect 1312 436 1344 438
rect 1278 434 1285 435
rect 1343 435 1344 436
rect 1348 435 1349 439
rect 1380 438 1382 452
rect 1390 451 1391 455
rect 1395 454 1396 455
rect 1415 455 1421 456
rect 1415 454 1416 455
rect 1395 452 1416 454
rect 1395 451 1396 452
rect 1390 450 1396 451
rect 1415 451 1416 452
rect 1420 451 1421 455
rect 1415 450 1421 451
rect 1495 455 1504 456
rect 1495 451 1496 455
rect 1503 451 1504 455
rect 1495 450 1504 451
rect 1558 455 1565 456
rect 1558 451 1559 455
rect 1564 451 1565 455
rect 1558 450 1565 451
rect 1398 445 1404 446
rect 1398 441 1399 445
rect 1403 441 1404 445
rect 1398 440 1404 441
rect 1478 445 1484 446
rect 1478 441 1479 445
rect 1483 441 1484 445
rect 1478 440 1484 441
rect 1542 445 1548 446
rect 1542 441 1543 445
rect 1547 441 1548 445
rect 1542 440 1548 441
rect 1582 444 1588 445
rect 1582 440 1583 444
rect 1587 440 1588 444
rect 1415 439 1421 440
rect 1415 438 1416 439
rect 1380 436 1416 438
rect 1343 434 1349 435
rect 1415 435 1416 436
rect 1420 435 1421 439
rect 1415 434 1421 435
rect 1486 439 1492 440
rect 1486 435 1487 439
rect 1491 438 1492 439
rect 1495 439 1501 440
rect 1495 438 1496 439
rect 1491 436 1496 438
rect 1491 435 1492 436
rect 1486 434 1492 435
rect 1495 435 1496 436
rect 1500 435 1501 439
rect 1495 434 1501 435
rect 1559 439 1565 440
rect 1559 435 1560 439
rect 1564 438 1565 439
rect 1567 439 1573 440
rect 1582 439 1588 440
rect 1567 438 1568 439
rect 1564 436 1568 438
rect 1564 435 1565 436
rect 1559 434 1565 435
rect 1567 435 1568 436
rect 1572 435 1573 439
rect 1567 434 1573 435
rect 1390 431 1396 432
rect 1390 430 1391 431
rect 1272 428 1391 430
rect 606 426 612 427
rect 1038 427 1044 428
rect 559 423 565 424
rect 559 422 560 423
rect 508 420 539 422
rect 552 420 560 422
rect 508 419 509 420
rect 503 418 509 419
rect 542 419 548 420
rect 486 414 492 415
rect 542 415 543 419
rect 547 415 548 419
rect 542 414 548 415
rect 377 412 418 414
rect 164 408 178 410
rect 216 408 242 410
rect 259 408 306 410
rect 416 410 418 412
rect 552 410 554 420
rect 559 419 560 420
rect 564 419 565 423
rect 607 423 613 424
rect 559 418 565 419
rect 590 419 596 420
rect 590 415 591 419
rect 595 415 596 419
rect 607 419 608 423
rect 612 419 613 423
rect 655 423 661 424
rect 607 418 613 419
rect 638 419 644 420
rect 590 414 596 415
rect 609 414 611 418
rect 638 415 639 419
rect 643 415 644 419
rect 655 419 656 423
rect 660 422 661 423
rect 695 423 701 424
rect 660 420 675 422
rect 660 419 661 420
rect 655 418 661 419
rect 638 414 644 415
rect 609 412 634 414
rect 416 408 434 410
rect 532 408 554 410
rect 632 410 634 412
rect 673 410 675 420
rect 678 419 684 420
rect 678 415 679 419
rect 683 415 684 419
rect 695 419 696 423
rect 700 422 701 423
rect 735 423 741 424
rect 700 420 714 422
rect 700 419 701 420
rect 695 418 701 419
rect 678 414 684 415
rect 712 410 714 420
rect 718 419 724 420
rect 718 415 719 419
rect 723 415 724 419
rect 735 419 736 423
rect 740 422 741 423
rect 743 423 749 424
rect 743 422 744 423
rect 740 420 744 422
rect 740 419 741 420
rect 735 418 741 419
rect 743 419 744 420
rect 748 419 749 423
rect 775 423 784 424
rect 743 418 749 419
rect 758 419 764 420
rect 718 414 724 415
rect 758 415 759 419
rect 763 415 764 419
rect 775 419 776 423
rect 783 419 784 423
rect 823 423 829 424
rect 823 422 824 423
rect 816 420 824 422
rect 775 418 784 419
rect 806 419 812 420
rect 758 414 764 415
rect 806 415 807 419
rect 811 415 812 419
rect 806 414 812 415
rect 816 410 818 420
rect 823 419 824 420
rect 828 419 829 423
rect 879 423 885 424
rect 879 422 880 423
rect 872 420 880 422
rect 823 418 829 419
rect 862 419 868 420
rect 862 415 863 419
rect 867 415 868 419
rect 862 414 868 415
rect 872 410 874 420
rect 879 419 880 420
rect 884 419 885 423
rect 935 423 941 424
rect 935 422 936 423
rect 928 420 936 422
rect 879 418 885 419
rect 918 419 924 420
rect 918 415 919 419
rect 923 415 924 419
rect 918 414 924 415
rect 928 410 930 420
rect 935 419 936 420
rect 940 419 941 423
rect 991 423 997 424
rect 991 422 992 423
rect 984 420 992 422
rect 935 418 941 419
rect 974 419 980 420
rect 974 415 975 419
rect 979 415 980 419
rect 974 414 980 415
rect 984 410 986 420
rect 991 419 992 420
rect 996 419 997 423
rect 1038 423 1039 427
rect 1043 423 1044 427
rect 1390 427 1391 428
rect 1395 427 1396 431
rect 1390 426 1396 427
rect 1038 422 1044 423
rect 1047 423 1053 424
rect 1047 422 1048 423
rect 1040 420 1048 422
rect 991 418 997 419
rect 1030 419 1036 420
rect 1030 415 1031 419
rect 1035 415 1036 419
rect 1047 419 1048 420
rect 1052 419 1053 423
rect 1103 423 1109 424
rect 1103 422 1104 423
rect 1099 420 1104 422
rect 1047 418 1053 419
rect 1086 419 1092 420
rect 1030 414 1036 415
rect 1086 415 1087 419
rect 1091 415 1092 419
rect 1086 414 1092 415
rect 1099 410 1101 420
rect 1103 419 1104 420
rect 1108 419 1109 423
rect 1167 423 1173 424
rect 1167 422 1168 423
rect 1160 420 1168 422
rect 1103 418 1109 419
rect 1150 419 1156 420
rect 1150 415 1151 419
rect 1155 415 1156 419
rect 1150 414 1156 415
rect 1160 410 1162 420
rect 1167 419 1168 420
rect 1172 419 1173 423
rect 1239 423 1245 424
rect 1239 422 1240 423
rect 1232 420 1240 422
rect 1167 418 1173 419
rect 1222 419 1228 420
rect 1222 415 1223 419
rect 1227 415 1228 419
rect 1222 414 1228 415
rect 1232 410 1234 420
rect 1239 419 1240 420
rect 1244 419 1245 423
rect 1319 423 1325 424
rect 1319 422 1320 423
rect 1312 420 1320 422
rect 1239 418 1245 419
rect 1302 419 1308 420
rect 1302 415 1303 419
rect 1307 415 1308 419
rect 1302 414 1308 415
rect 1312 410 1314 420
rect 1319 419 1320 420
rect 1324 419 1325 423
rect 1399 423 1405 424
rect 1399 422 1400 423
rect 1392 420 1400 422
rect 1319 418 1325 419
rect 1382 419 1388 420
rect 1382 415 1383 419
rect 1387 415 1388 419
rect 1382 414 1388 415
rect 1392 410 1394 420
rect 1399 419 1400 420
rect 1404 419 1405 423
rect 1487 423 1493 424
rect 1399 418 1405 419
rect 1470 419 1476 420
rect 1470 415 1471 419
rect 1475 415 1476 419
rect 1487 419 1488 423
rect 1492 422 1493 423
rect 1502 423 1508 424
rect 1502 422 1503 423
rect 1492 420 1503 422
rect 1492 419 1493 420
rect 1487 418 1493 419
rect 1502 419 1503 420
rect 1507 419 1508 423
rect 1558 423 1565 424
rect 1502 418 1508 419
rect 1542 419 1548 420
rect 1470 414 1476 415
rect 1542 415 1543 419
rect 1547 415 1548 419
rect 1558 419 1559 423
rect 1564 419 1565 423
rect 1558 418 1565 419
rect 1582 420 1588 421
rect 1582 416 1583 420
rect 1587 416 1588 420
rect 1582 415 1588 416
rect 1542 414 1548 415
rect 632 408 650 410
rect 673 408 690 410
rect 712 408 739 410
rect 800 408 818 410
rect 825 408 874 410
rect 908 408 930 410
rect 937 408 986 410
rect 1072 408 1101 410
rect 1136 408 1162 410
rect 1204 408 1234 410
rect 1280 408 1314 410
rect 1321 408 1394 410
rect 151 407 157 408
rect 110 403 116 404
rect 110 399 111 403
rect 115 399 116 403
rect 151 403 152 407
rect 156 406 157 407
rect 164 406 166 408
rect 156 404 166 406
rect 183 407 189 408
rect 156 403 157 404
rect 151 402 157 403
rect 183 403 184 407
rect 188 406 189 407
rect 216 406 218 408
rect 188 404 218 406
rect 247 407 253 408
rect 188 403 189 404
rect 183 402 189 403
rect 247 403 248 407
rect 252 406 253 407
rect 259 406 261 408
rect 252 404 261 406
rect 310 407 317 408
rect 252 403 253 404
rect 247 402 253 403
rect 310 403 311 407
rect 316 403 317 407
rect 310 402 317 403
rect 375 407 384 408
rect 375 403 376 407
rect 383 403 384 407
rect 432 406 434 408
rect 439 407 445 408
rect 439 406 440 407
rect 432 404 440 406
rect 375 402 384 403
rect 439 403 440 404
rect 444 403 445 407
rect 439 402 445 403
rect 503 407 509 408
rect 503 403 504 407
rect 508 406 509 407
rect 532 406 534 408
rect 508 404 534 406
rect 559 407 568 408
rect 508 403 509 404
rect 503 402 509 403
rect 559 403 560 407
rect 567 403 568 407
rect 559 402 568 403
rect 606 407 613 408
rect 606 403 607 407
rect 612 403 613 407
rect 648 406 650 408
rect 655 407 661 408
rect 655 406 656 407
rect 648 404 656 406
rect 606 402 613 403
rect 655 403 656 404
rect 660 403 661 407
rect 688 406 690 408
rect 695 407 701 408
rect 695 406 696 407
rect 688 404 696 406
rect 655 402 661 403
rect 695 403 696 404
rect 700 403 701 407
rect 695 402 701 403
rect 735 407 741 408
rect 735 403 736 407
rect 740 403 741 407
rect 735 402 741 403
rect 775 407 781 408
rect 775 403 776 407
rect 780 406 781 407
rect 800 406 802 408
rect 780 404 802 406
rect 823 407 829 408
rect 780 403 781 404
rect 775 402 781 403
rect 823 403 824 407
rect 828 403 829 407
rect 823 402 829 403
rect 879 407 885 408
rect 879 403 880 407
rect 884 406 885 407
rect 908 406 910 408
rect 884 404 910 406
rect 935 407 941 408
rect 884 403 885 404
rect 879 402 885 403
rect 935 403 936 407
rect 940 403 941 407
rect 991 407 997 408
rect 991 406 992 407
rect 935 402 941 403
rect 984 404 992 406
rect 110 398 116 399
rect 134 401 140 402
rect 134 397 135 401
rect 139 397 140 401
rect 134 396 140 397
rect 166 401 172 402
rect 166 397 167 401
rect 171 397 172 401
rect 166 396 172 397
rect 230 401 236 402
rect 230 397 231 401
rect 235 397 236 401
rect 230 396 236 397
rect 294 401 300 402
rect 294 397 295 401
rect 299 397 300 401
rect 294 396 300 397
rect 358 401 364 402
rect 358 397 359 401
rect 363 397 364 401
rect 358 396 364 397
rect 422 401 428 402
rect 422 397 423 401
rect 427 397 428 401
rect 422 396 428 397
rect 486 401 492 402
rect 486 397 487 401
rect 491 397 492 401
rect 486 396 492 397
rect 542 401 548 402
rect 542 397 543 401
rect 547 397 548 401
rect 542 396 548 397
rect 590 401 596 402
rect 590 397 591 401
rect 595 397 596 401
rect 590 396 596 397
rect 638 401 644 402
rect 638 397 639 401
rect 643 397 644 401
rect 638 396 644 397
rect 678 401 684 402
rect 678 397 679 401
rect 683 397 684 401
rect 678 396 684 397
rect 718 401 724 402
rect 718 397 719 401
rect 723 397 724 401
rect 718 396 724 397
rect 758 401 764 402
rect 758 397 759 401
rect 763 397 764 401
rect 758 396 764 397
rect 806 401 812 402
rect 806 397 807 401
rect 811 397 812 401
rect 806 396 812 397
rect 862 401 868 402
rect 862 397 863 401
rect 867 397 868 401
rect 862 396 868 397
rect 918 401 924 402
rect 918 397 919 401
rect 923 397 924 401
rect 918 396 924 397
rect 974 401 980 402
rect 974 397 975 401
rect 979 397 980 401
rect 974 396 980 397
rect 826 395 832 396
rect 826 391 827 395
rect 831 394 832 395
rect 984 394 986 404
rect 991 403 992 404
rect 996 403 997 407
rect 991 402 997 403
rect 1047 407 1053 408
rect 1047 403 1048 407
rect 1052 406 1053 407
rect 1072 406 1074 408
rect 1052 404 1074 406
rect 1103 407 1109 408
rect 1052 403 1053 404
rect 1047 402 1053 403
rect 1103 403 1104 407
rect 1108 406 1109 407
rect 1136 406 1138 408
rect 1108 404 1138 406
rect 1167 407 1173 408
rect 1108 403 1109 404
rect 1103 402 1109 403
rect 1167 403 1168 407
rect 1172 406 1173 407
rect 1204 406 1206 408
rect 1172 404 1206 406
rect 1239 407 1245 408
rect 1172 403 1173 404
rect 1167 402 1173 403
rect 1239 403 1240 407
rect 1244 406 1245 407
rect 1280 406 1282 408
rect 1244 404 1282 406
rect 1319 407 1325 408
rect 1244 403 1245 404
rect 1239 402 1245 403
rect 1319 403 1320 407
rect 1324 403 1325 407
rect 1399 407 1405 408
rect 1399 406 1400 407
rect 1319 402 1325 403
rect 1392 404 1400 406
rect 1030 401 1036 402
rect 1030 397 1031 401
rect 1035 397 1036 401
rect 1030 396 1036 397
rect 1086 401 1092 402
rect 1086 397 1087 401
rect 1091 397 1092 401
rect 1086 396 1092 397
rect 1150 401 1156 402
rect 1150 397 1151 401
rect 1155 397 1156 401
rect 1150 396 1156 397
rect 1222 401 1228 402
rect 1222 397 1223 401
rect 1227 397 1228 401
rect 1222 396 1228 397
rect 1302 401 1308 402
rect 1302 397 1303 401
rect 1307 397 1308 401
rect 1302 396 1308 397
rect 1382 401 1388 402
rect 1382 397 1383 401
rect 1387 397 1388 401
rect 1382 396 1388 397
rect 831 392 986 394
rect 1158 395 1164 396
rect 831 391 832 392
rect 826 390 832 391
rect 1158 391 1159 395
rect 1163 394 1164 395
rect 1392 394 1394 404
rect 1399 403 1400 404
rect 1404 403 1405 407
rect 1399 402 1405 403
rect 1486 407 1493 408
rect 1486 403 1487 407
rect 1492 403 1493 407
rect 1486 402 1493 403
rect 1558 407 1565 408
rect 1558 403 1559 407
rect 1564 403 1565 407
rect 1558 402 1565 403
rect 1582 403 1588 404
rect 1470 401 1476 402
rect 1470 397 1471 401
rect 1475 397 1476 401
rect 1470 396 1476 397
rect 1542 401 1548 402
rect 1542 397 1543 401
rect 1547 397 1548 401
rect 1582 399 1583 403
rect 1587 399 1588 403
rect 1582 398 1588 399
rect 1542 396 1548 397
rect 1163 392 1394 394
rect 1163 391 1164 392
rect 1158 390 1164 391
rect 134 387 140 388
rect 110 385 116 386
rect 110 381 111 385
rect 115 381 116 385
rect 134 383 135 387
rect 139 383 140 387
rect 134 382 140 383
rect 206 387 212 388
rect 206 383 207 387
rect 211 383 212 387
rect 206 382 212 383
rect 294 387 300 388
rect 294 383 295 387
rect 299 383 300 387
rect 294 382 300 383
rect 382 387 388 388
rect 382 383 383 387
rect 387 383 388 387
rect 382 382 388 383
rect 462 387 468 388
rect 462 383 463 387
rect 467 383 468 387
rect 462 382 468 383
rect 534 387 540 388
rect 534 383 535 387
rect 539 383 540 387
rect 534 382 540 383
rect 598 387 604 388
rect 598 383 599 387
rect 603 383 604 387
rect 598 382 604 383
rect 654 387 660 388
rect 654 383 655 387
rect 659 383 660 387
rect 654 382 660 383
rect 702 387 708 388
rect 702 383 703 387
rect 707 383 708 387
rect 702 382 708 383
rect 750 387 756 388
rect 750 383 751 387
rect 755 383 756 387
rect 750 382 756 383
rect 806 387 812 388
rect 806 383 807 387
rect 811 383 812 387
rect 806 382 812 383
rect 862 387 868 388
rect 862 383 863 387
rect 867 383 868 387
rect 862 382 868 383
rect 918 387 924 388
rect 918 383 919 387
rect 923 383 924 387
rect 918 382 924 383
rect 982 387 988 388
rect 982 383 983 387
rect 987 383 988 387
rect 982 382 988 383
rect 1054 387 1060 388
rect 1054 383 1055 387
rect 1059 383 1060 387
rect 1054 382 1060 383
rect 1126 387 1132 388
rect 1126 383 1127 387
rect 1131 383 1132 387
rect 1126 382 1132 383
rect 1198 387 1204 388
rect 1198 383 1199 387
rect 1203 383 1204 387
rect 1198 382 1204 383
rect 1270 387 1276 388
rect 1270 383 1271 387
rect 1275 383 1276 387
rect 1270 382 1276 383
rect 1342 387 1348 388
rect 1342 383 1343 387
rect 1347 383 1348 387
rect 1342 382 1348 383
rect 1414 387 1420 388
rect 1414 383 1415 387
rect 1419 383 1420 387
rect 1414 382 1420 383
rect 1486 387 1492 388
rect 1486 383 1487 387
rect 1491 383 1492 387
rect 1486 382 1492 383
rect 1542 387 1548 388
rect 1542 383 1543 387
rect 1547 383 1548 387
rect 1542 382 1548 383
rect 1582 385 1588 386
rect 110 380 116 381
rect 1582 381 1583 385
rect 1587 381 1588 385
rect 1582 380 1588 381
rect 150 379 157 380
rect 150 375 151 379
rect 156 375 157 379
rect 223 379 229 380
rect 223 378 224 379
rect 150 374 157 375
rect 192 376 224 378
rect 134 369 140 370
rect 110 368 116 369
rect 110 364 111 368
rect 115 364 116 368
rect 134 365 135 369
rect 139 365 140 369
rect 134 364 140 365
rect 110 363 116 364
rect 151 363 157 364
rect 151 359 152 363
rect 156 362 157 363
rect 192 362 194 376
rect 223 375 224 376
rect 228 375 229 379
rect 223 374 229 375
rect 311 379 317 380
rect 311 375 312 379
rect 316 378 317 379
rect 399 379 405 380
rect 316 376 394 378
rect 316 375 317 376
rect 311 374 317 375
rect 310 371 316 372
rect 310 370 311 371
rect 206 369 212 370
rect 206 365 207 369
rect 211 365 212 369
rect 206 364 212 365
rect 294 369 300 370
rect 294 365 295 369
rect 299 365 300 369
rect 294 364 300 365
rect 304 368 311 370
rect 156 360 194 362
rect 223 363 229 364
rect 156 359 157 360
rect 151 358 157 359
rect 223 359 224 363
rect 228 362 229 363
rect 304 362 306 368
rect 310 367 311 368
rect 315 367 316 371
rect 310 366 316 367
rect 382 369 388 370
rect 382 365 383 369
rect 387 365 388 369
rect 382 364 388 365
rect 228 360 306 362
rect 311 363 317 364
rect 228 359 229 360
rect 223 358 229 359
rect 311 359 312 363
rect 316 362 317 363
rect 350 363 356 364
rect 350 362 351 363
rect 316 360 351 362
rect 316 359 317 360
rect 311 358 317 359
rect 350 359 351 360
rect 355 359 356 363
rect 392 362 394 376
rect 399 375 400 379
rect 404 378 405 379
rect 455 379 461 380
rect 404 376 442 378
rect 404 375 405 376
rect 399 374 405 375
rect 399 363 405 364
rect 399 362 400 363
rect 392 360 400 362
rect 350 358 356 359
rect 399 359 400 360
rect 404 359 405 363
rect 440 362 442 376
rect 455 375 456 379
rect 460 378 461 379
rect 479 379 485 380
rect 479 378 480 379
rect 460 376 480 378
rect 460 375 461 376
rect 455 374 461 375
rect 479 375 480 376
rect 484 375 485 379
rect 479 374 485 375
rect 551 379 557 380
rect 551 375 552 379
rect 556 378 557 379
rect 615 379 621 380
rect 556 376 586 378
rect 556 375 557 376
rect 551 374 557 375
rect 462 369 468 370
rect 462 365 463 369
rect 467 365 468 369
rect 462 364 468 365
rect 534 369 540 370
rect 534 365 535 369
rect 539 365 540 369
rect 534 364 540 365
rect 479 363 485 364
rect 479 362 480 363
rect 440 360 480 362
rect 399 358 405 359
rect 479 359 480 360
rect 484 359 485 363
rect 479 358 485 359
rect 551 363 557 364
rect 551 359 552 363
rect 556 362 557 363
rect 574 363 580 364
rect 574 362 575 363
rect 556 360 575 362
rect 556 359 557 360
rect 551 358 557 359
rect 574 359 575 360
rect 579 359 580 363
rect 584 362 586 376
rect 615 375 616 379
rect 620 378 621 379
rect 671 379 677 380
rect 620 376 646 378
rect 620 375 621 376
rect 615 374 621 375
rect 598 369 604 370
rect 598 365 599 369
rect 603 365 604 369
rect 598 364 604 365
rect 615 363 621 364
rect 615 362 616 363
rect 584 360 616 362
rect 574 358 580 359
rect 615 359 616 360
rect 620 359 621 363
rect 644 362 646 376
rect 671 375 672 379
rect 676 378 677 379
rect 719 379 725 380
rect 676 376 714 378
rect 676 375 677 376
rect 671 374 677 375
rect 654 369 660 370
rect 654 365 655 369
rect 659 365 660 369
rect 654 364 660 365
rect 702 369 708 370
rect 702 365 703 369
rect 707 365 708 369
rect 702 364 708 365
rect 671 363 677 364
rect 671 362 672 363
rect 644 360 672 362
rect 615 358 621 359
rect 671 359 672 360
rect 676 359 677 363
rect 712 362 714 376
rect 719 375 720 379
rect 724 378 725 379
rect 743 379 749 380
rect 724 376 739 378
rect 724 375 725 376
rect 719 374 725 375
rect 719 363 725 364
rect 719 362 720 363
rect 712 360 720 362
rect 671 358 677 359
rect 719 359 720 360
rect 724 359 725 363
rect 737 362 739 376
rect 743 375 744 379
rect 748 378 749 379
rect 767 379 773 380
rect 767 378 768 379
rect 748 376 768 378
rect 748 375 749 376
rect 743 374 749 375
rect 767 375 768 376
rect 772 375 773 379
rect 767 374 773 375
rect 823 379 829 380
rect 823 375 824 379
rect 828 378 829 379
rect 879 379 885 380
rect 828 376 874 378
rect 828 375 829 376
rect 823 374 829 375
rect 750 369 756 370
rect 750 365 751 369
rect 755 365 756 369
rect 750 364 756 365
rect 806 369 812 370
rect 806 365 807 369
rect 811 365 812 369
rect 806 364 812 365
rect 862 369 868 370
rect 862 365 863 369
rect 867 365 868 369
rect 862 364 868 365
rect 767 363 773 364
rect 767 362 768 363
rect 737 360 768 362
rect 719 358 725 359
rect 767 359 768 360
rect 772 359 773 363
rect 767 358 773 359
rect 823 363 832 364
rect 823 359 824 363
rect 831 359 832 363
rect 872 362 874 376
rect 879 375 880 379
rect 884 378 885 379
rect 935 379 941 380
rect 884 376 910 378
rect 884 375 885 376
rect 879 374 885 375
rect 879 363 885 364
rect 879 362 880 363
rect 872 360 880 362
rect 823 358 832 359
rect 879 359 880 360
rect 884 359 885 363
rect 908 362 910 376
rect 935 375 936 379
rect 940 378 941 379
rect 999 379 1005 380
rect 940 376 994 378
rect 940 375 941 376
rect 935 374 941 375
rect 918 369 924 370
rect 918 365 919 369
rect 923 365 924 369
rect 918 364 924 365
rect 982 369 988 370
rect 982 365 983 369
rect 987 365 988 369
rect 982 364 988 365
rect 935 363 941 364
rect 935 362 936 363
rect 908 360 936 362
rect 879 358 885 359
rect 935 359 936 360
rect 940 359 941 363
rect 992 362 994 376
rect 999 375 1000 379
rect 1004 378 1005 379
rect 1070 379 1077 380
rect 1004 376 1066 378
rect 1004 375 1005 376
rect 999 374 1005 375
rect 1054 369 1060 370
rect 1054 365 1055 369
rect 1059 365 1060 369
rect 1054 364 1060 365
rect 999 363 1005 364
rect 999 362 1000 363
rect 992 360 1000 362
rect 935 358 941 359
rect 999 359 1000 360
rect 1004 359 1005 363
rect 1064 362 1066 376
rect 1070 375 1071 379
rect 1076 375 1077 379
rect 1070 374 1077 375
rect 1143 379 1149 380
rect 1143 375 1144 379
rect 1148 378 1149 379
rect 1215 379 1221 380
rect 1148 376 1182 378
rect 1148 375 1149 376
rect 1143 374 1149 375
rect 1126 369 1132 370
rect 1126 365 1127 369
rect 1131 365 1132 369
rect 1126 364 1132 365
rect 1071 363 1077 364
rect 1071 362 1072 363
rect 1064 360 1072 362
rect 999 358 1005 359
rect 1071 359 1072 360
rect 1076 359 1077 363
rect 1071 358 1077 359
rect 1143 363 1149 364
rect 1143 359 1144 363
rect 1148 362 1149 363
rect 1158 363 1164 364
rect 1158 362 1159 363
rect 1148 360 1159 362
rect 1148 359 1149 360
rect 1143 358 1149 359
rect 1158 359 1159 360
rect 1163 359 1164 363
rect 1180 362 1182 376
rect 1215 375 1216 379
rect 1220 378 1221 379
rect 1287 379 1293 380
rect 1220 376 1254 378
rect 1220 375 1221 376
rect 1215 374 1221 375
rect 1198 369 1204 370
rect 1198 365 1199 369
rect 1203 365 1204 369
rect 1198 364 1204 365
rect 1215 363 1221 364
rect 1215 362 1216 363
rect 1180 360 1216 362
rect 1158 358 1164 359
rect 1215 359 1216 360
rect 1220 359 1221 363
rect 1252 362 1254 376
rect 1287 375 1288 379
rect 1292 378 1293 379
rect 1354 379 1365 380
rect 1292 376 1326 378
rect 1292 375 1293 376
rect 1287 374 1293 375
rect 1270 369 1276 370
rect 1270 365 1271 369
rect 1275 365 1276 369
rect 1270 364 1276 365
rect 1287 363 1293 364
rect 1287 362 1288 363
rect 1252 360 1288 362
rect 1215 358 1221 359
rect 1287 359 1288 360
rect 1292 359 1293 363
rect 1324 362 1326 376
rect 1354 375 1355 379
rect 1359 375 1360 379
rect 1364 375 1365 379
rect 1354 374 1365 375
rect 1431 379 1437 380
rect 1431 375 1432 379
rect 1436 378 1437 379
rect 1502 379 1509 380
rect 1436 376 1461 378
rect 1436 375 1437 376
rect 1431 374 1437 375
rect 1342 369 1348 370
rect 1342 365 1343 369
rect 1347 365 1348 369
rect 1342 364 1348 365
rect 1414 369 1420 370
rect 1414 365 1415 369
rect 1419 365 1420 369
rect 1414 364 1420 365
rect 1359 363 1365 364
rect 1359 362 1360 363
rect 1324 360 1360 362
rect 1287 358 1293 359
rect 1359 359 1360 360
rect 1364 359 1365 363
rect 1359 358 1365 359
rect 1426 363 1437 364
rect 1426 359 1427 363
rect 1431 359 1432 363
rect 1436 359 1437 363
rect 1459 362 1461 376
rect 1502 375 1503 379
rect 1508 375 1509 379
rect 1502 374 1509 375
rect 1559 379 1565 380
rect 1559 375 1560 379
rect 1564 378 1565 379
rect 1567 379 1573 380
rect 1567 378 1568 379
rect 1564 376 1568 378
rect 1564 375 1565 376
rect 1559 374 1565 375
rect 1567 375 1568 376
rect 1572 375 1573 379
rect 1567 374 1573 375
rect 1486 369 1492 370
rect 1486 365 1487 369
rect 1491 365 1492 369
rect 1486 364 1492 365
rect 1542 369 1548 370
rect 1542 365 1543 369
rect 1547 365 1548 369
rect 1542 364 1548 365
rect 1582 368 1588 369
rect 1582 364 1583 368
rect 1587 364 1588 368
rect 1503 363 1509 364
rect 1503 362 1504 363
rect 1459 360 1504 362
rect 1426 358 1437 359
rect 1503 359 1504 360
rect 1508 359 1509 363
rect 1503 358 1509 359
rect 1558 363 1565 364
rect 1582 363 1588 364
rect 1558 359 1559 363
rect 1564 359 1565 363
rect 1558 358 1565 359
rect 888 356 906 358
rect 888 354 890 356
rect 873 352 890 354
rect 904 354 906 356
rect 944 356 978 358
rect 944 354 946 356
rect 904 352 946 354
rect 976 354 978 356
rect 1008 356 1058 358
rect 1008 354 1010 356
rect 976 352 1010 354
rect 1056 354 1058 356
rect 1070 355 1076 356
rect 1070 354 1071 355
rect 1056 352 1071 354
rect 150 351 157 352
rect 110 348 116 349
rect 110 344 111 348
rect 115 344 116 348
rect 110 343 116 344
rect 134 347 140 348
rect 134 343 135 347
rect 139 343 140 347
rect 150 347 151 351
rect 156 347 157 351
rect 191 351 197 352
rect 191 350 192 351
rect 184 348 192 350
rect 150 346 157 347
rect 174 347 180 348
rect 134 342 140 343
rect 174 343 175 347
rect 179 343 180 347
rect 174 342 180 343
rect 184 338 186 348
rect 191 347 192 348
rect 196 347 197 351
rect 239 351 245 352
rect 239 350 240 351
rect 232 348 240 350
rect 191 346 197 347
rect 222 347 228 348
rect 222 343 223 347
rect 227 343 228 347
rect 222 342 228 343
rect 232 338 234 348
rect 239 347 240 348
rect 244 347 245 351
rect 295 351 301 352
rect 295 350 296 351
rect 288 348 296 350
rect 239 346 245 347
rect 278 347 284 348
rect 278 343 279 347
rect 283 343 284 347
rect 278 342 284 343
rect 288 338 290 348
rect 295 347 296 348
rect 300 347 301 351
rect 351 351 357 352
rect 295 346 301 347
rect 334 347 340 348
rect 334 343 335 347
rect 339 343 340 347
rect 351 347 352 351
rect 356 350 357 351
rect 402 351 413 352
rect 356 348 387 350
rect 356 347 357 348
rect 351 346 357 347
rect 334 342 340 343
rect 172 336 186 338
rect 193 336 234 338
rect 259 336 290 338
rect 385 338 387 348
rect 390 347 396 348
rect 390 343 391 347
rect 395 343 396 347
rect 402 347 403 351
rect 407 347 408 351
rect 412 347 413 351
rect 463 351 469 352
rect 402 346 413 347
rect 446 347 452 348
rect 390 342 396 343
rect 446 343 447 347
rect 451 343 452 347
rect 463 347 464 351
rect 468 350 469 351
rect 494 351 500 352
rect 494 350 495 351
rect 468 348 495 350
rect 468 347 469 348
rect 463 346 469 347
rect 494 347 495 348
rect 499 347 500 351
rect 519 351 525 352
rect 519 350 520 351
rect 512 348 520 350
rect 494 346 500 347
rect 502 347 508 348
rect 446 342 452 343
rect 502 343 503 347
rect 507 343 508 347
rect 502 342 508 343
rect 512 338 514 348
rect 519 347 520 348
rect 524 347 525 351
rect 583 351 589 352
rect 583 350 584 351
rect 576 348 584 350
rect 519 346 525 347
rect 566 347 572 348
rect 566 343 567 347
rect 571 343 572 347
rect 566 342 572 343
rect 576 338 578 348
rect 583 347 584 348
rect 588 347 589 351
rect 647 351 653 352
rect 647 350 648 351
rect 640 348 648 350
rect 583 346 589 347
rect 630 347 636 348
rect 630 343 631 347
rect 635 343 636 347
rect 630 342 636 343
rect 640 338 642 348
rect 647 347 648 348
rect 652 347 653 351
rect 703 351 709 352
rect 703 350 704 351
rect 696 348 704 350
rect 647 346 653 347
rect 686 347 692 348
rect 686 343 687 347
rect 691 343 692 347
rect 686 342 692 343
rect 696 338 698 348
rect 703 347 704 348
rect 708 347 709 351
rect 767 351 773 352
rect 767 350 768 351
rect 760 348 768 350
rect 703 346 709 347
rect 750 347 756 348
rect 750 343 751 347
rect 755 343 756 347
rect 750 342 756 343
rect 760 338 762 348
rect 767 347 768 348
rect 772 347 773 351
rect 831 351 837 352
rect 767 346 773 347
rect 814 347 820 348
rect 814 343 815 347
rect 819 343 820 347
rect 831 347 832 351
rect 836 350 837 351
rect 873 350 875 352
rect 895 351 901 352
rect 895 350 896 351
rect 836 348 875 350
rect 888 348 896 350
rect 836 347 837 348
rect 831 346 837 347
rect 878 347 884 348
rect 814 342 820 343
rect 878 343 879 347
rect 883 343 884 347
rect 878 342 884 343
rect 888 338 890 348
rect 895 347 896 348
rect 900 347 901 351
rect 967 351 973 352
rect 967 350 968 351
rect 960 348 968 350
rect 895 346 901 347
rect 950 347 956 348
rect 950 343 951 347
rect 955 343 956 347
rect 950 342 956 343
rect 960 338 962 348
rect 967 347 968 348
rect 972 347 973 351
rect 1047 351 1053 352
rect 1047 350 1048 351
rect 1040 348 1048 350
rect 967 346 973 347
rect 1030 347 1036 348
rect 1030 343 1031 347
rect 1035 343 1036 347
rect 1030 342 1036 343
rect 1040 338 1042 348
rect 1047 347 1048 348
rect 1052 347 1053 351
rect 1070 351 1071 352
rect 1075 351 1076 355
rect 1228 352 1258 354
rect 1070 350 1076 351
rect 1119 351 1125 352
rect 1119 350 1120 351
rect 1112 348 1120 350
rect 1047 346 1053 347
rect 1102 347 1108 348
rect 1102 343 1103 347
rect 1107 343 1108 347
rect 1102 342 1108 343
rect 1112 338 1114 348
rect 1119 347 1120 348
rect 1124 347 1125 351
rect 1191 351 1197 352
rect 1119 346 1125 347
rect 1174 347 1180 348
rect 1174 343 1175 347
rect 1179 343 1180 347
rect 1191 347 1192 351
rect 1196 350 1197 351
rect 1228 350 1230 352
rect 1196 348 1230 350
rect 1196 347 1197 348
rect 1191 346 1197 347
rect 1246 347 1252 348
rect 1174 342 1180 343
rect 1246 343 1247 347
rect 1251 343 1252 347
rect 1246 342 1252 343
rect 385 336 402 338
rect 492 336 514 338
rect 552 336 578 338
rect 616 336 642 338
rect 676 336 698 338
rect 737 336 762 338
rect 864 336 890 338
rect 897 336 962 338
rect 969 336 1042 338
rect 1099 336 1114 338
rect 151 335 157 336
rect 110 331 116 332
rect 110 327 111 331
rect 115 327 116 331
rect 151 331 152 335
rect 156 334 157 335
rect 172 334 174 336
rect 156 332 174 334
rect 191 335 197 336
rect 156 331 157 332
rect 151 330 157 331
rect 191 331 192 335
rect 196 331 197 335
rect 191 330 197 331
rect 239 335 245 336
rect 239 331 240 335
rect 244 334 245 335
rect 259 334 261 336
rect 244 332 261 334
rect 295 335 301 336
rect 244 331 245 332
rect 239 330 245 331
rect 295 331 296 335
rect 300 334 301 335
rect 310 335 316 336
rect 310 334 311 335
rect 300 332 311 334
rect 300 331 301 332
rect 295 330 301 331
rect 310 331 311 332
rect 315 331 316 335
rect 310 330 316 331
rect 350 335 357 336
rect 350 331 351 335
rect 356 331 357 335
rect 400 334 402 336
rect 407 335 413 336
rect 407 334 408 335
rect 400 332 408 334
rect 350 330 357 331
rect 407 331 408 332
rect 412 331 413 335
rect 407 330 413 331
rect 463 335 469 336
rect 463 331 464 335
rect 468 334 469 335
rect 492 334 494 336
rect 468 332 494 334
rect 519 335 525 336
rect 468 331 469 332
rect 463 330 469 331
rect 519 331 520 335
rect 524 334 525 335
rect 552 334 554 336
rect 524 332 554 334
rect 583 335 589 336
rect 524 331 525 332
rect 519 330 525 331
rect 583 331 584 335
rect 588 334 589 335
rect 616 334 618 336
rect 588 332 618 334
rect 647 335 653 336
rect 588 331 589 332
rect 583 330 589 331
rect 647 331 648 335
rect 652 334 653 335
rect 676 334 678 336
rect 652 332 678 334
rect 703 335 709 336
rect 652 331 653 332
rect 647 330 653 331
rect 703 331 704 335
rect 708 334 709 335
rect 737 334 739 336
rect 767 335 773 336
rect 767 334 768 335
rect 708 332 739 334
rect 760 332 768 334
rect 708 331 709 332
rect 703 330 709 331
rect 110 326 116 327
rect 134 329 140 330
rect 134 325 135 329
rect 139 325 140 329
rect 134 324 140 325
rect 174 329 180 330
rect 174 325 175 329
rect 179 325 180 329
rect 174 324 180 325
rect 222 329 228 330
rect 222 325 223 329
rect 227 325 228 329
rect 222 324 228 325
rect 278 329 284 330
rect 278 325 279 329
rect 283 325 284 329
rect 278 324 284 325
rect 334 329 340 330
rect 334 325 335 329
rect 339 325 340 329
rect 334 324 340 325
rect 390 329 396 330
rect 390 325 391 329
rect 395 325 396 329
rect 390 324 396 325
rect 446 329 452 330
rect 446 325 447 329
rect 451 325 452 329
rect 446 324 452 325
rect 502 329 508 330
rect 502 325 503 329
rect 507 325 508 329
rect 502 324 508 325
rect 566 329 572 330
rect 566 325 567 329
rect 571 325 572 329
rect 566 324 572 325
rect 630 329 636 330
rect 630 325 631 329
rect 635 325 636 329
rect 630 324 636 325
rect 686 329 692 330
rect 686 325 687 329
rect 691 325 692 329
rect 686 324 692 325
rect 750 329 756 330
rect 750 325 751 329
rect 755 325 756 329
rect 750 324 756 325
rect 438 323 444 324
rect 438 319 439 323
rect 443 322 444 323
rect 574 323 580 324
rect 443 320 570 322
rect 443 319 444 320
rect 438 318 444 319
rect 190 315 196 316
rect 110 313 116 314
rect 110 309 111 313
rect 115 309 116 313
rect 190 311 191 315
rect 195 311 196 315
rect 190 310 196 311
rect 222 315 228 316
rect 222 311 223 315
rect 227 311 228 315
rect 222 310 228 311
rect 254 315 260 316
rect 254 311 255 315
rect 259 311 260 315
rect 254 310 260 311
rect 294 315 300 316
rect 294 311 295 315
rect 299 311 300 315
rect 294 310 300 311
rect 334 315 340 316
rect 334 311 335 315
rect 339 311 340 315
rect 334 310 340 311
rect 366 315 372 316
rect 366 311 367 315
rect 371 311 372 315
rect 366 310 372 311
rect 406 315 412 316
rect 406 311 407 315
rect 411 311 412 315
rect 406 310 412 311
rect 454 315 460 316
rect 454 311 455 315
rect 459 311 460 315
rect 454 310 460 311
rect 518 315 524 316
rect 518 311 519 315
rect 523 311 524 315
rect 518 310 524 311
rect 568 310 570 320
rect 574 319 575 323
rect 579 322 580 323
rect 760 322 762 332
rect 767 331 768 332
rect 772 331 773 335
rect 767 330 773 331
rect 831 335 837 336
rect 831 331 832 335
rect 836 334 837 335
rect 864 334 866 336
rect 836 332 866 334
rect 895 335 901 336
rect 836 331 837 332
rect 831 330 837 331
rect 895 331 896 335
rect 900 331 901 335
rect 895 330 901 331
rect 967 335 973 336
rect 967 331 968 335
rect 972 331 973 335
rect 967 330 973 331
rect 1047 335 1053 336
rect 1047 331 1048 335
rect 1052 334 1053 335
rect 1099 334 1101 336
rect 1119 335 1125 336
rect 1119 334 1120 335
rect 1052 332 1101 334
rect 1112 332 1120 334
rect 1052 331 1053 332
rect 1047 330 1053 331
rect 814 329 820 330
rect 814 325 815 329
rect 819 325 820 329
rect 814 324 820 325
rect 878 329 884 330
rect 878 325 879 329
rect 883 325 884 329
rect 878 324 884 325
rect 950 329 956 330
rect 950 325 951 329
rect 955 325 956 329
rect 950 324 956 325
rect 1030 329 1036 330
rect 1030 325 1031 329
rect 1035 325 1036 329
rect 1030 324 1036 325
rect 1102 329 1108 330
rect 1102 325 1103 329
rect 1107 325 1108 329
rect 1102 324 1108 325
rect 579 320 762 322
rect 826 323 832 324
rect 579 319 580 320
rect 574 318 580 319
rect 826 319 827 323
rect 831 322 832 323
rect 1112 322 1114 332
rect 1119 331 1120 332
rect 1124 331 1125 335
rect 1119 330 1125 331
rect 1191 335 1197 336
rect 1191 331 1192 335
rect 1196 334 1197 335
rect 1238 335 1244 336
rect 1238 334 1239 335
rect 1196 332 1239 334
rect 1196 331 1197 332
rect 1191 330 1197 331
rect 1238 331 1239 332
rect 1243 331 1244 335
rect 1256 334 1258 352
rect 1263 351 1269 352
rect 1263 347 1264 351
rect 1268 350 1269 351
rect 1343 351 1349 352
rect 1268 348 1323 350
rect 1268 347 1269 348
rect 1263 346 1269 347
rect 1321 338 1323 348
rect 1326 347 1332 348
rect 1326 343 1327 347
rect 1331 343 1332 347
rect 1343 347 1344 351
rect 1348 350 1349 351
rect 1354 351 1360 352
rect 1354 350 1355 351
rect 1348 348 1355 350
rect 1348 347 1349 348
rect 1343 346 1349 347
rect 1354 347 1355 348
rect 1359 347 1360 351
rect 1423 351 1429 352
rect 1354 346 1360 347
rect 1406 347 1412 348
rect 1326 342 1332 343
rect 1406 343 1407 347
rect 1411 343 1412 347
rect 1423 347 1424 351
rect 1428 350 1429 351
rect 1498 351 1509 352
rect 1428 348 1461 350
rect 1428 347 1429 348
rect 1423 346 1429 347
rect 1406 342 1412 343
rect 1459 338 1461 348
rect 1486 347 1492 348
rect 1486 343 1487 347
rect 1491 343 1492 347
rect 1498 347 1499 351
rect 1503 347 1504 351
rect 1508 347 1509 351
rect 1559 351 1565 352
rect 1498 346 1509 347
rect 1542 347 1548 348
rect 1486 342 1492 343
rect 1542 343 1543 347
rect 1547 343 1548 347
rect 1559 347 1560 351
rect 1564 350 1565 351
rect 1567 351 1573 352
rect 1567 350 1568 351
rect 1564 348 1568 350
rect 1564 347 1565 348
rect 1559 346 1565 347
rect 1567 347 1568 348
rect 1572 347 1573 351
rect 1567 346 1573 347
rect 1582 348 1588 349
rect 1582 344 1583 348
rect 1587 344 1588 348
rect 1582 343 1588 344
rect 1542 342 1548 343
rect 1530 339 1536 340
rect 1321 336 1338 338
rect 1459 336 1498 338
rect 1263 335 1269 336
rect 1263 334 1264 335
rect 1256 332 1264 334
rect 1238 330 1244 331
rect 1263 331 1264 332
rect 1268 331 1269 335
rect 1336 334 1338 336
rect 1343 335 1349 336
rect 1343 334 1344 335
rect 1336 332 1344 334
rect 1263 330 1269 331
rect 1343 331 1344 332
rect 1348 331 1349 335
rect 1343 330 1349 331
rect 1423 335 1432 336
rect 1423 331 1424 335
rect 1431 331 1432 335
rect 1496 334 1498 336
rect 1503 335 1509 336
rect 1503 334 1504 335
rect 1496 332 1504 334
rect 1423 330 1432 331
rect 1503 331 1504 332
rect 1508 331 1509 335
rect 1530 335 1531 339
rect 1535 338 1536 339
rect 1535 336 1554 338
rect 1535 335 1536 336
rect 1530 334 1536 335
rect 1552 334 1554 336
rect 1559 335 1565 336
rect 1559 334 1560 335
rect 1552 332 1560 334
rect 1503 330 1509 331
rect 1559 331 1560 332
rect 1564 331 1565 335
rect 1559 330 1565 331
rect 1582 331 1588 332
rect 1174 329 1180 330
rect 1174 325 1175 329
rect 1179 325 1180 329
rect 1174 324 1180 325
rect 1246 329 1252 330
rect 1246 325 1247 329
rect 1251 325 1252 329
rect 1246 324 1252 325
rect 1326 329 1332 330
rect 1326 325 1327 329
rect 1331 325 1332 329
rect 1326 324 1332 325
rect 1406 329 1412 330
rect 1406 325 1407 329
rect 1411 325 1412 329
rect 1406 324 1412 325
rect 1486 329 1492 330
rect 1486 325 1487 329
rect 1491 325 1492 329
rect 1486 324 1492 325
rect 1542 329 1548 330
rect 1542 325 1543 329
rect 1547 325 1548 329
rect 1582 327 1583 331
rect 1587 327 1588 331
rect 1582 326 1588 327
rect 1542 324 1548 325
rect 831 320 1114 322
rect 831 319 832 320
rect 826 318 832 319
rect 590 315 596 316
rect 590 311 591 315
rect 595 311 596 315
rect 590 310 596 311
rect 662 315 668 316
rect 662 311 663 315
rect 667 311 668 315
rect 662 310 668 311
rect 734 315 740 316
rect 734 311 735 315
rect 739 311 740 315
rect 734 310 740 311
rect 806 315 812 316
rect 806 311 807 315
rect 811 311 812 315
rect 806 310 812 311
rect 878 315 884 316
rect 878 311 879 315
rect 883 311 884 315
rect 878 310 884 311
rect 950 315 956 316
rect 950 311 951 315
rect 955 311 956 315
rect 950 310 956 311
rect 1022 315 1028 316
rect 1022 311 1023 315
rect 1027 311 1028 315
rect 1022 310 1028 311
rect 1094 315 1100 316
rect 1094 311 1095 315
rect 1099 311 1100 315
rect 1094 310 1100 311
rect 1110 315 1116 316
rect 1110 311 1111 315
rect 1115 314 1116 315
rect 1166 315 1172 316
rect 1115 312 1154 314
rect 1115 311 1116 312
rect 1110 310 1116 311
rect 110 308 116 309
rect 568 308 586 310
rect 170 307 176 308
rect 170 303 171 307
rect 175 306 176 307
rect 207 307 213 308
rect 207 306 208 307
rect 175 304 208 306
rect 175 303 176 304
rect 170 302 176 303
rect 207 303 208 304
rect 212 303 213 307
rect 239 307 245 308
rect 239 306 240 307
rect 207 302 213 303
rect 232 304 240 306
rect 190 297 196 298
rect 110 296 116 297
rect 110 292 111 296
rect 115 292 116 296
rect 190 293 191 297
rect 195 293 196 297
rect 190 292 196 293
rect 222 297 228 298
rect 222 293 223 297
rect 227 293 228 297
rect 222 292 228 293
rect 110 291 116 292
rect 207 291 213 292
rect 207 287 208 291
rect 212 290 213 291
rect 232 290 234 304
rect 239 303 240 304
rect 244 303 245 307
rect 271 307 277 308
rect 271 306 272 307
rect 239 302 245 303
rect 264 304 272 306
rect 254 297 260 298
rect 254 293 255 297
rect 259 293 260 297
rect 254 292 260 293
rect 212 288 234 290
rect 239 291 245 292
rect 212 287 213 288
rect 207 286 213 287
rect 239 287 240 291
rect 244 290 245 291
rect 264 290 266 304
rect 271 303 272 304
rect 276 303 277 307
rect 311 307 317 308
rect 311 306 312 307
rect 271 302 277 303
rect 288 304 312 306
rect 244 288 266 290
rect 271 291 277 292
rect 244 287 245 288
rect 239 286 245 287
rect 271 287 272 291
rect 276 290 277 291
rect 288 290 290 304
rect 311 303 312 304
rect 316 303 317 307
rect 311 302 317 303
rect 351 307 357 308
rect 351 303 352 307
rect 356 306 357 307
rect 383 307 389 308
rect 356 304 378 306
rect 356 303 357 304
rect 351 302 357 303
rect 294 297 300 298
rect 294 293 295 297
rect 299 293 300 297
rect 294 292 300 293
rect 334 297 340 298
rect 334 293 335 297
rect 339 293 340 297
rect 334 292 340 293
rect 366 297 372 298
rect 366 293 367 297
rect 371 293 372 297
rect 366 292 372 293
rect 276 288 290 290
rect 310 291 317 292
rect 276 287 277 288
rect 271 286 277 287
rect 310 287 311 291
rect 316 287 317 291
rect 310 286 317 287
rect 342 291 348 292
rect 342 287 343 291
rect 347 290 348 291
rect 351 291 357 292
rect 351 290 352 291
rect 347 288 352 290
rect 347 287 348 288
rect 342 286 348 287
rect 351 287 352 288
rect 356 287 357 291
rect 376 290 378 304
rect 383 303 384 307
rect 388 306 389 307
rect 398 307 404 308
rect 398 306 399 307
rect 388 304 399 306
rect 388 303 389 304
rect 383 302 389 303
rect 398 303 399 304
rect 403 303 404 307
rect 398 302 404 303
rect 423 307 429 308
rect 423 303 424 307
rect 428 306 429 307
rect 471 307 477 308
rect 428 304 450 306
rect 428 303 429 304
rect 423 302 429 303
rect 406 297 412 298
rect 406 293 407 297
rect 411 293 412 297
rect 406 292 412 293
rect 383 291 389 292
rect 383 290 384 291
rect 376 288 384 290
rect 351 286 357 287
rect 383 287 384 288
rect 388 287 389 291
rect 383 286 389 287
rect 423 291 429 292
rect 423 287 424 291
rect 428 290 429 291
rect 438 291 444 292
rect 438 290 439 291
rect 428 288 439 290
rect 428 287 429 288
rect 423 286 429 287
rect 438 287 439 288
rect 443 287 444 291
rect 448 290 450 304
rect 471 303 472 307
rect 476 306 477 307
rect 535 307 541 308
rect 476 304 506 306
rect 476 303 477 304
rect 471 302 477 303
rect 454 297 460 298
rect 454 293 455 297
rect 459 293 460 297
rect 454 292 460 293
rect 471 291 477 292
rect 471 290 472 291
rect 448 288 472 290
rect 438 286 444 287
rect 471 287 472 288
rect 476 287 477 291
rect 504 290 506 304
rect 535 303 536 307
rect 540 306 541 307
rect 584 306 586 308
rect 607 307 613 308
rect 540 304 574 306
rect 584 304 602 306
rect 540 303 541 304
rect 535 302 541 303
rect 518 297 524 298
rect 518 293 519 297
rect 523 293 524 297
rect 518 292 524 293
rect 535 291 541 292
rect 535 290 536 291
rect 504 288 536 290
rect 471 286 477 287
rect 535 287 536 288
rect 540 287 541 291
rect 572 290 574 304
rect 600 298 602 304
rect 607 303 608 307
rect 612 306 613 307
rect 679 307 685 308
rect 612 304 674 306
rect 612 303 613 304
rect 607 302 613 303
rect 654 299 660 300
rect 654 298 655 299
rect 590 297 596 298
rect 590 293 591 297
rect 595 293 596 297
rect 600 296 655 298
rect 654 295 655 296
rect 659 295 660 299
rect 654 294 660 295
rect 662 297 668 298
rect 590 292 596 293
rect 662 293 663 297
rect 667 293 668 297
rect 662 292 668 293
rect 607 291 613 292
rect 607 290 608 291
rect 572 288 608 290
rect 535 286 541 287
rect 607 287 608 288
rect 612 287 613 291
rect 672 290 674 304
rect 679 303 680 307
rect 684 306 685 307
rect 722 307 728 308
rect 684 304 718 306
rect 684 303 685 304
rect 679 302 685 303
rect 679 291 685 292
rect 679 290 680 291
rect 672 288 680 290
rect 607 286 613 287
rect 679 287 680 288
rect 684 287 685 291
rect 716 290 718 304
rect 722 303 723 307
rect 727 306 728 307
rect 751 307 757 308
rect 751 306 752 307
rect 727 304 752 306
rect 727 303 728 304
rect 722 302 728 303
rect 751 303 752 304
rect 756 303 757 307
rect 751 302 757 303
rect 823 307 829 308
rect 823 303 824 307
rect 828 306 829 307
rect 895 307 901 308
rect 828 304 862 306
rect 828 303 829 304
rect 823 302 829 303
rect 734 297 740 298
rect 734 293 735 297
rect 739 293 740 297
rect 734 292 740 293
rect 806 297 812 298
rect 806 293 807 297
rect 811 293 812 297
rect 806 292 812 293
rect 751 291 757 292
rect 751 290 752 291
rect 716 288 752 290
rect 679 286 685 287
rect 751 287 752 288
rect 756 287 757 291
rect 751 286 757 287
rect 823 291 832 292
rect 823 287 824 291
rect 831 287 832 291
rect 860 290 862 304
rect 895 303 896 307
rect 900 306 901 307
rect 967 307 973 308
rect 900 304 934 306
rect 900 303 901 304
rect 895 302 901 303
rect 878 297 884 298
rect 878 293 879 297
rect 883 293 884 297
rect 878 292 884 293
rect 895 291 901 292
rect 895 290 896 291
rect 860 288 896 290
rect 823 286 832 287
rect 895 287 896 288
rect 900 287 901 291
rect 932 290 934 304
rect 967 303 968 307
rect 972 306 973 307
rect 1039 307 1045 308
rect 972 304 1034 306
rect 972 303 973 304
rect 967 302 973 303
rect 950 297 956 298
rect 950 293 951 297
rect 955 293 956 297
rect 950 292 956 293
rect 1022 297 1028 298
rect 1022 293 1023 297
rect 1027 293 1028 297
rect 1022 292 1028 293
rect 967 291 973 292
rect 967 290 968 291
rect 932 288 968 290
rect 895 286 901 287
rect 967 287 968 288
rect 972 287 973 291
rect 1032 290 1034 304
rect 1039 303 1040 307
rect 1044 306 1045 307
rect 1111 307 1117 308
rect 1044 304 1078 306
rect 1044 303 1045 304
rect 1039 302 1045 303
rect 1039 291 1045 292
rect 1039 290 1040 291
rect 1032 288 1040 290
rect 967 286 973 287
rect 1039 287 1040 288
rect 1044 287 1045 291
rect 1076 290 1078 304
rect 1111 303 1112 307
rect 1116 306 1117 307
rect 1152 306 1154 312
rect 1166 311 1167 315
rect 1171 311 1172 315
rect 1166 310 1172 311
rect 1230 315 1236 316
rect 1230 311 1231 315
rect 1235 311 1236 315
rect 1230 310 1236 311
rect 1294 315 1300 316
rect 1294 311 1295 315
rect 1299 311 1300 315
rect 1294 310 1300 311
rect 1350 315 1356 316
rect 1350 311 1351 315
rect 1355 311 1356 315
rect 1350 310 1356 311
rect 1398 315 1404 316
rect 1398 311 1399 315
rect 1403 311 1404 315
rect 1398 310 1404 311
rect 1454 315 1460 316
rect 1454 311 1455 315
rect 1459 311 1460 315
rect 1454 310 1460 311
rect 1510 315 1516 316
rect 1510 311 1511 315
rect 1515 311 1516 315
rect 1510 310 1516 311
rect 1542 315 1548 316
rect 1542 311 1543 315
rect 1547 311 1548 315
rect 1542 310 1548 311
rect 1582 313 1588 314
rect 1582 309 1583 313
rect 1587 309 1588 313
rect 1582 308 1588 309
rect 1183 307 1189 308
rect 1183 306 1184 307
rect 1116 304 1150 306
rect 1152 304 1184 306
rect 1116 303 1117 304
rect 1111 302 1117 303
rect 1094 297 1100 298
rect 1094 293 1095 297
rect 1099 293 1100 297
rect 1094 292 1100 293
rect 1111 291 1117 292
rect 1111 290 1112 291
rect 1076 288 1112 290
rect 1039 286 1045 287
rect 1111 287 1112 288
rect 1116 287 1117 291
rect 1148 290 1150 304
rect 1183 303 1184 304
rect 1188 303 1189 307
rect 1183 302 1189 303
rect 1247 307 1253 308
rect 1247 303 1248 307
rect 1252 306 1253 307
rect 1286 307 1292 308
rect 1252 304 1282 306
rect 1252 303 1253 304
rect 1247 302 1253 303
rect 1166 297 1172 298
rect 1166 293 1167 297
rect 1171 293 1172 297
rect 1166 292 1172 293
rect 1230 297 1236 298
rect 1230 293 1231 297
rect 1235 293 1236 297
rect 1230 292 1236 293
rect 1183 291 1189 292
rect 1183 290 1184 291
rect 1148 288 1184 290
rect 1111 286 1117 287
rect 1183 287 1184 288
rect 1188 287 1189 291
rect 1183 286 1189 287
rect 1238 291 1244 292
rect 1238 287 1239 291
rect 1243 290 1244 291
rect 1247 291 1253 292
rect 1247 290 1248 291
rect 1243 288 1248 290
rect 1243 287 1244 288
rect 1238 286 1244 287
rect 1247 287 1248 288
rect 1252 287 1253 291
rect 1280 290 1282 304
rect 1286 303 1287 307
rect 1291 306 1292 307
rect 1311 307 1317 308
rect 1311 306 1312 307
rect 1291 304 1312 306
rect 1291 303 1292 304
rect 1286 302 1292 303
rect 1311 303 1312 304
rect 1316 303 1317 307
rect 1311 302 1317 303
rect 1367 307 1373 308
rect 1367 303 1368 307
rect 1372 306 1373 307
rect 1415 307 1421 308
rect 1372 304 1394 306
rect 1372 303 1373 304
rect 1367 302 1373 303
rect 1294 297 1300 298
rect 1294 293 1295 297
rect 1299 293 1300 297
rect 1294 292 1300 293
rect 1350 297 1356 298
rect 1350 293 1351 297
rect 1355 293 1356 297
rect 1350 292 1356 293
rect 1311 291 1317 292
rect 1311 290 1312 291
rect 1280 288 1312 290
rect 1247 286 1253 287
rect 1311 287 1312 288
rect 1316 287 1317 291
rect 1311 286 1317 287
rect 1367 291 1373 292
rect 1367 287 1368 291
rect 1372 290 1373 291
rect 1383 291 1389 292
rect 1383 290 1384 291
rect 1372 288 1384 290
rect 1372 287 1373 288
rect 1367 286 1373 287
rect 1383 287 1384 288
rect 1388 287 1389 291
rect 1392 290 1394 304
rect 1415 303 1416 307
rect 1420 306 1421 307
rect 1471 307 1477 308
rect 1420 304 1446 306
rect 1420 303 1421 304
rect 1415 302 1421 303
rect 1398 297 1404 298
rect 1398 293 1399 297
rect 1403 293 1404 297
rect 1398 292 1404 293
rect 1415 291 1421 292
rect 1415 290 1416 291
rect 1392 288 1416 290
rect 1383 286 1389 287
rect 1415 287 1416 288
rect 1420 287 1421 291
rect 1444 290 1446 304
rect 1471 303 1472 307
rect 1476 306 1477 307
rect 1498 307 1504 308
rect 1498 306 1499 307
rect 1476 304 1499 306
rect 1476 303 1477 304
rect 1471 302 1477 303
rect 1498 303 1499 304
rect 1503 303 1504 307
rect 1498 302 1504 303
rect 1527 307 1533 308
rect 1527 303 1528 307
rect 1532 306 1533 307
rect 1558 307 1565 308
rect 1532 304 1554 306
rect 1532 303 1533 304
rect 1527 302 1533 303
rect 1454 297 1460 298
rect 1454 293 1455 297
rect 1459 293 1460 297
rect 1454 292 1460 293
rect 1510 297 1516 298
rect 1510 293 1511 297
rect 1515 293 1516 297
rect 1510 292 1516 293
rect 1542 297 1548 298
rect 1542 293 1543 297
rect 1547 293 1548 297
rect 1542 292 1548 293
rect 1471 291 1477 292
rect 1471 290 1472 291
rect 1444 288 1472 290
rect 1415 286 1421 287
rect 1471 287 1472 288
rect 1476 287 1477 291
rect 1471 286 1477 287
rect 1527 291 1536 292
rect 1527 287 1528 291
rect 1535 287 1536 291
rect 1552 290 1554 304
rect 1558 303 1559 307
rect 1564 303 1565 307
rect 1558 302 1565 303
rect 1582 296 1588 297
rect 1582 292 1583 296
rect 1587 292 1588 296
rect 1559 291 1565 292
rect 1582 291 1588 292
rect 1559 290 1560 291
rect 1552 288 1560 290
rect 1527 286 1536 287
rect 1559 287 1560 288
rect 1564 287 1565 291
rect 1559 286 1565 287
rect 494 283 500 284
rect 494 279 495 283
rect 499 282 500 283
rect 722 283 728 284
rect 722 282 723 283
rect 499 280 723 282
rect 499 279 500 280
rect 494 278 500 279
rect 722 279 723 280
rect 727 279 728 283
rect 1110 283 1116 284
rect 1110 282 1111 283
rect 722 278 728 279
rect 841 280 1111 282
rect 208 276 226 278
rect 841 276 843 280
rect 1110 279 1111 280
rect 1115 279 1116 283
rect 1286 283 1292 284
rect 1286 282 1287 283
rect 1256 280 1287 282
rect 1110 278 1116 279
rect 1143 279 1149 280
rect 167 275 176 276
rect 110 272 116 273
rect 110 268 111 272
rect 115 268 116 272
rect 110 267 116 268
rect 150 271 156 272
rect 150 267 151 271
rect 155 267 156 271
rect 167 271 168 275
rect 175 271 176 275
rect 199 275 205 276
rect 199 274 200 275
rect 192 272 200 274
rect 167 270 176 271
rect 182 271 188 272
rect 150 266 156 267
rect 182 267 183 271
rect 187 267 188 271
rect 182 266 188 267
rect 192 262 194 272
rect 199 271 200 272
rect 204 271 205 275
rect 199 270 205 271
rect 172 260 194 262
rect 167 259 174 260
rect 110 255 116 256
rect 110 251 111 255
rect 115 251 116 255
rect 167 255 168 259
rect 172 256 174 259
rect 199 259 205 260
rect 172 255 173 256
rect 167 254 173 255
rect 199 255 200 259
rect 204 258 205 259
rect 208 258 210 276
rect 224 274 226 276
rect 231 275 237 276
rect 231 274 232 275
rect 224 272 232 274
rect 214 271 220 272
rect 214 267 215 271
rect 219 267 220 271
rect 231 271 232 272
rect 236 271 237 275
rect 263 275 272 276
rect 231 270 237 271
rect 246 271 252 272
rect 214 266 220 267
rect 246 267 247 271
rect 251 267 252 271
rect 263 271 264 275
rect 271 271 272 275
rect 295 275 301 276
rect 295 274 296 275
rect 288 272 296 274
rect 263 270 272 271
rect 278 271 284 272
rect 246 266 252 267
rect 278 267 279 271
rect 283 267 284 271
rect 278 266 284 267
rect 288 262 290 272
rect 295 271 296 272
rect 300 271 301 275
rect 327 275 333 276
rect 327 274 328 275
rect 320 272 328 274
rect 295 270 301 271
rect 310 271 316 272
rect 310 267 311 271
rect 315 267 316 271
rect 310 266 316 267
rect 320 262 322 272
rect 327 271 328 272
rect 332 271 333 275
rect 367 275 373 276
rect 327 270 333 271
rect 350 271 356 272
rect 350 267 351 271
rect 355 267 356 271
rect 367 271 368 275
rect 372 274 373 275
rect 398 275 404 276
rect 398 274 399 275
rect 372 272 399 274
rect 372 271 373 272
rect 367 270 373 271
rect 398 271 399 272
rect 403 271 404 275
rect 423 275 429 276
rect 423 274 424 275
rect 416 272 424 274
rect 398 270 404 271
rect 406 271 412 272
rect 350 266 356 267
rect 406 267 407 271
rect 411 267 412 271
rect 406 266 412 267
rect 416 262 418 272
rect 423 271 424 272
rect 428 271 429 275
rect 495 275 501 276
rect 495 274 496 275
rect 488 272 496 274
rect 423 270 429 271
rect 478 271 484 272
rect 478 267 479 271
rect 483 267 484 271
rect 478 266 484 267
rect 488 262 490 272
rect 495 271 496 272
rect 500 271 501 275
rect 575 275 581 276
rect 575 274 576 275
rect 568 272 576 274
rect 495 270 501 271
rect 558 271 564 272
rect 558 267 559 271
rect 563 267 564 271
rect 558 266 564 267
rect 568 262 570 272
rect 575 271 576 272
rect 580 271 581 275
rect 663 275 669 276
rect 663 274 664 275
rect 656 272 664 274
rect 575 270 581 271
rect 646 271 652 272
rect 646 267 647 271
rect 651 267 652 271
rect 646 266 652 267
rect 656 262 658 272
rect 663 271 664 272
rect 668 271 669 275
rect 751 275 757 276
rect 751 274 752 275
rect 744 272 752 274
rect 663 270 669 271
rect 734 271 740 272
rect 734 267 735 271
rect 739 267 740 271
rect 734 266 740 267
rect 744 262 746 272
rect 751 271 752 272
rect 756 271 757 275
rect 839 275 845 276
rect 751 270 757 271
rect 822 271 828 272
rect 822 267 823 271
rect 827 267 828 271
rect 839 271 840 275
rect 844 271 845 275
rect 919 275 925 276
rect 919 274 920 275
rect 912 272 920 274
rect 839 270 845 271
rect 902 271 908 272
rect 822 266 828 267
rect 902 267 903 271
rect 907 267 908 271
rect 902 266 908 267
rect 912 262 914 272
rect 919 271 920 272
rect 924 271 925 275
rect 999 275 1005 276
rect 999 274 1000 275
rect 992 272 1000 274
rect 919 270 925 271
rect 982 271 988 272
rect 982 267 983 271
rect 987 267 988 271
rect 982 266 988 267
rect 992 262 994 272
rect 999 271 1000 272
rect 1004 271 1005 275
rect 1071 275 1077 276
rect 1071 274 1072 275
rect 1064 272 1072 274
rect 999 270 1005 271
rect 1054 271 1060 272
rect 1054 267 1055 271
rect 1059 267 1060 271
rect 1054 266 1060 267
rect 1064 262 1066 272
rect 1071 271 1072 272
rect 1076 271 1077 275
rect 1135 275 1141 276
rect 1135 274 1136 275
rect 1128 272 1136 274
rect 1071 270 1077 271
rect 1118 271 1124 272
rect 1118 267 1119 271
rect 1123 267 1124 271
rect 1118 266 1124 267
rect 1128 262 1130 272
rect 1135 271 1136 272
rect 1140 271 1141 275
rect 1143 275 1144 279
rect 1148 278 1149 279
rect 1148 276 1195 278
rect 1148 275 1149 276
rect 1143 274 1149 275
rect 1191 275 1197 276
rect 1135 270 1141 271
rect 1174 271 1180 272
rect 1174 267 1175 271
rect 1179 267 1180 271
rect 1191 271 1192 275
rect 1196 271 1197 275
rect 1239 275 1245 276
rect 1191 270 1197 271
rect 1222 271 1228 272
rect 1174 266 1180 267
rect 1222 267 1223 271
rect 1227 267 1228 271
rect 1239 271 1240 275
rect 1244 274 1245 275
rect 1256 274 1258 280
rect 1286 279 1287 280
rect 1291 279 1292 283
rect 1286 278 1292 279
rect 1327 279 1333 280
rect 1279 275 1285 276
rect 1279 274 1280 275
rect 1244 272 1258 274
rect 1272 272 1280 274
rect 1244 271 1245 272
rect 1239 270 1245 271
rect 1262 271 1268 272
rect 1222 266 1228 267
rect 1262 267 1263 271
rect 1267 267 1268 271
rect 1262 266 1268 267
rect 1272 262 1274 272
rect 1279 271 1280 272
rect 1284 271 1285 275
rect 1319 275 1325 276
rect 1319 274 1320 275
rect 1312 272 1320 274
rect 1279 270 1285 271
rect 1302 271 1308 272
rect 1302 267 1303 271
rect 1307 267 1308 271
rect 1302 266 1308 267
rect 1312 262 1314 272
rect 1319 271 1320 272
rect 1324 271 1325 275
rect 1327 275 1328 279
rect 1332 278 1333 279
rect 1332 276 1362 278
rect 1332 275 1333 276
rect 1327 274 1333 275
rect 1360 274 1362 276
rect 1367 275 1373 276
rect 1367 274 1368 275
rect 1360 272 1368 274
rect 1319 270 1325 271
rect 1350 271 1356 272
rect 1350 267 1351 271
rect 1355 267 1356 271
rect 1367 271 1368 272
rect 1372 271 1373 275
rect 1415 275 1421 276
rect 1367 270 1373 271
rect 1398 271 1404 272
rect 1350 266 1356 267
rect 1398 267 1399 271
rect 1403 267 1404 271
rect 1415 271 1416 275
rect 1420 274 1421 275
rect 1463 275 1469 276
rect 1420 272 1442 274
rect 1420 271 1421 272
rect 1415 270 1421 271
rect 1398 266 1404 267
rect 276 260 290 262
rect 308 260 322 262
rect 396 260 418 262
rect 460 260 490 262
rect 536 260 570 262
rect 619 260 658 262
rect 708 260 746 262
rect 841 260 914 262
rect 960 260 994 262
rect 1036 260 1066 262
rect 1099 260 1130 262
rect 1260 260 1274 262
rect 1300 260 1314 262
rect 1383 263 1389 264
rect 204 256 210 258
rect 226 259 237 260
rect 204 255 205 256
rect 199 254 205 255
rect 226 255 227 259
rect 231 255 232 259
rect 236 255 237 259
rect 226 254 237 255
rect 263 259 269 260
rect 263 255 264 259
rect 268 258 269 259
rect 276 258 278 260
rect 268 256 278 258
rect 295 259 301 260
rect 268 255 269 256
rect 263 254 269 255
rect 295 255 296 259
rect 300 258 301 259
rect 308 258 310 260
rect 300 256 310 258
rect 327 259 333 260
rect 300 255 301 256
rect 295 254 301 255
rect 327 255 328 259
rect 332 258 333 259
rect 342 259 348 260
rect 342 258 343 259
rect 332 256 343 258
rect 332 255 333 256
rect 327 254 333 255
rect 342 255 343 256
rect 347 255 348 259
rect 342 254 348 255
rect 367 259 373 260
rect 367 255 368 259
rect 372 258 373 259
rect 396 258 398 260
rect 372 256 398 258
rect 423 259 429 260
rect 372 255 373 256
rect 367 254 373 255
rect 423 255 424 259
rect 428 258 429 259
rect 460 258 462 260
rect 428 256 462 258
rect 495 259 501 260
rect 428 255 429 256
rect 423 254 429 255
rect 495 255 496 259
rect 500 258 501 259
rect 536 258 538 260
rect 500 256 538 258
rect 575 259 581 260
rect 500 255 501 256
rect 495 254 501 255
rect 575 255 576 259
rect 580 258 581 259
rect 619 258 621 260
rect 580 256 621 258
rect 663 259 669 260
rect 580 255 581 256
rect 575 254 581 255
rect 663 255 664 259
rect 668 258 669 259
rect 708 258 710 260
rect 751 259 757 260
rect 751 258 752 259
rect 668 256 710 258
rect 744 256 752 258
rect 668 255 669 256
rect 663 254 669 255
rect 110 250 116 251
rect 150 253 156 254
rect 150 249 151 253
rect 155 249 156 253
rect 150 248 156 249
rect 182 253 188 254
rect 182 249 183 253
rect 187 249 188 253
rect 182 248 188 249
rect 214 253 220 254
rect 214 249 215 253
rect 219 249 220 253
rect 214 248 220 249
rect 246 253 252 254
rect 246 249 247 253
rect 251 249 252 253
rect 246 248 252 249
rect 278 253 284 254
rect 278 249 279 253
rect 283 249 284 253
rect 278 248 284 249
rect 310 253 316 254
rect 310 249 311 253
rect 315 249 316 253
rect 310 248 316 249
rect 350 253 356 254
rect 350 249 351 253
rect 355 249 356 253
rect 350 248 356 249
rect 406 253 412 254
rect 406 249 407 253
rect 411 249 412 253
rect 406 248 412 249
rect 478 253 484 254
rect 478 249 479 253
rect 483 249 484 253
rect 478 248 484 249
rect 558 253 564 254
rect 558 249 559 253
rect 563 249 564 253
rect 558 248 564 249
rect 646 253 652 254
rect 646 249 647 253
rect 651 249 652 253
rect 646 248 652 249
rect 734 253 740 254
rect 734 249 735 253
rect 739 249 740 253
rect 734 248 740 249
rect 462 247 468 248
rect 462 243 463 247
rect 467 246 468 247
rect 654 247 660 248
rect 467 244 621 246
rect 467 243 468 244
rect 462 242 468 243
rect 134 239 140 240
rect 110 237 116 238
rect 110 233 111 237
rect 115 233 116 237
rect 134 235 135 239
rect 139 235 140 239
rect 134 234 140 235
rect 166 239 172 240
rect 166 235 167 239
rect 171 235 172 239
rect 166 234 172 235
rect 206 239 212 240
rect 206 235 207 239
rect 211 235 212 239
rect 206 234 212 235
rect 254 239 260 240
rect 254 235 255 239
rect 259 235 260 239
rect 254 234 260 235
rect 302 239 308 240
rect 302 235 303 239
rect 307 235 308 239
rect 302 234 308 235
rect 342 239 348 240
rect 342 235 343 239
rect 347 235 348 239
rect 342 234 348 235
rect 382 239 388 240
rect 382 235 383 239
rect 387 235 388 239
rect 382 234 388 235
rect 438 239 444 240
rect 438 235 439 239
rect 443 235 444 239
rect 438 234 444 235
rect 510 239 516 240
rect 510 235 511 239
rect 515 235 516 239
rect 510 234 516 235
rect 590 239 596 240
rect 590 235 591 239
rect 595 235 596 239
rect 590 234 596 235
rect 619 234 621 244
rect 654 243 655 247
rect 659 246 660 247
rect 744 246 746 256
rect 751 255 752 256
rect 756 255 757 259
rect 751 254 757 255
rect 839 259 845 260
rect 839 255 840 259
rect 844 255 845 259
rect 839 254 845 255
rect 919 259 925 260
rect 919 255 920 259
rect 924 258 925 259
rect 960 258 962 260
rect 924 256 962 258
rect 999 259 1005 260
rect 924 255 925 256
rect 919 254 925 255
rect 999 255 1000 259
rect 1004 258 1005 259
rect 1036 258 1038 260
rect 1004 256 1038 258
rect 1071 259 1077 260
rect 1004 255 1005 256
rect 999 254 1005 255
rect 1071 255 1072 259
rect 1076 258 1077 259
rect 1099 258 1101 260
rect 1076 256 1101 258
rect 1135 259 1141 260
rect 1076 255 1077 256
rect 1071 254 1077 255
rect 1135 255 1136 259
rect 1140 258 1141 259
rect 1143 259 1149 260
rect 1143 258 1144 259
rect 1140 256 1144 258
rect 1140 255 1141 256
rect 1135 254 1141 255
rect 1143 255 1144 256
rect 1148 255 1149 259
rect 1143 254 1149 255
rect 1186 259 1197 260
rect 1186 255 1187 259
rect 1191 255 1192 259
rect 1196 255 1197 259
rect 1186 254 1197 255
rect 1239 259 1245 260
rect 1239 255 1240 259
rect 1244 258 1245 259
rect 1260 258 1262 260
rect 1244 256 1262 258
rect 1279 259 1285 260
rect 1244 255 1245 256
rect 1239 254 1245 255
rect 1279 255 1280 259
rect 1284 258 1285 259
rect 1300 258 1302 260
rect 1284 256 1302 258
rect 1319 259 1325 260
rect 1284 255 1285 256
rect 1279 254 1285 255
rect 1319 255 1320 259
rect 1324 258 1325 259
rect 1327 259 1333 260
rect 1327 258 1328 259
rect 1324 256 1328 258
rect 1324 255 1325 256
rect 1319 254 1325 255
rect 1327 255 1328 256
rect 1332 255 1333 259
rect 1327 254 1333 255
rect 1362 259 1373 260
rect 1362 255 1363 259
rect 1367 255 1368 259
rect 1372 255 1373 259
rect 1383 259 1384 263
rect 1388 262 1389 263
rect 1440 262 1442 272
rect 1446 271 1452 272
rect 1446 267 1447 271
rect 1451 267 1452 271
rect 1463 271 1464 275
rect 1468 274 1469 275
rect 1518 275 1525 276
rect 1468 272 1498 274
rect 1468 271 1469 272
rect 1463 270 1469 271
rect 1446 266 1452 267
rect 1496 262 1498 272
rect 1502 271 1508 272
rect 1502 267 1503 271
rect 1507 267 1508 271
rect 1518 271 1519 275
rect 1524 271 1525 275
rect 1558 275 1565 276
rect 1518 270 1525 271
rect 1542 271 1548 272
rect 1502 266 1508 267
rect 1542 267 1543 271
rect 1547 267 1548 271
rect 1558 271 1559 275
rect 1564 271 1565 275
rect 1558 270 1565 271
rect 1582 272 1588 273
rect 1582 268 1583 272
rect 1587 268 1588 272
rect 1582 267 1588 268
rect 1542 266 1548 267
rect 1388 260 1410 262
rect 1440 260 1458 262
rect 1496 260 1514 262
rect 1388 259 1389 260
rect 1383 258 1389 259
rect 1408 258 1410 260
rect 1415 259 1421 260
rect 1415 258 1416 259
rect 1408 256 1416 258
rect 1362 254 1373 255
rect 1415 255 1416 256
rect 1420 255 1421 259
rect 1456 258 1458 260
rect 1463 259 1469 260
rect 1463 258 1464 259
rect 1456 256 1464 258
rect 1415 254 1421 255
rect 1463 255 1464 256
rect 1468 255 1469 259
rect 1512 258 1514 260
rect 1519 259 1525 260
rect 1519 258 1520 259
rect 1512 256 1520 258
rect 1463 254 1469 255
rect 1519 255 1520 256
rect 1524 255 1525 259
rect 1519 254 1525 255
rect 1558 259 1565 260
rect 1558 255 1559 259
rect 1564 255 1565 259
rect 1558 254 1565 255
rect 1582 255 1588 256
rect 822 253 828 254
rect 822 249 823 253
rect 827 249 828 253
rect 822 248 828 249
rect 902 253 908 254
rect 902 249 903 253
rect 907 249 908 253
rect 902 248 908 249
rect 982 253 988 254
rect 982 249 983 253
rect 987 249 988 253
rect 982 248 988 249
rect 1054 253 1060 254
rect 1054 249 1055 253
rect 1059 249 1060 253
rect 1054 248 1060 249
rect 1118 253 1124 254
rect 1118 249 1119 253
rect 1123 249 1124 253
rect 1118 248 1124 249
rect 1174 253 1180 254
rect 1174 249 1175 253
rect 1179 249 1180 253
rect 1174 248 1180 249
rect 1222 253 1228 254
rect 1222 249 1223 253
rect 1227 249 1228 253
rect 1222 248 1228 249
rect 1262 253 1268 254
rect 1262 249 1263 253
rect 1267 249 1268 253
rect 1262 248 1268 249
rect 1302 253 1308 254
rect 1302 249 1303 253
rect 1307 249 1308 253
rect 1302 248 1308 249
rect 1350 253 1356 254
rect 1350 249 1351 253
rect 1355 249 1356 253
rect 1350 248 1356 249
rect 1398 253 1404 254
rect 1398 249 1399 253
rect 1403 249 1404 253
rect 1398 248 1404 249
rect 1446 253 1452 254
rect 1446 249 1447 253
rect 1451 249 1452 253
rect 1446 248 1452 249
rect 1502 253 1508 254
rect 1502 249 1503 253
rect 1507 249 1508 253
rect 1502 248 1508 249
rect 1542 253 1548 254
rect 1542 249 1543 253
rect 1547 249 1548 253
rect 1582 251 1583 255
rect 1587 251 1588 255
rect 1582 250 1588 251
rect 1542 248 1548 249
rect 659 244 746 246
rect 659 243 660 244
rect 654 242 660 243
rect 678 239 684 240
rect 678 235 679 239
rect 683 235 684 239
rect 758 239 764 240
rect 758 238 759 239
rect 678 234 684 235
rect 688 236 759 238
rect 110 232 116 233
rect 619 232 662 234
rect 150 231 157 232
rect 150 227 151 231
rect 156 227 157 231
rect 183 231 189 232
rect 183 230 184 231
rect 150 226 157 227
rect 176 228 184 230
rect 134 221 140 222
rect 110 220 116 221
rect 110 216 111 220
rect 115 216 116 220
rect 134 217 135 221
rect 139 217 140 221
rect 134 216 140 217
rect 166 221 172 222
rect 166 217 167 221
rect 171 217 172 221
rect 166 216 172 217
rect 110 215 116 216
rect 151 215 157 216
rect 151 211 152 215
rect 156 214 157 215
rect 176 214 178 228
rect 183 227 184 228
rect 188 227 189 231
rect 223 231 229 232
rect 223 230 224 231
rect 183 226 189 227
rect 196 228 224 230
rect 156 212 178 214
rect 183 215 189 216
rect 156 211 157 212
rect 151 210 157 211
rect 183 211 184 215
rect 188 214 189 215
rect 196 214 198 228
rect 223 227 224 228
rect 228 227 229 231
rect 223 226 229 227
rect 266 231 277 232
rect 266 227 267 231
rect 271 227 272 231
rect 276 227 277 231
rect 319 231 325 232
rect 319 230 320 231
rect 266 226 277 227
rect 296 228 320 230
rect 206 221 212 222
rect 206 217 207 221
rect 211 217 212 221
rect 206 216 212 217
rect 254 221 260 222
rect 254 217 255 221
rect 259 217 260 221
rect 254 216 260 217
rect 188 212 198 214
rect 223 215 232 216
rect 188 211 189 212
rect 183 210 189 211
rect 223 211 224 215
rect 231 211 232 215
rect 223 210 232 211
rect 271 215 277 216
rect 271 211 272 215
rect 276 214 277 215
rect 296 214 298 228
rect 319 227 320 228
rect 324 227 325 231
rect 359 231 365 232
rect 359 230 360 231
rect 319 226 325 227
rect 336 228 360 230
rect 302 221 308 222
rect 302 217 303 221
rect 307 217 308 221
rect 302 216 308 217
rect 276 212 298 214
rect 319 215 325 216
rect 276 211 277 212
rect 271 210 277 211
rect 319 211 320 215
rect 324 214 325 215
rect 336 214 338 228
rect 359 227 360 228
rect 364 227 365 231
rect 359 226 365 227
rect 398 231 405 232
rect 398 227 399 231
rect 404 227 405 231
rect 455 231 461 232
rect 455 230 456 231
rect 398 226 405 227
rect 432 228 456 230
rect 342 221 348 222
rect 342 217 343 221
rect 347 217 348 221
rect 342 216 348 217
rect 382 221 388 222
rect 382 217 383 221
rect 387 217 388 221
rect 382 216 388 217
rect 324 212 338 214
rect 359 215 365 216
rect 324 211 325 212
rect 319 210 325 211
rect 359 211 360 215
rect 364 214 365 215
rect 374 215 380 216
rect 374 214 375 215
rect 364 212 375 214
rect 364 211 365 212
rect 359 210 365 211
rect 374 211 375 212
rect 379 211 380 215
rect 374 210 380 211
rect 399 215 405 216
rect 399 211 400 215
rect 404 214 405 215
rect 432 214 434 228
rect 455 227 456 228
rect 460 227 461 231
rect 527 231 533 232
rect 527 230 528 231
rect 455 226 461 227
rect 492 228 528 230
rect 438 221 444 222
rect 438 217 439 221
rect 443 217 444 221
rect 438 216 444 217
rect 404 212 434 214
rect 455 215 461 216
rect 404 211 405 212
rect 399 210 405 211
rect 455 211 456 215
rect 460 214 461 215
rect 492 214 494 228
rect 527 227 528 228
rect 532 227 533 231
rect 527 226 533 227
rect 607 231 613 232
rect 607 227 608 231
rect 612 230 613 231
rect 660 230 662 232
rect 688 230 690 236
rect 758 235 759 236
rect 763 235 764 239
rect 758 234 764 235
rect 766 239 772 240
rect 766 235 767 239
rect 771 235 772 239
rect 766 234 772 235
rect 846 239 852 240
rect 846 235 847 239
rect 851 235 852 239
rect 846 234 852 235
rect 918 239 924 240
rect 918 235 919 239
rect 923 235 924 239
rect 918 234 924 235
rect 982 239 988 240
rect 982 235 983 239
rect 987 235 988 239
rect 982 234 988 235
rect 1046 239 1052 240
rect 1046 235 1047 239
rect 1051 235 1052 239
rect 1046 234 1052 235
rect 1102 239 1108 240
rect 1102 235 1103 239
rect 1107 235 1108 239
rect 1102 234 1108 235
rect 1158 239 1164 240
rect 1158 235 1159 239
rect 1163 235 1164 239
rect 1158 234 1164 235
rect 1214 239 1220 240
rect 1214 235 1215 239
rect 1219 235 1220 239
rect 1214 234 1220 235
rect 1270 239 1276 240
rect 1270 235 1271 239
rect 1275 235 1276 239
rect 1270 234 1276 235
rect 1326 239 1332 240
rect 1326 235 1327 239
rect 1331 235 1332 239
rect 1326 234 1332 235
rect 1382 239 1388 240
rect 1382 235 1383 239
rect 1387 235 1388 239
rect 1382 234 1388 235
rect 1438 239 1444 240
rect 1438 235 1439 239
rect 1443 235 1444 239
rect 1438 234 1444 235
rect 1502 239 1508 240
rect 1502 235 1503 239
rect 1507 235 1508 239
rect 1502 234 1508 235
rect 1542 239 1548 240
rect 1542 235 1543 239
rect 1547 235 1548 239
rect 1542 234 1548 235
rect 1582 237 1588 238
rect 1582 233 1583 237
rect 1587 233 1588 237
rect 1582 232 1588 233
rect 612 228 621 230
rect 660 228 690 230
rect 695 231 701 232
rect 612 227 613 228
rect 607 226 613 227
rect 510 221 516 222
rect 510 217 511 221
rect 515 217 516 221
rect 510 216 516 217
rect 590 221 596 222
rect 590 217 591 221
rect 595 217 596 221
rect 590 216 596 217
rect 460 212 494 214
rect 527 215 533 216
rect 460 211 461 212
rect 455 210 461 211
rect 527 211 528 215
rect 532 214 533 215
rect 554 215 560 216
rect 532 212 550 214
rect 532 211 533 212
rect 527 210 533 211
rect 548 206 550 212
rect 554 211 555 215
rect 559 214 560 215
rect 607 215 613 216
rect 607 214 608 215
rect 559 212 608 214
rect 559 211 560 212
rect 554 210 560 211
rect 607 211 608 212
rect 612 211 613 215
rect 619 214 621 228
rect 695 227 696 231
rect 700 230 701 231
rect 751 231 757 232
rect 700 228 742 230
rect 700 227 701 228
rect 695 226 701 227
rect 678 221 684 222
rect 678 217 679 221
rect 683 217 684 221
rect 678 216 684 217
rect 695 215 701 216
rect 695 214 696 215
rect 619 212 696 214
rect 607 210 613 211
rect 695 211 696 212
rect 700 211 701 215
rect 740 214 742 228
rect 751 227 752 231
rect 756 230 757 231
rect 783 231 789 232
rect 783 230 784 231
rect 756 228 784 230
rect 756 227 757 228
rect 751 226 757 227
rect 783 227 784 228
rect 788 227 789 231
rect 783 226 789 227
rect 863 231 869 232
rect 863 227 864 231
rect 868 230 869 231
rect 935 231 941 232
rect 868 228 902 230
rect 868 227 869 228
rect 863 226 869 227
rect 766 221 772 222
rect 766 217 767 221
rect 771 217 772 221
rect 766 216 772 217
rect 846 221 852 222
rect 846 217 847 221
rect 851 217 852 221
rect 846 216 852 217
rect 783 215 789 216
rect 783 214 784 215
rect 740 212 784 214
rect 695 210 701 211
rect 783 211 784 212
rect 788 211 789 215
rect 783 210 789 211
rect 863 215 869 216
rect 863 211 864 215
rect 868 214 869 215
rect 900 214 902 228
rect 935 227 936 231
rect 940 230 941 231
rect 999 231 1005 232
rect 940 228 970 230
rect 940 227 941 228
rect 935 226 941 227
rect 918 221 924 222
rect 918 217 919 221
rect 923 217 924 221
rect 918 216 924 217
rect 935 215 941 216
rect 935 214 936 215
rect 868 212 898 214
rect 900 212 936 214
rect 868 211 869 212
rect 863 210 869 211
rect 751 207 757 208
rect 751 206 752 207
rect 548 204 752 206
rect 239 203 245 204
rect 150 199 157 200
rect 110 196 116 197
rect 110 192 111 196
rect 115 192 116 196
rect 110 191 116 192
rect 134 195 140 196
rect 134 191 135 195
rect 139 191 140 195
rect 150 195 151 199
rect 156 195 157 199
rect 183 199 189 200
rect 183 198 184 199
rect 176 196 184 198
rect 150 194 157 195
rect 166 195 172 196
rect 134 190 140 191
rect 166 191 167 195
rect 171 191 172 195
rect 166 190 172 191
rect 176 186 178 196
rect 183 195 184 196
rect 188 195 189 199
rect 231 199 237 200
rect 231 198 232 199
rect 224 196 232 198
rect 183 194 189 195
rect 214 195 220 196
rect 214 191 215 195
rect 219 191 220 195
rect 214 190 220 191
rect 224 186 226 196
rect 231 195 232 196
rect 236 195 237 199
rect 239 199 240 203
rect 244 202 245 203
rect 751 203 752 204
rect 756 203 757 207
rect 896 206 898 212
rect 935 211 936 212
rect 940 211 941 215
rect 968 214 970 228
rect 999 227 1000 231
rect 1004 230 1005 231
rect 1022 231 1028 232
rect 1022 230 1023 231
rect 1004 228 1023 230
rect 1004 227 1005 228
rect 999 226 1005 227
rect 1022 227 1023 228
rect 1027 227 1028 231
rect 1022 226 1028 227
rect 1030 231 1036 232
rect 1030 227 1031 231
rect 1035 230 1036 231
rect 1063 231 1069 232
rect 1063 230 1064 231
rect 1035 228 1064 230
rect 1035 227 1036 228
rect 1030 226 1036 227
rect 1063 227 1064 228
rect 1068 227 1069 231
rect 1119 231 1125 232
rect 1119 230 1120 231
rect 1063 226 1069 227
rect 1092 228 1120 230
rect 982 221 988 222
rect 982 217 983 221
rect 987 217 988 221
rect 982 216 988 217
rect 1046 221 1052 222
rect 1046 217 1047 221
rect 1051 217 1052 221
rect 1046 216 1052 217
rect 999 215 1005 216
rect 999 214 1000 215
rect 968 212 1000 214
rect 935 210 941 211
rect 999 211 1000 212
rect 1004 211 1005 215
rect 999 210 1005 211
rect 1063 215 1069 216
rect 1063 211 1064 215
rect 1068 214 1069 215
rect 1092 214 1094 228
rect 1119 227 1120 228
rect 1124 227 1125 231
rect 1175 231 1181 232
rect 1175 230 1176 231
rect 1119 226 1125 227
rect 1148 228 1176 230
rect 1102 221 1108 222
rect 1102 217 1103 221
rect 1107 217 1108 221
rect 1102 216 1108 217
rect 1068 212 1094 214
rect 1119 215 1125 216
rect 1068 211 1069 212
rect 1063 210 1069 211
rect 1119 211 1120 215
rect 1124 214 1125 215
rect 1148 214 1150 228
rect 1175 227 1176 228
rect 1180 227 1181 231
rect 1175 226 1181 227
rect 1231 231 1237 232
rect 1231 227 1232 231
rect 1236 230 1237 231
rect 1246 231 1252 232
rect 1246 230 1247 231
rect 1236 228 1247 230
rect 1236 227 1237 228
rect 1231 226 1237 227
rect 1246 227 1247 228
rect 1251 227 1252 231
rect 1287 231 1293 232
rect 1287 230 1288 231
rect 1246 226 1252 227
rect 1260 228 1288 230
rect 1158 221 1164 222
rect 1158 217 1159 221
rect 1163 217 1164 221
rect 1158 216 1164 217
rect 1214 221 1220 222
rect 1214 217 1215 221
rect 1219 217 1220 221
rect 1214 216 1220 217
rect 1124 212 1150 214
rect 1175 215 1181 216
rect 1124 211 1125 212
rect 1119 210 1125 211
rect 1175 211 1176 215
rect 1180 214 1181 215
rect 1186 215 1192 216
rect 1186 214 1187 215
rect 1180 212 1187 214
rect 1180 211 1181 212
rect 1175 210 1181 211
rect 1186 211 1187 212
rect 1191 211 1192 215
rect 1186 210 1192 211
rect 1231 215 1237 216
rect 1231 211 1232 215
rect 1236 214 1237 215
rect 1260 214 1262 228
rect 1287 227 1288 228
rect 1292 227 1293 231
rect 1343 231 1349 232
rect 1343 230 1344 231
rect 1287 226 1293 227
rect 1320 228 1344 230
rect 1270 221 1276 222
rect 1270 217 1271 221
rect 1275 217 1276 221
rect 1270 216 1276 217
rect 1236 212 1262 214
rect 1287 215 1293 216
rect 1236 211 1237 212
rect 1231 210 1237 211
rect 1287 211 1288 215
rect 1292 214 1293 215
rect 1320 214 1322 228
rect 1343 227 1344 228
rect 1348 227 1349 231
rect 1343 226 1349 227
rect 1399 231 1405 232
rect 1399 227 1400 231
rect 1404 230 1405 231
rect 1455 231 1461 232
rect 1404 228 1430 230
rect 1404 227 1405 228
rect 1399 226 1405 227
rect 1326 221 1332 222
rect 1326 217 1327 221
rect 1331 217 1332 221
rect 1326 216 1332 217
rect 1382 221 1388 222
rect 1382 217 1383 221
rect 1387 217 1388 221
rect 1382 216 1388 217
rect 1292 212 1322 214
rect 1343 215 1349 216
rect 1292 211 1293 212
rect 1287 210 1293 211
rect 1343 211 1344 215
rect 1348 214 1349 215
rect 1362 215 1368 216
rect 1362 214 1363 215
rect 1348 212 1363 214
rect 1348 211 1349 212
rect 1343 210 1349 211
rect 1362 211 1363 212
rect 1367 211 1368 215
rect 1362 210 1368 211
rect 1399 215 1405 216
rect 1399 211 1400 215
rect 1404 214 1405 215
rect 1428 214 1430 228
rect 1455 227 1456 231
rect 1460 230 1461 231
rect 1518 231 1525 232
rect 1460 228 1490 230
rect 1460 227 1461 228
rect 1455 226 1461 227
rect 1438 221 1444 222
rect 1438 217 1439 221
rect 1443 217 1444 221
rect 1438 216 1444 217
rect 1455 215 1461 216
rect 1455 214 1456 215
rect 1404 212 1426 214
rect 1428 212 1456 214
rect 1404 211 1405 212
rect 1399 210 1405 211
rect 1030 207 1036 208
rect 1030 206 1031 207
rect 896 204 1031 206
rect 751 202 757 203
rect 1030 203 1031 204
rect 1035 203 1036 207
rect 1302 207 1308 208
rect 1302 206 1303 207
rect 1030 202 1036 203
rect 1193 204 1303 206
rect 244 200 274 202
rect 1193 200 1195 204
rect 1302 203 1303 204
rect 1307 203 1308 207
rect 1424 206 1426 212
rect 1455 211 1456 212
rect 1460 211 1461 215
rect 1488 214 1490 228
rect 1518 227 1519 231
rect 1524 227 1525 231
rect 1518 226 1525 227
rect 1559 231 1565 232
rect 1559 227 1560 231
rect 1564 230 1565 231
rect 1567 231 1573 232
rect 1567 230 1568 231
rect 1564 228 1568 230
rect 1564 227 1565 228
rect 1559 226 1565 227
rect 1567 227 1568 228
rect 1572 227 1573 231
rect 1567 226 1573 227
rect 1502 221 1508 222
rect 1502 217 1503 221
rect 1507 217 1508 221
rect 1502 216 1508 217
rect 1542 221 1548 222
rect 1542 217 1543 221
rect 1547 217 1548 221
rect 1542 216 1548 217
rect 1582 220 1588 221
rect 1582 216 1583 220
rect 1587 216 1588 220
rect 1519 215 1525 216
rect 1519 214 1520 215
rect 1488 212 1520 214
rect 1455 210 1461 211
rect 1519 211 1520 212
rect 1524 211 1525 215
rect 1519 210 1525 211
rect 1558 215 1565 216
rect 1582 215 1588 216
rect 1558 211 1559 215
rect 1564 211 1565 215
rect 1558 210 1565 211
rect 1470 207 1476 208
rect 1470 206 1471 207
rect 1424 204 1471 206
rect 1302 202 1308 203
rect 1470 203 1471 204
rect 1475 203 1476 207
rect 1470 202 1476 203
rect 244 199 245 200
rect 239 198 245 199
rect 272 198 274 200
rect 279 199 285 200
rect 279 198 280 199
rect 272 196 280 198
rect 231 194 237 195
rect 262 195 268 196
rect 262 191 263 195
rect 267 191 268 195
rect 279 195 280 196
rect 284 195 285 199
rect 322 199 333 200
rect 279 194 285 195
rect 310 195 316 196
rect 262 190 268 191
rect 310 191 311 195
rect 315 191 316 195
rect 322 195 323 199
rect 327 195 328 199
rect 332 195 333 199
rect 375 199 381 200
rect 375 198 376 199
rect 368 196 376 198
rect 322 194 333 195
rect 358 195 364 196
rect 310 190 316 191
rect 358 191 359 195
rect 363 191 364 195
rect 358 190 364 191
rect 368 186 370 196
rect 375 195 376 196
rect 380 195 381 199
rect 431 199 437 200
rect 375 194 381 195
rect 414 195 420 196
rect 414 191 415 195
rect 419 191 420 195
rect 431 195 432 199
rect 436 198 437 199
rect 462 199 468 200
rect 462 198 463 199
rect 436 196 463 198
rect 436 195 437 196
rect 431 194 437 195
rect 462 195 463 196
rect 467 195 468 199
rect 487 199 493 200
rect 487 198 488 199
rect 480 196 488 198
rect 462 194 468 195
rect 470 195 476 196
rect 414 190 420 191
rect 470 191 471 195
rect 475 191 476 195
rect 470 190 476 191
rect 480 186 482 196
rect 487 195 488 196
rect 492 195 493 199
rect 551 199 557 200
rect 551 198 552 199
rect 544 196 552 198
rect 487 194 493 195
rect 534 195 540 196
rect 534 191 535 195
rect 539 191 540 195
rect 534 190 540 191
rect 544 186 546 196
rect 551 195 552 196
rect 556 195 557 199
rect 618 199 629 200
rect 551 194 557 195
rect 606 195 612 196
rect 606 191 607 195
rect 611 191 612 195
rect 618 195 619 199
rect 623 195 624 199
rect 628 195 629 199
rect 695 199 701 200
rect 695 198 696 199
rect 688 196 696 198
rect 618 194 629 195
rect 678 195 684 196
rect 606 190 612 191
rect 678 191 679 195
rect 683 191 684 195
rect 678 190 684 191
rect 688 186 690 196
rect 695 195 696 196
rect 700 195 701 199
rect 767 199 773 200
rect 767 198 768 199
rect 760 196 768 198
rect 695 194 701 195
rect 750 195 756 196
rect 750 191 751 195
rect 755 191 756 195
rect 750 190 756 191
rect 760 186 762 196
rect 767 195 768 196
rect 772 195 773 199
rect 831 199 837 200
rect 767 194 773 195
rect 814 195 820 196
rect 814 191 815 195
rect 819 191 820 195
rect 831 195 832 199
rect 836 198 837 199
rect 870 199 876 200
rect 870 198 871 199
rect 836 196 871 198
rect 836 195 837 196
rect 831 194 837 195
rect 870 195 871 196
rect 875 195 876 199
rect 895 199 901 200
rect 895 198 896 199
rect 888 196 896 198
rect 870 194 876 195
rect 878 195 884 196
rect 814 190 820 191
rect 878 191 879 195
rect 883 191 884 195
rect 878 190 884 191
rect 888 186 890 196
rect 895 195 896 196
rect 900 195 901 199
rect 959 199 965 200
rect 959 198 960 199
rect 952 196 960 198
rect 895 194 901 195
rect 942 195 948 196
rect 942 191 943 195
rect 947 191 948 195
rect 942 190 948 191
rect 952 186 954 196
rect 959 195 960 196
rect 964 195 965 199
rect 1022 199 1029 200
rect 959 194 965 195
rect 1006 195 1012 196
rect 1006 191 1007 195
rect 1011 191 1012 195
rect 1022 195 1023 199
rect 1028 195 1029 199
rect 1079 199 1085 200
rect 1079 198 1080 199
rect 1072 196 1080 198
rect 1022 194 1029 195
rect 1062 195 1068 196
rect 1006 190 1012 191
rect 1062 191 1063 195
rect 1067 191 1068 195
rect 1062 190 1068 191
rect 1072 186 1074 196
rect 1079 195 1080 196
rect 1084 195 1085 199
rect 1135 199 1141 200
rect 1135 198 1136 199
rect 1128 196 1136 198
rect 1079 194 1085 195
rect 1118 195 1124 196
rect 1118 191 1119 195
rect 1123 191 1124 195
rect 1118 190 1124 191
rect 1128 186 1130 196
rect 1135 195 1136 196
rect 1140 195 1141 199
rect 1191 199 1197 200
rect 1135 194 1141 195
rect 1174 195 1180 196
rect 1174 191 1175 195
rect 1179 191 1180 195
rect 1191 195 1192 199
rect 1196 195 1197 199
rect 1246 199 1253 200
rect 1191 194 1197 195
rect 1230 195 1236 196
rect 1174 190 1180 191
rect 1230 191 1231 195
rect 1235 191 1236 195
rect 1246 195 1247 199
rect 1252 195 1253 199
rect 1303 199 1309 200
rect 1303 198 1304 199
rect 1296 196 1304 198
rect 1246 194 1253 195
rect 1286 195 1292 196
rect 1230 190 1236 191
rect 1286 191 1287 195
rect 1291 191 1292 195
rect 1286 190 1292 191
rect 1296 186 1298 196
rect 1303 195 1304 196
rect 1308 195 1309 199
rect 1359 199 1368 200
rect 1303 194 1309 195
rect 1342 195 1348 196
rect 1342 191 1343 195
rect 1347 191 1348 195
rect 1359 195 1360 199
rect 1367 195 1368 199
rect 1415 199 1421 200
rect 1415 198 1416 199
rect 1408 196 1416 198
rect 1359 194 1368 195
rect 1398 195 1404 196
rect 1342 190 1348 191
rect 1398 191 1399 195
rect 1403 191 1404 195
rect 1398 190 1404 191
rect 1408 186 1410 196
rect 1415 195 1416 196
rect 1420 195 1421 199
rect 1471 199 1477 200
rect 1471 198 1472 199
rect 1464 196 1472 198
rect 1415 194 1421 195
rect 1454 195 1460 196
rect 1454 191 1455 195
rect 1459 191 1460 195
rect 1454 190 1460 191
rect 1464 186 1466 196
rect 1471 195 1472 196
rect 1476 195 1477 199
rect 1527 199 1533 200
rect 1471 194 1477 195
rect 1510 195 1516 196
rect 1510 191 1511 195
rect 1515 191 1516 195
rect 1527 195 1528 199
rect 1532 198 1533 199
rect 1559 199 1565 200
rect 1532 196 1538 198
rect 1532 195 1533 196
rect 1527 194 1533 195
rect 1510 190 1516 191
rect 153 184 178 186
rect 208 184 226 186
rect 352 184 370 186
rect 460 184 482 186
rect 520 184 546 186
rect 660 184 690 186
rect 732 184 762 186
rect 864 184 890 186
rect 928 184 954 186
rect 1052 184 1074 186
rect 1099 184 1130 186
rect 1276 184 1298 186
rect 1388 184 1410 186
rect 1444 184 1466 186
rect 1536 186 1538 196
rect 1542 195 1548 196
rect 1542 191 1543 195
rect 1547 191 1548 195
rect 1559 195 1560 199
rect 1564 198 1565 199
rect 1567 199 1573 200
rect 1567 198 1568 199
rect 1564 196 1568 198
rect 1564 195 1565 196
rect 1559 194 1565 195
rect 1567 195 1568 196
rect 1572 195 1573 199
rect 1567 194 1573 195
rect 1582 196 1588 197
rect 1582 192 1583 196
rect 1587 192 1588 196
rect 1582 191 1588 192
rect 1542 190 1548 191
rect 1536 184 1563 186
rect 151 183 157 184
rect 110 179 116 180
rect 110 175 111 179
rect 115 175 116 179
rect 151 179 152 183
rect 156 179 157 183
rect 151 178 157 179
rect 183 183 189 184
rect 183 179 184 183
rect 188 182 189 183
rect 208 182 210 184
rect 188 180 210 182
rect 231 183 237 184
rect 188 179 189 180
rect 183 178 189 179
rect 231 179 232 183
rect 236 182 237 183
rect 239 183 245 184
rect 239 182 240 183
rect 236 180 240 182
rect 236 179 237 180
rect 231 178 237 179
rect 239 179 240 180
rect 244 179 245 183
rect 239 178 245 179
rect 274 183 285 184
rect 274 179 275 183
rect 279 179 280 183
rect 284 179 285 183
rect 274 178 285 179
rect 327 183 333 184
rect 327 179 328 183
rect 332 182 333 183
rect 352 182 354 184
rect 332 180 354 182
rect 374 183 381 184
rect 332 179 333 180
rect 327 178 333 179
rect 374 179 375 183
rect 380 179 381 183
rect 374 178 381 179
rect 431 183 437 184
rect 431 179 432 183
rect 436 182 437 183
rect 460 182 462 184
rect 436 180 462 182
rect 487 183 493 184
rect 436 179 437 180
rect 431 178 437 179
rect 487 179 488 183
rect 492 182 493 183
rect 520 182 522 184
rect 492 180 522 182
rect 551 183 560 184
rect 492 179 493 180
rect 487 178 493 179
rect 551 179 552 183
rect 559 179 560 183
rect 551 178 560 179
rect 623 183 629 184
rect 623 179 624 183
rect 628 182 629 183
rect 660 182 662 184
rect 628 180 662 182
rect 695 183 701 184
rect 628 179 629 180
rect 623 178 629 179
rect 695 179 696 183
rect 700 182 701 183
rect 732 182 734 184
rect 700 180 734 182
rect 766 183 773 184
rect 700 179 701 180
rect 695 178 701 179
rect 766 179 767 183
rect 772 179 773 183
rect 766 178 773 179
rect 831 183 837 184
rect 831 179 832 183
rect 836 182 837 183
rect 864 182 866 184
rect 836 180 866 182
rect 895 183 901 184
rect 836 179 837 180
rect 831 178 837 179
rect 895 179 896 183
rect 900 182 901 183
rect 928 182 930 184
rect 900 180 930 182
rect 959 183 965 184
rect 900 179 901 180
rect 895 178 901 179
rect 959 179 960 183
rect 964 182 965 183
rect 990 183 996 184
rect 990 182 991 183
rect 964 180 991 182
rect 964 179 965 180
rect 959 178 965 179
rect 990 179 991 180
rect 995 179 996 183
rect 990 178 996 179
rect 1023 183 1029 184
rect 1023 179 1024 183
rect 1028 182 1029 183
rect 1052 182 1054 184
rect 1028 180 1054 182
rect 1079 183 1085 184
rect 1028 179 1029 180
rect 1023 178 1029 179
rect 1079 179 1080 183
rect 1084 182 1085 183
rect 1099 182 1101 184
rect 1135 183 1141 184
rect 1135 182 1136 183
rect 1084 180 1101 182
rect 1128 180 1136 182
rect 1084 179 1085 180
rect 1079 178 1085 179
rect 110 174 116 175
rect 134 177 140 178
rect 134 173 135 177
rect 139 173 140 177
rect 134 172 140 173
rect 166 177 172 178
rect 166 173 167 177
rect 171 173 172 177
rect 166 172 172 173
rect 214 177 220 178
rect 214 173 215 177
rect 219 173 220 177
rect 214 172 220 173
rect 262 177 268 178
rect 262 173 263 177
rect 267 173 268 177
rect 262 172 268 173
rect 310 177 316 178
rect 310 173 311 177
rect 315 173 316 177
rect 310 172 316 173
rect 358 177 364 178
rect 358 173 359 177
rect 363 173 364 177
rect 358 172 364 173
rect 414 177 420 178
rect 414 173 415 177
rect 419 173 420 177
rect 414 172 420 173
rect 470 177 476 178
rect 470 173 471 177
rect 475 173 476 177
rect 470 172 476 173
rect 534 177 540 178
rect 534 173 535 177
rect 539 173 540 177
rect 534 172 540 173
rect 606 177 612 178
rect 606 173 607 177
rect 611 173 612 177
rect 606 172 612 173
rect 678 177 684 178
rect 678 173 679 177
rect 683 173 684 177
rect 678 172 684 173
rect 750 177 756 178
rect 750 173 751 177
rect 755 173 756 177
rect 750 172 756 173
rect 814 177 820 178
rect 814 173 815 177
rect 819 173 820 177
rect 814 172 820 173
rect 878 177 884 178
rect 878 173 879 177
rect 883 173 884 177
rect 878 172 884 173
rect 942 177 948 178
rect 942 173 943 177
rect 947 173 948 177
rect 942 172 948 173
rect 1006 177 1012 178
rect 1006 173 1007 177
rect 1011 173 1012 177
rect 1006 172 1012 173
rect 1062 177 1068 178
rect 1062 173 1063 177
rect 1067 173 1068 177
rect 1062 172 1068 173
rect 1118 177 1124 178
rect 1118 173 1119 177
rect 1123 173 1124 177
rect 1118 172 1124 173
rect 482 171 488 172
rect 482 167 483 171
rect 487 170 488 171
rect 870 171 876 172
rect 487 168 738 170
rect 487 167 488 168
rect 482 166 488 167
rect 142 163 148 164
rect 110 161 116 162
rect 110 157 111 161
rect 115 157 116 161
rect 142 159 143 163
rect 147 159 148 163
rect 142 158 148 159
rect 190 163 196 164
rect 190 159 191 163
rect 195 159 196 163
rect 190 158 196 159
rect 238 163 244 164
rect 238 159 239 163
rect 243 159 244 163
rect 238 158 244 159
rect 294 163 300 164
rect 294 159 295 163
rect 299 159 300 163
rect 294 158 300 159
rect 350 163 356 164
rect 350 159 351 163
rect 355 159 356 163
rect 350 158 356 159
rect 406 163 412 164
rect 406 159 407 163
rect 411 159 412 163
rect 406 158 412 159
rect 462 163 468 164
rect 462 159 463 163
rect 467 159 468 163
rect 462 158 468 159
rect 518 163 524 164
rect 518 159 519 163
rect 523 159 524 163
rect 518 158 524 159
rect 574 163 580 164
rect 574 159 575 163
rect 579 159 580 163
rect 574 158 580 159
rect 630 163 636 164
rect 630 159 631 163
rect 635 159 636 163
rect 630 158 636 159
rect 686 163 692 164
rect 686 159 687 163
rect 691 159 692 163
rect 686 158 692 159
rect 110 156 116 157
rect 154 155 165 156
rect 154 151 155 155
rect 159 151 160 155
rect 164 151 165 155
rect 207 155 213 156
rect 207 154 208 155
rect 154 150 165 151
rect 184 152 208 154
rect 142 145 148 146
rect 110 144 116 145
rect 110 140 111 144
rect 115 140 116 144
rect 142 141 143 145
rect 147 141 148 145
rect 142 140 148 141
rect 110 139 116 140
rect 159 139 165 140
rect 159 135 160 139
rect 164 138 165 139
rect 184 138 186 152
rect 207 151 208 152
rect 212 151 213 155
rect 255 155 261 156
rect 255 154 256 155
rect 207 150 213 151
rect 232 152 256 154
rect 190 145 196 146
rect 190 141 191 145
rect 195 141 196 145
rect 190 140 196 141
rect 164 136 186 138
rect 207 139 213 140
rect 164 135 165 136
rect 159 134 165 135
rect 207 135 208 139
rect 212 138 213 139
rect 232 138 234 152
rect 255 151 256 152
rect 260 151 261 155
rect 255 150 261 151
rect 311 155 317 156
rect 311 151 312 155
rect 316 154 317 155
rect 322 155 328 156
rect 322 154 323 155
rect 316 152 323 154
rect 316 151 317 152
rect 311 150 317 151
rect 322 151 323 152
rect 327 151 328 155
rect 367 155 373 156
rect 367 154 368 155
rect 322 150 328 151
rect 340 152 368 154
rect 238 145 244 146
rect 238 141 239 145
rect 243 141 244 145
rect 238 140 244 141
rect 294 145 300 146
rect 294 141 295 145
rect 299 141 300 145
rect 294 140 300 141
rect 212 136 234 138
rect 255 139 261 140
rect 212 135 213 136
rect 207 134 213 135
rect 255 135 256 139
rect 260 138 261 139
rect 274 139 280 140
rect 274 138 275 139
rect 260 136 275 138
rect 260 135 261 136
rect 255 134 261 135
rect 274 135 275 136
rect 279 135 280 139
rect 274 134 280 135
rect 311 139 317 140
rect 311 135 312 139
rect 316 138 317 139
rect 340 138 342 152
rect 367 151 368 152
rect 372 151 373 155
rect 423 155 429 156
rect 423 154 424 155
rect 367 150 373 151
rect 396 152 424 154
rect 350 145 356 146
rect 350 141 351 145
rect 355 141 356 145
rect 350 140 356 141
rect 316 136 342 138
rect 367 139 373 140
rect 316 135 317 136
rect 311 134 317 135
rect 367 135 368 139
rect 372 138 373 139
rect 396 138 398 152
rect 423 151 424 152
rect 428 151 429 155
rect 423 150 429 151
rect 479 155 485 156
rect 479 151 480 155
rect 484 154 485 155
rect 535 155 541 156
rect 484 152 510 154
rect 484 151 485 152
rect 479 150 485 151
rect 406 145 412 146
rect 406 141 407 145
rect 411 141 412 145
rect 406 140 412 141
rect 462 145 468 146
rect 462 141 463 145
rect 467 141 468 145
rect 462 140 468 141
rect 372 136 398 138
rect 423 139 429 140
rect 372 135 373 136
rect 367 134 373 135
rect 423 135 424 139
rect 428 138 429 139
rect 438 139 444 140
rect 438 138 439 139
rect 428 136 439 138
rect 428 135 429 136
rect 423 134 429 135
rect 438 135 439 136
rect 443 135 444 139
rect 438 134 444 135
rect 479 139 488 140
rect 479 135 480 139
rect 487 135 488 139
rect 508 138 510 152
rect 535 151 536 155
rect 540 154 541 155
rect 591 155 597 156
rect 540 152 566 154
rect 540 151 541 152
rect 535 150 541 151
rect 518 145 524 146
rect 518 141 519 145
rect 523 141 524 145
rect 518 140 524 141
rect 535 139 541 140
rect 535 138 536 139
rect 508 136 536 138
rect 479 134 488 135
rect 535 135 536 136
rect 540 135 541 139
rect 564 138 566 152
rect 591 151 592 155
rect 596 154 597 155
rect 618 155 624 156
rect 618 154 619 155
rect 596 152 619 154
rect 596 151 597 152
rect 591 150 597 151
rect 618 151 619 152
rect 623 151 624 155
rect 618 150 624 151
rect 647 155 653 156
rect 647 151 648 155
rect 652 154 653 155
rect 703 155 709 156
rect 652 152 678 154
rect 652 151 653 152
rect 647 150 653 151
rect 574 145 580 146
rect 574 141 575 145
rect 579 141 580 145
rect 574 140 580 141
rect 630 145 636 146
rect 630 141 631 145
rect 635 141 636 145
rect 630 140 636 141
rect 591 139 597 140
rect 591 138 592 139
rect 564 136 592 138
rect 535 134 541 135
rect 591 135 592 136
rect 596 135 597 139
rect 647 139 653 140
rect 647 138 648 139
rect 591 134 597 135
rect 600 136 648 138
rect 538 131 544 132
rect 538 127 539 131
rect 543 130 544 131
rect 600 130 602 136
rect 647 135 648 136
rect 652 135 653 139
rect 676 138 678 152
rect 703 151 704 155
rect 708 154 709 155
rect 736 154 738 168
rect 870 167 871 171
rect 875 170 876 171
rect 1128 170 1130 180
rect 1135 179 1136 180
rect 1140 179 1141 183
rect 1135 178 1141 179
rect 1186 183 1197 184
rect 1186 179 1187 183
rect 1191 179 1192 183
rect 1196 179 1197 183
rect 1186 178 1197 179
rect 1247 183 1253 184
rect 1247 179 1248 183
rect 1252 182 1253 183
rect 1276 182 1278 184
rect 1252 180 1278 182
rect 1302 183 1309 184
rect 1252 179 1253 180
rect 1247 178 1253 179
rect 1302 179 1303 183
rect 1308 179 1309 183
rect 1302 178 1309 179
rect 1359 183 1365 184
rect 1359 179 1360 183
rect 1364 182 1365 183
rect 1388 182 1390 184
rect 1364 180 1390 182
rect 1415 183 1421 184
rect 1364 179 1365 180
rect 1359 178 1365 179
rect 1415 179 1416 183
rect 1420 182 1421 183
rect 1444 182 1446 184
rect 1420 180 1446 182
rect 1470 183 1477 184
rect 1420 179 1421 180
rect 1415 178 1421 179
rect 1470 179 1471 183
rect 1476 179 1477 183
rect 1470 178 1477 179
rect 1526 183 1533 184
rect 1526 179 1527 183
rect 1532 179 1533 183
rect 1526 178 1533 179
rect 1559 183 1565 184
rect 1559 179 1560 183
rect 1564 179 1565 183
rect 1559 178 1565 179
rect 1582 179 1588 180
rect 1174 177 1180 178
rect 1174 173 1175 177
rect 1179 173 1180 177
rect 1174 172 1180 173
rect 1230 177 1236 178
rect 1230 173 1231 177
rect 1235 173 1236 177
rect 1230 172 1236 173
rect 1286 177 1292 178
rect 1286 173 1287 177
rect 1291 173 1292 177
rect 1286 172 1292 173
rect 1342 177 1348 178
rect 1342 173 1343 177
rect 1347 173 1348 177
rect 1342 172 1348 173
rect 1398 177 1404 178
rect 1398 173 1399 177
rect 1403 173 1404 177
rect 1398 172 1404 173
rect 1454 177 1460 178
rect 1454 173 1455 177
rect 1459 173 1460 177
rect 1454 172 1460 173
rect 1510 177 1516 178
rect 1510 173 1511 177
rect 1515 173 1516 177
rect 1510 172 1516 173
rect 1542 177 1548 178
rect 1542 173 1543 177
rect 1547 173 1548 177
rect 1582 175 1583 179
rect 1587 175 1588 179
rect 1582 174 1588 175
rect 1542 172 1548 173
rect 875 168 1130 170
rect 875 167 876 168
rect 870 166 876 167
rect 742 163 748 164
rect 742 159 743 163
rect 747 159 748 163
rect 742 158 748 159
rect 798 163 804 164
rect 798 159 799 163
rect 803 159 804 163
rect 798 158 804 159
rect 854 163 860 164
rect 854 159 855 163
rect 859 159 860 163
rect 854 158 860 159
rect 910 163 916 164
rect 910 159 911 163
rect 915 159 916 163
rect 910 158 916 159
rect 974 163 980 164
rect 974 159 975 163
rect 979 159 980 163
rect 974 158 980 159
rect 1038 163 1044 164
rect 1038 159 1039 163
rect 1043 159 1044 163
rect 1038 158 1044 159
rect 1094 163 1100 164
rect 1094 159 1095 163
rect 1099 159 1100 163
rect 1094 158 1100 159
rect 1150 163 1156 164
rect 1150 159 1151 163
rect 1155 159 1156 163
rect 1150 158 1156 159
rect 1206 163 1212 164
rect 1206 159 1207 163
rect 1211 159 1212 163
rect 1206 158 1212 159
rect 1254 163 1260 164
rect 1254 159 1255 163
rect 1259 159 1260 163
rect 1254 158 1260 159
rect 1302 163 1308 164
rect 1302 159 1303 163
rect 1307 159 1308 163
rect 1302 158 1308 159
rect 1350 163 1356 164
rect 1350 159 1351 163
rect 1355 159 1356 163
rect 1350 158 1356 159
rect 1398 163 1404 164
rect 1398 159 1399 163
rect 1403 159 1404 163
rect 1398 158 1404 159
rect 1454 163 1460 164
rect 1454 159 1455 163
rect 1459 159 1460 163
rect 1454 158 1460 159
rect 1510 163 1516 164
rect 1510 159 1511 163
rect 1515 159 1516 163
rect 1510 158 1516 159
rect 1542 163 1548 164
rect 1542 159 1543 163
rect 1547 159 1548 163
rect 1542 158 1548 159
rect 1582 161 1588 162
rect 1582 157 1583 161
rect 1587 157 1588 161
rect 1582 156 1588 157
rect 759 155 765 156
rect 759 154 760 155
rect 708 152 734 154
rect 736 152 760 154
rect 708 151 709 152
rect 703 150 709 151
rect 686 145 692 146
rect 686 141 687 145
rect 691 141 692 145
rect 686 140 692 141
rect 703 139 709 140
rect 703 138 704 139
rect 676 136 704 138
rect 647 134 653 135
rect 703 135 704 136
rect 708 135 709 139
rect 732 138 734 152
rect 759 151 760 152
rect 764 151 765 155
rect 759 150 765 151
rect 815 155 821 156
rect 815 151 816 155
rect 820 154 821 155
rect 871 155 877 156
rect 820 152 846 154
rect 820 151 821 152
rect 815 150 821 151
rect 742 145 748 146
rect 742 141 743 145
rect 747 141 748 145
rect 742 140 748 141
rect 798 145 804 146
rect 798 141 799 145
rect 803 141 804 145
rect 798 140 804 141
rect 759 139 765 140
rect 759 138 760 139
rect 732 136 760 138
rect 703 134 709 135
rect 759 135 760 136
rect 764 135 765 139
rect 759 134 765 135
rect 815 139 821 140
rect 815 135 816 139
rect 820 138 821 139
rect 844 138 846 152
rect 871 151 872 155
rect 876 154 877 155
rect 927 155 933 156
rect 876 152 902 154
rect 876 151 877 152
rect 871 150 877 151
rect 854 145 860 146
rect 854 141 855 145
rect 859 141 860 145
rect 854 140 860 141
rect 871 139 877 140
rect 871 138 872 139
rect 820 136 838 138
rect 844 136 872 138
rect 820 135 821 136
rect 815 134 821 135
rect 543 128 602 130
rect 836 130 838 136
rect 871 135 872 136
rect 876 135 877 139
rect 900 138 902 152
rect 927 151 928 155
rect 932 154 933 155
rect 967 155 973 156
rect 967 154 968 155
rect 932 152 968 154
rect 932 151 933 152
rect 927 150 933 151
rect 967 151 968 152
rect 972 151 973 155
rect 967 150 973 151
rect 991 155 997 156
rect 991 151 992 155
rect 996 154 997 155
rect 1055 155 1061 156
rect 996 152 1026 154
rect 996 151 997 152
rect 991 150 997 151
rect 910 145 916 146
rect 910 141 911 145
rect 915 141 916 145
rect 910 140 916 141
rect 974 145 980 146
rect 974 141 975 145
rect 979 141 980 145
rect 974 140 980 141
rect 927 139 933 140
rect 927 138 928 139
rect 900 136 928 138
rect 871 134 877 135
rect 927 135 928 136
rect 932 135 933 139
rect 927 134 933 135
rect 990 139 997 140
rect 990 135 991 139
rect 996 135 997 139
rect 1024 138 1026 152
rect 1055 151 1056 155
rect 1060 154 1061 155
rect 1106 155 1117 156
rect 1060 152 1086 154
rect 1060 151 1061 152
rect 1055 150 1061 151
rect 1038 145 1044 146
rect 1038 141 1039 145
rect 1043 141 1044 145
rect 1038 140 1044 141
rect 1055 139 1061 140
rect 1055 138 1056 139
rect 1024 136 1056 138
rect 990 134 997 135
rect 1055 135 1056 136
rect 1060 135 1061 139
rect 1084 138 1086 152
rect 1106 151 1107 155
rect 1111 151 1112 155
rect 1116 151 1117 155
rect 1106 150 1117 151
rect 1167 155 1173 156
rect 1167 151 1168 155
rect 1172 154 1173 155
rect 1223 155 1229 156
rect 1172 152 1198 154
rect 1172 151 1173 152
rect 1167 150 1173 151
rect 1094 145 1100 146
rect 1094 141 1095 145
rect 1099 141 1100 145
rect 1094 140 1100 141
rect 1150 145 1156 146
rect 1150 141 1151 145
rect 1155 141 1156 145
rect 1150 140 1156 141
rect 1111 139 1117 140
rect 1111 138 1112 139
rect 1084 136 1112 138
rect 1055 134 1061 135
rect 1111 135 1112 136
rect 1116 135 1117 139
rect 1111 134 1117 135
rect 1167 139 1173 140
rect 1167 135 1168 139
rect 1172 138 1173 139
rect 1186 139 1192 140
rect 1186 138 1187 139
rect 1172 136 1187 138
rect 1172 135 1173 136
rect 1167 134 1173 135
rect 1186 135 1187 136
rect 1191 135 1192 139
rect 1196 138 1198 152
rect 1223 151 1224 155
rect 1228 154 1229 155
rect 1271 155 1277 156
rect 1228 152 1250 154
rect 1228 151 1229 152
rect 1223 150 1229 151
rect 1206 145 1212 146
rect 1206 141 1207 145
rect 1211 141 1212 145
rect 1206 140 1212 141
rect 1223 139 1229 140
rect 1223 138 1224 139
rect 1196 136 1224 138
rect 1186 134 1192 135
rect 1223 135 1224 136
rect 1228 135 1229 139
rect 1248 138 1250 152
rect 1271 151 1272 155
rect 1276 154 1277 155
rect 1314 155 1325 156
rect 1276 152 1298 154
rect 1276 151 1277 152
rect 1271 150 1277 151
rect 1254 145 1260 146
rect 1254 141 1255 145
rect 1259 141 1260 145
rect 1254 140 1260 141
rect 1271 139 1277 140
rect 1271 138 1272 139
rect 1248 136 1272 138
rect 1223 134 1229 135
rect 1271 135 1272 136
rect 1276 135 1277 139
rect 1296 138 1298 152
rect 1314 151 1315 155
rect 1319 151 1320 155
rect 1324 151 1325 155
rect 1314 150 1325 151
rect 1362 155 1373 156
rect 1362 151 1363 155
rect 1367 151 1368 155
rect 1372 151 1373 155
rect 1415 155 1421 156
rect 1415 154 1416 155
rect 1362 150 1373 151
rect 1392 152 1416 154
rect 1302 145 1308 146
rect 1302 141 1303 145
rect 1307 141 1308 145
rect 1302 140 1308 141
rect 1350 145 1356 146
rect 1350 141 1351 145
rect 1355 141 1356 145
rect 1350 140 1356 141
rect 1319 139 1325 140
rect 1319 138 1320 139
rect 1296 136 1320 138
rect 1271 134 1277 135
rect 1319 135 1320 136
rect 1324 135 1325 139
rect 1319 134 1325 135
rect 1367 139 1373 140
rect 1367 135 1368 139
rect 1372 138 1373 139
rect 1392 138 1394 152
rect 1415 151 1416 152
rect 1420 151 1421 155
rect 1471 155 1477 156
rect 1471 154 1472 155
rect 1415 150 1421 151
rect 1444 152 1472 154
rect 1398 145 1404 146
rect 1398 141 1399 145
rect 1403 141 1404 145
rect 1398 140 1404 141
rect 1372 136 1394 138
rect 1415 139 1421 140
rect 1372 135 1373 136
rect 1367 134 1373 135
rect 1415 135 1416 139
rect 1420 138 1421 139
rect 1444 138 1446 152
rect 1471 151 1472 152
rect 1476 151 1477 155
rect 1471 150 1477 151
rect 1527 155 1533 156
rect 1527 151 1528 155
rect 1532 154 1533 155
rect 1558 155 1565 156
rect 1532 152 1554 154
rect 1532 151 1533 152
rect 1527 150 1533 151
rect 1454 145 1460 146
rect 1454 141 1455 145
rect 1459 141 1460 145
rect 1454 140 1460 141
rect 1510 145 1516 146
rect 1510 141 1511 145
rect 1515 141 1516 145
rect 1510 140 1516 141
rect 1542 145 1548 146
rect 1542 141 1543 145
rect 1547 141 1548 145
rect 1542 140 1548 141
rect 1420 136 1446 138
rect 1471 139 1477 140
rect 1420 135 1421 136
rect 1415 134 1421 135
rect 1471 135 1472 139
rect 1476 138 1477 139
rect 1486 139 1492 140
rect 1486 138 1487 139
rect 1476 136 1487 138
rect 1476 135 1477 136
rect 1471 134 1477 135
rect 1486 135 1487 136
rect 1491 135 1492 139
rect 1486 134 1492 135
rect 1526 139 1533 140
rect 1526 135 1527 139
rect 1532 135 1533 139
rect 1552 138 1554 152
rect 1558 151 1559 155
rect 1564 151 1565 155
rect 1558 150 1565 151
rect 1582 144 1588 145
rect 1582 140 1583 144
rect 1587 140 1588 144
rect 1559 139 1565 140
rect 1582 139 1588 140
rect 1559 138 1560 139
rect 1552 136 1560 138
rect 1526 134 1533 135
rect 1559 135 1560 136
rect 1564 135 1565 139
rect 1559 134 1565 135
rect 1106 131 1112 132
rect 1106 130 1107 131
rect 836 128 1107 130
rect 543 127 544 128
rect 538 126 544 127
rect 1106 127 1107 128
rect 1111 127 1112 131
rect 1106 126 1112 127
rect 562 123 568 124
rect 562 122 563 123
rect 480 120 563 122
rect 151 115 160 116
rect 110 112 116 113
rect 110 108 111 112
rect 115 108 116 112
rect 110 107 116 108
rect 134 111 140 112
rect 134 107 135 111
rect 139 107 140 111
rect 151 111 152 115
rect 159 111 160 115
rect 183 115 189 116
rect 183 114 184 115
rect 176 112 184 114
rect 151 110 160 111
rect 166 111 172 112
rect 134 106 140 107
rect 166 107 167 111
rect 171 107 172 111
rect 166 106 172 107
rect 176 102 178 112
rect 183 111 184 112
rect 188 111 189 115
rect 215 115 221 116
rect 215 114 216 115
rect 208 112 216 114
rect 183 110 189 111
rect 198 111 204 112
rect 198 107 199 111
rect 203 107 204 111
rect 198 106 204 107
rect 208 102 210 112
rect 215 111 216 112
rect 220 111 221 115
rect 247 115 253 116
rect 247 114 248 115
rect 240 112 248 114
rect 215 110 221 111
rect 230 111 236 112
rect 230 107 231 111
rect 235 107 236 111
rect 230 106 236 107
rect 240 102 242 112
rect 247 111 248 112
rect 252 111 253 115
rect 279 115 285 116
rect 279 114 280 115
rect 272 112 280 114
rect 247 110 253 111
rect 262 111 268 112
rect 262 107 263 111
rect 267 107 268 111
rect 262 106 268 107
rect 272 102 274 112
rect 279 111 280 112
rect 284 111 285 115
rect 311 115 317 116
rect 311 114 312 115
rect 304 112 312 114
rect 279 110 285 111
rect 294 111 300 112
rect 294 107 295 111
rect 299 107 300 111
rect 294 106 300 107
rect 304 102 306 112
rect 311 111 312 112
rect 316 111 317 115
rect 343 115 349 116
rect 343 114 344 115
rect 336 112 344 114
rect 311 110 317 111
rect 326 111 332 112
rect 326 107 327 111
rect 331 107 332 111
rect 326 106 332 107
rect 336 102 338 112
rect 343 111 344 112
rect 348 111 349 115
rect 375 115 381 116
rect 375 114 376 115
rect 368 112 376 114
rect 343 110 349 111
rect 358 111 364 112
rect 358 107 359 111
rect 363 107 364 111
rect 358 106 364 107
rect 368 102 370 112
rect 375 111 376 112
rect 380 111 381 115
rect 407 115 413 116
rect 407 114 408 115
rect 400 112 408 114
rect 375 110 381 111
rect 390 111 396 112
rect 390 107 391 111
rect 395 107 396 111
rect 390 106 396 107
rect 400 102 402 112
rect 407 111 408 112
rect 412 111 413 115
rect 439 115 445 116
rect 439 114 440 115
rect 432 112 440 114
rect 407 110 413 111
rect 422 111 428 112
rect 422 107 423 111
rect 427 107 428 111
rect 422 106 428 107
rect 432 102 434 112
rect 439 111 440 112
rect 444 111 445 115
rect 471 115 477 116
rect 439 110 445 111
rect 454 111 460 112
rect 454 107 455 111
rect 459 107 460 111
rect 471 111 472 115
rect 476 114 477 115
rect 480 114 482 120
rect 562 119 563 120
rect 567 119 568 123
rect 562 118 568 119
rect 967 123 973 124
rect 967 119 968 123
rect 972 122 973 123
rect 1314 123 1320 124
rect 1314 122 1315 123
rect 972 120 1042 122
rect 972 119 973 120
rect 967 118 973 119
rect 503 115 509 116
rect 503 114 504 115
rect 476 112 482 114
rect 496 112 504 114
rect 476 111 477 112
rect 471 110 477 111
rect 486 111 492 112
rect 454 106 460 107
rect 486 107 487 111
rect 491 107 492 111
rect 486 106 492 107
rect 496 102 498 112
rect 503 111 504 112
rect 508 111 509 115
rect 535 115 541 116
rect 535 114 536 115
rect 528 112 536 114
rect 503 110 509 111
rect 518 111 524 112
rect 518 107 519 111
rect 523 107 524 111
rect 518 106 524 107
rect 528 102 530 112
rect 535 111 536 112
rect 540 111 541 115
rect 567 115 573 116
rect 535 110 541 111
rect 550 111 556 112
rect 550 107 551 111
rect 555 107 556 111
rect 567 111 568 115
rect 572 114 573 115
rect 599 115 605 116
rect 572 112 578 114
rect 572 111 573 112
rect 567 110 573 111
rect 550 106 556 107
rect 153 100 178 102
rect 196 100 210 102
rect 228 100 242 102
rect 260 100 274 102
rect 292 100 306 102
rect 324 100 338 102
rect 356 100 370 102
rect 388 100 402 102
rect 420 100 434 102
rect 484 100 498 102
rect 516 100 530 102
rect 576 102 578 112
rect 582 111 588 112
rect 582 107 583 111
rect 587 107 588 111
rect 599 111 600 115
rect 604 114 605 115
rect 631 115 637 116
rect 604 112 610 114
rect 604 111 605 112
rect 599 110 605 111
rect 582 106 588 107
rect 608 102 610 112
rect 614 111 620 112
rect 614 107 615 111
rect 619 107 620 111
rect 631 111 632 115
rect 636 114 637 115
rect 663 115 669 116
rect 636 112 642 114
rect 636 111 637 112
rect 631 110 637 111
rect 614 106 620 107
rect 624 104 634 106
rect 624 102 626 104
rect 632 102 634 104
rect 640 102 642 112
rect 646 111 652 112
rect 646 107 647 111
rect 651 107 652 111
rect 663 111 664 115
rect 668 114 669 115
rect 695 115 701 116
rect 668 112 674 114
rect 668 111 669 112
rect 663 110 669 111
rect 646 106 652 107
rect 672 102 674 112
rect 678 111 684 112
rect 678 107 679 111
rect 683 107 684 111
rect 695 111 696 115
rect 700 114 701 115
rect 727 115 733 116
rect 700 112 706 114
rect 700 111 701 112
rect 695 110 701 111
rect 678 106 684 107
rect 704 102 706 112
rect 710 111 716 112
rect 710 107 711 111
rect 715 107 716 111
rect 727 111 728 115
rect 732 114 733 115
rect 759 115 765 116
rect 732 112 738 114
rect 732 111 733 112
rect 727 110 733 111
rect 710 106 716 107
rect 736 102 738 112
rect 742 111 748 112
rect 742 107 743 111
rect 747 107 748 111
rect 759 111 760 115
rect 764 114 765 115
rect 791 115 797 116
rect 764 112 770 114
rect 764 111 765 112
rect 759 110 765 111
rect 742 106 748 107
rect 768 102 770 112
rect 774 111 780 112
rect 774 107 775 111
rect 779 107 780 111
rect 791 111 792 115
rect 796 114 797 115
rect 823 115 829 116
rect 796 112 802 114
rect 796 111 797 112
rect 791 110 797 111
rect 774 106 780 107
rect 800 102 802 112
rect 806 111 812 112
rect 806 107 807 111
rect 811 107 812 111
rect 823 111 824 115
rect 828 114 829 115
rect 855 115 861 116
rect 828 112 834 114
rect 828 111 829 112
rect 823 110 829 111
rect 806 106 812 107
rect 832 102 834 112
rect 838 111 844 112
rect 838 107 839 111
rect 843 107 844 111
rect 855 111 856 115
rect 860 114 861 115
rect 887 115 893 116
rect 860 112 866 114
rect 860 111 861 112
rect 855 110 861 111
rect 838 106 844 107
rect 864 102 866 112
rect 870 111 876 112
rect 870 107 871 111
rect 875 107 876 111
rect 887 111 888 115
rect 892 114 893 115
rect 919 115 925 116
rect 892 112 898 114
rect 892 111 893 112
rect 887 110 893 111
rect 870 106 876 107
rect 896 102 898 112
rect 902 111 908 112
rect 902 107 903 111
rect 907 107 908 111
rect 919 111 920 115
rect 924 114 925 115
rect 959 115 965 116
rect 924 112 938 114
rect 924 111 925 112
rect 919 110 925 111
rect 902 106 908 107
rect 936 102 938 112
rect 942 111 948 112
rect 942 107 943 111
rect 947 107 948 111
rect 959 111 960 115
rect 964 114 965 115
rect 999 115 1005 116
rect 964 112 978 114
rect 964 111 965 112
rect 959 110 965 111
rect 942 106 948 107
rect 976 102 978 112
rect 982 111 988 112
rect 982 107 983 111
rect 987 107 988 111
rect 999 111 1000 115
rect 1004 114 1005 115
rect 1022 115 1028 116
rect 1022 114 1023 115
rect 1004 112 1023 114
rect 1004 111 1005 112
rect 999 110 1005 111
rect 1022 111 1023 112
rect 1027 111 1028 115
rect 1040 114 1042 120
rect 1193 120 1315 122
rect 1193 116 1195 120
rect 1314 119 1315 120
rect 1319 119 1320 123
rect 1314 118 1320 119
rect 1047 115 1053 116
rect 1047 114 1048 115
rect 1040 112 1048 114
rect 1022 110 1028 111
rect 1030 111 1036 112
rect 982 106 988 107
rect 1030 107 1031 111
rect 1035 107 1036 111
rect 1047 111 1048 112
rect 1052 111 1053 115
rect 1095 115 1101 116
rect 1095 114 1096 115
rect 1088 112 1096 114
rect 1047 110 1053 111
rect 1078 111 1084 112
rect 1030 106 1036 107
rect 1078 107 1079 111
rect 1083 107 1084 111
rect 1078 106 1084 107
rect 1088 102 1090 112
rect 1095 111 1096 112
rect 1100 111 1101 115
rect 1143 115 1149 116
rect 1143 114 1144 115
rect 1136 112 1144 114
rect 1095 110 1101 111
rect 1126 111 1132 112
rect 1126 107 1127 111
rect 1131 107 1132 111
rect 1126 106 1132 107
rect 1136 102 1138 112
rect 1143 111 1144 112
rect 1148 111 1149 115
rect 1191 115 1197 116
rect 1143 110 1149 111
rect 1174 111 1180 112
rect 1174 107 1175 111
rect 1179 107 1180 111
rect 1191 111 1192 115
rect 1196 111 1197 115
rect 1239 115 1245 116
rect 1239 114 1240 115
rect 1232 112 1240 114
rect 1191 110 1197 111
rect 1222 111 1228 112
rect 1174 106 1180 107
rect 1222 107 1223 111
rect 1227 107 1228 111
rect 1222 106 1228 107
rect 1232 102 1234 112
rect 1239 111 1240 112
rect 1244 111 1245 115
rect 1279 115 1285 116
rect 1279 114 1280 115
rect 1272 112 1280 114
rect 1239 110 1245 111
rect 1262 111 1268 112
rect 1262 107 1263 111
rect 1267 107 1268 111
rect 1262 106 1268 107
rect 1272 102 1274 112
rect 1279 111 1280 112
rect 1284 111 1285 115
rect 1319 115 1325 116
rect 1319 114 1320 115
rect 1312 112 1320 114
rect 1279 110 1285 111
rect 1302 111 1308 112
rect 1302 107 1303 111
rect 1307 107 1308 111
rect 1302 106 1308 107
rect 1312 102 1314 112
rect 1319 111 1320 112
rect 1324 111 1325 115
rect 1359 115 1365 116
rect 1359 114 1360 115
rect 1352 112 1360 114
rect 1319 110 1325 111
rect 1342 111 1348 112
rect 1342 107 1343 111
rect 1347 107 1348 111
rect 1342 106 1348 107
rect 1352 102 1354 112
rect 1359 111 1360 112
rect 1364 111 1365 115
rect 1399 115 1405 116
rect 1399 114 1400 115
rect 1392 112 1400 114
rect 1359 110 1365 111
rect 1382 111 1388 112
rect 1382 107 1383 111
rect 1387 107 1388 111
rect 1382 106 1388 107
rect 1392 102 1394 112
rect 1399 111 1400 112
rect 1404 111 1405 115
rect 1439 115 1445 116
rect 1439 114 1440 115
rect 1432 112 1440 114
rect 1399 110 1405 111
rect 1422 111 1428 112
rect 1422 107 1423 111
rect 1427 107 1428 111
rect 1422 106 1428 107
rect 1432 102 1434 112
rect 1439 111 1440 112
rect 1444 111 1445 115
rect 1487 115 1493 116
rect 1487 114 1488 115
rect 1480 112 1488 114
rect 1439 110 1445 111
rect 1470 111 1476 112
rect 1470 107 1471 111
rect 1475 107 1476 111
rect 1470 106 1476 107
rect 1480 102 1482 112
rect 1487 111 1488 112
rect 1492 111 1493 115
rect 1527 115 1533 116
rect 1487 110 1493 111
rect 1510 111 1516 112
rect 1510 107 1511 111
rect 1515 107 1516 111
rect 1527 111 1528 115
rect 1532 114 1533 115
rect 1558 115 1565 116
rect 1532 112 1538 114
rect 1532 111 1533 112
rect 1527 110 1533 111
rect 1510 106 1516 107
rect 576 100 594 102
rect 608 100 626 102
rect 631 101 637 102
rect 151 99 157 100
rect 110 95 116 96
rect 110 91 111 95
rect 115 91 116 95
rect 151 95 152 99
rect 156 95 157 99
rect 151 94 157 95
rect 183 99 189 100
rect 183 95 184 99
rect 188 98 189 99
rect 196 98 198 100
rect 188 96 198 98
rect 215 99 221 100
rect 188 95 189 96
rect 183 94 189 95
rect 215 95 216 99
rect 220 98 221 99
rect 228 98 230 100
rect 220 96 230 98
rect 247 99 253 100
rect 220 95 221 96
rect 215 94 221 95
rect 247 95 248 99
rect 252 98 253 99
rect 260 98 262 100
rect 252 96 262 98
rect 279 99 285 100
rect 252 95 253 96
rect 247 94 253 95
rect 279 95 280 99
rect 284 98 285 99
rect 292 98 294 100
rect 284 96 294 98
rect 311 99 317 100
rect 284 95 285 96
rect 279 94 285 95
rect 311 95 312 99
rect 316 98 317 99
rect 324 98 326 100
rect 316 96 326 98
rect 343 99 349 100
rect 316 95 317 96
rect 311 94 317 95
rect 343 95 344 99
rect 348 98 349 99
rect 356 98 358 100
rect 348 96 358 98
rect 375 99 381 100
rect 348 95 349 96
rect 343 94 349 95
rect 375 95 376 99
rect 380 98 381 99
rect 388 98 390 100
rect 380 96 390 98
rect 407 99 413 100
rect 380 95 381 96
rect 375 94 381 95
rect 407 95 408 99
rect 412 98 413 99
rect 420 98 422 100
rect 412 96 422 98
rect 438 99 445 100
rect 412 95 413 96
rect 407 94 413 95
rect 438 95 439 99
rect 444 95 445 99
rect 438 94 445 95
rect 471 99 477 100
rect 471 95 472 99
rect 476 98 477 99
rect 484 98 486 100
rect 476 96 486 98
rect 503 99 509 100
rect 476 95 477 96
rect 471 94 477 95
rect 503 95 504 99
rect 508 98 509 99
rect 516 98 518 100
rect 508 96 518 98
rect 535 99 544 100
rect 508 95 509 96
rect 503 94 509 95
rect 535 95 536 99
rect 543 95 544 99
rect 535 94 544 95
rect 562 99 573 100
rect 562 95 563 99
rect 567 95 568 99
rect 572 95 573 99
rect 592 98 594 100
rect 599 99 605 100
rect 599 98 600 99
rect 592 96 600 98
rect 562 94 573 95
rect 599 95 600 96
rect 604 95 605 99
rect 631 97 632 101
rect 636 97 637 101
rect 640 100 658 102
rect 672 100 690 102
rect 704 100 722 102
rect 736 100 754 102
rect 768 100 786 102
rect 800 100 818 102
rect 832 100 850 102
rect 864 100 882 102
rect 896 100 914 102
rect 936 100 954 102
rect 976 100 994 102
rect 1072 100 1090 102
rect 1097 100 1138 102
rect 1193 100 1234 102
rect 1260 100 1274 102
rect 1300 100 1314 102
rect 1321 100 1354 102
rect 1380 100 1394 102
rect 1420 100 1434 102
rect 1464 100 1482 102
rect 1536 102 1538 112
rect 1542 111 1548 112
rect 1542 107 1543 111
rect 1547 107 1548 111
rect 1558 111 1559 115
rect 1564 111 1565 115
rect 1558 110 1565 111
rect 1582 112 1588 113
rect 1582 108 1583 112
rect 1587 108 1588 112
rect 1582 107 1588 108
rect 1542 106 1548 107
rect 1536 100 1563 102
rect 631 96 637 97
rect 656 98 658 100
rect 663 99 669 100
rect 663 98 664 99
rect 656 96 664 98
rect 599 94 605 95
rect 663 95 664 96
rect 668 95 669 99
rect 688 98 690 100
rect 695 99 701 100
rect 695 98 696 99
rect 688 96 696 98
rect 663 94 669 95
rect 695 95 696 96
rect 700 95 701 99
rect 720 98 722 100
rect 727 99 733 100
rect 727 98 728 99
rect 720 96 728 98
rect 695 94 701 95
rect 727 95 728 96
rect 732 95 733 99
rect 752 98 754 100
rect 759 99 765 100
rect 759 98 760 99
rect 752 96 760 98
rect 727 94 733 95
rect 759 95 760 96
rect 764 95 765 99
rect 784 98 786 100
rect 791 99 797 100
rect 791 98 792 99
rect 784 96 792 98
rect 759 94 765 95
rect 791 95 792 96
rect 796 95 797 99
rect 816 98 818 100
rect 823 99 829 100
rect 823 98 824 99
rect 816 96 824 98
rect 791 94 797 95
rect 823 95 824 96
rect 828 95 829 99
rect 848 98 850 100
rect 855 99 861 100
rect 855 98 856 99
rect 848 96 856 98
rect 823 94 829 95
rect 855 95 856 96
rect 860 95 861 99
rect 880 98 882 100
rect 887 99 893 100
rect 887 98 888 99
rect 880 96 888 98
rect 855 94 861 95
rect 887 95 888 96
rect 892 95 893 99
rect 912 98 914 100
rect 919 99 925 100
rect 919 98 920 99
rect 912 96 920 98
rect 887 94 893 95
rect 919 95 920 96
rect 924 95 925 99
rect 952 98 954 100
rect 959 99 965 100
rect 959 98 960 99
rect 952 96 960 98
rect 919 94 925 95
rect 959 95 960 96
rect 964 95 965 99
rect 992 98 994 100
rect 999 99 1005 100
rect 999 98 1000 99
rect 992 96 1000 98
rect 959 94 965 95
rect 999 95 1000 96
rect 1004 95 1005 99
rect 999 94 1005 95
rect 1047 99 1053 100
rect 1047 95 1048 99
rect 1052 98 1053 99
rect 1072 98 1074 100
rect 1052 96 1074 98
rect 1095 99 1101 100
rect 1052 95 1053 96
rect 1047 94 1053 95
rect 1095 95 1096 99
rect 1100 95 1101 99
rect 1143 99 1149 100
rect 1143 98 1144 99
rect 1095 94 1101 95
rect 1136 96 1144 98
rect 110 90 116 91
rect 134 93 140 94
rect 134 89 135 93
rect 139 89 140 93
rect 134 88 140 89
rect 166 93 172 94
rect 166 89 167 93
rect 171 89 172 93
rect 166 88 172 89
rect 198 93 204 94
rect 198 89 199 93
rect 203 89 204 93
rect 198 88 204 89
rect 230 93 236 94
rect 230 89 231 93
rect 235 89 236 93
rect 230 88 236 89
rect 262 93 268 94
rect 262 89 263 93
rect 267 89 268 93
rect 262 88 268 89
rect 294 93 300 94
rect 294 89 295 93
rect 299 89 300 93
rect 294 88 300 89
rect 326 93 332 94
rect 326 89 327 93
rect 331 89 332 93
rect 326 88 332 89
rect 358 93 364 94
rect 358 89 359 93
rect 363 89 364 93
rect 358 88 364 89
rect 390 93 396 94
rect 390 89 391 93
rect 395 89 396 93
rect 390 88 396 89
rect 422 93 428 94
rect 422 89 423 93
rect 427 89 428 93
rect 422 88 428 89
rect 454 93 460 94
rect 454 89 455 93
rect 459 89 460 93
rect 454 88 460 89
rect 486 93 492 94
rect 486 89 487 93
rect 491 89 492 93
rect 486 88 492 89
rect 518 93 524 94
rect 518 89 519 93
rect 523 89 524 93
rect 518 88 524 89
rect 550 93 556 94
rect 550 89 551 93
rect 555 89 556 93
rect 550 88 556 89
rect 582 93 588 94
rect 582 89 583 93
rect 587 89 588 93
rect 582 88 588 89
rect 614 93 620 94
rect 614 89 615 93
rect 619 89 620 93
rect 614 88 620 89
rect 646 93 652 94
rect 646 89 647 93
rect 651 89 652 93
rect 646 88 652 89
rect 678 93 684 94
rect 678 89 679 93
rect 683 89 684 93
rect 678 88 684 89
rect 710 93 716 94
rect 710 89 711 93
rect 715 89 716 93
rect 710 88 716 89
rect 742 93 748 94
rect 742 89 743 93
rect 747 89 748 93
rect 742 88 748 89
rect 774 93 780 94
rect 774 89 775 93
rect 779 89 780 93
rect 774 88 780 89
rect 806 93 812 94
rect 806 89 807 93
rect 811 89 812 93
rect 806 88 812 89
rect 838 93 844 94
rect 838 89 839 93
rect 843 89 844 93
rect 838 88 844 89
rect 870 93 876 94
rect 870 89 871 93
rect 875 89 876 93
rect 870 88 876 89
rect 902 93 908 94
rect 902 89 903 93
rect 907 89 908 93
rect 902 88 908 89
rect 942 93 948 94
rect 942 89 943 93
rect 947 89 948 93
rect 942 88 948 89
rect 982 93 988 94
rect 982 89 983 93
rect 987 89 988 93
rect 982 88 988 89
rect 1030 93 1036 94
rect 1030 89 1031 93
rect 1035 89 1036 93
rect 1030 88 1036 89
rect 1078 93 1084 94
rect 1078 89 1079 93
rect 1083 89 1084 93
rect 1078 88 1084 89
rect 1126 93 1132 94
rect 1126 89 1127 93
rect 1131 89 1132 93
rect 1126 88 1132 89
rect 1022 87 1028 88
rect 1022 83 1023 87
rect 1027 86 1028 87
rect 1136 86 1138 96
rect 1143 95 1144 96
rect 1148 95 1149 99
rect 1143 94 1149 95
rect 1191 99 1197 100
rect 1191 95 1192 99
rect 1196 95 1197 99
rect 1191 94 1197 95
rect 1239 99 1245 100
rect 1239 95 1240 99
rect 1244 98 1245 99
rect 1260 98 1262 100
rect 1244 96 1262 98
rect 1279 99 1285 100
rect 1244 95 1245 96
rect 1239 94 1245 95
rect 1279 95 1280 99
rect 1284 98 1285 99
rect 1300 98 1302 100
rect 1284 96 1302 98
rect 1319 99 1325 100
rect 1284 95 1285 96
rect 1279 94 1285 95
rect 1319 95 1320 99
rect 1324 95 1325 99
rect 1319 94 1325 95
rect 1359 99 1365 100
rect 1359 95 1360 99
rect 1364 98 1365 99
rect 1380 98 1382 100
rect 1364 96 1382 98
rect 1399 99 1405 100
rect 1364 95 1365 96
rect 1359 94 1365 95
rect 1399 95 1400 99
rect 1404 98 1405 99
rect 1420 98 1422 100
rect 1404 96 1422 98
rect 1439 99 1445 100
rect 1404 95 1405 96
rect 1399 94 1405 95
rect 1439 95 1440 99
rect 1444 98 1445 99
rect 1464 98 1466 100
rect 1444 96 1466 98
rect 1486 99 1493 100
rect 1444 95 1445 96
rect 1439 94 1445 95
rect 1486 95 1487 99
rect 1492 95 1493 99
rect 1486 94 1493 95
rect 1559 99 1565 100
rect 1559 95 1560 99
rect 1564 95 1565 99
rect 1559 94 1565 95
rect 1582 95 1588 96
rect 1174 93 1180 94
rect 1174 89 1175 93
rect 1179 89 1180 93
rect 1174 88 1180 89
rect 1222 93 1228 94
rect 1222 89 1223 93
rect 1227 89 1228 93
rect 1222 88 1228 89
rect 1262 93 1268 94
rect 1262 89 1263 93
rect 1267 89 1268 93
rect 1262 88 1268 89
rect 1302 93 1308 94
rect 1302 89 1303 93
rect 1307 89 1308 93
rect 1302 88 1308 89
rect 1342 93 1348 94
rect 1342 89 1343 93
rect 1347 89 1348 93
rect 1342 88 1348 89
rect 1382 93 1388 94
rect 1382 89 1383 93
rect 1387 89 1388 93
rect 1382 88 1388 89
rect 1422 93 1428 94
rect 1422 89 1423 93
rect 1427 89 1428 93
rect 1422 88 1428 89
rect 1470 93 1476 94
rect 1470 89 1471 93
rect 1475 89 1476 93
rect 1470 88 1476 89
rect 1510 93 1516 94
rect 1510 89 1511 93
rect 1515 89 1516 93
rect 1510 88 1516 89
rect 1542 93 1548 94
rect 1542 89 1543 93
rect 1547 89 1548 93
rect 1582 91 1583 95
rect 1587 91 1588 95
rect 1582 90 1588 91
rect 1542 88 1548 89
rect 1027 84 1138 86
rect 1027 83 1028 84
rect 1022 82 1028 83
<< m3c >>
rect 111 1641 115 1645
rect 135 1643 139 1647
rect 167 1643 171 1647
rect 199 1643 203 1647
rect 1583 1641 1587 1645
rect 151 1635 152 1639
rect 152 1635 155 1639
rect 111 1624 115 1628
rect 135 1625 139 1629
rect 167 1625 171 1629
rect 199 1625 203 1629
rect 1583 1624 1587 1628
rect 111 1604 115 1608
rect 135 1603 139 1607
rect 151 1607 152 1611
rect 152 1607 155 1611
rect 175 1603 179 1607
rect 239 1603 243 1607
rect 295 1603 299 1607
rect 351 1603 355 1607
rect 399 1607 403 1611
rect 407 1603 411 1607
rect 455 1603 459 1607
rect 503 1603 507 1607
rect 551 1603 555 1607
rect 599 1603 603 1607
rect 647 1603 651 1607
rect 695 1603 699 1607
rect 743 1603 747 1607
rect 791 1603 795 1607
rect 831 1607 835 1611
rect 839 1603 843 1607
rect 887 1603 891 1607
rect 935 1603 939 1607
rect 991 1603 995 1607
rect 1047 1603 1051 1607
rect 1095 1603 1099 1607
rect 1143 1603 1147 1607
rect 1191 1603 1195 1607
rect 1203 1607 1207 1611
rect 1239 1603 1243 1607
rect 1287 1603 1291 1607
rect 1327 1603 1331 1607
rect 1367 1603 1371 1607
rect 1407 1603 1411 1607
rect 1447 1603 1451 1607
rect 1479 1603 1483 1607
rect 1511 1603 1515 1607
rect 1543 1603 1547 1607
rect 1583 1604 1587 1608
rect 111 1587 115 1591
rect 1159 1591 1160 1595
rect 1160 1591 1163 1595
rect 135 1585 139 1589
rect 175 1585 179 1589
rect 239 1585 243 1589
rect 295 1585 299 1589
rect 195 1579 199 1583
rect 351 1585 355 1589
rect 407 1585 411 1589
rect 455 1585 459 1589
rect 503 1585 507 1589
rect 551 1585 555 1589
rect 599 1585 603 1589
rect 647 1585 651 1589
rect 695 1585 699 1589
rect 743 1585 747 1589
rect 399 1579 403 1583
rect 111 1569 115 1573
rect 175 1571 179 1575
rect 215 1571 219 1575
rect 255 1571 259 1575
rect 295 1571 299 1575
rect 343 1571 347 1575
rect 391 1571 395 1575
rect 439 1571 443 1575
rect 487 1571 491 1575
rect 535 1571 539 1575
rect 111 1552 115 1556
rect 175 1553 179 1557
rect 195 1547 196 1551
rect 196 1547 199 1551
rect 247 1563 251 1567
rect 215 1553 219 1557
rect 255 1553 259 1557
rect 295 1553 299 1557
rect 343 1553 347 1557
rect 391 1553 395 1557
rect 439 1553 443 1557
rect 791 1585 795 1589
rect 839 1585 843 1589
rect 887 1585 891 1589
rect 935 1585 939 1589
rect 991 1585 995 1589
rect 1047 1585 1051 1589
rect 1095 1585 1099 1589
rect 1143 1585 1147 1589
rect 1191 1585 1195 1589
rect 1239 1585 1243 1589
rect 1287 1585 1291 1589
rect 1327 1585 1331 1589
rect 1367 1585 1371 1589
rect 1407 1585 1411 1589
rect 1447 1585 1451 1589
rect 1479 1585 1483 1589
rect 1511 1585 1515 1589
rect 1543 1585 1547 1589
rect 1499 1579 1503 1583
rect 1583 1587 1587 1591
rect 583 1571 587 1575
rect 639 1571 643 1575
rect 703 1571 707 1575
rect 775 1571 779 1575
rect 855 1571 859 1575
rect 935 1571 939 1575
rect 1015 1571 1019 1575
rect 1087 1571 1091 1575
rect 1159 1571 1163 1575
rect 1239 1571 1243 1575
rect 1319 1571 1323 1575
rect 487 1553 491 1557
rect 535 1553 539 1557
rect 583 1553 587 1557
rect 639 1553 643 1557
rect 703 1553 707 1557
rect 767 1563 771 1567
rect 831 1563 835 1567
rect 775 1553 779 1557
rect 855 1553 859 1557
rect 987 1563 991 1567
rect 935 1553 939 1557
rect 1015 1553 1019 1557
rect 1087 1553 1091 1557
rect 915 1547 919 1551
rect 1203 1563 1207 1567
rect 1159 1553 1163 1557
rect 1151 1547 1155 1551
rect 1239 1553 1243 1557
rect 1399 1571 1403 1575
rect 1479 1571 1483 1575
rect 1543 1571 1547 1575
rect 1583 1569 1587 1573
rect 1319 1553 1323 1557
rect 1327 1547 1331 1551
rect 1399 1553 1403 1557
rect 1479 1553 1483 1557
rect 1499 1553 1503 1555
rect 1499 1551 1500 1553
rect 1500 1551 1503 1553
rect 1543 1553 1547 1557
rect 1559 1563 1560 1567
rect 1560 1563 1563 1567
rect 1583 1552 1587 1556
rect 111 1532 115 1536
rect 159 1531 163 1535
rect 207 1531 211 1535
rect 247 1539 251 1543
rect 255 1531 259 1535
rect 311 1531 315 1535
rect 359 1531 363 1535
rect 371 1535 375 1539
rect 415 1531 419 1535
rect 111 1515 115 1519
rect 175 1519 176 1523
rect 176 1519 179 1523
rect 471 1531 475 1535
rect 159 1513 163 1517
rect 207 1513 211 1517
rect 255 1513 259 1517
rect 311 1513 315 1517
rect 359 1513 363 1517
rect 415 1513 419 1517
rect 527 1531 531 1535
rect 583 1531 587 1535
rect 639 1531 643 1535
rect 695 1531 699 1535
rect 767 1539 771 1543
rect 759 1531 763 1535
rect 775 1531 779 1535
rect 823 1531 827 1535
rect 895 1531 899 1535
rect 967 1531 971 1535
rect 987 1535 988 1539
rect 988 1535 991 1539
rect 1039 1531 1043 1535
rect 1103 1531 1107 1535
rect 1167 1531 1171 1535
rect 1223 1535 1227 1539
rect 1231 1531 1235 1535
rect 1295 1531 1299 1535
rect 1359 1531 1363 1535
rect 1423 1531 1427 1535
rect 1439 1535 1440 1539
rect 1440 1535 1443 1539
rect 1495 1531 1499 1535
rect 1543 1531 1547 1535
rect 1559 1535 1560 1539
rect 1560 1535 1563 1539
rect 1583 1532 1587 1536
rect 915 1519 916 1523
rect 916 1519 919 1523
rect 1115 1519 1119 1523
rect 1327 1519 1331 1523
rect 471 1513 475 1517
rect 527 1513 531 1517
rect 583 1513 587 1517
rect 639 1513 643 1517
rect 695 1513 699 1517
rect 759 1513 763 1517
rect 823 1513 827 1517
rect 895 1513 899 1517
rect 967 1513 971 1517
rect 1039 1513 1043 1517
rect 1103 1513 1107 1517
rect 1167 1513 1171 1517
rect 1231 1513 1235 1517
rect 1295 1513 1299 1517
rect 1359 1513 1363 1517
rect 483 1507 487 1511
rect 111 1497 115 1501
rect 159 1499 163 1503
rect 207 1499 211 1503
rect 255 1499 259 1503
rect 303 1499 307 1503
rect 351 1499 355 1503
rect 407 1499 411 1503
rect 463 1499 467 1503
rect 527 1499 531 1503
rect 591 1499 595 1503
rect 111 1480 115 1484
rect 159 1481 163 1485
rect 175 1475 176 1479
rect 176 1475 179 1479
rect 219 1491 223 1495
rect 207 1481 211 1485
rect 255 1481 259 1485
rect 275 1475 276 1479
rect 276 1475 279 1479
rect 303 1481 307 1485
rect 371 1491 372 1495
rect 372 1491 375 1495
rect 351 1481 355 1485
rect 407 1481 411 1485
rect 463 1481 467 1485
rect 527 1481 531 1485
rect 1223 1507 1227 1511
rect 1511 1519 1512 1523
rect 1512 1519 1515 1523
rect 1423 1513 1427 1517
rect 1495 1513 1499 1517
rect 1543 1513 1547 1517
rect 1583 1515 1587 1519
rect 655 1499 659 1503
rect 719 1499 723 1503
rect 783 1499 787 1503
rect 855 1499 859 1503
rect 935 1499 939 1503
rect 1007 1499 1011 1503
rect 1079 1499 1083 1503
rect 1151 1499 1155 1503
rect 1215 1499 1219 1503
rect 1279 1499 1283 1503
rect 1351 1499 1355 1503
rect 1423 1499 1427 1503
rect 1495 1499 1499 1503
rect 1543 1499 1547 1503
rect 1583 1497 1587 1501
rect 591 1481 595 1485
rect 775 1491 779 1495
rect 655 1481 659 1485
rect 719 1481 723 1485
rect 783 1481 787 1485
rect 899 1491 903 1495
rect 855 1481 859 1485
rect 935 1481 939 1485
rect 835 1475 839 1479
rect 1007 1481 1011 1485
rect 1079 1481 1083 1485
rect 1151 1481 1155 1485
rect 1115 1475 1119 1479
rect 1215 1481 1219 1485
rect 111 1460 115 1464
rect 135 1459 139 1463
rect 183 1459 187 1463
rect 219 1463 223 1467
rect 231 1459 235 1463
rect 259 1459 263 1463
rect 287 1459 291 1463
rect 343 1459 347 1463
rect 399 1459 403 1463
rect 455 1459 459 1463
rect 483 1463 487 1467
rect 511 1459 515 1463
rect 575 1459 579 1463
rect 1279 1481 1283 1485
rect 1351 1481 1355 1485
rect 1439 1491 1440 1495
rect 1440 1491 1443 1495
rect 1423 1481 1427 1485
rect 1495 1481 1499 1485
rect 1511 1475 1512 1479
rect 1512 1475 1515 1479
rect 1559 1491 1560 1495
rect 1560 1491 1563 1495
rect 1543 1481 1547 1485
rect 1583 1480 1587 1484
rect 631 1459 635 1463
rect 687 1459 691 1463
rect 699 1463 703 1467
rect 751 1459 755 1463
rect 815 1459 819 1463
rect 879 1459 883 1463
rect 899 1463 900 1467
rect 900 1463 903 1467
rect 943 1459 947 1463
rect 1015 1459 1019 1463
rect 1087 1459 1091 1463
rect 1159 1459 1163 1463
rect 1175 1463 1176 1467
rect 1176 1463 1179 1467
rect 1239 1459 1243 1463
rect 1319 1459 1323 1463
rect 1399 1459 1403 1463
rect 1479 1459 1483 1463
rect 1543 1459 1547 1463
rect 1559 1463 1560 1467
rect 1560 1463 1563 1467
rect 1583 1460 1587 1464
rect 111 1443 115 1447
rect 151 1447 152 1451
rect 152 1447 155 1451
rect 135 1441 139 1445
rect 183 1441 187 1445
rect 231 1441 235 1445
rect 287 1441 291 1445
rect 343 1441 347 1445
rect 399 1441 403 1445
rect 275 1435 279 1439
rect 643 1447 647 1451
rect 835 1447 836 1451
rect 836 1447 839 1451
rect 1103 1447 1104 1451
rect 1104 1447 1107 1451
rect 1527 1447 1531 1451
rect 455 1441 459 1445
rect 511 1441 515 1445
rect 575 1441 579 1445
rect 631 1441 635 1445
rect 687 1441 691 1445
rect 751 1441 755 1445
rect 815 1441 819 1445
rect 879 1441 883 1445
rect 943 1441 947 1445
rect 1015 1441 1019 1445
rect 1087 1441 1091 1445
rect 1159 1441 1163 1445
rect 1239 1441 1243 1445
rect 1319 1441 1323 1445
rect 1399 1441 1403 1445
rect 1479 1441 1483 1445
rect 1543 1441 1547 1445
rect 1583 1443 1587 1447
rect 911 1435 915 1439
rect 111 1425 115 1429
rect 135 1427 139 1431
rect 183 1427 187 1431
rect 255 1427 259 1431
rect 327 1427 331 1431
rect 399 1427 403 1431
rect 471 1427 475 1431
rect 543 1427 547 1431
rect 615 1427 619 1431
rect 679 1427 683 1431
rect 743 1427 747 1431
rect 815 1427 819 1431
rect 879 1427 883 1431
rect 951 1427 955 1431
rect 1023 1427 1027 1431
rect 195 1419 199 1423
rect 111 1408 115 1412
rect 135 1409 139 1413
rect 151 1403 152 1407
rect 152 1403 155 1407
rect 183 1409 187 1413
rect 255 1409 259 1413
rect 263 1403 267 1407
rect 327 1409 331 1413
rect 399 1409 403 1413
rect 415 1419 416 1423
rect 416 1419 419 1423
rect 483 1419 487 1423
rect 471 1409 475 1413
rect 543 1409 547 1413
rect 699 1419 700 1423
rect 700 1419 703 1423
rect 615 1409 619 1413
rect 643 1407 647 1411
rect 679 1409 683 1413
rect 743 1409 747 1413
rect 815 1409 819 1413
rect 879 1409 883 1413
rect 951 1409 955 1413
rect 855 1403 859 1407
rect 1023 1409 1027 1413
rect 1363 1435 1367 1439
rect 1095 1427 1099 1431
rect 1159 1427 1163 1431
rect 1223 1427 1227 1431
rect 1287 1427 1291 1431
rect 1343 1427 1347 1431
rect 1399 1427 1403 1431
rect 1455 1427 1459 1431
rect 1511 1427 1515 1431
rect 1543 1427 1547 1431
rect 1583 1425 1587 1429
rect 1175 1419 1176 1423
rect 1176 1419 1179 1423
rect 1095 1409 1099 1413
rect 1159 1409 1163 1413
rect 1223 1409 1227 1413
rect 1287 1409 1291 1413
rect 1343 1409 1347 1413
rect 1307 1403 1308 1407
rect 1308 1403 1311 1407
rect 1363 1403 1364 1407
rect 1364 1403 1367 1407
rect 1399 1409 1403 1413
rect 1455 1409 1459 1413
rect 1495 1419 1499 1423
rect 1511 1409 1515 1413
rect 1543 1409 1547 1413
rect 1527 1403 1528 1407
rect 1528 1403 1531 1407
rect 1583 1408 1587 1412
rect 111 1388 115 1392
rect 135 1387 139 1391
rect 175 1387 179 1391
rect 195 1391 196 1395
rect 196 1391 199 1395
rect 247 1387 251 1391
rect 319 1387 323 1391
rect 391 1387 395 1391
rect 447 1391 451 1395
rect 455 1387 459 1391
rect 483 1391 487 1395
rect 519 1387 523 1391
rect 583 1387 587 1391
rect 647 1387 651 1391
rect 711 1387 715 1391
rect 775 1387 779 1391
rect 839 1387 843 1391
rect 895 1387 899 1391
rect 911 1391 912 1395
rect 912 1391 915 1395
rect 951 1387 955 1391
rect 999 1387 1003 1391
rect 1055 1387 1059 1391
rect 1103 1395 1107 1399
rect 1111 1387 1115 1391
rect 1175 1387 1179 1391
rect 1187 1391 1191 1395
rect 1239 1387 1243 1391
rect 1295 1387 1299 1391
rect 1351 1387 1355 1391
rect 1407 1391 1411 1395
rect 1415 1387 1419 1391
rect 1479 1387 1483 1391
rect 1495 1391 1496 1395
rect 1496 1391 1499 1395
rect 1543 1387 1547 1391
rect 1583 1388 1587 1392
rect 111 1371 115 1375
rect 151 1375 152 1379
rect 152 1375 155 1379
rect 263 1375 264 1379
rect 264 1375 267 1379
rect 855 1375 856 1379
rect 856 1375 859 1379
rect 1127 1375 1128 1379
rect 1128 1375 1131 1379
rect 1307 1375 1311 1379
rect 1463 1375 1467 1379
rect 135 1369 139 1373
rect 175 1369 179 1373
rect 247 1369 251 1373
rect 319 1369 323 1373
rect 391 1369 395 1373
rect 455 1369 459 1373
rect 519 1369 523 1373
rect 583 1369 587 1373
rect 647 1369 651 1373
rect 711 1369 715 1373
rect 775 1369 779 1373
rect 839 1369 843 1373
rect 895 1369 899 1373
rect 951 1369 955 1373
rect 999 1369 1003 1373
rect 1055 1369 1059 1373
rect 1111 1369 1115 1373
rect 1175 1369 1179 1373
rect 1239 1369 1243 1373
rect 1295 1369 1299 1373
rect 1351 1369 1355 1373
rect 1415 1369 1419 1373
rect 1479 1369 1483 1373
rect 1543 1369 1547 1373
rect 447 1363 451 1367
rect 111 1353 115 1357
rect 135 1355 139 1359
rect 167 1355 171 1359
rect 215 1355 219 1359
rect 303 1355 307 1359
rect 415 1355 419 1359
rect 527 1355 531 1359
rect 111 1336 115 1340
rect 135 1337 139 1341
rect 167 1337 171 1341
rect 151 1331 152 1335
rect 152 1331 155 1335
rect 203 1347 207 1351
rect 215 1337 219 1341
rect 303 1337 307 1341
rect 267 1331 271 1335
rect 415 1337 419 1341
rect 639 1355 643 1359
rect 751 1355 755 1359
rect 863 1355 867 1359
rect 967 1355 971 1359
rect 1063 1355 1067 1359
rect 527 1337 531 1341
rect 639 1337 643 1341
rect 751 1337 755 1341
rect 903 1347 907 1351
rect 911 1347 915 1351
rect 863 1337 867 1341
rect 967 1337 971 1341
rect 1063 1337 1067 1341
rect 911 1327 915 1331
rect 1127 1355 1131 1359
rect 1151 1355 1155 1359
rect 1231 1355 1235 1359
rect 1187 1347 1191 1351
rect 1407 1363 1411 1367
rect 1583 1371 1587 1375
rect 1311 1355 1315 1359
rect 1383 1355 1387 1359
rect 1455 1355 1459 1359
rect 1151 1337 1155 1341
rect 1231 1337 1235 1341
rect 1311 1337 1315 1341
rect 1239 1331 1243 1335
rect 1355 1335 1359 1339
rect 1439 1347 1443 1351
rect 1447 1347 1451 1351
rect 1535 1355 1539 1359
rect 1583 1353 1587 1357
rect 1383 1337 1387 1341
rect 1455 1337 1459 1341
rect 1463 1331 1467 1335
rect 1535 1337 1539 1341
rect 1583 1336 1587 1340
rect 111 1316 115 1320
rect 135 1315 139 1319
rect 183 1315 187 1319
rect 203 1319 204 1323
rect 204 1319 207 1323
rect 247 1315 251 1319
rect 311 1315 315 1319
rect 375 1315 379 1319
rect 407 1319 411 1323
rect 439 1315 443 1319
rect 479 1319 483 1323
rect 495 1315 499 1319
rect 543 1315 547 1319
rect 591 1315 595 1319
rect 639 1315 643 1319
rect 687 1315 691 1319
rect 743 1315 747 1319
rect 791 1315 795 1319
rect 839 1315 843 1319
rect 887 1315 891 1319
rect 903 1319 904 1323
rect 904 1319 907 1323
rect 935 1315 939 1319
rect 991 1315 995 1319
rect 1055 1323 1059 1327
rect 1047 1315 1051 1319
rect 1103 1315 1107 1319
rect 1159 1315 1163 1319
rect 1215 1315 1219 1319
rect 1271 1315 1275 1319
rect 1327 1315 1331 1319
rect 1375 1315 1379 1319
rect 111 1299 115 1303
rect 151 1303 152 1307
rect 152 1303 155 1307
rect 267 1303 268 1307
rect 268 1303 271 1307
rect 855 1303 856 1307
rect 856 1303 859 1307
rect 1007 1303 1008 1307
rect 1008 1303 1011 1307
rect 1232 1303 1236 1307
rect 1359 1303 1363 1307
rect 1415 1319 1419 1323
rect 1423 1315 1427 1319
rect 1439 1319 1440 1323
rect 1440 1319 1443 1323
rect 1471 1315 1475 1319
rect 1527 1315 1531 1319
rect 1583 1316 1587 1320
rect 135 1297 139 1301
rect 183 1297 187 1301
rect 247 1297 251 1301
rect 311 1297 315 1301
rect 375 1297 379 1301
rect 439 1297 443 1301
rect 495 1297 499 1301
rect 543 1297 547 1301
rect 591 1297 595 1301
rect 639 1297 643 1301
rect 687 1297 691 1301
rect 743 1297 747 1301
rect 791 1297 795 1301
rect 839 1297 843 1301
rect 887 1297 891 1301
rect 935 1297 939 1301
rect 991 1297 995 1301
rect 1047 1297 1051 1301
rect 1103 1297 1107 1301
rect 1159 1297 1163 1301
rect 1215 1297 1219 1301
rect 1271 1297 1275 1301
rect 1327 1297 1331 1301
rect 1375 1297 1379 1301
rect 1423 1297 1427 1301
rect 1471 1297 1475 1301
rect 1527 1297 1531 1301
rect 111 1281 115 1285
rect 135 1283 139 1287
rect 191 1283 195 1287
rect 255 1283 259 1287
rect 327 1283 331 1287
rect 391 1283 395 1287
rect 463 1283 467 1287
rect 535 1283 539 1287
rect 599 1283 603 1287
rect 663 1283 667 1287
rect 727 1283 731 1287
rect 791 1283 795 1287
rect 1019 1291 1023 1295
rect 855 1283 859 1287
rect 927 1283 931 1287
rect 999 1283 1003 1287
rect 1063 1283 1067 1287
rect 1223 1291 1227 1295
rect 1127 1283 1131 1287
rect 1191 1283 1195 1287
rect 1247 1283 1251 1287
rect 111 1264 115 1268
rect 135 1265 139 1269
rect 191 1265 195 1269
rect 151 1259 152 1263
rect 152 1259 155 1263
rect 247 1275 251 1279
rect 255 1265 259 1269
rect 303 1259 307 1263
rect 327 1265 331 1269
rect 391 1265 395 1269
rect 407 1275 408 1279
rect 408 1275 411 1279
rect 479 1275 480 1279
rect 480 1275 483 1279
rect 463 1265 467 1269
rect 535 1265 539 1269
rect 599 1265 603 1269
rect 663 1265 667 1269
rect 619 1259 620 1263
rect 620 1259 623 1263
rect 875 1275 876 1279
rect 876 1275 879 1279
rect 727 1265 731 1269
rect 791 1265 795 1269
rect 815 1267 819 1271
rect 855 1265 859 1269
rect 847 1259 851 1263
rect 1055 1275 1059 1279
rect 927 1265 931 1269
rect 999 1265 1003 1269
rect 1063 1265 1067 1269
rect 1007 1259 1011 1263
rect 1019 1259 1020 1263
rect 1020 1259 1023 1263
rect 1075 1259 1079 1263
rect 1127 1265 1131 1269
rect 1191 1265 1195 1269
rect 1247 1265 1251 1269
rect 1223 1259 1227 1263
rect 1415 1291 1419 1295
rect 1583 1299 1587 1303
rect 1303 1283 1307 1287
rect 1367 1283 1371 1287
rect 111 1244 115 1248
rect 135 1243 139 1247
rect 175 1243 179 1247
rect 231 1243 235 1247
rect 247 1247 248 1251
rect 248 1247 251 1251
rect 287 1243 291 1247
rect 335 1251 339 1255
rect 351 1243 355 1247
rect 415 1243 419 1247
rect 431 1247 432 1251
rect 432 1247 435 1251
rect 479 1243 483 1247
rect 543 1243 547 1247
rect 571 1251 575 1255
rect 1303 1265 1307 1269
rect 1431 1283 1435 1287
rect 1583 1281 1587 1285
rect 1367 1265 1371 1269
rect 1359 1259 1363 1263
rect 1431 1265 1435 1269
rect 1583 1264 1587 1268
rect 607 1243 611 1247
rect 671 1243 675 1247
rect 735 1243 739 1247
rect 799 1243 803 1247
rect 815 1247 816 1251
rect 816 1247 819 1251
rect 863 1243 867 1247
rect 875 1247 879 1251
rect 927 1243 931 1247
rect 991 1243 995 1247
rect 1055 1243 1059 1247
rect 1119 1243 1123 1247
rect 1175 1247 1179 1251
rect 1183 1243 1187 1247
rect 1247 1243 1251 1247
rect 1311 1243 1315 1247
rect 1375 1243 1379 1247
rect 1439 1243 1443 1247
rect 1487 1247 1491 1251
rect 1503 1243 1507 1247
rect 1543 1243 1547 1247
rect 1583 1244 1587 1248
rect 111 1227 115 1231
rect 155 1231 156 1235
rect 156 1231 159 1235
rect 303 1231 304 1235
rect 304 1231 307 1235
rect 571 1231 575 1235
rect 619 1231 623 1235
rect 703 1231 707 1235
rect 947 1231 948 1235
rect 948 1231 951 1235
rect 1075 1231 1076 1235
rect 1076 1231 1079 1235
rect 1295 1231 1299 1235
rect 135 1225 139 1229
rect 175 1225 179 1229
rect 231 1225 235 1229
rect 287 1225 291 1229
rect 351 1225 355 1229
rect 415 1225 419 1229
rect 479 1225 483 1229
rect 543 1225 547 1229
rect 607 1225 611 1229
rect 671 1225 675 1229
rect 735 1225 739 1229
rect 799 1225 803 1229
rect 863 1225 867 1229
rect 927 1225 931 1229
rect 991 1225 995 1229
rect 1055 1225 1059 1229
rect 1119 1225 1123 1229
rect 1183 1225 1187 1229
rect 1247 1225 1251 1229
rect 1311 1225 1315 1229
rect 1375 1225 1379 1229
rect 295 1219 299 1223
rect 111 1209 115 1213
rect 143 1211 147 1215
rect 175 1211 179 1215
rect 215 1211 219 1215
rect 263 1211 267 1215
rect 311 1211 315 1215
rect 359 1211 363 1215
rect 415 1211 419 1215
rect 471 1211 475 1215
rect 527 1211 531 1215
rect 583 1211 587 1215
rect 639 1211 643 1215
rect 687 1211 691 1215
rect 735 1211 739 1215
rect 783 1211 787 1215
rect 831 1211 835 1215
rect 879 1211 883 1215
rect 935 1211 939 1215
rect 111 1192 115 1196
rect 143 1193 147 1197
rect 175 1193 179 1197
rect 155 1187 159 1191
rect 231 1203 232 1207
rect 232 1203 235 1207
rect 215 1193 219 1197
rect 263 1193 267 1197
rect 311 1193 315 1197
rect 295 1187 299 1191
rect 328 1203 332 1207
rect 431 1203 432 1207
rect 432 1203 435 1207
rect 359 1193 363 1197
rect 415 1193 419 1197
rect 423 1187 427 1191
rect 471 1193 475 1197
rect 527 1193 531 1197
rect 583 1193 587 1197
rect 639 1193 643 1197
rect 687 1193 691 1197
rect 611 1187 615 1191
rect 703 1187 704 1191
rect 704 1187 707 1191
rect 735 1193 739 1197
rect 783 1193 787 1197
rect 831 1193 835 1197
rect 1047 1219 1051 1223
rect 1175 1219 1179 1223
rect 1559 1231 1560 1235
rect 1560 1231 1563 1235
rect 1439 1225 1443 1229
rect 1503 1225 1507 1229
rect 1543 1225 1547 1229
rect 1583 1227 1587 1231
rect 983 1211 987 1215
rect 1039 1211 1043 1215
rect 1095 1211 1099 1215
rect 1159 1211 1163 1215
rect 1231 1211 1235 1215
rect 1303 1211 1307 1215
rect 879 1193 883 1197
rect 935 1193 939 1197
rect 947 1187 951 1191
rect 999 1203 1000 1207
rect 1000 1203 1003 1207
rect 983 1193 987 1197
rect 1039 1193 1043 1197
rect 1095 1193 1099 1197
rect 1047 1187 1051 1191
rect 1159 1193 1163 1197
rect 1231 1193 1235 1197
rect 1383 1211 1387 1215
rect 1471 1211 1475 1215
rect 1543 1211 1547 1215
rect 1583 1209 1587 1213
rect 1303 1193 1307 1197
rect 1295 1187 1299 1191
rect 1487 1203 1488 1207
rect 1488 1203 1491 1207
rect 1383 1193 1387 1197
rect 1471 1193 1475 1197
rect 1543 1193 1547 1197
rect 1583 1192 1587 1196
rect 1559 1187 1560 1191
rect 1560 1187 1563 1191
rect 111 1172 115 1176
rect 143 1171 147 1175
rect 175 1171 179 1175
rect 215 1171 219 1175
rect 231 1175 232 1179
rect 232 1175 235 1179
rect 255 1171 259 1175
rect 303 1171 307 1175
rect 359 1171 363 1175
rect 415 1171 419 1175
rect 471 1171 475 1175
rect 519 1175 523 1179
rect 527 1171 531 1175
rect 591 1171 595 1175
rect 655 1171 659 1175
rect 719 1171 723 1175
rect 791 1171 795 1175
rect 803 1175 807 1179
rect 855 1171 859 1175
rect 919 1171 923 1175
rect 983 1171 987 1175
rect 999 1175 1000 1179
rect 1000 1175 1003 1179
rect 1039 1171 1043 1175
rect 1103 1171 1107 1175
rect 1167 1171 1171 1175
rect 1239 1171 1243 1175
rect 1311 1171 1315 1175
rect 1391 1171 1395 1175
rect 1479 1171 1483 1175
rect 111 1155 115 1159
rect 155 1159 159 1163
rect 431 1159 432 1163
rect 432 1159 435 1163
rect 611 1159 612 1163
rect 612 1159 615 1163
rect 143 1153 147 1157
rect 175 1153 179 1157
rect 215 1153 219 1157
rect 255 1153 259 1157
rect 303 1153 307 1157
rect 359 1153 363 1157
rect 415 1153 419 1157
rect 471 1153 475 1157
rect 527 1153 531 1157
rect 591 1153 595 1157
rect 655 1153 659 1157
rect 111 1137 115 1141
rect 135 1139 139 1143
rect 167 1139 171 1143
rect 199 1139 203 1143
rect 231 1139 235 1143
rect 263 1139 267 1143
rect 295 1139 299 1143
rect 327 1139 331 1143
rect 359 1139 363 1143
rect 391 1139 395 1143
rect 447 1139 451 1143
rect 111 1120 115 1124
rect 135 1121 139 1125
rect 155 1119 159 1123
rect 167 1121 171 1125
rect 199 1121 203 1125
rect 231 1121 235 1125
rect 263 1121 267 1125
rect 295 1121 299 1125
rect 311 1131 312 1135
rect 312 1131 315 1135
rect 327 1121 331 1125
rect 359 1121 363 1125
rect 347 1115 348 1119
rect 348 1115 351 1119
rect 391 1121 395 1125
rect 519 1147 523 1151
rect 867 1159 871 1163
rect 1419 1159 1423 1163
rect 1495 1175 1496 1179
rect 1496 1175 1499 1179
rect 1543 1171 1547 1175
rect 1583 1172 1587 1176
rect 1559 1159 1560 1163
rect 1560 1159 1563 1163
rect 719 1153 723 1157
rect 791 1153 795 1157
rect 855 1153 859 1157
rect 919 1153 923 1157
rect 983 1153 987 1157
rect 1039 1153 1043 1157
rect 1103 1153 1107 1157
rect 1167 1153 1171 1157
rect 1239 1153 1243 1157
rect 1311 1153 1315 1157
rect 1391 1153 1395 1157
rect 1479 1153 1483 1157
rect 1543 1153 1547 1157
rect 1583 1155 1587 1159
rect 875 1147 879 1151
rect 503 1139 507 1143
rect 559 1139 563 1143
rect 615 1139 619 1143
rect 671 1139 675 1143
rect 727 1139 731 1143
rect 783 1139 787 1143
rect 839 1139 843 1143
rect 895 1139 899 1143
rect 951 1139 955 1143
rect 1007 1139 1011 1143
rect 447 1121 451 1125
rect 503 1121 507 1125
rect 559 1121 563 1125
rect 615 1121 619 1125
rect 607 1115 611 1119
rect 671 1121 675 1125
rect 727 1121 731 1125
rect 803 1131 804 1135
rect 804 1131 807 1135
rect 783 1121 787 1125
rect 839 1121 843 1125
rect 867 1115 871 1119
rect 895 1121 899 1125
rect 951 1121 955 1125
rect 1007 1121 1011 1125
rect 1227 1147 1231 1151
rect 1063 1139 1067 1143
rect 1127 1139 1131 1143
rect 1191 1139 1195 1143
rect 1255 1139 1259 1143
rect 1327 1139 1331 1143
rect 1063 1121 1067 1125
rect 1127 1121 1131 1125
rect 1159 1115 1163 1119
rect 1191 1121 1195 1125
rect 1255 1121 1259 1125
rect 1399 1139 1403 1143
rect 1479 1139 1483 1143
rect 1543 1139 1547 1143
rect 1583 1137 1587 1141
rect 1327 1121 1331 1125
rect 1495 1131 1496 1135
rect 1496 1131 1499 1135
rect 1399 1121 1403 1125
rect 1479 1121 1483 1125
rect 1543 1121 1547 1125
rect 1583 1120 1587 1124
rect 1519 1115 1523 1119
rect 1559 1115 1560 1119
rect 1560 1115 1563 1119
rect 111 1100 115 1104
rect 151 1099 155 1103
rect 167 1099 171 1103
rect 183 1099 187 1103
rect 223 1099 227 1103
rect 271 1099 275 1103
rect 327 1099 331 1103
rect 383 1099 387 1103
rect 439 1099 443 1103
rect 495 1103 499 1107
rect 503 1099 507 1103
rect 567 1099 571 1103
rect 639 1099 643 1103
rect 711 1099 715 1103
rect 783 1099 787 1103
rect 855 1099 859 1103
rect 875 1103 876 1107
rect 876 1103 879 1107
rect 919 1099 923 1103
rect 983 1099 987 1103
rect 1039 1099 1043 1103
rect 1095 1099 1099 1103
rect 1151 1099 1155 1103
rect 1207 1099 1211 1103
rect 1227 1103 1228 1107
rect 1228 1103 1231 1107
rect 1263 1099 1267 1103
rect 1319 1099 1323 1103
rect 1375 1099 1379 1103
rect 1411 1107 1415 1111
rect 1439 1099 1443 1103
rect 1503 1099 1507 1103
rect 1543 1099 1547 1103
rect 1583 1100 1587 1104
rect 111 1083 115 1087
rect 151 1081 155 1085
rect 183 1081 187 1085
rect 223 1081 227 1085
rect 271 1081 275 1085
rect 327 1081 331 1085
rect 383 1081 387 1085
rect 347 1075 351 1079
rect 439 1081 443 1085
rect 503 1081 507 1085
rect 567 1081 571 1085
rect 639 1081 643 1085
rect 711 1081 715 1085
rect 783 1081 787 1085
rect 607 1075 611 1079
rect 1167 1087 1168 1091
rect 1168 1087 1171 1091
rect 1391 1087 1392 1091
rect 1392 1087 1395 1091
rect 1519 1087 1520 1091
rect 1520 1087 1523 1091
rect 1559 1087 1560 1091
rect 1560 1087 1563 1091
rect 855 1081 859 1085
rect 919 1081 923 1085
rect 983 1081 987 1085
rect 1039 1081 1043 1085
rect 1095 1081 1099 1085
rect 1151 1081 1155 1085
rect 1207 1081 1211 1085
rect 1263 1081 1267 1085
rect 1319 1081 1323 1085
rect 1375 1081 1379 1085
rect 1439 1081 1443 1085
rect 1503 1081 1507 1085
rect 1543 1081 1547 1085
rect 1583 1083 1587 1087
rect 1159 1075 1163 1079
rect 1419 1075 1423 1079
rect 495 1067 499 1071
rect 111 1057 115 1061
rect 447 1059 451 1063
rect 487 1059 491 1063
rect 543 1059 547 1063
rect 599 1059 603 1063
rect 663 1059 667 1063
rect 727 1059 731 1063
rect 791 1059 795 1063
rect 863 1059 867 1063
rect 935 1059 939 1063
rect 1007 1059 1011 1063
rect 1079 1059 1083 1063
rect 1151 1059 1155 1063
rect 1215 1059 1219 1063
rect 1279 1059 1283 1063
rect 1335 1059 1339 1063
rect 1391 1059 1395 1063
rect 1447 1059 1451 1063
rect 1503 1059 1507 1063
rect 1543 1059 1547 1063
rect 1583 1057 1587 1061
rect 111 1040 115 1044
rect 447 1041 451 1045
rect 487 1041 491 1045
rect 543 1041 547 1045
rect 599 1041 603 1045
rect 663 1041 667 1045
rect 727 1041 731 1045
rect 791 1041 795 1045
rect 863 1041 867 1045
rect 987 1051 991 1055
rect 995 1051 999 1055
rect 935 1041 939 1045
rect 1007 1041 1011 1045
rect 719 1027 723 1031
rect 995 1031 999 1035
rect 1079 1041 1083 1045
rect 1187 1051 1191 1055
rect 1151 1041 1155 1045
rect 1215 1041 1219 1045
rect 1167 1035 1168 1039
rect 1168 1035 1171 1039
rect 1279 1041 1283 1045
rect 1411 1051 1412 1055
rect 1412 1051 1415 1055
rect 1335 1041 1339 1045
rect 1391 1041 1395 1045
rect 1447 1041 1451 1045
rect 1383 1035 1387 1039
rect 1531 1051 1535 1055
rect 1503 1041 1507 1045
rect 1543 1041 1547 1045
rect 1583 1040 1587 1044
rect 1475 1035 1479 1039
rect 1559 1035 1560 1039
rect 1560 1035 1563 1039
rect 111 1016 115 1020
rect 511 1015 515 1019
rect 543 1015 547 1019
rect 575 1015 579 1019
rect 615 1015 619 1019
rect 627 1019 631 1023
rect 663 1015 667 1019
rect 711 1015 715 1019
rect 775 1015 779 1019
rect 847 1015 851 1019
rect 927 1015 931 1019
rect 979 1019 983 1023
rect 987 1023 991 1027
rect 1007 1015 1011 1019
rect 1087 1015 1091 1019
rect 1167 1015 1171 1019
rect 1187 1019 1188 1023
rect 1188 1019 1191 1023
rect 1239 1015 1243 1019
rect 1303 1015 1307 1019
rect 1359 1015 1363 1019
rect 1407 1015 1411 1019
rect 1455 1015 1459 1019
rect 1511 1015 1515 1019
rect 1531 1019 1532 1023
rect 1532 1019 1535 1023
rect 1543 1015 1547 1019
rect 1583 1016 1587 1020
rect 111 999 115 1003
rect 727 1003 728 1007
rect 728 1003 731 1007
rect 791 1003 792 1007
rect 792 1003 795 1007
rect 511 997 515 1001
rect 543 997 547 1001
rect 575 997 579 1001
rect 615 997 619 1001
rect 663 997 667 1001
rect 711 997 715 1001
rect 775 997 779 1001
rect 847 997 851 1001
rect 927 997 931 1001
rect 1007 997 1011 1001
rect 1087 997 1091 1001
rect 979 991 983 995
rect 1475 1003 1476 1007
rect 1476 1003 1479 1007
rect 1559 1003 1560 1007
rect 1560 1003 1563 1007
rect 1167 997 1171 1001
rect 1239 997 1243 1001
rect 1303 997 1307 1001
rect 1359 997 1363 1001
rect 1407 997 1411 1001
rect 1455 997 1459 1001
rect 1511 997 1515 1001
rect 1543 997 1547 1001
rect 1583 999 1587 1003
rect 111 973 115 977
rect 159 975 163 979
rect 199 975 203 979
rect 255 975 259 979
rect 311 975 315 979
rect 375 975 379 979
rect 439 975 443 979
rect 503 975 507 979
rect 559 975 563 979
rect 627 983 631 987
rect 823 983 827 987
rect 615 975 619 979
rect 663 975 667 979
rect 703 975 707 979
rect 735 975 739 979
rect 775 975 779 979
rect 831 975 835 979
rect 895 975 899 979
rect 967 975 971 979
rect 1047 975 1051 979
rect 1127 975 1131 979
rect 1199 975 1203 979
rect 1271 975 1275 979
rect 1343 975 1347 979
rect 1415 975 1419 979
rect 1487 975 1491 979
rect 1543 975 1547 979
rect 1583 973 1587 977
rect 171 967 175 971
rect 111 956 115 960
rect 159 957 163 961
rect 199 957 203 961
rect 255 957 259 961
rect 311 957 315 961
rect 375 957 379 961
rect 439 957 443 961
rect 503 957 507 961
rect 559 957 563 961
rect 587 967 591 971
rect 615 957 619 961
rect 451 951 455 955
rect 523 951 524 955
rect 524 951 527 955
rect 663 957 667 961
rect 703 957 707 961
rect 735 957 739 961
rect 775 957 779 961
rect 783 951 787 955
rect 791 951 792 955
rect 792 951 795 955
rect 831 957 835 961
rect 895 957 899 961
rect 967 957 971 961
rect 1047 957 1051 961
rect 1127 957 1131 961
rect 1219 967 1220 971
rect 1220 967 1223 971
rect 1199 957 1203 961
rect 1271 957 1275 961
rect 1343 957 1347 961
rect 1415 957 1419 961
rect 1487 957 1491 961
rect 1543 957 1547 961
rect 1583 956 1587 960
rect 1499 951 1503 955
rect 1559 951 1560 955
rect 1560 951 1563 955
rect 111 936 115 940
rect 151 935 155 939
rect 171 939 172 943
rect 172 939 175 943
rect 191 935 195 939
rect 247 935 251 939
rect 303 935 307 939
rect 319 939 320 943
rect 320 939 323 943
rect 367 935 371 939
rect 431 935 435 939
rect 495 935 499 939
rect 551 939 555 943
rect 559 935 563 939
rect 615 935 619 939
rect 671 935 675 939
rect 719 935 723 939
rect 767 935 771 939
rect 823 943 827 947
rect 815 935 819 939
rect 871 935 875 939
rect 935 935 939 939
rect 1007 935 1011 939
rect 1079 935 1083 939
rect 1143 935 1147 939
rect 1207 935 1211 939
rect 1219 939 1223 943
rect 1271 935 1275 939
rect 1327 935 1331 939
rect 1375 935 1379 939
rect 1423 935 1427 939
rect 1471 935 1475 939
rect 1511 935 1515 939
rect 1543 935 1547 939
rect 1583 936 1587 940
rect 111 919 115 923
rect 263 923 264 927
rect 264 923 267 927
rect 451 923 452 927
rect 452 923 455 927
rect 783 923 784 927
rect 784 923 787 927
rect 151 917 155 921
rect 191 917 195 921
rect 247 917 251 921
rect 303 917 307 921
rect 367 917 371 921
rect 431 917 435 921
rect 495 917 499 921
rect 559 917 563 921
rect 615 917 619 921
rect 671 917 675 921
rect 719 917 723 921
rect 767 917 771 921
rect 815 917 819 921
rect 871 917 875 921
rect 935 917 939 921
rect 1007 917 1011 921
rect 1079 917 1083 921
rect 1143 917 1147 921
rect 551 907 555 911
rect 1367 923 1371 927
rect 1499 923 1503 927
rect 1207 917 1211 921
rect 1271 917 1275 921
rect 1327 917 1331 921
rect 1375 917 1379 921
rect 1423 917 1427 921
rect 1471 917 1475 921
rect 1511 917 1515 921
rect 1543 917 1547 921
rect 1583 919 1587 923
rect 111 897 115 901
rect 135 899 139 903
rect 167 899 171 903
rect 223 899 227 903
rect 279 899 283 903
rect 335 899 339 903
rect 391 899 395 903
rect 447 899 451 903
rect 503 899 507 903
rect 559 899 563 903
rect 623 899 627 903
rect 695 899 699 903
rect 151 891 152 895
rect 152 891 155 895
rect 111 880 115 884
rect 135 881 139 885
rect 167 881 171 885
rect 319 891 323 895
rect 223 881 227 885
rect 279 881 283 885
rect 263 875 267 879
rect 335 881 339 885
rect 391 881 395 885
rect 447 881 451 885
rect 111 860 115 864
rect 135 859 139 863
rect 151 863 152 867
rect 152 863 155 867
rect 167 859 171 863
rect 207 859 211 863
rect 255 859 259 863
rect 267 863 271 867
rect 303 859 307 863
rect 343 859 347 863
rect 483 875 487 879
rect 503 881 507 885
rect 559 881 563 885
rect 623 881 627 885
rect 759 899 763 903
rect 823 899 827 903
rect 887 899 891 903
rect 951 899 955 903
rect 1015 899 1019 903
rect 1079 899 1083 903
rect 1135 899 1139 903
rect 1527 907 1531 911
rect 1191 899 1195 903
rect 1247 899 1251 903
rect 1303 899 1307 903
rect 1359 899 1363 903
rect 1407 899 1411 903
rect 1455 899 1459 903
rect 1511 899 1515 903
rect 1543 899 1547 903
rect 1583 897 1587 901
rect 695 881 699 885
rect 759 881 763 885
rect 823 881 827 885
rect 887 881 891 885
rect 951 881 955 885
rect 1015 881 1019 885
rect 1079 881 1083 885
rect 1135 881 1139 885
rect 1191 881 1195 885
rect 1247 881 1251 885
rect 1279 891 1283 895
rect 1287 891 1291 895
rect 1303 881 1307 885
rect 1287 871 1291 875
rect 1359 881 1363 885
rect 1407 881 1411 885
rect 1367 875 1371 879
rect 1455 881 1459 885
rect 1511 881 1515 885
rect 1543 881 1547 885
rect 1495 875 1499 879
rect 1527 875 1528 879
rect 1528 875 1531 879
rect 1559 891 1560 895
rect 1560 891 1563 895
rect 1583 880 1587 884
rect 383 859 387 863
rect 439 859 443 863
rect 511 859 515 863
rect 591 859 595 863
rect 679 859 683 863
rect 767 859 771 863
rect 847 859 851 863
rect 919 859 923 863
rect 983 859 987 863
rect 1039 859 1043 863
rect 1095 859 1099 863
rect 1151 859 1155 863
rect 111 843 115 847
rect 223 847 224 851
rect 224 847 227 851
rect 135 841 139 845
rect 167 841 171 845
rect 207 841 211 845
rect 255 841 259 845
rect 303 841 307 845
rect 343 841 347 845
rect 383 841 387 845
rect 439 841 443 845
rect 483 839 487 843
rect 511 841 515 845
rect 591 841 595 845
rect 679 841 683 845
rect 767 841 771 845
rect 847 841 851 845
rect 919 841 923 845
rect 983 841 987 845
rect 1039 841 1043 845
rect 1095 841 1099 845
rect 1019 835 1023 839
rect 1207 859 1211 863
rect 1263 859 1267 863
rect 1279 863 1280 867
rect 1280 863 1283 867
rect 1327 859 1331 863
rect 1399 859 1403 863
rect 1479 859 1483 863
rect 1543 859 1547 863
rect 1559 863 1560 867
rect 1560 863 1563 867
rect 1583 860 1587 864
rect 1151 841 1155 845
rect 1207 841 1211 845
rect 1263 841 1267 845
rect 1327 841 1331 845
rect 1399 841 1403 845
rect 1495 847 1496 851
rect 1496 847 1499 851
rect 1479 841 1483 845
rect 1543 841 1547 845
rect 1583 843 1587 847
rect 111 821 115 825
rect 135 823 139 827
rect 167 823 171 827
rect 223 823 227 827
rect 287 823 291 827
rect 351 823 355 827
rect 423 823 427 827
rect 495 823 499 827
rect 151 815 152 819
rect 152 815 155 819
rect 111 804 115 808
rect 135 805 139 809
rect 167 805 171 809
rect 267 815 271 819
rect 223 805 227 809
rect 215 799 219 803
rect 287 805 291 809
rect 351 805 355 809
rect 423 805 427 809
rect 371 799 372 803
rect 372 799 375 803
rect 567 823 571 827
rect 639 823 643 827
rect 719 823 723 827
rect 791 823 795 827
rect 863 823 867 827
rect 935 823 939 827
rect 999 823 1003 827
rect 1055 823 1059 827
rect 1103 823 1107 827
rect 1143 823 1147 827
rect 1183 823 1187 827
rect 1231 823 1235 827
rect 1247 827 1251 831
rect 1279 823 1283 827
rect 1327 823 1331 827
rect 495 805 499 809
rect 567 805 571 809
rect 503 799 507 803
rect 751 815 755 819
rect 639 805 643 809
rect 719 805 723 809
rect 687 799 691 803
rect 791 805 795 809
rect 863 805 867 809
rect 935 805 939 809
rect 999 805 1003 809
rect 1007 799 1011 803
rect 1019 799 1020 803
rect 1020 799 1023 803
rect 1087 815 1091 819
rect 1055 805 1059 809
rect 1103 805 1107 809
rect 1143 805 1147 809
rect 111 784 115 788
rect 135 783 139 787
rect 151 787 152 791
rect 152 787 155 791
rect 167 783 171 787
rect 199 783 203 787
rect 247 783 251 787
rect 303 783 307 787
rect 359 783 363 787
rect 423 783 427 787
rect 487 783 491 787
rect 551 783 555 787
rect 599 787 603 791
rect 607 783 611 787
rect 671 783 675 787
rect 735 783 739 787
rect 751 787 752 791
rect 752 787 755 791
rect 1087 795 1091 799
rect 1183 805 1187 809
rect 1231 805 1235 809
rect 1279 805 1283 809
rect 1583 821 1587 825
rect 1327 805 1331 809
rect 1583 804 1587 808
rect 799 783 803 787
rect 871 783 875 787
rect 883 787 887 791
rect 935 783 939 787
rect 999 783 1003 787
rect 1063 783 1067 787
rect 1127 783 1131 787
rect 1191 783 1195 787
rect 1247 787 1251 791
rect 1255 783 1259 787
rect 1319 783 1323 787
rect 1383 783 1387 787
rect 1583 784 1587 788
rect 111 767 115 771
rect 215 771 216 775
rect 216 771 219 775
rect 371 771 375 775
rect 535 771 539 775
rect 687 771 688 775
rect 688 771 691 775
rect 811 771 815 775
rect 135 765 139 769
rect 167 765 171 769
rect 199 765 203 769
rect 247 765 251 769
rect 303 765 307 769
rect 359 765 363 769
rect 423 765 427 769
rect 487 765 491 769
rect 551 765 555 769
rect 607 765 611 769
rect 671 765 675 769
rect 735 765 739 769
rect 799 765 803 769
rect 871 765 875 769
rect 935 765 939 769
rect 999 765 1003 769
rect 1011 767 1015 771
rect 1079 771 1080 775
rect 1080 771 1083 775
rect 1063 765 1067 769
rect 1127 765 1131 769
rect 1191 765 1195 769
rect 1255 765 1259 769
rect 1319 765 1323 769
rect 1383 765 1387 769
rect 1291 759 1295 763
rect 1583 767 1587 771
rect 111 749 115 753
rect 135 751 139 755
rect 167 751 171 755
rect 199 751 203 755
rect 255 751 259 755
rect 319 751 323 755
rect 391 751 395 755
rect 463 751 467 755
rect 543 751 547 755
rect 623 751 627 755
rect 703 751 707 755
rect 775 751 779 755
rect 847 751 851 755
rect 919 751 923 755
rect 991 751 995 755
rect 1063 751 1067 755
rect 1135 751 1139 755
rect 1207 751 1211 755
rect 1271 751 1275 755
rect 1327 751 1331 755
rect 1375 751 1379 755
rect 1423 751 1427 755
rect 1471 751 1475 755
rect 1511 751 1515 755
rect 1543 751 1547 755
rect 1583 749 1587 753
rect 151 743 152 747
rect 152 743 155 747
rect 111 732 115 736
rect 135 733 139 737
rect 167 733 171 737
rect 199 733 203 737
rect 215 735 219 739
rect 255 733 259 737
rect 319 733 323 737
rect 503 743 507 747
rect 559 743 560 747
rect 560 743 563 747
rect 599 743 603 747
rect 767 743 771 747
rect 391 733 395 737
rect 463 733 467 737
rect 543 733 547 737
rect 623 733 627 737
rect 703 733 707 737
rect 775 733 779 737
rect 399 727 403 731
rect 443 727 447 731
rect 535 727 539 731
rect 635 727 639 731
rect 883 743 887 747
rect 847 733 851 737
rect 811 727 815 731
rect 919 733 923 737
rect 991 733 995 737
rect 1063 733 1067 737
rect 1023 727 1027 731
rect 1079 727 1080 731
rect 1080 727 1083 731
rect 1187 743 1191 747
rect 1135 733 1139 737
rect 1207 733 1211 737
rect 1271 733 1275 737
rect 1291 727 1292 731
rect 1292 727 1295 731
rect 1327 733 1331 737
rect 1375 733 1379 737
rect 1423 733 1427 737
rect 1471 733 1475 737
rect 1511 733 1515 737
rect 1543 733 1547 737
rect 1559 743 1560 747
rect 1560 743 1563 747
rect 1583 732 1587 736
rect 111 712 115 716
rect 135 711 139 715
rect 151 715 152 719
rect 152 715 155 719
rect 167 711 171 715
rect 207 711 211 715
rect 255 711 259 715
rect 271 715 272 719
rect 272 715 275 719
rect 311 711 315 715
rect 367 711 371 715
rect 423 711 427 715
rect 435 715 439 719
rect 479 711 483 715
rect 543 711 547 715
rect 111 695 115 699
rect 223 699 224 703
rect 224 699 227 703
rect 399 699 403 703
rect 443 699 444 703
rect 444 699 447 703
rect 535 699 539 703
rect 559 715 560 719
rect 560 715 563 719
rect 615 711 619 715
rect 659 719 663 723
rect 687 711 691 715
rect 767 719 771 723
rect 759 711 763 715
rect 839 711 843 715
rect 855 715 856 719
rect 856 715 859 719
rect 919 711 923 715
rect 635 699 636 703
rect 636 699 639 703
rect 715 703 719 707
rect 1007 711 1011 715
rect 1087 711 1091 715
rect 1023 699 1024 703
rect 1024 699 1027 703
rect 1035 703 1039 707
rect 1167 711 1171 715
rect 1187 715 1188 719
rect 1188 715 1191 719
rect 1239 711 1243 715
rect 1295 715 1299 719
rect 1303 711 1307 715
rect 1359 711 1363 715
rect 1407 711 1411 715
rect 1455 711 1459 715
rect 1511 711 1515 715
rect 1543 711 1547 715
rect 1559 715 1560 719
rect 1560 715 1563 719
rect 1583 712 1587 716
rect 1351 699 1355 703
rect 135 693 139 697
rect 167 693 171 697
rect 207 693 211 697
rect 255 693 259 697
rect 311 693 315 697
rect 367 693 371 697
rect 423 693 427 697
rect 479 693 483 697
rect 543 693 547 697
rect 615 693 619 697
rect 687 693 691 697
rect 759 693 763 697
rect 839 693 843 697
rect 919 693 923 697
rect 1007 693 1011 697
rect 1087 693 1091 697
rect 1167 693 1171 697
rect 1239 693 1243 697
rect 1303 693 1307 697
rect 1359 693 1363 697
rect 1295 687 1299 691
rect 1407 693 1411 697
rect 1455 693 1459 697
rect 1511 693 1515 697
rect 1543 693 1547 697
rect 1583 695 1587 699
rect 111 677 115 681
rect 159 679 163 683
rect 207 679 211 683
rect 255 679 259 683
rect 303 679 307 683
rect 359 679 363 683
rect 415 679 419 683
rect 471 679 475 683
rect 527 679 531 683
rect 583 679 587 683
rect 639 679 643 683
rect 695 679 699 683
rect 759 679 763 683
rect 823 679 827 683
rect 887 679 891 683
rect 951 679 955 683
rect 1015 679 1019 683
rect 1079 679 1083 683
rect 1135 679 1139 683
rect 1191 679 1195 683
rect 1247 679 1251 683
rect 1303 679 1307 683
rect 1359 679 1363 683
rect 1583 677 1587 681
rect 179 671 180 675
rect 180 671 183 675
rect 111 660 115 664
rect 159 661 163 665
rect 271 671 272 675
rect 272 671 275 675
rect 207 661 211 665
rect 255 661 259 665
rect 223 655 224 659
rect 224 655 227 659
rect 303 661 307 665
rect 435 671 436 675
rect 436 671 439 675
rect 443 671 447 675
rect 507 671 511 675
rect 359 661 363 665
rect 415 661 419 665
rect 471 661 475 665
rect 527 661 531 665
rect 583 661 587 665
rect 403 655 407 659
rect 451 655 455 659
rect 535 655 539 659
rect 603 655 604 659
rect 604 655 607 659
rect 659 671 660 675
rect 660 671 663 675
rect 639 661 643 665
rect 695 661 699 665
rect 715 655 716 659
rect 716 655 719 659
rect 775 671 776 675
rect 776 671 779 675
rect 855 671 859 675
rect 759 661 763 665
rect 823 661 827 665
rect 887 661 891 665
rect 951 661 955 665
rect 1015 661 1019 665
rect 1035 655 1036 659
rect 1036 655 1039 659
rect 1127 671 1131 675
rect 1183 671 1187 675
rect 1079 661 1083 665
rect 1135 661 1139 665
rect 1191 661 1195 665
rect 1247 661 1251 665
rect 1303 661 1307 665
rect 1359 661 1363 665
rect 1583 660 1587 664
rect 1351 655 1355 659
rect 443 647 447 651
rect 907 647 911 651
rect 111 636 115 640
rect 167 635 171 639
rect 179 639 183 643
rect 215 635 219 639
rect 271 635 275 639
rect 327 635 331 639
rect 339 639 343 643
rect 383 635 387 639
rect 431 635 435 639
rect 443 639 447 643
rect 487 635 491 639
rect 507 639 508 643
rect 508 639 511 643
rect 535 635 539 639
rect 591 635 595 639
rect 647 635 651 639
rect 703 635 707 639
rect 759 635 763 639
rect 775 639 776 643
rect 776 639 779 643
rect 823 635 827 639
rect 835 639 839 643
rect 887 635 891 639
rect 943 635 947 639
rect 999 635 1003 639
rect 111 619 115 623
rect 303 623 307 627
rect 403 623 404 627
rect 404 623 407 627
rect 451 623 452 627
rect 452 623 455 627
rect 575 623 579 627
rect 603 623 607 627
rect 907 623 908 627
rect 908 623 911 627
rect 991 623 995 627
rect 1055 635 1059 639
rect 1111 635 1115 639
rect 1127 639 1128 643
rect 1128 639 1131 643
rect 1167 635 1171 639
rect 1183 639 1184 643
rect 1184 639 1187 643
rect 1215 635 1219 639
rect 1271 635 1275 639
rect 1327 635 1331 639
rect 1383 635 1387 639
rect 1439 635 1443 639
rect 1503 635 1507 639
rect 1523 639 1524 643
rect 1524 639 1527 643
rect 1543 635 1547 639
rect 1583 636 1587 640
rect 167 617 171 621
rect 215 617 219 621
rect 271 617 275 621
rect 327 617 331 621
rect 383 617 387 621
rect 431 617 435 621
rect 487 617 491 621
rect 535 617 539 621
rect 591 617 595 621
rect 647 617 651 621
rect 703 617 707 621
rect 759 617 763 621
rect 823 617 827 621
rect 887 617 891 621
rect 943 617 947 621
rect 999 617 1003 621
rect 1055 617 1059 621
rect 1111 617 1115 621
rect 1167 617 1171 621
rect 1215 617 1219 621
rect 1271 617 1275 621
rect 1327 617 1331 621
rect 1383 617 1387 621
rect 1439 617 1443 621
rect 1231 611 1235 615
rect 1559 623 1560 627
rect 1560 623 1563 627
rect 1503 617 1507 621
rect 1543 617 1547 621
rect 1583 619 1587 623
rect 111 601 115 605
rect 223 603 227 607
rect 255 603 259 607
rect 287 603 291 607
rect 319 603 323 607
rect 339 601 343 603
rect 211 595 215 599
rect 111 584 115 588
rect 223 585 227 589
rect 255 585 259 589
rect 287 585 291 589
rect 339 599 340 601
rect 340 599 343 601
rect 351 603 355 607
rect 383 603 387 607
rect 423 603 427 607
rect 463 603 467 607
rect 519 603 523 607
rect 583 603 587 607
rect 319 585 323 589
rect 351 585 355 589
rect 303 579 304 583
rect 304 579 307 583
rect 383 585 387 589
rect 443 595 444 599
rect 444 595 447 599
rect 423 585 427 589
rect 415 579 419 583
rect 463 585 467 589
rect 519 585 523 589
rect 647 603 651 607
rect 719 603 723 607
rect 799 603 803 607
rect 887 603 891 607
rect 975 603 979 607
rect 1063 603 1067 607
rect 1143 603 1147 607
rect 1215 603 1219 607
rect 1287 603 1291 607
rect 1351 603 1355 607
rect 1407 603 1411 607
rect 1455 603 1459 607
rect 1511 603 1515 607
rect 1543 603 1547 607
rect 1583 601 1587 605
rect 583 585 587 589
rect 575 579 579 583
rect 647 585 651 589
rect 719 585 723 589
rect 799 585 803 589
rect 835 595 839 599
rect 847 595 851 599
rect 887 585 891 589
rect 975 585 979 589
rect 111 564 115 568
rect 191 563 195 567
rect 211 567 212 571
rect 212 567 215 571
rect 255 563 259 567
rect 327 563 331 567
rect 399 563 403 567
rect 847 575 851 579
rect 991 579 992 583
rect 992 579 995 583
rect 1063 585 1067 589
rect 1183 595 1187 599
rect 1143 585 1147 589
rect 1215 585 1219 589
rect 1231 585 1235 587
rect 1231 583 1232 585
rect 1232 583 1235 585
rect 1287 585 1291 589
rect 1351 585 1355 589
rect 1407 585 1411 589
rect 1487 595 1491 599
rect 1523 595 1527 599
rect 1455 585 1459 589
rect 1511 585 1515 589
rect 1543 585 1547 589
rect 1583 584 1587 588
rect 1527 579 1528 583
rect 1528 579 1531 583
rect 1559 579 1560 583
rect 1560 579 1563 583
rect 471 563 475 567
rect 535 563 539 567
rect 591 567 595 571
rect 599 563 603 567
rect 663 563 667 567
rect 727 563 731 567
rect 783 563 787 567
rect 839 563 843 567
rect 903 563 907 567
rect 967 563 971 567
rect 1039 563 1043 567
rect 1103 563 1107 567
rect 1167 563 1171 567
rect 1183 567 1184 571
rect 1184 567 1187 571
rect 1231 563 1235 567
rect 111 547 115 551
rect 339 551 343 555
rect 415 551 416 555
rect 416 551 419 555
rect 1287 563 1291 567
rect 1335 563 1339 567
rect 1383 563 1387 567
rect 1423 563 1427 567
rect 1471 563 1475 567
rect 1487 567 1488 571
rect 1488 567 1491 571
rect 1551 571 1555 575
rect 1511 563 1515 567
rect 1543 563 1547 567
rect 1583 564 1587 568
rect 1527 551 1528 555
rect 1528 551 1531 555
rect 1559 551 1560 555
rect 1560 551 1563 555
rect 191 545 195 549
rect 255 545 259 549
rect 327 545 331 549
rect 399 545 403 549
rect 471 545 475 549
rect 535 545 539 549
rect 599 545 603 549
rect 663 545 667 549
rect 727 545 731 549
rect 783 545 787 549
rect 839 545 843 549
rect 903 545 907 549
rect 967 545 971 549
rect 1039 545 1043 549
rect 1103 545 1107 549
rect 1167 545 1171 549
rect 1231 545 1235 549
rect 1287 545 1291 549
rect 1335 545 1339 549
rect 1383 545 1387 549
rect 1423 545 1427 549
rect 1471 545 1475 549
rect 1511 545 1515 549
rect 1543 545 1547 549
rect 1583 547 1587 551
rect 591 539 595 543
rect 111 529 115 533
rect 135 531 139 535
rect 175 531 179 535
rect 231 531 235 535
rect 295 531 299 535
rect 359 531 363 535
rect 423 531 427 535
rect 479 531 483 535
rect 543 531 547 535
rect 599 531 603 535
rect 655 531 659 535
rect 711 531 715 535
rect 151 523 152 527
rect 152 523 155 527
rect 111 512 115 516
rect 135 513 139 517
rect 175 513 179 517
rect 231 513 235 517
rect 295 513 299 517
rect 339 511 343 515
rect 359 513 363 517
rect 423 513 427 517
rect 367 507 371 511
rect 479 513 483 517
rect 543 513 547 517
rect 599 513 603 517
rect 655 513 659 517
rect 711 513 715 517
rect 911 539 915 543
rect 767 531 771 535
rect 831 531 835 535
rect 895 531 899 535
rect 967 531 971 535
rect 1031 531 1035 535
rect 695 503 699 507
rect 767 513 771 517
rect 831 513 835 517
rect 895 513 899 517
rect 967 513 971 517
rect 911 507 912 511
rect 912 507 915 511
rect 1095 531 1099 535
rect 1167 531 1171 535
rect 1239 531 1243 535
rect 1311 531 1315 535
rect 1391 531 1395 535
rect 1479 531 1483 535
rect 1543 531 1547 535
rect 1583 529 1587 533
rect 1031 513 1035 517
rect 1095 513 1099 517
rect 1167 513 1171 517
rect 1239 513 1243 517
rect 1311 513 1315 517
rect 1391 513 1395 517
rect 1479 513 1483 517
rect 1543 513 1547 517
rect 1583 512 1587 516
rect 1559 507 1560 511
rect 1560 507 1563 511
rect 111 492 115 496
rect 135 491 139 495
rect 151 495 152 499
rect 152 495 155 499
rect 167 491 171 495
rect 199 491 203 495
rect 247 491 251 495
rect 295 491 299 495
rect 327 495 331 499
rect 343 491 347 495
rect 399 491 403 495
rect 439 495 443 499
rect 455 491 459 495
rect 511 491 515 495
rect 567 491 571 495
rect 623 491 627 495
rect 679 491 683 495
rect 743 491 747 495
rect 815 491 819 495
rect 887 491 891 495
rect 959 491 963 495
rect 1039 491 1043 495
rect 1127 491 1131 495
rect 1215 495 1219 499
rect 1223 491 1227 495
rect 1327 491 1331 495
rect 1439 491 1443 495
rect 1499 499 1503 503
rect 1543 491 1547 495
rect 1583 492 1587 496
rect 111 475 115 479
rect 267 479 268 483
rect 268 479 271 483
rect 360 479 364 483
rect 695 479 696 483
rect 696 479 699 483
rect 1279 479 1283 483
rect 135 473 139 477
rect 167 473 171 477
rect 199 473 203 477
rect 247 473 251 477
rect 295 473 299 477
rect 343 473 347 477
rect 399 473 403 477
rect 455 473 459 477
rect 511 473 515 477
rect 567 473 571 477
rect 623 473 627 477
rect 679 473 683 477
rect 743 473 747 477
rect 815 473 819 477
rect 887 473 891 477
rect 959 473 963 477
rect 1039 473 1043 477
rect 555 467 559 471
rect 111 457 115 461
rect 135 459 139 463
rect 167 459 171 463
rect 199 459 203 463
rect 255 459 259 463
rect 311 459 315 463
rect 367 459 371 463
rect 423 459 427 463
rect 479 459 483 463
rect 535 459 539 463
rect 599 459 603 463
rect 663 459 667 463
rect 735 459 739 463
rect 895 467 899 471
rect 1127 473 1131 477
rect 1223 473 1227 477
rect 1327 473 1331 477
rect 1215 467 1219 471
rect 1555 479 1559 483
rect 1439 473 1443 477
rect 1543 473 1547 477
rect 1583 475 1587 479
rect 807 459 811 463
rect 871 459 875 463
rect 935 459 939 463
rect 991 459 995 463
rect 1047 459 1051 463
rect 1095 459 1099 463
rect 1143 459 1147 463
rect 1199 459 1203 463
rect 1263 459 1267 463
rect 1327 459 1331 463
rect 1399 459 1403 463
rect 1479 459 1483 463
rect 1543 459 1547 463
rect 1583 457 1587 461
rect 151 451 152 455
rect 152 451 155 455
rect 111 440 115 444
rect 135 441 139 445
rect 167 441 171 445
rect 199 441 203 445
rect 327 451 328 455
rect 328 451 331 455
rect 255 441 259 445
rect 311 441 315 445
rect 267 435 271 439
rect 439 451 440 455
rect 440 451 443 455
rect 367 441 371 445
rect 423 441 427 445
rect 379 435 383 439
rect 479 441 483 445
rect 535 441 539 445
rect 599 441 603 445
rect 555 435 556 439
rect 556 435 559 439
rect 563 435 567 439
rect 663 441 667 445
rect 735 441 739 445
rect 779 451 783 455
rect 807 441 811 445
rect 871 441 875 445
rect 935 441 939 445
rect 888 435 892 439
rect 1039 451 1043 455
rect 991 441 995 445
rect 1047 441 1051 445
rect 111 416 115 420
rect 135 415 139 419
rect 151 419 152 423
rect 152 419 155 423
rect 167 415 171 419
rect 231 415 235 419
rect 295 415 299 419
rect 359 415 363 419
rect 423 415 427 419
rect 487 415 491 419
rect 607 427 611 431
rect 1095 441 1099 445
rect 1143 441 1147 445
rect 1199 441 1203 445
rect 1263 441 1267 445
rect 1279 435 1280 439
rect 1280 435 1283 439
rect 1327 441 1331 445
rect 1391 451 1395 455
rect 1499 451 1500 455
rect 1500 451 1503 455
rect 1559 451 1560 455
rect 1560 451 1563 455
rect 1399 441 1403 445
rect 1479 441 1483 445
rect 1543 441 1547 445
rect 1583 440 1587 444
rect 1487 435 1491 439
rect 543 415 547 419
rect 591 415 595 419
rect 639 415 643 419
rect 679 415 683 419
rect 719 415 723 419
rect 759 415 763 419
rect 779 419 780 423
rect 780 419 783 423
rect 807 415 811 419
rect 863 415 867 419
rect 919 415 923 419
rect 975 415 979 419
rect 1039 423 1043 427
rect 1391 427 1395 431
rect 1031 415 1035 419
rect 1087 415 1091 419
rect 1151 415 1155 419
rect 1223 415 1227 419
rect 1303 415 1307 419
rect 1383 415 1387 419
rect 1471 415 1475 419
rect 1503 419 1507 423
rect 1543 415 1547 419
rect 1559 419 1560 423
rect 1560 419 1563 423
rect 1583 416 1587 420
rect 111 399 115 403
rect 311 403 312 407
rect 312 403 315 407
rect 379 403 380 407
rect 380 403 383 407
rect 563 403 564 407
rect 564 403 567 407
rect 607 403 608 407
rect 608 403 611 407
rect 135 397 139 401
rect 167 397 171 401
rect 231 397 235 401
rect 295 397 299 401
rect 359 397 363 401
rect 423 397 427 401
rect 487 397 491 401
rect 543 397 547 401
rect 591 397 595 401
rect 639 397 643 401
rect 679 397 683 401
rect 719 397 723 401
rect 759 397 763 401
rect 807 397 811 401
rect 863 397 867 401
rect 919 397 923 401
rect 975 397 979 401
rect 827 391 831 395
rect 1031 397 1035 401
rect 1087 397 1091 401
rect 1151 397 1155 401
rect 1223 397 1227 401
rect 1303 397 1307 401
rect 1383 397 1387 401
rect 1159 391 1163 395
rect 1487 403 1488 407
rect 1488 403 1491 407
rect 1559 403 1560 407
rect 1560 403 1563 407
rect 1471 397 1475 401
rect 1543 397 1547 401
rect 1583 399 1587 403
rect 111 381 115 385
rect 135 383 139 387
rect 207 383 211 387
rect 295 383 299 387
rect 383 383 387 387
rect 463 383 467 387
rect 535 383 539 387
rect 599 383 603 387
rect 655 383 659 387
rect 703 383 707 387
rect 751 383 755 387
rect 807 383 811 387
rect 863 383 867 387
rect 919 383 923 387
rect 983 383 987 387
rect 1055 383 1059 387
rect 1127 383 1131 387
rect 1199 383 1203 387
rect 1271 383 1275 387
rect 1343 383 1347 387
rect 1415 383 1419 387
rect 1487 383 1491 387
rect 1543 383 1547 387
rect 1583 381 1587 385
rect 151 375 152 379
rect 152 375 155 379
rect 111 364 115 368
rect 135 365 139 369
rect 207 365 211 369
rect 295 365 299 369
rect 311 367 315 371
rect 383 365 387 369
rect 351 359 355 363
rect 463 365 467 369
rect 535 365 539 369
rect 575 359 579 363
rect 599 365 603 369
rect 655 365 659 369
rect 703 365 707 369
rect 751 365 755 369
rect 807 365 811 369
rect 863 365 867 369
rect 827 359 828 363
rect 828 359 831 363
rect 919 365 923 369
rect 983 365 987 369
rect 1055 365 1059 369
rect 1071 375 1072 379
rect 1072 375 1075 379
rect 1127 365 1131 369
rect 1159 359 1163 363
rect 1199 365 1203 369
rect 1271 365 1275 369
rect 1355 375 1359 379
rect 1343 365 1347 369
rect 1415 365 1419 369
rect 1427 359 1431 363
rect 1503 375 1504 379
rect 1504 375 1507 379
rect 1487 365 1491 369
rect 1543 365 1547 369
rect 1583 364 1587 368
rect 1559 359 1560 363
rect 1560 359 1563 363
rect 111 344 115 348
rect 135 343 139 347
rect 151 347 152 351
rect 152 347 155 351
rect 175 343 179 347
rect 223 343 227 347
rect 279 343 283 347
rect 335 343 339 347
rect 391 343 395 347
rect 403 347 407 351
rect 447 343 451 347
rect 495 347 499 351
rect 503 343 507 347
rect 567 343 571 347
rect 631 343 635 347
rect 687 343 691 347
rect 751 343 755 347
rect 815 343 819 347
rect 879 343 883 347
rect 951 343 955 347
rect 1031 343 1035 347
rect 1071 351 1075 355
rect 1103 343 1107 347
rect 1175 343 1179 347
rect 1247 343 1251 347
rect 111 327 115 331
rect 311 331 315 335
rect 351 331 352 335
rect 352 331 355 335
rect 135 325 139 329
rect 175 325 179 329
rect 223 325 227 329
rect 279 325 283 329
rect 335 325 339 329
rect 391 325 395 329
rect 447 325 451 329
rect 503 325 507 329
rect 567 325 571 329
rect 631 325 635 329
rect 687 325 691 329
rect 751 325 755 329
rect 439 319 443 323
rect 111 309 115 313
rect 191 311 195 315
rect 223 311 227 315
rect 255 311 259 315
rect 295 311 299 315
rect 335 311 339 315
rect 367 311 371 315
rect 407 311 411 315
rect 455 311 459 315
rect 519 311 523 315
rect 575 319 579 323
rect 815 325 819 329
rect 879 325 883 329
rect 951 325 955 329
rect 1031 325 1035 329
rect 1103 325 1107 329
rect 827 319 831 323
rect 1239 331 1243 335
rect 1327 343 1331 347
rect 1355 347 1359 351
rect 1407 343 1411 347
rect 1487 343 1491 347
rect 1499 347 1503 351
rect 1543 343 1547 347
rect 1583 344 1587 348
rect 1427 331 1428 335
rect 1428 331 1431 335
rect 1531 335 1535 339
rect 1175 325 1179 329
rect 1247 325 1251 329
rect 1327 325 1331 329
rect 1407 325 1411 329
rect 1487 325 1491 329
rect 1543 325 1547 329
rect 1583 327 1587 331
rect 591 311 595 315
rect 663 311 667 315
rect 735 311 739 315
rect 807 311 811 315
rect 879 311 883 315
rect 951 311 955 315
rect 1023 311 1027 315
rect 1095 311 1099 315
rect 1111 311 1115 315
rect 171 303 175 307
rect 111 292 115 296
rect 191 293 195 297
rect 223 293 227 297
rect 255 293 259 297
rect 295 293 299 297
rect 335 293 339 297
rect 367 293 371 297
rect 311 287 312 291
rect 312 287 315 291
rect 343 287 347 291
rect 399 303 403 307
rect 407 293 411 297
rect 439 287 443 291
rect 455 293 459 297
rect 519 293 523 297
rect 591 293 595 297
rect 655 295 659 299
rect 663 293 667 297
rect 723 303 727 307
rect 735 293 739 297
rect 807 293 811 297
rect 827 287 828 291
rect 828 287 831 291
rect 879 293 883 297
rect 951 293 955 297
rect 1023 293 1027 297
rect 1167 311 1171 315
rect 1231 311 1235 315
rect 1295 311 1299 315
rect 1351 311 1355 315
rect 1399 311 1403 315
rect 1455 311 1459 315
rect 1511 311 1515 315
rect 1543 311 1547 315
rect 1583 309 1587 313
rect 1095 293 1099 297
rect 1167 293 1171 297
rect 1231 293 1235 297
rect 1239 287 1243 291
rect 1287 303 1291 307
rect 1295 293 1299 297
rect 1351 293 1355 297
rect 1399 293 1403 297
rect 1499 303 1503 307
rect 1455 293 1459 297
rect 1511 293 1515 297
rect 1543 293 1547 297
rect 1531 287 1532 291
rect 1532 287 1535 291
rect 1559 303 1560 307
rect 1560 303 1563 307
rect 1583 292 1587 296
rect 495 279 499 283
rect 723 279 727 283
rect 1111 279 1115 283
rect 111 268 115 272
rect 151 267 155 271
rect 171 271 172 275
rect 172 271 175 275
rect 183 267 187 271
rect 111 251 115 255
rect 215 267 219 271
rect 247 267 251 271
rect 267 271 268 275
rect 268 271 271 275
rect 279 267 283 271
rect 311 267 315 271
rect 351 267 355 271
rect 399 271 403 275
rect 407 267 411 271
rect 479 267 483 271
rect 559 267 563 271
rect 647 267 651 271
rect 735 267 739 271
rect 823 267 827 271
rect 903 267 907 271
rect 983 267 987 271
rect 1055 267 1059 271
rect 1119 267 1123 271
rect 1175 267 1179 271
rect 1223 267 1227 271
rect 1287 279 1291 283
rect 1263 267 1267 271
rect 1303 267 1307 271
rect 1351 267 1355 271
rect 1399 267 1403 271
rect 227 255 231 259
rect 343 255 347 259
rect 151 249 155 253
rect 183 249 187 253
rect 215 249 219 253
rect 247 249 251 253
rect 279 249 283 253
rect 311 249 315 253
rect 351 249 355 253
rect 407 249 411 253
rect 479 249 483 253
rect 559 249 563 253
rect 647 249 651 253
rect 735 249 739 253
rect 463 243 467 247
rect 111 233 115 237
rect 135 235 139 239
rect 167 235 171 239
rect 207 235 211 239
rect 255 235 259 239
rect 303 235 307 239
rect 343 235 347 239
rect 383 235 387 239
rect 439 235 443 239
rect 511 235 515 239
rect 591 235 595 239
rect 655 243 659 247
rect 1187 255 1191 259
rect 1363 255 1367 259
rect 1447 267 1451 271
rect 1503 267 1507 271
rect 1519 271 1520 275
rect 1520 271 1523 275
rect 1543 267 1547 271
rect 1559 271 1560 275
rect 1560 271 1563 275
rect 1583 268 1587 272
rect 1559 255 1560 259
rect 1560 255 1563 259
rect 823 249 827 253
rect 903 249 907 253
rect 983 249 987 253
rect 1055 249 1059 253
rect 1119 249 1123 253
rect 1175 249 1179 253
rect 1223 249 1227 253
rect 1263 249 1267 253
rect 1303 249 1307 253
rect 1351 249 1355 253
rect 1399 249 1403 253
rect 1447 249 1451 253
rect 1503 249 1507 253
rect 1543 249 1547 253
rect 1583 251 1587 255
rect 679 235 683 239
rect 151 227 152 231
rect 152 227 155 231
rect 111 216 115 220
rect 135 217 139 221
rect 167 217 171 221
rect 267 227 271 231
rect 207 217 211 221
rect 255 217 259 221
rect 227 211 228 215
rect 228 211 231 215
rect 303 217 307 221
rect 399 227 400 231
rect 400 227 403 231
rect 343 217 347 221
rect 383 217 387 221
rect 375 211 379 215
rect 439 217 443 221
rect 759 235 763 239
rect 767 235 771 239
rect 847 235 851 239
rect 919 235 923 239
rect 983 235 987 239
rect 1047 235 1051 239
rect 1103 235 1107 239
rect 1159 235 1163 239
rect 1215 235 1219 239
rect 1271 235 1275 239
rect 1327 235 1331 239
rect 1383 235 1387 239
rect 1439 235 1443 239
rect 1503 235 1507 239
rect 1543 235 1547 239
rect 1583 233 1587 237
rect 511 217 515 221
rect 591 217 595 221
rect 555 211 559 215
rect 679 217 683 221
rect 767 217 771 221
rect 847 217 851 221
rect 919 217 923 221
rect 111 192 115 196
rect 135 191 139 195
rect 151 195 152 199
rect 152 195 155 199
rect 167 191 171 195
rect 215 191 219 195
rect 1023 227 1027 231
rect 1031 227 1035 231
rect 983 217 987 221
rect 1047 217 1051 221
rect 1103 217 1107 221
rect 1247 227 1251 231
rect 1159 217 1163 221
rect 1215 217 1219 221
rect 1187 211 1191 215
rect 1271 217 1275 221
rect 1327 217 1331 221
rect 1383 217 1387 221
rect 1363 211 1367 215
rect 1439 217 1443 221
rect 1031 203 1035 207
rect 1303 203 1307 207
rect 1519 227 1520 231
rect 1520 227 1523 231
rect 1503 217 1507 221
rect 1543 217 1547 221
rect 1583 216 1587 220
rect 1559 211 1560 215
rect 1560 211 1563 215
rect 1471 203 1475 207
rect 263 191 267 195
rect 311 191 315 195
rect 323 195 327 199
rect 359 191 363 195
rect 415 191 419 195
rect 463 195 467 199
rect 471 191 475 195
rect 535 191 539 195
rect 607 191 611 195
rect 619 195 623 199
rect 679 191 683 195
rect 751 191 755 195
rect 815 191 819 195
rect 871 195 875 199
rect 879 191 883 195
rect 943 191 947 195
rect 1007 191 1011 195
rect 1023 195 1024 199
rect 1024 195 1027 199
rect 1063 191 1067 195
rect 1119 191 1123 195
rect 1175 191 1179 195
rect 1231 191 1235 195
rect 1247 195 1248 199
rect 1248 195 1251 199
rect 1287 191 1291 195
rect 1343 191 1347 195
rect 1363 195 1364 199
rect 1364 195 1367 199
rect 1399 191 1403 195
rect 1455 191 1459 195
rect 1511 191 1515 195
rect 1543 191 1547 195
rect 1583 192 1587 196
rect 111 175 115 179
rect 275 179 279 183
rect 375 179 376 183
rect 376 179 379 183
rect 555 179 556 183
rect 556 179 559 183
rect 767 179 768 183
rect 768 179 771 183
rect 991 179 995 183
rect 135 173 139 177
rect 167 173 171 177
rect 215 173 219 177
rect 263 173 267 177
rect 311 173 315 177
rect 359 173 363 177
rect 415 173 419 177
rect 471 173 475 177
rect 535 173 539 177
rect 607 173 611 177
rect 679 173 683 177
rect 751 173 755 177
rect 815 173 819 177
rect 879 173 883 177
rect 943 173 947 177
rect 1007 173 1011 177
rect 1063 173 1067 177
rect 1119 173 1123 177
rect 483 167 487 171
rect 111 157 115 161
rect 143 159 147 163
rect 191 159 195 163
rect 239 159 243 163
rect 295 159 299 163
rect 351 159 355 163
rect 407 159 411 163
rect 463 159 467 163
rect 519 159 523 163
rect 575 159 579 163
rect 631 159 635 163
rect 687 159 691 163
rect 155 151 159 155
rect 111 140 115 144
rect 143 141 147 145
rect 191 141 195 145
rect 323 151 327 155
rect 239 141 243 145
rect 295 141 299 145
rect 275 135 279 139
rect 351 141 355 145
rect 407 141 411 145
rect 463 141 467 145
rect 439 135 443 139
rect 483 135 484 139
rect 484 135 487 139
rect 519 141 523 145
rect 619 151 623 155
rect 575 141 579 145
rect 631 141 635 145
rect 539 127 543 131
rect 871 167 875 171
rect 1187 179 1191 183
rect 1303 179 1304 183
rect 1304 179 1307 183
rect 1471 179 1472 183
rect 1472 179 1475 183
rect 1527 179 1528 183
rect 1528 179 1531 183
rect 1175 173 1179 177
rect 1231 173 1235 177
rect 1287 173 1291 177
rect 1343 173 1347 177
rect 1399 173 1403 177
rect 1455 173 1459 177
rect 1511 173 1515 177
rect 1543 173 1547 177
rect 1583 175 1587 179
rect 743 159 747 163
rect 799 159 803 163
rect 855 159 859 163
rect 911 159 915 163
rect 975 159 979 163
rect 1039 159 1043 163
rect 1095 159 1099 163
rect 1151 159 1155 163
rect 1207 159 1211 163
rect 1255 159 1259 163
rect 1303 159 1307 163
rect 1351 159 1355 163
rect 1399 159 1403 163
rect 1455 159 1459 163
rect 1511 159 1515 163
rect 1543 159 1547 163
rect 1583 157 1587 161
rect 687 141 691 145
rect 743 141 747 145
rect 799 141 803 145
rect 855 141 859 145
rect 911 141 915 145
rect 975 141 979 145
rect 991 135 992 139
rect 992 135 995 139
rect 1039 141 1043 145
rect 1107 151 1111 155
rect 1095 141 1099 145
rect 1151 141 1155 145
rect 1187 135 1191 139
rect 1207 141 1211 145
rect 1255 141 1259 145
rect 1315 151 1319 155
rect 1363 151 1367 155
rect 1303 141 1307 145
rect 1351 141 1355 145
rect 1399 141 1403 145
rect 1455 141 1459 145
rect 1511 141 1515 145
rect 1543 141 1547 145
rect 1487 135 1491 139
rect 1527 135 1528 139
rect 1528 135 1531 139
rect 1559 151 1560 155
rect 1560 151 1563 155
rect 1583 140 1587 144
rect 1107 127 1111 131
rect 111 108 115 112
rect 135 107 139 111
rect 155 111 156 115
rect 156 111 159 115
rect 167 107 171 111
rect 199 107 203 111
rect 231 107 235 111
rect 263 107 267 111
rect 295 107 299 111
rect 327 107 331 111
rect 359 107 363 111
rect 391 107 395 111
rect 423 107 427 111
rect 455 107 459 111
rect 563 119 567 123
rect 487 107 491 111
rect 519 107 523 111
rect 551 107 555 111
rect 583 107 587 111
rect 615 107 619 111
rect 647 107 651 111
rect 679 107 683 111
rect 711 107 715 111
rect 743 107 747 111
rect 775 107 779 111
rect 807 107 811 111
rect 839 107 843 111
rect 871 107 875 111
rect 903 107 907 111
rect 943 107 947 111
rect 983 107 987 111
rect 1023 111 1027 115
rect 1315 119 1319 123
rect 1031 107 1035 111
rect 1079 107 1083 111
rect 1127 107 1131 111
rect 1175 107 1179 111
rect 1223 107 1227 111
rect 1263 107 1267 111
rect 1303 107 1307 111
rect 1343 107 1347 111
rect 1383 107 1387 111
rect 1423 107 1427 111
rect 1471 107 1475 111
rect 1511 107 1515 111
rect 111 91 115 95
rect 439 95 440 99
rect 440 95 443 99
rect 539 95 540 99
rect 540 95 543 99
rect 563 95 567 99
rect 1543 107 1547 111
rect 1559 111 1560 115
rect 1560 111 1563 115
rect 1583 108 1587 112
rect 135 89 139 93
rect 167 89 171 93
rect 199 89 203 93
rect 231 89 235 93
rect 263 89 267 93
rect 295 89 299 93
rect 327 89 331 93
rect 359 89 363 93
rect 391 89 395 93
rect 423 89 427 93
rect 455 89 459 93
rect 487 89 491 93
rect 519 89 523 93
rect 551 89 555 93
rect 583 89 587 93
rect 615 89 619 93
rect 647 89 651 93
rect 679 89 683 93
rect 711 89 715 93
rect 743 89 747 93
rect 775 89 779 93
rect 807 89 811 93
rect 839 89 843 93
rect 871 89 875 93
rect 903 89 907 93
rect 943 89 947 93
rect 983 89 987 93
rect 1031 89 1035 93
rect 1079 89 1083 93
rect 1127 89 1131 93
rect 1023 83 1027 87
rect 1487 95 1488 99
rect 1488 95 1491 99
rect 1175 89 1179 93
rect 1223 89 1227 93
rect 1263 89 1267 93
rect 1303 89 1307 93
rect 1343 89 1347 93
rect 1383 89 1387 93
rect 1423 89 1427 93
rect 1471 89 1475 93
rect 1511 89 1515 93
rect 1543 89 1547 93
rect 1583 91 1587 95
<< m3 >>
rect 111 1654 115 1655
rect 111 1649 115 1650
rect 135 1654 139 1655
rect 112 1646 114 1649
rect 135 1648 139 1650
rect 167 1654 171 1655
rect 167 1648 171 1650
rect 199 1654 203 1655
rect 199 1648 203 1650
rect 1583 1654 1587 1655
rect 1583 1649 1587 1650
rect 134 1647 140 1648
rect 110 1645 116 1646
rect 110 1641 111 1645
rect 115 1641 116 1645
rect 134 1643 135 1647
rect 139 1643 140 1647
rect 134 1642 140 1643
rect 166 1647 172 1648
rect 166 1643 167 1647
rect 171 1643 172 1647
rect 166 1642 172 1643
rect 198 1647 204 1648
rect 198 1643 199 1647
rect 203 1643 204 1647
rect 1584 1646 1586 1649
rect 198 1642 204 1643
rect 1582 1645 1588 1646
rect 110 1640 116 1641
rect 1582 1641 1583 1645
rect 1587 1641 1588 1645
rect 1582 1640 1588 1641
rect 150 1639 156 1640
rect 150 1635 151 1639
rect 155 1635 156 1639
rect 150 1634 156 1635
rect 134 1629 140 1630
rect 110 1628 116 1629
rect 110 1624 111 1628
rect 115 1624 116 1628
rect 134 1625 135 1629
rect 139 1625 140 1629
rect 134 1624 140 1625
rect 110 1623 116 1624
rect 112 1619 114 1623
rect 136 1619 138 1624
rect 111 1618 115 1619
rect 111 1613 115 1614
rect 135 1618 139 1619
rect 135 1613 139 1614
rect 112 1609 114 1613
rect 110 1608 116 1609
rect 136 1608 138 1613
rect 152 1612 154 1634
rect 166 1629 172 1630
rect 166 1625 167 1629
rect 171 1625 172 1629
rect 166 1624 172 1625
rect 198 1629 204 1630
rect 198 1625 199 1629
rect 203 1625 204 1629
rect 198 1624 204 1625
rect 1582 1628 1588 1629
rect 1582 1624 1583 1628
rect 1587 1624 1588 1628
rect 168 1619 170 1624
rect 200 1619 202 1624
rect 1582 1623 1588 1624
rect 1584 1619 1586 1623
rect 167 1618 171 1619
rect 167 1613 171 1614
rect 175 1618 179 1619
rect 175 1613 179 1614
rect 199 1618 203 1619
rect 199 1613 203 1614
rect 239 1618 243 1619
rect 239 1613 243 1614
rect 295 1618 299 1619
rect 295 1613 299 1614
rect 351 1618 355 1619
rect 351 1613 355 1614
rect 407 1618 411 1619
rect 407 1613 411 1614
rect 455 1618 459 1619
rect 455 1613 459 1614
rect 503 1618 507 1619
rect 503 1613 507 1614
rect 551 1618 555 1619
rect 551 1613 555 1614
rect 599 1618 603 1619
rect 599 1613 603 1614
rect 647 1618 651 1619
rect 647 1613 651 1614
rect 695 1618 699 1619
rect 695 1613 699 1614
rect 743 1618 747 1619
rect 743 1613 747 1614
rect 791 1618 795 1619
rect 791 1613 795 1614
rect 839 1618 843 1619
rect 839 1613 843 1614
rect 887 1618 891 1619
rect 887 1613 891 1614
rect 935 1618 939 1619
rect 935 1613 939 1614
rect 991 1618 995 1619
rect 991 1613 995 1614
rect 1047 1618 1051 1619
rect 1047 1613 1051 1614
rect 1095 1618 1099 1619
rect 1095 1613 1099 1614
rect 1143 1618 1147 1619
rect 1143 1613 1147 1614
rect 1191 1618 1195 1619
rect 1191 1613 1195 1614
rect 1239 1618 1243 1619
rect 1239 1613 1243 1614
rect 1287 1618 1291 1619
rect 1287 1613 1291 1614
rect 1327 1618 1331 1619
rect 1327 1613 1331 1614
rect 1367 1618 1371 1619
rect 1367 1613 1371 1614
rect 1407 1618 1411 1619
rect 1407 1613 1411 1614
rect 1447 1618 1451 1619
rect 1447 1613 1451 1614
rect 1479 1618 1483 1619
rect 1479 1613 1483 1614
rect 1511 1618 1515 1619
rect 1511 1613 1515 1614
rect 1543 1618 1547 1619
rect 1543 1613 1547 1614
rect 1583 1618 1587 1619
rect 1583 1613 1587 1614
rect 150 1611 156 1612
rect 110 1604 111 1608
rect 115 1604 116 1608
rect 110 1603 116 1604
rect 134 1607 140 1608
rect 134 1603 135 1607
rect 139 1603 140 1607
rect 150 1607 151 1611
rect 155 1607 156 1611
rect 176 1608 178 1613
rect 240 1608 242 1613
rect 296 1608 298 1613
rect 352 1608 354 1613
rect 398 1611 404 1612
rect 150 1606 156 1607
rect 174 1607 180 1608
rect 134 1602 140 1603
rect 174 1603 175 1607
rect 179 1603 180 1607
rect 174 1602 180 1603
rect 238 1607 244 1608
rect 238 1603 239 1607
rect 243 1603 244 1607
rect 238 1602 244 1603
rect 294 1607 300 1608
rect 294 1603 295 1607
rect 299 1603 300 1607
rect 294 1602 300 1603
rect 350 1607 356 1608
rect 350 1603 351 1607
rect 355 1603 356 1607
rect 398 1607 399 1611
rect 403 1607 404 1611
rect 408 1608 410 1613
rect 456 1608 458 1613
rect 504 1608 506 1613
rect 552 1608 554 1613
rect 600 1608 602 1613
rect 648 1608 650 1613
rect 696 1608 698 1613
rect 744 1608 746 1613
rect 792 1608 794 1613
rect 830 1611 836 1612
rect 398 1606 404 1607
rect 406 1607 412 1608
rect 350 1602 356 1603
rect 110 1591 116 1592
rect 110 1587 111 1591
rect 115 1587 116 1591
rect 110 1586 116 1587
rect 134 1589 140 1590
rect 112 1583 114 1586
rect 134 1585 135 1589
rect 139 1585 140 1589
rect 134 1584 140 1585
rect 174 1589 180 1590
rect 174 1585 175 1589
rect 179 1585 180 1589
rect 174 1584 180 1585
rect 238 1589 244 1590
rect 238 1585 239 1589
rect 243 1585 244 1589
rect 238 1584 244 1585
rect 294 1589 300 1590
rect 294 1585 295 1589
rect 299 1585 300 1589
rect 294 1584 300 1585
rect 350 1589 356 1590
rect 350 1585 351 1589
rect 355 1585 356 1589
rect 350 1584 356 1585
rect 400 1584 402 1606
rect 406 1603 407 1607
rect 411 1603 412 1607
rect 406 1602 412 1603
rect 454 1607 460 1608
rect 454 1603 455 1607
rect 459 1603 460 1607
rect 454 1602 460 1603
rect 502 1607 508 1608
rect 502 1603 503 1607
rect 507 1603 508 1607
rect 502 1602 508 1603
rect 550 1607 556 1608
rect 550 1603 551 1607
rect 555 1603 556 1607
rect 550 1602 556 1603
rect 598 1607 604 1608
rect 598 1603 599 1607
rect 603 1603 604 1607
rect 598 1602 604 1603
rect 646 1607 652 1608
rect 646 1603 647 1607
rect 651 1603 652 1607
rect 646 1602 652 1603
rect 694 1607 700 1608
rect 694 1603 695 1607
rect 699 1603 700 1607
rect 694 1602 700 1603
rect 742 1607 748 1608
rect 742 1603 743 1607
rect 747 1603 748 1607
rect 742 1602 748 1603
rect 790 1607 796 1608
rect 790 1603 791 1607
rect 795 1603 796 1607
rect 830 1607 831 1611
rect 835 1607 836 1611
rect 840 1608 842 1613
rect 888 1608 890 1613
rect 936 1608 938 1613
rect 992 1608 994 1613
rect 1048 1608 1050 1613
rect 1096 1608 1098 1613
rect 1144 1608 1146 1613
rect 1192 1608 1194 1613
rect 1202 1611 1208 1612
rect 830 1606 836 1607
rect 838 1607 844 1608
rect 790 1602 796 1603
rect 406 1589 412 1590
rect 406 1585 407 1589
rect 411 1585 412 1589
rect 406 1584 412 1585
rect 454 1589 460 1590
rect 454 1585 455 1589
rect 459 1585 460 1589
rect 454 1584 460 1585
rect 502 1589 508 1590
rect 502 1585 503 1589
rect 507 1585 508 1589
rect 502 1584 508 1585
rect 550 1589 556 1590
rect 550 1585 551 1589
rect 555 1585 556 1589
rect 550 1584 556 1585
rect 598 1589 604 1590
rect 598 1585 599 1589
rect 603 1585 604 1589
rect 598 1584 604 1585
rect 646 1589 652 1590
rect 646 1585 647 1589
rect 651 1585 652 1589
rect 646 1584 652 1585
rect 694 1589 700 1590
rect 694 1585 695 1589
rect 699 1585 700 1589
rect 694 1584 700 1585
rect 742 1589 748 1590
rect 742 1585 743 1589
rect 747 1585 748 1589
rect 742 1584 748 1585
rect 790 1589 796 1590
rect 790 1585 791 1589
rect 795 1585 796 1589
rect 790 1584 796 1585
rect 111 1582 115 1583
rect 111 1577 115 1578
rect 135 1582 139 1584
rect 135 1577 139 1578
rect 175 1582 179 1584
rect 194 1583 200 1584
rect 194 1579 195 1583
rect 199 1579 200 1583
rect 194 1578 200 1579
rect 215 1582 219 1583
rect 112 1574 114 1577
rect 175 1576 179 1578
rect 174 1575 180 1576
rect 110 1573 116 1574
rect 110 1569 111 1573
rect 115 1569 116 1573
rect 174 1571 175 1575
rect 179 1571 180 1575
rect 174 1570 180 1571
rect 110 1568 116 1569
rect 174 1557 180 1558
rect 110 1556 116 1557
rect 110 1552 111 1556
rect 115 1552 116 1556
rect 174 1553 175 1557
rect 179 1553 180 1557
rect 174 1552 180 1553
rect 196 1552 198 1578
rect 215 1576 219 1578
rect 239 1582 243 1584
rect 239 1577 243 1578
rect 255 1582 259 1583
rect 255 1576 259 1578
rect 295 1582 299 1584
rect 295 1576 299 1578
rect 343 1582 347 1583
rect 343 1576 347 1578
rect 351 1582 355 1584
rect 398 1583 404 1584
rect 351 1577 355 1578
rect 391 1582 395 1583
rect 398 1579 399 1583
rect 403 1579 404 1583
rect 398 1578 404 1579
rect 407 1582 411 1584
rect 391 1576 395 1578
rect 407 1577 411 1578
rect 439 1582 443 1583
rect 439 1576 443 1578
rect 455 1582 459 1584
rect 455 1577 459 1578
rect 487 1582 491 1583
rect 487 1576 491 1578
rect 503 1582 507 1584
rect 503 1577 507 1578
rect 535 1582 539 1583
rect 535 1576 539 1578
rect 551 1582 555 1584
rect 551 1577 555 1578
rect 583 1582 587 1583
rect 583 1576 587 1578
rect 599 1582 603 1584
rect 599 1577 603 1578
rect 639 1582 643 1583
rect 639 1576 643 1578
rect 647 1582 651 1584
rect 647 1577 651 1578
rect 695 1582 699 1584
rect 695 1577 699 1578
rect 703 1582 707 1583
rect 703 1576 707 1578
rect 743 1582 747 1584
rect 743 1577 747 1578
rect 775 1582 779 1583
rect 775 1576 779 1578
rect 791 1582 795 1584
rect 791 1577 795 1578
rect 214 1575 220 1576
rect 214 1571 215 1575
rect 219 1571 220 1575
rect 214 1570 220 1571
rect 254 1575 260 1576
rect 254 1571 255 1575
rect 259 1571 260 1575
rect 254 1570 260 1571
rect 294 1575 300 1576
rect 294 1571 295 1575
rect 299 1571 300 1575
rect 294 1570 300 1571
rect 342 1575 348 1576
rect 342 1571 343 1575
rect 347 1571 348 1575
rect 342 1570 348 1571
rect 390 1575 396 1576
rect 390 1571 391 1575
rect 395 1571 396 1575
rect 390 1570 396 1571
rect 438 1575 444 1576
rect 438 1571 439 1575
rect 443 1571 444 1575
rect 438 1570 444 1571
rect 486 1575 492 1576
rect 486 1571 487 1575
rect 491 1571 492 1575
rect 486 1570 492 1571
rect 534 1575 540 1576
rect 534 1571 535 1575
rect 539 1571 540 1575
rect 534 1570 540 1571
rect 582 1575 588 1576
rect 582 1571 583 1575
rect 587 1571 588 1575
rect 582 1570 588 1571
rect 638 1575 644 1576
rect 638 1571 639 1575
rect 643 1571 644 1575
rect 638 1570 644 1571
rect 702 1575 708 1576
rect 702 1571 703 1575
rect 707 1571 708 1575
rect 702 1570 708 1571
rect 774 1575 780 1576
rect 774 1571 775 1575
rect 779 1571 780 1575
rect 774 1570 780 1571
rect 832 1568 834 1606
rect 838 1603 839 1607
rect 843 1603 844 1607
rect 838 1602 844 1603
rect 886 1607 892 1608
rect 886 1603 887 1607
rect 891 1603 892 1607
rect 886 1602 892 1603
rect 934 1607 940 1608
rect 934 1603 935 1607
rect 939 1603 940 1607
rect 934 1602 940 1603
rect 990 1607 996 1608
rect 990 1603 991 1607
rect 995 1603 996 1607
rect 990 1602 996 1603
rect 1046 1607 1052 1608
rect 1046 1603 1047 1607
rect 1051 1603 1052 1607
rect 1046 1602 1052 1603
rect 1094 1607 1100 1608
rect 1094 1603 1095 1607
rect 1099 1603 1100 1607
rect 1094 1602 1100 1603
rect 1142 1607 1148 1608
rect 1142 1603 1143 1607
rect 1147 1603 1148 1607
rect 1142 1602 1148 1603
rect 1190 1607 1196 1608
rect 1190 1603 1191 1607
rect 1195 1603 1196 1607
rect 1202 1607 1203 1611
rect 1207 1607 1208 1611
rect 1240 1608 1242 1613
rect 1288 1608 1290 1613
rect 1328 1608 1330 1613
rect 1368 1608 1370 1613
rect 1408 1608 1410 1613
rect 1448 1608 1450 1613
rect 1480 1608 1482 1613
rect 1512 1608 1514 1613
rect 1544 1608 1546 1613
rect 1584 1609 1586 1613
rect 1582 1608 1588 1609
rect 1202 1606 1208 1607
rect 1238 1607 1244 1608
rect 1190 1602 1196 1603
rect 1158 1595 1164 1596
rect 1158 1591 1159 1595
rect 1163 1591 1164 1595
rect 1158 1590 1164 1591
rect 838 1589 844 1590
rect 838 1585 839 1589
rect 843 1585 844 1589
rect 838 1584 844 1585
rect 886 1589 892 1590
rect 886 1585 887 1589
rect 891 1585 892 1589
rect 886 1584 892 1585
rect 934 1589 940 1590
rect 934 1585 935 1589
rect 939 1585 940 1589
rect 934 1584 940 1585
rect 990 1589 996 1590
rect 990 1585 991 1589
rect 995 1585 996 1589
rect 990 1584 996 1585
rect 1046 1589 1052 1590
rect 1046 1585 1047 1589
rect 1051 1585 1052 1589
rect 1046 1584 1052 1585
rect 1094 1589 1100 1590
rect 1094 1585 1095 1589
rect 1099 1585 1100 1589
rect 1094 1584 1100 1585
rect 1142 1589 1148 1590
rect 1142 1585 1143 1589
rect 1147 1585 1148 1589
rect 1160 1587 1162 1590
rect 1142 1584 1148 1585
rect 1152 1585 1162 1587
rect 1190 1589 1196 1590
rect 1190 1585 1191 1589
rect 1195 1585 1196 1589
rect 839 1582 843 1584
rect 839 1577 843 1578
rect 855 1582 859 1583
rect 855 1576 859 1578
rect 887 1582 891 1584
rect 887 1577 891 1578
rect 935 1582 939 1584
rect 935 1576 939 1578
rect 991 1582 995 1584
rect 991 1577 995 1578
rect 1015 1582 1019 1583
rect 1015 1576 1019 1578
rect 1047 1582 1051 1584
rect 1047 1577 1051 1578
rect 1087 1582 1091 1583
rect 1087 1576 1091 1578
rect 1095 1582 1099 1584
rect 1095 1577 1099 1578
rect 1143 1582 1147 1584
rect 1143 1577 1147 1578
rect 854 1575 860 1576
rect 854 1571 855 1575
rect 859 1571 860 1575
rect 854 1570 860 1571
rect 934 1575 940 1576
rect 934 1571 935 1575
rect 939 1571 940 1575
rect 934 1570 940 1571
rect 1014 1575 1020 1576
rect 1014 1571 1015 1575
rect 1019 1571 1020 1575
rect 1014 1570 1020 1571
rect 1086 1575 1092 1576
rect 1086 1571 1087 1575
rect 1091 1571 1092 1575
rect 1086 1570 1092 1571
rect 246 1567 252 1568
rect 246 1563 247 1567
rect 251 1563 252 1567
rect 246 1562 252 1563
rect 766 1567 772 1568
rect 766 1563 767 1567
rect 771 1563 772 1567
rect 766 1562 772 1563
rect 830 1567 836 1568
rect 830 1563 831 1567
rect 835 1563 836 1567
rect 830 1562 836 1563
rect 986 1567 992 1568
rect 986 1563 987 1567
rect 991 1563 992 1567
rect 986 1562 992 1563
rect 214 1557 220 1558
rect 214 1553 215 1557
rect 219 1553 220 1557
rect 214 1552 220 1553
rect 110 1551 116 1552
rect 112 1547 114 1551
rect 176 1547 178 1552
rect 194 1551 200 1552
rect 194 1547 195 1551
rect 199 1547 200 1551
rect 216 1547 218 1552
rect 111 1546 115 1547
rect 111 1541 115 1542
rect 159 1546 163 1547
rect 159 1541 163 1542
rect 175 1546 179 1547
rect 194 1546 200 1547
rect 207 1546 211 1547
rect 175 1541 179 1542
rect 207 1541 211 1542
rect 215 1546 219 1547
rect 248 1544 250 1562
rect 254 1557 260 1558
rect 254 1553 255 1557
rect 259 1553 260 1557
rect 254 1552 260 1553
rect 294 1557 300 1558
rect 294 1553 295 1557
rect 299 1553 300 1557
rect 294 1552 300 1553
rect 342 1557 348 1558
rect 342 1553 343 1557
rect 347 1553 348 1557
rect 342 1552 348 1553
rect 390 1557 396 1558
rect 390 1553 391 1557
rect 395 1553 396 1557
rect 390 1552 396 1553
rect 438 1557 444 1558
rect 438 1553 439 1557
rect 443 1553 444 1557
rect 438 1552 444 1553
rect 486 1557 492 1558
rect 486 1553 487 1557
rect 491 1553 492 1557
rect 486 1552 492 1553
rect 534 1557 540 1558
rect 534 1553 535 1557
rect 539 1553 540 1557
rect 534 1552 540 1553
rect 582 1557 588 1558
rect 582 1553 583 1557
rect 587 1553 588 1557
rect 582 1552 588 1553
rect 638 1557 644 1558
rect 638 1553 639 1557
rect 643 1553 644 1557
rect 638 1552 644 1553
rect 702 1557 708 1558
rect 702 1553 703 1557
rect 707 1553 708 1557
rect 702 1552 708 1553
rect 256 1547 258 1552
rect 296 1547 298 1552
rect 344 1547 346 1552
rect 392 1547 394 1552
rect 440 1547 442 1552
rect 488 1547 490 1552
rect 536 1547 538 1552
rect 584 1547 586 1552
rect 640 1547 642 1552
rect 704 1547 706 1552
rect 255 1546 259 1547
rect 215 1541 219 1542
rect 246 1543 252 1544
rect 112 1537 114 1541
rect 110 1536 116 1537
rect 160 1536 162 1541
rect 208 1536 210 1541
rect 246 1539 247 1543
rect 251 1539 252 1543
rect 255 1541 259 1542
rect 295 1546 299 1547
rect 295 1541 299 1542
rect 311 1546 315 1547
rect 311 1541 315 1542
rect 343 1546 347 1547
rect 343 1541 347 1542
rect 359 1546 363 1547
rect 359 1541 363 1542
rect 391 1546 395 1547
rect 391 1541 395 1542
rect 415 1546 419 1547
rect 415 1541 419 1542
rect 439 1546 443 1547
rect 439 1541 443 1542
rect 471 1546 475 1547
rect 471 1541 475 1542
rect 487 1546 491 1547
rect 487 1541 491 1542
rect 527 1546 531 1547
rect 527 1541 531 1542
rect 535 1546 539 1547
rect 535 1541 539 1542
rect 583 1546 587 1547
rect 583 1541 587 1542
rect 639 1546 643 1547
rect 639 1541 643 1542
rect 695 1546 699 1547
rect 695 1541 699 1542
rect 703 1546 707 1547
rect 703 1541 707 1542
rect 759 1546 763 1547
rect 768 1544 770 1562
rect 774 1557 780 1558
rect 774 1553 775 1557
rect 779 1553 780 1557
rect 774 1552 780 1553
rect 854 1557 860 1558
rect 854 1553 855 1557
rect 859 1553 860 1557
rect 854 1552 860 1553
rect 934 1557 940 1558
rect 934 1553 935 1557
rect 939 1553 940 1557
rect 934 1552 940 1553
rect 776 1547 778 1552
rect 856 1547 858 1552
rect 914 1551 920 1552
rect 914 1547 915 1551
rect 919 1547 920 1551
rect 936 1547 938 1552
rect 775 1546 779 1547
rect 759 1541 763 1542
rect 766 1543 772 1544
rect 246 1538 252 1539
rect 256 1536 258 1541
rect 312 1536 314 1541
rect 360 1536 362 1541
rect 370 1539 376 1540
rect 110 1532 111 1536
rect 115 1532 116 1536
rect 110 1531 116 1532
rect 158 1535 164 1536
rect 158 1531 159 1535
rect 163 1531 164 1535
rect 158 1530 164 1531
rect 206 1535 212 1536
rect 206 1531 207 1535
rect 211 1531 212 1535
rect 206 1530 212 1531
rect 254 1535 260 1536
rect 254 1531 255 1535
rect 259 1531 260 1535
rect 254 1530 260 1531
rect 310 1535 316 1536
rect 310 1531 311 1535
rect 315 1531 316 1535
rect 310 1530 316 1531
rect 358 1535 364 1536
rect 358 1531 359 1535
rect 363 1531 364 1535
rect 370 1535 371 1539
rect 375 1535 376 1539
rect 416 1536 418 1541
rect 472 1536 474 1541
rect 528 1536 530 1541
rect 584 1536 586 1541
rect 640 1536 642 1541
rect 696 1536 698 1541
rect 760 1536 762 1541
rect 766 1539 767 1543
rect 771 1539 772 1543
rect 775 1541 779 1542
rect 823 1546 827 1547
rect 823 1541 827 1542
rect 855 1546 859 1547
rect 855 1541 859 1542
rect 895 1546 899 1547
rect 914 1546 920 1547
rect 935 1546 939 1547
rect 895 1541 899 1542
rect 766 1538 772 1539
rect 824 1536 826 1541
rect 896 1536 898 1541
rect 370 1534 376 1535
rect 414 1535 420 1536
rect 358 1530 364 1531
rect 174 1523 180 1524
rect 110 1519 116 1520
rect 110 1515 111 1519
rect 115 1515 116 1519
rect 174 1519 175 1523
rect 179 1519 180 1523
rect 174 1518 180 1519
rect 110 1514 116 1515
rect 158 1517 164 1518
rect 112 1511 114 1514
rect 158 1513 159 1517
rect 163 1513 164 1517
rect 158 1512 164 1513
rect 111 1510 115 1511
rect 111 1505 115 1506
rect 159 1510 163 1512
rect 112 1502 114 1505
rect 159 1504 163 1506
rect 158 1503 164 1504
rect 110 1501 116 1502
rect 110 1497 111 1501
rect 115 1497 116 1501
rect 158 1499 159 1503
rect 163 1499 164 1503
rect 158 1498 164 1499
rect 110 1496 116 1497
rect 158 1485 164 1486
rect 110 1484 116 1485
rect 110 1480 111 1484
rect 115 1480 116 1484
rect 158 1481 159 1485
rect 163 1481 164 1485
rect 158 1480 164 1481
rect 176 1480 178 1518
rect 206 1517 212 1518
rect 206 1513 207 1517
rect 211 1513 212 1517
rect 206 1512 212 1513
rect 254 1517 260 1518
rect 254 1513 255 1517
rect 259 1513 260 1517
rect 254 1512 260 1513
rect 310 1517 316 1518
rect 310 1513 311 1517
rect 315 1513 316 1517
rect 310 1512 316 1513
rect 358 1517 364 1518
rect 358 1513 359 1517
rect 363 1513 364 1517
rect 358 1512 364 1513
rect 207 1510 211 1512
rect 207 1504 211 1506
rect 255 1510 259 1512
rect 255 1504 259 1506
rect 303 1510 307 1511
rect 303 1504 307 1506
rect 311 1510 315 1512
rect 311 1505 315 1506
rect 351 1510 355 1511
rect 351 1504 355 1506
rect 359 1510 363 1512
rect 359 1505 363 1506
rect 206 1503 212 1504
rect 206 1499 207 1503
rect 211 1499 212 1503
rect 206 1498 212 1499
rect 254 1503 260 1504
rect 254 1499 255 1503
rect 259 1499 260 1503
rect 254 1498 260 1499
rect 302 1503 308 1504
rect 302 1499 303 1503
rect 307 1499 308 1503
rect 302 1498 308 1499
rect 350 1503 356 1504
rect 350 1499 351 1503
rect 355 1499 356 1503
rect 350 1498 356 1499
rect 372 1496 374 1534
rect 414 1531 415 1535
rect 419 1531 420 1535
rect 414 1530 420 1531
rect 470 1535 476 1536
rect 470 1531 471 1535
rect 475 1531 476 1535
rect 470 1530 476 1531
rect 526 1535 532 1536
rect 526 1531 527 1535
rect 531 1531 532 1535
rect 526 1530 532 1531
rect 582 1535 588 1536
rect 582 1531 583 1535
rect 587 1531 588 1535
rect 582 1530 588 1531
rect 638 1535 644 1536
rect 638 1531 639 1535
rect 643 1531 644 1535
rect 638 1530 644 1531
rect 694 1535 700 1536
rect 694 1531 695 1535
rect 699 1531 700 1535
rect 694 1530 700 1531
rect 758 1535 764 1536
rect 758 1531 759 1535
rect 763 1531 764 1535
rect 758 1530 764 1531
rect 774 1535 780 1536
rect 774 1531 775 1535
rect 779 1531 780 1535
rect 774 1530 780 1531
rect 822 1535 828 1536
rect 822 1531 823 1535
rect 827 1531 828 1535
rect 822 1530 828 1531
rect 894 1535 900 1536
rect 894 1531 895 1535
rect 899 1531 900 1535
rect 894 1530 900 1531
rect 414 1517 420 1518
rect 414 1513 415 1517
rect 419 1513 420 1517
rect 414 1512 420 1513
rect 470 1517 476 1518
rect 470 1513 471 1517
rect 475 1513 476 1517
rect 470 1512 476 1513
rect 526 1517 532 1518
rect 526 1513 527 1517
rect 531 1513 532 1517
rect 526 1512 532 1513
rect 582 1517 588 1518
rect 582 1513 583 1517
rect 587 1513 588 1517
rect 582 1512 588 1513
rect 638 1517 644 1518
rect 638 1513 639 1517
rect 643 1513 644 1517
rect 638 1512 644 1513
rect 694 1517 700 1518
rect 694 1513 695 1517
rect 699 1513 700 1517
rect 694 1512 700 1513
rect 758 1517 764 1518
rect 758 1513 759 1517
rect 763 1513 764 1517
rect 758 1512 764 1513
rect 407 1510 411 1511
rect 407 1504 411 1506
rect 415 1510 419 1512
rect 415 1505 419 1506
rect 463 1510 467 1511
rect 463 1504 467 1506
rect 471 1510 475 1512
rect 482 1511 488 1512
rect 482 1507 483 1511
rect 487 1507 488 1511
rect 482 1506 488 1507
rect 527 1510 531 1512
rect 471 1505 475 1506
rect 406 1503 412 1504
rect 406 1499 407 1503
rect 411 1499 412 1503
rect 406 1498 412 1499
rect 462 1503 468 1504
rect 462 1499 463 1503
rect 467 1499 468 1503
rect 462 1498 468 1499
rect 218 1495 224 1496
rect 218 1491 219 1495
rect 223 1491 224 1495
rect 218 1490 224 1491
rect 370 1495 376 1496
rect 370 1491 371 1495
rect 375 1491 376 1495
rect 370 1490 376 1491
rect 206 1485 212 1486
rect 206 1481 207 1485
rect 211 1481 212 1485
rect 206 1480 212 1481
rect 110 1479 116 1480
rect 112 1475 114 1479
rect 160 1475 162 1480
rect 174 1479 180 1480
rect 174 1475 175 1479
rect 179 1475 180 1479
rect 208 1475 210 1480
rect 111 1474 115 1475
rect 111 1469 115 1470
rect 135 1474 139 1475
rect 135 1469 139 1470
rect 159 1474 163 1475
rect 174 1474 180 1475
rect 183 1474 187 1475
rect 159 1469 163 1470
rect 183 1469 187 1470
rect 207 1474 211 1475
rect 207 1469 211 1470
rect 112 1465 114 1469
rect 110 1464 116 1465
rect 136 1464 138 1469
rect 184 1464 186 1469
rect 220 1468 222 1490
rect 254 1485 260 1486
rect 254 1481 255 1485
rect 259 1481 260 1485
rect 254 1480 260 1481
rect 302 1485 308 1486
rect 302 1481 303 1485
rect 307 1481 308 1485
rect 302 1480 308 1481
rect 350 1485 356 1486
rect 350 1481 351 1485
rect 355 1481 356 1485
rect 350 1480 356 1481
rect 406 1485 412 1486
rect 406 1481 407 1485
rect 411 1481 412 1485
rect 406 1480 412 1481
rect 462 1485 468 1486
rect 462 1481 463 1485
rect 467 1481 468 1485
rect 462 1480 468 1481
rect 256 1475 258 1480
rect 274 1479 280 1480
rect 274 1475 275 1479
rect 279 1475 280 1479
rect 304 1475 306 1480
rect 352 1475 354 1480
rect 408 1475 410 1480
rect 464 1475 466 1480
rect 231 1474 235 1475
rect 231 1469 235 1470
rect 255 1474 259 1475
rect 274 1474 280 1475
rect 287 1474 291 1475
rect 255 1469 259 1470
rect 218 1467 224 1468
rect 110 1460 111 1464
rect 115 1460 116 1464
rect 110 1459 116 1460
rect 134 1463 140 1464
rect 134 1459 135 1463
rect 139 1459 140 1463
rect 134 1458 140 1459
rect 182 1463 188 1464
rect 182 1459 183 1463
rect 187 1459 188 1463
rect 218 1463 219 1467
rect 223 1463 224 1467
rect 232 1464 234 1469
rect 218 1462 224 1463
rect 230 1463 236 1464
rect 182 1458 188 1459
rect 230 1459 231 1463
rect 235 1459 236 1463
rect 230 1458 236 1459
rect 258 1463 264 1464
rect 258 1458 259 1463
rect 263 1458 264 1463
rect 259 1455 263 1456
rect 150 1451 156 1452
rect 110 1447 116 1448
rect 110 1443 111 1447
rect 115 1443 116 1447
rect 150 1447 151 1451
rect 155 1447 156 1451
rect 150 1446 156 1447
rect 110 1442 116 1443
rect 134 1445 140 1446
rect 112 1439 114 1442
rect 134 1441 135 1445
rect 139 1441 140 1445
rect 134 1440 140 1441
rect 111 1438 115 1439
rect 111 1433 115 1434
rect 135 1438 139 1440
rect 112 1430 114 1433
rect 135 1432 139 1434
rect 134 1431 140 1432
rect 110 1429 116 1430
rect 110 1425 111 1429
rect 115 1425 116 1429
rect 134 1427 135 1431
rect 139 1427 140 1431
rect 134 1426 140 1427
rect 110 1424 116 1425
rect 134 1413 140 1414
rect 110 1412 116 1413
rect 110 1408 111 1412
rect 115 1408 116 1412
rect 134 1409 135 1413
rect 139 1409 140 1413
rect 134 1408 140 1409
rect 152 1408 154 1446
rect 182 1445 188 1446
rect 182 1441 183 1445
rect 187 1441 188 1445
rect 182 1440 188 1441
rect 230 1445 236 1446
rect 230 1441 231 1445
rect 235 1441 236 1445
rect 230 1440 236 1441
rect 276 1440 278 1474
rect 287 1469 291 1470
rect 303 1474 307 1475
rect 303 1469 307 1470
rect 343 1474 347 1475
rect 343 1469 347 1470
rect 351 1474 355 1475
rect 351 1469 355 1470
rect 399 1474 403 1475
rect 399 1469 403 1470
rect 407 1474 411 1475
rect 407 1469 411 1470
rect 455 1474 459 1475
rect 455 1469 459 1470
rect 463 1474 467 1475
rect 463 1469 467 1470
rect 288 1464 290 1469
rect 344 1464 346 1469
rect 400 1464 402 1469
rect 456 1464 458 1469
rect 484 1468 486 1506
rect 527 1504 531 1506
rect 583 1510 587 1512
rect 583 1505 587 1506
rect 591 1510 595 1511
rect 591 1504 595 1506
rect 639 1510 643 1512
rect 639 1505 643 1506
rect 655 1510 659 1511
rect 655 1504 659 1506
rect 695 1510 699 1512
rect 695 1505 699 1506
rect 719 1510 723 1511
rect 719 1504 723 1506
rect 759 1510 763 1512
rect 759 1505 763 1506
rect 526 1503 532 1504
rect 526 1499 527 1503
rect 531 1499 532 1503
rect 526 1498 532 1499
rect 590 1503 596 1504
rect 590 1499 591 1503
rect 595 1499 596 1503
rect 590 1498 596 1499
rect 654 1503 660 1504
rect 654 1499 655 1503
rect 659 1499 660 1503
rect 654 1498 660 1499
rect 718 1503 724 1504
rect 718 1499 719 1503
rect 723 1499 724 1503
rect 718 1498 724 1499
rect 776 1496 778 1530
rect 916 1524 918 1546
rect 935 1541 939 1542
rect 967 1546 971 1547
rect 967 1541 971 1542
rect 968 1536 970 1541
rect 988 1540 990 1562
rect 1014 1557 1020 1558
rect 1014 1553 1015 1557
rect 1019 1553 1020 1557
rect 1014 1552 1020 1553
rect 1086 1557 1092 1558
rect 1086 1553 1087 1557
rect 1091 1553 1092 1557
rect 1086 1552 1092 1553
rect 1152 1552 1154 1585
rect 1190 1584 1196 1585
rect 1159 1582 1163 1583
rect 1159 1576 1163 1578
rect 1191 1582 1195 1584
rect 1191 1577 1195 1578
rect 1158 1575 1164 1576
rect 1158 1571 1159 1575
rect 1163 1571 1164 1575
rect 1158 1570 1164 1571
rect 1204 1568 1206 1606
rect 1238 1603 1239 1607
rect 1243 1603 1244 1607
rect 1238 1602 1244 1603
rect 1286 1607 1292 1608
rect 1286 1603 1287 1607
rect 1291 1603 1292 1607
rect 1286 1602 1292 1603
rect 1326 1607 1332 1608
rect 1326 1603 1327 1607
rect 1331 1603 1332 1607
rect 1326 1602 1332 1603
rect 1366 1607 1372 1608
rect 1366 1603 1367 1607
rect 1371 1603 1372 1607
rect 1366 1602 1372 1603
rect 1406 1607 1412 1608
rect 1406 1603 1407 1607
rect 1411 1603 1412 1607
rect 1406 1602 1412 1603
rect 1446 1607 1452 1608
rect 1446 1603 1447 1607
rect 1451 1603 1452 1607
rect 1446 1602 1452 1603
rect 1478 1607 1484 1608
rect 1478 1603 1479 1607
rect 1483 1603 1484 1607
rect 1478 1602 1484 1603
rect 1510 1607 1516 1608
rect 1510 1603 1511 1607
rect 1515 1603 1516 1607
rect 1510 1602 1516 1603
rect 1542 1607 1548 1608
rect 1542 1603 1543 1607
rect 1547 1603 1548 1607
rect 1582 1604 1583 1608
rect 1587 1604 1588 1608
rect 1582 1603 1588 1604
rect 1542 1602 1548 1603
rect 1582 1591 1588 1592
rect 1238 1589 1244 1590
rect 1238 1585 1239 1589
rect 1243 1585 1244 1589
rect 1238 1584 1244 1585
rect 1286 1589 1292 1590
rect 1286 1585 1287 1589
rect 1291 1585 1292 1589
rect 1286 1584 1292 1585
rect 1326 1589 1332 1590
rect 1326 1585 1327 1589
rect 1331 1585 1332 1589
rect 1326 1584 1332 1585
rect 1366 1589 1372 1590
rect 1366 1585 1367 1589
rect 1371 1585 1372 1589
rect 1366 1584 1372 1585
rect 1406 1589 1412 1590
rect 1406 1585 1407 1589
rect 1411 1585 1412 1589
rect 1406 1584 1412 1585
rect 1446 1589 1452 1590
rect 1446 1585 1447 1589
rect 1451 1585 1452 1589
rect 1446 1584 1452 1585
rect 1478 1589 1484 1590
rect 1478 1585 1479 1589
rect 1483 1585 1484 1589
rect 1478 1584 1484 1585
rect 1510 1589 1516 1590
rect 1510 1585 1511 1589
rect 1515 1585 1516 1589
rect 1510 1584 1516 1585
rect 1542 1589 1548 1590
rect 1542 1585 1543 1589
rect 1547 1585 1548 1589
rect 1582 1587 1583 1591
rect 1587 1587 1588 1591
rect 1582 1586 1588 1587
rect 1542 1584 1548 1585
rect 1239 1582 1243 1584
rect 1239 1576 1243 1578
rect 1287 1582 1291 1584
rect 1287 1577 1291 1578
rect 1319 1582 1323 1583
rect 1319 1576 1323 1578
rect 1327 1582 1331 1584
rect 1327 1577 1331 1578
rect 1367 1582 1371 1584
rect 1367 1577 1371 1578
rect 1399 1582 1403 1583
rect 1399 1576 1403 1578
rect 1407 1582 1411 1584
rect 1407 1577 1411 1578
rect 1447 1582 1451 1584
rect 1447 1577 1451 1578
rect 1479 1582 1483 1584
rect 1498 1583 1504 1584
rect 1498 1579 1499 1583
rect 1503 1579 1504 1583
rect 1498 1578 1504 1579
rect 1511 1582 1515 1584
rect 1479 1576 1483 1578
rect 1238 1575 1244 1576
rect 1238 1571 1239 1575
rect 1243 1571 1244 1575
rect 1238 1570 1244 1571
rect 1318 1575 1324 1576
rect 1318 1571 1319 1575
rect 1323 1571 1324 1575
rect 1318 1570 1324 1571
rect 1398 1575 1404 1576
rect 1398 1571 1399 1575
rect 1403 1571 1404 1575
rect 1398 1570 1404 1571
rect 1478 1575 1484 1576
rect 1478 1571 1479 1575
rect 1483 1571 1484 1575
rect 1478 1570 1484 1571
rect 1202 1567 1208 1568
rect 1202 1563 1203 1567
rect 1207 1563 1208 1567
rect 1202 1562 1208 1563
rect 1158 1557 1164 1558
rect 1158 1553 1159 1557
rect 1163 1553 1164 1557
rect 1158 1552 1164 1553
rect 1238 1557 1244 1558
rect 1238 1553 1239 1557
rect 1243 1553 1244 1557
rect 1238 1552 1244 1553
rect 1318 1557 1324 1558
rect 1318 1553 1319 1557
rect 1323 1553 1324 1557
rect 1318 1552 1324 1553
rect 1398 1557 1404 1558
rect 1398 1553 1399 1557
rect 1403 1553 1404 1557
rect 1398 1552 1404 1553
rect 1478 1557 1484 1558
rect 1478 1553 1479 1557
rect 1483 1553 1484 1557
rect 1500 1556 1502 1578
rect 1511 1577 1515 1578
rect 1543 1582 1547 1584
rect 1584 1583 1586 1586
rect 1543 1576 1547 1578
rect 1583 1582 1587 1583
rect 1583 1577 1587 1578
rect 1542 1575 1548 1576
rect 1542 1571 1543 1575
rect 1547 1571 1548 1575
rect 1584 1574 1586 1577
rect 1542 1570 1548 1571
rect 1582 1573 1588 1574
rect 1582 1569 1583 1573
rect 1587 1569 1588 1573
rect 1582 1568 1588 1569
rect 1558 1567 1564 1568
rect 1558 1563 1559 1567
rect 1563 1563 1564 1567
rect 1558 1562 1564 1563
rect 1542 1557 1548 1558
rect 1478 1552 1484 1553
rect 1498 1555 1504 1556
rect 1016 1547 1018 1552
rect 1088 1547 1090 1552
rect 1150 1551 1156 1552
rect 1150 1547 1151 1551
rect 1155 1547 1156 1551
rect 1160 1547 1162 1552
rect 1240 1547 1242 1552
rect 1320 1547 1322 1552
rect 1326 1551 1332 1552
rect 1326 1547 1327 1551
rect 1331 1547 1332 1551
rect 1400 1547 1402 1552
rect 1480 1547 1482 1552
rect 1498 1551 1499 1555
rect 1503 1551 1504 1555
rect 1542 1553 1543 1557
rect 1547 1553 1548 1557
rect 1542 1552 1548 1553
rect 1498 1550 1504 1551
rect 1544 1547 1546 1552
rect 1015 1546 1019 1547
rect 1015 1541 1019 1542
rect 1039 1546 1043 1547
rect 1039 1541 1043 1542
rect 1087 1546 1091 1547
rect 1087 1541 1091 1542
rect 1103 1546 1107 1547
rect 1150 1546 1156 1547
rect 1159 1546 1163 1547
rect 1103 1541 1107 1542
rect 1159 1541 1163 1542
rect 1167 1546 1171 1547
rect 1167 1541 1171 1542
rect 1231 1546 1235 1547
rect 1231 1541 1235 1542
rect 1239 1546 1243 1547
rect 1239 1541 1243 1542
rect 1295 1546 1299 1547
rect 1295 1541 1299 1542
rect 1319 1546 1323 1547
rect 1326 1546 1332 1547
rect 1359 1546 1363 1547
rect 1319 1541 1323 1542
rect 986 1539 992 1540
rect 966 1535 972 1536
rect 966 1531 967 1535
rect 971 1531 972 1535
rect 986 1535 987 1539
rect 991 1535 992 1539
rect 1040 1536 1042 1541
rect 1104 1536 1106 1541
rect 1168 1536 1170 1541
rect 1222 1539 1228 1540
rect 986 1534 992 1535
rect 1038 1535 1044 1536
rect 966 1530 972 1531
rect 1038 1531 1039 1535
rect 1043 1531 1044 1535
rect 1038 1530 1044 1531
rect 1102 1535 1108 1536
rect 1102 1531 1103 1535
rect 1107 1531 1108 1535
rect 1102 1530 1108 1531
rect 1166 1535 1172 1536
rect 1166 1531 1167 1535
rect 1171 1531 1172 1535
rect 1222 1535 1223 1539
rect 1227 1535 1228 1539
rect 1232 1536 1234 1541
rect 1296 1536 1298 1541
rect 1222 1534 1228 1535
rect 1230 1535 1236 1536
rect 1166 1530 1172 1531
rect 914 1523 920 1524
rect 914 1519 915 1523
rect 919 1519 920 1523
rect 914 1518 920 1519
rect 1114 1523 1120 1524
rect 1114 1519 1115 1523
rect 1119 1519 1120 1523
rect 1114 1518 1120 1519
rect 822 1517 828 1518
rect 822 1513 823 1517
rect 827 1513 828 1517
rect 822 1512 828 1513
rect 894 1517 900 1518
rect 894 1513 895 1517
rect 899 1513 900 1517
rect 894 1512 900 1513
rect 966 1517 972 1518
rect 966 1513 967 1517
rect 971 1513 972 1517
rect 966 1512 972 1513
rect 1038 1517 1044 1518
rect 1038 1513 1039 1517
rect 1043 1513 1044 1517
rect 1038 1512 1044 1513
rect 1102 1517 1108 1518
rect 1102 1513 1103 1517
rect 1107 1513 1108 1517
rect 1102 1512 1108 1513
rect 783 1510 787 1511
rect 783 1504 787 1506
rect 823 1510 827 1512
rect 823 1505 827 1506
rect 855 1510 859 1511
rect 855 1504 859 1506
rect 895 1510 899 1512
rect 895 1505 899 1506
rect 935 1510 939 1511
rect 935 1504 939 1506
rect 967 1510 971 1512
rect 967 1505 971 1506
rect 1007 1510 1011 1511
rect 1007 1504 1011 1506
rect 1039 1510 1043 1512
rect 1039 1505 1043 1506
rect 1079 1510 1083 1511
rect 1079 1504 1083 1506
rect 1103 1510 1107 1512
rect 1103 1505 1107 1506
rect 782 1503 788 1504
rect 782 1499 783 1503
rect 787 1499 788 1503
rect 782 1498 788 1499
rect 854 1503 860 1504
rect 854 1499 855 1503
rect 859 1499 860 1503
rect 854 1498 860 1499
rect 934 1503 940 1504
rect 934 1499 935 1503
rect 939 1499 940 1503
rect 934 1498 940 1499
rect 1006 1503 1012 1504
rect 1006 1499 1007 1503
rect 1011 1499 1012 1503
rect 1006 1498 1012 1499
rect 1078 1503 1084 1504
rect 1078 1499 1079 1503
rect 1083 1499 1084 1503
rect 1078 1498 1084 1499
rect 774 1495 780 1496
rect 774 1491 775 1495
rect 779 1491 780 1495
rect 774 1490 780 1491
rect 898 1495 904 1496
rect 898 1491 899 1495
rect 903 1491 904 1495
rect 898 1490 904 1491
rect 526 1485 532 1486
rect 526 1481 527 1485
rect 531 1481 532 1485
rect 526 1480 532 1481
rect 590 1485 596 1486
rect 590 1481 591 1485
rect 595 1481 596 1485
rect 590 1480 596 1481
rect 654 1485 660 1486
rect 654 1481 655 1485
rect 659 1481 660 1485
rect 654 1480 660 1481
rect 718 1485 724 1486
rect 718 1481 719 1485
rect 723 1481 724 1485
rect 718 1480 724 1481
rect 782 1485 788 1486
rect 782 1481 783 1485
rect 787 1481 788 1485
rect 782 1480 788 1481
rect 854 1485 860 1486
rect 854 1481 855 1485
rect 859 1481 860 1485
rect 854 1480 860 1481
rect 528 1475 530 1480
rect 592 1475 594 1480
rect 656 1475 658 1480
rect 720 1475 722 1480
rect 784 1475 786 1480
rect 834 1479 840 1480
rect 834 1475 835 1479
rect 839 1475 840 1479
rect 856 1475 858 1480
rect 511 1474 515 1475
rect 511 1469 515 1470
rect 527 1474 531 1475
rect 527 1469 531 1470
rect 575 1474 579 1475
rect 575 1469 579 1470
rect 591 1474 595 1475
rect 591 1469 595 1470
rect 631 1474 635 1475
rect 631 1469 635 1470
rect 655 1474 659 1475
rect 655 1469 659 1470
rect 687 1474 691 1475
rect 687 1469 691 1470
rect 719 1474 723 1475
rect 719 1469 723 1470
rect 751 1474 755 1475
rect 751 1469 755 1470
rect 783 1474 787 1475
rect 783 1469 787 1470
rect 815 1474 819 1475
rect 834 1474 840 1475
rect 855 1474 859 1475
rect 815 1469 819 1470
rect 482 1467 488 1468
rect 286 1463 292 1464
rect 286 1459 287 1463
rect 291 1459 292 1463
rect 286 1458 292 1459
rect 342 1463 348 1464
rect 342 1459 343 1463
rect 347 1459 348 1463
rect 342 1458 348 1459
rect 398 1463 404 1464
rect 398 1459 399 1463
rect 403 1459 404 1463
rect 454 1463 460 1464
rect 398 1458 404 1459
rect 415 1460 419 1461
rect 454 1459 455 1463
rect 459 1459 460 1463
rect 482 1463 483 1467
rect 487 1463 488 1467
rect 512 1464 514 1469
rect 576 1464 578 1469
rect 632 1464 634 1469
rect 688 1464 690 1469
rect 698 1467 704 1468
rect 482 1462 488 1463
rect 510 1463 516 1464
rect 454 1458 460 1459
rect 510 1459 511 1463
rect 515 1459 516 1463
rect 510 1458 516 1459
rect 574 1463 580 1464
rect 574 1459 575 1463
rect 579 1459 580 1463
rect 574 1458 580 1459
rect 630 1463 636 1464
rect 630 1459 631 1463
rect 635 1459 636 1463
rect 630 1458 636 1459
rect 686 1463 692 1464
rect 686 1459 687 1463
rect 691 1459 692 1463
rect 698 1463 699 1467
rect 703 1463 704 1467
rect 752 1464 754 1469
rect 816 1464 818 1469
rect 698 1462 704 1463
rect 750 1463 756 1464
rect 686 1458 692 1459
rect 415 1455 419 1456
rect 286 1445 292 1446
rect 286 1441 287 1445
rect 291 1441 292 1445
rect 286 1440 292 1441
rect 342 1445 348 1446
rect 342 1441 343 1445
rect 347 1441 348 1445
rect 342 1440 348 1441
rect 398 1445 404 1446
rect 398 1441 399 1445
rect 403 1441 404 1445
rect 398 1440 404 1441
rect 183 1438 187 1440
rect 183 1432 187 1434
rect 231 1438 235 1440
rect 274 1439 280 1440
rect 231 1433 235 1434
rect 255 1438 259 1439
rect 274 1435 275 1439
rect 279 1435 280 1439
rect 274 1434 280 1435
rect 287 1438 291 1440
rect 255 1432 259 1434
rect 287 1433 291 1434
rect 327 1438 331 1439
rect 327 1432 331 1434
rect 343 1438 347 1440
rect 343 1433 347 1434
rect 399 1438 403 1440
rect 399 1432 403 1434
rect 182 1431 188 1432
rect 182 1427 183 1431
rect 187 1427 188 1431
rect 182 1426 188 1427
rect 254 1431 260 1432
rect 254 1427 255 1431
rect 259 1427 260 1431
rect 254 1426 260 1427
rect 326 1431 332 1432
rect 326 1427 327 1431
rect 331 1427 332 1431
rect 326 1426 332 1427
rect 398 1431 404 1432
rect 398 1427 399 1431
rect 403 1427 404 1431
rect 398 1426 404 1427
rect 416 1424 418 1455
rect 642 1451 648 1452
rect 642 1447 643 1451
rect 647 1447 648 1451
rect 642 1446 648 1447
rect 454 1445 460 1446
rect 454 1441 455 1445
rect 459 1441 460 1445
rect 454 1440 460 1441
rect 510 1445 516 1446
rect 510 1441 511 1445
rect 515 1441 516 1445
rect 510 1440 516 1441
rect 574 1445 580 1446
rect 574 1441 575 1445
rect 579 1441 580 1445
rect 574 1440 580 1441
rect 630 1445 636 1446
rect 630 1441 631 1445
rect 635 1441 636 1445
rect 630 1440 636 1441
rect 455 1438 459 1440
rect 455 1433 459 1434
rect 471 1438 475 1439
rect 471 1432 475 1434
rect 511 1438 515 1440
rect 511 1433 515 1434
rect 543 1438 547 1439
rect 543 1432 547 1434
rect 575 1438 579 1440
rect 575 1433 579 1434
rect 615 1438 619 1439
rect 615 1432 619 1434
rect 631 1438 635 1440
rect 631 1433 635 1434
rect 470 1431 476 1432
rect 470 1427 471 1431
rect 475 1427 476 1431
rect 470 1426 476 1427
rect 542 1431 548 1432
rect 542 1427 543 1431
rect 547 1427 548 1431
rect 542 1426 548 1427
rect 614 1431 620 1432
rect 614 1427 615 1431
rect 619 1427 620 1431
rect 614 1426 620 1427
rect 194 1423 200 1424
rect 194 1419 195 1423
rect 199 1419 200 1423
rect 194 1418 200 1419
rect 414 1423 420 1424
rect 414 1419 415 1423
rect 419 1419 420 1423
rect 414 1418 420 1419
rect 482 1423 488 1424
rect 482 1419 483 1423
rect 487 1419 488 1423
rect 482 1418 488 1419
rect 182 1413 188 1414
rect 182 1409 183 1413
rect 187 1409 188 1413
rect 182 1408 188 1409
rect 110 1407 116 1408
rect 112 1403 114 1407
rect 136 1403 138 1408
rect 150 1407 156 1408
rect 150 1403 151 1407
rect 155 1403 156 1407
rect 184 1403 186 1408
rect 111 1402 115 1403
rect 111 1397 115 1398
rect 135 1402 139 1403
rect 150 1402 156 1403
rect 175 1402 179 1403
rect 135 1397 139 1398
rect 175 1397 179 1398
rect 183 1402 187 1403
rect 183 1397 187 1398
rect 112 1393 114 1397
rect 110 1392 116 1393
rect 136 1392 138 1397
rect 176 1392 178 1397
rect 196 1396 198 1418
rect 254 1413 260 1414
rect 254 1409 255 1413
rect 259 1409 260 1413
rect 254 1408 260 1409
rect 326 1413 332 1414
rect 326 1409 327 1413
rect 331 1409 332 1413
rect 326 1408 332 1409
rect 398 1413 404 1414
rect 398 1409 399 1413
rect 403 1409 404 1413
rect 398 1408 404 1409
rect 470 1413 476 1414
rect 470 1409 471 1413
rect 475 1409 476 1413
rect 470 1408 476 1409
rect 256 1403 258 1408
rect 262 1407 268 1408
rect 262 1403 263 1407
rect 267 1403 268 1407
rect 328 1403 330 1408
rect 400 1403 402 1408
rect 472 1403 474 1408
rect 247 1402 251 1403
rect 247 1397 251 1398
rect 255 1402 259 1403
rect 262 1402 268 1403
rect 319 1402 323 1403
rect 255 1397 259 1398
rect 194 1395 200 1396
rect 110 1388 111 1392
rect 115 1388 116 1392
rect 110 1387 116 1388
rect 134 1391 140 1392
rect 134 1387 135 1391
rect 139 1387 140 1391
rect 134 1386 140 1387
rect 174 1391 180 1392
rect 174 1387 175 1391
rect 179 1387 180 1391
rect 194 1391 195 1395
rect 199 1391 200 1395
rect 248 1392 250 1397
rect 194 1390 200 1391
rect 246 1391 252 1392
rect 174 1386 180 1387
rect 246 1387 247 1391
rect 251 1387 252 1391
rect 246 1386 252 1387
rect 264 1380 266 1402
rect 319 1397 323 1398
rect 327 1402 331 1403
rect 327 1397 331 1398
rect 391 1402 395 1403
rect 391 1397 395 1398
rect 399 1402 403 1403
rect 399 1397 403 1398
rect 455 1402 459 1403
rect 455 1397 459 1398
rect 471 1402 475 1403
rect 471 1397 475 1398
rect 320 1392 322 1397
rect 392 1392 394 1397
rect 446 1395 452 1396
rect 318 1391 324 1392
rect 318 1387 319 1391
rect 323 1387 324 1391
rect 318 1386 324 1387
rect 390 1391 396 1392
rect 390 1387 391 1391
rect 395 1387 396 1391
rect 446 1391 447 1395
rect 451 1391 452 1395
rect 456 1392 458 1397
rect 484 1396 486 1418
rect 542 1413 548 1414
rect 542 1409 543 1413
rect 547 1409 548 1413
rect 542 1408 548 1409
rect 614 1413 620 1414
rect 614 1409 615 1413
rect 619 1409 620 1413
rect 644 1412 646 1446
rect 686 1445 692 1446
rect 686 1441 687 1445
rect 691 1441 692 1445
rect 686 1440 692 1441
rect 679 1438 683 1439
rect 679 1432 683 1434
rect 687 1438 691 1440
rect 687 1433 691 1434
rect 678 1431 684 1432
rect 678 1427 679 1431
rect 683 1427 684 1431
rect 678 1426 684 1427
rect 700 1424 702 1462
rect 750 1459 751 1463
rect 755 1459 756 1463
rect 750 1458 756 1459
rect 814 1463 820 1464
rect 814 1459 815 1463
rect 819 1459 820 1463
rect 814 1458 820 1459
rect 836 1452 838 1474
rect 855 1469 859 1470
rect 879 1474 883 1475
rect 879 1469 883 1470
rect 880 1464 882 1469
rect 900 1468 902 1490
rect 934 1485 940 1486
rect 934 1481 935 1485
rect 939 1481 940 1485
rect 934 1480 940 1481
rect 1006 1485 1012 1486
rect 1006 1481 1007 1485
rect 1011 1481 1012 1485
rect 1006 1480 1012 1481
rect 1078 1485 1084 1486
rect 1078 1481 1079 1485
rect 1083 1481 1084 1485
rect 1078 1480 1084 1481
rect 1116 1480 1118 1518
rect 1166 1517 1172 1518
rect 1166 1513 1167 1517
rect 1171 1513 1172 1517
rect 1166 1512 1172 1513
rect 1224 1512 1226 1534
rect 1230 1531 1231 1535
rect 1235 1531 1236 1535
rect 1230 1530 1236 1531
rect 1294 1535 1300 1536
rect 1294 1531 1295 1535
rect 1299 1531 1300 1535
rect 1294 1530 1300 1531
rect 1328 1524 1330 1546
rect 1359 1541 1363 1542
rect 1399 1546 1403 1547
rect 1399 1541 1403 1542
rect 1423 1546 1427 1547
rect 1423 1541 1427 1542
rect 1479 1546 1483 1547
rect 1479 1541 1483 1542
rect 1495 1546 1499 1547
rect 1495 1541 1499 1542
rect 1543 1546 1547 1547
rect 1543 1541 1547 1542
rect 1360 1536 1362 1541
rect 1424 1536 1426 1541
rect 1438 1539 1444 1540
rect 1358 1535 1364 1536
rect 1358 1531 1359 1535
rect 1363 1531 1364 1535
rect 1358 1530 1364 1531
rect 1422 1535 1428 1536
rect 1422 1531 1423 1535
rect 1427 1531 1428 1535
rect 1438 1535 1439 1539
rect 1443 1535 1444 1539
rect 1496 1536 1498 1541
rect 1544 1536 1546 1541
rect 1560 1540 1562 1562
rect 1582 1556 1588 1557
rect 1582 1552 1583 1556
rect 1587 1552 1588 1556
rect 1582 1551 1588 1552
rect 1584 1547 1586 1551
rect 1583 1546 1587 1547
rect 1583 1541 1587 1542
rect 1558 1539 1564 1540
rect 1438 1534 1444 1535
rect 1494 1535 1500 1536
rect 1422 1530 1428 1531
rect 1326 1523 1332 1524
rect 1326 1519 1327 1523
rect 1331 1519 1332 1523
rect 1326 1518 1332 1519
rect 1230 1517 1236 1518
rect 1230 1513 1231 1517
rect 1235 1513 1236 1517
rect 1230 1512 1236 1513
rect 1294 1517 1300 1518
rect 1294 1513 1295 1517
rect 1299 1513 1300 1517
rect 1294 1512 1300 1513
rect 1358 1517 1364 1518
rect 1358 1513 1359 1517
rect 1363 1513 1364 1517
rect 1358 1512 1364 1513
rect 1422 1517 1428 1518
rect 1422 1513 1423 1517
rect 1427 1513 1428 1517
rect 1422 1512 1428 1513
rect 1151 1510 1155 1511
rect 1151 1504 1155 1506
rect 1167 1510 1171 1512
rect 1222 1511 1228 1512
rect 1167 1505 1171 1506
rect 1215 1510 1219 1511
rect 1222 1507 1223 1511
rect 1227 1507 1228 1511
rect 1222 1506 1228 1507
rect 1231 1510 1235 1512
rect 1215 1504 1219 1506
rect 1231 1505 1235 1506
rect 1279 1510 1283 1511
rect 1279 1504 1283 1506
rect 1295 1510 1299 1512
rect 1295 1505 1299 1506
rect 1351 1510 1355 1511
rect 1351 1504 1355 1506
rect 1359 1510 1363 1512
rect 1359 1505 1363 1506
rect 1423 1510 1427 1512
rect 1423 1504 1427 1506
rect 1150 1503 1156 1504
rect 1150 1499 1151 1503
rect 1155 1499 1156 1503
rect 1150 1498 1156 1499
rect 1214 1503 1220 1504
rect 1214 1499 1215 1503
rect 1219 1499 1220 1503
rect 1214 1498 1220 1499
rect 1278 1503 1284 1504
rect 1278 1499 1279 1503
rect 1283 1499 1284 1503
rect 1278 1498 1284 1499
rect 1350 1503 1356 1504
rect 1350 1499 1351 1503
rect 1355 1499 1356 1503
rect 1350 1498 1356 1499
rect 1422 1503 1428 1504
rect 1422 1499 1423 1503
rect 1427 1499 1428 1503
rect 1422 1498 1428 1499
rect 1440 1496 1442 1534
rect 1494 1531 1495 1535
rect 1499 1531 1500 1535
rect 1494 1530 1500 1531
rect 1542 1535 1548 1536
rect 1542 1531 1543 1535
rect 1547 1531 1548 1535
rect 1558 1535 1559 1539
rect 1563 1535 1564 1539
rect 1584 1537 1586 1541
rect 1558 1534 1564 1535
rect 1582 1536 1588 1537
rect 1582 1532 1583 1536
rect 1587 1532 1588 1536
rect 1582 1531 1588 1532
rect 1542 1530 1548 1531
rect 1510 1523 1516 1524
rect 1510 1519 1511 1523
rect 1515 1519 1516 1523
rect 1510 1518 1516 1519
rect 1582 1519 1588 1520
rect 1494 1517 1500 1518
rect 1494 1513 1495 1517
rect 1499 1513 1500 1517
rect 1494 1512 1500 1513
rect 1495 1510 1499 1512
rect 1495 1504 1499 1506
rect 1494 1503 1500 1504
rect 1494 1499 1495 1503
rect 1499 1499 1500 1503
rect 1494 1498 1500 1499
rect 1438 1495 1444 1496
rect 1438 1491 1439 1495
rect 1443 1491 1444 1495
rect 1438 1490 1444 1491
rect 1150 1485 1156 1486
rect 1150 1481 1151 1485
rect 1155 1481 1156 1485
rect 1150 1480 1156 1481
rect 1214 1485 1220 1486
rect 1214 1481 1215 1485
rect 1219 1481 1220 1485
rect 1214 1480 1220 1481
rect 1278 1485 1284 1486
rect 1278 1481 1279 1485
rect 1283 1481 1284 1485
rect 1278 1480 1284 1481
rect 1350 1485 1356 1486
rect 1350 1481 1351 1485
rect 1355 1481 1356 1485
rect 1350 1480 1356 1481
rect 1422 1485 1428 1486
rect 1422 1481 1423 1485
rect 1427 1481 1428 1485
rect 1422 1480 1428 1481
rect 1494 1485 1500 1486
rect 1494 1481 1495 1485
rect 1499 1481 1500 1485
rect 1494 1480 1500 1481
rect 1512 1480 1514 1518
rect 1542 1517 1548 1518
rect 1542 1513 1543 1517
rect 1547 1513 1548 1517
rect 1582 1515 1583 1519
rect 1587 1515 1588 1519
rect 1582 1514 1588 1515
rect 1542 1512 1548 1513
rect 1543 1510 1547 1512
rect 1584 1511 1586 1514
rect 1543 1504 1547 1506
rect 1583 1510 1587 1511
rect 1583 1505 1587 1506
rect 1542 1503 1548 1504
rect 1542 1499 1543 1503
rect 1547 1499 1548 1503
rect 1584 1502 1586 1505
rect 1542 1498 1548 1499
rect 1582 1501 1588 1502
rect 1582 1497 1583 1501
rect 1587 1497 1588 1501
rect 1582 1496 1588 1497
rect 1558 1495 1564 1496
rect 1558 1491 1559 1495
rect 1563 1491 1564 1495
rect 1558 1490 1564 1491
rect 1542 1485 1548 1486
rect 1542 1481 1543 1485
rect 1547 1481 1548 1485
rect 1542 1480 1548 1481
rect 936 1475 938 1480
rect 1008 1475 1010 1480
rect 1080 1475 1082 1480
rect 1114 1479 1120 1480
rect 1114 1475 1115 1479
rect 1119 1475 1120 1479
rect 1152 1475 1154 1480
rect 1216 1475 1218 1480
rect 1280 1475 1282 1480
rect 1352 1475 1354 1480
rect 1424 1475 1426 1480
rect 1496 1475 1498 1480
rect 1510 1479 1516 1480
rect 1510 1475 1511 1479
rect 1515 1475 1516 1479
rect 1544 1475 1546 1480
rect 935 1474 939 1475
rect 935 1469 939 1470
rect 943 1474 947 1475
rect 943 1469 947 1470
rect 1007 1474 1011 1475
rect 1007 1469 1011 1470
rect 1015 1474 1019 1475
rect 1015 1469 1019 1470
rect 1079 1474 1083 1475
rect 1079 1469 1083 1470
rect 1087 1474 1091 1475
rect 1114 1474 1120 1475
rect 1151 1474 1155 1475
rect 1087 1469 1091 1470
rect 1151 1469 1155 1470
rect 1159 1474 1163 1475
rect 1159 1469 1163 1470
rect 1215 1474 1219 1475
rect 1215 1469 1219 1470
rect 1239 1474 1243 1475
rect 1239 1469 1243 1470
rect 1279 1474 1283 1475
rect 1279 1469 1283 1470
rect 1319 1474 1323 1475
rect 1319 1469 1323 1470
rect 1351 1474 1355 1475
rect 1351 1469 1355 1470
rect 1399 1474 1403 1475
rect 1399 1469 1403 1470
rect 1423 1474 1427 1475
rect 1423 1469 1427 1470
rect 1479 1474 1483 1475
rect 1479 1469 1483 1470
rect 1495 1474 1499 1475
rect 1510 1474 1516 1475
rect 1543 1474 1547 1475
rect 1495 1469 1499 1470
rect 1543 1469 1547 1470
rect 898 1467 904 1468
rect 878 1463 884 1464
rect 878 1459 879 1463
rect 883 1459 884 1463
rect 898 1463 899 1467
rect 903 1463 904 1467
rect 944 1464 946 1469
rect 1016 1464 1018 1469
rect 1088 1464 1090 1469
rect 1160 1464 1162 1469
rect 1174 1467 1180 1468
rect 898 1462 904 1463
rect 942 1463 948 1464
rect 878 1458 884 1459
rect 942 1459 943 1463
rect 947 1459 948 1463
rect 942 1458 948 1459
rect 1014 1463 1020 1464
rect 1014 1459 1015 1463
rect 1019 1459 1020 1463
rect 1014 1458 1020 1459
rect 1086 1463 1092 1464
rect 1086 1459 1087 1463
rect 1091 1459 1092 1463
rect 1086 1458 1092 1459
rect 1158 1463 1164 1464
rect 1158 1459 1159 1463
rect 1163 1459 1164 1463
rect 1174 1463 1175 1467
rect 1179 1463 1180 1467
rect 1240 1464 1242 1469
rect 1320 1464 1322 1469
rect 1400 1464 1402 1469
rect 1480 1464 1482 1469
rect 1544 1464 1546 1469
rect 1560 1468 1562 1490
rect 1582 1484 1588 1485
rect 1582 1480 1583 1484
rect 1587 1480 1588 1484
rect 1582 1479 1588 1480
rect 1584 1475 1586 1479
rect 1583 1474 1587 1475
rect 1583 1469 1587 1470
rect 1558 1467 1564 1468
rect 1174 1462 1180 1463
rect 1238 1463 1244 1464
rect 1158 1458 1164 1459
rect 834 1451 840 1452
rect 834 1447 835 1451
rect 839 1447 840 1451
rect 834 1446 840 1447
rect 1102 1451 1108 1452
rect 1102 1447 1103 1451
rect 1107 1447 1108 1451
rect 1102 1446 1108 1447
rect 750 1445 756 1446
rect 750 1441 751 1445
rect 755 1441 756 1445
rect 750 1440 756 1441
rect 814 1445 820 1446
rect 814 1441 815 1445
rect 819 1441 820 1445
rect 814 1440 820 1441
rect 878 1445 884 1446
rect 878 1441 879 1445
rect 883 1441 884 1445
rect 878 1440 884 1441
rect 942 1445 948 1446
rect 942 1441 943 1445
rect 947 1441 948 1445
rect 942 1440 948 1441
rect 1014 1445 1020 1446
rect 1014 1441 1015 1445
rect 1019 1441 1020 1445
rect 1014 1440 1020 1441
rect 1086 1445 1092 1446
rect 1086 1441 1087 1445
rect 1091 1441 1092 1445
rect 1086 1440 1092 1441
rect 743 1438 747 1439
rect 743 1432 747 1434
rect 751 1438 755 1440
rect 751 1433 755 1434
rect 815 1438 819 1440
rect 815 1432 819 1434
rect 879 1438 883 1440
rect 910 1439 916 1440
rect 910 1435 911 1439
rect 915 1435 916 1439
rect 910 1434 916 1435
rect 943 1438 947 1440
rect 879 1432 883 1434
rect 742 1431 748 1432
rect 742 1427 743 1431
rect 747 1427 748 1431
rect 742 1426 748 1427
rect 814 1431 820 1432
rect 814 1427 815 1431
rect 819 1427 820 1431
rect 814 1426 820 1427
rect 878 1431 884 1432
rect 878 1427 879 1431
rect 883 1427 884 1431
rect 878 1426 884 1427
rect 698 1423 704 1424
rect 698 1419 699 1423
rect 703 1419 704 1423
rect 698 1418 704 1419
rect 678 1413 684 1414
rect 614 1408 620 1409
rect 642 1411 648 1412
rect 544 1403 546 1408
rect 616 1403 618 1408
rect 642 1407 643 1411
rect 647 1407 648 1411
rect 678 1409 679 1413
rect 683 1409 684 1413
rect 678 1408 684 1409
rect 742 1413 748 1414
rect 742 1409 743 1413
rect 747 1409 748 1413
rect 742 1408 748 1409
rect 814 1413 820 1414
rect 814 1409 815 1413
rect 819 1409 820 1413
rect 814 1408 820 1409
rect 878 1413 884 1414
rect 878 1409 879 1413
rect 883 1409 884 1413
rect 878 1408 884 1409
rect 642 1406 648 1407
rect 680 1403 682 1408
rect 744 1403 746 1408
rect 816 1403 818 1408
rect 854 1407 860 1408
rect 854 1403 855 1407
rect 859 1403 860 1407
rect 880 1403 882 1408
rect 519 1402 523 1403
rect 519 1397 523 1398
rect 543 1402 547 1403
rect 543 1397 547 1398
rect 583 1402 587 1403
rect 583 1397 587 1398
rect 615 1402 619 1403
rect 615 1397 619 1398
rect 647 1402 651 1403
rect 647 1397 651 1398
rect 679 1402 683 1403
rect 679 1397 683 1398
rect 711 1402 715 1403
rect 711 1397 715 1398
rect 743 1402 747 1403
rect 743 1397 747 1398
rect 775 1402 779 1403
rect 775 1397 779 1398
rect 815 1402 819 1403
rect 815 1397 819 1398
rect 839 1402 843 1403
rect 854 1402 860 1403
rect 879 1402 883 1403
rect 839 1397 843 1398
rect 482 1395 488 1396
rect 446 1390 452 1391
rect 454 1391 460 1392
rect 390 1386 396 1387
rect 150 1379 156 1380
rect 110 1375 116 1376
rect 110 1371 111 1375
rect 115 1371 116 1375
rect 150 1375 151 1379
rect 155 1375 156 1379
rect 150 1374 156 1375
rect 262 1379 268 1380
rect 262 1375 263 1379
rect 267 1375 268 1379
rect 262 1374 268 1375
rect 110 1370 116 1371
rect 134 1373 140 1374
rect 112 1367 114 1370
rect 134 1369 135 1373
rect 139 1369 140 1373
rect 134 1368 140 1369
rect 111 1366 115 1367
rect 111 1361 115 1362
rect 135 1366 139 1368
rect 112 1358 114 1361
rect 135 1360 139 1362
rect 134 1359 140 1360
rect 110 1357 116 1358
rect 110 1353 111 1357
rect 115 1353 116 1357
rect 134 1355 135 1359
rect 139 1355 140 1359
rect 134 1354 140 1355
rect 110 1352 116 1353
rect 134 1341 140 1342
rect 110 1340 116 1341
rect 110 1336 111 1340
rect 115 1336 116 1340
rect 134 1337 135 1341
rect 139 1337 140 1341
rect 134 1336 140 1337
rect 152 1336 154 1374
rect 174 1373 180 1374
rect 174 1369 175 1373
rect 179 1369 180 1373
rect 174 1368 180 1369
rect 246 1373 252 1374
rect 246 1369 247 1373
rect 251 1369 252 1373
rect 246 1368 252 1369
rect 318 1373 324 1374
rect 318 1369 319 1373
rect 323 1369 324 1373
rect 318 1368 324 1369
rect 390 1373 396 1374
rect 390 1369 391 1373
rect 395 1369 396 1373
rect 390 1368 396 1369
rect 448 1368 450 1390
rect 454 1387 455 1391
rect 459 1387 460 1391
rect 482 1391 483 1395
rect 487 1391 488 1395
rect 520 1392 522 1397
rect 584 1392 586 1397
rect 648 1392 650 1397
rect 712 1392 714 1397
rect 776 1392 778 1397
rect 840 1392 842 1397
rect 482 1390 488 1391
rect 518 1391 524 1392
rect 454 1386 460 1387
rect 518 1387 519 1391
rect 523 1387 524 1391
rect 518 1386 524 1387
rect 582 1391 588 1392
rect 582 1387 583 1391
rect 587 1387 588 1391
rect 582 1386 588 1387
rect 646 1391 652 1392
rect 646 1387 647 1391
rect 651 1387 652 1391
rect 646 1386 652 1387
rect 710 1391 716 1392
rect 710 1387 711 1391
rect 715 1387 716 1391
rect 710 1386 716 1387
rect 774 1391 780 1392
rect 774 1387 775 1391
rect 779 1387 780 1391
rect 774 1386 780 1387
rect 838 1391 844 1392
rect 838 1387 839 1391
rect 843 1387 844 1391
rect 838 1386 844 1387
rect 856 1380 858 1402
rect 879 1397 883 1398
rect 895 1402 899 1403
rect 895 1397 899 1398
rect 896 1392 898 1397
rect 912 1396 914 1434
rect 943 1433 947 1434
rect 951 1438 955 1439
rect 951 1432 955 1434
rect 1015 1438 1019 1440
rect 1015 1433 1019 1434
rect 1023 1438 1027 1439
rect 1023 1432 1027 1434
rect 1087 1438 1091 1440
rect 1087 1433 1091 1434
rect 1095 1438 1099 1439
rect 1095 1432 1099 1434
rect 950 1431 956 1432
rect 950 1427 951 1431
rect 955 1427 956 1431
rect 950 1426 956 1427
rect 1022 1431 1028 1432
rect 1022 1427 1023 1431
rect 1027 1427 1028 1431
rect 1022 1426 1028 1427
rect 1094 1431 1100 1432
rect 1094 1427 1095 1431
rect 1099 1427 1100 1431
rect 1094 1426 1100 1427
rect 950 1413 956 1414
rect 950 1409 951 1413
rect 955 1409 956 1413
rect 950 1408 956 1409
rect 1022 1413 1028 1414
rect 1022 1409 1023 1413
rect 1027 1409 1028 1413
rect 1022 1408 1028 1409
rect 1094 1413 1100 1414
rect 1094 1409 1095 1413
rect 1099 1409 1100 1413
rect 1094 1408 1100 1409
rect 952 1403 954 1408
rect 1024 1403 1026 1408
rect 1096 1403 1098 1408
rect 951 1402 955 1403
rect 951 1397 955 1398
rect 999 1402 1003 1403
rect 999 1397 1003 1398
rect 1023 1402 1027 1403
rect 1023 1397 1027 1398
rect 1055 1402 1059 1403
rect 1055 1397 1059 1398
rect 1095 1402 1099 1403
rect 1104 1400 1106 1446
rect 1158 1445 1164 1446
rect 1158 1441 1159 1445
rect 1163 1441 1164 1445
rect 1158 1440 1164 1441
rect 1159 1438 1163 1440
rect 1159 1432 1163 1434
rect 1158 1431 1164 1432
rect 1158 1427 1159 1431
rect 1163 1427 1164 1431
rect 1158 1426 1164 1427
rect 1176 1424 1178 1462
rect 1238 1459 1239 1463
rect 1243 1459 1244 1463
rect 1238 1458 1244 1459
rect 1318 1463 1324 1464
rect 1318 1459 1319 1463
rect 1323 1459 1324 1463
rect 1318 1458 1324 1459
rect 1398 1463 1404 1464
rect 1398 1459 1399 1463
rect 1403 1459 1404 1463
rect 1398 1458 1404 1459
rect 1478 1463 1484 1464
rect 1478 1459 1479 1463
rect 1483 1459 1484 1463
rect 1478 1458 1484 1459
rect 1542 1463 1548 1464
rect 1542 1459 1543 1463
rect 1547 1459 1548 1463
rect 1558 1463 1559 1467
rect 1563 1463 1564 1467
rect 1584 1465 1586 1469
rect 1558 1462 1564 1463
rect 1582 1464 1588 1465
rect 1582 1460 1583 1464
rect 1587 1460 1588 1464
rect 1582 1459 1588 1460
rect 1542 1458 1548 1459
rect 1526 1451 1532 1452
rect 1526 1447 1527 1451
rect 1531 1447 1532 1451
rect 1526 1446 1532 1447
rect 1582 1447 1588 1448
rect 1238 1445 1244 1446
rect 1238 1441 1239 1445
rect 1243 1441 1244 1445
rect 1238 1440 1244 1441
rect 1318 1445 1324 1446
rect 1318 1441 1319 1445
rect 1323 1441 1324 1445
rect 1318 1440 1324 1441
rect 1398 1445 1404 1446
rect 1398 1441 1399 1445
rect 1403 1441 1404 1445
rect 1398 1440 1404 1441
rect 1478 1445 1484 1446
rect 1478 1441 1479 1445
rect 1483 1441 1484 1445
rect 1478 1440 1484 1441
rect 1223 1438 1227 1439
rect 1223 1432 1227 1434
rect 1239 1438 1243 1440
rect 1239 1433 1243 1434
rect 1287 1438 1291 1439
rect 1287 1432 1291 1434
rect 1319 1438 1323 1440
rect 1362 1439 1368 1440
rect 1319 1433 1323 1434
rect 1343 1438 1347 1439
rect 1362 1435 1363 1439
rect 1367 1435 1368 1439
rect 1362 1434 1368 1435
rect 1399 1438 1403 1440
rect 1343 1432 1347 1434
rect 1222 1431 1228 1432
rect 1222 1427 1223 1431
rect 1227 1427 1228 1431
rect 1222 1426 1228 1427
rect 1286 1431 1292 1432
rect 1286 1427 1287 1431
rect 1291 1427 1292 1431
rect 1286 1426 1292 1427
rect 1342 1431 1348 1432
rect 1342 1427 1343 1431
rect 1347 1427 1348 1431
rect 1342 1426 1348 1427
rect 1174 1423 1180 1424
rect 1174 1419 1175 1423
rect 1179 1419 1180 1423
rect 1174 1418 1180 1419
rect 1158 1413 1164 1414
rect 1158 1409 1159 1413
rect 1163 1409 1164 1413
rect 1158 1408 1164 1409
rect 1222 1413 1228 1414
rect 1222 1409 1223 1413
rect 1227 1409 1228 1413
rect 1222 1408 1228 1409
rect 1286 1413 1292 1414
rect 1286 1409 1287 1413
rect 1291 1409 1292 1413
rect 1286 1408 1292 1409
rect 1342 1413 1348 1414
rect 1342 1409 1343 1413
rect 1347 1409 1348 1413
rect 1342 1408 1348 1409
rect 1364 1408 1366 1434
rect 1399 1432 1403 1434
rect 1455 1438 1459 1439
rect 1455 1432 1459 1434
rect 1479 1438 1483 1440
rect 1479 1433 1483 1434
rect 1511 1438 1515 1439
rect 1511 1432 1515 1434
rect 1398 1431 1404 1432
rect 1398 1427 1399 1431
rect 1403 1427 1404 1431
rect 1398 1426 1404 1427
rect 1454 1431 1460 1432
rect 1454 1427 1455 1431
rect 1459 1427 1460 1431
rect 1454 1426 1460 1427
rect 1510 1431 1516 1432
rect 1510 1427 1511 1431
rect 1515 1427 1516 1431
rect 1510 1426 1516 1427
rect 1494 1423 1500 1424
rect 1494 1419 1495 1423
rect 1499 1419 1500 1423
rect 1494 1418 1500 1419
rect 1398 1413 1404 1414
rect 1398 1409 1399 1413
rect 1403 1409 1404 1413
rect 1398 1408 1404 1409
rect 1454 1413 1460 1414
rect 1454 1409 1455 1413
rect 1459 1409 1460 1413
rect 1454 1408 1460 1409
rect 1160 1403 1162 1408
rect 1224 1403 1226 1408
rect 1288 1403 1290 1408
rect 1306 1407 1312 1408
rect 1306 1403 1307 1407
rect 1311 1403 1312 1407
rect 1344 1403 1346 1408
rect 1362 1407 1368 1408
rect 1362 1403 1363 1407
rect 1367 1403 1368 1407
rect 1400 1403 1402 1408
rect 1456 1403 1458 1408
rect 1111 1402 1115 1403
rect 1095 1397 1099 1398
rect 1102 1399 1108 1400
rect 910 1395 916 1396
rect 894 1391 900 1392
rect 894 1387 895 1391
rect 899 1387 900 1391
rect 910 1391 911 1395
rect 915 1391 916 1395
rect 952 1392 954 1397
rect 1000 1392 1002 1397
rect 1056 1392 1058 1397
rect 1102 1395 1103 1399
rect 1107 1395 1108 1399
rect 1111 1397 1115 1398
rect 1159 1402 1163 1403
rect 1159 1397 1163 1398
rect 1175 1402 1179 1403
rect 1175 1397 1179 1398
rect 1223 1402 1227 1403
rect 1223 1397 1227 1398
rect 1239 1402 1243 1403
rect 1239 1397 1243 1398
rect 1287 1402 1291 1403
rect 1287 1397 1291 1398
rect 1295 1402 1299 1403
rect 1306 1402 1312 1403
rect 1343 1402 1347 1403
rect 1295 1397 1299 1398
rect 1102 1394 1108 1395
rect 1112 1392 1114 1397
rect 1176 1392 1178 1397
rect 1186 1395 1192 1396
rect 910 1390 916 1391
rect 950 1391 956 1392
rect 894 1386 900 1387
rect 950 1387 951 1391
rect 955 1387 956 1391
rect 950 1386 956 1387
rect 998 1391 1004 1392
rect 998 1387 999 1391
rect 1003 1387 1004 1391
rect 998 1386 1004 1387
rect 1054 1391 1060 1392
rect 1054 1387 1055 1391
rect 1059 1387 1060 1391
rect 1054 1386 1060 1387
rect 1110 1391 1116 1392
rect 1110 1387 1111 1391
rect 1115 1387 1116 1391
rect 1110 1386 1116 1387
rect 1174 1391 1180 1392
rect 1174 1387 1175 1391
rect 1179 1387 1180 1391
rect 1186 1391 1187 1395
rect 1191 1391 1192 1395
rect 1240 1392 1242 1397
rect 1296 1392 1298 1397
rect 1186 1390 1192 1391
rect 1238 1391 1244 1392
rect 1174 1386 1180 1387
rect 854 1379 860 1380
rect 854 1375 855 1379
rect 859 1375 860 1379
rect 854 1374 860 1375
rect 1126 1379 1132 1380
rect 1126 1375 1127 1379
rect 1131 1375 1132 1379
rect 1126 1374 1132 1375
rect 454 1373 460 1374
rect 454 1369 455 1373
rect 459 1369 460 1373
rect 454 1368 460 1369
rect 518 1373 524 1374
rect 518 1369 519 1373
rect 523 1369 524 1373
rect 518 1368 524 1369
rect 582 1373 588 1374
rect 582 1369 583 1373
rect 587 1369 588 1373
rect 582 1368 588 1369
rect 646 1373 652 1374
rect 646 1369 647 1373
rect 651 1369 652 1373
rect 646 1368 652 1369
rect 710 1373 716 1374
rect 710 1369 711 1373
rect 715 1369 716 1373
rect 710 1368 716 1369
rect 774 1373 780 1374
rect 774 1369 775 1373
rect 779 1369 780 1373
rect 774 1368 780 1369
rect 838 1373 844 1374
rect 838 1369 839 1373
rect 843 1369 844 1373
rect 838 1368 844 1369
rect 894 1373 900 1374
rect 894 1369 895 1373
rect 899 1369 900 1373
rect 894 1368 900 1369
rect 950 1373 956 1374
rect 950 1369 951 1373
rect 955 1369 956 1373
rect 950 1368 956 1369
rect 998 1373 1004 1374
rect 998 1369 999 1373
rect 1003 1369 1004 1373
rect 998 1368 1004 1369
rect 1054 1373 1060 1374
rect 1054 1369 1055 1373
rect 1059 1369 1060 1373
rect 1054 1368 1060 1369
rect 1110 1373 1116 1374
rect 1110 1369 1111 1373
rect 1115 1369 1116 1373
rect 1110 1368 1116 1369
rect 167 1366 171 1367
rect 167 1360 171 1362
rect 175 1366 179 1368
rect 175 1361 179 1362
rect 215 1366 219 1367
rect 215 1360 219 1362
rect 247 1366 251 1368
rect 247 1361 251 1362
rect 303 1366 307 1367
rect 303 1360 307 1362
rect 319 1366 323 1368
rect 319 1361 323 1362
rect 391 1366 395 1368
rect 446 1367 452 1368
rect 391 1361 395 1362
rect 415 1366 419 1367
rect 446 1363 447 1367
rect 451 1363 452 1367
rect 446 1362 452 1363
rect 455 1366 459 1368
rect 415 1360 419 1362
rect 455 1361 459 1362
rect 519 1366 523 1368
rect 519 1361 523 1362
rect 527 1366 531 1367
rect 527 1360 531 1362
rect 583 1366 587 1368
rect 583 1361 587 1362
rect 639 1366 643 1367
rect 639 1360 643 1362
rect 647 1366 651 1368
rect 647 1361 651 1362
rect 711 1366 715 1368
rect 711 1361 715 1362
rect 751 1366 755 1367
rect 751 1360 755 1362
rect 775 1366 779 1368
rect 775 1361 779 1362
rect 839 1366 843 1368
rect 839 1361 843 1362
rect 863 1366 867 1367
rect 863 1360 867 1362
rect 895 1366 899 1368
rect 895 1361 899 1362
rect 951 1366 955 1368
rect 951 1361 955 1362
rect 967 1366 971 1367
rect 967 1360 971 1362
rect 999 1366 1003 1368
rect 999 1361 1003 1362
rect 1055 1366 1059 1368
rect 1055 1361 1059 1362
rect 1063 1366 1067 1367
rect 1063 1360 1067 1362
rect 1111 1366 1115 1368
rect 1111 1361 1115 1362
rect 1128 1360 1130 1374
rect 1174 1373 1180 1374
rect 1174 1369 1175 1373
rect 1179 1369 1180 1373
rect 1174 1368 1180 1369
rect 1151 1366 1155 1367
rect 1151 1360 1155 1362
rect 1175 1366 1179 1368
rect 1175 1361 1179 1362
rect 166 1359 172 1360
rect 166 1355 167 1359
rect 171 1355 172 1359
rect 166 1354 172 1355
rect 214 1359 220 1360
rect 214 1355 215 1359
rect 219 1355 220 1359
rect 214 1354 220 1355
rect 302 1359 308 1360
rect 302 1355 303 1359
rect 307 1355 308 1359
rect 302 1354 308 1355
rect 414 1359 420 1360
rect 414 1355 415 1359
rect 419 1355 420 1359
rect 414 1354 420 1355
rect 526 1359 532 1360
rect 526 1355 527 1359
rect 531 1355 532 1359
rect 526 1354 532 1355
rect 638 1359 644 1360
rect 638 1355 639 1359
rect 643 1355 644 1359
rect 638 1354 644 1355
rect 750 1359 756 1360
rect 750 1355 751 1359
rect 755 1355 756 1359
rect 750 1354 756 1355
rect 862 1359 868 1360
rect 862 1355 863 1359
rect 867 1355 868 1359
rect 862 1354 868 1355
rect 966 1359 972 1360
rect 966 1355 967 1359
rect 971 1355 972 1359
rect 966 1354 972 1355
rect 1062 1359 1068 1360
rect 1062 1355 1063 1359
rect 1067 1355 1068 1359
rect 1062 1354 1068 1355
rect 1126 1359 1132 1360
rect 1126 1355 1127 1359
rect 1131 1355 1132 1359
rect 1126 1354 1132 1355
rect 1150 1359 1156 1360
rect 1150 1355 1151 1359
rect 1155 1355 1156 1359
rect 1150 1354 1156 1355
rect 1188 1352 1190 1390
rect 1238 1387 1239 1391
rect 1243 1387 1244 1391
rect 1238 1386 1244 1387
rect 1294 1391 1300 1392
rect 1294 1387 1295 1391
rect 1299 1387 1300 1391
rect 1294 1386 1300 1387
rect 1308 1380 1310 1402
rect 1343 1397 1347 1398
rect 1351 1402 1355 1403
rect 1362 1402 1368 1403
rect 1399 1402 1403 1403
rect 1351 1397 1355 1398
rect 1399 1397 1403 1398
rect 1415 1402 1419 1403
rect 1415 1397 1419 1398
rect 1455 1402 1459 1403
rect 1455 1397 1459 1398
rect 1479 1402 1483 1403
rect 1479 1397 1483 1398
rect 1352 1392 1354 1397
rect 1406 1395 1412 1396
rect 1350 1391 1356 1392
rect 1350 1387 1351 1391
rect 1355 1387 1356 1391
rect 1406 1391 1407 1395
rect 1411 1391 1412 1395
rect 1416 1392 1418 1397
rect 1480 1392 1482 1397
rect 1496 1396 1498 1418
rect 1510 1413 1516 1414
rect 1510 1409 1511 1413
rect 1515 1409 1516 1413
rect 1510 1408 1516 1409
rect 1528 1408 1530 1446
rect 1542 1445 1548 1446
rect 1542 1441 1543 1445
rect 1547 1441 1548 1445
rect 1582 1443 1583 1447
rect 1587 1443 1588 1447
rect 1582 1442 1588 1443
rect 1542 1440 1548 1441
rect 1543 1438 1547 1440
rect 1584 1439 1586 1442
rect 1543 1432 1547 1434
rect 1583 1438 1587 1439
rect 1583 1433 1587 1434
rect 1542 1431 1548 1432
rect 1542 1427 1543 1431
rect 1547 1427 1548 1431
rect 1584 1430 1586 1433
rect 1542 1426 1548 1427
rect 1582 1429 1588 1430
rect 1582 1425 1583 1429
rect 1587 1425 1588 1429
rect 1582 1424 1588 1425
rect 1542 1413 1548 1414
rect 1542 1409 1543 1413
rect 1547 1409 1548 1413
rect 1542 1408 1548 1409
rect 1582 1412 1588 1413
rect 1582 1408 1583 1412
rect 1587 1408 1588 1412
rect 1512 1403 1514 1408
rect 1526 1407 1532 1408
rect 1526 1403 1527 1407
rect 1531 1403 1532 1407
rect 1544 1403 1546 1408
rect 1582 1407 1588 1408
rect 1584 1403 1586 1407
rect 1511 1402 1515 1403
rect 1526 1402 1532 1403
rect 1543 1402 1547 1403
rect 1511 1397 1515 1398
rect 1543 1397 1547 1398
rect 1583 1402 1587 1403
rect 1583 1397 1587 1398
rect 1494 1395 1500 1396
rect 1406 1390 1412 1391
rect 1414 1391 1420 1392
rect 1350 1386 1356 1387
rect 1306 1379 1312 1380
rect 1306 1375 1307 1379
rect 1311 1375 1312 1379
rect 1306 1374 1312 1375
rect 1238 1373 1244 1374
rect 1238 1369 1239 1373
rect 1243 1369 1244 1373
rect 1238 1368 1244 1369
rect 1294 1373 1300 1374
rect 1294 1369 1295 1373
rect 1299 1369 1300 1373
rect 1294 1368 1300 1369
rect 1350 1373 1356 1374
rect 1350 1369 1351 1373
rect 1355 1369 1356 1373
rect 1350 1368 1356 1369
rect 1408 1368 1410 1390
rect 1414 1387 1415 1391
rect 1419 1387 1420 1391
rect 1414 1386 1420 1387
rect 1478 1391 1484 1392
rect 1478 1387 1479 1391
rect 1483 1387 1484 1391
rect 1494 1391 1495 1395
rect 1499 1391 1500 1395
rect 1544 1392 1546 1397
rect 1584 1393 1586 1397
rect 1582 1392 1588 1393
rect 1494 1390 1500 1391
rect 1542 1391 1548 1392
rect 1478 1386 1484 1387
rect 1542 1387 1543 1391
rect 1547 1387 1548 1391
rect 1582 1388 1583 1392
rect 1587 1388 1588 1392
rect 1582 1387 1588 1388
rect 1542 1386 1548 1387
rect 1462 1379 1468 1380
rect 1462 1375 1463 1379
rect 1467 1375 1468 1379
rect 1462 1374 1468 1375
rect 1582 1375 1588 1376
rect 1414 1373 1420 1374
rect 1414 1369 1415 1373
rect 1419 1369 1420 1373
rect 1414 1368 1420 1369
rect 1231 1366 1235 1367
rect 1231 1360 1235 1362
rect 1239 1366 1243 1368
rect 1239 1361 1243 1362
rect 1295 1366 1299 1368
rect 1295 1361 1299 1362
rect 1311 1366 1315 1367
rect 1311 1360 1315 1362
rect 1351 1366 1355 1368
rect 1406 1367 1412 1368
rect 1351 1361 1355 1362
rect 1383 1366 1387 1367
rect 1406 1363 1407 1367
rect 1411 1363 1412 1367
rect 1406 1362 1412 1363
rect 1415 1366 1419 1368
rect 1383 1360 1387 1362
rect 1415 1361 1419 1362
rect 1455 1366 1459 1367
rect 1455 1360 1459 1362
rect 1230 1359 1236 1360
rect 1230 1355 1231 1359
rect 1235 1355 1236 1359
rect 1230 1354 1236 1355
rect 1310 1359 1316 1360
rect 1310 1355 1311 1359
rect 1315 1355 1316 1359
rect 1310 1354 1316 1355
rect 1382 1359 1388 1360
rect 1382 1355 1383 1359
rect 1387 1355 1388 1359
rect 1382 1354 1388 1355
rect 1454 1359 1460 1360
rect 1454 1355 1455 1359
rect 1459 1355 1460 1359
rect 1454 1354 1460 1355
rect 202 1351 208 1352
rect 202 1347 203 1351
rect 207 1347 208 1351
rect 202 1346 208 1347
rect 902 1351 908 1352
rect 902 1347 903 1351
rect 907 1347 908 1351
rect 902 1346 908 1347
rect 910 1351 916 1352
rect 910 1347 911 1351
rect 915 1347 916 1351
rect 910 1346 916 1347
rect 1186 1351 1192 1352
rect 1186 1347 1187 1351
rect 1191 1347 1192 1351
rect 1186 1346 1192 1347
rect 1438 1351 1444 1352
rect 1438 1347 1439 1351
rect 1443 1347 1444 1351
rect 1438 1346 1444 1347
rect 1446 1351 1452 1352
rect 1446 1347 1447 1351
rect 1451 1347 1452 1351
rect 1446 1346 1452 1347
rect 166 1341 172 1342
rect 166 1337 167 1341
rect 171 1337 172 1341
rect 166 1336 172 1337
rect 110 1335 116 1336
rect 112 1331 114 1335
rect 136 1331 138 1336
rect 150 1335 156 1336
rect 150 1331 151 1335
rect 155 1331 156 1335
rect 168 1331 170 1336
rect 111 1330 115 1331
rect 111 1325 115 1326
rect 135 1330 139 1331
rect 150 1330 156 1331
rect 167 1330 171 1331
rect 135 1325 139 1326
rect 167 1325 171 1326
rect 183 1330 187 1331
rect 183 1325 187 1326
rect 112 1321 114 1325
rect 110 1320 116 1321
rect 136 1320 138 1325
rect 184 1320 186 1325
rect 204 1324 206 1346
rect 214 1341 220 1342
rect 214 1337 215 1341
rect 219 1337 220 1341
rect 214 1336 220 1337
rect 302 1341 308 1342
rect 302 1337 303 1341
rect 307 1337 308 1341
rect 302 1336 308 1337
rect 414 1341 420 1342
rect 414 1337 415 1341
rect 419 1337 420 1341
rect 414 1336 420 1337
rect 526 1341 532 1342
rect 526 1337 527 1341
rect 531 1337 532 1341
rect 526 1336 532 1337
rect 638 1341 644 1342
rect 638 1337 639 1341
rect 643 1337 644 1341
rect 638 1336 644 1337
rect 750 1341 756 1342
rect 750 1337 751 1341
rect 755 1337 756 1341
rect 750 1336 756 1337
rect 862 1341 868 1342
rect 862 1337 863 1341
rect 867 1337 868 1341
rect 862 1336 868 1337
rect 216 1331 218 1336
rect 266 1335 272 1336
rect 266 1331 267 1335
rect 271 1331 272 1335
rect 304 1331 306 1336
rect 416 1331 418 1336
rect 528 1331 530 1336
rect 640 1331 642 1336
rect 752 1331 754 1336
rect 864 1331 866 1336
rect 215 1330 219 1331
rect 215 1325 219 1326
rect 247 1330 251 1331
rect 266 1330 272 1331
rect 303 1330 307 1331
rect 247 1325 251 1326
rect 202 1323 208 1324
rect 110 1316 111 1320
rect 115 1316 116 1320
rect 110 1315 116 1316
rect 134 1319 140 1320
rect 134 1315 135 1319
rect 139 1315 140 1319
rect 134 1314 140 1315
rect 182 1319 188 1320
rect 182 1315 183 1319
rect 187 1315 188 1319
rect 202 1319 203 1323
rect 207 1319 208 1323
rect 248 1320 250 1325
rect 202 1318 208 1319
rect 246 1319 252 1320
rect 182 1314 188 1315
rect 246 1315 247 1319
rect 251 1315 252 1319
rect 246 1314 252 1315
rect 268 1308 270 1330
rect 303 1325 307 1326
rect 311 1330 315 1331
rect 311 1325 315 1326
rect 375 1330 379 1331
rect 375 1325 379 1326
rect 415 1330 419 1331
rect 415 1325 419 1326
rect 439 1330 443 1331
rect 439 1325 443 1326
rect 495 1330 499 1331
rect 495 1325 499 1326
rect 527 1330 531 1331
rect 527 1325 531 1326
rect 543 1330 547 1331
rect 543 1325 547 1326
rect 591 1330 595 1331
rect 591 1325 595 1326
rect 639 1330 643 1331
rect 639 1325 643 1326
rect 687 1330 691 1331
rect 687 1325 691 1326
rect 743 1330 747 1331
rect 743 1325 747 1326
rect 751 1330 755 1331
rect 751 1325 755 1326
rect 791 1330 795 1331
rect 791 1325 795 1326
rect 839 1330 843 1331
rect 839 1325 843 1326
rect 863 1330 867 1331
rect 863 1325 867 1326
rect 887 1330 891 1331
rect 887 1325 891 1326
rect 312 1320 314 1325
rect 376 1320 378 1325
rect 406 1323 412 1324
rect 310 1319 316 1320
rect 310 1315 311 1319
rect 315 1315 316 1319
rect 310 1314 316 1315
rect 374 1319 380 1320
rect 374 1315 375 1319
rect 379 1315 380 1319
rect 406 1319 407 1323
rect 411 1319 412 1323
rect 440 1320 442 1325
rect 478 1323 484 1324
rect 406 1318 412 1319
rect 438 1319 444 1320
rect 374 1314 380 1315
rect 150 1307 156 1308
rect 110 1303 116 1304
rect 110 1299 111 1303
rect 115 1299 116 1303
rect 150 1303 151 1307
rect 155 1303 156 1307
rect 150 1302 156 1303
rect 266 1307 272 1308
rect 266 1303 267 1307
rect 271 1303 272 1307
rect 266 1302 272 1303
rect 110 1298 116 1299
rect 134 1301 140 1302
rect 112 1295 114 1298
rect 134 1297 135 1301
rect 139 1297 140 1301
rect 134 1296 140 1297
rect 111 1294 115 1295
rect 111 1289 115 1290
rect 135 1294 139 1296
rect 112 1286 114 1289
rect 135 1288 139 1290
rect 134 1287 140 1288
rect 110 1285 116 1286
rect 110 1281 111 1285
rect 115 1281 116 1285
rect 134 1283 135 1287
rect 139 1283 140 1287
rect 134 1282 140 1283
rect 110 1280 116 1281
rect 134 1269 140 1270
rect 110 1268 116 1269
rect 110 1264 111 1268
rect 115 1264 116 1268
rect 134 1265 135 1269
rect 139 1265 140 1269
rect 134 1264 140 1265
rect 152 1264 154 1302
rect 182 1301 188 1302
rect 182 1297 183 1301
rect 187 1297 188 1301
rect 182 1296 188 1297
rect 246 1301 252 1302
rect 246 1297 247 1301
rect 251 1297 252 1301
rect 246 1296 252 1297
rect 310 1301 316 1302
rect 310 1297 311 1301
rect 315 1297 316 1301
rect 310 1296 316 1297
rect 374 1301 380 1302
rect 374 1297 375 1301
rect 379 1297 380 1301
rect 374 1296 380 1297
rect 183 1294 187 1296
rect 183 1289 187 1290
rect 191 1294 195 1295
rect 191 1288 195 1290
rect 247 1294 251 1296
rect 247 1289 251 1290
rect 255 1294 259 1295
rect 255 1288 259 1290
rect 311 1294 315 1296
rect 311 1289 315 1290
rect 327 1294 331 1295
rect 327 1288 331 1290
rect 375 1294 379 1296
rect 375 1289 379 1290
rect 391 1294 395 1295
rect 391 1288 395 1290
rect 190 1287 196 1288
rect 190 1283 191 1287
rect 195 1283 196 1287
rect 190 1282 196 1283
rect 254 1287 260 1288
rect 254 1283 255 1287
rect 259 1283 260 1287
rect 254 1282 260 1283
rect 326 1287 332 1288
rect 326 1283 327 1287
rect 331 1283 332 1287
rect 326 1282 332 1283
rect 390 1287 396 1288
rect 390 1283 391 1287
rect 395 1283 396 1287
rect 390 1282 396 1283
rect 408 1280 410 1318
rect 438 1315 439 1319
rect 443 1315 444 1319
rect 478 1319 479 1323
rect 483 1319 484 1323
rect 496 1320 498 1325
rect 544 1320 546 1325
rect 592 1320 594 1325
rect 640 1320 642 1325
rect 688 1320 690 1325
rect 744 1320 746 1325
rect 792 1320 794 1325
rect 840 1320 842 1325
rect 888 1320 890 1325
rect 904 1324 906 1346
rect 912 1332 914 1346
rect 966 1341 972 1342
rect 966 1337 967 1341
rect 971 1337 972 1341
rect 966 1336 972 1337
rect 1062 1341 1068 1342
rect 1062 1337 1063 1341
rect 1067 1337 1068 1341
rect 1062 1336 1068 1337
rect 1150 1341 1156 1342
rect 1150 1337 1151 1341
rect 1155 1337 1156 1341
rect 1150 1336 1156 1337
rect 1230 1341 1236 1342
rect 1230 1337 1231 1341
rect 1235 1337 1236 1341
rect 1230 1336 1236 1337
rect 1310 1341 1316 1342
rect 1382 1341 1388 1342
rect 1310 1337 1311 1341
rect 1315 1337 1316 1341
rect 1355 1340 1359 1341
rect 1310 1336 1316 1337
rect 910 1331 916 1332
rect 968 1331 970 1336
rect 1064 1331 1066 1336
rect 1152 1331 1154 1336
rect 1232 1331 1234 1336
rect 1238 1335 1244 1336
rect 1238 1331 1239 1335
rect 1243 1331 1244 1335
rect 1312 1331 1314 1336
rect 1354 1335 1355 1340
rect 1359 1335 1360 1340
rect 1382 1337 1383 1341
rect 1387 1337 1388 1341
rect 1382 1336 1388 1337
rect 1354 1334 1360 1335
rect 1384 1331 1386 1336
rect 910 1327 911 1331
rect 915 1327 916 1331
rect 910 1326 916 1327
rect 935 1330 939 1331
rect 935 1325 939 1326
rect 967 1330 971 1331
rect 967 1325 971 1326
rect 991 1330 995 1331
rect 991 1325 995 1326
rect 1047 1330 1051 1331
rect 1063 1330 1067 1331
rect 1047 1325 1051 1326
rect 1054 1327 1060 1328
rect 902 1323 908 1324
rect 478 1318 484 1319
rect 494 1319 500 1320
rect 438 1314 444 1315
rect 438 1301 444 1302
rect 438 1297 439 1301
rect 443 1297 444 1301
rect 438 1296 444 1297
rect 439 1294 443 1296
rect 439 1289 443 1290
rect 463 1294 467 1295
rect 463 1288 467 1290
rect 462 1287 468 1288
rect 462 1283 463 1287
rect 467 1283 468 1287
rect 462 1282 468 1283
rect 480 1280 482 1318
rect 494 1315 495 1319
rect 499 1315 500 1319
rect 494 1314 500 1315
rect 542 1319 548 1320
rect 542 1315 543 1319
rect 547 1315 548 1319
rect 542 1314 548 1315
rect 590 1319 596 1320
rect 590 1315 591 1319
rect 595 1315 596 1319
rect 590 1314 596 1315
rect 638 1319 644 1320
rect 638 1315 639 1319
rect 643 1315 644 1319
rect 638 1314 644 1315
rect 686 1319 692 1320
rect 686 1315 687 1319
rect 691 1315 692 1319
rect 686 1314 692 1315
rect 742 1319 748 1320
rect 742 1315 743 1319
rect 747 1315 748 1319
rect 742 1314 748 1315
rect 790 1319 796 1320
rect 790 1315 791 1319
rect 795 1315 796 1319
rect 790 1314 796 1315
rect 838 1319 844 1320
rect 838 1315 839 1319
rect 843 1315 844 1319
rect 838 1314 844 1315
rect 886 1319 892 1320
rect 886 1315 887 1319
rect 891 1315 892 1319
rect 902 1319 903 1323
rect 907 1319 908 1323
rect 936 1320 938 1325
rect 992 1320 994 1325
rect 1048 1320 1050 1325
rect 1054 1323 1055 1327
rect 1059 1323 1060 1327
rect 1063 1325 1067 1326
rect 1103 1330 1107 1331
rect 1103 1325 1107 1326
rect 1151 1330 1155 1331
rect 1151 1325 1155 1326
rect 1159 1330 1163 1331
rect 1159 1325 1163 1326
rect 1215 1330 1219 1331
rect 1215 1325 1219 1326
rect 1231 1330 1235 1331
rect 1238 1330 1244 1331
rect 1271 1330 1275 1331
rect 1231 1325 1235 1326
rect 1054 1322 1060 1323
rect 902 1318 908 1319
rect 934 1319 940 1320
rect 886 1314 892 1315
rect 934 1315 935 1319
rect 939 1315 940 1319
rect 934 1314 940 1315
rect 990 1319 996 1320
rect 990 1315 991 1319
rect 995 1315 996 1319
rect 990 1314 996 1315
rect 1046 1319 1052 1320
rect 1046 1315 1047 1319
rect 1051 1315 1052 1319
rect 1046 1314 1052 1315
rect 854 1307 860 1308
rect 854 1303 855 1307
rect 859 1303 860 1307
rect 854 1302 860 1303
rect 1006 1307 1012 1308
rect 1006 1303 1007 1307
rect 1011 1303 1012 1307
rect 1006 1302 1012 1303
rect 494 1301 500 1302
rect 494 1297 495 1301
rect 499 1297 500 1301
rect 494 1296 500 1297
rect 542 1301 548 1302
rect 542 1297 543 1301
rect 547 1297 548 1301
rect 542 1296 548 1297
rect 590 1301 596 1302
rect 590 1297 591 1301
rect 595 1297 596 1301
rect 590 1296 596 1297
rect 638 1301 644 1302
rect 638 1297 639 1301
rect 643 1297 644 1301
rect 638 1296 644 1297
rect 686 1301 692 1302
rect 686 1297 687 1301
rect 691 1297 692 1301
rect 686 1296 692 1297
rect 742 1301 748 1302
rect 742 1297 743 1301
rect 747 1297 748 1301
rect 742 1296 748 1297
rect 790 1301 796 1302
rect 790 1297 791 1301
rect 795 1297 796 1301
rect 790 1296 796 1297
rect 838 1301 844 1302
rect 838 1297 839 1301
rect 843 1297 844 1301
rect 856 1299 858 1302
rect 838 1296 844 1297
rect 848 1297 858 1299
rect 886 1301 892 1302
rect 886 1297 887 1301
rect 891 1297 892 1301
rect 495 1294 499 1296
rect 495 1289 499 1290
rect 535 1294 539 1295
rect 535 1288 539 1290
rect 543 1294 547 1296
rect 543 1289 547 1290
rect 591 1294 595 1296
rect 591 1289 595 1290
rect 599 1294 603 1295
rect 599 1288 603 1290
rect 639 1294 643 1296
rect 639 1289 643 1290
rect 663 1294 667 1295
rect 663 1288 667 1290
rect 687 1294 691 1296
rect 687 1289 691 1290
rect 727 1294 731 1295
rect 727 1288 731 1290
rect 743 1294 747 1296
rect 743 1289 747 1290
rect 791 1294 795 1296
rect 791 1288 795 1290
rect 839 1294 843 1296
rect 839 1289 843 1290
rect 534 1287 540 1288
rect 534 1283 535 1287
rect 539 1283 540 1287
rect 534 1282 540 1283
rect 598 1287 604 1288
rect 598 1283 599 1287
rect 603 1283 604 1287
rect 598 1282 604 1283
rect 662 1287 668 1288
rect 662 1283 663 1287
rect 667 1283 668 1287
rect 662 1282 668 1283
rect 726 1287 732 1288
rect 726 1283 727 1287
rect 731 1283 732 1287
rect 726 1282 732 1283
rect 790 1287 796 1288
rect 790 1283 791 1287
rect 795 1283 796 1287
rect 790 1282 796 1283
rect 246 1279 252 1280
rect 246 1275 247 1279
rect 251 1275 252 1279
rect 246 1274 252 1275
rect 406 1279 412 1280
rect 406 1275 407 1279
rect 411 1275 412 1279
rect 406 1274 412 1275
rect 478 1279 484 1280
rect 478 1275 479 1279
rect 483 1275 484 1279
rect 478 1274 484 1275
rect 190 1269 196 1270
rect 190 1265 191 1269
rect 195 1265 196 1269
rect 190 1264 196 1265
rect 110 1263 116 1264
rect 112 1259 114 1263
rect 136 1259 138 1264
rect 150 1263 156 1264
rect 150 1259 151 1263
rect 155 1259 156 1263
rect 192 1259 194 1264
rect 111 1258 115 1259
rect 111 1253 115 1254
rect 135 1258 139 1259
rect 150 1258 156 1259
rect 175 1258 179 1259
rect 135 1253 139 1254
rect 175 1253 179 1254
rect 191 1258 195 1259
rect 191 1253 195 1254
rect 231 1258 235 1259
rect 231 1253 235 1254
rect 112 1249 114 1253
rect 110 1248 116 1249
rect 136 1248 138 1253
rect 176 1248 178 1253
rect 232 1248 234 1253
rect 248 1252 250 1274
rect 814 1271 820 1272
rect 254 1269 260 1270
rect 254 1265 255 1269
rect 259 1265 260 1269
rect 254 1264 260 1265
rect 326 1269 332 1270
rect 326 1265 327 1269
rect 331 1265 332 1269
rect 326 1264 332 1265
rect 390 1269 396 1270
rect 390 1265 391 1269
rect 395 1265 396 1269
rect 390 1264 396 1265
rect 462 1269 468 1270
rect 462 1265 463 1269
rect 467 1265 468 1269
rect 462 1264 468 1265
rect 534 1269 540 1270
rect 534 1265 535 1269
rect 539 1265 540 1269
rect 534 1264 540 1265
rect 598 1269 604 1270
rect 598 1265 599 1269
rect 603 1265 604 1269
rect 598 1264 604 1265
rect 662 1269 668 1270
rect 662 1265 663 1269
rect 667 1265 668 1269
rect 662 1264 668 1265
rect 726 1269 732 1270
rect 726 1265 727 1269
rect 731 1265 732 1269
rect 726 1264 732 1265
rect 790 1269 796 1270
rect 790 1265 791 1269
rect 795 1265 796 1269
rect 814 1267 815 1271
rect 819 1267 820 1271
rect 814 1266 820 1267
rect 790 1264 796 1265
rect 256 1259 258 1264
rect 302 1263 308 1264
rect 302 1259 303 1263
rect 307 1259 308 1263
rect 328 1259 330 1264
rect 392 1259 394 1264
rect 464 1259 466 1264
rect 536 1259 538 1264
rect 600 1259 602 1264
rect 618 1263 624 1264
rect 618 1259 619 1263
rect 623 1259 624 1263
rect 664 1259 666 1264
rect 728 1259 730 1264
rect 792 1259 794 1264
rect 255 1258 259 1259
rect 255 1253 259 1254
rect 287 1258 291 1259
rect 302 1258 308 1259
rect 327 1258 331 1259
rect 287 1253 291 1254
rect 246 1251 252 1252
rect 110 1244 111 1248
rect 115 1244 116 1248
rect 110 1243 116 1244
rect 134 1247 140 1248
rect 134 1243 135 1247
rect 139 1243 140 1247
rect 134 1242 140 1243
rect 174 1247 180 1248
rect 174 1243 175 1247
rect 179 1243 180 1247
rect 174 1242 180 1243
rect 230 1247 236 1248
rect 230 1243 231 1247
rect 235 1243 236 1247
rect 246 1247 247 1251
rect 251 1247 252 1251
rect 288 1248 290 1253
rect 246 1246 252 1247
rect 286 1247 292 1248
rect 230 1242 236 1243
rect 286 1243 287 1247
rect 291 1243 292 1247
rect 286 1242 292 1243
rect 304 1236 306 1258
rect 351 1258 355 1259
rect 327 1253 331 1254
rect 334 1255 340 1256
rect 334 1251 335 1255
rect 339 1251 340 1255
rect 351 1253 355 1254
rect 391 1258 395 1259
rect 391 1253 395 1254
rect 415 1258 419 1259
rect 415 1253 419 1254
rect 463 1258 467 1259
rect 463 1253 467 1254
rect 479 1258 483 1259
rect 479 1253 483 1254
rect 535 1258 539 1259
rect 535 1253 539 1254
rect 543 1258 547 1259
rect 599 1258 603 1259
rect 543 1253 547 1254
rect 570 1255 576 1256
rect 334 1250 340 1251
rect 154 1235 160 1236
rect 110 1231 116 1232
rect 110 1227 111 1231
rect 115 1227 116 1231
rect 154 1231 155 1235
rect 159 1231 160 1235
rect 154 1230 160 1231
rect 302 1235 308 1236
rect 302 1231 303 1235
rect 307 1231 308 1235
rect 302 1230 308 1231
rect 110 1226 116 1227
rect 134 1229 140 1230
rect 112 1223 114 1226
rect 134 1225 135 1229
rect 139 1225 140 1229
rect 134 1224 140 1225
rect 111 1222 115 1223
rect 111 1217 115 1218
rect 135 1222 139 1224
rect 135 1217 139 1218
rect 143 1222 147 1223
rect 112 1214 114 1217
rect 143 1216 147 1218
rect 142 1215 148 1216
rect 110 1213 116 1214
rect 110 1209 111 1213
rect 115 1209 116 1213
rect 142 1211 143 1215
rect 147 1211 148 1215
rect 142 1210 148 1211
rect 110 1208 116 1209
rect 142 1197 148 1198
rect 110 1196 116 1197
rect 110 1192 111 1196
rect 115 1192 116 1196
rect 142 1193 143 1197
rect 147 1193 148 1197
rect 142 1192 148 1193
rect 156 1192 158 1230
rect 174 1229 180 1230
rect 174 1225 175 1229
rect 179 1225 180 1229
rect 174 1224 180 1225
rect 230 1229 236 1230
rect 230 1225 231 1229
rect 235 1225 236 1229
rect 230 1224 236 1225
rect 286 1229 292 1230
rect 286 1225 287 1229
rect 291 1225 292 1229
rect 286 1224 292 1225
rect 175 1222 179 1224
rect 175 1216 179 1218
rect 215 1222 219 1223
rect 215 1216 219 1218
rect 231 1222 235 1224
rect 231 1217 235 1218
rect 263 1222 267 1223
rect 263 1216 267 1218
rect 287 1222 291 1224
rect 294 1223 300 1224
rect 294 1219 295 1223
rect 299 1219 300 1223
rect 294 1218 300 1219
rect 311 1222 315 1223
rect 287 1217 291 1218
rect 174 1215 180 1216
rect 174 1211 175 1215
rect 179 1211 180 1215
rect 174 1210 180 1211
rect 214 1215 220 1216
rect 214 1211 215 1215
rect 219 1211 220 1215
rect 214 1210 220 1211
rect 262 1215 268 1216
rect 262 1211 263 1215
rect 267 1211 268 1215
rect 262 1210 268 1211
rect 230 1207 236 1208
rect 230 1203 231 1207
rect 235 1203 236 1207
rect 230 1202 236 1203
rect 174 1197 180 1198
rect 174 1193 175 1197
rect 179 1193 180 1197
rect 174 1192 180 1193
rect 214 1197 220 1198
rect 214 1193 215 1197
rect 219 1193 220 1197
rect 214 1192 220 1193
rect 110 1191 116 1192
rect 112 1187 114 1191
rect 144 1187 146 1192
rect 154 1191 160 1192
rect 154 1187 155 1191
rect 159 1187 160 1191
rect 176 1187 178 1192
rect 216 1187 218 1192
rect 111 1186 115 1187
rect 111 1181 115 1182
rect 143 1186 147 1187
rect 154 1186 160 1187
rect 175 1186 179 1187
rect 143 1181 147 1182
rect 175 1181 179 1182
rect 215 1186 219 1187
rect 215 1181 219 1182
rect 112 1177 114 1181
rect 110 1176 116 1177
rect 144 1176 146 1181
rect 176 1176 178 1181
rect 216 1176 218 1181
rect 232 1180 234 1202
rect 262 1197 268 1198
rect 262 1193 263 1197
rect 267 1193 268 1197
rect 262 1192 268 1193
rect 296 1192 298 1218
rect 311 1216 315 1218
rect 310 1215 316 1216
rect 310 1211 311 1215
rect 315 1211 316 1215
rect 310 1210 316 1211
rect 327 1207 333 1208
rect 327 1203 328 1207
rect 332 1206 333 1207
rect 336 1206 338 1250
rect 352 1248 354 1253
rect 416 1248 418 1253
rect 430 1251 436 1252
rect 350 1247 356 1248
rect 350 1243 351 1247
rect 355 1243 356 1247
rect 350 1242 356 1243
rect 414 1247 420 1248
rect 414 1243 415 1247
rect 419 1243 420 1247
rect 430 1247 431 1251
rect 435 1247 436 1251
rect 480 1248 482 1253
rect 544 1248 546 1253
rect 570 1251 571 1255
rect 575 1251 576 1255
rect 599 1253 603 1254
rect 607 1258 611 1259
rect 618 1258 624 1259
rect 663 1258 667 1259
rect 607 1253 611 1254
rect 570 1250 576 1251
rect 430 1246 436 1247
rect 478 1247 484 1248
rect 414 1242 420 1243
rect 350 1229 356 1230
rect 350 1225 351 1229
rect 355 1225 356 1229
rect 350 1224 356 1225
rect 414 1229 420 1230
rect 414 1225 415 1229
rect 419 1225 420 1229
rect 414 1224 420 1225
rect 351 1222 355 1224
rect 351 1217 355 1218
rect 359 1222 363 1223
rect 359 1216 363 1218
rect 415 1222 419 1224
rect 415 1216 419 1218
rect 358 1215 364 1216
rect 358 1211 359 1215
rect 363 1211 364 1215
rect 358 1210 364 1211
rect 414 1215 420 1216
rect 414 1211 415 1215
rect 419 1211 420 1215
rect 414 1210 420 1211
rect 432 1208 434 1246
rect 478 1243 479 1247
rect 483 1243 484 1247
rect 478 1242 484 1243
rect 542 1247 548 1248
rect 542 1243 543 1247
rect 547 1243 548 1247
rect 542 1242 548 1243
rect 572 1236 574 1250
rect 608 1248 610 1253
rect 606 1247 612 1248
rect 606 1243 607 1247
rect 611 1243 612 1247
rect 606 1242 612 1243
rect 620 1236 622 1258
rect 663 1253 667 1254
rect 671 1258 675 1259
rect 671 1253 675 1254
rect 727 1258 731 1259
rect 727 1253 731 1254
rect 735 1258 739 1259
rect 735 1253 739 1254
rect 791 1258 795 1259
rect 791 1253 795 1254
rect 799 1258 803 1259
rect 799 1253 803 1254
rect 672 1248 674 1253
rect 736 1248 738 1253
rect 800 1248 802 1253
rect 816 1252 818 1266
rect 848 1264 850 1297
rect 886 1296 892 1297
rect 934 1301 940 1302
rect 934 1297 935 1301
rect 939 1297 940 1301
rect 934 1296 940 1297
rect 990 1301 996 1302
rect 990 1297 991 1301
rect 995 1297 996 1301
rect 990 1296 996 1297
rect 855 1294 859 1295
rect 855 1288 859 1290
rect 887 1294 891 1296
rect 887 1289 891 1290
rect 927 1294 931 1295
rect 927 1288 931 1290
rect 935 1294 939 1296
rect 935 1289 939 1290
rect 991 1294 995 1296
rect 991 1289 995 1290
rect 999 1294 1003 1295
rect 999 1288 1003 1290
rect 854 1287 860 1288
rect 854 1283 855 1287
rect 859 1283 860 1287
rect 854 1282 860 1283
rect 926 1287 932 1288
rect 926 1283 927 1287
rect 931 1283 932 1287
rect 926 1282 932 1283
rect 998 1287 1004 1288
rect 998 1283 999 1287
rect 1003 1283 1004 1287
rect 998 1282 1004 1283
rect 874 1279 880 1280
rect 874 1275 875 1279
rect 879 1275 880 1279
rect 874 1274 880 1275
rect 854 1269 860 1270
rect 854 1265 855 1269
rect 859 1265 860 1269
rect 854 1264 860 1265
rect 846 1263 852 1264
rect 846 1259 847 1263
rect 851 1259 852 1263
rect 856 1259 858 1264
rect 846 1258 852 1259
rect 855 1258 859 1259
rect 855 1253 859 1254
rect 863 1258 867 1259
rect 863 1253 867 1254
rect 814 1251 820 1252
rect 670 1247 676 1248
rect 670 1243 671 1247
rect 675 1243 676 1247
rect 670 1242 676 1243
rect 734 1247 740 1248
rect 734 1243 735 1247
rect 739 1243 740 1247
rect 734 1242 740 1243
rect 798 1247 804 1248
rect 798 1243 799 1247
rect 803 1243 804 1247
rect 814 1247 815 1251
rect 819 1247 820 1251
rect 864 1248 866 1253
rect 876 1252 878 1274
rect 926 1269 932 1270
rect 926 1265 927 1269
rect 931 1265 932 1269
rect 926 1264 932 1265
rect 998 1269 1004 1270
rect 998 1265 999 1269
rect 1003 1265 1004 1269
rect 998 1264 1004 1265
rect 1008 1264 1010 1302
rect 1046 1301 1052 1302
rect 1046 1297 1047 1301
rect 1051 1297 1052 1301
rect 1046 1296 1052 1297
rect 1018 1295 1024 1296
rect 1018 1291 1019 1295
rect 1023 1291 1024 1295
rect 1018 1290 1024 1291
rect 1047 1294 1051 1296
rect 1020 1264 1022 1290
rect 1047 1289 1051 1290
rect 1056 1280 1058 1322
rect 1104 1320 1106 1325
rect 1160 1320 1162 1325
rect 1216 1320 1218 1325
rect 1102 1319 1108 1320
rect 1102 1315 1103 1319
rect 1107 1315 1108 1319
rect 1102 1314 1108 1315
rect 1158 1319 1164 1320
rect 1158 1315 1159 1319
rect 1163 1315 1164 1319
rect 1158 1314 1164 1315
rect 1214 1319 1220 1320
rect 1214 1315 1215 1319
rect 1219 1315 1220 1319
rect 1214 1314 1220 1315
rect 1231 1307 1237 1308
rect 1231 1303 1232 1307
rect 1236 1306 1237 1307
rect 1240 1306 1242 1330
rect 1271 1325 1275 1326
rect 1311 1330 1315 1331
rect 1311 1325 1315 1326
rect 1327 1330 1331 1331
rect 1327 1325 1331 1326
rect 1375 1330 1379 1331
rect 1375 1325 1379 1326
rect 1383 1330 1387 1331
rect 1383 1325 1387 1326
rect 1423 1330 1427 1331
rect 1423 1325 1427 1326
rect 1272 1320 1274 1325
rect 1328 1320 1330 1325
rect 1376 1320 1378 1325
rect 1414 1323 1420 1324
rect 1270 1319 1276 1320
rect 1270 1315 1271 1319
rect 1275 1315 1276 1319
rect 1270 1314 1276 1315
rect 1326 1319 1332 1320
rect 1326 1315 1327 1319
rect 1331 1315 1332 1319
rect 1326 1314 1332 1315
rect 1374 1319 1380 1320
rect 1374 1315 1375 1319
rect 1379 1315 1380 1319
rect 1414 1319 1415 1323
rect 1419 1319 1420 1323
rect 1424 1320 1426 1325
rect 1440 1324 1442 1346
rect 1448 1341 1450 1346
rect 1454 1341 1460 1342
rect 1447 1340 1451 1341
rect 1454 1337 1455 1341
rect 1459 1337 1460 1341
rect 1454 1336 1460 1337
rect 1464 1336 1466 1374
rect 1478 1373 1484 1374
rect 1478 1369 1479 1373
rect 1483 1369 1484 1373
rect 1478 1368 1484 1369
rect 1542 1373 1548 1374
rect 1542 1369 1543 1373
rect 1547 1369 1548 1373
rect 1582 1371 1583 1375
rect 1587 1371 1588 1375
rect 1582 1370 1588 1371
rect 1542 1368 1548 1369
rect 1479 1366 1483 1368
rect 1479 1361 1483 1362
rect 1535 1366 1539 1367
rect 1535 1360 1539 1362
rect 1543 1366 1547 1368
rect 1584 1367 1586 1370
rect 1543 1361 1547 1362
rect 1583 1366 1587 1367
rect 1583 1361 1587 1362
rect 1534 1359 1540 1360
rect 1534 1355 1535 1359
rect 1539 1355 1540 1359
rect 1584 1358 1586 1361
rect 1534 1354 1540 1355
rect 1582 1357 1588 1358
rect 1582 1353 1583 1357
rect 1587 1353 1588 1357
rect 1582 1352 1588 1353
rect 1534 1341 1540 1342
rect 1534 1337 1535 1341
rect 1539 1337 1540 1341
rect 1534 1336 1540 1337
rect 1582 1340 1588 1341
rect 1582 1336 1583 1340
rect 1587 1336 1588 1340
rect 1447 1335 1451 1336
rect 1456 1331 1458 1336
rect 1462 1335 1468 1336
rect 1462 1331 1463 1335
rect 1467 1331 1468 1335
rect 1536 1331 1538 1336
rect 1582 1335 1588 1336
rect 1584 1331 1586 1335
rect 1455 1330 1459 1331
rect 1462 1330 1468 1331
rect 1471 1330 1475 1331
rect 1455 1325 1459 1326
rect 1471 1325 1475 1326
rect 1527 1330 1531 1331
rect 1527 1325 1531 1326
rect 1535 1330 1539 1331
rect 1535 1325 1539 1326
rect 1583 1330 1587 1331
rect 1583 1325 1587 1326
rect 1438 1323 1444 1324
rect 1414 1318 1420 1319
rect 1422 1319 1428 1320
rect 1374 1314 1380 1315
rect 1236 1304 1242 1306
rect 1358 1307 1364 1308
rect 1236 1303 1237 1304
rect 1231 1302 1237 1303
rect 1358 1303 1359 1307
rect 1363 1303 1364 1307
rect 1358 1302 1364 1303
rect 1102 1301 1108 1302
rect 1102 1297 1103 1301
rect 1107 1297 1108 1301
rect 1102 1296 1108 1297
rect 1158 1301 1164 1302
rect 1158 1297 1159 1301
rect 1163 1297 1164 1301
rect 1158 1296 1164 1297
rect 1214 1301 1220 1302
rect 1214 1297 1215 1301
rect 1219 1297 1220 1301
rect 1214 1296 1220 1297
rect 1270 1301 1276 1302
rect 1270 1297 1271 1301
rect 1275 1297 1276 1301
rect 1270 1296 1276 1297
rect 1326 1301 1332 1302
rect 1326 1297 1327 1301
rect 1331 1297 1332 1301
rect 1326 1296 1332 1297
rect 1063 1294 1067 1295
rect 1063 1288 1067 1290
rect 1103 1294 1107 1296
rect 1103 1289 1107 1290
rect 1127 1294 1131 1295
rect 1127 1288 1131 1290
rect 1159 1294 1163 1296
rect 1159 1289 1163 1290
rect 1191 1294 1195 1295
rect 1191 1288 1195 1290
rect 1215 1294 1219 1296
rect 1222 1295 1228 1296
rect 1222 1291 1223 1295
rect 1227 1291 1228 1295
rect 1222 1290 1228 1291
rect 1247 1294 1251 1295
rect 1215 1289 1219 1290
rect 1062 1287 1068 1288
rect 1062 1283 1063 1287
rect 1067 1283 1068 1287
rect 1062 1282 1068 1283
rect 1126 1287 1132 1288
rect 1126 1283 1127 1287
rect 1131 1283 1132 1287
rect 1126 1282 1132 1283
rect 1190 1287 1196 1288
rect 1190 1283 1191 1287
rect 1195 1283 1196 1287
rect 1190 1282 1196 1283
rect 1054 1279 1060 1280
rect 1054 1275 1055 1279
rect 1059 1275 1060 1279
rect 1054 1274 1060 1275
rect 1062 1269 1068 1270
rect 1062 1265 1063 1269
rect 1067 1265 1068 1269
rect 1062 1264 1068 1265
rect 1126 1269 1132 1270
rect 1126 1265 1127 1269
rect 1131 1265 1132 1269
rect 1126 1264 1132 1265
rect 1190 1269 1196 1270
rect 1190 1265 1191 1269
rect 1195 1265 1196 1269
rect 1190 1264 1196 1265
rect 1224 1264 1226 1290
rect 1247 1288 1251 1290
rect 1271 1294 1275 1296
rect 1271 1289 1275 1290
rect 1303 1294 1307 1295
rect 1303 1288 1307 1290
rect 1327 1294 1331 1296
rect 1327 1289 1331 1290
rect 1246 1287 1252 1288
rect 1246 1283 1247 1287
rect 1251 1283 1252 1287
rect 1246 1282 1252 1283
rect 1302 1287 1308 1288
rect 1302 1283 1303 1287
rect 1307 1283 1308 1287
rect 1302 1282 1308 1283
rect 1246 1269 1252 1270
rect 1246 1265 1247 1269
rect 1251 1265 1252 1269
rect 1246 1264 1252 1265
rect 1302 1269 1308 1270
rect 1302 1265 1303 1269
rect 1307 1265 1308 1269
rect 1302 1264 1308 1265
rect 1360 1264 1362 1302
rect 1374 1301 1380 1302
rect 1374 1297 1375 1301
rect 1379 1297 1380 1301
rect 1374 1296 1380 1297
rect 1416 1296 1418 1318
rect 1422 1315 1423 1319
rect 1427 1315 1428 1319
rect 1438 1319 1439 1323
rect 1443 1319 1444 1323
rect 1472 1320 1474 1325
rect 1528 1320 1530 1325
rect 1584 1321 1586 1325
rect 1582 1320 1588 1321
rect 1438 1318 1444 1319
rect 1470 1319 1476 1320
rect 1422 1314 1428 1315
rect 1470 1315 1471 1319
rect 1475 1315 1476 1319
rect 1470 1314 1476 1315
rect 1526 1319 1532 1320
rect 1526 1315 1527 1319
rect 1531 1315 1532 1319
rect 1582 1316 1583 1320
rect 1587 1316 1588 1320
rect 1582 1315 1588 1316
rect 1526 1314 1532 1315
rect 1582 1303 1588 1304
rect 1422 1301 1428 1302
rect 1422 1297 1423 1301
rect 1427 1297 1428 1301
rect 1422 1296 1428 1297
rect 1470 1301 1476 1302
rect 1470 1297 1471 1301
rect 1475 1297 1476 1301
rect 1470 1296 1476 1297
rect 1526 1301 1532 1302
rect 1526 1297 1527 1301
rect 1531 1297 1532 1301
rect 1582 1299 1583 1303
rect 1587 1299 1588 1303
rect 1582 1298 1588 1299
rect 1526 1296 1532 1297
rect 1367 1294 1371 1295
rect 1367 1288 1371 1290
rect 1375 1294 1379 1296
rect 1414 1295 1420 1296
rect 1414 1291 1415 1295
rect 1419 1291 1420 1295
rect 1414 1290 1420 1291
rect 1423 1294 1427 1296
rect 1375 1289 1379 1290
rect 1423 1289 1427 1290
rect 1431 1294 1435 1295
rect 1431 1288 1435 1290
rect 1471 1294 1475 1296
rect 1471 1289 1475 1290
rect 1527 1294 1531 1296
rect 1584 1295 1586 1298
rect 1527 1289 1531 1290
rect 1583 1294 1587 1295
rect 1583 1289 1587 1290
rect 1366 1287 1372 1288
rect 1366 1283 1367 1287
rect 1371 1283 1372 1287
rect 1366 1282 1372 1283
rect 1430 1287 1436 1288
rect 1430 1283 1431 1287
rect 1435 1283 1436 1287
rect 1584 1286 1586 1289
rect 1430 1282 1436 1283
rect 1582 1285 1588 1286
rect 1582 1281 1583 1285
rect 1587 1281 1588 1285
rect 1582 1280 1588 1281
rect 1366 1269 1372 1270
rect 1366 1265 1367 1269
rect 1371 1265 1372 1269
rect 1366 1264 1372 1265
rect 1430 1269 1436 1270
rect 1430 1265 1431 1269
rect 1435 1265 1436 1269
rect 1430 1264 1436 1265
rect 1582 1268 1588 1269
rect 1582 1264 1583 1268
rect 1587 1264 1588 1268
rect 928 1259 930 1264
rect 1000 1259 1002 1264
rect 1006 1263 1012 1264
rect 1006 1259 1007 1263
rect 1011 1259 1012 1263
rect 927 1258 931 1259
rect 927 1253 931 1254
rect 991 1258 995 1259
rect 991 1253 995 1254
rect 999 1258 1003 1259
rect 1006 1258 1012 1259
rect 1018 1263 1024 1264
rect 1018 1259 1019 1263
rect 1023 1259 1024 1263
rect 1064 1259 1066 1264
rect 1074 1263 1080 1264
rect 1074 1259 1075 1263
rect 1079 1259 1080 1263
rect 1128 1259 1130 1264
rect 1192 1259 1194 1264
rect 1222 1263 1228 1264
rect 1222 1259 1223 1263
rect 1227 1259 1228 1263
rect 1248 1259 1250 1264
rect 1304 1259 1306 1264
rect 1358 1263 1364 1264
rect 1358 1259 1359 1263
rect 1363 1259 1364 1263
rect 1368 1259 1370 1264
rect 1432 1259 1434 1264
rect 1582 1263 1588 1264
rect 1584 1259 1586 1263
rect 1018 1258 1024 1259
rect 1055 1258 1059 1259
rect 999 1253 1003 1254
rect 1055 1253 1059 1254
rect 1063 1258 1067 1259
rect 1074 1258 1080 1259
rect 1119 1258 1123 1259
rect 1063 1253 1067 1254
rect 874 1251 880 1252
rect 814 1246 820 1247
rect 862 1247 868 1248
rect 798 1242 804 1243
rect 862 1243 863 1247
rect 867 1243 868 1247
rect 874 1247 875 1251
rect 879 1247 880 1251
rect 928 1248 930 1253
rect 992 1248 994 1253
rect 1056 1248 1058 1253
rect 874 1246 880 1247
rect 926 1247 932 1248
rect 862 1242 868 1243
rect 926 1243 927 1247
rect 931 1243 932 1247
rect 926 1242 932 1243
rect 990 1247 996 1248
rect 990 1243 991 1247
rect 995 1243 996 1247
rect 990 1242 996 1243
rect 1054 1247 1060 1248
rect 1054 1243 1055 1247
rect 1059 1243 1060 1247
rect 1054 1242 1060 1243
rect 1076 1236 1078 1258
rect 1119 1253 1123 1254
rect 1127 1258 1131 1259
rect 1127 1253 1131 1254
rect 1183 1258 1187 1259
rect 1183 1253 1187 1254
rect 1191 1258 1195 1259
rect 1222 1258 1228 1259
rect 1247 1258 1251 1259
rect 1191 1253 1195 1254
rect 1247 1253 1251 1254
rect 1303 1258 1307 1259
rect 1303 1253 1307 1254
rect 1311 1258 1315 1259
rect 1358 1258 1364 1259
rect 1367 1258 1371 1259
rect 1311 1253 1315 1254
rect 1367 1253 1371 1254
rect 1375 1258 1379 1259
rect 1375 1253 1379 1254
rect 1431 1258 1435 1259
rect 1431 1253 1435 1254
rect 1439 1258 1443 1259
rect 1439 1253 1443 1254
rect 1503 1258 1507 1259
rect 1503 1253 1507 1254
rect 1543 1258 1547 1259
rect 1543 1253 1547 1254
rect 1583 1258 1587 1259
rect 1583 1253 1587 1254
rect 1120 1248 1122 1253
rect 1174 1251 1180 1252
rect 1118 1247 1124 1248
rect 1118 1243 1119 1247
rect 1123 1243 1124 1247
rect 1174 1247 1175 1251
rect 1179 1247 1180 1251
rect 1184 1248 1186 1253
rect 1248 1248 1250 1253
rect 1312 1248 1314 1253
rect 1376 1248 1378 1253
rect 1440 1248 1442 1253
rect 1486 1251 1492 1252
rect 1174 1246 1180 1247
rect 1182 1247 1188 1248
rect 1118 1242 1124 1243
rect 570 1235 576 1236
rect 570 1231 571 1235
rect 575 1231 576 1235
rect 570 1230 576 1231
rect 618 1235 624 1236
rect 618 1231 619 1235
rect 623 1231 624 1235
rect 618 1230 624 1231
rect 702 1235 708 1236
rect 702 1231 703 1235
rect 707 1231 708 1235
rect 702 1230 708 1231
rect 946 1235 952 1236
rect 946 1231 947 1235
rect 951 1231 952 1235
rect 946 1230 952 1231
rect 1074 1235 1080 1236
rect 1074 1231 1075 1235
rect 1079 1231 1080 1235
rect 1074 1230 1080 1231
rect 478 1229 484 1230
rect 478 1225 479 1229
rect 483 1225 484 1229
rect 478 1224 484 1225
rect 542 1229 548 1230
rect 542 1225 543 1229
rect 547 1225 548 1229
rect 542 1224 548 1225
rect 606 1229 612 1230
rect 606 1225 607 1229
rect 611 1225 612 1229
rect 606 1224 612 1225
rect 670 1229 676 1230
rect 670 1225 671 1229
rect 675 1225 676 1229
rect 670 1224 676 1225
rect 471 1222 475 1223
rect 471 1216 475 1218
rect 479 1222 483 1224
rect 479 1217 483 1218
rect 527 1222 531 1223
rect 527 1216 531 1218
rect 543 1222 547 1224
rect 543 1217 547 1218
rect 583 1222 587 1223
rect 583 1216 587 1218
rect 607 1222 611 1224
rect 607 1217 611 1218
rect 639 1222 643 1223
rect 639 1216 643 1218
rect 671 1222 675 1224
rect 671 1217 675 1218
rect 687 1222 691 1223
rect 687 1216 691 1218
rect 470 1215 476 1216
rect 470 1211 471 1215
rect 475 1211 476 1215
rect 470 1210 476 1211
rect 526 1215 532 1216
rect 526 1211 527 1215
rect 531 1211 532 1215
rect 526 1210 532 1211
rect 582 1215 588 1216
rect 582 1211 583 1215
rect 587 1211 588 1215
rect 582 1210 588 1211
rect 638 1215 644 1216
rect 638 1211 639 1215
rect 643 1211 644 1215
rect 638 1210 644 1211
rect 686 1215 692 1216
rect 686 1211 687 1215
rect 691 1211 692 1215
rect 686 1210 692 1211
rect 332 1204 338 1206
rect 430 1207 436 1208
rect 332 1203 333 1204
rect 327 1202 333 1203
rect 430 1203 431 1207
rect 435 1203 436 1207
rect 430 1202 436 1203
rect 310 1197 316 1198
rect 310 1193 311 1197
rect 315 1193 316 1197
rect 310 1192 316 1193
rect 358 1197 364 1198
rect 358 1193 359 1197
rect 363 1193 364 1197
rect 358 1192 364 1193
rect 414 1197 420 1198
rect 414 1193 415 1197
rect 419 1193 420 1197
rect 414 1192 420 1193
rect 470 1197 476 1198
rect 470 1193 471 1197
rect 475 1193 476 1197
rect 470 1192 476 1193
rect 526 1197 532 1198
rect 526 1193 527 1197
rect 531 1193 532 1197
rect 526 1192 532 1193
rect 582 1197 588 1198
rect 582 1193 583 1197
rect 587 1193 588 1197
rect 582 1192 588 1193
rect 638 1197 644 1198
rect 638 1193 639 1197
rect 643 1193 644 1197
rect 638 1192 644 1193
rect 686 1197 692 1198
rect 686 1193 687 1197
rect 691 1193 692 1197
rect 686 1192 692 1193
rect 704 1192 706 1230
rect 734 1229 740 1230
rect 734 1225 735 1229
rect 739 1225 740 1229
rect 734 1224 740 1225
rect 798 1229 804 1230
rect 798 1225 799 1229
rect 803 1225 804 1229
rect 798 1224 804 1225
rect 862 1229 868 1230
rect 862 1225 863 1229
rect 867 1225 868 1229
rect 862 1224 868 1225
rect 926 1229 932 1230
rect 926 1225 927 1229
rect 931 1225 932 1229
rect 926 1224 932 1225
rect 735 1222 739 1224
rect 735 1216 739 1218
rect 783 1222 787 1223
rect 783 1216 787 1218
rect 799 1222 803 1224
rect 799 1217 803 1218
rect 831 1222 835 1223
rect 831 1216 835 1218
rect 863 1222 867 1224
rect 863 1217 867 1218
rect 879 1222 883 1223
rect 879 1216 883 1218
rect 927 1222 931 1224
rect 927 1217 931 1218
rect 935 1222 939 1223
rect 935 1216 939 1218
rect 734 1215 740 1216
rect 734 1211 735 1215
rect 739 1211 740 1215
rect 734 1210 740 1211
rect 782 1215 788 1216
rect 782 1211 783 1215
rect 787 1211 788 1215
rect 782 1210 788 1211
rect 830 1215 836 1216
rect 830 1211 831 1215
rect 835 1211 836 1215
rect 830 1210 836 1211
rect 878 1215 884 1216
rect 878 1211 879 1215
rect 883 1211 884 1215
rect 878 1210 884 1211
rect 934 1215 940 1216
rect 934 1211 935 1215
rect 939 1211 940 1215
rect 934 1210 940 1211
rect 734 1197 740 1198
rect 734 1193 735 1197
rect 739 1193 740 1197
rect 734 1192 740 1193
rect 782 1197 788 1198
rect 782 1193 783 1197
rect 787 1193 788 1197
rect 782 1192 788 1193
rect 830 1197 836 1198
rect 830 1193 831 1197
rect 835 1193 836 1197
rect 830 1192 836 1193
rect 878 1197 884 1198
rect 878 1193 879 1197
rect 883 1193 884 1197
rect 878 1192 884 1193
rect 934 1197 940 1198
rect 934 1193 935 1197
rect 939 1193 940 1197
rect 934 1192 940 1193
rect 948 1192 950 1230
rect 990 1229 996 1230
rect 990 1225 991 1229
rect 995 1225 996 1229
rect 990 1224 996 1225
rect 1054 1229 1060 1230
rect 1054 1225 1055 1229
rect 1059 1225 1060 1229
rect 1054 1224 1060 1225
rect 1118 1229 1124 1230
rect 1118 1225 1119 1229
rect 1123 1225 1124 1229
rect 1118 1224 1124 1225
rect 1176 1224 1178 1246
rect 1182 1243 1183 1247
rect 1187 1243 1188 1247
rect 1182 1242 1188 1243
rect 1246 1247 1252 1248
rect 1246 1243 1247 1247
rect 1251 1243 1252 1247
rect 1246 1242 1252 1243
rect 1310 1247 1316 1248
rect 1310 1243 1311 1247
rect 1315 1243 1316 1247
rect 1310 1242 1316 1243
rect 1374 1247 1380 1248
rect 1374 1243 1375 1247
rect 1379 1243 1380 1247
rect 1374 1242 1380 1243
rect 1438 1247 1444 1248
rect 1438 1243 1439 1247
rect 1443 1243 1444 1247
rect 1486 1247 1487 1251
rect 1491 1247 1492 1251
rect 1504 1248 1506 1253
rect 1544 1248 1546 1253
rect 1584 1249 1586 1253
rect 1582 1248 1588 1249
rect 1486 1246 1492 1247
rect 1502 1247 1508 1248
rect 1438 1242 1444 1243
rect 1294 1235 1300 1236
rect 1294 1231 1295 1235
rect 1299 1231 1300 1235
rect 1294 1230 1300 1231
rect 1182 1229 1188 1230
rect 1182 1225 1183 1229
rect 1187 1225 1188 1229
rect 1182 1224 1188 1225
rect 1246 1229 1252 1230
rect 1246 1225 1247 1229
rect 1251 1225 1252 1229
rect 1246 1224 1252 1225
rect 983 1222 987 1223
rect 983 1216 987 1218
rect 991 1222 995 1224
rect 1046 1223 1052 1224
rect 991 1217 995 1218
rect 1039 1222 1043 1223
rect 1046 1219 1047 1223
rect 1051 1219 1052 1223
rect 1046 1218 1052 1219
rect 1055 1222 1059 1224
rect 1039 1216 1043 1218
rect 982 1215 988 1216
rect 982 1211 983 1215
rect 987 1211 988 1215
rect 982 1210 988 1211
rect 1038 1215 1044 1216
rect 1038 1211 1039 1215
rect 1043 1211 1044 1215
rect 1038 1210 1044 1211
rect 998 1207 1004 1208
rect 998 1203 999 1207
rect 1003 1203 1004 1207
rect 998 1202 1004 1203
rect 982 1197 988 1198
rect 982 1193 983 1197
rect 987 1193 988 1197
rect 982 1192 988 1193
rect 264 1187 266 1192
rect 294 1191 300 1192
rect 294 1187 295 1191
rect 299 1187 300 1191
rect 312 1187 314 1192
rect 360 1187 362 1192
rect 416 1187 418 1192
rect 422 1191 428 1192
rect 422 1187 423 1191
rect 427 1187 428 1191
rect 472 1187 474 1192
rect 528 1187 530 1192
rect 584 1187 586 1192
rect 610 1191 616 1192
rect 610 1187 611 1191
rect 615 1187 616 1191
rect 640 1187 642 1192
rect 688 1187 690 1192
rect 702 1191 708 1192
rect 702 1187 703 1191
rect 707 1187 708 1191
rect 736 1187 738 1192
rect 784 1187 786 1192
rect 832 1187 834 1192
rect 880 1187 882 1192
rect 936 1187 938 1192
rect 946 1191 952 1192
rect 946 1187 947 1191
rect 951 1187 952 1191
rect 984 1187 986 1192
rect 255 1186 259 1187
rect 255 1181 259 1182
rect 263 1186 267 1187
rect 294 1186 300 1187
rect 303 1186 307 1187
rect 263 1181 267 1182
rect 303 1181 307 1182
rect 311 1186 315 1187
rect 311 1181 315 1182
rect 359 1186 363 1187
rect 359 1181 363 1182
rect 415 1186 419 1187
rect 422 1186 428 1187
rect 471 1186 475 1187
rect 415 1181 419 1182
rect 230 1179 236 1180
rect 110 1172 111 1176
rect 115 1172 116 1176
rect 110 1171 116 1172
rect 142 1175 148 1176
rect 142 1171 143 1175
rect 147 1171 148 1175
rect 142 1170 148 1171
rect 174 1175 180 1176
rect 174 1171 175 1175
rect 179 1171 180 1175
rect 174 1170 180 1171
rect 214 1175 220 1176
rect 214 1171 215 1175
rect 219 1171 220 1175
rect 230 1175 231 1179
rect 235 1175 236 1179
rect 256 1176 258 1181
rect 304 1176 306 1181
rect 360 1176 362 1181
rect 416 1176 418 1181
rect 230 1174 236 1175
rect 254 1175 260 1176
rect 214 1170 220 1171
rect 254 1171 255 1175
rect 259 1171 260 1175
rect 254 1170 260 1171
rect 302 1175 308 1176
rect 302 1171 303 1175
rect 307 1171 308 1175
rect 302 1170 308 1171
rect 358 1175 364 1176
rect 358 1171 359 1175
rect 363 1171 364 1175
rect 358 1170 364 1171
rect 414 1175 420 1176
rect 414 1171 415 1175
rect 419 1171 420 1175
rect 414 1170 420 1171
rect 424 1171 426 1186
rect 471 1181 475 1182
rect 527 1186 531 1187
rect 527 1181 531 1182
rect 583 1186 587 1187
rect 583 1181 587 1182
rect 591 1186 595 1187
rect 610 1186 616 1187
rect 639 1186 643 1187
rect 591 1181 595 1182
rect 472 1176 474 1181
rect 518 1179 524 1180
rect 470 1175 476 1176
rect 470 1171 471 1175
rect 475 1171 476 1175
rect 518 1175 519 1179
rect 523 1175 524 1179
rect 528 1176 530 1181
rect 592 1176 594 1181
rect 518 1174 524 1175
rect 526 1175 532 1176
rect 424 1169 434 1171
rect 470 1170 476 1171
rect 432 1164 434 1169
rect 154 1163 160 1164
rect 110 1159 116 1160
rect 110 1155 111 1159
rect 115 1155 116 1159
rect 154 1159 155 1163
rect 159 1159 160 1163
rect 154 1158 160 1159
rect 430 1163 436 1164
rect 430 1159 431 1163
rect 435 1159 436 1163
rect 430 1158 436 1159
rect 110 1154 116 1155
rect 142 1157 148 1158
rect 112 1151 114 1154
rect 142 1153 143 1157
rect 147 1153 148 1157
rect 142 1152 148 1153
rect 111 1150 115 1151
rect 111 1145 115 1146
rect 135 1150 139 1151
rect 112 1142 114 1145
rect 135 1144 139 1146
rect 143 1150 147 1152
rect 143 1145 147 1146
rect 134 1143 140 1144
rect 110 1141 116 1142
rect 110 1137 111 1141
rect 115 1137 116 1141
rect 134 1139 135 1143
rect 139 1139 140 1143
rect 134 1138 140 1139
rect 110 1136 116 1137
rect 134 1125 140 1126
rect 110 1124 116 1125
rect 110 1120 111 1124
rect 115 1120 116 1124
rect 134 1121 135 1125
rect 139 1121 140 1125
rect 156 1124 158 1158
rect 174 1157 180 1158
rect 174 1153 175 1157
rect 179 1153 180 1157
rect 174 1152 180 1153
rect 214 1157 220 1158
rect 214 1153 215 1157
rect 219 1153 220 1157
rect 214 1152 220 1153
rect 254 1157 260 1158
rect 254 1153 255 1157
rect 259 1153 260 1157
rect 254 1152 260 1153
rect 302 1157 308 1158
rect 302 1153 303 1157
rect 307 1153 308 1157
rect 302 1152 308 1153
rect 358 1157 364 1158
rect 358 1153 359 1157
rect 363 1153 364 1157
rect 358 1152 364 1153
rect 414 1157 420 1158
rect 414 1153 415 1157
rect 419 1153 420 1157
rect 414 1152 420 1153
rect 470 1157 476 1158
rect 470 1153 471 1157
rect 475 1153 476 1157
rect 470 1152 476 1153
rect 520 1152 522 1174
rect 526 1171 527 1175
rect 531 1171 532 1175
rect 526 1170 532 1171
rect 590 1175 596 1176
rect 590 1171 591 1175
rect 595 1171 596 1175
rect 590 1170 596 1171
rect 612 1164 614 1186
rect 639 1181 643 1182
rect 655 1186 659 1187
rect 655 1181 659 1182
rect 687 1186 691 1187
rect 702 1186 708 1187
rect 719 1186 723 1187
rect 687 1181 691 1182
rect 719 1181 723 1182
rect 735 1186 739 1187
rect 735 1181 739 1182
rect 783 1186 787 1187
rect 783 1181 787 1182
rect 791 1186 795 1187
rect 791 1181 795 1182
rect 831 1186 835 1187
rect 831 1181 835 1182
rect 855 1186 859 1187
rect 855 1181 859 1182
rect 879 1186 883 1187
rect 879 1181 883 1182
rect 919 1186 923 1187
rect 919 1181 923 1182
rect 935 1186 939 1187
rect 946 1186 952 1187
rect 983 1186 987 1187
rect 935 1181 939 1182
rect 983 1181 987 1182
rect 656 1176 658 1181
rect 720 1176 722 1181
rect 792 1176 794 1181
rect 802 1179 808 1180
rect 654 1175 660 1176
rect 654 1171 655 1175
rect 659 1171 660 1175
rect 654 1170 660 1171
rect 718 1175 724 1176
rect 718 1171 719 1175
rect 723 1171 724 1175
rect 718 1170 724 1171
rect 790 1175 796 1176
rect 790 1171 791 1175
rect 795 1171 796 1175
rect 802 1175 803 1179
rect 807 1175 808 1179
rect 856 1176 858 1181
rect 920 1176 922 1181
rect 984 1176 986 1181
rect 1000 1180 1002 1202
rect 1038 1197 1044 1198
rect 1038 1193 1039 1197
rect 1043 1193 1044 1197
rect 1038 1192 1044 1193
rect 1048 1192 1050 1218
rect 1055 1217 1059 1218
rect 1095 1222 1099 1223
rect 1095 1216 1099 1218
rect 1119 1222 1123 1224
rect 1174 1223 1180 1224
rect 1119 1217 1123 1218
rect 1159 1222 1163 1223
rect 1174 1219 1175 1223
rect 1179 1219 1180 1223
rect 1174 1218 1180 1219
rect 1183 1222 1187 1224
rect 1159 1216 1163 1218
rect 1183 1217 1187 1218
rect 1231 1222 1235 1223
rect 1231 1216 1235 1218
rect 1247 1222 1251 1224
rect 1247 1217 1251 1218
rect 1094 1215 1100 1216
rect 1094 1211 1095 1215
rect 1099 1211 1100 1215
rect 1094 1210 1100 1211
rect 1158 1215 1164 1216
rect 1158 1211 1159 1215
rect 1163 1211 1164 1215
rect 1158 1210 1164 1211
rect 1230 1215 1236 1216
rect 1230 1211 1231 1215
rect 1235 1211 1236 1215
rect 1230 1210 1236 1211
rect 1094 1197 1100 1198
rect 1094 1193 1095 1197
rect 1099 1193 1100 1197
rect 1094 1192 1100 1193
rect 1158 1197 1164 1198
rect 1158 1193 1159 1197
rect 1163 1193 1164 1197
rect 1158 1192 1164 1193
rect 1230 1197 1236 1198
rect 1230 1193 1231 1197
rect 1235 1193 1236 1197
rect 1230 1192 1236 1193
rect 1296 1192 1298 1230
rect 1310 1229 1316 1230
rect 1310 1225 1311 1229
rect 1315 1225 1316 1229
rect 1310 1224 1316 1225
rect 1374 1229 1380 1230
rect 1374 1225 1375 1229
rect 1379 1225 1380 1229
rect 1374 1224 1380 1225
rect 1438 1229 1444 1230
rect 1438 1225 1439 1229
rect 1443 1225 1444 1229
rect 1438 1224 1444 1225
rect 1303 1222 1307 1223
rect 1303 1216 1307 1218
rect 1311 1222 1315 1224
rect 1311 1217 1315 1218
rect 1375 1222 1379 1224
rect 1375 1217 1379 1218
rect 1383 1222 1387 1223
rect 1383 1216 1387 1218
rect 1439 1222 1443 1224
rect 1439 1217 1443 1218
rect 1471 1222 1475 1223
rect 1471 1216 1475 1218
rect 1302 1215 1308 1216
rect 1302 1211 1303 1215
rect 1307 1211 1308 1215
rect 1302 1210 1308 1211
rect 1382 1215 1388 1216
rect 1382 1211 1383 1215
rect 1387 1211 1388 1215
rect 1382 1210 1388 1211
rect 1470 1215 1476 1216
rect 1470 1211 1471 1215
rect 1475 1211 1476 1215
rect 1470 1210 1476 1211
rect 1488 1208 1490 1246
rect 1502 1243 1503 1247
rect 1507 1243 1508 1247
rect 1502 1242 1508 1243
rect 1542 1247 1548 1248
rect 1542 1243 1543 1247
rect 1547 1243 1548 1247
rect 1582 1244 1583 1248
rect 1587 1244 1588 1248
rect 1582 1243 1588 1244
rect 1542 1242 1548 1243
rect 1558 1235 1564 1236
rect 1558 1231 1559 1235
rect 1563 1231 1564 1235
rect 1558 1230 1564 1231
rect 1582 1231 1588 1232
rect 1502 1229 1508 1230
rect 1502 1225 1503 1229
rect 1507 1225 1508 1229
rect 1502 1224 1508 1225
rect 1542 1229 1548 1230
rect 1542 1225 1543 1229
rect 1547 1225 1548 1229
rect 1542 1224 1548 1225
rect 1503 1222 1507 1224
rect 1503 1217 1507 1218
rect 1543 1222 1547 1224
rect 1543 1216 1547 1218
rect 1542 1215 1548 1216
rect 1542 1211 1543 1215
rect 1547 1211 1548 1215
rect 1542 1210 1548 1211
rect 1486 1207 1492 1208
rect 1486 1203 1487 1207
rect 1491 1203 1492 1207
rect 1486 1202 1492 1203
rect 1302 1197 1308 1198
rect 1302 1193 1303 1197
rect 1307 1193 1308 1197
rect 1302 1192 1308 1193
rect 1382 1197 1388 1198
rect 1382 1193 1383 1197
rect 1387 1193 1388 1197
rect 1382 1192 1388 1193
rect 1470 1197 1476 1198
rect 1470 1193 1471 1197
rect 1475 1193 1476 1197
rect 1470 1192 1476 1193
rect 1542 1197 1548 1198
rect 1542 1193 1543 1197
rect 1547 1193 1548 1197
rect 1542 1192 1548 1193
rect 1560 1192 1562 1230
rect 1582 1227 1583 1231
rect 1587 1227 1588 1231
rect 1582 1226 1588 1227
rect 1584 1223 1586 1226
rect 1583 1222 1587 1223
rect 1583 1217 1587 1218
rect 1584 1214 1586 1217
rect 1582 1213 1588 1214
rect 1582 1209 1583 1213
rect 1587 1209 1588 1213
rect 1582 1208 1588 1209
rect 1582 1196 1588 1197
rect 1582 1192 1583 1196
rect 1587 1192 1588 1196
rect 1040 1187 1042 1192
rect 1046 1191 1052 1192
rect 1046 1187 1047 1191
rect 1051 1187 1052 1191
rect 1096 1187 1098 1192
rect 1160 1187 1162 1192
rect 1232 1187 1234 1192
rect 1294 1191 1300 1192
rect 1294 1187 1295 1191
rect 1299 1187 1300 1191
rect 1304 1187 1306 1192
rect 1384 1187 1386 1192
rect 1472 1187 1474 1192
rect 1544 1187 1546 1192
rect 1558 1191 1564 1192
rect 1582 1191 1588 1192
rect 1558 1187 1559 1191
rect 1563 1187 1564 1191
rect 1584 1187 1586 1191
rect 1039 1186 1043 1187
rect 1046 1186 1052 1187
rect 1095 1186 1099 1187
rect 1039 1181 1043 1182
rect 1095 1181 1099 1182
rect 1103 1186 1107 1187
rect 1103 1181 1107 1182
rect 1159 1186 1163 1187
rect 1159 1181 1163 1182
rect 1167 1186 1171 1187
rect 1167 1181 1171 1182
rect 1231 1186 1235 1187
rect 1231 1181 1235 1182
rect 1239 1186 1243 1187
rect 1294 1186 1300 1187
rect 1303 1186 1307 1187
rect 1239 1181 1243 1182
rect 1303 1181 1307 1182
rect 1311 1186 1315 1187
rect 1311 1181 1315 1182
rect 1383 1186 1387 1187
rect 1383 1181 1387 1182
rect 1391 1186 1395 1187
rect 1391 1181 1395 1182
rect 1471 1186 1475 1187
rect 1471 1181 1475 1182
rect 1479 1186 1483 1187
rect 1479 1181 1483 1182
rect 1543 1186 1547 1187
rect 1558 1186 1564 1187
rect 1583 1186 1587 1187
rect 1543 1181 1547 1182
rect 1583 1181 1587 1182
rect 998 1179 1004 1180
rect 802 1174 808 1175
rect 854 1175 860 1176
rect 790 1170 796 1171
rect 610 1163 616 1164
rect 610 1159 611 1163
rect 615 1159 616 1163
rect 610 1158 616 1159
rect 526 1157 532 1158
rect 526 1153 527 1157
rect 531 1153 532 1157
rect 526 1152 532 1153
rect 590 1157 596 1158
rect 590 1153 591 1157
rect 595 1153 596 1157
rect 590 1152 596 1153
rect 654 1157 660 1158
rect 654 1153 655 1157
rect 659 1153 660 1157
rect 654 1152 660 1153
rect 718 1157 724 1158
rect 718 1153 719 1157
rect 723 1153 724 1157
rect 718 1152 724 1153
rect 790 1157 796 1158
rect 790 1153 791 1157
rect 795 1153 796 1157
rect 790 1152 796 1153
rect 167 1150 171 1151
rect 167 1144 171 1146
rect 175 1150 179 1152
rect 175 1145 179 1146
rect 199 1150 203 1151
rect 199 1144 203 1146
rect 215 1150 219 1152
rect 215 1145 219 1146
rect 231 1150 235 1151
rect 231 1144 235 1146
rect 255 1150 259 1152
rect 255 1145 259 1146
rect 263 1150 267 1151
rect 263 1144 267 1146
rect 295 1150 299 1151
rect 295 1144 299 1146
rect 303 1150 307 1152
rect 303 1145 307 1146
rect 327 1150 331 1151
rect 327 1144 331 1146
rect 359 1150 363 1152
rect 359 1144 363 1146
rect 391 1150 395 1151
rect 391 1144 395 1146
rect 415 1150 419 1152
rect 415 1145 419 1146
rect 447 1150 451 1151
rect 447 1144 451 1146
rect 471 1150 475 1152
rect 518 1151 524 1152
rect 471 1145 475 1146
rect 503 1150 507 1151
rect 518 1147 519 1151
rect 523 1147 524 1151
rect 518 1146 524 1147
rect 527 1150 531 1152
rect 503 1144 507 1146
rect 527 1145 531 1146
rect 559 1150 563 1151
rect 559 1144 563 1146
rect 591 1150 595 1152
rect 591 1145 595 1146
rect 615 1150 619 1151
rect 615 1144 619 1146
rect 655 1150 659 1152
rect 655 1145 659 1146
rect 671 1150 675 1151
rect 671 1144 675 1146
rect 719 1150 723 1152
rect 719 1145 723 1146
rect 727 1150 731 1151
rect 727 1144 731 1146
rect 783 1150 787 1151
rect 783 1144 787 1146
rect 791 1150 795 1152
rect 791 1145 795 1146
rect 166 1143 172 1144
rect 166 1139 167 1143
rect 171 1139 172 1143
rect 166 1138 172 1139
rect 198 1143 204 1144
rect 198 1139 199 1143
rect 203 1139 204 1143
rect 198 1138 204 1139
rect 230 1143 236 1144
rect 230 1139 231 1143
rect 235 1139 236 1143
rect 230 1138 236 1139
rect 262 1143 268 1144
rect 262 1139 263 1143
rect 267 1139 268 1143
rect 262 1138 268 1139
rect 294 1143 300 1144
rect 294 1139 295 1143
rect 299 1139 300 1143
rect 294 1138 300 1139
rect 326 1143 332 1144
rect 326 1139 327 1143
rect 331 1139 332 1143
rect 326 1138 332 1139
rect 358 1143 364 1144
rect 358 1139 359 1143
rect 363 1139 364 1143
rect 358 1138 364 1139
rect 390 1143 396 1144
rect 390 1139 391 1143
rect 395 1139 396 1143
rect 390 1138 396 1139
rect 446 1143 452 1144
rect 446 1139 447 1143
rect 451 1139 452 1143
rect 446 1138 452 1139
rect 502 1143 508 1144
rect 502 1139 503 1143
rect 507 1139 508 1143
rect 502 1138 508 1139
rect 558 1143 564 1144
rect 558 1139 559 1143
rect 563 1139 564 1143
rect 558 1138 564 1139
rect 614 1143 620 1144
rect 614 1139 615 1143
rect 619 1139 620 1143
rect 614 1138 620 1139
rect 670 1143 676 1144
rect 670 1139 671 1143
rect 675 1139 676 1143
rect 670 1138 676 1139
rect 726 1143 732 1144
rect 726 1139 727 1143
rect 731 1139 732 1143
rect 726 1138 732 1139
rect 782 1143 788 1144
rect 782 1139 783 1143
rect 787 1139 788 1143
rect 782 1138 788 1139
rect 804 1136 806 1174
rect 854 1171 855 1175
rect 859 1171 860 1175
rect 854 1170 860 1171
rect 918 1175 924 1176
rect 918 1171 919 1175
rect 923 1171 924 1175
rect 918 1170 924 1171
rect 982 1175 988 1176
rect 982 1171 983 1175
rect 987 1171 988 1175
rect 998 1175 999 1179
rect 1003 1175 1004 1179
rect 1040 1176 1042 1181
rect 1104 1176 1106 1181
rect 1168 1176 1170 1181
rect 1240 1176 1242 1181
rect 1312 1176 1314 1181
rect 1392 1176 1394 1181
rect 1480 1176 1482 1181
rect 1494 1179 1500 1180
rect 998 1174 1004 1175
rect 1038 1175 1044 1176
rect 982 1170 988 1171
rect 1038 1171 1039 1175
rect 1043 1171 1044 1175
rect 1038 1170 1044 1171
rect 1102 1175 1108 1176
rect 1102 1171 1103 1175
rect 1107 1171 1108 1175
rect 1102 1170 1108 1171
rect 1166 1175 1172 1176
rect 1166 1171 1167 1175
rect 1171 1171 1172 1175
rect 1166 1170 1172 1171
rect 1238 1175 1244 1176
rect 1238 1171 1239 1175
rect 1243 1171 1244 1175
rect 1238 1170 1244 1171
rect 1310 1175 1316 1176
rect 1310 1171 1311 1175
rect 1315 1171 1316 1175
rect 1310 1170 1316 1171
rect 1390 1175 1396 1176
rect 1390 1171 1391 1175
rect 1395 1171 1396 1175
rect 1390 1170 1396 1171
rect 1478 1175 1484 1176
rect 1478 1171 1479 1175
rect 1483 1171 1484 1175
rect 1494 1175 1495 1179
rect 1499 1175 1500 1179
rect 1544 1176 1546 1181
rect 1584 1177 1586 1181
rect 1582 1176 1588 1177
rect 1494 1174 1500 1175
rect 1542 1175 1548 1176
rect 1478 1170 1484 1171
rect 866 1163 872 1164
rect 866 1159 867 1163
rect 871 1159 872 1163
rect 866 1158 872 1159
rect 1418 1163 1424 1164
rect 1418 1159 1419 1163
rect 1423 1159 1424 1163
rect 1418 1158 1424 1159
rect 854 1157 860 1158
rect 854 1153 855 1157
rect 859 1153 860 1157
rect 854 1152 860 1153
rect 839 1150 843 1151
rect 839 1144 843 1146
rect 855 1150 859 1152
rect 855 1145 859 1146
rect 838 1143 844 1144
rect 838 1139 839 1143
rect 843 1139 844 1143
rect 838 1138 844 1139
rect 310 1135 316 1136
rect 310 1131 311 1135
rect 315 1131 316 1135
rect 310 1130 316 1131
rect 802 1135 808 1136
rect 802 1131 803 1135
rect 807 1131 808 1135
rect 802 1130 808 1131
rect 166 1125 172 1126
rect 134 1120 140 1121
rect 154 1123 160 1124
rect 110 1119 116 1120
rect 112 1115 114 1119
rect 136 1115 138 1120
rect 154 1119 155 1123
rect 159 1119 160 1123
rect 166 1121 167 1125
rect 171 1121 172 1125
rect 166 1120 172 1121
rect 198 1125 204 1126
rect 198 1121 199 1125
rect 203 1121 204 1125
rect 198 1120 204 1121
rect 230 1125 236 1126
rect 230 1121 231 1125
rect 235 1121 236 1125
rect 230 1120 236 1121
rect 262 1125 268 1126
rect 262 1121 263 1125
rect 267 1121 268 1125
rect 262 1120 268 1121
rect 294 1125 300 1126
rect 294 1121 295 1125
rect 299 1121 300 1125
rect 294 1120 300 1121
rect 154 1118 160 1119
rect 168 1115 170 1120
rect 200 1115 202 1120
rect 232 1115 234 1120
rect 264 1115 266 1120
rect 296 1115 298 1120
rect 111 1114 115 1115
rect 111 1109 115 1110
rect 135 1114 139 1115
rect 135 1109 139 1110
rect 151 1114 155 1115
rect 151 1109 155 1110
rect 167 1114 171 1115
rect 167 1109 171 1110
rect 183 1114 187 1115
rect 183 1109 187 1110
rect 199 1114 203 1115
rect 199 1109 203 1110
rect 223 1114 227 1115
rect 223 1109 227 1110
rect 231 1114 235 1115
rect 231 1109 235 1110
rect 263 1114 267 1115
rect 263 1109 267 1110
rect 271 1114 275 1115
rect 271 1109 275 1110
rect 295 1114 299 1115
rect 295 1109 299 1110
rect 112 1105 114 1109
rect 110 1104 116 1105
rect 152 1104 154 1109
rect 184 1104 186 1109
rect 224 1104 226 1109
rect 272 1104 274 1109
rect 110 1100 111 1104
rect 115 1100 116 1104
rect 110 1099 116 1100
rect 150 1103 156 1104
rect 150 1099 151 1103
rect 155 1099 156 1103
rect 150 1098 156 1099
rect 166 1103 172 1104
rect 166 1098 167 1103
rect 171 1098 172 1103
rect 182 1103 188 1104
rect 182 1099 183 1103
rect 187 1099 188 1103
rect 182 1098 188 1099
rect 222 1103 228 1104
rect 222 1099 223 1103
rect 227 1099 228 1103
rect 222 1098 228 1099
rect 270 1103 276 1104
rect 270 1099 271 1103
rect 275 1099 276 1103
rect 312 1101 314 1130
rect 326 1125 332 1126
rect 326 1121 327 1125
rect 331 1121 332 1125
rect 326 1120 332 1121
rect 358 1125 364 1126
rect 358 1121 359 1125
rect 363 1121 364 1125
rect 358 1120 364 1121
rect 390 1125 396 1126
rect 390 1121 391 1125
rect 395 1121 396 1125
rect 390 1120 396 1121
rect 446 1125 452 1126
rect 446 1121 447 1125
rect 451 1121 452 1125
rect 446 1120 452 1121
rect 502 1125 508 1126
rect 502 1121 503 1125
rect 507 1121 508 1125
rect 502 1120 508 1121
rect 558 1125 564 1126
rect 558 1121 559 1125
rect 563 1121 564 1125
rect 558 1120 564 1121
rect 614 1125 620 1126
rect 614 1121 615 1125
rect 619 1121 620 1125
rect 614 1120 620 1121
rect 670 1125 676 1126
rect 670 1121 671 1125
rect 675 1121 676 1125
rect 670 1120 676 1121
rect 726 1125 732 1126
rect 726 1121 727 1125
rect 731 1121 732 1125
rect 726 1120 732 1121
rect 782 1125 788 1126
rect 782 1121 783 1125
rect 787 1121 788 1125
rect 782 1120 788 1121
rect 838 1125 844 1126
rect 838 1121 839 1125
rect 843 1121 844 1125
rect 838 1120 844 1121
rect 868 1120 870 1158
rect 918 1157 924 1158
rect 918 1153 919 1157
rect 923 1153 924 1157
rect 918 1152 924 1153
rect 982 1157 988 1158
rect 982 1153 983 1157
rect 987 1153 988 1157
rect 982 1152 988 1153
rect 1038 1157 1044 1158
rect 1038 1153 1039 1157
rect 1043 1153 1044 1157
rect 1038 1152 1044 1153
rect 1102 1157 1108 1158
rect 1102 1153 1103 1157
rect 1107 1153 1108 1157
rect 1102 1152 1108 1153
rect 1166 1157 1172 1158
rect 1166 1153 1167 1157
rect 1171 1153 1172 1157
rect 1166 1152 1172 1153
rect 1238 1157 1244 1158
rect 1238 1153 1239 1157
rect 1243 1153 1244 1157
rect 1238 1152 1244 1153
rect 1310 1157 1316 1158
rect 1310 1153 1311 1157
rect 1315 1153 1316 1157
rect 1310 1152 1316 1153
rect 1390 1157 1396 1158
rect 1390 1153 1391 1157
rect 1395 1153 1396 1157
rect 1390 1152 1396 1153
rect 874 1151 880 1152
rect 874 1147 875 1151
rect 879 1147 880 1151
rect 874 1146 880 1147
rect 895 1150 899 1151
rect 328 1115 330 1120
rect 346 1119 352 1120
rect 346 1115 347 1119
rect 351 1115 352 1119
rect 360 1115 362 1120
rect 392 1115 394 1120
rect 448 1115 450 1120
rect 504 1115 506 1120
rect 560 1115 562 1120
rect 606 1119 612 1120
rect 606 1115 607 1119
rect 611 1115 612 1119
rect 616 1115 618 1120
rect 672 1115 674 1120
rect 728 1115 730 1120
rect 784 1115 786 1120
rect 840 1115 842 1120
rect 866 1119 872 1120
rect 866 1115 867 1119
rect 871 1115 872 1119
rect 327 1114 331 1115
rect 346 1114 352 1115
rect 359 1114 363 1115
rect 327 1109 331 1110
rect 328 1104 330 1109
rect 326 1103 332 1104
rect 270 1098 276 1099
rect 311 1100 315 1101
rect 167 1095 171 1096
rect 326 1099 327 1103
rect 331 1099 332 1103
rect 326 1098 332 1099
rect 311 1095 315 1096
rect 110 1087 116 1088
rect 110 1083 111 1087
rect 115 1083 116 1087
rect 110 1082 116 1083
rect 150 1085 156 1086
rect 112 1071 114 1082
rect 150 1081 151 1085
rect 155 1081 156 1085
rect 150 1080 156 1081
rect 182 1085 188 1086
rect 182 1081 183 1085
rect 187 1081 188 1085
rect 182 1080 188 1081
rect 222 1085 228 1086
rect 222 1081 223 1085
rect 227 1081 228 1085
rect 222 1080 228 1081
rect 270 1085 276 1086
rect 270 1081 271 1085
rect 275 1081 276 1085
rect 270 1080 276 1081
rect 326 1085 332 1086
rect 326 1081 327 1085
rect 331 1081 332 1085
rect 326 1080 332 1081
rect 348 1080 350 1114
rect 359 1109 363 1110
rect 383 1114 387 1115
rect 383 1109 387 1110
rect 391 1114 395 1115
rect 391 1109 395 1110
rect 439 1114 443 1115
rect 439 1109 443 1110
rect 447 1114 451 1115
rect 447 1109 451 1110
rect 503 1114 507 1115
rect 503 1109 507 1110
rect 559 1114 563 1115
rect 559 1109 563 1110
rect 567 1114 571 1115
rect 606 1114 612 1115
rect 615 1114 619 1115
rect 567 1109 571 1110
rect 384 1104 386 1109
rect 440 1104 442 1109
rect 494 1107 500 1108
rect 382 1103 388 1104
rect 382 1099 383 1103
rect 387 1099 388 1103
rect 382 1098 388 1099
rect 438 1103 444 1104
rect 438 1099 439 1103
rect 443 1099 444 1103
rect 494 1103 495 1107
rect 499 1103 500 1107
rect 504 1104 506 1109
rect 568 1104 570 1109
rect 494 1102 500 1103
rect 502 1103 508 1104
rect 438 1098 444 1099
rect 382 1085 388 1086
rect 382 1081 383 1085
rect 387 1081 388 1085
rect 382 1080 388 1081
rect 438 1085 444 1086
rect 438 1081 439 1085
rect 443 1081 444 1085
rect 438 1080 444 1081
rect 152 1071 154 1080
rect 184 1071 186 1080
rect 224 1071 226 1080
rect 272 1071 274 1080
rect 328 1071 330 1080
rect 346 1079 352 1080
rect 346 1075 347 1079
rect 351 1075 352 1079
rect 346 1074 352 1075
rect 384 1071 386 1080
rect 440 1071 442 1080
rect 496 1072 498 1102
rect 502 1099 503 1103
rect 507 1099 508 1103
rect 502 1098 508 1099
rect 566 1103 572 1104
rect 566 1099 567 1103
rect 571 1099 572 1103
rect 566 1098 572 1099
rect 502 1085 508 1086
rect 502 1081 503 1085
rect 507 1081 508 1085
rect 502 1080 508 1081
rect 566 1085 572 1086
rect 566 1081 567 1085
rect 571 1081 572 1085
rect 566 1080 572 1081
rect 608 1080 610 1114
rect 615 1109 619 1110
rect 639 1114 643 1115
rect 639 1109 643 1110
rect 671 1114 675 1115
rect 671 1109 675 1110
rect 711 1114 715 1115
rect 711 1109 715 1110
rect 727 1114 731 1115
rect 727 1109 731 1110
rect 783 1114 787 1115
rect 783 1109 787 1110
rect 839 1114 843 1115
rect 839 1109 843 1110
rect 855 1114 859 1115
rect 866 1114 872 1115
rect 855 1109 859 1110
rect 640 1104 642 1109
rect 712 1104 714 1109
rect 784 1104 786 1109
rect 856 1104 858 1109
rect 876 1108 878 1146
rect 895 1144 899 1146
rect 919 1150 923 1152
rect 919 1145 923 1146
rect 951 1150 955 1151
rect 951 1144 955 1146
rect 983 1150 987 1152
rect 983 1145 987 1146
rect 1007 1150 1011 1151
rect 1007 1144 1011 1146
rect 1039 1150 1043 1152
rect 1039 1145 1043 1146
rect 1063 1150 1067 1151
rect 1063 1144 1067 1146
rect 1103 1150 1107 1152
rect 1103 1145 1107 1146
rect 1127 1150 1131 1151
rect 1127 1144 1131 1146
rect 1167 1150 1171 1152
rect 1226 1151 1232 1152
rect 1167 1145 1171 1146
rect 1191 1150 1195 1151
rect 1226 1147 1227 1151
rect 1231 1147 1232 1151
rect 1226 1146 1232 1147
rect 1239 1150 1243 1152
rect 1191 1144 1195 1146
rect 894 1143 900 1144
rect 894 1139 895 1143
rect 899 1139 900 1143
rect 894 1138 900 1139
rect 950 1143 956 1144
rect 950 1139 951 1143
rect 955 1139 956 1143
rect 950 1138 956 1139
rect 1006 1143 1012 1144
rect 1006 1139 1007 1143
rect 1011 1139 1012 1143
rect 1006 1138 1012 1139
rect 1062 1143 1068 1144
rect 1062 1139 1063 1143
rect 1067 1139 1068 1143
rect 1062 1138 1068 1139
rect 1126 1143 1132 1144
rect 1126 1139 1127 1143
rect 1131 1139 1132 1143
rect 1126 1138 1132 1139
rect 1190 1143 1196 1144
rect 1190 1139 1191 1143
rect 1195 1139 1196 1143
rect 1190 1138 1196 1139
rect 894 1125 900 1126
rect 894 1121 895 1125
rect 899 1121 900 1125
rect 894 1120 900 1121
rect 950 1125 956 1126
rect 950 1121 951 1125
rect 955 1121 956 1125
rect 950 1120 956 1121
rect 1006 1125 1012 1126
rect 1006 1121 1007 1125
rect 1011 1121 1012 1125
rect 1006 1120 1012 1121
rect 1062 1125 1068 1126
rect 1062 1121 1063 1125
rect 1067 1121 1068 1125
rect 1062 1120 1068 1121
rect 1126 1125 1132 1126
rect 1126 1121 1127 1125
rect 1131 1121 1132 1125
rect 1126 1120 1132 1121
rect 1190 1125 1196 1126
rect 1190 1121 1191 1125
rect 1195 1121 1196 1125
rect 1190 1120 1196 1121
rect 896 1115 898 1120
rect 952 1115 954 1120
rect 1008 1115 1010 1120
rect 1064 1115 1066 1120
rect 1128 1115 1130 1120
rect 1158 1119 1164 1120
rect 1158 1115 1159 1119
rect 1163 1115 1164 1119
rect 1192 1115 1194 1120
rect 895 1114 899 1115
rect 895 1109 899 1110
rect 919 1114 923 1115
rect 919 1109 923 1110
rect 951 1114 955 1115
rect 951 1109 955 1110
rect 983 1114 987 1115
rect 983 1109 987 1110
rect 1007 1114 1011 1115
rect 1007 1109 1011 1110
rect 1039 1114 1043 1115
rect 1039 1109 1043 1110
rect 1063 1114 1067 1115
rect 1063 1109 1067 1110
rect 1095 1114 1099 1115
rect 1095 1109 1099 1110
rect 1127 1114 1131 1115
rect 1127 1109 1131 1110
rect 1151 1114 1155 1115
rect 1158 1114 1164 1115
rect 1191 1114 1195 1115
rect 1151 1109 1155 1110
rect 874 1107 880 1108
rect 638 1103 644 1104
rect 638 1099 639 1103
rect 643 1099 644 1103
rect 638 1098 644 1099
rect 710 1103 716 1104
rect 710 1099 711 1103
rect 715 1099 716 1103
rect 710 1098 716 1099
rect 782 1103 788 1104
rect 782 1099 783 1103
rect 787 1099 788 1103
rect 782 1098 788 1099
rect 854 1103 860 1104
rect 854 1099 855 1103
rect 859 1099 860 1103
rect 874 1103 875 1107
rect 879 1103 880 1107
rect 920 1104 922 1109
rect 984 1104 986 1109
rect 1040 1104 1042 1109
rect 1096 1104 1098 1109
rect 1152 1104 1154 1109
rect 874 1102 880 1103
rect 918 1103 924 1104
rect 854 1098 860 1099
rect 918 1099 919 1103
rect 923 1099 924 1103
rect 918 1098 924 1099
rect 982 1103 988 1104
rect 982 1099 983 1103
rect 987 1099 988 1103
rect 982 1098 988 1099
rect 1038 1103 1044 1104
rect 1038 1099 1039 1103
rect 1043 1099 1044 1103
rect 1038 1098 1044 1099
rect 1094 1103 1100 1104
rect 1094 1099 1095 1103
rect 1099 1099 1100 1103
rect 1094 1098 1100 1099
rect 1150 1103 1156 1104
rect 1150 1099 1151 1103
rect 1155 1099 1156 1103
rect 1150 1098 1156 1099
rect 638 1085 644 1086
rect 638 1081 639 1085
rect 643 1081 644 1085
rect 638 1080 644 1081
rect 710 1085 716 1086
rect 710 1081 711 1085
rect 715 1081 716 1085
rect 710 1080 716 1081
rect 782 1085 788 1086
rect 782 1081 783 1085
rect 787 1081 788 1085
rect 782 1080 788 1081
rect 854 1085 860 1086
rect 854 1081 855 1085
rect 859 1081 860 1085
rect 854 1080 860 1081
rect 918 1085 924 1086
rect 918 1081 919 1085
rect 923 1081 924 1085
rect 918 1080 924 1081
rect 982 1085 988 1086
rect 982 1081 983 1085
rect 987 1081 988 1085
rect 982 1080 988 1081
rect 1038 1085 1044 1086
rect 1038 1081 1039 1085
rect 1043 1081 1044 1085
rect 1038 1080 1044 1081
rect 1094 1085 1100 1086
rect 1094 1081 1095 1085
rect 1099 1081 1100 1085
rect 1094 1080 1100 1081
rect 1150 1085 1156 1086
rect 1150 1081 1151 1085
rect 1155 1081 1156 1085
rect 1150 1080 1156 1081
rect 1160 1080 1162 1114
rect 1191 1109 1195 1110
rect 1207 1114 1211 1115
rect 1207 1109 1211 1110
rect 1208 1104 1210 1109
rect 1228 1108 1230 1146
rect 1239 1145 1243 1146
rect 1255 1150 1259 1151
rect 1255 1144 1259 1146
rect 1311 1150 1315 1152
rect 1311 1145 1315 1146
rect 1327 1150 1331 1151
rect 1327 1144 1331 1146
rect 1391 1150 1395 1152
rect 1391 1145 1395 1146
rect 1399 1150 1403 1151
rect 1399 1144 1403 1146
rect 1254 1143 1260 1144
rect 1254 1139 1255 1143
rect 1259 1139 1260 1143
rect 1254 1138 1260 1139
rect 1326 1143 1332 1144
rect 1326 1139 1327 1143
rect 1331 1139 1332 1143
rect 1326 1138 1332 1139
rect 1398 1143 1404 1144
rect 1398 1139 1399 1143
rect 1403 1139 1404 1143
rect 1398 1138 1404 1139
rect 1254 1125 1260 1126
rect 1254 1121 1255 1125
rect 1259 1121 1260 1125
rect 1254 1120 1260 1121
rect 1326 1125 1332 1126
rect 1326 1121 1327 1125
rect 1331 1121 1332 1125
rect 1326 1120 1332 1121
rect 1398 1125 1404 1126
rect 1398 1121 1399 1125
rect 1403 1121 1404 1125
rect 1398 1120 1404 1121
rect 1256 1115 1258 1120
rect 1328 1115 1330 1120
rect 1400 1115 1402 1120
rect 1255 1114 1259 1115
rect 1255 1109 1259 1110
rect 1263 1114 1267 1115
rect 1263 1109 1267 1110
rect 1319 1114 1323 1115
rect 1319 1109 1323 1110
rect 1327 1114 1331 1115
rect 1327 1109 1331 1110
rect 1375 1114 1379 1115
rect 1375 1109 1379 1110
rect 1399 1114 1403 1115
rect 1399 1109 1403 1110
rect 1410 1111 1416 1112
rect 1226 1107 1232 1108
rect 1206 1103 1212 1104
rect 1206 1099 1207 1103
rect 1211 1099 1212 1103
rect 1226 1103 1227 1107
rect 1231 1103 1232 1107
rect 1264 1104 1266 1109
rect 1320 1104 1322 1109
rect 1376 1104 1378 1109
rect 1410 1107 1411 1111
rect 1415 1107 1416 1111
rect 1410 1106 1416 1107
rect 1226 1102 1232 1103
rect 1262 1103 1268 1104
rect 1206 1098 1212 1099
rect 1262 1099 1263 1103
rect 1267 1099 1268 1103
rect 1262 1098 1268 1099
rect 1318 1103 1324 1104
rect 1318 1099 1319 1103
rect 1323 1099 1324 1103
rect 1318 1098 1324 1099
rect 1374 1103 1380 1104
rect 1374 1099 1375 1103
rect 1379 1099 1380 1103
rect 1374 1098 1380 1099
rect 1166 1091 1172 1092
rect 1166 1087 1167 1091
rect 1171 1087 1172 1091
rect 1166 1086 1172 1087
rect 1390 1091 1396 1092
rect 1390 1087 1391 1091
rect 1395 1087 1396 1091
rect 1390 1086 1396 1087
rect 494 1071 500 1072
rect 504 1071 506 1080
rect 568 1071 570 1080
rect 606 1079 612 1080
rect 606 1075 607 1079
rect 611 1075 612 1079
rect 606 1074 612 1075
rect 640 1071 642 1080
rect 712 1071 714 1080
rect 784 1071 786 1080
rect 856 1071 858 1080
rect 920 1071 922 1080
rect 984 1071 986 1080
rect 1040 1071 1042 1080
rect 1096 1071 1098 1080
rect 1152 1071 1154 1080
rect 1158 1079 1164 1080
rect 1158 1075 1159 1079
rect 1163 1075 1164 1079
rect 1158 1074 1164 1075
rect 111 1070 115 1071
rect 111 1065 115 1066
rect 151 1070 155 1071
rect 151 1065 155 1066
rect 183 1070 187 1071
rect 183 1065 187 1066
rect 223 1070 227 1071
rect 223 1065 227 1066
rect 271 1070 275 1071
rect 271 1065 275 1066
rect 327 1070 331 1071
rect 327 1065 331 1066
rect 383 1070 387 1071
rect 383 1065 387 1066
rect 439 1070 443 1071
rect 439 1065 443 1066
rect 447 1070 451 1071
rect 112 1062 114 1065
rect 447 1064 451 1066
rect 487 1070 491 1071
rect 494 1067 495 1071
rect 499 1067 500 1071
rect 494 1066 500 1067
rect 503 1070 507 1071
rect 487 1064 491 1066
rect 503 1065 507 1066
rect 543 1070 547 1071
rect 543 1064 547 1066
rect 567 1070 571 1071
rect 567 1065 571 1066
rect 599 1070 603 1071
rect 599 1064 603 1066
rect 639 1070 643 1071
rect 639 1065 643 1066
rect 663 1070 667 1071
rect 663 1064 667 1066
rect 711 1070 715 1071
rect 711 1065 715 1066
rect 727 1070 731 1071
rect 727 1064 731 1066
rect 783 1070 787 1071
rect 783 1065 787 1066
rect 791 1070 795 1071
rect 791 1064 795 1066
rect 855 1070 859 1071
rect 855 1065 859 1066
rect 863 1070 867 1071
rect 863 1064 867 1066
rect 919 1070 923 1071
rect 919 1065 923 1066
rect 935 1070 939 1071
rect 935 1064 939 1066
rect 983 1070 987 1071
rect 983 1065 987 1066
rect 1007 1070 1011 1071
rect 1007 1064 1011 1066
rect 1039 1070 1043 1071
rect 1039 1065 1043 1066
rect 1079 1070 1083 1071
rect 1079 1064 1083 1066
rect 1095 1070 1099 1071
rect 1095 1065 1099 1066
rect 1151 1070 1155 1071
rect 1151 1064 1155 1066
rect 446 1063 452 1064
rect 110 1061 116 1062
rect 110 1057 111 1061
rect 115 1057 116 1061
rect 446 1059 447 1063
rect 451 1059 452 1063
rect 446 1058 452 1059
rect 486 1063 492 1064
rect 486 1059 487 1063
rect 491 1059 492 1063
rect 486 1058 492 1059
rect 542 1063 548 1064
rect 542 1059 543 1063
rect 547 1059 548 1063
rect 542 1058 548 1059
rect 598 1063 604 1064
rect 598 1059 599 1063
rect 603 1059 604 1063
rect 598 1058 604 1059
rect 662 1063 668 1064
rect 662 1059 663 1063
rect 667 1059 668 1063
rect 662 1058 668 1059
rect 726 1063 732 1064
rect 726 1059 727 1063
rect 731 1059 732 1063
rect 726 1058 732 1059
rect 790 1063 796 1064
rect 790 1059 791 1063
rect 795 1059 796 1063
rect 790 1058 796 1059
rect 862 1063 868 1064
rect 862 1059 863 1063
rect 867 1059 868 1063
rect 862 1058 868 1059
rect 934 1063 940 1064
rect 934 1059 935 1063
rect 939 1059 940 1063
rect 934 1058 940 1059
rect 1006 1063 1012 1064
rect 1006 1059 1007 1063
rect 1011 1059 1012 1063
rect 1006 1058 1012 1059
rect 1078 1063 1084 1064
rect 1078 1059 1079 1063
rect 1083 1059 1084 1063
rect 1078 1058 1084 1059
rect 1150 1063 1156 1064
rect 1150 1059 1151 1063
rect 1155 1059 1156 1063
rect 1150 1058 1156 1059
rect 110 1056 116 1057
rect 986 1055 992 1056
rect 986 1051 987 1055
rect 991 1051 992 1055
rect 986 1050 992 1051
rect 994 1055 1000 1056
rect 994 1051 995 1055
rect 999 1051 1000 1055
rect 994 1050 1000 1051
rect 446 1045 452 1046
rect 110 1044 116 1045
rect 110 1040 111 1044
rect 115 1040 116 1044
rect 446 1041 447 1045
rect 451 1041 452 1045
rect 446 1040 452 1041
rect 486 1045 492 1046
rect 486 1041 487 1045
rect 491 1041 492 1045
rect 486 1040 492 1041
rect 542 1045 548 1046
rect 542 1041 543 1045
rect 547 1041 548 1045
rect 542 1040 548 1041
rect 598 1045 604 1046
rect 598 1041 599 1045
rect 603 1041 604 1045
rect 598 1040 604 1041
rect 662 1045 668 1046
rect 662 1041 663 1045
rect 667 1041 668 1045
rect 662 1040 668 1041
rect 726 1045 732 1046
rect 726 1041 727 1045
rect 731 1041 732 1045
rect 726 1040 732 1041
rect 790 1045 796 1046
rect 790 1041 791 1045
rect 795 1041 796 1045
rect 790 1040 796 1041
rect 862 1045 868 1046
rect 862 1041 863 1045
rect 867 1041 868 1045
rect 862 1040 868 1041
rect 934 1045 940 1046
rect 934 1041 935 1045
rect 939 1041 940 1045
rect 934 1040 940 1041
rect 110 1039 116 1040
rect 112 1031 114 1039
rect 448 1031 450 1040
rect 488 1031 490 1040
rect 544 1031 546 1040
rect 600 1031 602 1040
rect 664 1031 666 1040
rect 718 1031 724 1032
rect 728 1031 730 1040
rect 792 1031 794 1040
rect 864 1031 866 1040
rect 936 1031 938 1040
rect 111 1030 115 1031
rect 111 1025 115 1026
rect 447 1030 451 1031
rect 447 1025 451 1026
rect 487 1030 491 1031
rect 487 1025 491 1026
rect 511 1030 515 1031
rect 511 1025 515 1026
rect 543 1030 547 1031
rect 543 1025 547 1026
rect 575 1030 579 1031
rect 575 1025 579 1026
rect 599 1030 603 1031
rect 599 1025 603 1026
rect 615 1030 619 1031
rect 615 1025 619 1026
rect 663 1030 667 1031
rect 663 1025 667 1026
rect 711 1030 715 1031
rect 718 1027 719 1031
rect 723 1027 724 1031
rect 718 1026 724 1027
rect 727 1030 731 1031
rect 711 1025 715 1026
rect 112 1021 114 1025
rect 110 1020 116 1021
rect 512 1020 514 1025
rect 544 1020 546 1025
rect 576 1020 578 1025
rect 616 1020 618 1025
rect 626 1023 632 1024
rect 110 1016 111 1020
rect 115 1016 116 1020
rect 110 1015 116 1016
rect 510 1019 516 1020
rect 510 1015 511 1019
rect 515 1015 516 1019
rect 510 1014 516 1015
rect 542 1019 548 1020
rect 542 1015 543 1019
rect 547 1015 548 1019
rect 542 1014 548 1015
rect 574 1019 580 1020
rect 574 1015 575 1019
rect 579 1015 580 1019
rect 574 1014 580 1015
rect 614 1019 620 1020
rect 614 1015 615 1019
rect 619 1015 620 1019
rect 626 1019 627 1023
rect 631 1019 632 1023
rect 664 1020 666 1025
rect 712 1020 714 1025
rect 626 1018 632 1019
rect 662 1019 668 1020
rect 614 1014 620 1015
rect 110 1003 116 1004
rect 110 999 111 1003
rect 115 999 116 1003
rect 110 998 116 999
rect 510 1001 516 1002
rect 112 987 114 998
rect 510 997 511 1001
rect 515 997 516 1001
rect 510 996 516 997
rect 542 1001 548 1002
rect 542 997 543 1001
rect 547 997 548 1001
rect 542 996 548 997
rect 574 1001 580 1002
rect 574 997 575 1001
rect 579 997 580 1001
rect 574 996 580 997
rect 614 1001 620 1002
rect 614 997 615 1001
rect 619 997 620 1001
rect 614 996 620 997
rect 512 987 514 996
rect 544 987 546 996
rect 576 987 578 996
rect 616 987 618 996
rect 628 988 630 1018
rect 662 1015 663 1019
rect 667 1015 668 1019
rect 662 1014 668 1015
rect 710 1019 716 1020
rect 710 1015 711 1019
rect 715 1015 716 1019
rect 710 1014 716 1015
rect 720 1006 722 1026
rect 727 1025 731 1026
rect 775 1030 779 1031
rect 775 1025 779 1026
rect 791 1030 795 1031
rect 791 1025 795 1026
rect 847 1030 851 1031
rect 847 1025 851 1026
rect 863 1030 867 1031
rect 863 1025 867 1026
rect 927 1030 931 1031
rect 927 1025 931 1026
rect 935 1030 939 1031
rect 988 1028 990 1050
rect 996 1036 998 1050
rect 1006 1045 1012 1046
rect 1006 1041 1007 1045
rect 1011 1041 1012 1045
rect 1006 1040 1012 1041
rect 1078 1045 1084 1046
rect 1078 1041 1079 1045
rect 1083 1041 1084 1045
rect 1078 1040 1084 1041
rect 1150 1045 1156 1046
rect 1150 1041 1151 1045
rect 1155 1041 1156 1045
rect 1150 1040 1156 1041
rect 1168 1040 1170 1086
rect 1206 1085 1212 1086
rect 1206 1081 1207 1085
rect 1211 1081 1212 1085
rect 1206 1080 1212 1081
rect 1262 1085 1268 1086
rect 1262 1081 1263 1085
rect 1267 1081 1268 1085
rect 1262 1080 1268 1081
rect 1318 1085 1324 1086
rect 1318 1081 1319 1085
rect 1323 1081 1324 1085
rect 1318 1080 1324 1081
rect 1374 1085 1380 1086
rect 1374 1081 1375 1085
rect 1379 1081 1380 1085
rect 1374 1080 1380 1081
rect 1208 1071 1210 1080
rect 1264 1071 1266 1080
rect 1320 1071 1322 1080
rect 1376 1071 1378 1080
rect 1392 1075 1394 1086
rect 1384 1073 1394 1075
rect 1207 1070 1211 1071
rect 1207 1065 1211 1066
rect 1215 1070 1219 1071
rect 1215 1064 1219 1066
rect 1263 1070 1267 1071
rect 1263 1065 1267 1066
rect 1279 1070 1283 1071
rect 1279 1064 1283 1066
rect 1319 1070 1323 1071
rect 1319 1065 1323 1066
rect 1335 1070 1339 1071
rect 1335 1064 1339 1066
rect 1375 1070 1379 1071
rect 1375 1065 1379 1066
rect 1214 1063 1220 1064
rect 1214 1059 1215 1063
rect 1219 1059 1220 1063
rect 1214 1058 1220 1059
rect 1278 1063 1284 1064
rect 1278 1059 1279 1063
rect 1283 1059 1284 1063
rect 1278 1058 1284 1059
rect 1334 1063 1340 1064
rect 1334 1059 1335 1063
rect 1339 1059 1340 1063
rect 1334 1058 1340 1059
rect 1186 1055 1192 1056
rect 1186 1051 1187 1055
rect 1191 1051 1192 1055
rect 1186 1050 1192 1051
rect 994 1035 1000 1036
rect 994 1031 995 1035
rect 999 1031 1000 1035
rect 1008 1031 1010 1040
rect 1080 1031 1082 1040
rect 1152 1031 1154 1040
rect 1166 1039 1172 1040
rect 1166 1035 1167 1039
rect 1171 1035 1172 1039
rect 1166 1034 1172 1035
rect 994 1030 1000 1031
rect 1007 1030 1011 1031
rect 935 1025 939 1026
rect 986 1027 992 1028
rect 776 1020 778 1025
rect 848 1020 850 1025
rect 928 1020 930 1025
rect 978 1023 984 1024
rect 774 1019 780 1020
rect 774 1015 775 1019
rect 779 1015 780 1019
rect 774 1014 780 1015
rect 846 1019 852 1020
rect 846 1015 847 1019
rect 851 1015 852 1019
rect 846 1014 852 1015
rect 926 1019 932 1020
rect 926 1015 927 1019
rect 931 1015 932 1019
rect 978 1019 979 1023
rect 983 1019 984 1023
rect 986 1023 987 1027
rect 991 1023 992 1027
rect 1007 1025 1011 1026
rect 1079 1030 1083 1031
rect 1079 1025 1083 1026
rect 1087 1030 1091 1031
rect 1087 1025 1091 1026
rect 1151 1030 1155 1031
rect 1151 1025 1155 1026
rect 1167 1030 1171 1031
rect 1167 1025 1171 1026
rect 986 1022 992 1023
rect 1008 1020 1010 1025
rect 1088 1020 1090 1025
rect 1168 1020 1170 1025
rect 1188 1024 1190 1050
rect 1214 1045 1220 1046
rect 1214 1041 1215 1045
rect 1219 1041 1220 1045
rect 1214 1040 1220 1041
rect 1278 1045 1284 1046
rect 1278 1041 1279 1045
rect 1283 1041 1284 1045
rect 1278 1040 1284 1041
rect 1334 1045 1340 1046
rect 1334 1041 1335 1045
rect 1339 1041 1340 1045
rect 1334 1040 1340 1041
rect 1384 1040 1386 1073
rect 1391 1070 1395 1071
rect 1391 1064 1395 1066
rect 1390 1063 1396 1064
rect 1390 1059 1391 1063
rect 1395 1059 1396 1063
rect 1390 1058 1396 1059
rect 1412 1056 1414 1106
rect 1420 1080 1422 1158
rect 1478 1157 1484 1158
rect 1478 1153 1479 1157
rect 1483 1153 1484 1157
rect 1478 1152 1484 1153
rect 1479 1150 1483 1152
rect 1479 1144 1483 1146
rect 1478 1143 1484 1144
rect 1478 1139 1479 1143
rect 1483 1139 1484 1143
rect 1478 1138 1484 1139
rect 1496 1136 1498 1174
rect 1542 1171 1543 1175
rect 1547 1171 1548 1175
rect 1582 1172 1583 1176
rect 1587 1172 1588 1176
rect 1582 1171 1588 1172
rect 1542 1170 1548 1171
rect 1558 1163 1564 1164
rect 1558 1159 1559 1163
rect 1563 1159 1564 1163
rect 1558 1158 1564 1159
rect 1582 1159 1588 1160
rect 1542 1157 1548 1158
rect 1542 1153 1543 1157
rect 1547 1153 1548 1157
rect 1542 1152 1548 1153
rect 1543 1150 1547 1152
rect 1543 1144 1547 1146
rect 1542 1143 1548 1144
rect 1542 1139 1543 1143
rect 1547 1139 1548 1143
rect 1542 1138 1548 1139
rect 1494 1135 1500 1136
rect 1494 1131 1495 1135
rect 1499 1131 1500 1135
rect 1494 1130 1500 1131
rect 1478 1125 1484 1126
rect 1478 1121 1479 1125
rect 1483 1121 1484 1125
rect 1478 1120 1484 1121
rect 1542 1125 1548 1126
rect 1542 1121 1543 1125
rect 1547 1121 1548 1125
rect 1542 1120 1548 1121
rect 1560 1120 1562 1158
rect 1582 1155 1583 1159
rect 1587 1155 1588 1159
rect 1582 1154 1588 1155
rect 1584 1151 1586 1154
rect 1583 1150 1587 1151
rect 1583 1145 1587 1146
rect 1584 1142 1586 1145
rect 1582 1141 1588 1142
rect 1582 1137 1583 1141
rect 1587 1137 1588 1141
rect 1582 1136 1588 1137
rect 1582 1124 1588 1125
rect 1582 1120 1583 1124
rect 1587 1120 1588 1124
rect 1480 1115 1482 1120
rect 1518 1119 1524 1120
rect 1518 1115 1519 1119
rect 1523 1115 1524 1119
rect 1544 1115 1546 1120
rect 1558 1119 1564 1120
rect 1582 1119 1588 1120
rect 1558 1115 1559 1119
rect 1563 1115 1564 1119
rect 1584 1115 1586 1119
rect 1439 1114 1443 1115
rect 1439 1109 1443 1110
rect 1479 1114 1483 1115
rect 1479 1109 1483 1110
rect 1503 1114 1507 1115
rect 1518 1114 1524 1115
rect 1543 1114 1547 1115
rect 1558 1114 1564 1115
rect 1583 1114 1587 1115
rect 1503 1109 1507 1110
rect 1440 1104 1442 1109
rect 1504 1104 1506 1109
rect 1438 1103 1444 1104
rect 1438 1099 1439 1103
rect 1443 1099 1444 1103
rect 1438 1098 1444 1099
rect 1502 1103 1508 1104
rect 1502 1099 1503 1103
rect 1507 1099 1508 1103
rect 1502 1098 1508 1099
rect 1520 1092 1522 1114
rect 1543 1109 1547 1110
rect 1583 1109 1587 1110
rect 1544 1104 1546 1109
rect 1584 1105 1586 1109
rect 1582 1104 1588 1105
rect 1542 1103 1548 1104
rect 1542 1099 1543 1103
rect 1547 1099 1548 1103
rect 1582 1100 1583 1104
rect 1587 1100 1588 1104
rect 1582 1099 1588 1100
rect 1542 1098 1548 1099
rect 1518 1091 1524 1092
rect 1518 1087 1519 1091
rect 1523 1087 1524 1091
rect 1518 1086 1524 1087
rect 1558 1091 1564 1092
rect 1558 1087 1559 1091
rect 1563 1087 1564 1091
rect 1558 1086 1564 1087
rect 1582 1087 1588 1088
rect 1438 1085 1444 1086
rect 1438 1081 1439 1085
rect 1443 1081 1444 1085
rect 1438 1080 1444 1081
rect 1502 1085 1508 1086
rect 1502 1081 1503 1085
rect 1507 1081 1508 1085
rect 1502 1080 1508 1081
rect 1542 1085 1548 1086
rect 1542 1081 1543 1085
rect 1547 1081 1548 1085
rect 1542 1080 1548 1081
rect 1418 1079 1424 1080
rect 1418 1075 1419 1079
rect 1423 1075 1424 1079
rect 1418 1074 1424 1075
rect 1440 1071 1442 1080
rect 1504 1071 1506 1080
rect 1544 1071 1546 1080
rect 1439 1070 1443 1071
rect 1439 1065 1443 1066
rect 1447 1070 1451 1071
rect 1447 1064 1451 1066
rect 1503 1070 1507 1071
rect 1503 1064 1507 1066
rect 1543 1070 1547 1071
rect 1543 1064 1547 1066
rect 1446 1063 1452 1064
rect 1446 1059 1447 1063
rect 1451 1059 1452 1063
rect 1446 1058 1452 1059
rect 1502 1063 1508 1064
rect 1502 1059 1503 1063
rect 1507 1059 1508 1063
rect 1502 1058 1508 1059
rect 1542 1063 1548 1064
rect 1542 1059 1543 1063
rect 1547 1059 1548 1063
rect 1542 1058 1548 1059
rect 1410 1055 1416 1056
rect 1410 1051 1411 1055
rect 1415 1051 1416 1055
rect 1410 1050 1416 1051
rect 1530 1055 1536 1056
rect 1530 1051 1531 1055
rect 1535 1051 1536 1055
rect 1530 1050 1536 1051
rect 1390 1045 1396 1046
rect 1390 1041 1391 1045
rect 1395 1041 1396 1045
rect 1390 1040 1396 1041
rect 1446 1045 1452 1046
rect 1446 1041 1447 1045
rect 1451 1041 1452 1045
rect 1446 1040 1452 1041
rect 1502 1045 1508 1046
rect 1502 1041 1503 1045
rect 1507 1041 1508 1045
rect 1502 1040 1508 1041
rect 1216 1031 1218 1040
rect 1280 1031 1282 1040
rect 1336 1031 1338 1040
rect 1382 1039 1388 1040
rect 1382 1035 1383 1039
rect 1387 1035 1388 1039
rect 1382 1034 1388 1035
rect 1392 1031 1394 1040
rect 1448 1031 1450 1040
rect 1474 1039 1480 1040
rect 1474 1035 1475 1039
rect 1479 1035 1480 1039
rect 1474 1034 1480 1035
rect 1215 1030 1219 1031
rect 1215 1025 1219 1026
rect 1239 1030 1243 1031
rect 1239 1025 1243 1026
rect 1279 1030 1283 1031
rect 1279 1025 1283 1026
rect 1303 1030 1307 1031
rect 1303 1025 1307 1026
rect 1335 1030 1339 1031
rect 1335 1025 1339 1026
rect 1359 1030 1363 1031
rect 1359 1025 1363 1026
rect 1391 1030 1395 1031
rect 1391 1025 1395 1026
rect 1407 1030 1411 1031
rect 1407 1025 1411 1026
rect 1447 1030 1451 1031
rect 1447 1025 1451 1026
rect 1455 1030 1459 1031
rect 1455 1025 1459 1026
rect 1186 1023 1192 1024
rect 978 1018 984 1019
rect 1006 1019 1012 1020
rect 926 1014 932 1015
rect 726 1007 732 1008
rect 726 1006 727 1007
rect 720 1004 727 1006
rect 726 1003 727 1004
rect 731 1003 732 1007
rect 726 1002 732 1003
rect 790 1007 796 1008
rect 790 1003 791 1007
rect 795 1003 796 1007
rect 790 1002 796 1003
rect 662 1001 668 1002
rect 662 997 663 1001
rect 667 997 668 1001
rect 662 996 668 997
rect 710 1001 716 1002
rect 710 997 711 1001
rect 715 997 716 1001
rect 710 996 716 997
rect 774 1001 780 1002
rect 774 997 775 1001
rect 779 997 780 1001
rect 774 996 780 997
rect 626 987 632 988
rect 664 987 666 996
rect 712 987 714 996
rect 776 987 778 996
rect 111 986 115 987
rect 111 981 115 982
rect 159 986 163 987
rect 112 978 114 981
rect 159 980 163 982
rect 199 986 203 987
rect 199 980 203 982
rect 255 986 259 987
rect 255 980 259 982
rect 311 986 315 987
rect 311 980 315 982
rect 375 986 379 987
rect 375 980 379 982
rect 439 986 443 987
rect 439 980 443 982
rect 503 986 507 987
rect 503 980 507 982
rect 511 986 515 987
rect 511 981 515 982
rect 543 986 547 987
rect 543 981 547 982
rect 559 986 563 987
rect 559 980 563 982
rect 575 986 579 987
rect 575 981 579 982
rect 615 986 619 987
rect 626 983 627 987
rect 631 983 632 987
rect 626 982 632 983
rect 663 986 667 987
rect 615 980 619 982
rect 663 980 667 982
rect 703 986 707 987
rect 703 980 707 982
rect 711 986 715 987
rect 711 981 715 982
rect 735 986 739 987
rect 735 980 739 982
rect 775 986 779 987
rect 775 980 779 982
rect 158 979 164 980
rect 110 977 116 978
rect 110 973 111 977
rect 115 973 116 977
rect 158 975 159 979
rect 163 975 164 979
rect 158 974 164 975
rect 198 979 204 980
rect 198 975 199 979
rect 203 975 204 979
rect 198 974 204 975
rect 254 979 260 980
rect 254 975 255 979
rect 259 975 260 979
rect 254 974 260 975
rect 310 979 316 980
rect 310 975 311 979
rect 315 975 316 979
rect 310 974 316 975
rect 374 979 380 980
rect 374 975 375 979
rect 379 975 380 979
rect 374 974 380 975
rect 438 979 444 980
rect 438 975 439 979
rect 443 975 444 979
rect 438 974 444 975
rect 502 979 508 980
rect 502 975 503 979
rect 507 975 508 979
rect 502 974 508 975
rect 558 979 564 980
rect 558 975 559 979
rect 563 975 564 979
rect 558 974 564 975
rect 614 979 620 980
rect 614 975 615 979
rect 619 975 620 979
rect 614 974 620 975
rect 662 979 668 980
rect 662 975 663 979
rect 667 975 668 979
rect 662 974 668 975
rect 702 979 708 980
rect 702 975 703 979
rect 707 975 708 979
rect 702 974 708 975
rect 734 979 740 980
rect 734 975 735 979
rect 739 975 740 979
rect 734 974 740 975
rect 774 979 780 980
rect 774 975 775 979
rect 779 975 780 979
rect 774 974 780 975
rect 110 972 116 973
rect 523 972 527 973
rect 587 972 591 973
rect 170 971 176 972
rect 170 967 171 971
rect 175 967 176 971
rect 523 967 527 968
rect 586 967 587 972
rect 591 967 592 972
rect 170 966 176 967
rect 158 961 164 962
rect 110 960 116 961
rect 110 956 111 960
rect 115 956 116 960
rect 158 957 159 961
rect 163 957 164 961
rect 158 956 164 957
rect 110 955 116 956
rect 112 951 114 955
rect 160 951 162 956
rect 111 950 115 951
rect 111 945 115 946
rect 151 950 155 951
rect 151 945 155 946
rect 159 950 163 951
rect 159 945 163 946
rect 112 941 114 945
rect 110 940 116 941
rect 152 940 154 945
rect 172 944 174 966
rect 198 961 204 962
rect 198 957 199 961
rect 203 957 204 961
rect 198 956 204 957
rect 254 961 260 962
rect 254 957 255 961
rect 259 957 260 961
rect 254 956 260 957
rect 310 961 316 962
rect 310 957 311 961
rect 315 957 316 961
rect 310 956 316 957
rect 374 961 380 962
rect 374 957 375 961
rect 379 957 380 961
rect 374 956 380 957
rect 438 961 444 962
rect 438 957 439 961
rect 443 957 444 961
rect 438 956 444 957
rect 502 961 508 962
rect 502 957 503 961
rect 507 957 508 961
rect 502 956 508 957
rect 524 956 526 967
rect 586 966 592 967
rect 558 961 564 962
rect 558 957 559 961
rect 563 957 564 961
rect 558 956 564 957
rect 614 961 620 962
rect 614 957 615 961
rect 619 957 620 961
rect 614 956 620 957
rect 662 961 668 962
rect 662 957 663 961
rect 667 957 668 961
rect 662 956 668 957
rect 702 961 708 962
rect 702 957 703 961
rect 707 957 708 961
rect 702 956 708 957
rect 734 961 740 962
rect 734 957 735 961
rect 739 957 740 961
rect 734 956 740 957
rect 774 961 780 962
rect 774 957 775 961
rect 779 957 780 961
rect 774 956 780 957
rect 792 956 794 1002
rect 846 1001 852 1002
rect 846 997 847 1001
rect 851 997 852 1001
rect 846 996 852 997
rect 926 1001 932 1002
rect 926 997 927 1001
rect 931 997 932 1001
rect 926 996 932 997
rect 980 996 982 1018
rect 1006 1015 1007 1019
rect 1011 1015 1012 1019
rect 1006 1014 1012 1015
rect 1086 1019 1092 1020
rect 1086 1015 1087 1019
rect 1091 1015 1092 1019
rect 1086 1014 1092 1015
rect 1166 1019 1172 1020
rect 1166 1015 1167 1019
rect 1171 1015 1172 1019
rect 1186 1019 1187 1023
rect 1191 1019 1192 1023
rect 1240 1020 1242 1025
rect 1304 1020 1306 1025
rect 1360 1020 1362 1025
rect 1408 1020 1410 1025
rect 1456 1020 1458 1025
rect 1186 1018 1192 1019
rect 1238 1019 1244 1020
rect 1166 1014 1172 1015
rect 1238 1015 1239 1019
rect 1243 1015 1244 1019
rect 1238 1014 1244 1015
rect 1302 1019 1308 1020
rect 1302 1015 1303 1019
rect 1307 1015 1308 1019
rect 1302 1014 1308 1015
rect 1358 1019 1364 1020
rect 1358 1015 1359 1019
rect 1363 1015 1364 1019
rect 1358 1014 1364 1015
rect 1406 1019 1412 1020
rect 1406 1015 1407 1019
rect 1411 1015 1412 1019
rect 1406 1014 1412 1015
rect 1454 1019 1460 1020
rect 1454 1015 1455 1019
rect 1459 1015 1460 1019
rect 1454 1014 1460 1015
rect 1476 1008 1478 1034
rect 1504 1031 1506 1040
rect 1503 1030 1507 1031
rect 1503 1025 1507 1026
rect 1511 1030 1515 1031
rect 1511 1025 1515 1026
rect 1512 1020 1514 1025
rect 1532 1024 1534 1050
rect 1542 1045 1548 1046
rect 1542 1041 1543 1045
rect 1547 1041 1548 1045
rect 1542 1040 1548 1041
rect 1560 1040 1562 1086
rect 1582 1083 1583 1087
rect 1587 1083 1588 1087
rect 1582 1082 1588 1083
rect 1584 1071 1586 1082
rect 1583 1070 1587 1071
rect 1583 1065 1587 1066
rect 1584 1062 1586 1065
rect 1582 1061 1588 1062
rect 1582 1057 1583 1061
rect 1587 1057 1588 1061
rect 1582 1056 1588 1057
rect 1582 1044 1588 1045
rect 1582 1040 1583 1044
rect 1587 1040 1588 1044
rect 1544 1031 1546 1040
rect 1558 1039 1564 1040
rect 1582 1039 1588 1040
rect 1558 1035 1559 1039
rect 1563 1035 1564 1039
rect 1558 1034 1564 1035
rect 1584 1031 1586 1039
rect 1543 1030 1547 1031
rect 1543 1025 1547 1026
rect 1583 1030 1587 1031
rect 1583 1025 1587 1026
rect 1530 1023 1536 1024
rect 1510 1019 1516 1020
rect 1510 1015 1511 1019
rect 1515 1015 1516 1019
rect 1530 1019 1531 1023
rect 1535 1019 1536 1023
rect 1544 1020 1546 1025
rect 1584 1021 1586 1025
rect 1582 1020 1588 1021
rect 1530 1018 1536 1019
rect 1542 1019 1548 1020
rect 1510 1014 1516 1015
rect 1542 1015 1543 1019
rect 1547 1015 1548 1019
rect 1582 1016 1583 1020
rect 1587 1016 1588 1020
rect 1582 1015 1588 1016
rect 1542 1014 1548 1015
rect 1474 1007 1480 1008
rect 1474 1003 1475 1007
rect 1479 1003 1480 1007
rect 1474 1002 1480 1003
rect 1558 1007 1564 1008
rect 1558 1003 1559 1007
rect 1563 1003 1564 1007
rect 1558 1002 1564 1003
rect 1582 1003 1588 1004
rect 1006 1001 1012 1002
rect 1006 997 1007 1001
rect 1011 997 1012 1001
rect 1006 996 1012 997
rect 1086 1001 1092 1002
rect 1086 997 1087 1001
rect 1091 997 1092 1001
rect 1086 996 1092 997
rect 1166 1001 1172 1002
rect 1166 997 1167 1001
rect 1171 997 1172 1001
rect 1166 996 1172 997
rect 1238 1001 1244 1002
rect 1238 997 1239 1001
rect 1243 997 1244 1001
rect 1238 996 1244 997
rect 1302 1001 1308 1002
rect 1302 997 1303 1001
rect 1307 997 1308 1001
rect 1302 996 1308 997
rect 1358 1001 1364 1002
rect 1358 997 1359 1001
rect 1363 997 1364 1001
rect 1358 996 1364 997
rect 1406 1001 1412 1002
rect 1406 997 1407 1001
rect 1411 997 1412 1001
rect 1406 996 1412 997
rect 1454 1001 1460 1002
rect 1454 997 1455 1001
rect 1459 997 1460 1001
rect 1454 996 1460 997
rect 1510 1001 1516 1002
rect 1510 997 1511 1001
rect 1515 997 1516 1001
rect 1510 996 1516 997
rect 1542 1001 1548 1002
rect 1542 997 1543 1001
rect 1547 997 1548 1001
rect 1542 996 1548 997
rect 822 987 828 988
rect 848 987 850 996
rect 928 987 930 996
rect 978 995 984 996
rect 978 991 979 995
rect 983 991 984 995
rect 978 990 984 991
rect 1008 987 1010 996
rect 1088 987 1090 996
rect 1168 987 1170 996
rect 1240 987 1242 996
rect 1304 987 1306 996
rect 1360 987 1362 996
rect 1408 987 1410 996
rect 1456 987 1458 996
rect 1512 987 1514 996
rect 1544 987 1546 996
rect 822 983 823 987
rect 827 983 828 987
rect 822 982 828 983
rect 831 986 835 987
rect 200 951 202 956
rect 256 951 258 956
rect 312 951 314 956
rect 376 951 378 956
rect 440 951 442 956
rect 450 955 456 956
rect 450 951 451 955
rect 455 951 456 955
rect 504 951 506 956
rect 522 955 528 956
rect 522 951 523 955
rect 527 951 528 955
rect 560 951 562 956
rect 616 951 618 956
rect 664 951 666 956
rect 704 951 706 956
rect 736 951 738 956
rect 776 951 778 956
rect 782 955 788 956
rect 782 951 783 955
rect 787 951 788 955
rect 191 950 195 951
rect 191 945 195 946
rect 199 950 203 951
rect 199 945 203 946
rect 247 950 251 951
rect 247 945 251 946
rect 255 950 259 951
rect 255 945 259 946
rect 303 950 307 951
rect 303 945 307 946
rect 311 950 315 951
rect 311 945 315 946
rect 367 950 371 951
rect 367 945 371 946
rect 375 950 379 951
rect 375 945 379 946
rect 431 950 435 951
rect 431 945 435 946
rect 439 950 443 951
rect 450 950 456 951
rect 495 950 499 951
rect 439 945 443 946
rect 170 943 176 944
rect 110 936 111 940
rect 115 936 116 940
rect 110 935 116 936
rect 150 939 156 940
rect 150 935 151 939
rect 155 935 156 939
rect 170 939 171 943
rect 175 939 176 943
rect 192 940 194 945
rect 248 940 250 945
rect 304 940 306 945
rect 318 943 324 944
rect 170 938 176 939
rect 190 939 196 940
rect 150 934 156 935
rect 190 935 191 939
rect 195 935 196 939
rect 190 934 196 935
rect 246 939 252 940
rect 246 935 247 939
rect 251 935 252 939
rect 246 934 252 935
rect 302 939 308 940
rect 302 935 303 939
rect 307 935 308 939
rect 318 939 319 943
rect 323 939 324 943
rect 368 940 370 945
rect 432 940 434 945
rect 318 938 324 939
rect 366 939 372 940
rect 302 934 308 935
rect 262 927 268 928
rect 110 923 116 924
rect 110 919 111 923
rect 115 919 116 923
rect 262 923 263 927
rect 267 923 268 927
rect 262 922 268 923
rect 110 918 116 919
rect 150 921 156 922
rect 112 911 114 918
rect 150 917 151 921
rect 155 917 156 921
rect 150 916 156 917
rect 190 921 196 922
rect 190 917 191 921
rect 195 917 196 921
rect 190 916 196 917
rect 246 921 252 922
rect 246 917 247 921
rect 251 917 252 921
rect 246 916 252 917
rect 152 911 154 916
rect 192 911 194 916
rect 248 911 250 916
rect 111 910 115 911
rect 111 905 115 906
rect 135 910 139 911
rect 112 902 114 905
rect 135 904 139 906
rect 151 910 155 911
rect 151 905 155 906
rect 167 910 171 911
rect 167 904 171 906
rect 191 910 195 911
rect 191 905 195 906
rect 223 910 227 911
rect 223 904 227 906
rect 247 910 251 911
rect 247 905 251 906
rect 134 903 140 904
rect 110 901 116 902
rect 110 897 111 901
rect 115 897 116 901
rect 134 899 135 903
rect 139 899 140 903
rect 134 898 140 899
rect 166 903 172 904
rect 166 899 167 903
rect 171 899 172 903
rect 166 898 172 899
rect 222 903 228 904
rect 222 899 223 903
rect 227 899 228 903
rect 222 898 228 899
rect 110 896 116 897
rect 150 895 156 896
rect 150 891 151 895
rect 155 891 156 895
rect 150 890 156 891
rect 134 885 140 886
rect 110 884 116 885
rect 110 880 111 884
rect 115 880 116 884
rect 134 881 135 885
rect 139 881 140 885
rect 134 880 140 881
rect 110 879 116 880
rect 112 875 114 879
rect 136 875 138 880
rect 111 874 115 875
rect 111 869 115 870
rect 135 874 139 875
rect 135 869 139 870
rect 112 865 114 869
rect 110 864 116 865
rect 136 864 138 869
rect 152 868 154 890
rect 166 885 172 886
rect 166 881 167 885
rect 171 881 172 885
rect 166 880 172 881
rect 222 885 228 886
rect 222 881 223 885
rect 227 881 228 885
rect 222 880 228 881
rect 264 880 266 922
rect 302 921 308 922
rect 302 917 303 921
rect 307 917 308 921
rect 302 916 308 917
rect 304 911 306 916
rect 279 910 283 911
rect 279 904 283 906
rect 303 910 307 911
rect 303 905 307 906
rect 278 903 284 904
rect 278 899 279 903
rect 283 899 284 903
rect 278 898 284 899
rect 320 896 322 938
rect 366 935 367 939
rect 371 935 372 939
rect 366 934 372 935
rect 430 939 436 940
rect 430 935 431 939
rect 435 935 436 939
rect 430 934 436 935
rect 452 928 454 950
rect 495 945 499 946
rect 503 950 507 951
rect 522 950 528 951
rect 559 950 563 951
rect 503 945 507 946
rect 559 945 563 946
rect 615 950 619 951
rect 615 945 619 946
rect 663 950 667 951
rect 663 945 667 946
rect 671 950 675 951
rect 671 945 675 946
rect 703 950 707 951
rect 703 945 707 946
rect 719 950 723 951
rect 719 945 723 946
rect 735 950 739 951
rect 735 945 739 946
rect 767 950 771 951
rect 767 945 771 946
rect 775 950 779 951
rect 782 950 788 951
rect 790 955 796 956
rect 790 951 791 955
rect 795 951 796 955
rect 790 950 796 951
rect 815 950 819 951
rect 775 945 779 946
rect 496 940 498 945
rect 550 943 556 944
rect 494 939 500 940
rect 494 935 495 939
rect 499 935 500 939
rect 550 939 551 943
rect 555 939 556 943
rect 560 940 562 945
rect 616 940 618 945
rect 672 940 674 945
rect 720 940 722 945
rect 768 940 770 945
rect 550 938 556 939
rect 558 939 564 940
rect 494 934 500 935
rect 450 927 456 928
rect 450 923 451 927
rect 455 923 456 927
rect 450 922 456 923
rect 366 921 372 922
rect 366 917 367 921
rect 371 917 372 921
rect 366 916 372 917
rect 430 921 436 922
rect 430 917 431 921
rect 435 917 436 921
rect 430 916 436 917
rect 494 921 500 922
rect 494 917 495 921
rect 499 917 500 921
rect 494 916 500 917
rect 368 911 370 916
rect 432 911 434 916
rect 496 911 498 916
rect 552 912 554 938
rect 558 935 559 939
rect 563 935 564 939
rect 558 934 564 935
rect 614 939 620 940
rect 614 935 615 939
rect 619 935 620 939
rect 614 934 620 935
rect 670 939 676 940
rect 670 935 671 939
rect 675 935 676 939
rect 670 934 676 935
rect 718 939 724 940
rect 718 935 719 939
rect 723 935 724 939
rect 718 934 724 935
rect 766 939 772 940
rect 766 935 767 939
rect 771 935 772 939
rect 766 934 772 935
rect 784 928 786 950
rect 824 948 826 982
rect 831 980 835 982
rect 847 986 851 987
rect 847 981 851 982
rect 895 986 899 987
rect 895 980 899 982
rect 927 986 931 987
rect 927 981 931 982
rect 967 986 971 987
rect 967 980 971 982
rect 1007 986 1011 987
rect 1007 981 1011 982
rect 1047 986 1051 987
rect 1047 980 1051 982
rect 1087 986 1091 987
rect 1087 981 1091 982
rect 1127 986 1131 987
rect 1127 980 1131 982
rect 1167 986 1171 987
rect 1167 981 1171 982
rect 1199 986 1203 987
rect 1199 980 1203 982
rect 1239 986 1243 987
rect 1239 981 1243 982
rect 1271 986 1275 987
rect 1271 980 1275 982
rect 1303 986 1307 987
rect 1303 981 1307 982
rect 1343 986 1347 987
rect 1343 980 1347 982
rect 1359 986 1363 987
rect 1359 981 1363 982
rect 1407 986 1411 987
rect 1407 981 1411 982
rect 1415 986 1419 987
rect 1415 980 1419 982
rect 1455 986 1459 987
rect 1455 981 1459 982
rect 1487 986 1491 987
rect 1487 980 1491 982
rect 1511 986 1515 987
rect 1511 981 1515 982
rect 1543 986 1547 987
rect 1543 980 1547 982
rect 830 979 836 980
rect 830 975 831 979
rect 835 975 836 979
rect 830 974 836 975
rect 894 979 900 980
rect 894 975 895 979
rect 899 975 900 979
rect 894 974 900 975
rect 966 979 972 980
rect 966 975 967 979
rect 971 975 972 979
rect 966 974 972 975
rect 1046 979 1052 980
rect 1046 975 1047 979
rect 1051 975 1052 979
rect 1046 974 1052 975
rect 1126 979 1132 980
rect 1126 975 1127 979
rect 1131 975 1132 979
rect 1126 974 1132 975
rect 1198 979 1204 980
rect 1198 975 1199 979
rect 1203 975 1204 979
rect 1198 974 1204 975
rect 1270 979 1276 980
rect 1270 975 1271 979
rect 1275 975 1276 979
rect 1270 974 1276 975
rect 1342 979 1348 980
rect 1342 975 1343 979
rect 1347 975 1348 979
rect 1342 974 1348 975
rect 1414 979 1420 980
rect 1414 975 1415 979
rect 1419 975 1420 979
rect 1414 974 1420 975
rect 1486 979 1492 980
rect 1486 975 1487 979
rect 1491 975 1492 979
rect 1486 974 1492 975
rect 1542 979 1548 980
rect 1542 975 1543 979
rect 1547 975 1548 979
rect 1542 974 1548 975
rect 1218 971 1224 972
rect 1218 967 1219 971
rect 1223 967 1224 971
rect 1218 966 1224 967
rect 830 961 836 962
rect 830 957 831 961
rect 835 957 836 961
rect 830 956 836 957
rect 894 961 900 962
rect 894 957 895 961
rect 899 957 900 961
rect 894 956 900 957
rect 966 961 972 962
rect 966 957 967 961
rect 971 957 972 961
rect 966 956 972 957
rect 1046 961 1052 962
rect 1046 957 1047 961
rect 1051 957 1052 961
rect 1046 956 1052 957
rect 1126 961 1132 962
rect 1126 957 1127 961
rect 1131 957 1132 961
rect 1126 956 1132 957
rect 1198 961 1204 962
rect 1198 957 1199 961
rect 1203 957 1204 961
rect 1198 956 1204 957
rect 832 951 834 956
rect 896 951 898 956
rect 968 951 970 956
rect 1048 951 1050 956
rect 1128 951 1130 956
rect 1200 951 1202 956
rect 831 950 835 951
rect 815 945 819 946
rect 822 947 828 948
rect 816 940 818 945
rect 822 943 823 947
rect 827 943 828 947
rect 831 945 835 946
rect 871 950 875 951
rect 871 945 875 946
rect 895 950 899 951
rect 895 945 899 946
rect 935 950 939 951
rect 935 945 939 946
rect 967 950 971 951
rect 967 945 971 946
rect 1007 950 1011 951
rect 1007 945 1011 946
rect 1047 950 1051 951
rect 1047 945 1051 946
rect 1079 950 1083 951
rect 1079 945 1083 946
rect 1127 950 1131 951
rect 1127 945 1131 946
rect 1143 950 1147 951
rect 1143 945 1147 946
rect 1199 950 1203 951
rect 1199 945 1203 946
rect 1207 950 1211 951
rect 1207 945 1211 946
rect 822 942 828 943
rect 872 940 874 945
rect 936 940 938 945
rect 1008 940 1010 945
rect 1080 940 1082 945
rect 1144 940 1146 945
rect 1208 940 1210 945
rect 1220 944 1222 966
rect 1270 961 1276 962
rect 1270 957 1271 961
rect 1275 957 1276 961
rect 1270 956 1276 957
rect 1342 961 1348 962
rect 1342 957 1343 961
rect 1347 957 1348 961
rect 1342 956 1348 957
rect 1414 961 1420 962
rect 1414 957 1415 961
rect 1419 957 1420 961
rect 1414 956 1420 957
rect 1486 961 1492 962
rect 1486 957 1487 961
rect 1491 957 1492 961
rect 1486 956 1492 957
rect 1542 961 1548 962
rect 1542 957 1543 961
rect 1547 957 1548 961
rect 1542 956 1548 957
rect 1560 956 1562 1002
rect 1582 999 1583 1003
rect 1587 999 1588 1003
rect 1582 998 1588 999
rect 1584 987 1586 998
rect 1583 986 1587 987
rect 1583 981 1587 982
rect 1584 978 1586 981
rect 1582 977 1588 978
rect 1582 973 1583 977
rect 1587 973 1588 977
rect 1582 972 1588 973
rect 1582 960 1588 961
rect 1582 956 1583 960
rect 1587 956 1588 960
rect 1272 951 1274 956
rect 1344 951 1346 956
rect 1416 951 1418 956
rect 1488 951 1490 956
rect 1498 955 1504 956
rect 1498 951 1499 955
rect 1503 951 1504 955
rect 1544 951 1546 956
rect 1558 955 1564 956
rect 1582 955 1588 956
rect 1558 951 1559 955
rect 1563 951 1564 955
rect 1584 951 1586 955
rect 1271 950 1275 951
rect 1271 945 1275 946
rect 1327 950 1331 951
rect 1327 945 1331 946
rect 1343 950 1347 951
rect 1343 945 1347 946
rect 1375 950 1379 951
rect 1375 945 1379 946
rect 1415 950 1419 951
rect 1415 945 1419 946
rect 1423 950 1427 951
rect 1423 945 1427 946
rect 1471 950 1475 951
rect 1471 945 1475 946
rect 1487 950 1491 951
rect 1498 950 1504 951
rect 1511 950 1515 951
rect 1487 945 1491 946
rect 1218 943 1224 944
rect 814 939 820 940
rect 814 935 815 939
rect 819 935 820 939
rect 814 934 820 935
rect 870 939 876 940
rect 870 935 871 939
rect 875 935 876 939
rect 870 934 876 935
rect 934 939 940 940
rect 934 935 935 939
rect 939 935 940 939
rect 934 934 940 935
rect 1006 939 1012 940
rect 1006 935 1007 939
rect 1011 935 1012 939
rect 1006 934 1012 935
rect 1078 939 1084 940
rect 1078 935 1079 939
rect 1083 935 1084 939
rect 1078 934 1084 935
rect 1142 939 1148 940
rect 1142 935 1143 939
rect 1147 935 1148 939
rect 1142 934 1148 935
rect 1206 939 1212 940
rect 1206 935 1207 939
rect 1211 935 1212 939
rect 1218 939 1219 943
rect 1223 939 1224 943
rect 1272 940 1274 945
rect 1328 940 1330 945
rect 1376 940 1378 945
rect 1424 940 1426 945
rect 1472 940 1474 945
rect 1218 938 1224 939
rect 1270 939 1276 940
rect 1206 934 1212 935
rect 1270 935 1271 939
rect 1275 935 1276 939
rect 1270 934 1276 935
rect 1326 939 1332 940
rect 1326 935 1327 939
rect 1331 935 1332 939
rect 1326 934 1332 935
rect 1374 939 1380 940
rect 1374 935 1375 939
rect 1379 935 1380 939
rect 1374 934 1380 935
rect 1422 939 1428 940
rect 1422 935 1423 939
rect 1427 935 1428 939
rect 1422 934 1428 935
rect 1470 939 1476 940
rect 1470 935 1471 939
rect 1475 935 1476 939
rect 1470 934 1476 935
rect 1500 928 1502 950
rect 1511 945 1515 946
rect 1543 950 1547 951
rect 1558 950 1564 951
rect 1583 950 1587 951
rect 1543 945 1547 946
rect 1583 945 1587 946
rect 1512 940 1514 945
rect 1544 940 1546 945
rect 1584 941 1586 945
rect 1582 940 1588 941
rect 1510 939 1516 940
rect 1510 935 1511 939
rect 1515 935 1516 939
rect 1510 934 1516 935
rect 1542 939 1548 940
rect 1542 935 1543 939
rect 1547 935 1548 939
rect 1582 936 1583 940
rect 1587 936 1588 940
rect 1582 935 1588 936
rect 1542 934 1548 935
rect 782 927 788 928
rect 782 923 783 927
rect 787 923 788 927
rect 782 922 788 923
rect 1366 927 1372 928
rect 1366 923 1367 927
rect 1371 923 1372 927
rect 1366 922 1372 923
rect 1498 927 1504 928
rect 1498 923 1499 927
rect 1503 923 1504 927
rect 1498 922 1504 923
rect 1582 923 1588 924
rect 558 921 564 922
rect 558 917 559 921
rect 563 917 564 921
rect 558 916 564 917
rect 614 921 620 922
rect 614 917 615 921
rect 619 917 620 921
rect 614 916 620 917
rect 670 921 676 922
rect 670 917 671 921
rect 675 917 676 921
rect 670 916 676 917
rect 718 921 724 922
rect 718 917 719 921
rect 723 917 724 921
rect 718 916 724 917
rect 766 921 772 922
rect 766 917 767 921
rect 771 917 772 921
rect 766 916 772 917
rect 814 921 820 922
rect 814 917 815 921
rect 819 917 820 921
rect 814 916 820 917
rect 870 921 876 922
rect 870 917 871 921
rect 875 917 876 921
rect 870 916 876 917
rect 934 921 940 922
rect 934 917 935 921
rect 939 917 940 921
rect 934 916 940 917
rect 1006 921 1012 922
rect 1006 917 1007 921
rect 1011 917 1012 921
rect 1006 916 1012 917
rect 1078 921 1084 922
rect 1078 917 1079 921
rect 1083 917 1084 921
rect 1078 916 1084 917
rect 1142 921 1148 922
rect 1142 917 1143 921
rect 1147 917 1148 921
rect 1142 916 1148 917
rect 1206 921 1212 922
rect 1206 917 1207 921
rect 1211 917 1212 921
rect 1206 916 1212 917
rect 1270 921 1276 922
rect 1270 917 1271 921
rect 1275 917 1276 921
rect 1270 916 1276 917
rect 1326 921 1332 922
rect 1326 917 1327 921
rect 1331 917 1332 921
rect 1326 916 1332 917
rect 550 911 556 912
rect 560 911 562 916
rect 616 911 618 916
rect 672 911 674 916
rect 720 911 722 916
rect 768 911 770 916
rect 816 911 818 916
rect 872 911 874 916
rect 936 911 938 916
rect 1008 911 1010 916
rect 1080 911 1082 916
rect 1144 911 1146 916
rect 1208 911 1210 916
rect 1272 911 1274 916
rect 1328 911 1330 916
rect 335 910 339 911
rect 335 904 339 906
rect 367 910 371 911
rect 367 905 371 906
rect 391 910 395 911
rect 391 904 395 906
rect 431 910 435 911
rect 431 905 435 906
rect 447 910 451 911
rect 447 904 451 906
rect 495 910 499 911
rect 495 905 499 906
rect 503 910 507 911
rect 550 907 551 911
rect 555 907 556 911
rect 550 906 556 907
rect 559 910 563 911
rect 503 904 507 906
rect 559 904 563 906
rect 615 910 619 911
rect 615 905 619 906
rect 623 910 627 911
rect 623 904 627 906
rect 671 910 675 911
rect 671 905 675 906
rect 695 910 699 911
rect 695 904 699 906
rect 719 910 723 911
rect 719 905 723 906
rect 759 910 763 911
rect 759 904 763 906
rect 767 910 771 911
rect 767 905 771 906
rect 815 910 819 911
rect 815 905 819 906
rect 823 910 827 911
rect 823 904 827 906
rect 871 910 875 911
rect 871 905 875 906
rect 887 910 891 911
rect 887 904 891 906
rect 935 910 939 911
rect 935 905 939 906
rect 951 910 955 911
rect 951 904 955 906
rect 1007 910 1011 911
rect 1007 905 1011 906
rect 1015 910 1019 911
rect 1015 904 1019 906
rect 1079 910 1083 911
rect 1079 904 1083 906
rect 1135 910 1139 911
rect 1135 904 1139 906
rect 1143 910 1147 911
rect 1143 905 1147 906
rect 1191 910 1195 911
rect 1191 904 1195 906
rect 1207 910 1211 911
rect 1207 905 1211 906
rect 1247 910 1251 911
rect 1247 904 1251 906
rect 1271 910 1275 911
rect 1271 905 1275 906
rect 1303 910 1307 911
rect 1303 904 1307 906
rect 1327 910 1331 911
rect 1327 905 1331 906
rect 1359 910 1363 911
rect 1359 904 1363 906
rect 334 903 340 904
rect 334 899 335 903
rect 339 899 340 903
rect 334 898 340 899
rect 390 903 396 904
rect 390 899 391 903
rect 395 899 396 903
rect 390 898 396 899
rect 446 903 452 904
rect 446 899 447 903
rect 451 899 452 903
rect 446 898 452 899
rect 502 903 508 904
rect 502 899 503 903
rect 507 899 508 903
rect 502 898 508 899
rect 558 903 564 904
rect 558 899 559 903
rect 563 899 564 903
rect 558 898 564 899
rect 622 903 628 904
rect 622 899 623 903
rect 627 899 628 903
rect 622 898 628 899
rect 694 903 700 904
rect 694 899 695 903
rect 699 899 700 903
rect 694 898 700 899
rect 758 903 764 904
rect 758 899 759 903
rect 763 899 764 903
rect 758 898 764 899
rect 822 903 828 904
rect 822 899 823 903
rect 827 899 828 903
rect 822 898 828 899
rect 886 903 892 904
rect 886 899 887 903
rect 891 899 892 903
rect 886 898 892 899
rect 950 903 956 904
rect 950 899 951 903
rect 955 899 956 903
rect 950 898 956 899
rect 1014 903 1020 904
rect 1014 899 1015 903
rect 1019 899 1020 903
rect 1014 898 1020 899
rect 1078 903 1084 904
rect 1078 899 1079 903
rect 1083 899 1084 903
rect 1078 898 1084 899
rect 1134 903 1140 904
rect 1134 899 1135 903
rect 1139 899 1140 903
rect 1134 898 1140 899
rect 1190 903 1196 904
rect 1190 899 1191 903
rect 1195 899 1196 903
rect 1190 898 1196 899
rect 1246 903 1252 904
rect 1246 899 1247 903
rect 1251 899 1252 903
rect 1246 898 1252 899
rect 1302 903 1308 904
rect 1302 899 1303 903
rect 1307 899 1308 903
rect 1302 898 1308 899
rect 1358 903 1364 904
rect 1358 899 1359 903
rect 1363 899 1364 903
rect 1358 898 1364 899
rect 318 895 324 896
rect 318 891 319 895
rect 323 891 324 895
rect 318 890 324 891
rect 1278 895 1284 896
rect 1278 891 1279 895
rect 1283 891 1284 895
rect 1278 890 1284 891
rect 1286 895 1292 896
rect 1286 891 1287 895
rect 1291 891 1292 895
rect 1286 890 1292 891
rect 278 885 284 886
rect 278 881 279 885
rect 283 881 284 885
rect 278 880 284 881
rect 334 885 340 886
rect 334 881 335 885
rect 339 881 340 885
rect 334 880 340 881
rect 390 885 396 886
rect 390 881 391 885
rect 395 881 396 885
rect 390 880 396 881
rect 446 885 452 886
rect 446 881 447 885
rect 451 881 452 885
rect 446 880 452 881
rect 502 885 508 886
rect 502 881 503 885
rect 507 881 508 885
rect 502 880 508 881
rect 558 885 564 886
rect 558 881 559 885
rect 563 881 564 885
rect 558 880 564 881
rect 622 885 628 886
rect 622 881 623 885
rect 627 881 628 885
rect 622 880 628 881
rect 694 885 700 886
rect 694 881 695 885
rect 699 881 700 885
rect 694 880 700 881
rect 758 885 764 886
rect 758 881 759 885
rect 763 881 764 885
rect 758 880 764 881
rect 822 885 828 886
rect 822 881 823 885
rect 827 881 828 885
rect 822 880 828 881
rect 886 885 892 886
rect 886 881 887 885
rect 891 881 892 885
rect 886 880 892 881
rect 950 885 956 886
rect 950 881 951 885
rect 955 881 956 885
rect 950 880 956 881
rect 1014 885 1020 886
rect 1014 881 1015 885
rect 1019 881 1020 885
rect 1014 880 1020 881
rect 1078 885 1084 886
rect 1078 881 1079 885
rect 1083 881 1084 885
rect 1078 880 1084 881
rect 1134 885 1140 886
rect 1134 881 1135 885
rect 1139 881 1140 885
rect 1134 880 1140 881
rect 1190 885 1196 886
rect 1190 881 1191 885
rect 1195 881 1196 885
rect 1190 880 1196 881
rect 1246 885 1252 886
rect 1246 881 1247 885
rect 1251 881 1252 885
rect 1246 880 1252 881
rect 168 875 170 880
rect 224 875 226 880
rect 262 879 268 880
rect 262 875 263 879
rect 267 875 268 879
rect 280 875 282 880
rect 336 875 338 880
rect 392 875 394 880
rect 448 875 450 880
rect 482 879 488 880
rect 482 875 483 879
rect 487 875 488 879
rect 504 875 506 880
rect 560 875 562 880
rect 624 875 626 880
rect 696 875 698 880
rect 760 875 762 880
rect 824 875 826 880
rect 888 875 890 880
rect 952 875 954 880
rect 1016 875 1018 880
rect 1080 875 1082 880
rect 1136 875 1138 880
rect 1192 875 1194 880
rect 1248 875 1250 880
rect 167 874 171 875
rect 167 869 171 870
rect 207 874 211 875
rect 207 869 211 870
rect 223 874 227 875
rect 223 869 227 870
rect 255 874 259 875
rect 262 874 268 875
rect 279 874 283 875
rect 255 869 259 870
rect 279 869 283 870
rect 303 874 307 875
rect 303 869 307 870
rect 335 874 339 875
rect 335 869 339 870
rect 343 874 347 875
rect 343 869 347 870
rect 383 874 387 875
rect 383 869 387 870
rect 391 874 395 875
rect 391 869 395 870
rect 439 874 443 875
rect 439 869 443 870
rect 447 874 451 875
rect 482 874 488 875
rect 503 874 507 875
rect 447 869 451 870
rect 150 867 156 868
rect 110 860 111 864
rect 115 860 116 864
rect 110 859 116 860
rect 134 863 140 864
rect 134 859 135 863
rect 139 859 140 863
rect 150 863 151 867
rect 155 863 156 867
rect 168 864 170 869
rect 208 864 210 869
rect 256 864 258 869
rect 266 867 272 868
rect 150 862 156 863
rect 166 863 172 864
rect 134 858 140 859
rect 166 859 167 863
rect 171 859 172 863
rect 166 858 172 859
rect 206 863 212 864
rect 206 859 207 863
rect 211 859 212 863
rect 206 858 212 859
rect 254 863 260 864
rect 254 859 255 863
rect 259 859 260 863
rect 266 863 267 867
rect 271 863 272 867
rect 304 864 306 869
rect 344 864 346 869
rect 384 864 386 869
rect 440 864 442 869
rect 266 862 272 863
rect 302 863 308 864
rect 254 858 260 859
rect 222 851 228 852
rect 110 847 116 848
rect 110 843 111 847
rect 115 843 116 847
rect 222 847 223 851
rect 227 847 228 851
rect 222 846 228 847
rect 110 842 116 843
rect 134 845 140 846
rect 112 835 114 842
rect 134 841 135 845
rect 139 841 140 845
rect 134 840 140 841
rect 166 845 172 846
rect 166 841 167 845
rect 171 841 172 845
rect 166 840 172 841
rect 206 845 212 846
rect 206 841 207 845
rect 211 841 212 845
rect 224 843 226 846
rect 206 840 212 841
rect 216 841 226 843
rect 254 845 260 846
rect 254 841 255 845
rect 259 841 260 845
rect 136 835 138 840
rect 168 835 170 840
rect 208 835 210 840
rect 111 834 115 835
rect 111 829 115 830
rect 135 834 139 835
rect 112 826 114 829
rect 135 828 139 830
rect 167 834 171 835
rect 167 828 171 830
rect 207 834 211 835
rect 207 829 211 830
rect 134 827 140 828
rect 110 825 116 826
rect 110 821 111 825
rect 115 821 116 825
rect 134 823 135 827
rect 139 823 140 827
rect 134 822 140 823
rect 166 827 172 828
rect 166 823 167 827
rect 171 823 172 827
rect 166 822 172 823
rect 110 820 116 821
rect 150 819 156 820
rect 150 815 151 819
rect 155 815 156 819
rect 150 814 156 815
rect 134 809 140 810
rect 110 808 116 809
rect 110 804 111 808
rect 115 804 116 808
rect 134 805 135 809
rect 139 805 140 809
rect 134 804 140 805
rect 110 803 116 804
rect 112 799 114 803
rect 136 799 138 804
rect 111 798 115 799
rect 111 793 115 794
rect 135 798 139 799
rect 135 793 139 794
rect 112 789 114 793
rect 110 788 116 789
rect 136 788 138 793
rect 152 792 154 814
rect 166 809 172 810
rect 166 805 167 809
rect 171 805 172 809
rect 166 804 172 805
rect 216 804 218 841
rect 254 840 260 841
rect 256 835 258 840
rect 223 834 227 835
rect 223 828 227 830
rect 255 834 259 835
rect 255 829 259 830
rect 222 827 228 828
rect 222 823 223 827
rect 227 823 228 827
rect 222 822 228 823
rect 268 820 270 862
rect 302 859 303 863
rect 307 859 308 863
rect 302 858 308 859
rect 342 863 348 864
rect 342 859 343 863
rect 347 859 348 863
rect 342 858 348 859
rect 382 863 388 864
rect 382 859 383 863
rect 387 859 388 863
rect 382 858 388 859
rect 438 863 444 864
rect 438 859 439 863
rect 443 859 444 863
rect 438 858 444 859
rect 302 845 308 846
rect 302 841 303 845
rect 307 841 308 845
rect 302 840 308 841
rect 342 845 348 846
rect 342 841 343 845
rect 347 841 348 845
rect 342 840 348 841
rect 382 845 388 846
rect 382 841 383 845
rect 387 841 388 845
rect 382 840 388 841
rect 438 845 444 846
rect 438 841 439 845
rect 443 841 444 845
rect 484 844 486 874
rect 503 869 507 870
rect 511 874 515 875
rect 511 869 515 870
rect 559 874 563 875
rect 559 869 563 870
rect 591 874 595 875
rect 591 869 595 870
rect 623 874 627 875
rect 623 869 627 870
rect 679 874 683 875
rect 679 869 683 870
rect 695 874 699 875
rect 695 869 699 870
rect 759 874 763 875
rect 759 869 763 870
rect 767 874 771 875
rect 767 869 771 870
rect 823 874 827 875
rect 823 869 827 870
rect 847 874 851 875
rect 847 869 851 870
rect 887 874 891 875
rect 887 869 891 870
rect 919 874 923 875
rect 919 869 923 870
rect 951 874 955 875
rect 951 869 955 870
rect 983 874 987 875
rect 983 869 987 870
rect 1015 874 1019 875
rect 1015 869 1019 870
rect 1039 874 1043 875
rect 1039 869 1043 870
rect 1079 874 1083 875
rect 1079 869 1083 870
rect 1095 874 1099 875
rect 1095 869 1099 870
rect 1135 874 1139 875
rect 1135 869 1139 870
rect 1151 874 1155 875
rect 1151 869 1155 870
rect 1191 874 1195 875
rect 1191 869 1195 870
rect 1207 874 1211 875
rect 1207 869 1211 870
rect 1247 874 1251 875
rect 1247 869 1251 870
rect 1263 874 1267 875
rect 1263 869 1267 870
rect 512 864 514 869
rect 592 864 594 869
rect 680 864 682 869
rect 768 864 770 869
rect 848 864 850 869
rect 920 864 922 869
rect 984 864 986 869
rect 1040 864 1042 869
rect 1096 864 1098 869
rect 1152 864 1154 869
rect 1208 864 1210 869
rect 1264 864 1266 869
rect 1280 868 1282 890
rect 1288 876 1290 890
rect 1302 885 1308 886
rect 1302 881 1303 885
rect 1307 881 1308 885
rect 1302 880 1308 881
rect 1358 885 1364 886
rect 1358 881 1359 885
rect 1363 881 1364 885
rect 1358 880 1364 881
rect 1368 880 1370 922
rect 1374 921 1380 922
rect 1374 917 1375 921
rect 1379 917 1380 921
rect 1374 916 1380 917
rect 1422 921 1428 922
rect 1422 917 1423 921
rect 1427 917 1428 921
rect 1422 916 1428 917
rect 1470 921 1476 922
rect 1470 917 1471 921
rect 1475 917 1476 921
rect 1470 916 1476 917
rect 1510 921 1516 922
rect 1510 917 1511 921
rect 1515 917 1516 921
rect 1510 916 1516 917
rect 1542 921 1548 922
rect 1542 917 1543 921
rect 1547 917 1548 921
rect 1582 919 1583 923
rect 1587 919 1588 923
rect 1582 918 1588 919
rect 1542 916 1548 917
rect 1376 911 1378 916
rect 1424 911 1426 916
rect 1472 911 1474 916
rect 1512 911 1514 916
rect 1526 911 1532 912
rect 1544 911 1546 916
rect 1584 911 1586 918
rect 1375 910 1379 911
rect 1375 905 1379 906
rect 1407 910 1411 911
rect 1407 904 1411 906
rect 1423 910 1427 911
rect 1423 905 1427 906
rect 1455 910 1459 911
rect 1455 904 1459 906
rect 1471 910 1475 911
rect 1471 905 1475 906
rect 1511 910 1515 911
rect 1526 907 1527 911
rect 1531 907 1532 911
rect 1526 906 1532 907
rect 1543 910 1547 911
rect 1511 904 1515 906
rect 1406 903 1412 904
rect 1406 899 1407 903
rect 1411 899 1412 903
rect 1406 898 1412 899
rect 1454 903 1460 904
rect 1454 899 1455 903
rect 1459 899 1460 903
rect 1454 898 1460 899
rect 1510 903 1516 904
rect 1510 899 1511 903
rect 1515 899 1516 903
rect 1510 898 1516 899
rect 1406 885 1412 886
rect 1406 881 1407 885
rect 1411 881 1412 885
rect 1406 880 1412 881
rect 1454 885 1460 886
rect 1454 881 1455 885
rect 1459 881 1460 885
rect 1454 880 1460 881
rect 1510 885 1516 886
rect 1510 881 1511 885
rect 1515 881 1516 885
rect 1510 880 1516 881
rect 1528 880 1530 906
rect 1543 904 1547 906
rect 1583 910 1587 911
rect 1583 905 1587 906
rect 1542 903 1548 904
rect 1542 899 1543 903
rect 1547 899 1548 903
rect 1584 902 1586 905
rect 1542 898 1548 899
rect 1582 901 1588 902
rect 1582 897 1583 901
rect 1587 897 1588 901
rect 1582 896 1588 897
rect 1558 895 1564 896
rect 1558 891 1559 895
rect 1563 891 1564 895
rect 1558 890 1564 891
rect 1542 885 1548 886
rect 1542 881 1543 885
rect 1547 881 1548 885
rect 1542 880 1548 881
rect 1286 875 1292 876
rect 1304 875 1306 880
rect 1360 875 1362 880
rect 1366 879 1372 880
rect 1366 875 1367 879
rect 1371 875 1372 879
rect 1408 875 1410 880
rect 1456 875 1458 880
rect 1494 879 1500 880
rect 1494 875 1495 879
rect 1499 875 1500 879
rect 1512 875 1514 880
rect 1526 879 1532 880
rect 1526 875 1527 879
rect 1531 875 1532 879
rect 1544 875 1546 880
rect 1286 871 1287 875
rect 1291 871 1292 875
rect 1286 870 1292 871
rect 1303 874 1307 875
rect 1303 869 1307 870
rect 1327 874 1331 875
rect 1327 869 1331 870
rect 1359 874 1363 875
rect 1366 874 1372 875
rect 1399 874 1403 875
rect 1359 869 1363 870
rect 1399 869 1403 870
rect 1407 874 1411 875
rect 1407 869 1411 870
rect 1455 874 1459 875
rect 1455 869 1459 870
rect 1479 874 1483 875
rect 1494 874 1500 875
rect 1511 874 1515 875
rect 1526 874 1532 875
rect 1543 874 1547 875
rect 1479 869 1483 870
rect 1278 867 1284 868
rect 510 863 516 864
rect 510 859 511 863
rect 515 859 516 863
rect 510 858 516 859
rect 590 863 596 864
rect 590 859 591 863
rect 595 859 596 863
rect 590 858 596 859
rect 678 863 684 864
rect 678 859 679 863
rect 683 859 684 863
rect 678 858 684 859
rect 766 863 772 864
rect 766 859 767 863
rect 771 859 772 863
rect 766 858 772 859
rect 846 863 852 864
rect 846 859 847 863
rect 851 859 852 863
rect 846 858 852 859
rect 918 863 924 864
rect 918 859 919 863
rect 923 859 924 863
rect 918 858 924 859
rect 982 863 988 864
rect 982 859 983 863
rect 987 859 988 863
rect 982 858 988 859
rect 1038 863 1044 864
rect 1038 859 1039 863
rect 1043 859 1044 863
rect 1038 858 1044 859
rect 1094 863 1100 864
rect 1094 859 1095 863
rect 1099 859 1100 863
rect 1094 858 1100 859
rect 1150 863 1156 864
rect 1150 859 1151 863
rect 1155 859 1156 863
rect 1150 858 1156 859
rect 1206 863 1212 864
rect 1206 859 1207 863
rect 1211 859 1212 863
rect 1206 858 1212 859
rect 1262 863 1268 864
rect 1262 859 1263 863
rect 1267 859 1268 863
rect 1278 863 1279 867
rect 1283 863 1284 867
rect 1328 864 1330 869
rect 1400 864 1402 869
rect 1480 864 1482 869
rect 1278 862 1284 863
rect 1326 863 1332 864
rect 1262 858 1268 859
rect 1326 859 1327 863
rect 1331 859 1332 863
rect 1326 858 1332 859
rect 1398 863 1404 864
rect 1398 859 1399 863
rect 1403 859 1404 863
rect 1398 858 1404 859
rect 1478 863 1484 864
rect 1478 859 1479 863
rect 1483 859 1484 863
rect 1478 858 1484 859
rect 1496 852 1498 874
rect 1511 869 1515 870
rect 1543 869 1547 870
rect 1544 864 1546 869
rect 1560 868 1562 890
rect 1582 884 1588 885
rect 1582 880 1583 884
rect 1587 880 1588 884
rect 1582 879 1588 880
rect 1584 875 1586 879
rect 1583 874 1587 875
rect 1583 869 1587 870
rect 1558 867 1564 868
rect 1542 863 1548 864
rect 1542 859 1543 863
rect 1547 859 1548 863
rect 1558 863 1559 867
rect 1563 863 1564 867
rect 1584 865 1586 869
rect 1558 862 1564 863
rect 1582 864 1588 865
rect 1582 860 1583 864
rect 1587 860 1588 864
rect 1582 859 1588 860
rect 1542 858 1548 859
rect 1494 851 1500 852
rect 1494 847 1495 851
rect 1499 847 1500 851
rect 1494 846 1500 847
rect 1582 847 1588 848
rect 510 845 516 846
rect 438 840 444 841
rect 482 843 488 844
rect 304 835 306 840
rect 344 835 346 840
rect 384 835 386 840
rect 440 835 442 840
rect 482 839 483 843
rect 487 839 488 843
rect 510 841 511 845
rect 515 841 516 845
rect 510 840 516 841
rect 590 845 596 846
rect 590 841 591 845
rect 595 841 596 845
rect 590 840 596 841
rect 678 845 684 846
rect 678 841 679 845
rect 683 841 684 845
rect 678 840 684 841
rect 766 845 772 846
rect 766 841 767 845
rect 771 841 772 845
rect 766 840 772 841
rect 846 845 852 846
rect 846 841 847 845
rect 851 841 852 845
rect 846 840 852 841
rect 918 845 924 846
rect 918 841 919 845
rect 923 841 924 845
rect 918 840 924 841
rect 982 845 988 846
rect 982 841 983 845
rect 987 841 988 845
rect 982 840 988 841
rect 1038 845 1044 846
rect 1038 841 1039 845
rect 1043 841 1044 845
rect 1038 840 1044 841
rect 1094 845 1100 846
rect 1094 841 1095 845
rect 1099 841 1100 845
rect 1094 840 1100 841
rect 1150 845 1156 846
rect 1150 841 1151 845
rect 1155 841 1156 845
rect 1150 840 1156 841
rect 1206 845 1212 846
rect 1206 841 1207 845
rect 1211 841 1212 845
rect 1206 840 1212 841
rect 1262 845 1268 846
rect 1262 841 1263 845
rect 1267 841 1268 845
rect 1262 840 1268 841
rect 1326 845 1332 846
rect 1326 841 1327 845
rect 1331 841 1332 845
rect 1326 840 1332 841
rect 1398 845 1404 846
rect 1398 841 1399 845
rect 1403 841 1404 845
rect 1398 840 1404 841
rect 1478 845 1484 846
rect 1478 841 1479 845
rect 1483 841 1484 845
rect 1478 840 1484 841
rect 1542 845 1548 846
rect 1542 841 1543 845
rect 1547 841 1548 845
rect 1582 843 1583 847
rect 1587 843 1588 847
rect 1582 842 1588 843
rect 1542 840 1548 841
rect 482 838 488 839
rect 512 835 514 840
rect 592 835 594 840
rect 680 835 682 840
rect 768 835 770 840
rect 848 835 850 840
rect 920 835 922 840
rect 984 835 986 840
rect 1018 839 1024 840
rect 1018 835 1019 839
rect 1023 835 1024 839
rect 1040 835 1042 840
rect 1096 835 1098 840
rect 1152 835 1154 840
rect 1208 835 1210 840
rect 1264 835 1266 840
rect 1328 835 1330 840
rect 1400 835 1402 840
rect 1480 835 1482 840
rect 1544 835 1546 840
rect 1584 835 1586 842
rect 287 834 291 835
rect 287 828 291 830
rect 303 834 307 835
rect 303 829 307 830
rect 343 834 347 835
rect 343 829 347 830
rect 351 834 355 835
rect 351 828 355 830
rect 383 834 387 835
rect 383 829 387 830
rect 423 834 427 835
rect 423 828 427 830
rect 439 834 443 835
rect 439 829 443 830
rect 495 834 499 835
rect 495 828 499 830
rect 511 834 515 835
rect 511 829 515 830
rect 567 834 571 835
rect 567 828 571 830
rect 591 834 595 835
rect 591 829 595 830
rect 639 834 643 835
rect 639 828 643 830
rect 679 834 683 835
rect 679 829 683 830
rect 719 834 723 835
rect 719 828 723 830
rect 767 834 771 835
rect 767 829 771 830
rect 791 834 795 835
rect 791 828 795 830
rect 847 834 851 835
rect 847 829 851 830
rect 863 834 867 835
rect 863 828 867 830
rect 919 834 923 835
rect 919 829 923 830
rect 935 834 939 835
rect 935 828 939 830
rect 983 834 987 835
rect 983 829 987 830
rect 999 834 1003 835
rect 1018 834 1024 835
rect 1039 834 1043 835
rect 999 828 1003 830
rect 286 827 292 828
rect 286 823 287 827
rect 291 823 292 827
rect 286 822 292 823
rect 350 827 356 828
rect 350 823 351 827
rect 355 823 356 827
rect 350 822 356 823
rect 422 827 428 828
rect 422 823 423 827
rect 427 823 428 827
rect 422 822 428 823
rect 494 827 500 828
rect 494 823 495 827
rect 499 823 500 827
rect 494 822 500 823
rect 566 827 572 828
rect 566 823 567 827
rect 571 823 572 827
rect 566 822 572 823
rect 638 827 644 828
rect 638 823 639 827
rect 643 823 644 827
rect 638 822 644 823
rect 718 827 724 828
rect 718 823 719 827
rect 723 823 724 827
rect 718 822 724 823
rect 790 827 796 828
rect 790 823 791 827
rect 795 823 796 827
rect 790 822 796 823
rect 862 827 868 828
rect 862 823 863 827
rect 867 823 868 827
rect 862 822 868 823
rect 934 827 940 828
rect 934 823 935 827
rect 939 823 940 827
rect 934 822 940 823
rect 998 827 1004 828
rect 998 823 999 827
rect 1003 823 1004 827
rect 998 822 1004 823
rect 266 819 272 820
rect 266 815 267 819
rect 271 815 272 819
rect 266 814 272 815
rect 750 819 756 820
rect 750 815 751 819
rect 755 815 756 819
rect 750 814 756 815
rect 222 809 228 810
rect 222 805 223 809
rect 227 805 228 809
rect 222 804 228 805
rect 286 809 292 810
rect 286 805 287 809
rect 291 805 292 809
rect 286 804 292 805
rect 350 809 356 810
rect 350 805 351 809
rect 355 805 356 809
rect 350 804 356 805
rect 422 809 428 810
rect 422 805 423 809
rect 427 805 428 809
rect 422 804 428 805
rect 494 809 500 810
rect 494 805 495 809
rect 499 805 500 809
rect 494 804 500 805
rect 566 809 572 810
rect 566 805 567 809
rect 571 805 572 809
rect 566 804 572 805
rect 638 809 644 810
rect 638 805 639 809
rect 643 805 644 809
rect 638 804 644 805
rect 718 809 724 810
rect 718 805 719 809
rect 723 805 724 809
rect 718 804 724 805
rect 168 799 170 804
rect 214 803 220 804
rect 214 799 215 803
rect 219 799 220 803
rect 224 799 226 804
rect 288 799 290 804
rect 352 799 354 804
rect 370 803 376 804
rect 370 799 371 803
rect 375 799 376 803
rect 424 799 426 804
rect 496 799 498 804
rect 502 803 508 804
rect 502 799 503 803
rect 507 799 508 803
rect 568 799 570 804
rect 640 799 642 804
rect 686 803 692 804
rect 686 799 687 803
rect 691 799 692 803
rect 720 799 722 804
rect 167 798 171 799
rect 167 793 171 794
rect 199 798 203 799
rect 214 798 220 799
rect 223 798 227 799
rect 199 793 203 794
rect 223 793 227 794
rect 247 798 251 799
rect 247 793 251 794
rect 287 798 291 799
rect 287 793 291 794
rect 303 798 307 799
rect 303 793 307 794
rect 351 798 355 799
rect 351 793 355 794
rect 359 798 363 799
rect 370 798 376 799
rect 423 798 427 799
rect 359 793 363 794
rect 150 791 156 792
rect 110 784 111 788
rect 115 784 116 788
rect 110 783 116 784
rect 134 787 140 788
rect 134 783 135 787
rect 139 783 140 787
rect 150 787 151 791
rect 155 787 156 791
rect 168 788 170 793
rect 200 788 202 793
rect 248 788 250 793
rect 304 788 306 793
rect 360 788 362 793
rect 150 786 156 787
rect 166 787 172 788
rect 134 782 140 783
rect 166 783 167 787
rect 171 783 172 787
rect 166 782 172 783
rect 198 787 204 788
rect 198 783 199 787
rect 203 783 204 787
rect 198 782 204 783
rect 246 787 252 788
rect 246 783 247 787
rect 251 783 252 787
rect 246 782 252 783
rect 302 787 308 788
rect 302 783 303 787
rect 307 783 308 787
rect 302 782 308 783
rect 358 787 364 788
rect 358 783 359 787
rect 363 783 364 787
rect 358 782 364 783
rect 372 776 374 798
rect 423 793 427 794
rect 487 798 491 799
rect 487 793 491 794
rect 495 798 499 799
rect 502 798 508 799
rect 551 798 555 799
rect 495 793 499 794
rect 424 788 426 793
rect 488 788 490 793
rect 422 787 428 788
rect 422 783 423 787
rect 427 783 428 787
rect 422 782 428 783
rect 486 787 492 788
rect 486 783 487 787
rect 491 783 492 787
rect 486 782 492 783
rect 214 775 220 776
rect 110 771 116 772
rect 110 767 111 771
rect 115 767 116 771
rect 214 771 215 775
rect 219 771 220 775
rect 214 770 220 771
rect 370 775 376 776
rect 370 771 371 775
rect 375 771 376 775
rect 370 770 376 771
rect 110 766 116 767
rect 134 769 140 770
rect 112 763 114 766
rect 134 765 135 769
rect 139 765 140 769
rect 134 764 140 765
rect 166 769 172 770
rect 166 765 167 769
rect 171 765 172 769
rect 166 764 172 765
rect 198 769 204 770
rect 198 765 199 769
rect 203 765 204 769
rect 198 764 204 765
rect 111 762 115 763
rect 111 757 115 758
rect 135 762 139 764
rect 112 754 114 757
rect 135 756 139 758
rect 167 762 171 764
rect 167 756 171 758
rect 199 762 203 764
rect 199 756 203 758
rect 134 755 140 756
rect 110 753 116 754
rect 110 749 111 753
rect 115 749 116 753
rect 134 751 135 755
rect 139 751 140 755
rect 134 750 140 751
rect 166 755 172 756
rect 166 751 167 755
rect 171 751 172 755
rect 166 750 172 751
rect 198 755 204 756
rect 198 751 199 755
rect 203 751 204 755
rect 198 750 204 751
rect 110 748 116 749
rect 150 747 156 748
rect 150 743 151 747
rect 155 743 156 747
rect 150 742 156 743
rect 134 737 140 738
rect 110 736 116 737
rect 110 732 111 736
rect 115 732 116 736
rect 134 733 135 737
rect 139 733 140 737
rect 134 732 140 733
rect 110 731 116 732
rect 112 727 114 731
rect 136 727 138 732
rect 111 726 115 727
rect 111 721 115 722
rect 135 726 139 727
rect 135 721 139 722
rect 112 717 114 721
rect 110 716 116 717
rect 136 716 138 721
rect 152 720 154 742
rect 216 740 218 770
rect 246 769 252 770
rect 246 765 247 769
rect 251 765 252 769
rect 246 764 252 765
rect 302 769 308 770
rect 302 765 303 769
rect 307 765 308 769
rect 302 764 308 765
rect 358 769 364 770
rect 358 765 359 769
rect 363 765 364 769
rect 358 764 364 765
rect 422 769 428 770
rect 422 765 423 769
rect 427 765 428 769
rect 422 764 428 765
rect 486 769 492 770
rect 486 765 487 769
rect 491 765 492 769
rect 486 764 492 765
rect 247 762 251 764
rect 247 757 251 758
rect 255 762 259 763
rect 255 756 259 758
rect 303 762 307 764
rect 303 757 307 758
rect 319 762 323 763
rect 319 756 323 758
rect 359 762 363 764
rect 359 757 363 758
rect 391 762 395 763
rect 391 756 395 758
rect 423 762 427 764
rect 423 757 427 758
rect 463 762 467 763
rect 463 756 467 758
rect 487 762 491 764
rect 487 757 491 758
rect 254 755 260 756
rect 254 751 255 755
rect 259 751 260 755
rect 254 750 260 751
rect 318 755 324 756
rect 318 751 319 755
rect 323 751 324 755
rect 318 750 324 751
rect 390 755 396 756
rect 390 751 391 755
rect 395 751 396 755
rect 390 750 396 751
rect 462 755 468 756
rect 462 751 463 755
rect 467 751 468 755
rect 462 750 468 751
rect 504 748 506 798
rect 551 793 555 794
rect 567 798 571 799
rect 567 793 571 794
rect 607 798 611 799
rect 607 793 611 794
rect 639 798 643 799
rect 639 793 643 794
rect 671 798 675 799
rect 686 798 692 799
rect 719 798 723 799
rect 671 793 675 794
rect 552 788 554 793
rect 598 791 604 792
rect 550 787 556 788
rect 550 783 551 787
rect 555 783 556 787
rect 598 787 599 791
rect 603 787 604 791
rect 608 788 610 793
rect 672 788 674 793
rect 598 786 604 787
rect 606 787 612 788
rect 550 782 556 783
rect 534 775 540 776
rect 534 771 535 775
rect 539 771 540 775
rect 534 770 540 771
rect 502 747 508 748
rect 502 743 503 747
rect 507 743 508 747
rect 502 742 508 743
rect 214 739 220 740
rect 166 737 172 738
rect 166 733 167 737
rect 171 733 172 737
rect 166 732 172 733
rect 198 737 204 738
rect 198 733 199 737
rect 203 733 204 737
rect 214 735 215 739
rect 219 735 220 739
rect 214 734 220 735
rect 254 737 260 738
rect 198 732 204 733
rect 254 733 255 737
rect 259 733 260 737
rect 254 732 260 733
rect 318 737 324 738
rect 318 733 319 737
rect 323 733 324 737
rect 318 732 324 733
rect 390 737 396 738
rect 390 733 391 737
rect 395 733 396 737
rect 390 732 396 733
rect 462 737 468 738
rect 462 733 463 737
rect 467 733 468 737
rect 462 732 468 733
rect 536 732 538 770
rect 550 769 556 770
rect 550 765 551 769
rect 555 765 556 769
rect 550 764 556 765
rect 543 762 547 763
rect 543 756 547 758
rect 551 762 555 764
rect 551 757 555 758
rect 542 755 548 756
rect 542 751 543 755
rect 547 751 548 755
rect 542 750 548 751
rect 600 748 602 786
rect 606 783 607 787
rect 611 783 612 787
rect 606 782 612 783
rect 670 787 676 788
rect 670 783 671 787
rect 675 783 676 787
rect 670 782 676 783
rect 688 776 690 798
rect 719 793 723 794
rect 735 798 739 799
rect 735 793 739 794
rect 736 788 738 793
rect 752 792 754 814
rect 790 809 796 810
rect 790 805 791 809
rect 795 805 796 809
rect 790 804 796 805
rect 862 809 868 810
rect 862 805 863 809
rect 867 805 868 809
rect 862 804 868 805
rect 934 809 940 810
rect 934 805 935 809
rect 939 805 940 809
rect 934 804 940 805
rect 998 809 1004 810
rect 998 805 999 809
rect 1003 805 1004 809
rect 998 804 1004 805
rect 1020 804 1022 834
rect 1039 829 1043 830
rect 1055 834 1059 835
rect 1055 828 1059 830
rect 1095 834 1099 835
rect 1095 829 1099 830
rect 1103 834 1107 835
rect 1103 828 1107 830
rect 1143 834 1147 835
rect 1143 828 1147 830
rect 1151 834 1155 835
rect 1151 829 1155 830
rect 1183 834 1187 835
rect 1183 828 1187 830
rect 1207 834 1211 835
rect 1207 829 1211 830
rect 1231 834 1235 835
rect 1263 834 1267 835
rect 1231 828 1235 830
rect 1246 831 1252 832
rect 1054 827 1060 828
rect 1054 823 1055 827
rect 1059 823 1060 827
rect 1054 822 1060 823
rect 1102 827 1108 828
rect 1102 823 1103 827
rect 1107 823 1108 827
rect 1102 822 1108 823
rect 1142 827 1148 828
rect 1142 823 1143 827
rect 1147 823 1148 827
rect 1142 822 1148 823
rect 1182 827 1188 828
rect 1182 823 1183 827
rect 1187 823 1188 827
rect 1182 822 1188 823
rect 1230 827 1236 828
rect 1230 823 1231 827
rect 1235 823 1236 827
rect 1246 827 1247 831
rect 1251 827 1252 831
rect 1263 829 1267 830
rect 1279 834 1283 835
rect 1279 828 1283 830
rect 1327 834 1331 835
rect 1327 828 1331 830
rect 1399 834 1403 835
rect 1399 829 1403 830
rect 1479 834 1483 835
rect 1479 829 1483 830
rect 1543 834 1547 835
rect 1543 829 1547 830
rect 1583 834 1587 835
rect 1583 829 1587 830
rect 1246 826 1252 827
rect 1278 827 1284 828
rect 1230 822 1236 823
rect 1086 819 1092 820
rect 1086 815 1087 819
rect 1091 815 1092 819
rect 1086 814 1092 815
rect 1054 809 1060 810
rect 1054 805 1055 809
rect 1059 805 1060 809
rect 1054 804 1060 805
rect 792 799 794 804
rect 864 799 866 804
rect 936 799 938 804
rect 1000 799 1002 804
rect 1006 803 1012 804
rect 1006 799 1007 803
rect 1011 799 1012 803
rect 791 798 795 799
rect 791 793 795 794
rect 799 798 803 799
rect 799 793 803 794
rect 863 798 867 799
rect 863 793 867 794
rect 871 798 875 799
rect 871 793 875 794
rect 935 798 939 799
rect 935 793 939 794
rect 999 798 1003 799
rect 1006 798 1012 799
rect 1018 803 1024 804
rect 1018 799 1019 803
rect 1023 799 1024 803
rect 1056 799 1058 804
rect 1088 800 1090 814
rect 1102 809 1108 810
rect 1102 805 1103 809
rect 1107 805 1108 809
rect 1102 804 1108 805
rect 1142 809 1148 810
rect 1142 805 1143 809
rect 1147 805 1148 809
rect 1142 804 1148 805
rect 1182 809 1188 810
rect 1182 805 1183 809
rect 1187 805 1188 809
rect 1182 804 1188 805
rect 1230 809 1236 810
rect 1230 805 1231 809
rect 1235 805 1236 809
rect 1230 804 1236 805
rect 1086 799 1092 800
rect 1104 799 1106 804
rect 1144 799 1146 804
rect 1184 799 1186 804
rect 1232 799 1234 804
rect 1018 798 1024 799
rect 1055 798 1059 799
rect 999 793 1003 794
rect 750 791 756 792
rect 734 787 740 788
rect 734 783 735 787
rect 739 783 740 787
rect 750 787 751 791
rect 755 787 756 791
rect 800 788 802 793
rect 872 788 874 793
rect 882 791 888 792
rect 750 786 756 787
rect 798 787 804 788
rect 734 782 740 783
rect 798 783 799 787
rect 803 783 804 787
rect 798 782 804 783
rect 870 787 876 788
rect 870 783 871 787
rect 875 783 876 787
rect 882 787 883 791
rect 887 787 888 791
rect 936 788 938 793
rect 1000 788 1002 793
rect 882 786 888 787
rect 934 787 940 788
rect 870 782 876 783
rect 686 775 692 776
rect 686 771 687 775
rect 691 771 692 775
rect 686 770 692 771
rect 810 775 816 776
rect 810 771 811 775
rect 815 771 816 775
rect 810 770 816 771
rect 606 769 612 770
rect 606 765 607 769
rect 611 765 612 769
rect 606 764 612 765
rect 670 769 676 770
rect 670 765 671 769
rect 675 765 676 769
rect 670 764 676 765
rect 734 769 740 770
rect 734 765 735 769
rect 739 765 740 769
rect 734 764 740 765
rect 798 769 804 770
rect 798 765 799 769
rect 803 765 804 769
rect 798 764 804 765
rect 607 762 611 764
rect 607 757 611 758
rect 623 762 627 763
rect 623 756 627 758
rect 671 762 675 764
rect 671 757 675 758
rect 703 762 707 763
rect 703 756 707 758
rect 735 762 739 764
rect 735 757 739 758
rect 775 762 779 763
rect 775 756 779 758
rect 799 762 803 764
rect 799 757 803 758
rect 622 755 628 756
rect 622 751 623 755
rect 627 751 628 755
rect 622 750 628 751
rect 702 755 708 756
rect 702 751 703 755
rect 707 751 708 755
rect 702 750 708 751
rect 774 755 780 756
rect 774 751 775 755
rect 779 751 780 755
rect 774 750 780 751
rect 558 747 564 748
rect 558 743 559 747
rect 563 743 564 747
rect 558 742 564 743
rect 598 747 604 748
rect 598 743 599 747
rect 603 743 604 747
rect 598 742 604 743
rect 766 747 772 748
rect 766 743 767 747
rect 771 743 772 747
rect 766 742 772 743
rect 542 737 548 738
rect 542 733 543 737
rect 547 733 548 737
rect 542 732 548 733
rect 168 727 170 732
rect 200 727 202 732
rect 256 727 258 732
rect 320 727 322 732
rect 392 727 394 732
rect 398 731 404 732
rect 398 727 399 731
rect 403 727 404 731
rect 442 731 448 732
rect 442 727 443 731
rect 447 727 448 731
rect 464 727 466 732
rect 534 731 540 732
rect 534 727 535 731
rect 539 727 540 731
rect 544 727 546 732
rect 167 726 171 727
rect 167 721 171 722
rect 199 726 203 727
rect 199 721 203 722
rect 207 726 211 727
rect 207 721 211 722
rect 255 726 259 727
rect 255 721 259 722
rect 311 726 315 727
rect 311 721 315 722
rect 319 726 323 727
rect 319 721 323 722
rect 367 726 371 727
rect 367 721 371 722
rect 391 726 395 727
rect 398 726 404 727
rect 423 726 427 727
rect 442 726 448 727
rect 463 726 467 727
rect 391 721 395 722
rect 150 719 156 720
rect 110 712 111 716
rect 115 712 116 716
rect 110 711 116 712
rect 134 715 140 716
rect 134 711 135 715
rect 139 711 140 715
rect 150 715 151 719
rect 155 715 156 719
rect 168 716 170 721
rect 208 716 210 721
rect 256 716 258 721
rect 270 719 276 720
rect 150 714 156 715
rect 166 715 172 716
rect 134 710 140 711
rect 166 711 167 715
rect 171 711 172 715
rect 166 710 172 711
rect 206 715 212 716
rect 206 711 207 715
rect 211 711 212 715
rect 206 710 212 711
rect 254 715 260 716
rect 254 711 255 715
rect 259 711 260 715
rect 270 715 271 719
rect 275 715 276 719
rect 312 716 314 721
rect 368 716 370 721
rect 270 714 276 715
rect 310 715 316 716
rect 254 710 260 711
rect 222 703 228 704
rect 110 699 116 700
rect 110 695 111 699
rect 115 695 116 699
rect 222 699 223 703
rect 227 699 228 703
rect 222 698 228 699
rect 110 694 116 695
rect 134 697 140 698
rect 112 691 114 694
rect 134 693 135 697
rect 139 693 140 697
rect 134 692 140 693
rect 166 697 172 698
rect 166 693 167 697
rect 171 693 172 697
rect 166 692 172 693
rect 206 697 212 698
rect 206 693 207 697
rect 211 693 212 697
rect 206 692 212 693
rect 111 690 115 691
rect 111 685 115 686
rect 135 690 139 692
rect 135 685 139 686
rect 159 690 163 691
rect 112 682 114 685
rect 159 684 163 686
rect 167 690 171 692
rect 167 685 171 686
rect 207 690 211 692
rect 207 684 211 686
rect 158 683 164 684
rect 110 681 116 682
rect 110 677 111 681
rect 115 677 116 681
rect 158 679 159 683
rect 163 679 164 683
rect 158 678 164 679
rect 206 683 212 684
rect 206 679 207 683
rect 211 679 212 683
rect 206 678 212 679
rect 110 676 116 677
rect 178 675 184 676
rect 178 671 179 675
rect 183 671 184 675
rect 178 670 184 671
rect 158 665 164 666
rect 110 664 116 665
rect 110 660 111 664
rect 115 660 116 664
rect 158 661 159 665
rect 163 661 164 665
rect 158 660 164 661
rect 110 659 116 660
rect 112 651 114 659
rect 160 651 162 660
rect 111 650 115 651
rect 111 645 115 646
rect 159 650 163 651
rect 159 645 163 646
rect 167 650 171 651
rect 167 645 171 646
rect 112 641 114 645
rect 110 640 116 641
rect 168 640 170 645
rect 180 644 182 670
rect 206 665 212 666
rect 206 661 207 665
rect 211 661 212 665
rect 206 660 212 661
rect 224 660 226 698
rect 254 697 260 698
rect 254 693 255 697
rect 259 693 260 697
rect 254 692 260 693
rect 255 690 259 692
rect 255 684 259 686
rect 254 683 260 684
rect 254 679 255 683
rect 259 679 260 683
rect 254 678 260 679
rect 272 676 274 714
rect 310 711 311 715
rect 315 711 316 715
rect 310 710 316 711
rect 366 715 372 716
rect 366 711 367 715
rect 371 711 372 715
rect 366 710 372 711
rect 400 704 402 726
rect 423 721 427 722
rect 424 716 426 721
rect 434 719 440 720
rect 422 715 428 716
rect 422 711 423 715
rect 427 711 428 715
rect 434 715 435 719
rect 439 715 440 719
rect 434 714 440 715
rect 422 710 428 711
rect 398 703 404 704
rect 398 699 399 703
rect 403 699 404 703
rect 398 698 404 699
rect 310 697 316 698
rect 310 693 311 697
rect 315 693 316 697
rect 310 692 316 693
rect 366 697 372 698
rect 366 693 367 697
rect 371 693 372 697
rect 366 692 372 693
rect 422 697 428 698
rect 422 693 423 697
rect 427 693 428 697
rect 422 692 428 693
rect 303 690 307 691
rect 303 684 307 686
rect 311 690 315 692
rect 311 685 315 686
rect 359 690 363 691
rect 359 684 363 686
rect 367 690 371 692
rect 367 685 371 686
rect 415 690 419 691
rect 415 684 419 686
rect 423 690 427 692
rect 423 685 427 686
rect 302 683 308 684
rect 302 679 303 683
rect 307 679 308 683
rect 302 678 308 679
rect 358 683 364 684
rect 358 679 359 683
rect 363 679 364 683
rect 358 678 364 679
rect 414 683 420 684
rect 414 679 415 683
rect 419 679 420 683
rect 414 678 420 679
rect 436 676 438 714
rect 444 704 446 726
rect 463 721 467 722
rect 479 726 483 727
rect 534 726 540 727
rect 543 726 547 727
rect 479 721 483 722
rect 543 721 547 722
rect 480 716 482 721
rect 544 716 546 721
rect 560 720 562 742
rect 622 737 628 738
rect 622 733 623 737
rect 627 733 628 737
rect 622 732 628 733
rect 702 737 708 738
rect 702 733 703 737
rect 707 733 708 737
rect 702 732 708 733
rect 624 727 626 732
rect 634 731 640 732
rect 634 727 635 731
rect 639 727 640 731
rect 704 727 706 732
rect 615 726 619 727
rect 615 721 619 722
rect 623 726 627 727
rect 634 726 640 727
rect 687 726 691 727
rect 623 721 627 722
rect 558 719 564 720
rect 478 715 484 716
rect 478 711 479 715
rect 483 711 484 715
rect 478 710 484 711
rect 542 715 548 716
rect 542 711 543 715
rect 547 711 548 715
rect 558 715 559 719
rect 563 715 564 719
rect 616 716 618 721
rect 558 714 564 715
rect 614 715 620 716
rect 542 710 548 711
rect 614 711 615 715
rect 619 711 620 715
rect 614 710 620 711
rect 636 704 638 726
rect 658 723 664 724
rect 658 719 659 723
rect 663 719 664 723
rect 687 721 691 722
rect 703 726 707 727
rect 703 721 707 722
rect 759 726 763 727
rect 768 724 770 742
rect 774 737 780 738
rect 774 733 775 737
rect 779 733 780 737
rect 774 732 780 733
rect 812 732 814 770
rect 870 769 876 770
rect 870 765 871 769
rect 875 765 876 769
rect 870 764 876 765
rect 847 762 851 763
rect 847 756 851 758
rect 871 762 875 764
rect 871 757 875 758
rect 846 755 852 756
rect 846 751 847 755
rect 851 751 852 755
rect 846 750 852 751
rect 884 748 886 786
rect 934 783 935 787
rect 939 783 940 787
rect 934 782 940 783
rect 998 787 1004 788
rect 998 783 999 787
rect 1003 783 1004 787
rect 998 782 1004 783
rect 1008 772 1010 798
rect 1055 793 1059 794
rect 1063 798 1067 799
rect 1086 795 1087 799
rect 1091 795 1092 799
rect 1086 794 1092 795
rect 1103 798 1107 799
rect 1063 793 1067 794
rect 1103 793 1107 794
rect 1127 798 1131 799
rect 1127 793 1131 794
rect 1143 798 1147 799
rect 1143 793 1147 794
rect 1183 798 1187 799
rect 1183 793 1187 794
rect 1191 798 1195 799
rect 1191 793 1195 794
rect 1231 798 1235 799
rect 1231 793 1235 794
rect 1064 788 1066 793
rect 1128 788 1130 793
rect 1192 788 1194 793
rect 1248 792 1250 826
rect 1278 823 1279 827
rect 1283 823 1284 827
rect 1278 822 1284 823
rect 1326 827 1332 828
rect 1326 823 1327 827
rect 1331 823 1332 827
rect 1584 826 1586 829
rect 1326 822 1332 823
rect 1582 825 1588 826
rect 1582 821 1583 825
rect 1587 821 1588 825
rect 1582 820 1588 821
rect 1278 809 1284 810
rect 1278 805 1279 809
rect 1283 805 1284 809
rect 1278 804 1284 805
rect 1326 809 1332 810
rect 1326 805 1327 809
rect 1331 805 1332 809
rect 1326 804 1332 805
rect 1582 808 1588 809
rect 1582 804 1583 808
rect 1587 804 1588 808
rect 1280 799 1282 804
rect 1328 799 1330 804
rect 1582 803 1588 804
rect 1584 799 1586 803
rect 1255 798 1259 799
rect 1255 793 1259 794
rect 1279 798 1283 799
rect 1279 793 1283 794
rect 1319 798 1323 799
rect 1319 793 1323 794
rect 1327 798 1331 799
rect 1327 793 1331 794
rect 1383 798 1387 799
rect 1383 793 1387 794
rect 1583 798 1587 799
rect 1583 793 1587 794
rect 1246 791 1252 792
rect 1062 787 1068 788
rect 1062 783 1063 787
rect 1067 783 1068 787
rect 1062 782 1068 783
rect 1126 787 1132 788
rect 1126 783 1127 787
rect 1131 783 1132 787
rect 1126 782 1132 783
rect 1190 787 1196 788
rect 1190 783 1191 787
rect 1195 783 1196 787
rect 1246 787 1247 791
rect 1251 787 1252 791
rect 1256 788 1258 793
rect 1320 788 1322 793
rect 1384 788 1386 793
rect 1584 789 1586 793
rect 1582 788 1588 789
rect 1246 786 1252 787
rect 1254 787 1260 788
rect 1190 782 1196 783
rect 1254 783 1255 787
rect 1259 783 1260 787
rect 1254 782 1260 783
rect 1318 787 1324 788
rect 1318 783 1319 787
rect 1323 783 1324 787
rect 1318 782 1324 783
rect 1382 787 1388 788
rect 1382 783 1383 787
rect 1387 783 1388 787
rect 1582 784 1583 788
rect 1587 784 1588 788
rect 1582 783 1588 784
rect 1382 782 1388 783
rect 1078 775 1084 776
rect 1008 771 1016 772
rect 934 769 940 770
rect 934 765 935 769
rect 939 765 940 769
rect 934 764 940 765
rect 998 769 1004 770
rect 1008 769 1011 771
rect 998 765 999 769
rect 1003 765 1004 769
rect 1010 767 1011 769
rect 1015 767 1016 771
rect 1078 771 1079 775
rect 1083 771 1084 775
rect 1078 770 1084 771
rect 1582 771 1588 772
rect 1010 766 1016 767
rect 1062 769 1068 770
rect 998 764 1004 765
rect 1062 765 1063 769
rect 1067 765 1068 769
rect 1062 764 1068 765
rect 919 762 923 763
rect 919 756 923 758
rect 935 762 939 764
rect 935 757 939 758
rect 991 762 995 763
rect 991 756 995 758
rect 999 762 1003 764
rect 999 757 1003 758
rect 1063 762 1067 764
rect 1063 756 1067 758
rect 918 755 924 756
rect 918 751 919 755
rect 923 751 924 755
rect 918 750 924 751
rect 990 755 996 756
rect 990 751 991 755
rect 995 751 996 755
rect 990 750 996 751
rect 1062 755 1068 756
rect 1062 751 1063 755
rect 1067 751 1068 755
rect 1062 750 1068 751
rect 882 747 888 748
rect 882 743 883 747
rect 887 743 888 747
rect 882 742 888 743
rect 846 737 852 738
rect 846 733 847 737
rect 851 733 852 737
rect 846 732 852 733
rect 918 737 924 738
rect 918 733 919 737
rect 923 733 924 737
rect 918 732 924 733
rect 990 737 996 738
rect 990 733 991 737
rect 995 733 996 737
rect 990 732 996 733
rect 1062 737 1068 738
rect 1062 733 1063 737
rect 1067 733 1068 737
rect 1062 732 1068 733
rect 1080 732 1082 770
rect 1126 769 1132 770
rect 1126 765 1127 769
rect 1131 765 1132 769
rect 1126 764 1132 765
rect 1190 769 1196 770
rect 1190 765 1191 769
rect 1195 765 1196 769
rect 1190 764 1196 765
rect 1254 769 1260 770
rect 1254 765 1255 769
rect 1259 765 1260 769
rect 1254 764 1260 765
rect 1318 769 1324 770
rect 1318 765 1319 769
rect 1323 765 1324 769
rect 1318 764 1324 765
rect 1382 769 1388 770
rect 1382 765 1383 769
rect 1387 765 1388 769
rect 1582 767 1583 771
rect 1587 767 1588 771
rect 1582 766 1588 767
rect 1382 764 1388 765
rect 1127 762 1131 764
rect 1127 757 1131 758
rect 1135 762 1139 763
rect 1135 756 1139 758
rect 1191 762 1195 764
rect 1191 757 1195 758
rect 1207 762 1211 763
rect 1207 756 1211 758
rect 1255 762 1259 764
rect 1290 763 1296 764
rect 1255 757 1259 758
rect 1271 762 1275 763
rect 1290 759 1291 763
rect 1295 759 1296 763
rect 1290 758 1296 759
rect 1319 762 1323 764
rect 1271 756 1275 758
rect 1134 755 1140 756
rect 1134 751 1135 755
rect 1139 751 1140 755
rect 1134 750 1140 751
rect 1206 755 1212 756
rect 1206 751 1207 755
rect 1211 751 1212 755
rect 1206 750 1212 751
rect 1270 755 1276 756
rect 1270 751 1271 755
rect 1275 751 1276 755
rect 1270 750 1276 751
rect 1186 747 1192 748
rect 1186 743 1187 747
rect 1191 743 1192 747
rect 1186 742 1192 743
rect 1134 737 1140 738
rect 1134 733 1135 737
rect 1139 733 1140 737
rect 1134 732 1140 733
rect 776 727 778 732
rect 810 731 816 732
rect 810 727 811 731
rect 815 727 816 731
rect 848 727 850 732
rect 920 727 922 732
rect 992 727 994 732
rect 1022 731 1028 732
rect 1022 727 1023 731
rect 1027 727 1028 731
rect 1064 727 1066 732
rect 1078 731 1084 732
rect 1078 727 1079 731
rect 1083 727 1084 731
rect 1136 727 1138 732
rect 775 726 779 727
rect 810 726 816 727
rect 839 726 843 727
rect 759 721 763 722
rect 766 723 772 724
rect 658 718 664 719
rect 442 703 448 704
rect 442 699 443 703
rect 447 699 448 703
rect 442 698 448 699
rect 534 703 540 704
rect 534 699 535 703
rect 539 699 540 703
rect 534 698 540 699
rect 634 703 640 704
rect 634 699 635 703
rect 639 699 640 703
rect 634 698 640 699
rect 478 697 484 698
rect 478 693 479 697
rect 483 693 484 697
rect 478 692 484 693
rect 471 690 475 691
rect 471 684 475 686
rect 479 690 483 692
rect 479 685 483 686
rect 527 690 531 691
rect 527 684 531 686
rect 470 683 476 684
rect 470 679 471 683
rect 475 679 476 683
rect 470 678 476 679
rect 526 683 532 684
rect 526 679 527 683
rect 531 679 532 683
rect 526 678 532 679
rect 270 675 276 676
rect 270 671 271 675
rect 275 671 276 675
rect 270 670 276 671
rect 434 675 440 676
rect 434 671 435 675
rect 439 671 440 675
rect 434 670 440 671
rect 442 675 448 676
rect 442 671 443 675
rect 447 671 448 675
rect 442 670 448 671
rect 506 675 512 676
rect 506 671 507 675
rect 511 671 512 675
rect 506 670 512 671
rect 254 665 260 666
rect 254 661 255 665
rect 259 661 260 665
rect 254 660 260 661
rect 302 665 308 666
rect 302 661 303 665
rect 307 661 308 665
rect 302 660 308 661
rect 358 665 364 666
rect 358 661 359 665
rect 363 661 364 665
rect 358 660 364 661
rect 414 665 420 666
rect 414 661 415 665
rect 419 661 420 665
rect 414 660 420 661
rect 208 651 210 660
rect 222 659 228 660
rect 222 655 223 659
rect 227 655 228 659
rect 222 654 228 655
rect 256 651 258 660
rect 304 651 306 660
rect 360 651 362 660
rect 402 659 408 660
rect 402 655 403 659
rect 407 655 408 659
rect 402 654 408 655
rect 207 650 211 651
rect 207 645 211 646
rect 215 650 219 651
rect 215 645 219 646
rect 255 650 259 651
rect 255 645 259 646
rect 271 650 275 651
rect 271 645 275 646
rect 303 650 307 651
rect 303 645 307 646
rect 327 650 331 651
rect 327 645 331 646
rect 359 650 363 651
rect 359 645 363 646
rect 383 650 387 651
rect 383 645 387 646
rect 178 643 184 644
rect 110 636 111 640
rect 115 636 116 640
rect 110 635 116 636
rect 166 639 172 640
rect 166 635 167 639
rect 171 635 172 639
rect 178 639 179 643
rect 183 639 184 643
rect 216 640 218 645
rect 272 640 274 645
rect 328 640 330 645
rect 338 643 344 644
rect 178 638 184 639
rect 214 639 220 640
rect 166 634 172 635
rect 214 635 215 639
rect 219 635 220 639
rect 214 634 220 635
rect 270 639 276 640
rect 270 635 271 639
rect 275 635 276 639
rect 270 634 276 635
rect 326 639 332 640
rect 326 635 327 639
rect 331 635 332 639
rect 338 639 339 643
rect 343 639 344 643
rect 384 640 386 645
rect 338 638 344 639
rect 382 639 388 640
rect 326 634 332 635
rect 302 627 308 628
rect 110 623 116 624
rect 110 619 111 623
rect 115 619 116 623
rect 302 623 303 627
rect 307 623 308 627
rect 302 622 308 623
rect 110 618 116 619
rect 166 621 172 622
rect 112 615 114 618
rect 166 617 167 621
rect 171 617 172 621
rect 166 616 172 617
rect 214 621 220 622
rect 214 617 215 621
rect 219 617 220 621
rect 214 616 220 617
rect 270 621 276 622
rect 270 617 271 621
rect 275 617 276 621
rect 270 616 276 617
rect 111 614 115 615
rect 111 609 115 610
rect 167 614 171 616
rect 167 609 171 610
rect 215 614 219 616
rect 215 609 219 610
rect 223 614 227 615
rect 112 606 114 609
rect 223 608 227 610
rect 255 614 259 615
rect 255 608 259 610
rect 271 614 275 616
rect 271 609 275 610
rect 287 614 291 615
rect 287 608 291 610
rect 222 607 228 608
rect 110 605 116 606
rect 110 601 111 605
rect 115 601 116 605
rect 222 603 223 607
rect 227 603 228 607
rect 222 602 228 603
rect 254 607 260 608
rect 254 603 255 607
rect 259 603 260 607
rect 254 602 260 603
rect 286 607 292 608
rect 286 603 287 607
rect 291 603 292 607
rect 286 602 292 603
rect 110 600 116 601
rect 210 599 216 600
rect 210 595 211 599
rect 215 595 216 599
rect 210 594 216 595
rect 110 588 116 589
rect 110 584 111 588
rect 115 584 116 588
rect 110 583 116 584
rect 112 579 114 583
rect 111 578 115 579
rect 111 573 115 574
rect 191 578 195 579
rect 191 573 195 574
rect 112 569 114 573
rect 110 568 116 569
rect 192 568 194 573
rect 212 572 214 594
rect 222 589 228 590
rect 222 585 223 589
rect 227 585 228 589
rect 222 584 228 585
rect 254 589 260 590
rect 254 585 255 589
rect 259 585 260 589
rect 254 584 260 585
rect 286 589 292 590
rect 286 585 287 589
rect 291 585 292 589
rect 286 584 292 585
rect 304 584 306 622
rect 326 621 332 622
rect 326 617 327 621
rect 331 617 332 621
rect 326 616 332 617
rect 319 614 323 615
rect 319 608 323 610
rect 327 614 331 616
rect 327 609 331 610
rect 318 607 324 608
rect 318 603 319 607
rect 323 603 324 607
rect 340 604 342 638
rect 382 635 383 639
rect 387 635 388 639
rect 382 634 388 635
rect 404 628 406 654
rect 416 651 418 660
rect 444 652 446 670
rect 470 665 476 666
rect 470 661 471 665
rect 475 661 476 665
rect 470 660 476 661
rect 450 659 456 660
rect 450 655 451 659
rect 455 655 456 659
rect 450 654 456 655
rect 442 651 448 652
rect 415 650 419 651
rect 415 645 419 646
rect 431 650 435 651
rect 442 647 443 651
rect 447 647 448 651
rect 442 646 448 647
rect 431 645 435 646
rect 432 640 434 645
rect 442 643 448 644
rect 430 639 436 640
rect 430 635 431 639
rect 435 635 436 639
rect 442 639 443 643
rect 447 639 448 643
rect 442 638 448 639
rect 430 634 436 635
rect 402 627 408 628
rect 402 623 403 627
rect 407 623 408 627
rect 402 622 408 623
rect 382 621 388 622
rect 382 617 383 621
rect 387 617 388 621
rect 382 616 388 617
rect 430 621 436 622
rect 430 617 431 621
rect 435 617 436 621
rect 430 616 436 617
rect 351 614 355 615
rect 351 608 355 610
rect 383 614 387 616
rect 383 608 387 610
rect 423 614 427 615
rect 423 608 427 610
rect 431 614 435 616
rect 431 609 435 610
rect 350 607 356 608
rect 318 602 324 603
rect 338 603 344 604
rect 338 599 339 603
rect 343 599 344 603
rect 350 603 351 607
rect 355 603 356 607
rect 350 602 356 603
rect 382 607 388 608
rect 382 603 383 607
rect 387 603 388 607
rect 382 602 388 603
rect 422 607 428 608
rect 422 603 423 607
rect 427 603 428 607
rect 422 602 428 603
rect 444 600 446 638
rect 452 628 454 654
rect 472 651 474 660
rect 471 650 475 651
rect 471 645 475 646
rect 487 650 491 651
rect 487 645 491 646
rect 488 640 490 645
rect 508 644 510 670
rect 526 665 532 666
rect 526 661 527 665
rect 531 661 532 665
rect 526 660 532 661
rect 536 660 538 698
rect 542 697 548 698
rect 542 693 543 697
rect 547 693 548 697
rect 542 692 548 693
rect 614 697 620 698
rect 614 693 615 697
rect 619 693 620 697
rect 614 692 620 693
rect 543 690 547 692
rect 543 685 547 686
rect 583 690 587 691
rect 583 684 587 686
rect 615 690 619 692
rect 615 685 619 686
rect 639 690 643 691
rect 639 684 643 686
rect 582 683 588 684
rect 582 679 583 683
rect 587 679 588 683
rect 582 678 588 679
rect 638 683 644 684
rect 638 679 639 683
rect 643 679 644 683
rect 638 678 644 679
rect 660 676 662 718
rect 688 716 690 721
rect 760 716 762 721
rect 766 719 767 723
rect 771 719 772 723
rect 775 721 779 722
rect 839 721 843 722
rect 847 726 851 727
rect 847 721 851 722
rect 919 726 923 727
rect 919 721 923 722
rect 991 726 995 727
rect 991 721 995 722
rect 1007 726 1011 727
rect 1022 726 1028 727
rect 1063 726 1067 727
rect 1078 726 1084 727
rect 1087 726 1091 727
rect 1007 721 1011 722
rect 766 718 772 719
rect 840 716 842 721
rect 854 719 860 720
rect 686 715 692 716
rect 686 711 687 715
rect 691 711 692 715
rect 686 710 692 711
rect 758 715 764 716
rect 758 711 759 715
rect 763 711 764 715
rect 758 710 764 711
rect 838 715 844 716
rect 838 711 839 715
rect 843 711 844 715
rect 854 715 855 719
rect 859 715 860 719
rect 920 716 922 721
rect 1008 716 1010 721
rect 854 714 860 715
rect 918 715 924 716
rect 838 710 844 711
rect 714 707 720 708
rect 714 703 715 707
rect 719 703 720 707
rect 714 702 720 703
rect 686 697 692 698
rect 686 693 687 697
rect 691 693 692 697
rect 686 692 692 693
rect 687 690 691 692
rect 687 685 691 686
rect 695 690 699 691
rect 695 684 699 686
rect 694 683 700 684
rect 694 679 695 683
rect 699 679 700 683
rect 694 678 700 679
rect 658 675 664 676
rect 658 671 659 675
rect 663 671 664 675
rect 658 670 664 671
rect 582 665 588 666
rect 582 661 583 665
rect 587 661 588 665
rect 582 660 588 661
rect 638 665 644 666
rect 638 661 639 665
rect 643 661 644 665
rect 638 660 644 661
rect 694 665 700 666
rect 694 661 695 665
rect 699 661 700 665
rect 694 660 700 661
rect 716 660 718 702
rect 758 697 764 698
rect 758 693 759 697
rect 763 693 764 697
rect 758 692 764 693
rect 838 697 844 698
rect 838 693 839 697
rect 843 693 844 697
rect 838 692 844 693
rect 759 690 763 692
rect 759 684 763 686
rect 823 690 827 691
rect 823 684 827 686
rect 839 690 843 692
rect 839 685 843 686
rect 758 683 764 684
rect 758 679 759 683
rect 763 679 764 683
rect 758 678 764 679
rect 822 683 828 684
rect 822 679 823 683
rect 827 679 828 683
rect 822 678 828 679
rect 856 676 858 714
rect 918 711 919 715
rect 923 711 924 715
rect 918 710 924 711
rect 1006 715 1012 716
rect 1006 711 1007 715
rect 1011 711 1012 715
rect 1006 710 1012 711
rect 1024 704 1026 726
rect 1063 721 1067 722
rect 1087 721 1091 722
rect 1135 726 1139 727
rect 1135 721 1139 722
rect 1167 726 1171 727
rect 1167 721 1171 722
rect 1088 716 1090 721
rect 1168 716 1170 721
rect 1188 720 1190 742
rect 1206 737 1212 738
rect 1206 733 1207 737
rect 1211 733 1212 737
rect 1206 732 1212 733
rect 1270 737 1276 738
rect 1270 733 1271 737
rect 1275 733 1276 737
rect 1270 732 1276 733
rect 1292 732 1294 758
rect 1319 757 1323 758
rect 1327 762 1331 763
rect 1327 756 1331 758
rect 1375 762 1379 763
rect 1375 756 1379 758
rect 1383 762 1387 764
rect 1584 763 1586 766
rect 1383 757 1387 758
rect 1423 762 1427 763
rect 1423 756 1427 758
rect 1471 762 1475 763
rect 1471 756 1475 758
rect 1511 762 1515 763
rect 1511 756 1515 758
rect 1543 762 1547 763
rect 1543 756 1547 758
rect 1583 762 1587 763
rect 1583 757 1587 758
rect 1326 755 1332 756
rect 1326 751 1327 755
rect 1331 751 1332 755
rect 1326 750 1332 751
rect 1374 755 1380 756
rect 1374 751 1375 755
rect 1379 751 1380 755
rect 1374 750 1380 751
rect 1422 755 1428 756
rect 1422 751 1423 755
rect 1427 751 1428 755
rect 1422 750 1428 751
rect 1470 755 1476 756
rect 1470 751 1471 755
rect 1475 751 1476 755
rect 1470 750 1476 751
rect 1510 755 1516 756
rect 1510 751 1511 755
rect 1515 751 1516 755
rect 1510 750 1516 751
rect 1542 755 1548 756
rect 1542 751 1543 755
rect 1547 751 1548 755
rect 1584 754 1586 757
rect 1542 750 1548 751
rect 1582 753 1588 754
rect 1582 749 1583 753
rect 1587 749 1588 753
rect 1582 748 1588 749
rect 1558 747 1564 748
rect 1558 743 1559 747
rect 1563 743 1564 747
rect 1558 742 1564 743
rect 1326 737 1332 738
rect 1326 733 1327 737
rect 1331 733 1332 737
rect 1326 732 1332 733
rect 1374 737 1380 738
rect 1374 733 1375 737
rect 1379 733 1380 737
rect 1374 732 1380 733
rect 1422 737 1428 738
rect 1422 733 1423 737
rect 1427 733 1428 737
rect 1422 732 1428 733
rect 1470 737 1476 738
rect 1470 733 1471 737
rect 1475 733 1476 737
rect 1470 732 1476 733
rect 1510 737 1516 738
rect 1510 733 1511 737
rect 1515 733 1516 737
rect 1510 732 1516 733
rect 1542 737 1548 738
rect 1542 733 1543 737
rect 1547 733 1548 737
rect 1542 732 1548 733
rect 1208 727 1210 732
rect 1272 727 1274 732
rect 1290 731 1296 732
rect 1290 727 1291 731
rect 1295 727 1296 731
rect 1328 727 1330 732
rect 1376 727 1378 732
rect 1424 727 1426 732
rect 1472 727 1474 732
rect 1512 727 1514 732
rect 1544 727 1546 732
rect 1207 726 1211 727
rect 1207 721 1211 722
rect 1239 726 1243 727
rect 1239 721 1243 722
rect 1271 726 1275 727
rect 1290 726 1296 727
rect 1303 726 1307 727
rect 1271 721 1275 722
rect 1303 721 1307 722
rect 1327 726 1331 727
rect 1327 721 1331 722
rect 1359 726 1363 727
rect 1359 721 1363 722
rect 1375 726 1379 727
rect 1375 721 1379 722
rect 1407 726 1411 727
rect 1407 721 1411 722
rect 1423 726 1427 727
rect 1423 721 1427 722
rect 1455 726 1459 727
rect 1455 721 1459 722
rect 1471 726 1475 727
rect 1471 721 1475 722
rect 1511 726 1515 727
rect 1511 721 1515 722
rect 1543 726 1547 727
rect 1543 721 1547 722
rect 1186 719 1192 720
rect 1086 715 1092 716
rect 1086 711 1087 715
rect 1091 711 1092 715
rect 1086 710 1092 711
rect 1166 715 1172 716
rect 1166 711 1167 715
rect 1171 711 1172 715
rect 1186 715 1187 719
rect 1191 715 1192 719
rect 1240 716 1242 721
rect 1294 719 1300 720
rect 1186 714 1192 715
rect 1238 715 1244 716
rect 1166 710 1172 711
rect 1238 711 1239 715
rect 1243 711 1244 715
rect 1294 715 1295 719
rect 1299 715 1300 719
rect 1304 716 1306 721
rect 1360 716 1362 721
rect 1408 716 1410 721
rect 1456 716 1458 721
rect 1512 716 1514 721
rect 1544 716 1546 721
rect 1560 720 1562 742
rect 1582 736 1588 737
rect 1582 732 1583 736
rect 1587 732 1588 736
rect 1582 731 1588 732
rect 1584 727 1586 731
rect 1583 726 1587 727
rect 1583 721 1587 722
rect 1558 719 1564 720
rect 1294 714 1300 715
rect 1302 715 1308 716
rect 1238 710 1244 711
rect 1034 707 1040 708
rect 1022 703 1028 704
rect 1022 699 1023 703
rect 1027 699 1028 703
rect 1034 703 1035 707
rect 1039 703 1040 707
rect 1034 702 1040 703
rect 1022 698 1028 699
rect 918 697 924 698
rect 918 693 919 697
rect 923 693 924 697
rect 918 692 924 693
rect 1006 697 1012 698
rect 1006 693 1007 697
rect 1011 693 1012 697
rect 1006 692 1012 693
rect 887 690 891 691
rect 887 684 891 686
rect 919 690 923 692
rect 919 685 923 686
rect 951 690 955 691
rect 951 684 955 686
rect 1007 690 1011 692
rect 1007 685 1011 686
rect 1015 690 1019 691
rect 1015 684 1019 686
rect 886 683 892 684
rect 886 679 887 683
rect 891 679 892 683
rect 886 678 892 679
rect 950 683 956 684
rect 950 679 951 683
rect 955 679 956 683
rect 950 678 956 679
rect 1014 683 1020 684
rect 1014 679 1015 683
rect 1019 679 1020 683
rect 1014 678 1020 679
rect 774 675 780 676
rect 774 671 775 675
rect 779 671 780 675
rect 774 670 780 671
rect 854 675 860 676
rect 854 671 855 675
rect 859 671 860 675
rect 854 670 860 671
rect 758 665 764 666
rect 758 661 759 665
rect 763 661 764 665
rect 758 660 764 661
rect 528 651 530 660
rect 534 659 540 660
rect 534 655 535 659
rect 539 655 540 659
rect 534 654 540 655
rect 584 651 586 660
rect 602 659 608 660
rect 602 655 603 659
rect 607 655 608 659
rect 602 654 608 655
rect 527 650 531 651
rect 527 645 531 646
rect 535 650 539 651
rect 535 645 539 646
rect 583 650 587 651
rect 583 645 587 646
rect 591 650 595 651
rect 591 645 595 646
rect 506 643 512 644
rect 486 639 492 640
rect 486 635 487 639
rect 491 635 492 639
rect 506 639 507 643
rect 511 639 512 643
rect 536 640 538 645
rect 592 640 594 645
rect 506 638 512 639
rect 534 639 540 640
rect 486 634 492 635
rect 534 635 535 639
rect 539 635 540 639
rect 534 634 540 635
rect 590 639 596 640
rect 590 635 591 639
rect 595 635 596 639
rect 590 634 596 635
rect 604 628 606 654
rect 640 651 642 660
rect 696 651 698 660
rect 714 659 720 660
rect 714 655 715 659
rect 719 655 720 659
rect 714 654 720 655
rect 760 651 762 660
rect 639 650 643 651
rect 639 645 643 646
rect 647 650 651 651
rect 647 645 651 646
rect 695 650 699 651
rect 695 645 699 646
rect 703 650 707 651
rect 703 645 707 646
rect 759 650 763 651
rect 759 645 763 646
rect 648 640 650 645
rect 704 640 706 645
rect 760 640 762 645
rect 776 644 778 670
rect 822 665 828 666
rect 822 661 823 665
rect 827 661 828 665
rect 822 660 828 661
rect 886 665 892 666
rect 886 661 887 665
rect 891 661 892 665
rect 886 660 892 661
rect 950 665 956 666
rect 950 661 951 665
rect 955 661 956 665
rect 950 660 956 661
rect 1014 665 1020 666
rect 1014 661 1015 665
rect 1019 661 1020 665
rect 1014 660 1020 661
rect 1036 660 1038 702
rect 1086 697 1092 698
rect 1086 693 1087 697
rect 1091 693 1092 697
rect 1086 692 1092 693
rect 1166 697 1172 698
rect 1166 693 1167 697
rect 1171 693 1172 697
rect 1166 692 1172 693
rect 1238 697 1244 698
rect 1238 693 1239 697
rect 1243 693 1244 697
rect 1238 692 1244 693
rect 1296 692 1298 714
rect 1302 711 1303 715
rect 1307 711 1308 715
rect 1302 710 1308 711
rect 1358 715 1364 716
rect 1358 711 1359 715
rect 1363 711 1364 715
rect 1358 710 1364 711
rect 1406 715 1412 716
rect 1406 711 1407 715
rect 1411 711 1412 715
rect 1406 710 1412 711
rect 1454 715 1460 716
rect 1454 711 1455 715
rect 1459 711 1460 715
rect 1454 710 1460 711
rect 1510 715 1516 716
rect 1510 711 1511 715
rect 1515 711 1516 715
rect 1510 710 1516 711
rect 1542 715 1548 716
rect 1542 711 1543 715
rect 1547 711 1548 715
rect 1558 715 1559 719
rect 1563 715 1564 719
rect 1584 717 1586 721
rect 1558 714 1564 715
rect 1582 716 1588 717
rect 1582 712 1583 716
rect 1587 712 1588 716
rect 1582 711 1588 712
rect 1542 710 1548 711
rect 1350 703 1356 704
rect 1350 699 1351 703
rect 1355 699 1356 703
rect 1350 698 1356 699
rect 1582 699 1588 700
rect 1302 697 1308 698
rect 1302 693 1303 697
rect 1307 693 1308 697
rect 1302 692 1308 693
rect 1079 690 1083 691
rect 1079 684 1083 686
rect 1087 690 1091 692
rect 1087 685 1091 686
rect 1135 690 1139 691
rect 1135 684 1139 686
rect 1167 690 1171 692
rect 1167 685 1171 686
rect 1191 690 1195 691
rect 1191 684 1195 686
rect 1239 690 1243 692
rect 1294 691 1300 692
rect 1239 685 1243 686
rect 1247 690 1251 691
rect 1294 687 1295 691
rect 1299 687 1300 691
rect 1294 686 1300 687
rect 1303 690 1307 692
rect 1247 684 1251 686
rect 1303 684 1307 686
rect 1078 683 1084 684
rect 1078 679 1079 683
rect 1083 679 1084 683
rect 1078 678 1084 679
rect 1134 683 1140 684
rect 1134 679 1135 683
rect 1139 679 1140 683
rect 1134 678 1140 679
rect 1190 683 1196 684
rect 1190 679 1191 683
rect 1195 679 1196 683
rect 1190 678 1196 679
rect 1246 683 1252 684
rect 1246 679 1247 683
rect 1251 679 1252 683
rect 1246 678 1252 679
rect 1302 683 1308 684
rect 1302 679 1303 683
rect 1307 679 1308 683
rect 1302 678 1308 679
rect 1126 675 1132 676
rect 1126 671 1127 675
rect 1131 671 1132 675
rect 1126 670 1132 671
rect 1182 675 1188 676
rect 1182 671 1183 675
rect 1187 671 1188 675
rect 1182 670 1188 671
rect 1078 665 1084 666
rect 1078 661 1079 665
rect 1083 661 1084 665
rect 1078 660 1084 661
rect 824 651 826 660
rect 888 651 890 660
rect 906 651 912 652
rect 952 651 954 660
rect 1016 651 1018 660
rect 1034 659 1040 660
rect 1034 655 1035 659
rect 1039 655 1040 659
rect 1034 654 1040 655
rect 1080 651 1082 660
rect 823 650 827 651
rect 823 645 827 646
rect 887 650 891 651
rect 906 647 907 651
rect 911 647 912 651
rect 906 646 912 647
rect 943 650 947 651
rect 887 645 891 646
rect 774 643 780 644
rect 646 639 652 640
rect 646 635 647 639
rect 651 635 652 639
rect 646 634 652 635
rect 702 639 708 640
rect 702 635 703 639
rect 707 635 708 639
rect 702 634 708 635
rect 758 639 764 640
rect 758 635 759 639
rect 763 635 764 639
rect 774 639 775 643
rect 779 639 780 643
rect 824 640 826 645
rect 834 643 840 644
rect 774 638 780 639
rect 822 639 828 640
rect 758 634 764 635
rect 822 635 823 639
rect 827 635 828 639
rect 834 639 835 643
rect 839 639 840 643
rect 888 640 890 645
rect 834 638 840 639
rect 886 639 892 640
rect 822 634 828 635
rect 450 627 456 628
rect 450 623 451 627
rect 455 623 456 627
rect 450 622 456 623
rect 574 627 580 628
rect 574 623 575 627
rect 579 623 580 627
rect 574 622 580 623
rect 602 627 608 628
rect 602 623 603 627
rect 607 623 608 627
rect 602 622 608 623
rect 486 621 492 622
rect 486 617 487 621
rect 491 617 492 621
rect 486 616 492 617
rect 534 621 540 622
rect 534 617 535 621
rect 539 617 540 621
rect 534 616 540 617
rect 463 614 467 615
rect 463 608 467 610
rect 487 614 491 616
rect 487 609 491 610
rect 519 614 523 615
rect 519 608 523 610
rect 535 614 539 616
rect 535 609 539 610
rect 462 607 468 608
rect 462 603 463 607
rect 467 603 468 607
rect 462 602 468 603
rect 518 607 524 608
rect 518 603 519 607
rect 523 603 524 607
rect 518 602 524 603
rect 338 598 344 599
rect 442 599 448 600
rect 442 595 443 599
rect 447 595 448 599
rect 442 594 448 595
rect 318 589 324 590
rect 318 585 319 589
rect 323 585 324 589
rect 318 584 324 585
rect 350 589 356 590
rect 350 585 351 589
rect 355 585 356 589
rect 350 584 356 585
rect 382 589 388 590
rect 382 585 383 589
rect 387 585 388 589
rect 382 584 388 585
rect 422 589 428 590
rect 422 585 423 589
rect 427 585 428 589
rect 422 584 428 585
rect 462 589 468 590
rect 462 585 463 589
rect 467 585 468 589
rect 462 584 468 585
rect 518 589 524 590
rect 518 585 519 589
rect 523 585 524 589
rect 518 584 524 585
rect 576 584 578 622
rect 590 621 596 622
rect 590 617 591 621
rect 595 617 596 621
rect 590 616 596 617
rect 646 621 652 622
rect 646 617 647 621
rect 651 617 652 621
rect 646 616 652 617
rect 702 621 708 622
rect 702 617 703 621
rect 707 617 708 621
rect 702 616 708 617
rect 758 621 764 622
rect 758 617 759 621
rect 763 617 764 621
rect 758 616 764 617
rect 822 621 828 622
rect 822 617 823 621
rect 827 617 828 621
rect 822 616 828 617
rect 583 614 587 615
rect 583 608 587 610
rect 591 614 595 616
rect 591 609 595 610
rect 647 614 651 616
rect 647 608 651 610
rect 703 614 707 616
rect 703 609 707 610
rect 719 614 723 615
rect 719 608 723 610
rect 759 614 763 616
rect 759 609 763 610
rect 799 614 803 615
rect 799 608 803 610
rect 823 614 827 616
rect 823 609 827 610
rect 582 607 588 608
rect 582 603 583 607
rect 587 603 588 607
rect 582 602 588 603
rect 646 607 652 608
rect 646 603 647 607
rect 651 603 652 607
rect 646 602 652 603
rect 718 607 724 608
rect 718 603 719 607
rect 723 603 724 607
rect 718 602 724 603
rect 798 607 804 608
rect 798 603 799 607
rect 803 603 804 607
rect 798 602 804 603
rect 836 600 838 638
rect 886 635 887 639
rect 891 635 892 639
rect 886 634 892 635
rect 908 628 910 646
rect 943 645 947 646
rect 951 650 955 651
rect 951 645 955 646
rect 999 650 1003 651
rect 999 645 1003 646
rect 1015 650 1019 651
rect 1015 645 1019 646
rect 1055 650 1059 651
rect 1055 645 1059 646
rect 1079 650 1083 651
rect 1079 645 1083 646
rect 1111 650 1115 651
rect 1111 645 1115 646
rect 944 640 946 645
rect 1000 640 1002 645
rect 1056 640 1058 645
rect 1112 640 1114 645
rect 1128 644 1130 670
rect 1134 665 1140 666
rect 1134 661 1135 665
rect 1139 661 1140 665
rect 1134 660 1140 661
rect 1136 651 1138 660
rect 1135 650 1139 651
rect 1135 645 1139 646
rect 1167 650 1171 651
rect 1167 645 1171 646
rect 1126 643 1132 644
rect 942 639 948 640
rect 942 635 943 639
rect 947 635 948 639
rect 942 634 948 635
rect 998 639 1004 640
rect 998 635 999 639
rect 1003 635 1004 639
rect 998 634 1004 635
rect 1054 639 1060 640
rect 1054 635 1055 639
rect 1059 635 1060 639
rect 1054 634 1060 635
rect 1110 639 1116 640
rect 1110 635 1111 639
rect 1115 635 1116 639
rect 1126 639 1127 643
rect 1131 639 1132 643
rect 1168 640 1170 645
rect 1184 644 1186 670
rect 1190 665 1196 666
rect 1190 661 1191 665
rect 1195 661 1196 665
rect 1190 660 1196 661
rect 1246 665 1252 666
rect 1246 661 1247 665
rect 1251 661 1252 665
rect 1246 660 1252 661
rect 1302 665 1308 666
rect 1302 661 1303 665
rect 1307 661 1308 665
rect 1302 660 1308 661
rect 1352 660 1354 698
rect 1358 697 1364 698
rect 1358 693 1359 697
rect 1363 693 1364 697
rect 1358 692 1364 693
rect 1406 697 1412 698
rect 1406 693 1407 697
rect 1411 693 1412 697
rect 1406 692 1412 693
rect 1454 697 1460 698
rect 1454 693 1455 697
rect 1459 693 1460 697
rect 1454 692 1460 693
rect 1510 697 1516 698
rect 1510 693 1511 697
rect 1515 693 1516 697
rect 1510 692 1516 693
rect 1542 697 1548 698
rect 1542 693 1543 697
rect 1547 693 1548 697
rect 1582 695 1583 699
rect 1587 695 1588 699
rect 1582 694 1588 695
rect 1542 692 1548 693
rect 1359 690 1363 692
rect 1359 684 1363 686
rect 1407 690 1411 692
rect 1407 685 1411 686
rect 1455 690 1459 692
rect 1455 685 1459 686
rect 1511 690 1515 692
rect 1511 685 1515 686
rect 1543 690 1547 692
rect 1584 691 1586 694
rect 1543 685 1547 686
rect 1583 690 1587 691
rect 1583 685 1587 686
rect 1358 683 1364 684
rect 1358 679 1359 683
rect 1363 679 1364 683
rect 1584 682 1586 685
rect 1358 678 1364 679
rect 1582 681 1588 682
rect 1582 677 1583 681
rect 1587 677 1588 681
rect 1582 676 1588 677
rect 1358 665 1364 666
rect 1358 661 1359 665
rect 1363 661 1364 665
rect 1358 660 1364 661
rect 1582 664 1588 665
rect 1582 660 1583 664
rect 1587 660 1588 664
rect 1192 651 1194 660
rect 1248 651 1250 660
rect 1304 651 1306 660
rect 1350 659 1356 660
rect 1350 655 1351 659
rect 1355 655 1356 659
rect 1350 654 1356 655
rect 1360 651 1362 660
rect 1582 659 1588 660
rect 1584 651 1586 659
rect 1191 650 1195 651
rect 1191 645 1195 646
rect 1215 650 1219 651
rect 1215 645 1219 646
rect 1247 650 1251 651
rect 1247 645 1251 646
rect 1271 650 1275 651
rect 1271 645 1275 646
rect 1303 650 1307 651
rect 1303 645 1307 646
rect 1327 650 1331 651
rect 1327 645 1331 646
rect 1359 650 1363 651
rect 1359 645 1363 646
rect 1383 650 1387 651
rect 1383 645 1387 646
rect 1439 650 1443 651
rect 1439 645 1443 646
rect 1503 650 1507 651
rect 1503 645 1507 646
rect 1543 650 1547 651
rect 1543 645 1547 646
rect 1583 650 1587 651
rect 1583 645 1587 646
rect 1182 643 1188 644
rect 1126 638 1132 639
rect 1166 639 1172 640
rect 1110 634 1116 635
rect 1166 635 1167 639
rect 1171 635 1172 639
rect 1182 639 1183 643
rect 1187 639 1188 643
rect 1216 640 1218 645
rect 1272 640 1274 645
rect 1328 640 1330 645
rect 1384 640 1386 645
rect 1440 640 1442 645
rect 1504 640 1506 645
rect 1522 643 1528 644
rect 1182 638 1188 639
rect 1214 639 1220 640
rect 1166 634 1172 635
rect 1214 635 1215 639
rect 1219 635 1220 639
rect 1214 634 1220 635
rect 1270 639 1276 640
rect 1270 635 1271 639
rect 1275 635 1276 639
rect 1270 634 1276 635
rect 1326 639 1332 640
rect 1326 635 1327 639
rect 1331 635 1332 639
rect 1326 634 1332 635
rect 1382 639 1388 640
rect 1382 635 1383 639
rect 1387 635 1388 639
rect 1382 634 1388 635
rect 1438 639 1444 640
rect 1438 635 1439 639
rect 1443 635 1444 639
rect 1438 634 1444 635
rect 1502 639 1508 640
rect 1502 635 1503 639
rect 1507 635 1508 639
rect 1522 639 1523 643
rect 1527 639 1528 643
rect 1544 640 1546 645
rect 1584 641 1586 645
rect 1582 640 1588 641
rect 1522 638 1528 639
rect 1542 639 1548 640
rect 1502 634 1508 635
rect 906 627 912 628
rect 906 623 907 627
rect 911 623 912 627
rect 906 622 912 623
rect 990 627 996 628
rect 990 623 991 627
rect 995 623 996 627
rect 990 622 996 623
rect 886 621 892 622
rect 886 617 887 621
rect 891 617 892 621
rect 886 616 892 617
rect 942 621 948 622
rect 942 617 943 621
rect 947 617 948 621
rect 942 616 948 617
rect 887 614 891 616
rect 887 608 891 610
rect 943 614 947 616
rect 943 609 947 610
rect 975 614 979 615
rect 975 608 979 610
rect 886 607 892 608
rect 886 603 887 607
rect 891 603 892 607
rect 886 602 892 603
rect 974 607 980 608
rect 974 603 975 607
rect 979 603 980 607
rect 974 602 980 603
rect 834 599 840 600
rect 834 595 835 599
rect 839 595 840 599
rect 834 594 840 595
rect 846 599 852 600
rect 846 595 847 599
rect 851 595 852 599
rect 846 594 852 595
rect 582 589 588 590
rect 582 585 583 589
rect 587 585 588 589
rect 582 584 588 585
rect 646 589 652 590
rect 646 585 647 589
rect 651 585 652 589
rect 646 584 652 585
rect 718 589 724 590
rect 718 585 719 589
rect 723 585 724 589
rect 718 584 724 585
rect 798 589 804 590
rect 798 585 799 589
rect 803 585 804 589
rect 798 584 804 585
rect 224 579 226 584
rect 256 579 258 584
rect 288 579 290 584
rect 302 583 308 584
rect 302 579 303 583
rect 307 579 308 583
rect 320 579 322 584
rect 352 579 354 584
rect 384 579 386 584
rect 414 583 420 584
rect 414 579 415 583
rect 419 579 420 583
rect 424 579 426 584
rect 464 579 466 584
rect 520 579 522 584
rect 574 583 580 584
rect 574 579 575 583
rect 579 579 580 583
rect 584 579 586 584
rect 648 579 650 584
rect 720 579 722 584
rect 800 579 802 584
rect 848 580 850 594
rect 886 589 892 590
rect 886 585 887 589
rect 891 585 892 589
rect 886 584 892 585
rect 974 589 980 590
rect 974 585 975 589
rect 979 585 980 589
rect 974 584 980 585
rect 992 584 994 622
rect 998 621 1004 622
rect 998 617 999 621
rect 1003 617 1004 621
rect 998 616 1004 617
rect 1054 621 1060 622
rect 1054 617 1055 621
rect 1059 617 1060 621
rect 1054 616 1060 617
rect 1110 621 1116 622
rect 1110 617 1111 621
rect 1115 617 1116 621
rect 1110 616 1116 617
rect 1166 621 1172 622
rect 1166 617 1167 621
rect 1171 617 1172 621
rect 1166 616 1172 617
rect 1214 621 1220 622
rect 1214 617 1215 621
rect 1219 617 1220 621
rect 1214 616 1220 617
rect 1270 621 1276 622
rect 1270 617 1271 621
rect 1275 617 1276 621
rect 1270 616 1276 617
rect 1326 621 1332 622
rect 1326 617 1327 621
rect 1331 617 1332 621
rect 1326 616 1332 617
rect 1382 621 1388 622
rect 1382 617 1383 621
rect 1387 617 1388 621
rect 1382 616 1388 617
rect 1438 621 1444 622
rect 1438 617 1439 621
rect 1443 617 1444 621
rect 1438 616 1444 617
rect 1502 621 1508 622
rect 1502 617 1503 621
rect 1507 617 1508 621
rect 1502 616 1508 617
rect 999 614 1003 616
rect 999 609 1003 610
rect 1055 614 1059 616
rect 1055 609 1059 610
rect 1063 614 1067 615
rect 1063 608 1067 610
rect 1111 614 1115 616
rect 1111 609 1115 610
rect 1143 614 1147 615
rect 1143 608 1147 610
rect 1167 614 1171 616
rect 1167 609 1171 610
rect 1215 614 1219 616
rect 1230 615 1236 616
rect 1230 611 1231 615
rect 1235 611 1236 615
rect 1230 610 1236 611
rect 1271 614 1275 616
rect 1215 608 1219 610
rect 1062 607 1068 608
rect 1062 603 1063 607
rect 1067 603 1068 607
rect 1062 602 1068 603
rect 1142 607 1148 608
rect 1142 603 1143 607
rect 1147 603 1148 607
rect 1142 602 1148 603
rect 1214 607 1220 608
rect 1214 603 1215 607
rect 1219 603 1220 607
rect 1214 602 1220 603
rect 1182 599 1188 600
rect 1182 595 1183 599
rect 1187 595 1188 599
rect 1182 594 1188 595
rect 1062 589 1068 590
rect 1062 585 1063 589
rect 1067 585 1068 589
rect 1062 584 1068 585
rect 1142 589 1148 590
rect 1142 585 1143 589
rect 1147 585 1148 589
rect 1142 584 1148 585
rect 846 579 852 580
rect 888 579 890 584
rect 976 579 978 584
rect 990 583 996 584
rect 990 579 991 583
rect 995 579 996 583
rect 1064 579 1066 584
rect 1144 579 1146 584
rect 223 578 227 579
rect 223 573 227 574
rect 255 578 259 579
rect 255 573 259 574
rect 287 578 291 579
rect 302 578 308 579
rect 319 578 323 579
rect 287 573 291 574
rect 319 573 323 574
rect 327 578 331 579
rect 327 573 331 574
rect 351 578 355 579
rect 351 573 355 574
rect 383 578 387 579
rect 383 573 387 574
rect 399 578 403 579
rect 414 578 420 579
rect 423 578 427 579
rect 399 573 403 574
rect 210 571 216 572
rect 110 564 111 568
rect 115 564 116 568
rect 110 563 116 564
rect 190 567 196 568
rect 190 563 191 567
rect 195 563 196 567
rect 210 567 211 571
rect 215 567 216 571
rect 256 568 258 573
rect 328 568 330 573
rect 400 568 402 573
rect 210 566 216 567
rect 254 567 260 568
rect 190 562 196 563
rect 254 563 255 567
rect 259 563 260 567
rect 254 562 260 563
rect 326 567 332 568
rect 326 563 327 567
rect 331 563 332 567
rect 326 562 332 563
rect 398 567 404 568
rect 398 563 399 567
rect 403 563 404 567
rect 398 562 404 563
rect 416 556 418 578
rect 423 573 427 574
rect 463 578 467 579
rect 463 573 467 574
rect 471 578 475 579
rect 471 573 475 574
rect 519 578 523 579
rect 519 573 523 574
rect 535 578 539 579
rect 574 578 580 579
rect 583 578 587 579
rect 535 573 539 574
rect 583 573 587 574
rect 599 578 603 579
rect 599 573 603 574
rect 647 578 651 579
rect 647 573 651 574
rect 663 578 667 579
rect 663 573 667 574
rect 719 578 723 579
rect 719 573 723 574
rect 727 578 731 579
rect 727 573 731 574
rect 783 578 787 579
rect 783 573 787 574
rect 799 578 803 579
rect 799 573 803 574
rect 839 578 843 579
rect 846 575 847 579
rect 851 575 852 579
rect 846 574 852 575
rect 887 578 891 579
rect 839 573 843 574
rect 887 573 891 574
rect 903 578 907 579
rect 903 573 907 574
rect 967 578 971 579
rect 967 573 971 574
rect 975 578 979 579
rect 990 578 996 579
rect 1039 578 1043 579
rect 975 573 979 574
rect 1039 573 1043 574
rect 1063 578 1067 579
rect 1063 573 1067 574
rect 1103 578 1107 579
rect 1103 573 1107 574
rect 1143 578 1147 579
rect 1143 573 1147 574
rect 1167 578 1171 579
rect 1167 573 1171 574
rect 472 568 474 573
rect 536 568 538 573
rect 590 571 596 572
rect 470 567 476 568
rect 470 563 471 567
rect 475 563 476 567
rect 470 562 476 563
rect 534 567 540 568
rect 534 563 535 567
rect 539 563 540 567
rect 590 567 591 571
rect 595 567 596 571
rect 600 568 602 573
rect 664 568 666 573
rect 728 568 730 573
rect 784 568 786 573
rect 840 568 842 573
rect 904 568 906 573
rect 968 568 970 573
rect 1040 568 1042 573
rect 1104 568 1106 573
rect 1168 568 1170 573
rect 1184 572 1186 594
rect 1214 589 1220 590
rect 1214 585 1215 589
rect 1219 585 1220 589
rect 1232 588 1234 610
rect 1271 609 1275 610
rect 1287 614 1291 615
rect 1287 608 1291 610
rect 1327 614 1331 616
rect 1327 609 1331 610
rect 1351 614 1355 615
rect 1351 608 1355 610
rect 1383 614 1387 616
rect 1383 609 1387 610
rect 1407 614 1411 615
rect 1407 608 1411 610
rect 1439 614 1443 616
rect 1439 609 1443 610
rect 1455 614 1459 615
rect 1455 608 1459 610
rect 1503 614 1507 616
rect 1503 609 1507 610
rect 1511 614 1515 615
rect 1511 608 1515 610
rect 1286 607 1292 608
rect 1286 603 1287 607
rect 1291 603 1292 607
rect 1286 602 1292 603
rect 1350 607 1356 608
rect 1350 603 1351 607
rect 1355 603 1356 607
rect 1350 602 1356 603
rect 1406 607 1412 608
rect 1406 603 1407 607
rect 1411 603 1412 607
rect 1406 602 1412 603
rect 1454 607 1460 608
rect 1454 603 1455 607
rect 1459 603 1460 607
rect 1454 602 1460 603
rect 1510 607 1516 608
rect 1510 603 1511 607
rect 1515 603 1516 607
rect 1510 602 1516 603
rect 1524 600 1526 638
rect 1542 635 1543 639
rect 1547 635 1548 639
rect 1582 636 1583 640
rect 1587 636 1588 640
rect 1582 635 1588 636
rect 1542 634 1548 635
rect 1558 627 1564 628
rect 1558 623 1559 627
rect 1563 623 1564 627
rect 1558 622 1564 623
rect 1582 623 1588 624
rect 1542 621 1548 622
rect 1542 617 1543 621
rect 1547 617 1548 621
rect 1542 616 1548 617
rect 1543 614 1547 616
rect 1543 608 1547 610
rect 1542 607 1548 608
rect 1542 603 1543 607
rect 1547 603 1548 607
rect 1542 602 1548 603
rect 1486 599 1492 600
rect 1486 595 1487 599
rect 1491 595 1492 599
rect 1486 594 1492 595
rect 1522 599 1528 600
rect 1522 595 1523 599
rect 1527 595 1528 599
rect 1522 594 1528 595
rect 1286 589 1292 590
rect 1214 584 1220 585
rect 1230 587 1236 588
rect 1216 579 1218 584
rect 1230 583 1231 587
rect 1235 583 1236 587
rect 1286 585 1287 589
rect 1291 585 1292 589
rect 1286 584 1292 585
rect 1350 589 1356 590
rect 1350 585 1351 589
rect 1355 585 1356 589
rect 1350 584 1356 585
rect 1406 589 1412 590
rect 1406 585 1407 589
rect 1411 585 1412 589
rect 1406 584 1412 585
rect 1454 589 1460 590
rect 1454 585 1455 589
rect 1459 585 1460 589
rect 1454 584 1460 585
rect 1230 582 1236 583
rect 1288 579 1290 584
rect 1352 579 1354 584
rect 1408 579 1410 584
rect 1456 579 1458 584
rect 1215 578 1219 579
rect 1215 573 1219 574
rect 1231 578 1235 579
rect 1231 573 1235 574
rect 1287 578 1291 579
rect 1287 573 1291 574
rect 1335 578 1339 579
rect 1335 573 1339 574
rect 1351 578 1355 579
rect 1351 573 1355 574
rect 1383 578 1387 579
rect 1383 573 1387 574
rect 1407 578 1411 579
rect 1407 573 1411 574
rect 1423 578 1427 579
rect 1423 573 1427 574
rect 1455 578 1459 579
rect 1455 573 1459 574
rect 1471 578 1475 579
rect 1471 573 1475 574
rect 1182 571 1188 572
rect 590 566 596 567
rect 598 567 604 568
rect 534 562 540 563
rect 338 555 344 556
rect 110 551 116 552
rect 110 547 111 551
rect 115 547 116 551
rect 338 551 339 555
rect 343 551 344 555
rect 338 550 344 551
rect 414 555 420 556
rect 414 551 415 555
rect 419 551 420 555
rect 414 550 420 551
rect 110 546 116 547
rect 190 549 196 550
rect 112 543 114 546
rect 190 545 191 549
rect 195 545 196 549
rect 190 544 196 545
rect 254 549 260 550
rect 254 545 255 549
rect 259 545 260 549
rect 254 544 260 545
rect 326 549 332 550
rect 326 545 327 549
rect 331 545 332 549
rect 326 544 332 545
rect 111 542 115 543
rect 111 537 115 538
rect 135 542 139 543
rect 112 534 114 537
rect 135 536 139 538
rect 175 542 179 543
rect 175 536 179 538
rect 191 542 195 544
rect 191 537 195 538
rect 231 542 235 543
rect 231 536 235 538
rect 255 542 259 544
rect 255 537 259 538
rect 295 542 299 543
rect 295 536 299 538
rect 327 542 331 544
rect 327 537 331 538
rect 134 535 140 536
rect 110 533 116 534
rect 110 529 111 533
rect 115 529 116 533
rect 134 531 135 535
rect 139 531 140 535
rect 134 530 140 531
rect 174 535 180 536
rect 174 531 175 535
rect 179 531 180 535
rect 174 530 180 531
rect 230 535 236 536
rect 230 531 231 535
rect 235 531 236 535
rect 230 530 236 531
rect 294 535 300 536
rect 294 531 295 535
rect 299 531 300 535
rect 294 530 300 531
rect 110 528 116 529
rect 150 527 156 528
rect 150 523 151 527
rect 155 523 156 527
rect 150 522 156 523
rect 134 517 140 518
rect 110 516 116 517
rect 110 512 111 516
rect 115 512 116 516
rect 134 513 135 517
rect 139 513 140 517
rect 134 512 140 513
rect 110 511 116 512
rect 112 507 114 511
rect 136 507 138 512
rect 111 506 115 507
rect 111 501 115 502
rect 135 506 139 507
rect 135 501 139 502
rect 112 497 114 501
rect 110 496 116 497
rect 136 496 138 501
rect 152 500 154 522
rect 174 517 180 518
rect 174 513 175 517
rect 179 513 180 517
rect 174 512 180 513
rect 230 517 236 518
rect 230 513 231 517
rect 235 513 236 517
rect 230 512 236 513
rect 294 517 300 518
rect 294 513 295 517
rect 299 513 300 517
rect 340 516 342 550
rect 398 549 404 550
rect 398 545 399 549
rect 403 545 404 549
rect 398 544 404 545
rect 470 549 476 550
rect 470 545 471 549
rect 475 545 476 549
rect 470 544 476 545
rect 534 549 540 550
rect 534 545 535 549
rect 539 545 540 549
rect 534 544 540 545
rect 592 544 594 566
rect 598 563 599 567
rect 603 563 604 567
rect 598 562 604 563
rect 662 567 668 568
rect 662 563 663 567
rect 667 563 668 567
rect 662 562 668 563
rect 726 567 732 568
rect 726 563 727 567
rect 731 563 732 567
rect 726 562 732 563
rect 782 567 788 568
rect 782 563 783 567
rect 787 563 788 567
rect 782 562 788 563
rect 838 567 844 568
rect 838 563 839 567
rect 843 563 844 567
rect 838 562 844 563
rect 902 567 908 568
rect 902 563 903 567
rect 907 563 908 567
rect 902 562 908 563
rect 966 567 972 568
rect 966 563 967 567
rect 971 563 972 567
rect 966 562 972 563
rect 1038 567 1044 568
rect 1038 563 1039 567
rect 1043 563 1044 567
rect 1038 562 1044 563
rect 1102 567 1108 568
rect 1102 563 1103 567
rect 1107 563 1108 567
rect 1102 562 1108 563
rect 1166 567 1172 568
rect 1166 563 1167 567
rect 1171 563 1172 567
rect 1182 567 1183 571
rect 1187 567 1188 571
rect 1232 568 1234 573
rect 1288 568 1290 573
rect 1336 568 1338 573
rect 1384 568 1386 573
rect 1424 568 1426 573
rect 1472 568 1474 573
rect 1488 572 1490 594
rect 1510 589 1516 590
rect 1510 585 1511 589
rect 1515 585 1516 589
rect 1510 584 1516 585
rect 1542 589 1548 590
rect 1542 585 1543 589
rect 1547 585 1548 589
rect 1542 584 1548 585
rect 1560 584 1562 622
rect 1582 619 1583 623
rect 1587 619 1588 623
rect 1582 618 1588 619
rect 1584 615 1586 618
rect 1583 614 1587 615
rect 1583 609 1587 610
rect 1584 606 1586 609
rect 1582 605 1588 606
rect 1582 601 1583 605
rect 1587 601 1588 605
rect 1582 600 1588 601
rect 1582 588 1588 589
rect 1582 584 1583 588
rect 1587 584 1588 588
rect 1512 579 1514 584
rect 1526 583 1532 584
rect 1526 579 1527 583
rect 1531 579 1532 583
rect 1544 579 1546 584
rect 1558 583 1564 584
rect 1582 583 1588 584
rect 1558 579 1559 583
rect 1563 579 1564 583
rect 1584 579 1586 583
rect 1511 578 1515 579
rect 1526 578 1532 579
rect 1543 578 1547 579
rect 1558 578 1564 579
rect 1583 578 1587 579
rect 1511 573 1515 574
rect 1486 571 1492 572
rect 1182 566 1188 567
rect 1230 567 1236 568
rect 1166 562 1172 563
rect 1230 563 1231 567
rect 1235 563 1236 567
rect 1230 562 1236 563
rect 1286 567 1292 568
rect 1286 563 1287 567
rect 1291 563 1292 567
rect 1286 562 1292 563
rect 1334 567 1340 568
rect 1334 563 1335 567
rect 1339 563 1340 567
rect 1334 562 1340 563
rect 1382 567 1388 568
rect 1382 563 1383 567
rect 1387 563 1388 567
rect 1382 562 1388 563
rect 1422 567 1428 568
rect 1422 563 1423 567
rect 1427 563 1428 567
rect 1422 562 1428 563
rect 1470 567 1476 568
rect 1470 563 1471 567
rect 1475 563 1476 567
rect 1486 567 1487 571
rect 1491 567 1492 571
rect 1512 568 1514 573
rect 1486 566 1492 567
rect 1510 567 1516 568
rect 1470 562 1476 563
rect 1510 563 1511 567
rect 1515 563 1516 567
rect 1510 562 1516 563
rect 1528 556 1530 578
rect 1543 573 1547 574
rect 1550 575 1556 576
rect 1544 568 1546 573
rect 1550 571 1551 575
rect 1555 571 1556 575
rect 1583 573 1587 574
rect 1550 570 1556 571
rect 1542 567 1548 568
rect 1542 563 1543 567
rect 1547 563 1548 567
rect 1542 562 1548 563
rect 1526 555 1532 556
rect 1526 551 1527 555
rect 1531 551 1532 555
rect 1526 550 1532 551
rect 598 549 604 550
rect 598 545 599 549
rect 603 545 604 549
rect 598 544 604 545
rect 662 549 668 550
rect 662 545 663 549
rect 667 545 668 549
rect 662 544 668 545
rect 726 549 732 550
rect 726 545 727 549
rect 731 545 732 549
rect 726 544 732 545
rect 782 549 788 550
rect 782 545 783 549
rect 787 545 788 549
rect 782 544 788 545
rect 838 549 844 550
rect 838 545 839 549
rect 843 545 844 549
rect 838 544 844 545
rect 902 549 908 550
rect 902 545 903 549
rect 907 545 908 549
rect 902 544 908 545
rect 966 549 972 550
rect 966 545 967 549
rect 971 545 972 549
rect 966 544 972 545
rect 1038 549 1044 550
rect 1038 545 1039 549
rect 1043 545 1044 549
rect 1038 544 1044 545
rect 1102 549 1108 550
rect 1102 545 1103 549
rect 1107 545 1108 549
rect 1102 544 1108 545
rect 1166 549 1172 550
rect 1166 545 1167 549
rect 1171 545 1172 549
rect 1166 544 1172 545
rect 1230 549 1236 550
rect 1230 545 1231 549
rect 1235 545 1236 549
rect 1230 544 1236 545
rect 1286 549 1292 550
rect 1286 545 1287 549
rect 1291 545 1292 549
rect 1286 544 1292 545
rect 1334 549 1340 550
rect 1334 545 1335 549
rect 1339 545 1340 549
rect 1334 544 1340 545
rect 1382 549 1388 550
rect 1382 545 1383 549
rect 1387 545 1388 549
rect 1382 544 1388 545
rect 1422 549 1428 550
rect 1422 545 1423 549
rect 1427 545 1428 549
rect 1422 544 1428 545
rect 1470 549 1476 550
rect 1470 545 1471 549
rect 1475 545 1476 549
rect 1470 544 1476 545
rect 1510 549 1516 550
rect 1510 545 1511 549
rect 1515 545 1516 549
rect 1510 544 1516 545
rect 1542 549 1548 550
rect 1542 545 1543 549
rect 1547 545 1548 549
rect 1542 544 1548 545
rect 359 542 363 543
rect 359 536 363 538
rect 399 542 403 544
rect 399 537 403 538
rect 423 542 427 543
rect 423 536 427 538
rect 471 542 475 544
rect 471 537 475 538
rect 479 542 483 543
rect 479 536 483 538
rect 535 542 539 544
rect 590 543 596 544
rect 535 537 539 538
rect 543 542 547 543
rect 590 539 591 543
rect 595 539 596 543
rect 590 538 596 539
rect 599 542 603 544
rect 543 536 547 538
rect 599 536 603 538
rect 655 542 659 543
rect 655 536 659 538
rect 663 542 667 544
rect 663 537 667 538
rect 711 542 715 543
rect 711 536 715 538
rect 727 542 731 544
rect 727 537 731 538
rect 767 542 771 543
rect 767 536 771 538
rect 783 542 787 544
rect 783 537 787 538
rect 831 542 835 543
rect 831 536 835 538
rect 839 542 843 544
rect 839 537 843 538
rect 895 542 899 543
rect 895 536 899 538
rect 903 542 907 544
rect 910 543 916 544
rect 910 539 911 543
rect 915 539 916 543
rect 910 538 916 539
rect 967 542 971 544
rect 903 537 907 538
rect 358 535 364 536
rect 358 531 359 535
rect 363 531 364 535
rect 358 530 364 531
rect 422 535 428 536
rect 422 531 423 535
rect 427 531 428 535
rect 422 530 428 531
rect 478 535 484 536
rect 478 531 479 535
rect 483 531 484 535
rect 478 530 484 531
rect 542 535 548 536
rect 542 531 543 535
rect 547 531 548 535
rect 542 530 548 531
rect 598 535 604 536
rect 598 531 599 535
rect 603 531 604 535
rect 598 530 604 531
rect 654 535 660 536
rect 654 531 655 535
rect 659 531 660 535
rect 654 530 660 531
rect 710 535 716 536
rect 710 531 711 535
rect 715 531 716 535
rect 710 530 716 531
rect 766 535 772 536
rect 766 531 767 535
rect 771 531 772 535
rect 766 530 772 531
rect 830 535 836 536
rect 830 531 831 535
rect 835 531 836 535
rect 830 530 836 531
rect 894 535 900 536
rect 894 531 895 535
rect 899 531 900 535
rect 894 530 900 531
rect 358 517 364 518
rect 294 512 300 513
rect 338 515 344 516
rect 176 507 178 512
rect 232 507 234 512
rect 296 507 298 512
rect 338 511 339 515
rect 343 511 344 515
rect 358 513 359 517
rect 363 513 364 517
rect 358 512 364 513
rect 422 517 428 518
rect 422 513 423 517
rect 427 513 428 517
rect 422 512 428 513
rect 478 517 484 518
rect 478 513 479 517
rect 483 513 484 517
rect 478 512 484 513
rect 542 517 548 518
rect 542 513 543 517
rect 547 513 548 517
rect 542 512 548 513
rect 598 517 604 518
rect 598 513 599 517
rect 603 513 604 517
rect 598 512 604 513
rect 654 517 660 518
rect 654 513 655 517
rect 659 513 660 517
rect 654 512 660 513
rect 710 517 716 518
rect 710 513 711 517
rect 715 513 716 517
rect 710 512 716 513
rect 766 517 772 518
rect 766 513 767 517
rect 771 513 772 517
rect 766 512 772 513
rect 830 517 836 518
rect 830 513 831 517
rect 835 513 836 517
rect 830 512 836 513
rect 894 517 900 518
rect 894 513 895 517
rect 899 513 900 517
rect 894 512 900 513
rect 912 512 914 538
rect 967 536 971 538
rect 1031 542 1035 543
rect 1031 536 1035 538
rect 1039 542 1043 544
rect 1039 537 1043 538
rect 1095 542 1099 543
rect 1095 536 1099 538
rect 1103 542 1107 544
rect 1103 537 1107 538
rect 1167 542 1171 544
rect 1167 536 1171 538
rect 1231 542 1235 544
rect 1231 537 1235 538
rect 1239 542 1243 543
rect 1239 536 1243 538
rect 1287 542 1291 544
rect 1287 537 1291 538
rect 1311 542 1315 543
rect 1311 536 1315 538
rect 1335 542 1339 544
rect 1335 537 1339 538
rect 1383 542 1387 544
rect 1383 537 1387 538
rect 1391 542 1395 543
rect 1391 536 1395 538
rect 1423 542 1427 544
rect 1423 537 1427 538
rect 1471 542 1475 544
rect 1471 537 1475 538
rect 1479 542 1483 543
rect 1479 536 1483 538
rect 1511 542 1515 544
rect 1511 537 1515 538
rect 1543 542 1547 544
rect 1543 536 1547 538
rect 966 535 972 536
rect 966 531 967 535
rect 971 531 972 535
rect 966 530 972 531
rect 1030 535 1036 536
rect 1030 531 1031 535
rect 1035 531 1036 535
rect 1030 530 1036 531
rect 1094 535 1100 536
rect 1094 531 1095 535
rect 1099 531 1100 535
rect 1094 530 1100 531
rect 1166 535 1172 536
rect 1166 531 1167 535
rect 1171 531 1172 535
rect 1166 530 1172 531
rect 1238 535 1244 536
rect 1238 531 1239 535
rect 1243 531 1244 535
rect 1238 530 1244 531
rect 1310 535 1316 536
rect 1310 531 1311 535
rect 1315 531 1316 535
rect 1310 530 1316 531
rect 1390 535 1396 536
rect 1390 531 1391 535
rect 1395 531 1396 535
rect 1390 530 1396 531
rect 1478 535 1484 536
rect 1478 531 1479 535
rect 1483 531 1484 535
rect 1478 530 1484 531
rect 1542 535 1548 536
rect 1542 531 1543 535
rect 1547 531 1548 535
rect 1542 530 1548 531
rect 966 517 972 518
rect 966 513 967 517
rect 971 513 972 517
rect 966 512 972 513
rect 1030 517 1036 518
rect 1030 513 1031 517
rect 1035 513 1036 517
rect 1030 512 1036 513
rect 1094 517 1100 518
rect 1094 513 1095 517
rect 1099 513 1100 517
rect 1094 512 1100 513
rect 1166 517 1172 518
rect 1166 513 1167 517
rect 1171 513 1172 517
rect 1166 512 1172 513
rect 1238 517 1244 518
rect 1238 513 1239 517
rect 1243 513 1244 517
rect 1238 512 1244 513
rect 1310 517 1316 518
rect 1310 513 1311 517
rect 1315 513 1316 517
rect 1310 512 1316 513
rect 1390 517 1396 518
rect 1390 513 1391 517
rect 1395 513 1396 517
rect 1390 512 1396 513
rect 1478 517 1484 518
rect 1478 513 1479 517
rect 1483 513 1484 517
rect 1478 512 1484 513
rect 1542 517 1548 518
rect 1542 513 1543 517
rect 1547 513 1548 517
rect 1542 512 1548 513
rect 338 510 344 511
rect 360 507 362 512
rect 366 511 372 512
rect 366 507 367 511
rect 371 507 372 511
rect 424 507 426 512
rect 480 507 482 512
rect 544 507 546 512
rect 600 507 602 512
rect 656 507 658 512
rect 694 507 700 508
rect 712 507 714 512
rect 768 507 770 512
rect 832 507 834 512
rect 896 507 898 512
rect 910 511 916 512
rect 910 507 911 511
rect 915 507 916 511
rect 968 507 970 512
rect 1032 507 1034 512
rect 1096 507 1098 512
rect 1168 507 1170 512
rect 1240 507 1242 512
rect 1312 507 1314 512
rect 1392 507 1394 512
rect 1480 507 1482 512
rect 1544 507 1546 512
rect 167 506 171 507
rect 167 501 171 502
rect 175 506 179 507
rect 175 501 179 502
rect 199 506 203 507
rect 199 501 203 502
rect 231 506 235 507
rect 231 501 235 502
rect 247 506 251 507
rect 247 501 251 502
rect 295 506 299 507
rect 295 501 299 502
rect 343 506 347 507
rect 343 501 347 502
rect 359 506 363 507
rect 366 506 372 507
rect 399 506 403 507
rect 359 501 363 502
rect 150 499 156 500
rect 110 492 111 496
rect 115 492 116 496
rect 110 491 116 492
rect 134 495 140 496
rect 134 491 135 495
rect 139 491 140 495
rect 150 495 151 499
rect 155 495 156 499
rect 168 496 170 501
rect 200 496 202 501
rect 248 496 250 501
rect 296 496 298 501
rect 326 499 332 500
rect 150 494 156 495
rect 166 495 172 496
rect 134 490 140 491
rect 166 491 167 495
rect 171 491 172 495
rect 166 490 172 491
rect 198 495 204 496
rect 198 491 199 495
rect 203 491 204 495
rect 198 490 204 491
rect 246 495 252 496
rect 246 491 247 495
rect 251 491 252 495
rect 246 490 252 491
rect 294 495 300 496
rect 294 491 295 495
rect 299 491 300 495
rect 326 495 327 499
rect 331 495 332 499
rect 344 496 346 501
rect 326 494 332 495
rect 342 495 348 496
rect 294 490 300 491
rect 266 483 272 484
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 266 479 267 483
rect 271 479 272 483
rect 266 478 272 479
rect 110 474 116 475
rect 134 477 140 478
rect 112 471 114 474
rect 134 473 135 477
rect 139 473 140 477
rect 134 472 140 473
rect 166 477 172 478
rect 166 473 167 477
rect 171 473 172 477
rect 166 472 172 473
rect 198 477 204 478
rect 198 473 199 477
rect 203 473 204 477
rect 198 472 204 473
rect 246 477 252 478
rect 246 473 247 477
rect 251 473 252 477
rect 246 472 252 473
rect 111 470 115 471
rect 111 465 115 466
rect 135 470 139 472
rect 112 462 114 465
rect 135 464 139 466
rect 167 470 171 472
rect 167 464 171 466
rect 199 470 203 472
rect 199 464 203 466
rect 247 470 251 472
rect 247 465 251 466
rect 255 470 259 471
rect 255 464 259 466
rect 134 463 140 464
rect 110 461 116 462
rect 110 457 111 461
rect 115 457 116 461
rect 134 459 135 463
rect 139 459 140 463
rect 134 458 140 459
rect 166 463 172 464
rect 166 459 167 463
rect 171 459 172 463
rect 166 458 172 459
rect 198 463 204 464
rect 198 459 199 463
rect 203 459 204 463
rect 198 458 204 459
rect 254 463 260 464
rect 254 459 255 463
rect 259 459 260 463
rect 254 458 260 459
rect 110 456 116 457
rect 150 455 156 456
rect 150 451 151 455
rect 155 451 156 455
rect 150 450 156 451
rect 134 445 140 446
rect 110 444 116 445
rect 110 440 111 444
rect 115 440 116 444
rect 134 441 135 445
rect 139 441 140 445
rect 134 440 140 441
rect 110 439 116 440
rect 112 431 114 439
rect 136 431 138 440
rect 111 430 115 431
rect 111 425 115 426
rect 135 430 139 431
rect 135 425 139 426
rect 112 421 114 425
rect 110 420 116 421
rect 136 420 138 425
rect 152 424 154 450
rect 166 445 172 446
rect 166 441 167 445
rect 171 441 172 445
rect 166 440 172 441
rect 198 445 204 446
rect 198 441 199 445
rect 203 441 204 445
rect 198 440 204 441
rect 254 445 260 446
rect 254 441 255 445
rect 259 441 260 445
rect 254 440 260 441
rect 268 440 270 478
rect 294 477 300 478
rect 294 473 295 477
rect 299 473 300 477
rect 294 472 300 473
rect 295 470 299 472
rect 295 465 299 466
rect 311 470 315 471
rect 311 464 315 466
rect 310 463 316 464
rect 310 459 311 463
rect 315 459 316 463
rect 310 458 316 459
rect 328 456 330 494
rect 342 491 343 495
rect 347 491 348 495
rect 342 490 348 491
rect 359 483 365 484
rect 359 479 360 483
rect 364 482 365 483
rect 368 482 370 506
rect 399 501 403 502
rect 423 506 427 507
rect 423 501 427 502
rect 455 506 459 507
rect 455 501 459 502
rect 479 506 483 507
rect 479 501 483 502
rect 511 506 515 507
rect 511 501 515 502
rect 543 506 547 507
rect 543 501 547 502
rect 567 506 571 507
rect 567 501 571 502
rect 599 506 603 507
rect 599 501 603 502
rect 623 506 627 507
rect 623 501 627 502
rect 655 506 659 507
rect 655 501 659 502
rect 679 506 683 507
rect 694 503 695 507
rect 699 503 700 507
rect 694 502 700 503
rect 711 506 715 507
rect 679 501 683 502
rect 400 496 402 501
rect 438 499 444 500
rect 398 495 404 496
rect 398 491 399 495
rect 403 491 404 495
rect 438 495 439 499
rect 443 495 444 499
rect 456 496 458 501
rect 512 496 514 501
rect 568 496 570 501
rect 624 496 626 501
rect 680 496 682 501
rect 438 494 444 495
rect 454 495 460 496
rect 398 490 404 491
rect 364 480 370 482
rect 364 479 365 480
rect 359 478 365 479
rect 342 477 348 478
rect 342 473 343 477
rect 347 473 348 477
rect 342 472 348 473
rect 398 477 404 478
rect 398 473 399 477
rect 403 473 404 477
rect 398 472 404 473
rect 343 470 347 472
rect 343 465 347 466
rect 367 470 371 471
rect 367 464 371 466
rect 399 470 403 472
rect 399 465 403 466
rect 423 470 427 471
rect 423 464 427 466
rect 366 463 372 464
rect 366 459 367 463
rect 371 459 372 463
rect 366 458 372 459
rect 422 463 428 464
rect 422 459 423 463
rect 427 459 428 463
rect 422 458 428 459
rect 440 456 442 494
rect 454 491 455 495
rect 459 491 460 495
rect 454 490 460 491
rect 510 495 516 496
rect 510 491 511 495
rect 515 491 516 495
rect 510 490 516 491
rect 566 495 572 496
rect 566 491 567 495
rect 571 491 572 495
rect 566 490 572 491
rect 622 495 628 496
rect 622 491 623 495
rect 627 491 628 495
rect 622 490 628 491
rect 678 495 684 496
rect 678 491 679 495
rect 683 491 684 495
rect 678 490 684 491
rect 696 484 698 502
rect 711 501 715 502
rect 743 506 747 507
rect 743 501 747 502
rect 767 506 771 507
rect 767 501 771 502
rect 815 506 819 507
rect 815 501 819 502
rect 831 506 835 507
rect 831 501 835 502
rect 887 506 891 507
rect 887 501 891 502
rect 895 506 899 507
rect 910 506 916 507
rect 959 506 963 507
rect 895 501 899 502
rect 959 501 963 502
rect 967 506 971 507
rect 967 501 971 502
rect 1031 506 1035 507
rect 1031 501 1035 502
rect 1039 506 1043 507
rect 1039 501 1043 502
rect 1095 506 1099 507
rect 1095 501 1099 502
rect 1127 506 1131 507
rect 1127 501 1131 502
rect 1167 506 1171 507
rect 1167 501 1171 502
rect 1223 506 1227 507
rect 1223 501 1227 502
rect 1239 506 1243 507
rect 1239 501 1243 502
rect 1311 506 1315 507
rect 1311 501 1315 502
rect 1327 506 1331 507
rect 1327 501 1331 502
rect 1391 506 1395 507
rect 1391 501 1395 502
rect 1439 506 1443 507
rect 1439 501 1443 502
rect 1479 506 1483 507
rect 1543 506 1547 507
rect 1479 501 1483 502
rect 1498 503 1504 504
rect 744 496 746 501
rect 816 496 818 501
rect 888 496 890 501
rect 960 496 962 501
rect 1040 496 1042 501
rect 1128 496 1130 501
rect 1214 499 1220 500
rect 742 495 748 496
rect 742 491 743 495
rect 747 491 748 495
rect 742 490 748 491
rect 814 495 820 496
rect 814 491 815 495
rect 819 491 820 495
rect 814 490 820 491
rect 886 495 892 496
rect 886 491 887 495
rect 891 491 892 495
rect 886 490 892 491
rect 958 495 964 496
rect 958 491 959 495
rect 963 491 964 495
rect 958 490 964 491
rect 1038 495 1044 496
rect 1038 491 1039 495
rect 1043 491 1044 495
rect 1038 490 1044 491
rect 1126 495 1132 496
rect 1126 491 1127 495
rect 1131 491 1132 495
rect 1214 495 1215 499
rect 1219 495 1220 499
rect 1224 496 1226 501
rect 1328 496 1330 501
rect 1440 496 1442 501
rect 1498 499 1499 503
rect 1503 499 1504 503
rect 1543 501 1547 502
rect 1498 498 1504 499
rect 1214 494 1220 495
rect 1222 495 1228 496
rect 1126 490 1132 491
rect 694 483 700 484
rect 694 479 695 483
rect 699 479 700 483
rect 694 478 700 479
rect 454 477 460 478
rect 454 473 455 477
rect 459 473 460 477
rect 454 472 460 473
rect 510 477 516 478
rect 510 473 511 477
rect 515 473 516 477
rect 510 472 516 473
rect 566 477 572 478
rect 566 473 567 477
rect 571 473 572 477
rect 566 472 572 473
rect 622 477 628 478
rect 622 473 623 477
rect 627 473 628 477
rect 622 472 628 473
rect 678 477 684 478
rect 678 473 679 477
rect 683 473 684 477
rect 678 472 684 473
rect 742 477 748 478
rect 742 473 743 477
rect 747 473 748 477
rect 742 472 748 473
rect 814 477 820 478
rect 814 473 815 477
rect 819 473 820 477
rect 814 472 820 473
rect 886 477 892 478
rect 886 473 887 477
rect 891 473 892 477
rect 886 472 892 473
rect 958 477 964 478
rect 958 473 959 477
rect 963 473 964 477
rect 958 472 964 473
rect 1038 477 1044 478
rect 1038 473 1039 477
rect 1043 473 1044 477
rect 1038 472 1044 473
rect 1126 477 1132 478
rect 1126 473 1127 477
rect 1131 473 1132 477
rect 1126 472 1132 473
rect 1216 472 1218 494
rect 1222 491 1223 495
rect 1227 491 1228 495
rect 1222 490 1228 491
rect 1326 495 1332 496
rect 1326 491 1327 495
rect 1331 491 1332 495
rect 1326 490 1332 491
rect 1438 495 1444 496
rect 1438 491 1439 495
rect 1443 491 1444 495
rect 1438 490 1444 491
rect 1278 483 1284 484
rect 1278 479 1279 483
rect 1283 479 1284 483
rect 1278 478 1284 479
rect 1222 477 1228 478
rect 1222 473 1223 477
rect 1227 473 1228 477
rect 1222 472 1228 473
rect 455 470 459 472
rect 455 465 459 466
rect 479 470 483 471
rect 479 464 483 466
rect 511 470 515 472
rect 554 471 560 472
rect 511 465 515 466
rect 535 470 539 471
rect 554 467 555 471
rect 559 467 560 471
rect 554 466 560 467
rect 567 470 571 472
rect 535 464 539 466
rect 478 463 484 464
rect 478 459 479 463
rect 483 459 484 463
rect 478 458 484 459
rect 534 463 540 464
rect 534 459 535 463
rect 539 459 540 463
rect 534 458 540 459
rect 326 455 332 456
rect 326 451 327 455
rect 331 451 332 455
rect 326 450 332 451
rect 438 455 444 456
rect 438 451 439 455
rect 443 451 444 455
rect 438 450 444 451
rect 310 445 316 446
rect 310 441 311 445
rect 315 441 316 445
rect 310 440 316 441
rect 366 445 372 446
rect 366 441 367 445
rect 371 441 372 445
rect 366 440 372 441
rect 422 445 428 446
rect 422 441 423 445
rect 427 441 428 445
rect 422 440 428 441
rect 478 445 484 446
rect 478 441 479 445
rect 483 441 484 445
rect 478 440 484 441
rect 534 445 540 446
rect 534 441 535 445
rect 539 441 540 445
rect 534 440 540 441
rect 556 440 558 466
rect 567 465 571 466
rect 599 470 603 471
rect 599 464 603 466
rect 623 470 627 472
rect 623 465 627 466
rect 663 470 667 471
rect 663 464 667 466
rect 679 470 683 472
rect 679 465 683 466
rect 735 470 739 471
rect 735 464 739 466
rect 743 470 747 472
rect 743 465 747 466
rect 807 470 811 471
rect 807 464 811 466
rect 815 470 819 472
rect 815 465 819 466
rect 871 470 875 471
rect 871 464 875 466
rect 887 470 891 472
rect 894 471 900 472
rect 894 467 895 471
rect 899 467 900 471
rect 894 466 900 467
rect 935 470 939 471
rect 887 465 891 466
rect 598 463 604 464
rect 598 459 599 463
rect 603 459 604 463
rect 598 458 604 459
rect 662 463 668 464
rect 662 459 663 463
rect 667 459 668 463
rect 662 458 668 459
rect 734 463 740 464
rect 734 459 735 463
rect 739 459 740 463
rect 734 458 740 459
rect 806 463 812 464
rect 806 459 807 463
rect 811 459 812 463
rect 806 458 812 459
rect 870 463 876 464
rect 870 459 871 463
rect 875 459 876 463
rect 870 458 876 459
rect 778 455 784 456
rect 778 451 779 455
rect 783 451 784 455
rect 778 450 784 451
rect 598 445 604 446
rect 598 441 599 445
rect 603 441 604 445
rect 598 440 604 441
rect 662 445 668 446
rect 662 441 663 445
rect 667 441 668 445
rect 662 440 668 441
rect 734 445 740 446
rect 734 441 735 445
rect 739 441 740 445
rect 734 440 740 441
rect 168 431 170 440
rect 200 431 202 440
rect 256 431 258 440
rect 266 439 272 440
rect 266 435 267 439
rect 271 435 272 439
rect 266 434 272 435
rect 312 431 314 440
rect 368 431 370 440
rect 378 439 384 440
rect 378 435 379 439
rect 383 435 384 439
rect 378 434 384 435
rect 167 430 171 431
rect 167 425 171 426
rect 199 430 203 431
rect 199 425 203 426
rect 231 430 235 431
rect 231 425 235 426
rect 255 430 259 431
rect 255 425 259 426
rect 295 430 299 431
rect 295 425 299 426
rect 311 430 315 431
rect 311 425 315 426
rect 359 430 363 431
rect 359 425 363 426
rect 367 430 371 431
rect 367 425 371 426
rect 150 423 156 424
rect 110 416 111 420
rect 115 416 116 420
rect 110 415 116 416
rect 134 419 140 420
rect 134 415 135 419
rect 139 415 140 419
rect 150 419 151 423
rect 155 419 156 423
rect 168 420 170 425
rect 232 420 234 425
rect 296 420 298 425
rect 360 420 362 425
rect 150 418 156 419
rect 166 419 172 420
rect 134 414 140 415
rect 166 415 167 419
rect 171 415 172 419
rect 166 414 172 415
rect 230 419 236 420
rect 230 415 231 419
rect 235 415 236 419
rect 230 414 236 415
rect 294 419 300 420
rect 294 415 295 419
rect 299 415 300 419
rect 294 414 300 415
rect 358 419 364 420
rect 358 415 359 419
rect 363 415 364 419
rect 358 414 364 415
rect 380 408 382 434
rect 424 431 426 440
rect 480 431 482 440
rect 536 431 538 440
rect 554 439 560 440
rect 554 435 555 439
rect 559 435 560 439
rect 554 434 560 435
rect 562 439 568 440
rect 562 435 563 439
rect 567 435 568 439
rect 562 434 568 435
rect 423 430 427 431
rect 423 425 427 426
rect 479 430 483 431
rect 479 425 483 426
rect 487 430 491 431
rect 487 425 491 426
rect 535 430 539 431
rect 535 425 539 426
rect 543 430 547 431
rect 543 425 547 426
rect 424 420 426 425
rect 488 420 490 425
rect 544 420 546 425
rect 422 419 428 420
rect 422 415 423 419
rect 427 415 428 419
rect 422 414 428 415
rect 486 419 492 420
rect 486 415 487 419
rect 491 415 492 419
rect 486 414 492 415
rect 542 419 548 420
rect 542 415 543 419
rect 547 415 548 419
rect 542 414 548 415
rect 564 408 566 434
rect 600 431 602 440
rect 606 431 612 432
rect 664 431 666 440
rect 736 431 738 440
rect 591 430 595 431
rect 591 425 595 426
rect 599 430 603 431
rect 606 427 607 431
rect 611 427 612 431
rect 606 426 612 427
rect 639 430 643 431
rect 599 425 603 426
rect 592 420 594 425
rect 590 419 596 420
rect 590 415 591 419
rect 595 415 596 419
rect 590 414 596 415
rect 608 408 610 426
rect 639 425 643 426
rect 663 430 667 431
rect 663 425 667 426
rect 679 430 683 431
rect 679 425 683 426
rect 719 430 723 431
rect 719 425 723 426
rect 735 430 739 431
rect 735 425 739 426
rect 759 430 763 431
rect 759 425 763 426
rect 640 420 642 425
rect 680 420 682 425
rect 720 420 722 425
rect 760 420 762 425
rect 780 424 782 450
rect 806 445 812 446
rect 806 441 807 445
rect 811 441 812 445
rect 806 440 812 441
rect 870 445 876 446
rect 870 441 871 445
rect 875 441 876 445
rect 870 440 876 441
rect 808 431 810 440
rect 872 431 874 440
rect 887 439 893 440
rect 887 435 888 439
rect 892 438 893 439
rect 896 438 898 466
rect 935 464 939 466
rect 959 470 963 472
rect 959 465 963 466
rect 991 470 995 471
rect 991 464 995 466
rect 1039 470 1043 472
rect 1039 465 1043 466
rect 1047 470 1051 471
rect 1047 464 1051 466
rect 1095 470 1099 471
rect 1095 464 1099 466
rect 1127 470 1131 472
rect 1214 471 1220 472
rect 1127 465 1131 466
rect 1143 470 1147 471
rect 1143 464 1147 466
rect 1199 470 1203 471
rect 1214 467 1215 471
rect 1219 467 1220 471
rect 1214 466 1220 467
rect 1223 470 1227 472
rect 1199 464 1203 466
rect 1223 465 1227 466
rect 1263 470 1267 471
rect 1263 464 1267 466
rect 934 463 940 464
rect 934 459 935 463
rect 939 459 940 463
rect 934 458 940 459
rect 990 463 996 464
rect 990 459 991 463
rect 995 459 996 463
rect 990 458 996 459
rect 1046 463 1052 464
rect 1046 459 1047 463
rect 1051 459 1052 463
rect 1046 458 1052 459
rect 1094 463 1100 464
rect 1094 459 1095 463
rect 1099 459 1100 463
rect 1094 458 1100 459
rect 1142 463 1148 464
rect 1142 459 1143 463
rect 1147 459 1148 463
rect 1142 458 1148 459
rect 1198 463 1204 464
rect 1198 459 1199 463
rect 1203 459 1204 463
rect 1198 458 1204 459
rect 1262 463 1268 464
rect 1262 459 1263 463
rect 1267 459 1268 463
rect 1262 458 1268 459
rect 1038 455 1044 456
rect 1038 451 1039 455
rect 1043 451 1044 455
rect 1038 450 1044 451
rect 934 445 940 446
rect 934 441 935 445
rect 939 441 940 445
rect 934 440 940 441
rect 990 445 996 446
rect 990 441 991 445
rect 995 441 996 445
rect 990 440 996 441
rect 892 436 898 438
rect 892 435 893 436
rect 887 434 893 435
rect 936 431 938 440
rect 992 431 994 440
rect 807 430 811 431
rect 807 425 811 426
rect 863 430 867 431
rect 863 425 867 426
rect 871 430 875 431
rect 871 425 875 426
rect 919 430 923 431
rect 919 425 923 426
rect 935 430 939 431
rect 935 425 939 426
rect 975 430 979 431
rect 975 425 979 426
rect 991 430 995 431
rect 991 425 995 426
rect 1031 430 1035 431
rect 1040 428 1042 450
rect 1046 445 1052 446
rect 1046 441 1047 445
rect 1051 441 1052 445
rect 1046 440 1052 441
rect 1094 445 1100 446
rect 1094 441 1095 445
rect 1099 441 1100 445
rect 1094 440 1100 441
rect 1142 445 1148 446
rect 1142 441 1143 445
rect 1147 441 1148 445
rect 1142 440 1148 441
rect 1198 445 1204 446
rect 1198 441 1199 445
rect 1203 441 1204 445
rect 1198 440 1204 441
rect 1262 445 1268 446
rect 1262 441 1263 445
rect 1267 441 1268 445
rect 1262 440 1268 441
rect 1280 440 1282 478
rect 1326 477 1332 478
rect 1326 473 1327 477
rect 1331 473 1332 477
rect 1326 472 1332 473
rect 1438 477 1444 478
rect 1438 473 1439 477
rect 1443 473 1444 477
rect 1438 472 1444 473
rect 1327 470 1331 472
rect 1327 464 1331 466
rect 1399 470 1403 471
rect 1399 464 1403 466
rect 1439 470 1443 472
rect 1439 465 1443 466
rect 1479 470 1483 471
rect 1479 464 1483 466
rect 1326 463 1332 464
rect 1326 459 1327 463
rect 1331 459 1332 463
rect 1326 458 1332 459
rect 1398 463 1404 464
rect 1398 459 1399 463
rect 1403 459 1404 463
rect 1398 458 1404 459
rect 1478 463 1484 464
rect 1478 459 1479 463
rect 1483 459 1484 463
rect 1478 458 1484 459
rect 1500 456 1502 498
rect 1544 496 1546 501
rect 1542 495 1548 496
rect 1542 491 1543 495
rect 1547 491 1548 495
rect 1542 490 1548 491
rect 1552 484 1554 570
rect 1584 569 1586 573
rect 1582 568 1588 569
rect 1582 564 1583 568
rect 1587 564 1588 568
rect 1582 563 1588 564
rect 1558 555 1564 556
rect 1558 551 1559 555
rect 1563 551 1564 555
rect 1558 550 1564 551
rect 1582 551 1588 552
rect 1560 512 1562 550
rect 1582 547 1583 551
rect 1587 547 1588 551
rect 1582 546 1588 547
rect 1584 543 1586 546
rect 1583 542 1587 543
rect 1583 537 1587 538
rect 1584 534 1586 537
rect 1582 533 1588 534
rect 1582 529 1583 533
rect 1587 529 1588 533
rect 1582 528 1588 529
rect 1582 516 1588 517
rect 1582 512 1583 516
rect 1587 512 1588 516
rect 1558 511 1564 512
rect 1582 511 1588 512
rect 1558 507 1559 511
rect 1563 507 1564 511
rect 1584 507 1586 511
rect 1558 506 1564 507
rect 1583 506 1587 507
rect 1583 501 1587 502
rect 1584 497 1586 501
rect 1582 496 1588 497
rect 1582 492 1583 496
rect 1587 492 1588 496
rect 1582 491 1588 492
rect 1552 483 1560 484
rect 1552 481 1555 483
rect 1554 479 1555 481
rect 1559 479 1560 483
rect 1554 478 1560 479
rect 1582 479 1588 480
rect 1542 477 1548 478
rect 1542 473 1543 477
rect 1547 473 1548 477
rect 1582 475 1583 479
rect 1587 475 1588 479
rect 1582 474 1588 475
rect 1542 472 1548 473
rect 1543 470 1547 472
rect 1584 471 1586 474
rect 1543 464 1547 466
rect 1583 470 1587 471
rect 1583 465 1587 466
rect 1542 463 1548 464
rect 1542 459 1543 463
rect 1547 459 1548 463
rect 1584 462 1586 465
rect 1542 458 1548 459
rect 1582 461 1588 462
rect 1582 457 1583 461
rect 1587 457 1588 461
rect 1582 456 1588 457
rect 1390 455 1396 456
rect 1390 451 1391 455
rect 1395 451 1396 455
rect 1390 450 1396 451
rect 1498 455 1504 456
rect 1498 451 1499 455
rect 1503 451 1504 455
rect 1498 450 1504 451
rect 1558 455 1564 456
rect 1558 451 1559 455
rect 1563 451 1564 455
rect 1558 450 1564 451
rect 1326 445 1332 446
rect 1326 441 1327 445
rect 1331 441 1332 445
rect 1326 440 1332 441
rect 1048 431 1050 440
rect 1096 431 1098 440
rect 1144 431 1146 440
rect 1200 431 1202 440
rect 1264 431 1266 440
rect 1278 439 1284 440
rect 1278 435 1279 439
rect 1283 435 1284 439
rect 1278 434 1284 435
rect 1328 431 1330 440
rect 1392 432 1394 450
rect 1398 445 1404 446
rect 1398 441 1399 445
rect 1403 441 1404 445
rect 1398 440 1404 441
rect 1478 445 1484 446
rect 1478 441 1479 445
rect 1483 441 1484 445
rect 1478 440 1484 441
rect 1542 445 1548 446
rect 1542 441 1543 445
rect 1547 441 1548 445
rect 1542 440 1548 441
rect 1390 431 1396 432
rect 1400 431 1402 440
rect 1480 431 1482 440
rect 1486 439 1492 440
rect 1486 435 1487 439
rect 1491 435 1492 439
rect 1486 434 1492 435
rect 1047 430 1051 431
rect 1031 425 1035 426
rect 1038 427 1044 428
rect 778 423 784 424
rect 638 419 644 420
rect 638 415 639 419
rect 643 415 644 419
rect 638 414 644 415
rect 678 419 684 420
rect 678 415 679 419
rect 683 415 684 419
rect 678 414 684 415
rect 718 419 724 420
rect 718 415 719 419
rect 723 415 724 419
rect 718 414 724 415
rect 758 419 764 420
rect 758 415 759 419
rect 763 415 764 419
rect 778 419 779 423
rect 783 419 784 423
rect 808 420 810 425
rect 864 420 866 425
rect 920 420 922 425
rect 976 420 978 425
rect 1032 420 1034 425
rect 1038 423 1039 427
rect 1043 423 1044 427
rect 1047 425 1051 426
rect 1087 430 1091 431
rect 1087 425 1091 426
rect 1095 430 1099 431
rect 1095 425 1099 426
rect 1143 430 1147 431
rect 1143 425 1147 426
rect 1151 430 1155 431
rect 1151 425 1155 426
rect 1199 430 1203 431
rect 1199 425 1203 426
rect 1223 430 1227 431
rect 1223 425 1227 426
rect 1263 430 1267 431
rect 1263 425 1267 426
rect 1303 430 1307 431
rect 1303 425 1307 426
rect 1327 430 1331 431
rect 1327 425 1331 426
rect 1383 430 1387 431
rect 1390 427 1391 431
rect 1395 427 1396 431
rect 1390 426 1396 427
rect 1399 430 1403 431
rect 1383 425 1387 426
rect 1399 425 1403 426
rect 1471 430 1475 431
rect 1471 425 1475 426
rect 1479 430 1483 431
rect 1479 425 1483 426
rect 1038 422 1044 423
rect 1088 420 1090 425
rect 1152 420 1154 425
rect 1224 420 1226 425
rect 1304 420 1306 425
rect 1384 420 1386 425
rect 1472 420 1474 425
rect 778 418 784 419
rect 806 419 812 420
rect 758 414 764 415
rect 806 415 807 419
rect 811 415 812 419
rect 806 414 812 415
rect 862 419 868 420
rect 862 415 863 419
rect 867 415 868 419
rect 862 414 868 415
rect 918 419 924 420
rect 918 415 919 419
rect 923 415 924 419
rect 918 414 924 415
rect 974 419 980 420
rect 974 415 975 419
rect 979 415 980 419
rect 974 414 980 415
rect 1030 419 1036 420
rect 1030 415 1031 419
rect 1035 415 1036 419
rect 1030 414 1036 415
rect 1086 419 1092 420
rect 1086 415 1087 419
rect 1091 415 1092 419
rect 1086 414 1092 415
rect 1150 419 1156 420
rect 1150 415 1151 419
rect 1155 415 1156 419
rect 1150 414 1156 415
rect 1222 419 1228 420
rect 1222 415 1223 419
rect 1227 415 1228 419
rect 1222 414 1228 415
rect 1302 419 1308 420
rect 1302 415 1303 419
rect 1307 415 1308 419
rect 1302 414 1308 415
rect 1382 419 1388 420
rect 1382 415 1383 419
rect 1387 415 1388 419
rect 1382 414 1388 415
rect 1470 419 1476 420
rect 1470 415 1471 419
rect 1475 415 1476 419
rect 1470 414 1476 415
rect 1488 408 1490 434
rect 1544 431 1546 440
rect 1543 430 1547 431
rect 1543 425 1547 426
rect 1502 423 1508 424
rect 1502 419 1503 423
rect 1507 419 1508 423
rect 1544 420 1546 425
rect 1560 424 1562 450
rect 1582 444 1588 445
rect 1582 440 1583 444
rect 1587 440 1588 444
rect 1582 439 1588 440
rect 1584 431 1586 439
rect 1583 430 1587 431
rect 1583 425 1587 426
rect 1558 423 1564 424
rect 1502 418 1508 419
rect 1542 419 1548 420
rect 310 407 316 408
rect 110 403 116 404
rect 110 399 111 403
rect 115 399 116 403
rect 310 403 311 407
rect 315 403 316 407
rect 310 402 316 403
rect 378 407 384 408
rect 378 403 379 407
rect 383 403 384 407
rect 378 402 384 403
rect 562 407 568 408
rect 562 403 563 407
rect 567 403 568 407
rect 562 402 568 403
rect 606 407 612 408
rect 606 403 607 407
rect 611 403 612 407
rect 606 402 612 403
rect 1486 407 1492 408
rect 1486 403 1487 407
rect 1491 403 1492 407
rect 1486 402 1492 403
rect 110 398 116 399
rect 134 401 140 402
rect 112 395 114 398
rect 134 397 135 401
rect 139 397 140 401
rect 134 396 140 397
rect 166 401 172 402
rect 166 397 167 401
rect 171 397 172 401
rect 166 396 172 397
rect 230 401 236 402
rect 230 397 231 401
rect 235 397 236 401
rect 230 396 236 397
rect 294 401 300 402
rect 294 397 295 401
rect 299 397 300 401
rect 294 396 300 397
rect 111 394 115 395
rect 111 389 115 390
rect 135 394 139 396
rect 112 386 114 389
rect 135 388 139 390
rect 167 394 171 396
rect 167 389 171 390
rect 207 394 211 395
rect 207 388 211 390
rect 231 394 235 396
rect 231 389 235 390
rect 295 394 299 396
rect 295 388 299 390
rect 134 387 140 388
rect 110 385 116 386
rect 110 381 111 385
rect 115 381 116 385
rect 134 383 135 387
rect 139 383 140 387
rect 134 382 140 383
rect 206 387 212 388
rect 206 383 207 387
rect 211 383 212 387
rect 206 382 212 383
rect 294 387 300 388
rect 294 383 295 387
rect 299 383 300 387
rect 294 382 300 383
rect 110 380 116 381
rect 150 379 156 380
rect 150 375 151 379
rect 155 375 156 379
rect 150 374 156 375
rect 134 369 140 370
rect 110 368 116 369
rect 110 364 111 368
rect 115 364 116 368
rect 134 365 135 369
rect 139 365 140 369
rect 134 364 140 365
rect 110 363 116 364
rect 112 359 114 363
rect 136 359 138 364
rect 111 358 115 359
rect 111 353 115 354
rect 135 358 139 359
rect 135 353 139 354
rect 112 349 114 353
rect 110 348 116 349
rect 136 348 138 353
rect 152 352 154 374
rect 312 372 314 402
rect 358 401 364 402
rect 358 397 359 401
rect 363 397 364 401
rect 358 396 364 397
rect 422 401 428 402
rect 422 397 423 401
rect 427 397 428 401
rect 422 396 428 397
rect 486 401 492 402
rect 486 397 487 401
rect 491 397 492 401
rect 486 396 492 397
rect 542 401 548 402
rect 542 397 543 401
rect 547 397 548 401
rect 542 396 548 397
rect 590 401 596 402
rect 590 397 591 401
rect 595 397 596 401
rect 590 396 596 397
rect 638 401 644 402
rect 638 397 639 401
rect 643 397 644 401
rect 638 396 644 397
rect 678 401 684 402
rect 678 397 679 401
rect 683 397 684 401
rect 678 396 684 397
rect 718 401 724 402
rect 718 397 719 401
rect 723 397 724 401
rect 718 396 724 397
rect 758 401 764 402
rect 758 397 759 401
rect 763 397 764 401
rect 758 396 764 397
rect 806 401 812 402
rect 806 397 807 401
rect 811 397 812 401
rect 806 396 812 397
rect 862 401 868 402
rect 862 397 863 401
rect 867 397 868 401
rect 862 396 868 397
rect 918 401 924 402
rect 918 397 919 401
rect 923 397 924 401
rect 918 396 924 397
rect 974 401 980 402
rect 974 397 975 401
rect 979 397 980 401
rect 974 396 980 397
rect 1030 401 1036 402
rect 1030 397 1031 401
rect 1035 397 1036 401
rect 1030 396 1036 397
rect 1086 401 1092 402
rect 1086 397 1087 401
rect 1091 397 1092 401
rect 1086 396 1092 397
rect 1150 401 1156 402
rect 1150 397 1151 401
rect 1155 397 1156 401
rect 1150 396 1156 397
rect 1222 401 1228 402
rect 1222 397 1223 401
rect 1227 397 1228 401
rect 1222 396 1228 397
rect 1302 401 1308 402
rect 1302 397 1303 401
rect 1307 397 1308 401
rect 1302 396 1308 397
rect 1382 401 1388 402
rect 1382 397 1383 401
rect 1387 397 1388 401
rect 1382 396 1388 397
rect 1470 401 1476 402
rect 1470 397 1471 401
rect 1475 397 1476 401
rect 1470 396 1476 397
rect 359 394 363 396
rect 359 389 363 390
rect 383 394 387 395
rect 383 388 387 390
rect 423 394 427 396
rect 423 389 427 390
rect 463 394 467 395
rect 463 388 467 390
rect 487 394 491 396
rect 487 389 491 390
rect 535 394 539 395
rect 535 388 539 390
rect 543 394 547 396
rect 543 389 547 390
rect 591 394 595 396
rect 591 389 595 390
rect 599 394 603 395
rect 599 388 603 390
rect 639 394 643 396
rect 639 389 643 390
rect 655 394 659 395
rect 655 388 659 390
rect 679 394 683 396
rect 679 389 683 390
rect 703 394 707 395
rect 703 388 707 390
rect 719 394 723 396
rect 719 389 723 390
rect 751 394 755 395
rect 751 388 755 390
rect 759 394 763 396
rect 759 389 763 390
rect 807 394 811 396
rect 826 395 832 396
rect 826 391 827 395
rect 831 391 832 395
rect 826 390 832 391
rect 863 394 867 396
rect 807 388 811 390
rect 382 387 388 388
rect 382 383 383 387
rect 387 383 388 387
rect 382 382 388 383
rect 462 387 468 388
rect 462 383 463 387
rect 467 383 468 387
rect 462 382 468 383
rect 534 387 540 388
rect 534 383 535 387
rect 539 383 540 387
rect 534 382 540 383
rect 598 387 604 388
rect 598 383 599 387
rect 603 383 604 387
rect 598 382 604 383
rect 654 387 660 388
rect 654 383 655 387
rect 659 383 660 387
rect 654 382 660 383
rect 702 387 708 388
rect 702 383 703 387
rect 707 383 708 387
rect 702 382 708 383
rect 750 387 756 388
rect 750 383 751 387
rect 755 383 756 387
rect 750 382 756 383
rect 806 387 812 388
rect 806 383 807 387
rect 811 383 812 387
rect 806 382 812 383
rect 310 371 316 372
rect 206 369 212 370
rect 206 365 207 369
rect 211 365 212 369
rect 206 364 212 365
rect 294 369 300 370
rect 294 365 295 369
rect 299 365 300 369
rect 310 367 311 371
rect 315 367 316 371
rect 310 366 316 367
rect 382 369 388 370
rect 294 364 300 365
rect 382 365 383 369
rect 387 365 388 369
rect 382 364 388 365
rect 462 369 468 370
rect 462 365 463 369
rect 467 365 468 369
rect 462 364 468 365
rect 534 369 540 370
rect 534 365 535 369
rect 539 365 540 369
rect 534 364 540 365
rect 598 369 604 370
rect 598 365 599 369
rect 603 365 604 369
rect 598 364 604 365
rect 654 369 660 370
rect 654 365 655 369
rect 659 365 660 369
rect 654 364 660 365
rect 702 369 708 370
rect 702 365 703 369
rect 707 365 708 369
rect 702 364 708 365
rect 750 369 756 370
rect 750 365 751 369
rect 755 365 756 369
rect 750 364 756 365
rect 806 369 812 370
rect 806 365 807 369
rect 811 365 812 369
rect 806 364 812 365
rect 828 364 830 390
rect 863 388 867 390
rect 919 394 923 396
rect 919 388 923 390
rect 975 394 979 396
rect 975 389 979 390
rect 983 394 987 395
rect 983 388 987 390
rect 1031 394 1035 396
rect 1031 389 1035 390
rect 1055 394 1059 395
rect 1055 388 1059 390
rect 1087 394 1091 396
rect 1087 389 1091 390
rect 1127 394 1131 395
rect 1127 388 1131 390
rect 1151 394 1155 396
rect 1158 395 1164 396
rect 1158 391 1159 395
rect 1163 391 1164 395
rect 1158 390 1164 391
rect 1199 394 1203 395
rect 1151 389 1155 390
rect 862 387 868 388
rect 862 383 863 387
rect 867 383 868 387
rect 862 382 868 383
rect 918 387 924 388
rect 918 383 919 387
rect 923 383 924 387
rect 918 382 924 383
rect 982 387 988 388
rect 982 383 983 387
rect 987 383 988 387
rect 982 382 988 383
rect 1054 387 1060 388
rect 1054 383 1055 387
rect 1059 383 1060 387
rect 1054 382 1060 383
rect 1126 387 1132 388
rect 1126 383 1127 387
rect 1131 383 1132 387
rect 1126 382 1132 383
rect 1070 379 1076 380
rect 1070 375 1071 379
rect 1075 375 1076 379
rect 1070 374 1076 375
rect 862 369 868 370
rect 862 365 863 369
rect 867 365 868 369
rect 862 364 868 365
rect 918 369 924 370
rect 918 365 919 369
rect 923 365 924 369
rect 918 364 924 365
rect 982 369 988 370
rect 982 365 983 369
rect 987 365 988 369
rect 982 364 988 365
rect 1054 369 1060 370
rect 1054 365 1055 369
rect 1059 365 1060 369
rect 1054 364 1060 365
rect 208 359 210 364
rect 296 359 298 364
rect 350 363 356 364
rect 350 359 351 363
rect 355 359 356 363
rect 384 359 386 364
rect 464 359 466 364
rect 536 359 538 364
rect 574 363 580 364
rect 574 359 575 363
rect 579 359 580 363
rect 600 359 602 364
rect 656 359 658 364
rect 704 359 706 364
rect 752 359 754 364
rect 808 359 810 364
rect 826 363 832 364
rect 826 359 827 363
rect 831 359 832 363
rect 864 359 866 364
rect 920 359 922 364
rect 984 359 986 364
rect 1056 359 1058 364
rect 175 358 179 359
rect 175 353 179 354
rect 207 358 211 359
rect 207 353 211 354
rect 223 358 227 359
rect 223 353 227 354
rect 279 358 283 359
rect 279 353 283 354
rect 295 358 299 359
rect 295 353 299 354
rect 335 358 339 359
rect 350 358 356 359
rect 383 358 387 359
rect 335 353 339 354
rect 150 351 156 352
rect 110 344 111 348
rect 115 344 116 348
rect 110 343 116 344
rect 134 347 140 348
rect 134 343 135 347
rect 139 343 140 347
rect 150 347 151 351
rect 155 347 156 351
rect 176 348 178 353
rect 224 348 226 353
rect 280 348 282 353
rect 336 348 338 353
rect 150 346 156 347
rect 174 347 180 348
rect 134 342 140 343
rect 174 343 175 347
rect 179 343 180 347
rect 174 342 180 343
rect 222 347 228 348
rect 222 343 223 347
rect 227 343 228 347
rect 222 342 228 343
rect 278 347 284 348
rect 278 343 279 347
rect 283 343 284 347
rect 278 342 284 343
rect 334 347 340 348
rect 334 343 335 347
rect 339 343 340 347
rect 334 342 340 343
rect 352 336 354 358
rect 383 353 387 354
rect 391 358 395 359
rect 391 353 395 354
rect 447 358 451 359
rect 447 353 451 354
rect 463 358 467 359
rect 463 353 467 354
rect 503 358 507 359
rect 503 353 507 354
rect 535 358 539 359
rect 535 353 539 354
rect 567 358 571 359
rect 574 358 580 359
rect 599 358 603 359
rect 567 353 571 354
rect 392 348 394 353
rect 402 351 408 352
rect 390 347 396 348
rect 390 343 391 347
rect 395 343 396 347
rect 402 347 403 351
rect 407 347 408 351
rect 448 348 450 353
rect 494 351 500 352
rect 402 346 408 347
rect 446 347 452 348
rect 390 342 396 343
rect 310 335 316 336
rect 110 331 116 332
rect 110 327 111 331
rect 115 327 116 331
rect 310 331 311 335
rect 315 331 316 335
rect 310 330 316 331
rect 350 335 356 336
rect 350 331 351 335
rect 355 331 356 335
rect 404 331 406 346
rect 446 343 447 347
rect 451 343 452 347
rect 494 347 495 351
rect 499 347 500 351
rect 504 348 506 353
rect 568 348 570 353
rect 494 346 500 347
rect 502 347 508 348
rect 446 342 452 343
rect 350 330 356 331
rect 110 326 116 327
rect 134 329 140 330
rect 112 323 114 326
rect 134 325 135 329
rect 139 325 140 329
rect 134 324 140 325
rect 174 329 180 330
rect 174 325 175 329
rect 179 325 180 329
rect 174 324 180 325
rect 222 329 228 330
rect 222 325 223 329
rect 227 325 228 329
rect 222 324 228 325
rect 278 329 284 330
rect 278 325 279 329
rect 283 325 284 329
rect 278 324 284 325
rect 111 322 115 323
rect 111 317 115 318
rect 135 322 139 324
rect 135 317 139 318
rect 175 322 179 324
rect 175 317 179 318
rect 191 322 195 323
rect 112 314 114 317
rect 191 316 195 318
rect 223 322 227 324
rect 223 316 227 318
rect 255 322 259 323
rect 255 316 259 318
rect 279 322 283 324
rect 279 317 283 318
rect 295 322 299 323
rect 295 316 299 318
rect 190 315 196 316
rect 110 313 116 314
rect 110 309 111 313
rect 115 309 116 313
rect 190 311 191 315
rect 195 311 196 315
rect 190 310 196 311
rect 222 315 228 316
rect 222 311 223 315
rect 227 311 228 315
rect 222 310 228 311
rect 254 315 260 316
rect 254 311 255 315
rect 259 311 260 315
rect 254 310 260 311
rect 294 315 300 316
rect 294 311 295 315
rect 299 311 300 315
rect 294 310 300 311
rect 110 308 116 309
rect 170 307 176 308
rect 170 303 171 307
rect 175 303 176 307
rect 170 302 176 303
rect 110 296 116 297
rect 110 292 111 296
rect 115 292 116 296
rect 110 291 116 292
rect 112 283 114 291
rect 111 282 115 283
rect 111 277 115 278
rect 151 282 155 283
rect 151 277 155 278
rect 112 273 114 277
rect 110 272 116 273
rect 152 272 154 277
rect 172 276 174 302
rect 190 297 196 298
rect 190 293 191 297
rect 195 293 196 297
rect 190 292 196 293
rect 222 297 228 298
rect 222 293 223 297
rect 227 293 228 297
rect 222 292 228 293
rect 254 297 260 298
rect 254 293 255 297
rect 259 293 260 297
rect 254 292 260 293
rect 294 297 300 298
rect 294 293 295 297
rect 299 293 300 297
rect 294 292 300 293
rect 312 292 314 330
rect 334 329 340 330
rect 334 325 335 329
rect 339 325 340 329
rect 334 324 340 325
rect 390 329 396 330
rect 390 325 391 329
rect 395 325 396 329
rect 390 324 396 325
rect 400 329 406 331
rect 446 329 452 330
rect 335 322 339 324
rect 335 316 339 318
rect 367 322 371 323
rect 367 316 371 318
rect 391 322 395 324
rect 391 317 395 318
rect 334 315 340 316
rect 334 311 335 315
rect 339 311 340 315
rect 334 310 340 311
rect 366 315 372 316
rect 366 311 367 315
rect 371 311 372 315
rect 366 310 372 311
rect 400 308 402 329
rect 446 325 447 329
rect 451 325 452 329
rect 446 324 452 325
rect 438 323 444 324
rect 407 322 411 323
rect 438 319 439 323
rect 443 319 444 323
rect 438 318 444 319
rect 447 322 451 324
rect 407 316 411 318
rect 406 315 412 316
rect 406 311 407 315
rect 411 311 412 315
rect 406 310 412 311
rect 398 307 404 308
rect 398 303 399 307
rect 403 303 404 307
rect 398 302 404 303
rect 334 297 340 298
rect 334 293 335 297
rect 339 293 340 297
rect 334 292 340 293
rect 366 297 372 298
rect 366 293 367 297
rect 371 293 372 297
rect 366 292 372 293
rect 406 297 412 298
rect 406 293 407 297
rect 411 293 412 297
rect 406 292 412 293
rect 440 292 442 318
rect 447 317 451 318
rect 455 322 459 323
rect 455 316 459 318
rect 454 315 460 316
rect 454 311 455 315
rect 459 311 460 315
rect 454 310 460 311
rect 454 297 460 298
rect 454 293 455 297
rect 459 293 460 297
rect 454 292 460 293
rect 192 283 194 292
rect 224 283 226 292
rect 256 283 258 292
rect 296 283 298 292
rect 310 291 316 292
rect 310 287 311 291
rect 315 287 316 291
rect 310 286 316 287
rect 336 283 338 292
rect 342 291 348 292
rect 342 287 343 291
rect 347 287 348 291
rect 342 286 348 287
rect 183 282 187 283
rect 183 277 187 278
rect 191 282 195 283
rect 191 277 195 278
rect 215 282 219 283
rect 215 277 219 278
rect 223 282 227 283
rect 223 277 227 278
rect 247 282 251 283
rect 247 277 251 278
rect 255 282 259 283
rect 255 277 259 278
rect 279 282 283 283
rect 279 277 283 278
rect 295 282 299 283
rect 295 277 299 278
rect 311 282 315 283
rect 311 277 315 278
rect 335 282 339 283
rect 335 277 339 278
rect 170 275 176 276
rect 110 268 111 272
rect 115 268 116 272
rect 110 267 116 268
rect 150 271 156 272
rect 150 267 151 271
rect 155 267 156 271
rect 170 271 171 275
rect 175 271 176 275
rect 184 272 186 277
rect 216 272 218 277
rect 248 272 250 277
rect 266 275 272 276
rect 170 270 176 271
rect 182 271 188 272
rect 150 266 156 267
rect 182 267 183 271
rect 187 267 188 271
rect 182 266 188 267
rect 214 271 220 272
rect 214 267 215 271
rect 219 267 220 271
rect 214 266 220 267
rect 246 271 252 272
rect 246 267 247 271
rect 251 267 252 271
rect 266 271 267 275
rect 271 271 272 275
rect 280 272 282 277
rect 312 272 314 277
rect 266 270 272 271
rect 278 271 284 272
rect 246 266 252 267
rect 226 259 232 260
rect 110 255 116 256
rect 110 251 111 255
rect 115 251 116 255
rect 226 255 227 259
rect 231 255 232 259
rect 226 254 232 255
rect 110 250 116 251
rect 150 253 156 254
rect 112 247 114 250
rect 150 249 151 253
rect 155 249 156 253
rect 150 248 156 249
rect 182 253 188 254
rect 182 249 183 253
rect 187 249 188 253
rect 182 248 188 249
rect 214 253 220 254
rect 214 249 215 253
rect 219 249 220 253
rect 214 248 220 249
rect 111 246 115 247
rect 111 241 115 242
rect 135 246 139 247
rect 112 238 114 241
rect 135 240 139 242
rect 151 246 155 248
rect 151 241 155 242
rect 167 246 171 247
rect 167 240 171 242
rect 183 246 187 248
rect 183 241 187 242
rect 207 246 211 247
rect 207 240 211 242
rect 215 246 219 248
rect 215 241 219 242
rect 134 239 140 240
rect 110 237 116 238
rect 110 233 111 237
rect 115 233 116 237
rect 134 235 135 239
rect 139 235 140 239
rect 134 234 140 235
rect 166 239 172 240
rect 166 235 167 239
rect 171 235 172 239
rect 166 234 172 235
rect 206 239 212 240
rect 206 235 207 239
rect 211 235 212 239
rect 206 234 212 235
rect 110 232 116 233
rect 150 231 156 232
rect 150 227 151 231
rect 155 227 156 231
rect 150 226 156 227
rect 134 221 140 222
rect 110 220 116 221
rect 110 216 111 220
rect 115 216 116 220
rect 134 217 135 221
rect 139 217 140 221
rect 134 216 140 217
rect 110 215 116 216
rect 112 207 114 215
rect 136 207 138 216
rect 111 206 115 207
rect 111 201 115 202
rect 135 206 139 207
rect 135 201 139 202
rect 112 197 114 201
rect 110 196 116 197
rect 136 196 138 201
rect 152 200 154 226
rect 166 221 172 222
rect 166 217 167 221
rect 171 217 172 221
rect 166 216 172 217
rect 206 221 212 222
rect 206 217 207 221
rect 211 217 212 221
rect 206 216 212 217
rect 228 216 230 254
rect 246 253 252 254
rect 246 249 247 253
rect 251 249 252 253
rect 246 248 252 249
rect 247 246 251 248
rect 247 241 251 242
rect 255 246 259 247
rect 255 240 259 242
rect 254 239 260 240
rect 254 235 255 239
rect 259 235 260 239
rect 254 234 260 235
rect 268 232 270 270
rect 278 267 279 271
rect 283 267 284 271
rect 278 266 284 267
rect 310 271 316 272
rect 310 267 311 271
rect 315 267 316 271
rect 310 266 316 267
rect 344 260 346 286
rect 368 283 370 292
rect 408 283 410 292
rect 438 291 444 292
rect 438 287 439 291
rect 443 287 444 291
rect 438 286 444 287
rect 456 283 458 292
rect 496 284 498 346
rect 502 343 503 347
rect 507 343 508 347
rect 502 342 508 343
rect 566 347 572 348
rect 566 343 567 347
rect 571 343 572 347
rect 566 342 572 343
rect 502 329 508 330
rect 502 325 503 329
rect 507 325 508 329
rect 502 324 508 325
rect 566 329 572 330
rect 566 325 567 329
rect 571 325 572 329
rect 566 324 572 325
rect 576 324 578 358
rect 599 353 603 354
rect 631 358 635 359
rect 631 353 635 354
rect 655 358 659 359
rect 655 353 659 354
rect 687 358 691 359
rect 687 353 691 354
rect 703 358 707 359
rect 703 353 707 354
rect 751 358 755 359
rect 751 353 755 354
rect 807 358 811 359
rect 807 353 811 354
rect 815 358 819 359
rect 826 358 832 359
rect 863 358 867 359
rect 815 353 819 354
rect 863 353 867 354
rect 879 358 883 359
rect 879 353 883 354
rect 919 358 923 359
rect 919 353 923 354
rect 951 358 955 359
rect 951 353 955 354
rect 983 358 987 359
rect 983 353 987 354
rect 1031 358 1035 359
rect 1031 353 1035 354
rect 1055 358 1059 359
rect 1072 356 1074 374
rect 1126 369 1132 370
rect 1126 365 1127 369
rect 1131 365 1132 369
rect 1126 364 1132 365
rect 1160 364 1162 390
rect 1199 388 1203 390
rect 1223 394 1227 396
rect 1223 389 1227 390
rect 1271 394 1275 395
rect 1271 388 1275 390
rect 1303 394 1307 396
rect 1303 389 1307 390
rect 1343 394 1347 395
rect 1343 388 1347 390
rect 1383 394 1387 396
rect 1383 389 1387 390
rect 1415 394 1419 395
rect 1415 388 1419 390
rect 1471 394 1475 396
rect 1471 389 1475 390
rect 1487 394 1491 395
rect 1487 388 1491 390
rect 1198 387 1204 388
rect 1198 383 1199 387
rect 1203 383 1204 387
rect 1198 382 1204 383
rect 1270 387 1276 388
rect 1270 383 1271 387
rect 1275 383 1276 387
rect 1270 382 1276 383
rect 1342 387 1348 388
rect 1342 383 1343 387
rect 1347 383 1348 387
rect 1342 382 1348 383
rect 1414 387 1420 388
rect 1414 383 1415 387
rect 1419 383 1420 387
rect 1414 382 1420 383
rect 1486 387 1492 388
rect 1486 383 1487 387
rect 1491 383 1492 387
rect 1486 382 1492 383
rect 1504 380 1506 418
rect 1542 415 1543 419
rect 1547 415 1548 419
rect 1558 419 1559 423
rect 1563 419 1564 423
rect 1584 421 1586 425
rect 1558 418 1564 419
rect 1582 420 1588 421
rect 1582 416 1583 420
rect 1587 416 1588 420
rect 1582 415 1588 416
rect 1542 414 1548 415
rect 1558 407 1564 408
rect 1558 403 1559 407
rect 1563 403 1564 407
rect 1558 402 1564 403
rect 1582 403 1588 404
rect 1542 401 1548 402
rect 1542 397 1543 401
rect 1547 397 1548 401
rect 1542 396 1548 397
rect 1543 394 1547 396
rect 1543 388 1547 390
rect 1542 387 1548 388
rect 1542 383 1543 387
rect 1547 383 1548 387
rect 1542 382 1548 383
rect 1354 379 1360 380
rect 1354 375 1355 379
rect 1359 375 1360 379
rect 1354 374 1360 375
rect 1502 379 1508 380
rect 1502 375 1503 379
rect 1507 375 1508 379
rect 1502 374 1508 375
rect 1198 369 1204 370
rect 1198 365 1199 369
rect 1203 365 1204 369
rect 1198 364 1204 365
rect 1270 369 1276 370
rect 1270 365 1271 369
rect 1275 365 1276 369
rect 1270 364 1276 365
rect 1342 369 1348 370
rect 1342 365 1343 369
rect 1347 365 1348 369
rect 1342 364 1348 365
rect 1128 359 1130 364
rect 1158 363 1164 364
rect 1158 359 1159 363
rect 1163 359 1164 363
rect 1200 359 1202 364
rect 1272 359 1274 364
rect 1344 359 1346 364
rect 1103 358 1107 359
rect 1055 353 1059 354
rect 1070 355 1076 356
rect 632 348 634 353
rect 688 348 690 353
rect 752 348 754 353
rect 816 348 818 353
rect 880 348 882 353
rect 952 348 954 353
rect 1032 348 1034 353
rect 1070 351 1071 355
rect 1075 351 1076 355
rect 1103 353 1107 354
rect 1127 358 1131 359
rect 1158 358 1164 359
rect 1175 358 1179 359
rect 1127 353 1131 354
rect 1175 353 1179 354
rect 1199 358 1203 359
rect 1199 353 1203 354
rect 1247 358 1251 359
rect 1247 353 1251 354
rect 1271 358 1275 359
rect 1271 353 1275 354
rect 1327 358 1331 359
rect 1327 353 1331 354
rect 1343 358 1347 359
rect 1343 353 1347 354
rect 1070 350 1076 351
rect 1104 348 1106 353
rect 1176 348 1178 353
rect 1248 348 1250 353
rect 1328 348 1330 353
rect 1356 352 1358 374
rect 1414 369 1420 370
rect 1414 365 1415 369
rect 1419 365 1420 369
rect 1414 364 1420 365
rect 1486 369 1492 370
rect 1486 365 1487 369
rect 1491 365 1492 369
rect 1486 364 1492 365
rect 1542 369 1548 370
rect 1542 365 1543 369
rect 1547 365 1548 369
rect 1542 364 1548 365
rect 1560 364 1562 402
rect 1582 399 1583 403
rect 1587 399 1588 403
rect 1582 398 1588 399
rect 1584 395 1586 398
rect 1583 394 1587 395
rect 1583 389 1587 390
rect 1584 386 1586 389
rect 1582 385 1588 386
rect 1582 381 1583 385
rect 1587 381 1588 385
rect 1582 380 1588 381
rect 1582 368 1588 369
rect 1582 364 1583 368
rect 1587 364 1588 368
rect 1416 359 1418 364
rect 1426 363 1432 364
rect 1426 359 1427 363
rect 1431 359 1432 363
rect 1488 359 1490 364
rect 1544 359 1546 364
rect 1558 363 1564 364
rect 1582 363 1588 364
rect 1558 359 1559 363
rect 1563 359 1564 363
rect 1584 359 1586 363
rect 1407 358 1411 359
rect 1407 353 1411 354
rect 1415 358 1419 359
rect 1426 358 1432 359
rect 1487 358 1491 359
rect 1415 353 1419 354
rect 1354 351 1360 352
rect 630 347 636 348
rect 630 343 631 347
rect 635 343 636 347
rect 630 342 636 343
rect 686 347 692 348
rect 686 343 687 347
rect 691 343 692 347
rect 686 342 692 343
rect 750 347 756 348
rect 750 343 751 347
rect 755 343 756 347
rect 750 342 756 343
rect 814 347 820 348
rect 814 343 815 347
rect 819 343 820 347
rect 814 342 820 343
rect 878 347 884 348
rect 878 343 879 347
rect 883 343 884 347
rect 878 342 884 343
rect 950 347 956 348
rect 950 343 951 347
rect 955 343 956 347
rect 950 342 956 343
rect 1030 347 1036 348
rect 1030 343 1031 347
rect 1035 343 1036 347
rect 1030 342 1036 343
rect 1102 347 1108 348
rect 1102 343 1103 347
rect 1107 343 1108 347
rect 1102 342 1108 343
rect 1174 347 1180 348
rect 1174 343 1175 347
rect 1179 343 1180 347
rect 1174 342 1180 343
rect 1246 347 1252 348
rect 1246 343 1247 347
rect 1251 343 1252 347
rect 1246 342 1252 343
rect 1326 347 1332 348
rect 1326 343 1327 347
rect 1331 343 1332 347
rect 1354 347 1355 351
rect 1359 347 1360 351
rect 1408 348 1410 353
rect 1354 346 1360 347
rect 1406 347 1412 348
rect 1326 342 1332 343
rect 1406 343 1407 347
rect 1411 343 1412 347
rect 1406 342 1412 343
rect 1428 336 1430 358
rect 1487 353 1491 354
rect 1543 358 1547 359
rect 1558 358 1564 359
rect 1583 358 1587 359
rect 1543 353 1547 354
rect 1583 353 1587 354
rect 1488 348 1490 353
rect 1498 351 1504 352
rect 1486 347 1492 348
rect 1486 343 1487 347
rect 1491 343 1492 347
rect 1498 347 1499 351
rect 1503 347 1504 351
rect 1544 348 1546 353
rect 1584 349 1586 353
rect 1582 348 1588 349
rect 1498 346 1504 347
rect 1542 347 1548 348
rect 1486 342 1492 343
rect 1238 335 1244 336
rect 1238 331 1239 335
rect 1243 331 1244 335
rect 1238 330 1244 331
rect 1426 335 1432 336
rect 1426 331 1427 335
rect 1431 331 1432 335
rect 1426 330 1432 331
rect 630 329 636 330
rect 630 325 631 329
rect 635 325 636 329
rect 630 324 636 325
rect 686 329 692 330
rect 686 325 687 329
rect 691 325 692 329
rect 686 324 692 325
rect 750 329 756 330
rect 750 325 751 329
rect 755 325 756 329
rect 750 324 756 325
rect 814 329 820 330
rect 814 325 815 329
rect 819 325 820 329
rect 814 324 820 325
rect 878 329 884 330
rect 878 325 879 329
rect 883 325 884 329
rect 878 324 884 325
rect 950 329 956 330
rect 950 325 951 329
rect 955 325 956 329
rect 950 324 956 325
rect 1030 329 1036 330
rect 1030 325 1031 329
rect 1035 325 1036 329
rect 1030 324 1036 325
rect 1102 329 1108 330
rect 1102 325 1103 329
rect 1107 325 1108 329
rect 1102 324 1108 325
rect 1174 329 1180 330
rect 1174 325 1175 329
rect 1179 325 1180 329
rect 1174 324 1180 325
rect 503 322 507 324
rect 503 317 507 318
rect 519 322 523 323
rect 519 316 523 318
rect 567 322 571 324
rect 574 323 580 324
rect 574 319 575 323
rect 579 319 580 323
rect 574 318 580 319
rect 591 322 595 323
rect 567 317 571 318
rect 591 316 595 318
rect 631 322 635 324
rect 631 317 635 318
rect 663 322 667 323
rect 663 316 667 318
rect 687 322 691 324
rect 687 317 691 318
rect 735 322 739 323
rect 735 316 739 318
rect 751 322 755 324
rect 751 317 755 318
rect 807 322 811 323
rect 807 316 811 318
rect 815 322 819 324
rect 826 323 832 324
rect 826 319 827 323
rect 831 319 832 323
rect 826 318 832 319
rect 879 322 883 324
rect 815 317 819 318
rect 518 315 524 316
rect 518 311 519 315
rect 523 311 524 315
rect 518 310 524 311
rect 590 315 596 316
rect 590 311 591 315
rect 595 311 596 315
rect 590 310 596 311
rect 662 315 668 316
rect 662 311 663 315
rect 667 311 668 315
rect 662 310 668 311
rect 734 315 740 316
rect 734 311 735 315
rect 739 311 740 315
rect 734 310 740 311
rect 806 315 812 316
rect 806 311 807 315
rect 811 311 812 315
rect 806 310 812 311
rect 722 307 728 308
rect 722 303 723 307
rect 727 303 728 307
rect 722 302 728 303
rect 654 299 660 300
rect 518 297 524 298
rect 518 293 519 297
rect 523 293 524 297
rect 518 292 524 293
rect 590 297 596 298
rect 590 293 591 297
rect 595 293 596 297
rect 654 295 655 299
rect 659 295 660 299
rect 654 294 660 295
rect 662 297 668 298
rect 590 292 596 293
rect 494 283 500 284
rect 520 283 522 292
rect 592 283 594 292
rect 351 282 355 283
rect 351 277 355 278
rect 367 282 371 283
rect 367 277 371 278
rect 407 282 411 283
rect 407 277 411 278
rect 455 282 459 283
rect 455 277 459 278
rect 479 282 483 283
rect 494 279 495 283
rect 499 279 500 283
rect 494 278 500 279
rect 519 282 523 283
rect 479 277 483 278
rect 519 277 523 278
rect 559 282 563 283
rect 559 277 563 278
rect 591 282 595 283
rect 591 277 595 278
rect 647 282 651 283
rect 647 277 651 278
rect 352 272 354 277
rect 398 275 404 276
rect 350 271 356 272
rect 350 267 351 271
rect 355 267 356 271
rect 398 271 399 275
rect 403 271 404 275
rect 408 272 410 277
rect 480 272 482 277
rect 560 272 562 277
rect 648 272 650 277
rect 398 270 404 271
rect 406 271 412 272
rect 350 266 356 267
rect 342 259 348 260
rect 342 255 343 259
rect 347 255 348 259
rect 342 254 348 255
rect 278 253 284 254
rect 278 249 279 253
rect 283 249 284 253
rect 278 248 284 249
rect 310 253 316 254
rect 310 249 311 253
rect 315 249 316 253
rect 310 248 316 249
rect 350 253 356 254
rect 350 249 351 253
rect 355 249 356 253
rect 350 248 356 249
rect 279 246 283 248
rect 279 241 283 242
rect 303 246 307 247
rect 303 240 307 242
rect 311 246 315 248
rect 311 241 315 242
rect 343 246 347 247
rect 343 240 347 242
rect 351 246 355 248
rect 351 241 355 242
rect 383 246 387 247
rect 383 240 387 242
rect 302 239 308 240
rect 302 235 303 239
rect 307 235 308 239
rect 302 234 308 235
rect 342 239 348 240
rect 342 235 343 239
rect 347 235 348 239
rect 342 234 348 235
rect 382 239 388 240
rect 382 235 383 239
rect 387 235 388 239
rect 382 234 388 235
rect 400 232 402 270
rect 406 267 407 271
rect 411 267 412 271
rect 406 266 412 267
rect 478 271 484 272
rect 478 267 479 271
rect 483 267 484 271
rect 478 266 484 267
rect 558 271 564 272
rect 558 267 559 271
rect 563 267 564 271
rect 558 266 564 267
rect 646 271 652 272
rect 646 267 647 271
rect 651 267 652 271
rect 646 266 652 267
rect 406 253 412 254
rect 406 249 407 253
rect 411 249 412 253
rect 406 248 412 249
rect 478 253 484 254
rect 478 249 479 253
rect 483 249 484 253
rect 478 248 484 249
rect 558 253 564 254
rect 558 249 559 253
rect 563 249 564 253
rect 558 248 564 249
rect 646 253 652 254
rect 646 249 647 253
rect 651 249 652 253
rect 646 248 652 249
rect 656 248 658 294
rect 662 293 663 297
rect 667 293 668 297
rect 662 292 668 293
rect 664 283 666 292
rect 724 284 726 302
rect 734 297 740 298
rect 734 293 735 297
rect 739 293 740 297
rect 734 292 740 293
rect 806 297 812 298
rect 806 293 807 297
rect 811 293 812 297
rect 806 292 812 293
rect 828 292 830 318
rect 879 316 883 318
rect 951 322 955 324
rect 951 316 955 318
rect 1023 322 1027 323
rect 1023 316 1027 318
rect 1031 322 1035 324
rect 1031 317 1035 318
rect 1095 322 1099 323
rect 1095 316 1099 318
rect 1103 322 1107 324
rect 1103 317 1107 318
rect 1167 322 1171 323
rect 1167 316 1171 318
rect 1175 322 1179 324
rect 1175 317 1179 318
rect 1231 322 1235 323
rect 1231 316 1235 318
rect 878 315 884 316
rect 878 311 879 315
rect 883 311 884 315
rect 878 310 884 311
rect 950 315 956 316
rect 950 311 951 315
rect 955 311 956 315
rect 950 310 956 311
rect 1022 315 1028 316
rect 1022 311 1023 315
rect 1027 311 1028 315
rect 1022 310 1028 311
rect 1094 315 1100 316
rect 1094 311 1095 315
rect 1099 311 1100 315
rect 1094 310 1100 311
rect 1110 315 1116 316
rect 1110 311 1111 315
rect 1115 311 1116 315
rect 1110 310 1116 311
rect 1166 315 1172 316
rect 1166 311 1167 315
rect 1171 311 1172 315
rect 1166 310 1172 311
rect 1230 315 1236 316
rect 1230 311 1231 315
rect 1235 311 1236 315
rect 1230 310 1236 311
rect 878 297 884 298
rect 878 293 879 297
rect 883 293 884 297
rect 878 292 884 293
rect 950 297 956 298
rect 950 293 951 297
rect 955 293 956 297
rect 950 292 956 293
rect 1022 297 1028 298
rect 1022 293 1023 297
rect 1027 293 1028 297
rect 1022 292 1028 293
rect 1094 297 1100 298
rect 1094 293 1095 297
rect 1099 293 1100 297
rect 1094 292 1100 293
rect 722 283 728 284
rect 736 283 738 292
rect 808 283 810 292
rect 826 291 832 292
rect 826 287 827 291
rect 831 287 832 291
rect 826 286 832 287
rect 880 283 882 292
rect 952 283 954 292
rect 1024 283 1026 292
rect 1096 283 1098 292
rect 1112 284 1114 310
rect 1166 297 1172 298
rect 1166 293 1167 297
rect 1171 293 1172 297
rect 1166 292 1172 293
rect 1230 297 1236 298
rect 1230 293 1231 297
rect 1235 293 1236 297
rect 1230 292 1236 293
rect 1240 292 1242 330
rect 1246 329 1252 330
rect 1246 325 1247 329
rect 1251 325 1252 329
rect 1246 324 1252 325
rect 1326 329 1332 330
rect 1326 325 1327 329
rect 1331 325 1332 329
rect 1326 324 1332 325
rect 1406 329 1412 330
rect 1406 325 1407 329
rect 1411 325 1412 329
rect 1406 324 1412 325
rect 1486 329 1492 330
rect 1486 325 1487 329
rect 1491 325 1492 329
rect 1486 324 1492 325
rect 1247 322 1251 324
rect 1247 317 1251 318
rect 1295 322 1299 323
rect 1295 316 1299 318
rect 1327 322 1331 324
rect 1327 317 1331 318
rect 1351 322 1355 323
rect 1351 316 1355 318
rect 1399 322 1403 323
rect 1399 316 1403 318
rect 1407 322 1411 324
rect 1407 317 1411 318
rect 1455 322 1459 323
rect 1455 316 1459 318
rect 1487 322 1491 324
rect 1487 317 1491 318
rect 1294 315 1300 316
rect 1294 311 1295 315
rect 1299 311 1300 315
rect 1294 310 1300 311
rect 1350 315 1356 316
rect 1350 311 1351 315
rect 1355 311 1356 315
rect 1350 310 1356 311
rect 1398 315 1404 316
rect 1398 311 1399 315
rect 1403 311 1404 315
rect 1398 310 1404 311
rect 1454 315 1460 316
rect 1454 311 1455 315
rect 1459 311 1460 315
rect 1454 310 1460 311
rect 1500 308 1502 346
rect 1542 343 1543 347
rect 1547 343 1548 347
rect 1582 344 1583 348
rect 1587 344 1588 348
rect 1582 343 1588 344
rect 1542 342 1548 343
rect 1530 339 1536 340
rect 1530 335 1531 339
rect 1535 335 1536 339
rect 1530 334 1536 335
rect 1511 322 1515 323
rect 1511 316 1515 318
rect 1510 315 1516 316
rect 1510 311 1511 315
rect 1515 311 1516 315
rect 1510 310 1516 311
rect 1286 307 1292 308
rect 1286 303 1287 307
rect 1291 303 1292 307
rect 1286 302 1292 303
rect 1498 307 1504 308
rect 1498 303 1499 307
rect 1503 303 1504 307
rect 1498 302 1504 303
rect 1110 283 1116 284
rect 1168 283 1170 292
rect 1232 283 1234 292
rect 1238 291 1244 292
rect 1238 287 1239 291
rect 1243 287 1244 291
rect 1238 286 1244 287
rect 1288 284 1290 302
rect 1294 297 1300 298
rect 1294 293 1295 297
rect 1299 293 1300 297
rect 1294 292 1300 293
rect 1350 297 1356 298
rect 1350 293 1351 297
rect 1355 293 1356 297
rect 1350 292 1356 293
rect 1398 297 1404 298
rect 1398 293 1399 297
rect 1403 293 1404 297
rect 1398 292 1404 293
rect 1454 297 1460 298
rect 1454 293 1455 297
rect 1459 293 1460 297
rect 1454 292 1460 293
rect 1510 297 1516 298
rect 1510 293 1511 297
rect 1515 293 1516 297
rect 1510 292 1516 293
rect 1532 292 1534 334
rect 1582 331 1588 332
rect 1542 329 1548 330
rect 1542 325 1543 329
rect 1547 325 1548 329
rect 1582 327 1583 331
rect 1587 327 1588 331
rect 1582 326 1588 327
rect 1542 324 1548 325
rect 1543 322 1547 324
rect 1584 323 1586 326
rect 1543 316 1547 318
rect 1583 322 1587 323
rect 1583 317 1587 318
rect 1542 315 1548 316
rect 1542 311 1543 315
rect 1547 311 1548 315
rect 1584 314 1586 317
rect 1542 310 1548 311
rect 1582 313 1588 314
rect 1582 309 1583 313
rect 1587 309 1588 313
rect 1582 308 1588 309
rect 1558 307 1564 308
rect 1558 303 1559 307
rect 1563 303 1564 307
rect 1558 302 1564 303
rect 1542 297 1548 298
rect 1542 293 1543 297
rect 1547 293 1548 297
rect 1542 292 1548 293
rect 1286 283 1292 284
rect 1296 283 1298 292
rect 1352 283 1354 292
rect 1400 283 1402 292
rect 1456 283 1458 292
rect 1512 283 1514 292
rect 1530 291 1536 292
rect 1530 287 1531 291
rect 1535 287 1536 291
rect 1530 286 1536 287
rect 1544 283 1546 292
rect 663 282 667 283
rect 722 279 723 283
rect 727 279 728 283
rect 722 278 728 279
rect 735 282 739 283
rect 663 277 667 278
rect 735 277 739 278
rect 807 282 811 283
rect 807 277 811 278
rect 823 282 827 283
rect 823 277 827 278
rect 879 282 883 283
rect 879 277 883 278
rect 903 282 907 283
rect 903 277 907 278
rect 951 282 955 283
rect 951 277 955 278
rect 983 282 987 283
rect 983 277 987 278
rect 1023 282 1027 283
rect 1023 277 1027 278
rect 1055 282 1059 283
rect 1055 277 1059 278
rect 1095 282 1099 283
rect 1110 279 1111 283
rect 1115 279 1116 283
rect 1110 278 1116 279
rect 1119 282 1123 283
rect 1095 277 1099 278
rect 1119 277 1123 278
rect 1167 282 1171 283
rect 1167 277 1171 278
rect 1175 282 1179 283
rect 1175 277 1179 278
rect 1223 282 1227 283
rect 1223 277 1227 278
rect 1231 282 1235 283
rect 1231 277 1235 278
rect 1263 282 1267 283
rect 1286 279 1287 283
rect 1291 279 1292 283
rect 1286 278 1292 279
rect 1295 282 1299 283
rect 1263 277 1267 278
rect 1295 277 1299 278
rect 1303 282 1307 283
rect 1303 277 1307 278
rect 1351 282 1355 283
rect 1351 277 1355 278
rect 1399 282 1403 283
rect 1399 277 1403 278
rect 1447 282 1451 283
rect 1447 277 1451 278
rect 1455 282 1459 283
rect 1455 277 1459 278
rect 1503 282 1507 283
rect 1503 277 1507 278
rect 1511 282 1515 283
rect 1511 277 1515 278
rect 1543 282 1547 283
rect 1543 277 1547 278
rect 736 272 738 277
rect 824 272 826 277
rect 904 272 906 277
rect 984 272 986 277
rect 1056 272 1058 277
rect 1120 272 1122 277
rect 1176 272 1178 277
rect 1224 272 1226 277
rect 1264 272 1266 277
rect 1304 272 1306 277
rect 1352 272 1354 277
rect 1400 272 1402 277
rect 1448 272 1450 277
rect 1504 272 1506 277
rect 1518 275 1524 276
rect 734 271 740 272
rect 734 267 735 271
rect 739 267 740 271
rect 734 266 740 267
rect 822 271 828 272
rect 822 267 823 271
rect 827 267 828 271
rect 822 266 828 267
rect 902 271 908 272
rect 902 267 903 271
rect 907 267 908 271
rect 902 266 908 267
rect 982 271 988 272
rect 982 267 983 271
rect 987 267 988 271
rect 982 266 988 267
rect 1054 271 1060 272
rect 1054 267 1055 271
rect 1059 267 1060 271
rect 1054 266 1060 267
rect 1118 271 1124 272
rect 1118 267 1119 271
rect 1123 267 1124 271
rect 1118 266 1124 267
rect 1174 271 1180 272
rect 1174 267 1175 271
rect 1179 267 1180 271
rect 1174 266 1180 267
rect 1222 271 1228 272
rect 1222 267 1223 271
rect 1227 267 1228 271
rect 1222 266 1228 267
rect 1262 271 1268 272
rect 1262 267 1263 271
rect 1267 267 1268 271
rect 1262 266 1268 267
rect 1302 271 1308 272
rect 1302 267 1303 271
rect 1307 267 1308 271
rect 1302 266 1308 267
rect 1350 271 1356 272
rect 1350 267 1351 271
rect 1355 267 1356 271
rect 1350 266 1356 267
rect 1398 271 1404 272
rect 1398 267 1399 271
rect 1403 267 1404 271
rect 1398 266 1404 267
rect 1446 271 1452 272
rect 1446 267 1447 271
rect 1451 267 1452 271
rect 1446 266 1452 267
rect 1502 271 1508 272
rect 1502 267 1503 271
rect 1507 267 1508 271
rect 1518 271 1519 275
rect 1523 271 1524 275
rect 1544 272 1546 277
rect 1560 276 1562 302
rect 1582 296 1588 297
rect 1582 292 1583 296
rect 1587 292 1588 296
rect 1582 291 1588 292
rect 1584 283 1586 291
rect 1583 282 1587 283
rect 1583 277 1587 278
rect 1558 275 1564 276
rect 1518 270 1524 271
rect 1542 271 1548 272
rect 1502 266 1508 267
rect 1186 259 1192 260
rect 1186 255 1187 259
rect 1191 255 1192 259
rect 1186 254 1192 255
rect 1362 259 1368 260
rect 1362 255 1363 259
rect 1367 255 1368 259
rect 1362 254 1368 255
rect 734 253 740 254
rect 734 249 735 253
rect 739 249 740 253
rect 734 248 740 249
rect 822 253 828 254
rect 822 249 823 253
rect 827 249 828 253
rect 822 248 828 249
rect 902 253 908 254
rect 902 249 903 253
rect 907 249 908 253
rect 902 248 908 249
rect 982 253 988 254
rect 982 249 983 253
rect 987 249 988 253
rect 982 248 988 249
rect 1054 253 1060 254
rect 1054 249 1055 253
rect 1059 249 1060 253
rect 1054 248 1060 249
rect 1118 253 1124 254
rect 1118 249 1119 253
rect 1123 249 1124 253
rect 1118 248 1124 249
rect 1174 253 1180 254
rect 1174 249 1175 253
rect 1179 249 1180 253
rect 1174 248 1180 249
rect 407 246 411 248
rect 462 247 468 248
rect 407 241 411 242
rect 439 246 443 247
rect 462 243 463 247
rect 467 243 468 247
rect 462 242 468 243
rect 479 246 483 248
rect 439 240 443 242
rect 438 239 444 240
rect 438 235 439 239
rect 443 235 444 239
rect 438 234 444 235
rect 266 231 272 232
rect 266 227 267 231
rect 271 227 272 231
rect 266 226 272 227
rect 398 231 404 232
rect 398 227 399 231
rect 403 227 404 231
rect 398 226 404 227
rect 254 221 260 222
rect 254 217 255 221
rect 259 217 260 221
rect 254 216 260 217
rect 302 221 308 222
rect 302 217 303 221
rect 307 217 308 221
rect 302 216 308 217
rect 342 221 348 222
rect 342 217 343 221
rect 347 217 348 221
rect 342 216 348 217
rect 382 221 388 222
rect 382 217 383 221
rect 387 217 388 221
rect 382 216 388 217
rect 438 221 444 222
rect 438 217 439 221
rect 443 217 444 221
rect 438 216 444 217
rect 168 207 170 216
rect 208 207 210 216
rect 226 215 232 216
rect 226 211 227 215
rect 231 211 232 215
rect 226 210 232 211
rect 256 207 258 216
rect 304 207 306 216
rect 344 207 346 216
rect 374 215 380 216
rect 374 211 375 215
rect 379 211 380 215
rect 374 210 380 211
rect 167 206 171 207
rect 167 201 171 202
rect 207 206 211 207
rect 207 201 211 202
rect 215 206 219 207
rect 215 201 219 202
rect 255 206 259 207
rect 255 201 259 202
rect 263 206 267 207
rect 263 201 267 202
rect 303 206 307 207
rect 303 201 307 202
rect 311 206 315 207
rect 311 201 315 202
rect 343 206 347 207
rect 343 201 347 202
rect 359 206 363 207
rect 359 201 363 202
rect 150 199 156 200
rect 110 192 111 196
rect 115 192 116 196
rect 110 191 116 192
rect 134 195 140 196
rect 134 191 135 195
rect 139 191 140 195
rect 150 195 151 199
rect 155 195 156 199
rect 168 196 170 201
rect 216 196 218 201
rect 264 196 266 201
rect 312 196 314 201
rect 322 199 328 200
rect 150 194 156 195
rect 166 195 172 196
rect 134 190 140 191
rect 166 191 167 195
rect 171 191 172 195
rect 166 190 172 191
rect 214 195 220 196
rect 214 191 215 195
rect 219 191 220 195
rect 214 190 220 191
rect 262 195 268 196
rect 262 191 263 195
rect 267 191 268 195
rect 262 190 268 191
rect 310 195 316 196
rect 310 191 311 195
rect 315 191 316 195
rect 322 195 323 199
rect 327 195 328 199
rect 360 196 362 201
rect 322 194 328 195
rect 358 195 364 196
rect 310 190 316 191
rect 274 183 280 184
rect 110 179 116 180
rect 110 175 111 179
rect 115 175 116 179
rect 274 179 275 183
rect 279 179 280 183
rect 274 178 280 179
rect 110 174 116 175
rect 134 177 140 178
rect 112 171 114 174
rect 134 173 135 177
rect 139 173 140 177
rect 134 172 140 173
rect 166 177 172 178
rect 166 173 167 177
rect 171 173 172 177
rect 166 172 172 173
rect 214 177 220 178
rect 214 173 215 177
rect 219 173 220 177
rect 214 172 220 173
rect 262 177 268 178
rect 262 173 263 177
rect 267 173 268 177
rect 262 172 268 173
rect 111 170 115 171
rect 111 165 115 166
rect 135 170 139 172
rect 135 165 139 166
rect 143 170 147 171
rect 112 162 114 165
rect 143 164 147 166
rect 167 170 171 172
rect 167 165 171 166
rect 191 170 195 171
rect 191 164 195 166
rect 215 170 219 172
rect 215 165 219 166
rect 239 170 243 171
rect 239 164 243 166
rect 263 170 267 172
rect 263 165 267 166
rect 142 163 148 164
rect 110 161 116 162
rect 110 157 111 161
rect 115 157 116 161
rect 142 159 143 163
rect 147 159 148 163
rect 142 158 148 159
rect 190 163 196 164
rect 190 159 191 163
rect 195 159 196 163
rect 190 158 196 159
rect 238 163 244 164
rect 238 159 239 163
rect 243 159 244 163
rect 238 158 244 159
rect 110 156 116 157
rect 154 155 160 156
rect 154 151 155 155
rect 159 151 160 155
rect 154 150 160 151
rect 142 145 148 146
rect 110 144 116 145
rect 110 140 111 144
rect 115 140 116 144
rect 142 141 143 145
rect 147 141 148 145
rect 142 140 148 141
rect 110 139 116 140
rect 112 123 114 139
rect 144 123 146 140
rect 111 122 115 123
rect 111 117 115 118
rect 135 122 139 123
rect 135 117 139 118
rect 143 122 147 123
rect 143 117 147 118
rect 112 113 114 117
rect 110 112 116 113
rect 136 112 138 117
rect 156 116 158 150
rect 190 145 196 146
rect 190 141 191 145
rect 195 141 196 145
rect 190 140 196 141
rect 238 145 244 146
rect 238 141 239 145
rect 243 141 244 145
rect 238 140 244 141
rect 276 140 278 178
rect 310 177 316 178
rect 310 173 311 177
rect 315 173 316 177
rect 310 172 316 173
rect 295 170 299 171
rect 295 164 299 166
rect 311 170 315 172
rect 311 165 315 166
rect 294 163 300 164
rect 294 159 295 163
rect 299 159 300 163
rect 294 158 300 159
rect 324 156 326 194
rect 358 191 359 195
rect 363 191 364 195
rect 358 190 364 191
rect 376 184 378 210
rect 384 207 386 216
rect 440 207 442 216
rect 383 206 387 207
rect 383 201 387 202
rect 415 206 419 207
rect 415 201 419 202
rect 439 206 443 207
rect 439 201 443 202
rect 416 196 418 201
rect 464 200 466 242
rect 479 241 483 242
rect 511 246 515 247
rect 511 240 515 242
rect 559 246 563 248
rect 559 241 563 242
rect 591 246 595 247
rect 591 240 595 242
rect 647 246 651 248
rect 654 247 660 248
rect 654 243 655 247
rect 659 243 660 247
rect 654 242 660 243
rect 679 246 683 247
rect 647 241 651 242
rect 679 240 683 242
rect 735 246 739 248
rect 735 241 739 242
rect 767 246 771 247
rect 767 240 771 242
rect 823 246 827 248
rect 823 241 827 242
rect 847 246 851 247
rect 847 240 851 242
rect 903 246 907 248
rect 903 241 907 242
rect 919 246 923 247
rect 919 240 923 242
rect 983 246 987 248
rect 983 240 987 242
rect 1047 246 1051 247
rect 1047 240 1051 242
rect 1055 246 1059 248
rect 1055 241 1059 242
rect 1103 246 1107 247
rect 1103 240 1107 242
rect 1119 246 1123 248
rect 1119 241 1123 242
rect 1159 246 1163 247
rect 1159 240 1163 242
rect 1175 246 1179 248
rect 1175 241 1179 242
rect 510 239 516 240
rect 510 235 511 239
rect 515 235 516 239
rect 510 234 516 235
rect 590 239 596 240
rect 590 235 591 239
rect 595 235 596 239
rect 590 234 596 235
rect 678 239 684 240
rect 678 235 679 239
rect 683 235 684 239
rect 678 234 684 235
rect 758 239 764 240
rect 758 235 759 239
rect 763 235 764 239
rect 758 234 764 235
rect 766 239 772 240
rect 766 235 767 239
rect 771 235 772 239
rect 766 234 772 235
rect 846 239 852 240
rect 846 235 847 239
rect 851 235 852 239
rect 846 234 852 235
rect 918 239 924 240
rect 918 235 919 239
rect 923 235 924 239
rect 918 234 924 235
rect 982 239 988 240
rect 982 235 983 239
rect 987 235 988 239
rect 982 234 988 235
rect 1046 239 1052 240
rect 1046 235 1047 239
rect 1051 235 1052 239
rect 1046 234 1052 235
rect 1102 239 1108 240
rect 1102 235 1103 239
rect 1107 235 1108 239
rect 1102 234 1108 235
rect 1158 239 1164 240
rect 1158 235 1159 239
rect 1163 235 1164 239
rect 1158 234 1164 235
rect 510 221 516 222
rect 510 217 511 221
rect 515 217 516 221
rect 510 216 516 217
rect 590 221 596 222
rect 590 217 591 221
rect 595 217 596 221
rect 590 216 596 217
rect 678 221 684 222
rect 678 217 679 221
rect 683 217 684 221
rect 678 216 684 217
rect 512 207 514 216
rect 554 215 560 216
rect 554 211 555 215
rect 559 211 560 215
rect 554 210 560 211
rect 471 206 475 207
rect 471 201 475 202
rect 511 206 515 207
rect 511 201 515 202
rect 535 206 539 207
rect 535 201 539 202
rect 462 199 468 200
rect 414 195 420 196
rect 414 191 415 195
rect 419 191 420 195
rect 462 195 463 199
rect 467 195 468 199
rect 472 196 474 201
rect 536 196 538 201
rect 462 194 468 195
rect 470 195 476 196
rect 414 190 420 191
rect 470 191 471 195
rect 475 191 476 195
rect 470 190 476 191
rect 534 195 540 196
rect 534 191 535 195
rect 539 191 540 195
rect 534 190 540 191
rect 556 184 558 210
rect 592 207 594 216
rect 680 207 682 216
rect 591 206 595 207
rect 591 201 595 202
rect 607 206 611 207
rect 607 201 611 202
rect 679 206 683 207
rect 679 201 683 202
rect 751 206 755 207
rect 751 201 755 202
rect 608 196 610 201
rect 618 199 624 200
rect 606 195 612 196
rect 606 191 607 195
rect 611 191 612 195
rect 618 195 619 199
rect 623 195 624 199
rect 680 196 682 201
rect 752 196 754 201
rect 618 194 624 195
rect 678 195 684 196
rect 606 190 612 191
rect 374 183 380 184
rect 374 179 375 183
rect 379 179 380 183
rect 374 178 380 179
rect 554 183 560 184
rect 554 179 555 183
rect 559 179 560 183
rect 554 178 560 179
rect 358 177 364 178
rect 358 173 359 177
rect 363 173 364 177
rect 358 172 364 173
rect 414 177 420 178
rect 414 173 415 177
rect 419 173 420 177
rect 414 172 420 173
rect 470 177 476 178
rect 470 173 471 177
rect 475 173 476 177
rect 470 172 476 173
rect 534 177 540 178
rect 534 173 535 177
rect 539 173 540 177
rect 534 172 540 173
rect 606 177 612 178
rect 606 173 607 177
rect 611 173 612 177
rect 606 172 612 173
rect 351 170 355 171
rect 351 164 355 166
rect 359 170 363 172
rect 359 165 363 166
rect 407 170 411 171
rect 407 164 411 166
rect 415 170 419 172
rect 415 165 419 166
rect 463 170 467 171
rect 463 164 467 166
rect 471 170 475 172
rect 482 171 488 172
rect 482 167 483 171
rect 487 167 488 171
rect 482 166 488 167
rect 519 170 523 171
rect 471 165 475 166
rect 350 163 356 164
rect 350 159 351 163
rect 355 159 356 163
rect 350 158 356 159
rect 406 163 412 164
rect 406 159 407 163
rect 411 159 412 163
rect 406 158 412 159
rect 462 163 468 164
rect 462 159 463 163
rect 467 159 468 163
rect 462 158 468 159
rect 322 155 328 156
rect 322 151 323 155
rect 327 151 328 155
rect 322 150 328 151
rect 294 145 300 146
rect 294 141 295 145
rect 299 141 300 145
rect 294 140 300 141
rect 350 145 356 146
rect 350 141 351 145
rect 355 141 356 145
rect 350 140 356 141
rect 406 145 412 146
rect 406 141 407 145
rect 411 141 412 145
rect 406 140 412 141
rect 462 145 468 146
rect 462 141 463 145
rect 467 141 468 145
rect 462 140 468 141
rect 484 140 486 166
rect 519 164 523 166
rect 535 170 539 172
rect 535 165 539 166
rect 575 170 579 171
rect 575 164 579 166
rect 607 170 611 172
rect 607 165 611 166
rect 518 163 524 164
rect 518 159 519 163
rect 523 159 524 163
rect 518 158 524 159
rect 574 163 580 164
rect 574 159 575 163
rect 579 159 580 163
rect 574 158 580 159
rect 620 156 622 194
rect 678 191 679 195
rect 683 191 684 195
rect 678 190 684 191
rect 750 195 756 196
rect 750 191 751 195
rect 755 191 756 195
rect 750 190 756 191
rect 760 182 762 234
rect 1022 231 1028 232
rect 1022 227 1023 231
rect 1027 227 1028 231
rect 1022 226 1028 227
rect 1030 231 1036 232
rect 1030 227 1031 231
rect 1035 227 1036 231
rect 1030 226 1036 227
rect 766 221 772 222
rect 766 217 767 221
rect 771 217 772 221
rect 766 216 772 217
rect 846 221 852 222
rect 846 217 847 221
rect 851 217 852 221
rect 846 216 852 217
rect 918 221 924 222
rect 918 217 919 221
rect 923 217 924 221
rect 918 216 924 217
rect 982 221 988 222
rect 982 217 983 221
rect 987 217 988 221
rect 982 216 988 217
rect 768 207 770 216
rect 848 207 850 216
rect 920 207 922 216
rect 984 207 986 216
rect 767 206 771 207
rect 767 201 771 202
rect 815 206 819 207
rect 815 201 819 202
rect 847 206 851 207
rect 847 201 851 202
rect 879 206 883 207
rect 879 201 883 202
rect 919 206 923 207
rect 919 201 923 202
rect 943 206 947 207
rect 943 201 947 202
rect 983 206 987 207
rect 983 201 987 202
rect 1007 206 1011 207
rect 1007 201 1011 202
rect 816 196 818 201
rect 870 199 876 200
rect 814 195 820 196
rect 814 191 815 195
rect 819 191 820 195
rect 870 195 871 199
rect 875 195 876 199
rect 880 196 882 201
rect 944 196 946 201
rect 1008 196 1010 201
rect 1024 200 1026 226
rect 1032 208 1034 226
rect 1046 221 1052 222
rect 1046 217 1047 221
rect 1051 217 1052 221
rect 1046 216 1052 217
rect 1102 221 1108 222
rect 1102 217 1103 221
rect 1107 217 1108 221
rect 1102 216 1108 217
rect 1158 221 1164 222
rect 1158 217 1159 221
rect 1163 217 1164 221
rect 1158 216 1164 217
rect 1188 216 1190 254
rect 1222 253 1228 254
rect 1222 249 1223 253
rect 1227 249 1228 253
rect 1222 248 1228 249
rect 1262 253 1268 254
rect 1262 249 1263 253
rect 1267 249 1268 253
rect 1262 248 1268 249
rect 1302 253 1308 254
rect 1302 249 1303 253
rect 1307 249 1308 253
rect 1302 248 1308 249
rect 1350 253 1356 254
rect 1350 249 1351 253
rect 1355 249 1356 253
rect 1350 248 1356 249
rect 1215 246 1219 247
rect 1215 240 1219 242
rect 1223 246 1227 248
rect 1223 241 1227 242
rect 1263 246 1267 248
rect 1263 241 1267 242
rect 1271 246 1275 247
rect 1271 240 1275 242
rect 1303 246 1307 248
rect 1303 241 1307 242
rect 1327 246 1331 247
rect 1327 240 1331 242
rect 1351 246 1355 248
rect 1351 241 1355 242
rect 1214 239 1220 240
rect 1214 235 1215 239
rect 1219 235 1220 239
rect 1214 234 1220 235
rect 1270 239 1276 240
rect 1270 235 1271 239
rect 1275 235 1276 239
rect 1270 234 1276 235
rect 1326 239 1332 240
rect 1326 235 1327 239
rect 1331 235 1332 239
rect 1326 234 1332 235
rect 1246 231 1252 232
rect 1246 227 1247 231
rect 1251 227 1252 231
rect 1246 226 1252 227
rect 1214 221 1220 222
rect 1214 217 1215 221
rect 1219 217 1220 221
rect 1214 216 1220 217
rect 1030 207 1036 208
rect 1048 207 1050 216
rect 1104 207 1106 216
rect 1160 207 1162 216
rect 1186 215 1192 216
rect 1186 211 1187 215
rect 1191 211 1192 215
rect 1186 210 1192 211
rect 1216 207 1218 216
rect 1030 203 1031 207
rect 1035 203 1036 207
rect 1030 202 1036 203
rect 1047 206 1051 207
rect 1047 201 1051 202
rect 1063 206 1067 207
rect 1063 201 1067 202
rect 1103 206 1107 207
rect 1103 201 1107 202
rect 1119 206 1123 207
rect 1119 201 1123 202
rect 1159 206 1163 207
rect 1159 201 1163 202
rect 1175 206 1179 207
rect 1175 201 1179 202
rect 1215 206 1219 207
rect 1215 201 1219 202
rect 1231 206 1235 207
rect 1231 201 1235 202
rect 1022 199 1028 200
rect 870 194 876 195
rect 878 195 884 196
rect 814 190 820 191
rect 766 183 772 184
rect 766 182 767 183
rect 760 180 767 182
rect 766 179 767 180
rect 771 179 772 183
rect 766 178 772 179
rect 678 177 684 178
rect 678 173 679 177
rect 683 173 684 177
rect 678 172 684 173
rect 750 177 756 178
rect 750 173 751 177
rect 755 173 756 177
rect 750 172 756 173
rect 814 177 820 178
rect 814 173 815 177
rect 819 173 820 177
rect 814 172 820 173
rect 872 172 874 194
rect 878 191 879 195
rect 883 191 884 195
rect 878 190 884 191
rect 942 195 948 196
rect 942 191 943 195
rect 947 191 948 195
rect 942 190 948 191
rect 1006 195 1012 196
rect 1006 191 1007 195
rect 1011 191 1012 195
rect 1022 195 1023 199
rect 1027 195 1028 199
rect 1064 196 1066 201
rect 1120 196 1122 201
rect 1176 196 1178 201
rect 1232 196 1234 201
rect 1248 200 1250 226
rect 1270 221 1276 222
rect 1270 217 1271 221
rect 1275 217 1276 221
rect 1270 216 1276 217
rect 1326 221 1332 222
rect 1326 217 1327 221
rect 1331 217 1332 221
rect 1326 216 1332 217
rect 1364 216 1366 254
rect 1398 253 1404 254
rect 1398 249 1399 253
rect 1403 249 1404 253
rect 1398 248 1404 249
rect 1446 253 1452 254
rect 1446 249 1447 253
rect 1451 249 1452 253
rect 1446 248 1452 249
rect 1502 253 1508 254
rect 1502 249 1503 253
rect 1507 249 1508 253
rect 1502 248 1508 249
rect 1383 246 1387 247
rect 1383 240 1387 242
rect 1399 246 1403 248
rect 1399 241 1403 242
rect 1439 246 1443 247
rect 1439 240 1443 242
rect 1447 246 1451 248
rect 1447 241 1451 242
rect 1503 246 1507 248
rect 1503 240 1507 242
rect 1382 239 1388 240
rect 1382 235 1383 239
rect 1387 235 1388 239
rect 1382 234 1388 235
rect 1438 239 1444 240
rect 1438 235 1439 239
rect 1443 235 1444 239
rect 1438 234 1444 235
rect 1502 239 1508 240
rect 1502 235 1503 239
rect 1507 235 1508 239
rect 1502 234 1508 235
rect 1520 232 1522 270
rect 1542 267 1543 271
rect 1547 267 1548 271
rect 1558 271 1559 275
rect 1563 271 1564 275
rect 1584 273 1586 277
rect 1558 270 1564 271
rect 1582 272 1588 273
rect 1582 268 1583 272
rect 1587 268 1588 272
rect 1582 267 1588 268
rect 1542 266 1548 267
rect 1558 259 1564 260
rect 1558 255 1559 259
rect 1563 255 1564 259
rect 1558 254 1564 255
rect 1582 255 1588 256
rect 1542 253 1548 254
rect 1542 249 1543 253
rect 1547 249 1548 253
rect 1542 248 1548 249
rect 1543 246 1547 248
rect 1543 240 1547 242
rect 1542 239 1548 240
rect 1542 235 1543 239
rect 1547 235 1548 239
rect 1542 234 1548 235
rect 1518 231 1524 232
rect 1518 227 1519 231
rect 1523 227 1524 231
rect 1518 226 1524 227
rect 1382 221 1388 222
rect 1382 217 1383 221
rect 1387 217 1388 221
rect 1382 216 1388 217
rect 1438 221 1444 222
rect 1438 217 1439 221
rect 1443 217 1444 221
rect 1438 216 1444 217
rect 1502 221 1508 222
rect 1502 217 1503 221
rect 1507 217 1508 221
rect 1502 216 1508 217
rect 1542 221 1548 222
rect 1542 217 1543 221
rect 1547 217 1548 221
rect 1542 216 1548 217
rect 1560 216 1562 254
rect 1582 251 1583 255
rect 1587 251 1588 255
rect 1582 250 1588 251
rect 1584 247 1586 250
rect 1583 246 1587 247
rect 1583 241 1587 242
rect 1584 238 1586 241
rect 1582 237 1588 238
rect 1582 233 1583 237
rect 1587 233 1588 237
rect 1582 232 1588 233
rect 1582 220 1588 221
rect 1582 216 1583 220
rect 1587 216 1588 220
rect 1272 207 1274 216
rect 1302 207 1308 208
rect 1328 207 1330 216
rect 1362 215 1368 216
rect 1362 211 1363 215
rect 1367 211 1368 215
rect 1362 210 1368 211
rect 1384 207 1386 216
rect 1440 207 1442 216
rect 1470 207 1476 208
rect 1504 207 1506 216
rect 1544 207 1546 216
rect 1558 215 1564 216
rect 1582 215 1588 216
rect 1558 211 1559 215
rect 1563 211 1564 215
rect 1558 210 1564 211
rect 1584 207 1586 215
rect 1271 206 1275 207
rect 1271 201 1275 202
rect 1287 206 1291 207
rect 1302 203 1303 207
rect 1307 203 1308 207
rect 1302 202 1308 203
rect 1327 206 1331 207
rect 1287 201 1291 202
rect 1246 199 1252 200
rect 1022 194 1028 195
rect 1062 195 1068 196
rect 1006 190 1012 191
rect 1062 191 1063 195
rect 1067 191 1068 195
rect 1062 190 1068 191
rect 1118 195 1124 196
rect 1118 191 1119 195
rect 1123 191 1124 195
rect 1118 190 1124 191
rect 1174 195 1180 196
rect 1174 191 1175 195
rect 1179 191 1180 195
rect 1174 190 1180 191
rect 1230 195 1236 196
rect 1230 191 1231 195
rect 1235 191 1236 195
rect 1246 195 1247 199
rect 1251 195 1252 199
rect 1288 196 1290 201
rect 1246 194 1252 195
rect 1286 195 1292 196
rect 1230 190 1236 191
rect 1286 191 1287 195
rect 1291 191 1292 195
rect 1286 190 1292 191
rect 1304 184 1306 202
rect 1327 201 1331 202
rect 1343 206 1347 207
rect 1343 201 1347 202
rect 1383 206 1387 207
rect 1383 201 1387 202
rect 1399 206 1403 207
rect 1399 201 1403 202
rect 1439 206 1443 207
rect 1439 201 1443 202
rect 1455 206 1459 207
rect 1470 203 1471 207
rect 1475 203 1476 207
rect 1470 202 1476 203
rect 1503 206 1507 207
rect 1455 201 1459 202
rect 1344 196 1346 201
rect 1362 199 1368 200
rect 1342 195 1348 196
rect 1342 191 1343 195
rect 1347 191 1348 195
rect 1362 195 1363 199
rect 1367 195 1368 199
rect 1400 196 1402 201
rect 1456 196 1458 201
rect 1362 194 1368 195
rect 1398 195 1404 196
rect 1342 190 1348 191
rect 990 183 996 184
rect 990 179 991 183
rect 995 179 996 183
rect 990 178 996 179
rect 1186 183 1192 184
rect 1186 179 1187 183
rect 1191 179 1192 183
rect 1186 178 1192 179
rect 1302 183 1308 184
rect 1302 179 1303 183
rect 1307 179 1308 183
rect 1302 178 1308 179
rect 878 177 884 178
rect 878 173 879 177
rect 883 173 884 177
rect 878 172 884 173
rect 942 177 948 178
rect 942 173 943 177
rect 947 173 948 177
rect 942 172 948 173
rect 631 170 635 171
rect 631 164 635 166
rect 679 170 683 172
rect 679 165 683 166
rect 687 170 691 171
rect 687 164 691 166
rect 743 170 747 171
rect 743 164 747 166
rect 751 170 755 172
rect 751 165 755 166
rect 799 170 803 171
rect 799 164 803 166
rect 815 170 819 172
rect 870 171 876 172
rect 815 165 819 166
rect 855 170 859 171
rect 870 167 871 171
rect 875 167 876 171
rect 870 166 876 167
rect 879 170 883 172
rect 855 164 859 166
rect 879 165 883 166
rect 911 170 915 171
rect 911 164 915 166
rect 943 170 947 172
rect 943 165 947 166
rect 975 170 979 171
rect 975 164 979 166
rect 630 163 636 164
rect 630 159 631 163
rect 635 159 636 163
rect 630 158 636 159
rect 686 163 692 164
rect 686 159 687 163
rect 691 159 692 163
rect 686 158 692 159
rect 742 163 748 164
rect 742 159 743 163
rect 747 159 748 163
rect 742 158 748 159
rect 798 163 804 164
rect 798 159 799 163
rect 803 159 804 163
rect 798 158 804 159
rect 854 163 860 164
rect 854 159 855 163
rect 859 159 860 163
rect 854 158 860 159
rect 910 163 916 164
rect 910 159 911 163
rect 915 159 916 163
rect 910 158 916 159
rect 974 163 980 164
rect 974 159 975 163
rect 979 159 980 163
rect 974 158 980 159
rect 618 155 624 156
rect 618 151 619 155
rect 623 151 624 155
rect 618 150 624 151
rect 518 145 524 146
rect 518 141 519 145
rect 523 141 524 145
rect 518 140 524 141
rect 574 145 580 146
rect 574 141 575 145
rect 579 141 580 145
rect 574 140 580 141
rect 630 145 636 146
rect 630 141 631 145
rect 635 141 636 145
rect 630 140 636 141
rect 686 145 692 146
rect 686 141 687 145
rect 691 141 692 145
rect 686 140 692 141
rect 742 145 748 146
rect 742 141 743 145
rect 747 141 748 145
rect 742 140 748 141
rect 798 145 804 146
rect 798 141 799 145
rect 803 141 804 145
rect 798 140 804 141
rect 854 145 860 146
rect 854 141 855 145
rect 859 141 860 145
rect 854 140 860 141
rect 910 145 916 146
rect 910 141 911 145
rect 915 141 916 145
rect 910 140 916 141
rect 974 145 980 146
rect 974 141 975 145
rect 979 141 980 145
rect 974 140 980 141
rect 992 140 994 178
rect 1006 177 1012 178
rect 1006 173 1007 177
rect 1011 173 1012 177
rect 1006 172 1012 173
rect 1062 177 1068 178
rect 1062 173 1063 177
rect 1067 173 1068 177
rect 1062 172 1068 173
rect 1118 177 1124 178
rect 1118 173 1119 177
rect 1123 173 1124 177
rect 1118 172 1124 173
rect 1174 177 1180 178
rect 1174 173 1175 177
rect 1179 173 1180 177
rect 1174 172 1180 173
rect 1007 170 1011 172
rect 1007 165 1011 166
rect 1039 170 1043 171
rect 1039 164 1043 166
rect 1063 170 1067 172
rect 1063 165 1067 166
rect 1095 170 1099 171
rect 1095 164 1099 166
rect 1119 170 1123 172
rect 1119 165 1123 166
rect 1151 170 1155 171
rect 1151 164 1155 166
rect 1175 170 1179 172
rect 1175 165 1179 166
rect 1038 163 1044 164
rect 1038 159 1039 163
rect 1043 159 1044 163
rect 1038 158 1044 159
rect 1094 163 1100 164
rect 1094 159 1095 163
rect 1099 159 1100 163
rect 1094 158 1100 159
rect 1150 163 1156 164
rect 1150 159 1151 163
rect 1155 159 1156 163
rect 1150 158 1156 159
rect 1106 155 1112 156
rect 1106 151 1107 155
rect 1111 151 1112 155
rect 1106 150 1112 151
rect 1038 145 1044 146
rect 1038 141 1039 145
rect 1043 141 1044 145
rect 1038 140 1044 141
rect 1094 145 1100 146
rect 1094 141 1095 145
rect 1099 141 1100 145
rect 1094 140 1100 141
rect 192 123 194 140
rect 240 123 242 140
rect 274 139 280 140
rect 274 135 275 139
rect 279 135 280 139
rect 274 134 280 135
rect 296 123 298 140
rect 352 123 354 140
rect 408 123 410 140
rect 438 139 444 140
rect 438 135 439 139
rect 443 135 444 139
rect 438 134 444 135
rect 167 122 171 123
rect 167 117 171 118
rect 191 122 195 123
rect 191 117 195 118
rect 199 122 203 123
rect 199 117 203 118
rect 231 122 235 123
rect 231 117 235 118
rect 239 122 243 123
rect 239 117 243 118
rect 263 122 267 123
rect 263 117 267 118
rect 295 122 299 123
rect 295 117 299 118
rect 327 122 331 123
rect 327 117 331 118
rect 351 122 355 123
rect 351 117 355 118
rect 359 122 363 123
rect 359 117 363 118
rect 391 122 395 123
rect 391 117 395 118
rect 407 122 411 123
rect 407 117 411 118
rect 423 122 427 123
rect 423 117 427 118
rect 154 115 160 116
rect 110 108 111 112
rect 115 108 116 112
rect 110 107 116 108
rect 134 111 140 112
rect 134 107 135 111
rect 139 107 140 111
rect 154 111 155 115
rect 159 111 160 115
rect 168 112 170 117
rect 200 112 202 117
rect 232 112 234 117
rect 264 112 266 117
rect 296 112 298 117
rect 328 112 330 117
rect 360 112 362 117
rect 392 112 394 117
rect 424 112 426 117
rect 154 110 160 111
rect 166 111 172 112
rect 134 106 140 107
rect 166 107 167 111
rect 171 107 172 111
rect 166 106 172 107
rect 198 111 204 112
rect 198 107 199 111
rect 203 107 204 111
rect 198 106 204 107
rect 230 111 236 112
rect 230 107 231 111
rect 235 107 236 111
rect 230 106 236 107
rect 262 111 268 112
rect 262 107 263 111
rect 267 107 268 111
rect 262 106 268 107
rect 294 111 300 112
rect 294 107 295 111
rect 299 107 300 111
rect 294 106 300 107
rect 326 111 332 112
rect 326 107 327 111
rect 331 107 332 111
rect 326 106 332 107
rect 358 111 364 112
rect 358 107 359 111
rect 363 107 364 111
rect 358 106 364 107
rect 390 111 396 112
rect 390 107 391 111
rect 395 107 396 111
rect 390 106 396 107
rect 422 111 428 112
rect 422 107 423 111
rect 427 107 428 111
rect 422 106 428 107
rect 440 100 442 134
rect 464 123 466 140
rect 482 139 488 140
rect 482 135 483 139
rect 487 135 488 139
rect 482 134 488 135
rect 520 123 522 140
rect 538 131 544 132
rect 538 127 539 131
rect 543 127 544 131
rect 538 126 544 127
rect 455 122 459 123
rect 455 117 459 118
rect 463 122 467 123
rect 463 117 467 118
rect 487 122 491 123
rect 487 117 491 118
rect 519 122 523 123
rect 519 117 523 118
rect 456 112 458 117
rect 488 112 490 117
rect 520 112 522 117
rect 454 111 460 112
rect 454 107 455 111
rect 459 107 460 111
rect 454 106 460 107
rect 486 111 492 112
rect 486 107 487 111
rect 491 107 492 111
rect 486 106 492 107
rect 518 111 524 112
rect 518 107 519 111
rect 523 107 524 111
rect 518 106 524 107
rect 540 100 542 126
rect 562 123 568 124
rect 576 123 578 140
rect 632 123 634 140
rect 688 123 690 140
rect 744 123 746 140
rect 800 123 802 140
rect 856 123 858 140
rect 912 123 914 140
rect 976 123 978 140
rect 990 139 996 140
rect 990 135 991 139
rect 995 135 996 139
rect 990 134 996 135
rect 1040 123 1042 140
rect 1096 123 1098 140
rect 1108 132 1110 150
rect 1150 145 1156 146
rect 1150 141 1151 145
rect 1155 141 1156 145
rect 1150 140 1156 141
rect 1188 140 1190 178
rect 1230 177 1236 178
rect 1230 173 1231 177
rect 1235 173 1236 177
rect 1230 172 1236 173
rect 1286 177 1292 178
rect 1286 173 1287 177
rect 1291 173 1292 177
rect 1286 172 1292 173
rect 1342 177 1348 178
rect 1342 173 1343 177
rect 1347 173 1348 177
rect 1342 172 1348 173
rect 1207 170 1211 171
rect 1207 164 1211 166
rect 1231 170 1235 172
rect 1231 165 1235 166
rect 1255 170 1259 171
rect 1255 164 1259 166
rect 1287 170 1291 172
rect 1287 165 1291 166
rect 1303 170 1307 171
rect 1303 164 1307 166
rect 1343 170 1347 172
rect 1343 165 1347 166
rect 1351 170 1355 171
rect 1351 164 1355 166
rect 1206 163 1212 164
rect 1206 159 1207 163
rect 1211 159 1212 163
rect 1206 158 1212 159
rect 1254 163 1260 164
rect 1254 159 1255 163
rect 1259 159 1260 163
rect 1254 158 1260 159
rect 1302 163 1308 164
rect 1302 159 1303 163
rect 1307 159 1308 163
rect 1302 158 1308 159
rect 1350 163 1356 164
rect 1350 159 1351 163
rect 1355 159 1356 163
rect 1350 158 1356 159
rect 1364 156 1366 194
rect 1398 191 1399 195
rect 1403 191 1404 195
rect 1398 190 1404 191
rect 1454 195 1460 196
rect 1454 191 1455 195
rect 1459 191 1460 195
rect 1454 190 1460 191
rect 1472 184 1474 202
rect 1503 201 1507 202
rect 1511 206 1515 207
rect 1511 201 1515 202
rect 1543 206 1547 207
rect 1543 201 1547 202
rect 1583 206 1587 207
rect 1583 201 1587 202
rect 1512 196 1514 201
rect 1544 196 1546 201
rect 1584 197 1586 201
rect 1582 196 1588 197
rect 1510 195 1516 196
rect 1510 191 1511 195
rect 1515 191 1516 195
rect 1510 190 1516 191
rect 1542 195 1548 196
rect 1542 191 1543 195
rect 1547 191 1548 195
rect 1582 192 1583 196
rect 1587 192 1588 196
rect 1582 191 1588 192
rect 1542 190 1548 191
rect 1470 183 1476 184
rect 1470 179 1471 183
rect 1475 179 1476 183
rect 1470 178 1476 179
rect 1526 183 1532 184
rect 1526 179 1527 183
rect 1531 179 1532 183
rect 1526 178 1532 179
rect 1582 179 1588 180
rect 1398 177 1404 178
rect 1398 173 1399 177
rect 1403 173 1404 177
rect 1398 172 1404 173
rect 1454 177 1460 178
rect 1454 173 1455 177
rect 1459 173 1460 177
rect 1454 172 1460 173
rect 1510 177 1516 178
rect 1510 173 1511 177
rect 1515 173 1516 177
rect 1510 172 1516 173
rect 1399 170 1403 172
rect 1399 164 1403 166
rect 1455 170 1459 172
rect 1455 164 1459 166
rect 1511 170 1515 172
rect 1511 164 1515 166
rect 1398 163 1404 164
rect 1398 159 1399 163
rect 1403 159 1404 163
rect 1398 158 1404 159
rect 1454 163 1460 164
rect 1454 159 1455 163
rect 1459 159 1460 163
rect 1454 158 1460 159
rect 1510 163 1516 164
rect 1510 159 1511 163
rect 1515 159 1516 163
rect 1510 158 1516 159
rect 1314 155 1320 156
rect 1314 151 1315 155
rect 1319 151 1320 155
rect 1314 150 1320 151
rect 1362 155 1368 156
rect 1362 151 1363 155
rect 1367 151 1368 155
rect 1362 150 1368 151
rect 1206 145 1212 146
rect 1206 141 1207 145
rect 1211 141 1212 145
rect 1206 140 1212 141
rect 1254 145 1260 146
rect 1254 141 1255 145
rect 1259 141 1260 145
rect 1254 140 1260 141
rect 1302 145 1308 146
rect 1302 141 1303 145
rect 1307 141 1308 145
rect 1302 140 1308 141
rect 1106 131 1112 132
rect 1106 127 1107 131
rect 1111 127 1112 131
rect 1106 126 1112 127
rect 1152 123 1154 140
rect 1186 139 1192 140
rect 1186 135 1187 139
rect 1191 135 1192 139
rect 1186 134 1192 135
rect 1208 123 1210 140
rect 1256 123 1258 140
rect 1304 123 1306 140
rect 1316 124 1318 150
rect 1350 145 1356 146
rect 1350 141 1351 145
rect 1355 141 1356 145
rect 1350 140 1356 141
rect 1398 145 1404 146
rect 1398 141 1399 145
rect 1403 141 1404 145
rect 1398 140 1404 141
rect 1454 145 1460 146
rect 1454 141 1455 145
rect 1459 141 1460 145
rect 1454 140 1460 141
rect 1510 145 1516 146
rect 1510 141 1511 145
rect 1515 141 1516 145
rect 1510 140 1516 141
rect 1528 140 1530 178
rect 1542 177 1548 178
rect 1542 173 1543 177
rect 1547 173 1548 177
rect 1582 175 1583 179
rect 1587 175 1588 179
rect 1582 174 1588 175
rect 1542 172 1548 173
rect 1543 170 1547 172
rect 1584 171 1586 174
rect 1543 164 1547 166
rect 1583 170 1587 171
rect 1583 165 1587 166
rect 1542 163 1548 164
rect 1542 159 1543 163
rect 1547 159 1548 163
rect 1584 162 1586 165
rect 1542 158 1548 159
rect 1582 161 1588 162
rect 1582 157 1583 161
rect 1587 157 1588 161
rect 1582 156 1588 157
rect 1558 155 1564 156
rect 1558 151 1559 155
rect 1563 151 1564 155
rect 1558 150 1564 151
rect 1542 145 1548 146
rect 1542 141 1543 145
rect 1547 141 1548 145
rect 1542 140 1548 141
rect 1314 123 1320 124
rect 1352 123 1354 140
rect 1400 123 1402 140
rect 1456 123 1458 140
rect 1486 139 1492 140
rect 1486 135 1487 139
rect 1491 135 1492 139
rect 1486 134 1492 135
rect 551 122 555 123
rect 562 119 563 123
rect 567 119 568 123
rect 562 118 568 119
rect 575 122 579 123
rect 551 117 555 118
rect 552 112 554 117
rect 550 111 556 112
rect 550 107 551 111
rect 555 107 556 111
rect 550 106 556 107
rect 564 100 566 118
rect 575 117 579 118
rect 583 122 587 123
rect 583 117 587 118
rect 615 122 619 123
rect 615 117 619 118
rect 631 122 635 123
rect 631 117 635 118
rect 647 122 651 123
rect 647 117 651 118
rect 679 122 683 123
rect 679 117 683 118
rect 687 122 691 123
rect 687 117 691 118
rect 711 122 715 123
rect 711 117 715 118
rect 743 122 747 123
rect 743 117 747 118
rect 775 122 779 123
rect 775 117 779 118
rect 799 122 803 123
rect 799 117 803 118
rect 807 122 811 123
rect 807 117 811 118
rect 839 122 843 123
rect 839 117 843 118
rect 855 122 859 123
rect 855 117 859 118
rect 871 122 875 123
rect 871 117 875 118
rect 903 122 907 123
rect 903 117 907 118
rect 911 122 915 123
rect 911 117 915 118
rect 943 122 947 123
rect 943 117 947 118
rect 975 122 979 123
rect 975 117 979 118
rect 983 122 987 123
rect 983 117 987 118
rect 1031 122 1035 123
rect 1031 117 1035 118
rect 1039 122 1043 123
rect 1039 117 1043 118
rect 1079 122 1083 123
rect 1079 117 1083 118
rect 1095 122 1099 123
rect 1095 117 1099 118
rect 1127 122 1131 123
rect 1127 117 1131 118
rect 1151 122 1155 123
rect 1151 117 1155 118
rect 1175 122 1179 123
rect 1175 117 1179 118
rect 1207 122 1211 123
rect 1207 117 1211 118
rect 1223 122 1227 123
rect 1223 117 1227 118
rect 1255 122 1259 123
rect 1255 117 1259 118
rect 1263 122 1267 123
rect 1263 117 1267 118
rect 1303 122 1307 123
rect 1314 119 1315 123
rect 1319 119 1320 123
rect 1314 118 1320 119
rect 1343 122 1347 123
rect 1303 117 1307 118
rect 1343 117 1347 118
rect 1351 122 1355 123
rect 1351 117 1355 118
rect 1383 122 1387 123
rect 1383 117 1387 118
rect 1399 122 1403 123
rect 1399 117 1403 118
rect 1423 122 1427 123
rect 1423 117 1427 118
rect 1455 122 1459 123
rect 1455 117 1459 118
rect 1471 122 1475 123
rect 1471 117 1475 118
rect 584 112 586 117
rect 616 112 618 117
rect 648 112 650 117
rect 680 112 682 117
rect 712 112 714 117
rect 744 112 746 117
rect 776 112 778 117
rect 808 112 810 117
rect 840 112 842 117
rect 872 112 874 117
rect 904 112 906 117
rect 944 112 946 117
rect 984 112 986 117
rect 1022 115 1028 116
rect 582 111 588 112
rect 582 107 583 111
rect 587 107 588 111
rect 582 106 588 107
rect 614 111 620 112
rect 614 107 615 111
rect 619 107 620 111
rect 614 106 620 107
rect 646 111 652 112
rect 646 107 647 111
rect 651 107 652 111
rect 646 106 652 107
rect 678 111 684 112
rect 678 107 679 111
rect 683 107 684 111
rect 678 106 684 107
rect 710 111 716 112
rect 710 107 711 111
rect 715 107 716 111
rect 710 106 716 107
rect 742 111 748 112
rect 742 107 743 111
rect 747 107 748 111
rect 742 106 748 107
rect 774 111 780 112
rect 774 107 775 111
rect 779 107 780 111
rect 774 106 780 107
rect 806 111 812 112
rect 806 107 807 111
rect 811 107 812 111
rect 806 106 812 107
rect 838 111 844 112
rect 838 107 839 111
rect 843 107 844 111
rect 838 106 844 107
rect 870 111 876 112
rect 870 107 871 111
rect 875 107 876 111
rect 870 106 876 107
rect 902 111 908 112
rect 902 107 903 111
rect 907 107 908 111
rect 902 106 908 107
rect 942 111 948 112
rect 942 107 943 111
rect 947 107 948 111
rect 942 106 948 107
rect 982 111 988 112
rect 982 107 983 111
rect 987 107 988 111
rect 1022 111 1023 115
rect 1027 111 1028 115
rect 1032 112 1034 117
rect 1080 112 1082 117
rect 1128 112 1130 117
rect 1176 112 1178 117
rect 1224 112 1226 117
rect 1264 112 1266 117
rect 1304 112 1306 117
rect 1344 112 1346 117
rect 1384 112 1386 117
rect 1424 112 1426 117
rect 1472 112 1474 117
rect 1022 110 1028 111
rect 1030 111 1036 112
rect 982 106 988 107
rect 438 99 444 100
rect 110 95 116 96
rect 110 91 111 95
rect 115 91 116 95
rect 438 95 439 99
rect 443 95 444 99
rect 438 94 444 95
rect 538 99 544 100
rect 538 95 539 99
rect 543 95 544 99
rect 538 94 544 95
rect 562 99 568 100
rect 562 95 563 99
rect 567 95 568 99
rect 562 94 568 95
rect 110 90 116 91
rect 134 93 140 94
rect 112 87 114 90
rect 134 89 135 93
rect 139 89 140 93
rect 134 88 140 89
rect 166 93 172 94
rect 166 89 167 93
rect 171 89 172 93
rect 166 88 172 89
rect 198 93 204 94
rect 198 89 199 93
rect 203 89 204 93
rect 198 88 204 89
rect 230 93 236 94
rect 230 89 231 93
rect 235 89 236 93
rect 230 88 236 89
rect 262 93 268 94
rect 262 89 263 93
rect 267 89 268 93
rect 262 88 268 89
rect 294 93 300 94
rect 294 89 295 93
rect 299 89 300 93
rect 294 88 300 89
rect 326 93 332 94
rect 326 89 327 93
rect 331 89 332 93
rect 326 88 332 89
rect 358 93 364 94
rect 358 89 359 93
rect 363 89 364 93
rect 358 88 364 89
rect 390 93 396 94
rect 390 89 391 93
rect 395 89 396 93
rect 390 88 396 89
rect 422 93 428 94
rect 422 89 423 93
rect 427 89 428 93
rect 422 88 428 89
rect 454 93 460 94
rect 454 89 455 93
rect 459 89 460 93
rect 454 88 460 89
rect 486 93 492 94
rect 486 89 487 93
rect 491 89 492 93
rect 486 88 492 89
rect 518 93 524 94
rect 518 89 519 93
rect 523 89 524 93
rect 518 88 524 89
rect 550 93 556 94
rect 550 89 551 93
rect 555 89 556 93
rect 550 88 556 89
rect 582 93 588 94
rect 582 89 583 93
rect 587 89 588 93
rect 582 88 588 89
rect 614 93 620 94
rect 614 89 615 93
rect 619 89 620 93
rect 614 88 620 89
rect 646 93 652 94
rect 646 89 647 93
rect 651 89 652 93
rect 646 88 652 89
rect 678 93 684 94
rect 678 89 679 93
rect 683 89 684 93
rect 678 88 684 89
rect 710 93 716 94
rect 710 89 711 93
rect 715 89 716 93
rect 710 88 716 89
rect 742 93 748 94
rect 742 89 743 93
rect 747 89 748 93
rect 742 88 748 89
rect 774 93 780 94
rect 774 89 775 93
rect 779 89 780 93
rect 774 88 780 89
rect 806 93 812 94
rect 806 89 807 93
rect 811 89 812 93
rect 806 88 812 89
rect 838 93 844 94
rect 838 89 839 93
rect 843 89 844 93
rect 838 88 844 89
rect 870 93 876 94
rect 870 89 871 93
rect 875 89 876 93
rect 870 88 876 89
rect 902 93 908 94
rect 902 89 903 93
rect 907 89 908 93
rect 902 88 908 89
rect 942 93 948 94
rect 942 89 943 93
rect 947 89 948 93
rect 942 88 948 89
rect 982 93 988 94
rect 982 89 983 93
rect 987 89 988 93
rect 982 88 988 89
rect 1024 88 1026 110
rect 1030 107 1031 111
rect 1035 107 1036 111
rect 1030 106 1036 107
rect 1078 111 1084 112
rect 1078 107 1079 111
rect 1083 107 1084 111
rect 1078 106 1084 107
rect 1126 111 1132 112
rect 1126 107 1127 111
rect 1131 107 1132 111
rect 1126 106 1132 107
rect 1174 111 1180 112
rect 1174 107 1175 111
rect 1179 107 1180 111
rect 1174 106 1180 107
rect 1222 111 1228 112
rect 1222 107 1223 111
rect 1227 107 1228 111
rect 1222 106 1228 107
rect 1262 111 1268 112
rect 1262 107 1263 111
rect 1267 107 1268 111
rect 1262 106 1268 107
rect 1302 111 1308 112
rect 1302 107 1303 111
rect 1307 107 1308 111
rect 1302 106 1308 107
rect 1342 111 1348 112
rect 1342 107 1343 111
rect 1347 107 1348 111
rect 1342 106 1348 107
rect 1382 111 1388 112
rect 1382 107 1383 111
rect 1387 107 1388 111
rect 1382 106 1388 107
rect 1422 111 1428 112
rect 1422 107 1423 111
rect 1427 107 1428 111
rect 1422 106 1428 107
rect 1470 111 1476 112
rect 1470 107 1471 111
rect 1475 107 1476 111
rect 1470 106 1476 107
rect 1488 100 1490 134
rect 1512 123 1514 140
rect 1526 139 1532 140
rect 1526 135 1527 139
rect 1531 135 1532 139
rect 1526 134 1532 135
rect 1544 123 1546 140
rect 1511 122 1515 123
rect 1511 117 1515 118
rect 1543 122 1547 123
rect 1543 117 1547 118
rect 1512 112 1514 117
rect 1544 112 1546 117
rect 1560 116 1562 150
rect 1582 144 1588 145
rect 1582 140 1583 144
rect 1587 140 1588 144
rect 1582 139 1588 140
rect 1584 123 1586 139
rect 1583 122 1587 123
rect 1583 117 1587 118
rect 1558 115 1564 116
rect 1510 111 1516 112
rect 1510 107 1511 111
rect 1515 107 1516 111
rect 1510 106 1516 107
rect 1542 111 1548 112
rect 1542 107 1543 111
rect 1547 107 1548 111
rect 1558 111 1559 115
rect 1563 111 1564 115
rect 1584 113 1586 117
rect 1558 110 1564 111
rect 1582 112 1588 113
rect 1582 108 1583 112
rect 1587 108 1588 112
rect 1582 107 1588 108
rect 1542 106 1548 107
rect 1486 99 1492 100
rect 1486 95 1487 99
rect 1491 95 1492 99
rect 1486 94 1492 95
rect 1582 95 1588 96
rect 1030 93 1036 94
rect 1030 89 1031 93
rect 1035 89 1036 93
rect 1030 88 1036 89
rect 1078 93 1084 94
rect 1078 89 1079 93
rect 1083 89 1084 93
rect 1078 88 1084 89
rect 1126 93 1132 94
rect 1126 89 1127 93
rect 1131 89 1132 93
rect 1126 88 1132 89
rect 1174 93 1180 94
rect 1174 89 1175 93
rect 1179 89 1180 93
rect 1174 88 1180 89
rect 1222 93 1228 94
rect 1222 89 1223 93
rect 1227 89 1228 93
rect 1222 88 1228 89
rect 1262 93 1268 94
rect 1262 89 1263 93
rect 1267 89 1268 93
rect 1262 88 1268 89
rect 1302 93 1308 94
rect 1302 89 1303 93
rect 1307 89 1308 93
rect 1302 88 1308 89
rect 1342 93 1348 94
rect 1342 89 1343 93
rect 1347 89 1348 93
rect 1342 88 1348 89
rect 1382 93 1388 94
rect 1382 89 1383 93
rect 1387 89 1388 93
rect 1382 88 1388 89
rect 1422 93 1428 94
rect 1422 89 1423 93
rect 1427 89 1428 93
rect 1422 88 1428 89
rect 1470 93 1476 94
rect 1470 89 1471 93
rect 1475 89 1476 93
rect 1470 88 1476 89
rect 1510 93 1516 94
rect 1510 89 1511 93
rect 1515 89 1516 93
rect 1510 88 1516 89
rect 1542 93 1548 94
rect 1542 89 1543 93
rect 1547 89 1548 93
rect 1582 91 1583 95
rect 1587 91 1588 95
rect 1582 90 1588 91
rect 1542 88 1548 89
rect 111 86 115 87
rect 111 81 115 82
rect 135 86 139 88
rect 135 81 139 82
rect 167 86 171 88
rect 167 81 171 82
rect 199 86 203 88
rect 199 81 203 82
rect 231 86 235 88
rect 231 81 235 82
rect 263 86 267 88
rect 263 81 267 82
rect 295 86 299 88
rect 295 81 299 82
rect 327 86 331 88
rect 327 81 331 82
rect 359 86 363 88
rect 359 81 363 82
rect 391 86 395 88
rect 391 81 395 82
rect 423 86 427 88
rect 423 81 427 82
rect 455 86 459 88
rect 455 81 459 82
rect 487 86 491 88
rect 487 81 491 82
rect 519 86 523 88
rect 519 81 523 82
rect 551 86 555 88
rect 551 81 555 82
rect 583 86 587 88
rect 583 81 587 82
rect 615 86 619 88
rect 615 81 619 82
rect 647 86 651 88
rect 647 81 651 82
rect 679 86 683 88
rect 679 81 683 82
rect 711 86 715 88
rect 711 81 715 82
rect 743 86 747 88
rect 743 81 747 82
rect 775 86 779 88
rect 775 81 779 82
rect 807 86 811 88
rect 807 81 811 82
rect 839 86 843 88
rect 839 81 843 82
rect 871 86 875 88
rect 871 81 875 82
rect 903 86 907 88
rect 903 81 907 82
rect 943 86 947 88
rect 943 81 947 82
rect 983 86 987 88
rect 1022 87 1028 88
rect 1022 83 1023 87
rect 1027 83 1028 87
rect 1022 82 1028 83
rect 1031 86 1035 88
rect 983 81 987 82
rect 1031 81 1035 82
rect 1079 86 1083 88
rect 1079 81 1083 82
rect 1127 86 1131 88
rect 1127 81 1131 82
rect 1175 86 1179 88
rect 1175 81 1179 82
rect 1223 86 1227 88
rect 1223 81 1227 82
rect 1263 86 1267 88
rect 1263 81 1267 82
rect 1303 86 1307 88
rect 1303 81 1307 82
rect 1343 86 1347 88
rect 1343 81 1347 82
rect 1383 86 1387 88
rect 1383 81 1387 82
rect 1423 86 1427 88
rect 1423 81 1427 82
rect 1471 86 1475 88
rect 1471 81 1475 82
rect 1511 86 1515 88
rect 1511 81 1515 82
rect 1543 86 1547 88
rect 1584 87 1586 90
rect 1543 81 1547 82
rect 1583 86 1587 87
rect 1583 81 1587 82
<< m4c >>
rect 111 1650 115 1654
rect 135 1650 139 1654
rect 167 1650 171 1654
rect 199 1650 203 1654
rect 1583 1650 1587 1654
rect 111 1614 115 1618
rect 135 1614 139 1618
rect 167 1614 171 1618
rect 175 1614 179 1618
rect 199 1614 203 1618
rect 239 1614 243 1618
rect 295 1614 299 1618
rect 351 1614 355 1618
rect 407 1614 411 1618
rect 455 1614 459 1618
rect 503 1614 507 1618
rect 551 1614 555 1618
rect 599 1614 603 1618
rect 647 1614 651 1618
rect 695 1614 699 1618
rect 743 1614 747 1618
rect 791 1614 795 1618
rect 839 1614 843 1618
rect 887 1614 891 1618
rect 935 1614 939 1618
rect 991 1614 995 1618
rect 1047 1614 1051 1618
rect 1095 1614 1099 1618
rect 1143 1614 1147 1618
rect 1191 1614 1195 1618
rect 1239 1614 1243 1618
rect 1287 1614 1291 1618
rect 1327 1614 1331 1618
rect 1367 1614 1371 1618
rect 1407 1614 1411 1618
rect 1447 1614 1451 1618
rect 1479 1614 1483 1618
rect 1511 1614 1515 1618
rect 1543 1614 1547 1618
rect 1583 1614 1587 1618
rect 111 1578 115 1582
rect 135 1578 139 1582
rect 175 1578 179 1582
rect 215 1578 219 1582
rect 239 1578 243 1582
rect 255 1578 259 1582
rect 295 1578 299 1582
rect 343 1578 347 1582
rect 351 1578 355 1582
rect 391 1578 395 1582
rect 407 1578 411 1582
rect 439 1578 443 1582
rect 455 1578 459 1582
rect 487 1578 491 1582
rect 503 1578 507 1582
rect 535 1578 539 1582
rect 551 1578 555 1582
rect 583 1578 587 1582
rect 599 1578 603 1582
rect 639 1578 643 1582
rect 647 1578 651 1582
rect 695 1578 699 1582
rect 703 1578 707 1582
rect 743 1578 747 1582
rect 775 1578 779 1582
rect 791 1578 795 1582
rect 839 1578 843 1582
rect 855 1578 859 1582
rect 887 1578 891 1582
rect 935 1578 939 1582
rect 991 1578 995 1582
rect 1015 1578 1019 1582
rect 1047 1578 1051 1582
rect 1087 1578 1091 1582
rect 1095 1578 1099 1582
rect 1143 1578 1147 1582
rect 111 1542 115 1546
rect 159 1542 163 1546
rect 175 1542 179 1546
rect 207 1542 211 1546
rect 215 1542 219 1546
rect 255 1542 259 1546
rect 295 1542 299 1546
rect 311 1542 315 1546
rect 343 1542 347 1546
rect 359 1542 363 1546
rect 391 1542 395 1546
rect 415 1542 419 1546
rect 439 1542 443 1546
rect 471 1542 475 1546
rect 487 1542 491 1546
rect 527 1542 531 1546
rect 535 1542 539 1546
rect 583 1542 587 1546
rect 639 1542 643 1546
rect 695 1542 699 1546
rect 703 1542 707 1546
rect 759 1542 763 1546
rect 775 1542 779 1546
rect 823 1542 827 1546
rect 855 1542 859 1546
rect 895 1542 899 1546
rect 111 1506 115 1510
rect 159 1506 163 1510
rect 207 1506 211 1510
rect 255 1506 259 1510
rect 303 1506 307 1510
rect 311 1506 315 1510
rect 351 1506 355 1510
rect 359 1506 363 1510
rect 407 1506 411 1510
rect 415 1506 419 1510
rect 463 1506 467 1510
rect 471 1506 475 1510
rect 527 1506 531 1510
rect 111 1470 115 1474
rect 135 1470 139 1474
rect 159 1470 163 1474
rect 183 1470 187 1474
rect 207 1470 211 1474
rect 231 1470 235 1474
rect 255 1470 259 1474
rect 259 1459 263 1460
rect 259 1456 263 1459
rect 111 1434 115 1438
rect 135 1434 139 1438
rect 287 1470 291 1474
rect 303 1470 307 1474
rect 343 1470 347 1474
rect 351 1470 355 1474
rect 399 1470 403 1474
rect 407 1470 411 1474
rect 455 1470 459 1474
rect 463 1470 467 1474
rect 583 1506 587 1510
rect 591 1506 595 1510
rect 639 1506 643 1510
rect 655 1506 659 1510
rect 695 1506 699 1510
rect 719 1506 723 1510
rect 759 1506 763 1510
rect 935 1542 939 1546
rect 967 1542 971 1546
rect 1159 1578 1163 1582
rect 1191 1578 1195 1582
rect 1239 1578 1243 1582
rect 1287 1578 1291 1582
rect 1319 1578 1323 1582
rect 1327 1578 1331 1582
rect 1367 1578 1371 1582
rect 1399 1578 1403 1582
rect 1407 1578 1411 1582
rect 1447 1578 1451 1582
rect 1479 1578 1483 1582
rect 1511 1578 1515 1582
rect 1543 1578 1547 1582
rect 1583 1578 1587 1582
rect 1015 1542 1019 1546
rect 1039 1542 1043 1546
rect 1087 1542 1091 1546
rect 1103 1542 1107 1546
rect 1159 1542 1163 1546
rect 1167 1542 1171 1546
rect 1231 1542 1235 1546
rect 1239 1542 1243 1546
rect 1295 1542 1299 1546
rect 1319 1542 1323 1546
rect 783 1506 787 1510
rect 823 1506 827 1510
rect 855 1506 859 1510
rect 895 1506 899 1510
rect 935 1506 939 1510
rect 967 1506 971 1510
rect 1007 1506 1011 1510
rect 1039 1506 1043 1510
rect 1079 1506 1083 1510
rect 1103 1506 1107 1510
rect 511 1470 515 1474
rect 527 1470 531 1474
rect 575 1470 579 1474
rect 591 1470 595 1474
rect 631 1470 635 1474
rect 655 1470 659 1474
rect 687 1470 691 1474
rect 719 1470 723 1474
rect 751 1470 755 1474
rect 783 1470 787 1474
rect 815 1470 819 1474
rect 415 1456 419 1460
rect 183 1434 187 1438
rect 231 1434 235 1438
rect 255 1434 259 1438
rect 287 1434 291 1438
rect 327 1434 331 1438
rect 343 1434 347 1438
rect 399 1434 403 1438
rect 455 1434 459 1438
rect 471 1434 475 1438
rect 511 1434 515 1438
rect 543 1434 547 1438
rect 575 1434 579 1438
rect 615 1434 619 1438
rect 631 1434 635 1438
rect 111 1398 115 1402
rect 135 1398 139 1402
rect 175 1398 179 1402
rect 183 1398 187 1402
rect 247 1398 251 1402
rect 255 1398 259 1402
rect 319 1398 323 1402
rect 327 1398 331 1402
rect 391 1398 395 1402
rect 399 1398 403 1402
rect 455 1398 459 1402
rect 471 1398 475 1402
rect 679 1434 683 1438
rect 687 1434 691 1438
rect 855 1470 859 1474
rect 879 1470 883 1474
rect 1359 1542 1363 1546
rect 1399 1542 1403 1546
rect 1423 1542 1427 1546
rect 1479 1542 1483 1546
rect 1495 1542 1499 1546
rect 1543 1542 1547 1546
rect 1583 1542 1587 1546
rect 1151 1506 1155 1510
rect 1167 1506 1171 1510
rect 1215 1506 1219 1510
rect 1231 1506 1235 1510
rect 1279 1506 1283 1510
rect 1295 1506 1299 1510
rect 1351 1506 1355 1510
rect 1359 1506 1363 1510
rect 1423 1506 1427 1510
rect 1495 1506 1499 1510
rect 1543 1506 1547 1510
rect 1583 1506 1587 1510
rect 935 1470 939 1474
rect 943 1470 947 1474
rect 1007 1470 1011 1474
rect 1015 1470 1019 1474
rect 1079 1470 1083 1474
rect 1087 1470 1091 1474
rect 1151 1470 1155 1474
rect 1159 1470 1163 1474
rect 1215 1470 1219 1474
rect 1239 1470 1243 1474
rect 1279 1470 1283 1474
rect 1319 1470 1323 1474
rect 1351 1470 1355 1474
rect 1399 1470 1403 1474
rect 1423 1470 1427 1474
rect 1479 1470 1483 1474
rect 1495 1470 1499 1474
rect 1543 1470 1547 1474
rect 1583 1470 1587 1474
rect 743 1434 747 1438
rect 751 1434 755 1438
rect 815 1434 819 1438
rect 879 1434 883 1438
rect 943 1434 947 1438
rect 519 1398 523 1402
rect 543 1398 547 1402
rect 583 1398 587 1402
rect 615 1398 619 1402
rect 647 1398 651 1402
rect 679 1398 683 1402
rect 711 1398 715 1402
rect 743 1398 747 1402
rect 775 1398 779 1402
rect 815 1398 819 1402
rect 839 1398 843 1402
rect 111 1362 115 1366
rect 135 1362 139 1366
rect 879 1398 883 1402
rect 895 1398 899 1402
rect 951 1434 955 1438
rect 1015 1434 1019 1438
rect 1023 1434 1027 1438
rect 1087 1434 1091 1438
rect 1095 1434 1099 1438
rect 951 1398 955 1402
rect 999 1398 1003 1402
rect 1023 1398 1027 1402
rect 1055 1398 1059 1402
rect 1095 1398 1099 1402
rect 1159 1434 1163 1438
rect 1223 1434 1227 1438
rect 1239 1434 1243 1438
rect 1287 1434 1291 1438
rect 1319 1434 1323 1438
rect 1343 1434 1347 1438
rect 1399 1434 1403 1438
rect 1455 1434 1459 1438
rect 1479 1434 1483 1438
rect 1511 1434 1515 1438
rect 1111 1398 1115 1402
rect 1159 1398 1163 1402
rect 1175 1398 1179 1402
rect 1223 1398 1227 1402
rect 1239 1398 1243 1402
rect 1287 1398 1291 1402
rect 1295 1398 1299 1402
rect 167 1362 171 1366
rect 175 1362 179 1366
rect 215 1362 219 1366
rect 247 1362 251 1366
rect 303 1362 307 1366
rect 319 1362 323 1366
rect 391 1362 395 1366
rect 415 1362 419 1366
rect 455 1362 459 1366
rect 519 1362 523 1366
rect 527 1362 531 1366
rect 583 1362 587 1366
rect 639 1362 643 1366
rect 647 1362 651 1366
rect 711 1362 715 1366
rect 751 1362 755 1366
rect 775 1362 779 1366
rect 839 1362 843 1366
rect 863 1362 867 1366
rect 895 1362 899 1366
rect 951 1362 955 1366
rect 967 1362 971 1366
rect 999 1362 1003 1366
rect 1055 1362 1059 1366
rect 1063 1362 1067 1366
rect 1111 1362 1115 1366
rect 1151 1362 1155 1366
rect 1175 1362 1179 1366
rect 1343 1398 1347 1402
rect 1351 1398 1355 1402
rect 1399 1398 1403 1402
rect 1415 1398 1419 1402
rect 1455 1398 1459 1402
rect 1479 1398 1483 1402
rect 1543 1434 1547 1438
rect 1583 1434 1587 1438
rect 1511 1398 1515 1402
rect 1543 1398 1547 1402
rect 1583 1398 1587 1402
rect 1231 1362 1235 1366
rect 1239 1362 1243 1366
rect 1295 1362 1299 1366
rect 1311 1362 1315 1366
rect 1351 1362 1355 1366
rect 1383 1362 1387 1366
rect 1415 1362 1419 1366
rect 1455 1362 1459 1366
rect 111 1326 115 1330
rect 135 1326 139 1330
rect 167 1326 171 1330
rect 183 1326 187 1330
rect 215 1326 219 1330
rect 247 1326 251 1330
rect 303 1326 307 1330
rect 311 1326 315 1330
rect 375 1326 379 1330
rect 415 1326 419 1330
rect 439 1326 443 1330
rect 495 1326 499 1330
rect 527 1326 531 1330
rect 543 1326 547 1330
rect 591 1326 595 1330
rect 639 1326 643 1330
rect 687 1326 691 1330
rect 743 1326 747 1330
rect 751 1326 755 1330
rect 791 1326 795 1330
rect 839 1326 843 1330
rect 863 1326 867 1330
rect 887 1326 891 1330
rect 111 1290 115 1294
rect 135 1290 139 1294
rect 183 1290 187 1294
rect 191 1290 195 1294
rect 247 1290 251 1294
rect 255 1290 259 1294
rect 311 1290 315 1294
rect 327 1290 331 1294
rect 375 1290 379 1294
rect 391 1290 395 1294
rect 1355 1339 1359 1340
rect 1355 1336 1359 1339
rect 935 1326 939 1330
rect 967 1326 971 1330
rect 991 1326 995 1330
rect 1047 1326 1051 1330
rect 439 1290 443 1294
rect 463 1290 467 1294
rect 1063 1326 1067 1330
rect 1103 1326 1107 1330
rect 1151 1326 1155 1330
rect 1159 1326 1163 1330
rect 1215 1326 1219 1330
rect 1231 1326 1235 1330
rect 495 1290 499 1294
rect 535 1290 539 1294
rect 543 1290 547 1294
rect 591 1290 595 1294
rect 599 1290 603 1294
rect 639 1290 643 1294
rect 663 1290 667 1294
rect 687 1290 691 1294
rect 727 1290 731 1294
rect 743 1290 747 1294
rect 791 1290 795 1294
rect 839 1290 843 1294
rect 111 1254 115 1258
rect 135 1254 139 1258
rect 175 1254 179 1258
rect 191 1254 195 1258
rect 231 1254 235 1258
rect 255 1254 259 1258
rect 287 1254 291 1258
rect 327 1254 331 1258
rect 351 1254 355 1258
rect 391 1254 395 1258
rect 415 1254 419 1258
rect 463 1254 467 1258
rect 479 1254 483 1258
rect 535 1254 539 1258
rect 543 1254 547 1258
rect 111 1218 115 1222
rect 135 1218 139 1222
rect 143 1218 147 1222
rect 175 1218 179 1222
rect 215 1218 219 1222
rect 231 1218 235 1222
rect 263 1218 267 1222
rect 287 1218 291 1222
rect 311 1218 315 1222
rect 111 1182 115 1186
rect 143 1182 147 1186
rect 175 1182 179 1186
rect 215 1182 219 1186
rect 599 1254 603 1258
rect 607 1254 611 1258
rect 351 1218 355 1222
rect 359 1218 363 1222
rect 415 1218 419 1222
rect 663 1254 667 1258
rect 671 1254 675 1258
rect 727 1254 731 1258
rect 735 1254 739 1258
rect 791 1254 795 1258
rect 799 1254 803 1258
rect 855 1290 859 1294
rect 887 1290 891 1294
rect 927 1290 931 1294
rect 935 1290 939 1294
rect 991 1290 995 1294
rect 999 1290 1003 1294
rect 855 1254 859 1258
rect 863 1254 867 1258
rect 1047 1290 1051 1294
rect 1271 1326 1275 1330
rect 1311 1326 1315 1330
rect 1327 1326 1331 1330
rect 1375 1326 1379 1330
rect 1383 1326 1387 1330
rect 1423 1326 1427 1330
rect 1447 1336 1451 1340
rect 1479 1362 1483 1366
rect 1535 1362 1539 1366
rect 1543 1362 1547 1366
rect 1583 1362 1587 1366
rect 1455 1326 1459 1330
rect 1471 1326 1475 1330
rect 1527 1326 1531 1330
rect 1535 1326 1539 1330
rect 1583 1326 1587 1330
rect 1063 1290 1067 1294
rect 1103 1290 1107 1294
rect 1127 1290 1131 1294
rect 1159 1290 1163 1294
rect 1191 1290 1195 1294
rect 1215 1290 1219 1294
rect 1247 1290 1251 1294
rect 1271 1290 1275 1294
rect 1303 1290 1307 1294
rect 1327 1290 1331 1294
rect 1367 1290 1371 1294
rect 1375 1290 1379 1294
rect 1423 1290 1427 1294
rect 1431 1290 1435 1294
rect 1471 1290 1475 1294
rect 1527 1290 1531 1294
rect 1583 1290 1587 1294
rect 927 1254 931 1258
rect 991 1254 995 1258
rect 999 1254 1003 1258
rect 1055 1254 1059 1258
rect 1063 1254 1067 1258
rect 1119 1254 1123 1258
rect 1127 1254 1131 1258
rect 1183 1254 1187 1258
rect 1191 1254 1195 1258
rect 1247 1254 1251 1258
rect 1303 1254 1307 1258
rect 1311 1254 1315 1258
rect 1367 1254 1371 1258
rect 1375 1254 1379 1258
rect 1431 1254 1435 1258
rect 1439 1254 1443 1258
rect 1503 1254 1507 1258
rect 1543 1254 1547 1258
rect 1583 1254 1587 1258
rect 471 1218 475 1222
rect 479 1218 483 1222
rect 527 1218 531 1222
rect 543 1218 547 1222
rect 583 1218 587 1222
rect 607 1218 611 1222
rect 639 1218 643 1222
rect 671 1218 675 1222
rect 687 1218 691 1222
rect 735 1218 739 1222
rect 783 1218 787 1222
rect 799 1218 803 1222
rect 831 1218 835 1222
rect 863 1218 867 1222
rect 879 1218 883 1222
rect 927 1218 931 1222
rect 935 1218 939 1222
rect 983 1218 987 1222
rect 991 1218 995 1222
rect 1039 1218 1043 1222
rect 1055 1218 1059 1222
rect 255 1182 259 1186
rect 263 1182 267 1186
rect 303 1182 307 1186
rect 311 1182 315 1186
rect 359 1182 363 1186
rect 415 1182 419 1186
rect 471 1182 475 1186
rect 527 1182 531 1186
rect 583 1182 587 1186
rect 591 1182 595 1186
rect 111 1146 115 1150
rect 135 1146 139 1150
rect 143 1146 147 1150
rect 639 1182 643 1186
rect 655 1182 659 1186
rect 687 1182 691 1186
rect 719 1182 723 1186
rect 735 1182 739 1186
rect 783 1182 787 1186
rect 791 1182 795 1186
rect 831 1182 835 1186
rect 855 1182 859 1186
rect 879 1182 883 1186
rect 919 1182 923 1186
rect 935 1182 939 1186
rect 983 1182 987 1186
rect 1095 1218 1099 1222
rect 1119 1218 1123 1222
rect 1159 1218 1163 1222
rect 1183 1218 1187 1222
rect 1231 1218 1235 1222
rect 1247 1218 1251 1222
rect 1303 1218 1307 1222
rect 1311 1218 1315 1222
rect 1375 1218 1379 1222
rect 1383 1218 1387 1222
rect 1439 1218 1443 1222
rect 1471 1218 1475 1222
rect 1503 1218 1507 1222
rect 1543 1218 1547 1222
rect 1583 1218 1587 1222
rect 1039 1182 1043 1186
rect 1095 1182 1099 1186
rect 1103 1182 1107 1186
rect 1159 1182 1163 1186
rect 1167 1182 1171 1186
rect 1231 1182 1235 1186
rect 1239 1182 1243 1186
rect 1303 1182 1307 1186
rect 1311 1182 1315 1186
rect 1383 1182 1387 1186
rect 1391 1182 1395 1186
rect 1471 1182 1475 1186
rect 1479 1182 1483 1186
rect 1543 1182 1547 1186
rect 1583 1182 1587 1186
rect 167 1146 171 1150
rect 175 1146 179 1150
rect 199 1146 203 1150
rect 215 1146 219 1150
rect 231 1146 235 1150
rect 255 1146 259 1150
rect 263 1146 267 1150
rect 295 1146 299 1150
rect 303 1146 307 1150
rect 327 1146 331 1150
rect 359 1146 363 1150
rect 391 1146 395 1150
rect 415 1146 419 1150
rect 447 1146 451 1150
rect 471 1146 475 1150
rect 503 1146 507 1150
rect 527 1146 531 1150
rect 559 1146 563 1150
rect 591 1146 595 1150
rect 615 1146 619 1150
rect 655 1146 659 1150
rect 671 1146 675 1150
rect 719 1146 723 1150
rect 727 1146 731 1150
rect 783 1146 787 1150
rect 791 1146 795 1150
rect 839 1146 843 1150
rect 855 1146 859 1150
rect 111 1110 115 1114
rect 135 1110 139 1114
rect 151 1110 155 1114
rect 167 1110 171 1114
rect 183 1110 187 1114
rect 199 1110 203 1114
rect 223 1110 227 1114
rect 231 1110 235 1114
rect 263 1110 267 1114
rect 271 1110 275 1114
rect 295 1110 299 1114
rect 167 1099 171 1100
rect 167 1096 171 1099
rect 895 1146 899 1150
rect 327 1110 331 1114
rect 311 1096 315 1100
rect 359 1110 363 1114
rect 383 1110 387 1114
rect 391 1110 395 1114
rect 439 1110 443 1114
rect 447 1110 451 1114
rect 503 1110 507 1114
rect 559 1110 563 1114
rect 567 1110 571 1114
rect 615 1110 619 1114
rect 639 1110 643 1114
rect 671 1110 675 1114
rect 711 1110 715 1114
rect 727 1110 731 1114
rect 783 1110 787 1114
rect 839 1110 843 1114
rect 855 1110 859 1114
rect 919 1146 923 1150
rect 951 1146 955 1150
rect 983 1146 987 1150
rect 1007 1146 1011 1150
rect 1039 1146 1043 1150
rect 1063 1146 1067 1150
rect 1103 1146 1107 1150
rect 1127 1146 1131 1150
rect 1167 1146 1171 1150
rect 1191 1146 1195 1150
rect 1239 1146 1243 1150
rect 895 1110 899 1114
rect 919 1110 923 1114
rect 951 1110 955 1114
rect 983 1110 987 1114
rect 1007 1110 1011 1114
rect 1039 1110 1043 1114
rect 1063 1110 1067 1114
rect 1095 1110 1099 1114
rect 1127 1110 1131 1114
rect 1151 1110 1155 1114
rect 1191 1110 1195 1114
rect 1207 1110 1211 1114
rect 1255 1146 1259 1150
rect 1311 1146 1315 1150
rect 1327 1146 1331 1150
rect 1391 1146 1395 1150
rect 1399 1146 1403 1150
rect 1255 1110 1259 1114
rect 1263 1110 1267 1114
rect 1319 1110 1323 1114
rect 1327 1110 1331 1114
rect 1375 1110 1379 1114
rect 1399 1110 1403 1114
rect 111 1066 115 1070
rect 151 1066 155 1070
rect 183 1066 187 1070
rect 223 1066 227 1070
rect 271 1066 275 1070
rect 327 1066 331 1070
rect 383 1066 387 1070
rect 439 1066 443 1070
rect 447 1066 451 1070
rect 487 1066 491 1070
rect 503 1066 507 1070
rect 543 1066 547 1070
rect 567 1066 571 1070
rect 599 1066 603 1070
rect 639 1066 643 1070
rect 663 1066 667 1070
rect 711 1066 715 1070
rect 727 1066 731 1070
rect 783 1066 787 1070
rect 791 1066 795 1070
rect 855 1066 859 1070
rect 863 1066 867 1070
rect 919 1066 923 1070
rect 935 1066 939 1070
rect 983 1066 987 1070
rect 1007 1066 1011 1070
rect 1039 1066 1043 1070
rect 1079 1066 1083 1070
rect 1095 1066 1099 1070
rect 1151 1066 1155 1070
rect 111 1026 115 1030
rect 447 1026 451 1030
rect 487 1026 491 1030
rect 511 1026 515 1030
rect 543 1026 547 1030
rect 575 1026 579 1030
rect 599 1026 603 1030
rect 615 1026 619 1030
rect 663 1026 667 1030
rect 711 1026 715 1030
rect 727 1026 731 1030
rect 775 1026 779 1030
rect 791 1026 795 1030
rect 847 1026 851 1030
rect 863 1026 867 1030
rect 927 1026 931 1030
rect 935 1026 939 1030
rect 1207 1066 1211 1070
rect 1215 1066 1219 1070
rect 1263 1066 1267 1070
rect 1279 1066 1283 1070
rect 1319 1066 1323 1070
rect 1335 1066 1339 1070
rect 1375 1066 1379 1070
rect 1007 1026 1011 1030
rect 1079 1026 1083 1030
rect 1087 1026 1091 1030
rect 1151 1026 1155 1030
rect 1167 1026 1171 1030
rect 1391 1066 1395 1070
rect 1479 1146 1483 1150
rect 1543 1146 1547 1150
rect 1583 1146 1587 1150
rect 1439 1110 1443 1114
rect 1479 1110 1483 1114
rect 1503 1110 1507 1114
rect 1543 1110 1547 1114
rect 1583 1110 1587 1114
rect 1439 1066 1443 1070
rect 1447 1066 1451 1070
rect 1503 1066 1507 1070
rect 1543 1066 1547 1070
rect 1215 1026 1219 1030
rect 1239 1026 1243 1030
rect 1279 1026 1283 1030
rect 1303 1026 1307 1030
rect 1335 1026 1339 1030
rect 1359 1026 1363 1030
rect 1391 1026 1395 1030
rect 1407 1026 1411 1030
rect 1447 1026 1451 1030
rect 1455 1026 1459 1030
rect 111 982 115 986
rect 159 982 163 986
rect 199 982 203 986
rect 255 982 259 986
rect 311 982 315 986
rect 375 982 379 986
rect 439 982 443 986
rect 503 982 507 986
rect 511 982 515 986
rect 543 982 547 986
rect 559 982 563 986
rect 575 982 579 986
rect 615 982 619 986
rect 663 982 667 986
rect 703 982 707 986
rect 711 982 715 986
rect 735 982 739 986
rect 775 982 779 986
rect 523 968 527 972
rect 587 971 591 972
rect 587 968 591 971
rect 111 946 115 950
rect 151 946 155 950
rect 159 946 163 950
rect 1503 1026 1507 1030
rect 1511 1026 1515 1030
rect 1583 1066 1587 1070
rect 1543 1026 1547 1030
rect 1583 1026 1587 1030
rect 831 982 835 986
rect 191 946 195 950
rect 199 946 203 950
rect 247 946 251 950
rect 255 946 259 950
rect 303 946 307 950
rect 311 946 315 950
rect 367 946 371 950
rect 375 946 379 950
rect 431 946 435 950
rect 439 946 443 950
rect 111 906 115 910
rect 135 906 139 910
rect 151 906 155 910
rect 167 906 171 910
rect 191 906 195 910
rect 223 906 227 910
rect 247 906 251 910
rect 111 870 115 874
rect 135 870 139 874
rect 279 906 283 910
rect 303 906 307 910
rect 495 946 499 950
rect 503 946 507 950
rect 559 946 563 950
rect 615 946 619 950
rect 663 946 667 950
rect 671 946 675 950
rect 703 946 707 950
rect 719 946 723 950
rect 735 946 739 950
rect 767 946 771 950
rect 775 946 779 950
rect 815 946 819 950
rect 847 982 851 986
rect 895 982 899 986
rect 927 982 931 986
rect 967 982 971 986
rect 1007 982 1011 986
rect 1047 982 1051 986
rect 1087 982 1091 986
rect 1127 982 1131 986
rect 1167 982 1171 986
rect 1199 982 1203 986
rect 1239 982 1243 986
rect 1271 982 1275 986
rect 1303 982 1307 986
rect 1343 982 1347 986
rect 1359 982 1363 986
rect 1407 982 1411 986
rect 1415 982 1419 986
rect 1455 982 1459 986
rect 1487 982 1491 986
rect 1511 982 1515 986
rect 1543 982 1547 986
rect 831 946 835 950
rect 871 946 875 950
rect 895 946 899 950
rect 935 946 939 950
rect 967 946 971 950
rect 1007 946 1011 950
rect 1047 946 1051 950
rect 1079 946 1083 950
rect 1127 946 1131 950
rect 1143 946 1147 950
rect 1199 946 1203 950
rect 1207 946 1211 950
rect 1583 982 1587 986
rect 1271 946 1275 950
rect 1327 946 1331 950
rect 1343 946 1347 950
rect 1375 946 1379 950
rect 1415 946 1419 950
rect 1423 946 1427 950
rect 1471 946 1475 950
rect 1487 946 1491 950
rect 1511 946 1515 950
rect 1543 946 1547 950
rect 1583 946 1587 950
rect 335 906 339 910
rect 367 906 371 910
rect 391 906 395 910
rect 431 906 435 910
rect 447 906 451 910
rect 495 906 499 910
rect 503 906 507 910
rect 559 906 563 910
rect 615 906 619 910
rect 623 906 627 910
rect 671 906 675 910
rect 695 906 699 910
rect 719 906 723 910
rect 759 906 763 910
rect 767 906 771 910
rect 815 906 819 910
rect 823 906 827 910
rect 871 906 875 910
rect 887 906 891 910
rect 935 906 939 910
rect 951 906 955 910
rect 1007 906 1011 910
rect 1015 906 1019 910
rect 1079 906 1083 910
rect 1135 906 1139 910
rect 1143 906 1147 910
rect 1191 906 1195 910
rect 1207 906 1211 910
rect 1247 906 1251 910
rect 1271 906 1275 910
rect 1303 906 1307 910
rect 1327 906 1331 910
rect 1359 906 1363 910
rect 167 870 171 874
rect 207 870 211 874
rect 223 870 227 874
rect 255 870 259 874
rect 279 870 283 874
rect 303 870 307 874
rect 335 870 339 874
rect 343 870 347 874
rect 383 870 387 874
rect 391 870 395 874
rect 439 870 443 874
rect 447 870 451 874
rect 111 830 115 834
rect 135 830 139 834
rect 167 830 171 834
rect 207 830 211 834
rect 111 794 115 798
rect 135 794 139 798
rect 223 830 227 834
rect 255 830 259 834
rect 503 870 507 874
rect 511 870 515 874
rect 559 870 563 874
rect 591 870 595 874
rect 623 870 627 874
rect 679 870 683 874
rect 695 870 699 874
rect 759 870 763 874
rect 767 870 771 874
rect 823 870 827 874
rect 847 870 851 874
rect 887 870 891 874
rect 919 870 923 874
rect 951 870 955 874
rect 983 870 987 874
rect 1015 870 1019 874
rect 1039 870 1043 874
rect 1079 870 1083 874
rect 1095 870 1099 874
rect 1135 870 1139 874
rect 1151 870 1155 874
rect 1191 870 1195 874
rect 1207 870 1211 874
rect 1247 870 1251 874
rect 1263 870 1267 874
rect 1375 906 1379 910
rect 1407 906 1411 910
rect 1423 906 1427 910
rect 1455 906 1459 910
rect 1471 906 1475 910
rect 1511 906 1515 910
rect 1543 906 1547 910
rect 1583 906 1587 910
rect 1303 870 1307 874
rect 1327 870 1331 874
rect 1359 870 1363 874
rect 1399 870 1403 874
rect 1407 870 1411 874
rect 1455 870 1459 874
rect 1479 870 1483 874
rect 1511 870 1515 874
rect 1543 870 1547 874
rect 1583 870 1587 874
rect 287 830 291 834
rect 303 830 307 834
rect 343 830 347 834
rect 351 830 355 834
rect 383 830 387 834
rect 423 830 427 834
rect 439 830 443 834
rect 495 830 499 834
rect 511 830 515 834
rect 567 830 571 834
rect 591 830 595 834
rect 639 830 643 834
rect 679 830 683 834
rect 719 830 723 834
rect 767 830 771 834
rect 791 830 795 834
rect 847 830 851 834
rect 863 830 867 834
rect 919 830 923 834
rect 935 830 939 834
rect 983 830 987 834
rect 999 830 1003 834
rect 167 794 171 798
rect 199 794 203 798
rect 223 794 227 798
rect 247 794 251 798
rect 287 794 291 798
rect 303 794 307 798
rect 351 794 355 798
rect 359 794 363 798
rect 423 794 427 798
rect 487 794 491 798
rect 495 794 499 798
rect 111 758 115 762
rect 135 758 139 762
rect 167 758 171 762
rect 199 758 203 762
rect 111 722 115 726
rect 135 722 139 726
rect 247 758 251 762
rect 255 758 259 762
rect 303 758 307 762
rect 319 758 323 762
rect 359 758 363 762
rect 391 758 395 762
rect 423 758 427 762
rect 463 758 467 762
rect 487 758 491 762
rect 551 794 555 798
rect 567 794 571 798
rect 607 794 611 798
rect 639 794 643 798
rect 671 794 675 798
rect 543 758 547 762
rect 551 758 555 762
rect 719 794 723 798
rect 735 794 739 798
rect 1039 830 1043 834
rect 1055 830 1059 834
rect 1095 830 1099 834
rect 1103 830 1107 834
rect 1143 830 1147 834
rect 1151 830 1155 834
rect 1183 830 1187 834
rect 1207 830 1211 834
rect 1231 830 1235 834
rect 1263 830 1267 834
rect 1279 830 1283 834
rect 1327 830 1331 834
rect 1399 830 1403 834
rect 1479 830 1483 834
rect 1543 830 1547 834
rect 1583 830 1587 834
rect 791 794 795 798
rect 799 794 803 798
rect 863 794 867 798
rect 871 794 875 798
rect 935 794 939 798
rect 999 794 1003 798
rect 607 758 611 762
rect 623 758 627 762
rect 671 758 675 762
rect 703 758 707 762
rect 735 758 739 762
rect 775 758 779 762
rect 799 758 803 762
rect 167 722 171 726
rect 199 722 203 726
rect 207 722 211 726
rect 255 722 259 726
rect 311 722 315 726
rect 319 722 323 726
rect 367 722 371 726
rect 391 722 395 726
rect 111 686 115 690
rect 135 686 139 690
rect 159 686 163 690
rect 167 686 171 690
rect 207 686 211 690
rect 111 646 115 650
rect 159 646 163 650
rect 167 646 171 650
rect 255 686 259 690
rect 423 722 427 726
rect 303 686 307 690
rect 311 686 315 690
rect 359 686 363 690
rect 367 686 371 690
rect 415 686 419 690
rect 423 686 427 690
rect 463 722 467 726
rect 479 722 483 726
rect 543 722 547 726
rect 615 722 619 726
rect 623 722 627 726
rect 687 722 691 726
rect 703 722 707 726
rect 759 722 763 726
rect 847 758 851 762
rect 871 758 875 762
rect 1055 794 1059 798
rect 1063 794 1067 798
rect 1103 794 1107 798
rect 1127 794 1131 798
rect 1143 794 1147 798
rect 1183 794 1187 798
rect 1191 794 1195 798
rect 1231 794 1235 798
rect 1255 794 1259 798
rect 1279 794 1283 798
rect 1319 794 1323 798
rect 1327 794 1331 798
rect 1383 794 1387 798
rect 1583 794 1587 798
rect 919 758 923 762
rect 935 758 939 762
rect 991 758 995 762
rect 999 758 1003 762
rect 1063 758 1067 762
rect 1127 758 1131 762
rect 1135 758 1139 762
rect 1191 758 1195 762
rect 1207 758 1211 762
rect 1255 758 1259 762
rect 1271 758 1275 762
rect 1319 758 1323 762
rect 471 686 475 690
rect 479 686 483 690
rect 527 686 531 690
rect 207 646 211 650
rect 215 646 219 650
rect 255 646 259 650
rect 271 646 275 650
rect 303 646 307 650
rect 327 646 331 650
rect 359 646 363 650
rect 383 646 387 650
rect 111 610 115 614
rect 167 610 171 614
rect 215 610 219 614
rect 223 610 227 614
rect 255 610 259 614
rect 271 610 275 614
rect 287 610 291 614
rect 111 574 115 578
rect 191 574 195 578
rect 319 610 323 614
rect 327 610 331 614
rect 415 646 419 650
rect 431 646 435 650
rect 351 610 355 614
rect 383 610 387 614
rect 423 610 427 614
rect 431 610 435 614
rect 471 646 475 650
rect 487 646 491 650
rect 543 686 547 690
rect 583 686 587 690
rect 615 686 619 690
rect 639 686 643 690
rect 775 722 779 726
rect 839 722 843 726
rect 847 722 851 726
rect 919 722 923 726
rect 991 722 995 726
rect 1007 722 1011 726
rect 687 686 691 690
rect 695 686 699 690
rect 759 686 763 690
rect 823 686 827 690
rect 839 686 843 690
rect 1063 722 1067 726
rect 1087 722 1091 726
rect 1135 722 1139 726
rect 1167 722 1171 726
rect 1327 758 1331 762
rect 1375 758 1379 762
rect 1383 758 1387 762
rect 1423 758 1427 762
rect 1471 758 1475 762
rect 1511 758 1515 762
rect 1543 758 1547 762
rect 1583 758 1587 762
rect 1207 722 1211 726
rect 1239 722 1243 726
rect 1271 722 1275 726
rect 1303 722 1307 726
rect 1327 722 1331 726
rect 1359 722 1363 726
rect 1375 722 1379 726
rect 1407 722 1411 726
rect 1423 722 1427 726
rect 1455 722 1459 726
rect 1471 722 1475 726
rect 1511 722 1515 726
rect 1543 722 1547 726
rect 1583 722 1587 726
rect 887 686 891 690
rect 919 686 923 690
rect 951 686 955 690
rect 1007 686 1011 690
rect 1015 686 1019 690
rect 527 646 531 650
rect 535 646 539 650
rect 583 646 587 650
rect 591 646 595 650
rect 639 646 643 650
rect 647 646 651 650
rect 695 646 699 650
rect 703 646 707 650
rect 759 646 763 650
rect 1079 686 1083 690
rect 1087 686 1091 690
rect 1135 686 1139 690
rect 1167 686 1171 690
rect 1191 686 1195 690
rect 1239 686 1243 690
rect 1247 686 1251 690
rect 1303 686 1307 690
rect 823 646 827 650
rect 887 646 891 650
rect 943 646 947 650
rect 463 610 467 614
rect 487 610 491 614
rect 519 610 523 614
rect 535 610 539 614
rect 583 610 587 614
rect 591 610 595 614
rect 647 610 651 614
rect 703 610 707 614
rect 719 610 723 614
rect 759 610 763 614
rect 799 610 803 614
rect 823 610 827 614
rect 951 646 955 650
rect 999 646 1003 650
rect 1015 646 1019 650
rect 1055 646 1059 650
rect 1079 646 1083 650
rect 1111 646 1115 650
rect 1135 646 1139 650
rect 1167 646 1171 650
rect 1359 686 1363 690
rect 1407 686 1411 690
rect 1455 686 1459 690
rect 1511 686 1515 690
rect 1543 686 1547 690
rect 1583 686 1587 690
rect 1191 646 1195 650
rect 1215 646 1219 650
rect 1247 646 1251 650
rect 1271 646 1275 650
rect 1303 646 1307 650
rect 1327 646 1331 650
rect 1359 646 1363 650
rect 1383 646 1387 650
rect 1439 646 1443 650
rect 1503 646 1507 650
rect 1543 646 1547 650
rect 1583 646 1587 650
rect 887 610 891 614
rect 943 610 947 614
rect 975 610 979 614
rect 999 610 1003 614
rect 1055 610 1059 614
rect 1063 610 1067 614
rect 1111 610 1115 614
rect 1143 610 1147 614
rect 1167 610 1171 614
rect 1215 610 1219 614
rect 1271 610 1275 614
rect 223 574 227 578
rect 255 574 259 578
rect 287 574 291 578
rect 319 574 323 578
rect 327 574 331 578
rect 351 574 355 578
rect 383 574 387 578
rect 399 574 403 578
rect 423 574 427 578
rect 463 574 467 578
rect 471 574 475 578
rect 519 574 523 578
rect 535 574 539 578
rect 583 574 587 578
rect 599 574 603 578
rect 647 574 651 578
rect 663 574 667 578
rect 719 574 723 578
rect 727 574 731 578
rect 783 574 787 578
rect 799 574 803 578
rect 839 574 843 578
rect 887 574 891 578
rect 903 574 907 578
rect 967 574 971 578
rect 975 574 979 578
rect 1039 574 1043 578
rect 1063 574 1067 578
rect 1103 574 1107 578
rect 1143 574 1147 578
rect 1167 574 1171 578
rect 1287 610 1291 614
rect 1327 610 1331 614
rect 1351 610 1355 614
rect 1383 610 1387 614
rect 1407 610 1411 614
rect 1439 610 1443 614
rect 1455 610 1459 614
rect 1503 610 1507 614
rect 1511 610 1515 614
rect 1543 610 1547 614
rect 1215 574 1219 578
rect 1231 574 1235 578
rect 1287 574 1291 578
rect 1335 574 1339 578
rect 1351 574 1355 578
rect 1383 574 1387 578
rect 1407 574 1411 578
rect 1423 574 1427 578
rect 1455 574 1459 578
rect 1471 574 1475 578
rect 111 538 115 542
rect 135 538 139 542
rect 175 538 179 542
rect 191 538 195 542
rect 231 538 235 542
rect 255 538 259 542
rect 295 538 299 542
rect 327 538 331 542
rect 111 502 115 506
rect 135 502 139 506
rect 1583 610 1587 614
rect 1511 574 1515 578
rect 1543 574 1547 578
rect 1583 574 1587 578
rect 359 538 363 542
rect 399 538 403 542
rect 423 538 427 542
rect 471 538 475 542
rect 479 538 483 542
rect 535 538 539 542
rect 543 538 547 542
rect 599 538 603 542
rect 655 538 659 542
rect 663 538 667 542
rect 711 538 715 542
rect 727 538 731 542
rect 767 538 771 542
rect 783 538 787 542
rect 831 538 835 542
rect 839 538 843 542
rect 895 538 899 542
rect 903 538 907 542
rect 967 538 971 542
rect 1031 538 1035 542
rect 1039 538 1043 542
rect 1095 538 1099 542
rect 1103 538 1107 542
rect 1167 538 1171 542
rect 1231 538 1235 542
rect 1239 538 1243 542
rect 1287 538 1291 542
rect 1311 538 1315 542
rect 1335 538 1339 542
rect 1383 538 1387 542
rect 1391 538 1395 542
rect 1423 538 1427 542
rect 1471 538 1475 542
rect 1479 538 1483 542
rect 1511 538 1515 542
rect 1543 538 1547 542
rect 167 502 171 506
rect 175 502 179 506
rect 199 502 203 506
rect 231 502 235 506
rect 247 502 251 506
rect 295 502 299 506
rect 343 502 347 506
rect 359 502 363 506
rect 111 466 115 470
rect 135 466 139 470
rect 167 466 171 470
rect 199 466 203 470
rect 247 466 251 470
rect 255 466 259 470
rect 111 426 115 430
rect 135 426 139 430
rect 295 466 299 470
rect 311 466 315 470
rect 399 502 403 506
rect 423 502 427 506
rect 455 502 459 506
rect 479 502 483 506
rect 511 502 515 506
rect 543 502 547 506
rect 567 502 571 506
rect 599 502 603 506
rect 623 502 627 506
rect 655 502 659 506
rect 679 502 683 506
rect 711 502 715 506
rect 343 466 347 470
rect 367 466 371 470
rect 399 466 403 470
rect 423 466 427 470
rect 743 502 747 506
rect 767 502 771 506
rect 815 502 819 506
rect 831 502 835 506
rect 887 502 891 506
rect 895 502 899 506
rect 959 502 963 506
rect 967 502 971 506
rect 1031 502 1035 506
rect 1039 502 1043 506
rect 1095 502 1099 506
rect 1127 502 1131 506
rect 1167 502 1171 506
rect 1223 502 1227 506
rect 1239 502 1243 506
rect 1311 502 1315 506
rect 1327 502 1331 506
rect 1391 502 1395 506
rect 1439 502 1443 506
rect 1479 502 1483 506
rect 1543 502 1547 506
rect 455 466 459 470
rect 479 466 483 470
rect 511 466 515 470
rect 535 466 539 470
rect 567 466 571 470
rect 599 466 603 470
rect 623 466 627 470
rect 663 466 667 470
rect 679 466 683 470
rect 735 466 739 470
rect 743 466 747 470
rect 807 466 811 470
rect 815 466 819 470
rect 871 466 875 470
rect 887 466 891 470
rect 935 466 939 470
rect 167 426 171 430
rect 199 426 203 430
rect 231 426 235 430
rect 255 426 259 430
rect 295 426 299 430
rect 311 426 315 430
rect 359 426 363 430
rect 367 426 371 430
rect 423 426 427 430
rect 479 426 483 430
rect 487 426 491 430
rect 535 426 539 430
rect 543 426 547 430
rect 591 426 595 430
rect 599 426 603 430
rect 639 426 643 430
rect 663 426 667 430
rect 679 426 683 430
rect 719 426 723 430
rect 735 426 739 430
rect 759 426 763 430
rect 959 466 963 470
rect 991 466 995 470
rect 1039 466 1043 470
rect 1047 466 1051 470
rect 1095 466 1099 470
rect 1127 466 1131 470
rect 1143 466 1147 470
rect 1199 466 1203 470
rect 1223 466 1227 470
rect 1263 466 1267 470
rect 807 426 811 430
rect 863 426 867 430
rect 871 426 875 430
rect 919 426 923 430
rect 935 426 939 430
rect 975 426 979 430
rect 991 426 995 430
rect 1031 426 1035 430
rect 1327 466 1331 470
rect 1399 466 1403 470
rect 1439 466 1443 470
rect 1479 466 1483 470
rect 1583 538 1587 542
rect 1583 502 1587 506
rect 1543 466 1547 470
rect 1583 466 1587 470
rect 1047 426 1051 430
rect 1087 426 1091 430
rect 1095 426 1099 430
rect 1143 426 1147 430
rect 1151 426 1155 430
rect 1199 426 1203 430
rect 1223 426 1227 430
rect 1263 426 1267 430
rect 1303 426 1307 430
rect 1327 426 1331 430
rect 1383 426 1387 430
rect 1399 426 1403 430
rect 1471 426 1475 430
rect 1479 426 1483 430
rect 1543 426 1547 430
rect 1583 426 1587 430
rect 111 390 115 394
rect 135 390 139 394
rect 167 390 171 394
rect 207 390 211 394
rect 231 390 235 394
rect 295 390 299 394
rect 111 354 115 358
rect 135 354 139 358
rect 359 390 363 394
rect 383 390 387 394
rect 423 390 427 394
rect 463 390 467 394
rect 487 390 491 394
rect 535 390 539 394
rect 543 390 547 394
rect 591 390 595 394
rect 599 390 603 394
rect 639 390 643 394
rect 655 390 659 394
rect 679 390 683 394
rect 703 390 707 394
rect 719 390 723 394
rect 751 390 755 394
rect 759 390 763 394
rect 807 390 811 394
rect 863 390 867 394
rect 919 390 923 394
rect 975 390 979 394
rect 983 390 987 394
rect 1031 390 1035 394
rect 1055 390 1059 394
rect 1087 390 1091 394
rect 1127 390 1131 394
rect 1151 390 1155 394
rect 1199 390 1203 394
rect 175 354 179 358
rect 207 354 211 358
rect 223 354 227 358
rect 279 354 283 358
rect 295 354 299 358
rect 335 354 339 358
rect 383 354 387 358
rect 391 354 395 358
rect 447 354 451 358
rect 463 354 467 358
rect 503 354 507 358
rect 535 354 539 358
rect 567 354 571 358
rect 111 318 115 322
rect 135 318 139 322
rect 175 318 179 322
rect 191 318 195 322
rect 223 318 227 322
rect 255 318 259 322
rect 279 318 283 322
rect 295 318 299 322
rect 111 278 115 282
rect 151 278 155 282
rect 335 318 339 322
rect 367 318 371 322
rect 391 318 395 322
rect 407 318 411 322
rect 447 318 451 322
rect 455 318 459 322
rect 183 278 187 282
rect 191 278 195 282
rect 215 278 219 282
rect 223 278 227 282
rect 247 278 251 282
rect 255 278 259 282
rect 279 278 283 282
rect 295 278 299 282
rect 311 278 315 282
rect 335 278 339 282
rect 111 242 115 246
rect 135 242 139 246
rect 151 242 155 246
rect 167 242 171 246
rect 183 242 187 246
rect 207 242 211 246
rect 215 242 219 246
rect 111 202 115 206
rect 135 202 139 206
rect 247 242 251 246
rect 255 242 259 246
rect 599 354 603 358
rect 631 354 635 358
rect 655 354 659 358
rect 687 354 691 358
rect 703 354 707 358
rect 751 354 755 358
rect 807 354 811 358
rect 815 354 819 358
rect 863 354 867 358
rect 879 354 883 358
rect 919 354 923 358
rect 951 354 955 358
rect 983 354 987 358
rect 1031 354 1035 358
rect 1055 354 1059 358
rect 1223 390 1227 394
rect 1271 390 1275 394
rect 1303 390 1307 394
rect 1343 390 1347 394
rect 1383 390 1387 394
rect 1415 390 1419 394
rect 1471 390 1475 394
rect 1487 390 1491 394
rect 1543 390 1547 394
rect 1103 354 1107 358
rect 1127 354 1131 358
rect 1175 354 1179 358
rect 1199 354 1203 358
rect 1247 354 1251 358
rect 1271 354 1275 358
rect 1327 354 1331 358
rect 1343 354 1347 358
rect 1583 390 1587 394
rect 1407 354 1411 358
rect 1415 354 1419 358
rect 1487 354 1491 358
rect 1543 354 1547 358
rect 1583 354 1587 358
rect 503 318 507 322
rect 519 318 523 322
rect 567 318 571 322
rect 591 318 595 322
rect 631 318 635 322
rect 663 318 667 322
rect 687 318 691 322
rect 735 318 739 322
rect 751 318 755 322
rect 807 318 811 322
rect 815 318 819 322
rect 879 318 883 322
rect 351 278 355 282
rect 367 278 371 282
rect 407 278 411 282
rect 455 278 459 282
rect 479 278 483 282
rect 519 278 523 282
rect 559 278 563 282
rect 591 278 595 282
rect 647 278 651 282
rect 279 242 283 246
rect 303 242 307 246
rect 311 242 315 246
rect 343 242 347 246
rect 351 242 355 246
rect 383 242 387 246
rect 951 318 955 322
rect 1023 318 1027 322
rect 1031 318 1035 322
rect 1095 318 1099 322
rect 1103 318 1107 322
rect 1167 318 1171 322
rect 1175 318 1179 322
rect 1231 318 1235 322
rect 1247 318 1251 322
rect 1295 318 1299 322
rect 1327 318 1331 322
rect 1351 318 1355 322
rect 1399 318 1403 322
rect 1407 318 1411 322
rect 1455 318 1459 322
rect 1487 318 1491 322
rect 1511 318 1515 322
rect 1543 318 1547 322
rect 1583 318 1587 322
rect 663 278 667 282
rect 735 278 739 282
rect 807 278 811 282
rect 823 278 827 282
rect 879 278 883 282
rect 903 278 907 282
rect 951 278 955 282
rect 983 278 987 282
rect 1023 278 1027 282
rect 1055 278 1059 282
rect 1095 278 1099 282
rect 1119 278 1123 282
rect 1167 278 1171 282
rect 1175 278 1179 282
rect 1223 278 1227 282
rect 1231 278 1235 282
rect 1263 278 1267 282
rect 1295 278 1299 282
rect 1303 278 1307 282
rect 1351 278 1355 282
rect 1399 278 1403 282
rect 1447 278 1451 282
rect 1455 278 1459 282
rect 1503 278 1507 282
rect 1511 278 1515 282
rect 1543 278 1547 282
rect 1583 278 1587 282
rect 407 242 411 246
rect 439 242 443 246
rect 479 242 483 246
rect 167 202 171 206
rect 207 202 211 206
rect 215 202 219 206
rect 255 202 259 206
rect 263 202 267 206
rect 303 202 307 206
rect 311 202 315 206
rect 343 202 347 206
rect 359 202 363 206
rect 111 166 115 170
rect 135 166 139 170
rect 143 166 147 170
rect 167 166 171 170
rect 191 166 195 170
rect 215 166 219 170
rect 239 166 243 170
rect 263 166 267 170
rect 111 118 115 122
rect 135 118 139 122
rect 143 118 147 122
rect 295 166 299 170
rect 311 166 315 170
rect 383 202 387 206
rect 415 202 419 206
rect 439 202 443 206
rect 511 242 515 246
rect 559 242 563 246
rect 591 242 595 246
rect 647 242 651 246
rect 679 242 683 246
rect 735 242 739 246
rect 767 242 771 246
rect 823 242 827 246
rect 847 242 851 246
rect 903 242 907 246
rect 919 242 923 246
rect 983 242 987 246
rect 1047 242 1051 246
rect 1055 242 1059 246
rect 1103 242 1107 246
rect 1119 242 1123 246
rect 1159 242 1163 246
rect 1175 242 1179 246
rect 471 202 475 206
rect 511 202 515 206
rect 535 202 539 206
rect 591 202 595 206
rect 607 202 611 206
rect 679 202 683 206
rect 751 202 755 206
rect 351 166 355 170
rect 359 166 363 170
rect 407 166 411 170
rect 415 166 419 170
rect 463 166 467 170
rect 471 166 475 170
rect 519 166 523 170
rect 535 166 539 170
rect 575 166 579 170
rect 607 166 611 170
rect 767 202 771 206
rect 815 202 819 206
rect 847 202 851 206
rect 879 202 883 206
rect 919 202 923 206
rect 943 202 947 206
rect 983 202 987 206
rect 1007 202 1011 206
rect 1215 242 1219 246
rect 1223 242 1227 246
rect 1263 242 1267 246
rect 1271 242 1275 246
rect 1303 242 1307 246
rect 1327 242 1331 246
rect 1351 242 1355 246
rect 1047 202 1051 206
rect 1063 202 1067 206
rect 1103 202 1107 206
rect 1119 202 1123 206
rect 1159 202 1163 206
rect 1175 202 1179 206
rect 1215 202 1219 206
rect 1231 202 1235 206
rect 1383 242 1387 246
rect 1399 242 1403 246
rect 1439 242 1443 246
rect 1447 242 1451 246
rect 1503 242 1507 246
rect 1543 242 1547 246
rect 1583 242 1587 246
rect 1271 202 1275 206
rect 1287 202 1291 206
rect 1327 202 1331 206
rect 1343 202 1347 206
rect 1383 202 1387 206
rect 1399 202 1403 206
rect 1439 202 1443 206
rect 1455 202 1459 206
rect 1503 202 1507 206
rect 631 166 635 170
rect 679 166 683 170
rect 687 166 691 170
rect 743 166 747 170
rect 751 166 755 170
rect 799 166 803 170
rect 815 166 819 170
rect 855 166 859 170
rect 879 166 883 170
rect 911 166 915 170
rect 943 166 947 170
rect 975 166 979 170
rect 1007 166 1011 170
rect 1039 166 1043 170
rect 1063 166 1067 170
rect 1095 166 1099 170
rect 1119 166 1123 170
rect 1151 166 1155 170
rect 1175 166 1179 170
rect 167 118 171 122
rect 191 118 195 122
rect 199 118 203 122
rect 231 118 235 122
rect 239 118 243 122
rect 263 118 267 122
rect 295 118 299 122
rect 327 118 331 122
rect 351 118 355 122
rect 359 118 363 122
rect 391 118 395 122
rect 407 118 411 122
rect 423 118 427 122
rect 455 118 459 122
rect 463 118 467 122
rect 487 118 491 122
rect 519 118 523 122
rect 1207 166 1211 170
rect 1231 166 1235 170
rect 1255 166 1259 170
rect 1287 166 1291 170
rect 1303 166 1307 170
rect 1343 166 1347 170
rect 1351 166 1355 170
rect 1511 202 1515 206
rect 1543 202 1547 206
rect 1583 202 1587 206
rect 1399 166 1403 170
rect 1455 166 1459 170
rect 1511 166 1515 170
rect 1543 166 1547 170
rect 1583 166 1587 170
rect 551 118 555 122
rect 575 118 579 122
rect 583 118 587 122
rect 615 118 619 122
rect 631 118 635 122
rect 647 118 651 122
rect 679 118 683 122
rect 687 118 691 122
rect 711 118 715 122
rect 743 118 747 122
rect 775 118 779 122
rect 799 118 803 122
rect 807 118 811 122
rect 839 118 843 122
rect 855 118 859 122
rect 871 118 875 122
rect 903 118 907 122
rect 911 118 915 122
rect 943 118 947 122
rect 975 118 979 122
rect 983 118 987 122
rect 1031 118 1035 122
rect 1039 118 1043 122
rect 1079 118 1083 122
rect 1095 118 1099 122
rect 1127 118 1131 122
rect 1151 118 1155 122
rect 1175 118 1179 122
rect 1207 118 1211 122
rect 1223 118 1227 122
rect 1255 118 1259 122
rect 1263 118 1267 122
rect 1303 118 1307 122
rect 1343 118 1347 122
rect 1351 118 1355 122
rect 1383 118 1387 122
rect 1399 118 1403 122
rect 1423 118 1427 122
rect 1455 118 1459 122
rect 1471 118 1475 122
rect 1511 118 1515 122
rect 1543 118 1547 122
rect 1583 118 1587 122
rect 111 82 115 86
rect 135 82 139 86
rect 167 82 171 86
rect 199 82 203 86
rect 231 82 235 86
rect 263 82 267 86
rect 295 82 299 86
rect 327 82 331 86
rect 359 82 363 86
rect 391 82 395 86
rect 423 82 427 86
rect 455 82 459 86
rect 487 82 491 86
rect 519 82 523 86
rect 551 82 555 86
rect 583 82 587 86
rect 615 82 619 86
rect 647 82 651 86
rect 679 82 683 86
rect 711 82 715 86
rect 743 82 747 86
rect 775 82 779 86
rect 807 82 811 86
rect 839 82 843 86
rect 871 82 875 86
rect 903 82 907 86
rect 943 82 947 86
rect 983 82 987 86
rect 1031 82 1035 86
rect 1079 82 1083 86
rect 1127 82 1131 86
rect 1175 82 1179 86
rect 1223 82 1227 86
rect 1263 82 1267 86
rect 1303 82 1307 86
rect 1343 82 1347 86
rect 1383 82 1387 86
rect 1423 82 1427 86
rect 1471 82 1475 86
rect 1511 82 1515 86
rect 1543 82 1547 86
rect 1583 82 1587 86
<< m4 >>
rect 84 1649 85 1655
rect 91 1654 1607 1655
rect 91 1650 111 1654
rect 115 1650 135 1654
rect 139 1650 167 1654
rect 171 1650 199 1654
rect 203 1650 1583 1654
rect 1587 1650 1607 1654
rect 91 1649 1607 1650
rect 1613 1649 1614 1655
rect 96 1613 97 1619
rect 103 1618 1619 1619
rect 103 1614 111 1618
rect 115 1614 135 1618
rect 139 1614 167 1618
rect 171 1614 175 1618
rect 179 1614 199 1618
rect 203 1614 239 1618
rect 243 1614 295 1618
rect 299 1614 351 1618
rect 355 1614 407 1618
rect 411 1614 455 1618
rect 459 1614 503 1618
rect 507 1614 551 1618
rect 555 1614 599 1618
rect 603 1614 647 1618
rect 651 1614 695 1618
rect 699 1614 743 1618
rect 747 1614 791 1618
rect 795 1614 839 1618
rect 843 1614 887 1618
rect 891 1614 935 1618
rect 939 1614 991 1618
rect 995 1614 1047 1618
rect 1051 1614 1095 1618
rect 1099 1614 1143 1618
rect 1147 1614 1191 1618
rect 1195 1614 1239 1618
rect 1243 1614 1287 1618
rect 1291 1614 1327 1618
rect 1331 1614 1367 1618
rect 1371 1614 1407 1618
rect 1411 1614 1447 1618
rect 1451 1614 1479 1618
rect 1483 1614 1511 1618
rect 1515 1614 1543 1618
rect 1547 1614 1583 1618
rect 1587 1614 1619 1618
rect 103 1613 1619 1614
rect 1625 1613 1626 1619
rect 84 1577 85 1583
rect 91 1582 1607 1583
rect 91 1578 111 1582
rect 115 1578 135 1582
rect 139 1578 175 1582
rect 179 1578 215 1582
rect 219 1578 239 1582
rect 243 1578 255 1582
rect 259 1578 295 1582
rect 299 1578 343 1582
rect 347 1578 351 1582
rect 355 1578 391 1582
rect 395 1578 407 1582
rect 411 1578 439 1582
rect 443 1578 455 1582
rect 459 1578 487 1582
rect 491 1578 503 1582
rect 507 1578 535 1582
rect 539 1578 551 1582
rect 555 1578 583 1582
rect 587 1578 599 1582
rect 603 1578 639 1582
rect 643 1578 647 1582
rect 651 1578 695 1582
rect 699 1578 703 1582
rect 707 1578 743 1582
rect 747 1578 775 1582
rect 779 1578 791 1582
rect 795 1578 839 1582
rect 843 1578 855 1582
rect 859 1578 887 1582
rect 891 1578 935 1582
rect 939 1578 991 1582
rect 995 1578 1015 1582
rect 1019 1578 1047 1582
rect 1051 1578 1087 1582
rect 1091 1578 1095 1582
rect 1099 1578 1143 1582
rect 1147 1578 1159 1582
rect 1163 1578 1191 1582
rect 1195 1578 1239 1582
rect 1243 1578 1287 1582
rect 1291 1578 1319 1582
rect 1323 1578 1327 1582
rect 1331 1578 1367 1582
rect 1371 1578 1399 1582
rect 1403 1578 1407 1582
rect 1411 1578 1447 1582
rect 1451 1578 1479 1582
rect 1483 1578 1511 1582
rect 1515 1578 1543 1582
rect 1547 1578 1583 1582
rect 1587 1578 1607 1582
rect 91 1577 1607 1578
rect 1613 1577 1614 1583
rect 96 1541 97 1547
rect 103 1546 1619 1547
rect 103 1542 111 1546
rect 115 1542 159 1546
rect 163 1542 175 1546
rect 179 1542 207 1546
rect 211 1542 215 1546
rect 219 1542 255 1546
rect 259 1542 295 1546
rect 299 1542 311 1546
rect 315 1542 343 1546
rect 347 1542 359 1546
rect 363 1542 391 1546
rect 395 1542 415 1546
rect 419 1542 439 1546
rect 443 1542 471 1546
rect 475 1542 487 1546
rect 491 1542 527 1546
rect 531 1542 535 1546
rect 539 1542 583 1546
rect 587 1542 639 1546
rect 643 1542 695 1546
rect 699 1542 703 1546
rect 707 1542 759 1546
rect 763 1542 775 1546
rect 779 1542 823 1546
rect 827 1542 855 1546
rect 859 1542 895 1546
rect 899 1542 935 1546
rect 939 1542 967 1546
rect 971 1542 1015 1546
rect 1019 1542 1039 1546
rect 1043 1542 1087 1546
rect 1091 1542 1103 1546
rect 1107 1542 1159 1546
rect 1163 1542 1167 1546
rect 1171 1542 1231 1546
rect 1235 1542 1239 1546
rect 1243 1542 1295 1546
rect 1299 1542 1319 1546
rect 1323 1542 1359 1546
rect 1363 1542 1399 1546
rect 1403 1542 1423 1546
rect 1427 1542 1479 1546
rect 1483 1542 1495 1546
rect 1499 1542 1543 1546
rect 1547 1542 1583 1546
rect 1587 1542 1619 1546
rect 103 1541 1619 1542
rect 1625 1541 1626 1547
rect 84 1505 85 1511
rect 91 1510 1607 1511
rect 91 1506 111 1510
rect 115 1506 159 1510
rect 163 1506 207 1510
rect 211 1506 255 1510
rect 259 1506 303 1510
rect 307 1506 311 1510
rect 315 1506 351 1510
rect 355 1506 359 1510
rect 363 1506 407 1510
rect 411 1506 415 1510
rect 419 1506 463 1510
rect 467 1506 471 1510
rect 475 1506 527 1510
rect 531 1506 583 1510
rect 587 1506 591 1510
rect 595 1506 639 1510
rect 643 1506 655 1510
rect 659 1506 695 1510
rect 699 1506 719 1510
rect 723 1506 759 1510
rect 763 1506 783 1510
rect 787 1506 823 1510
rect 827 1506 855 1510
rect 859 1506 895 1510
rect 899 1506 935 1510
rect 939 1506 967 1510
rect 971 1506 1007 1510
rect 1011 1506 1039 1510
rect 1043 1506 1079 1510
rect 1083 1506 1103 1510
rect 1107 1506 1151 1510
rect 1155 1506 1167 1510
rect 1171 1506 1215 1510
rect 1219 1506 1231 1510
rect 1235 1506 1279 1510
rect 1283 1506 1295 1510
rect 1299 1506 1351 1510
rect 1355 1506 1359 1510
rect 1363 1506 1423 1510
rect 1427 1506 1495 1510
rect 1499 1506 1543 1510
rect 1547 1506 1583 1510
rect 1587 1506 1607 1510
rect 91 1505 1607 1506
rect 1613 1505 1614 1511
rect 96 1469 97 1475
rect 103 1474 1619 1475
rect 103 1470 111 1474
rect 115 1470 135 1474
rect 139 1470 159 1474
rect 163 1470 183 1474
rect 187 1470 207 1474
rect 211 1470 231 1474
rect 235 1470 255 1474
rect 259 1470 287 1474
rect 291 1470 303 1474
rect 307 1470 343 1474
rect 347 1470 351 1474
rect 355 1470 399 1474
rect 403 1470 407 1474
rect 411 1470 455 1474
rect 459 1470 463 1474
rect 467 1470 511 1474
rect 515 1470 527 1474
rect 531 1470 575 1474
rect 579 1470 591 1474
rect 595 1470 631 1474
rect 635 1470 655 1474
rect 659 1470 687 1474
rect 691 1470 719 1474
rect 723 1470 751 1474
rect 755 1470 783 1474
rect 787 1470 815 1474
rect 819 1470 855 1474
rect 859 1470 879 1474
rect 883 1470 935 1474
rect 939 1470 943 1474
rect 947 1470 1007 1474
rect 1011 1470 1015 1474
rect 1019 1470 1079 1474
rect 1083 1470 1087 1474
rect 1091 1470 1151 1474
rect 1155 1470 1159 1474
rect 1163 1470 1215 1474
rect 1219 1470 1239 1474
rect 1243 1470 1279 1474
rect 1283 1470 1319 1474
rect 1323 1470 1351 1474
rect 1355 1470 1399 1474
rect 1403 1470 1423 1474
rect 1427 1470 1479 1474
rect 1483 1470 1495 1474
rect 1499 1470 1543 1474
rect 1547 1470 1583 1474
rect 1587 1470 1619 1474
rect 103 1469 1619 1470
rect 1625 1469 1626 1475
rect 258 1460 264 1461
rect 414 1460 420 1461
rect 258 1456 259 1460
rect 263 1456 415 1460
rect 419 1456 420 1460
rect 258 1455 264 1456
rect 414 1455 420 1456
rect 84 1433 85 1439
rect 91 1438 1607 1439
rect 91 1434 111 1438
rect 115 1434 135 1438
rect 139 1434 183 1438
rect 187 1434 231 1438
rect 235 1434 255 1438
rect 259 1434 287 1438
rect 291 1434 327 1438
rect 331 1434 343 1438
rect 347 1434 399 1438
rect 403 1434 455 1438
rect 459 1434 471 1438
rect 475 1434 511 1438
rect 515 1434 543 1438
rect 547 1434 575 1438
rect 579 1434 615 1438
rect 619 1434 631 1438
rect 635 1434 679 1438
rect 683 1434 687 1438
rect 691 1434 743 1438
rect 747 1434 751 1438
rect 755 1434 815 1438
rect 819 1434 879 1438
rect 883 1434 943 1438
rect 947 1434 951 1438
rect 955 1434 1015 1438
rect 1019 1434 1023 1438
rect 1027 1434 1087 1438
rect 1091 1434 1095 1438
rect 1099 1434 1159 1438
rect 1163 1434 1223 1438
rect 1227 1434 1239 1438
rect 1243 1434 1287 1438
rect 1291 1434 1319 1438
rect 1323 1434 1343 1438
rect 1347 1434 1399 1438
rect 1403 1434 1455 1438
rect 1459 1434 1479 1438
rect 1483 1434 1511 1438
rect 1515 1434 1543 1438
rect 1547 1434 1583 1438
rect 1587 1434 1607 1438
rect 91 1433 1607 1434
rect 1613 1433 1614 1439
rect 96 1397 97 1403
rect 103 1402 1619 1403
rect 103 1398 111 1402
rect 115 1398 135 1402
rect 139 1398 175 1402
rect 179 1398 183 1402
rect 187 1398 247 1402
rect 251 1398 255 1402
rect 259 1398 319 1402
rect 323 1398 327 1402
rect 331 1398 391 1402
rect 395 1398 399 1402
rect 403 1398 455 1402
rect 459 1398 471 1402
rect 475 1398 519 1402
rect 523 1398 543 1402
rect 547 1398 583 1402
rect 587 1398 615 1402
rect 619 1398 647 1402
rect 651 1398 679 1402
rect 683 1398 711 1402
rect 715 1398 743 1402
rect 747 1398 775 1402
rect 779 1398 815 1402
rect 819 1398 839 1402
rect 843 1398 879 1402
rect 883 1398 895 1402
rect 899 1398 951 1402
rect 955 1398 999 1402
rect 1003 1398 1023 1402
rect 1027 1398 1055 1402
rect 1059 1398 1095 1402
rect 1099 1398 1111 1402
rect 1115 1398 1159 1402
rect 1163 1398 1175 1402
rect 1179 1398 1223 1402
rect 1227 1398 1239 1402
rect 1243 1398 1287 1402
rect 1291 1398 1295 1402
rect 1299 1398 1343 1402
rect 1347 1398 1351 1402
rect 1355 1398 1399 1402
rect 1403 1398 1415 1402
rect 1419 1398 1455 1402
rect 1459 1398 1479 1402
rect 1483 1398 1511 1402
rect 1515 1398 1543 1402
rect 1547 1398 1583 1402
rect 1587 1398 1619 1402
rect 103 1397 1619 1398
rect 1625 1397 1626 1403
rect 84 1361 85 1367
rect 91 1366 1607 1367
rect 91 1362 111 1366
rect 115 1362 135 1366
rect 139 1362 167 1366
rect 171 1362 175 1366
rect 179 1362 215 1366
rect 219 1362 247 1366
rect 251 1362 303 1366
rect 307 1362 319 1366
rect 323 1362 391 1366
rect 395 1362 415 1366
rect 419 1362 455 1366
rect 459 1362 519 1366
rect 523 1362 527 1366
rect 531 1362 583 1366
rect 587 1362 639 1366
rect 643 1362 647 1366
rect 651 1362 711 1366
rect 715 1362 751 1366
rect 755 1362 775 1366
rect 779 1362 839 1366
rect 843 1362 863 1366
rect 867 1362 895 1366
rect 899 1362 951 1366
rect 955 1362 967 1366
rect 971 1362 999 1366
rect 1003 1362 1055 1366
rect 1059 1362 1063 1366
rect 1067 1362 1111 1366
rect 1115 1362 1151 1366
rect 1155 1362 1175 1366
rect 1179 1362 1231 1366
rect 1235 1362 1239 1366
rect 1243 1362 1295 1366
rect 1299 1362 1311 1366
rect 1315 1362 1351 1366
rect 1355 1362 1383 1366
rect 1387 1362 1415 1366
rect 1419 1362 1455 1366
rect 1459 1362 1479 1366
rect 1483 1362 1535 1366
rect 1539 1362 1543 1366
rect 1547 1362 1583 1366
rect 1587 1362 1607 1366
rect 91 1361 1607 1362
rect 1613 1361 1614 1367
rect 1354 1340 1360 1341
rect 1446 1340 1452 1341
rect 1354 1336 1355 1340
rect 1359 1336 1447 1340
rect 1451 1336 1452 1340
rect 1354 1335 1360 1336
rect 1446 1335 1452 1336
rect 96 1325 97 1331
rect 103 1330 1619 1331
rect 103 1326 111 1330
rect 115 1326 135 1330
rect 139 1326 167 1330
rect 171 1326 183 1330
rect 187 1326 215 1330
rect 219 1326 247 1330
rect 251 1326 303 1330
rect 307 1326 311 1330
rect 315 1326 375 1330
rect 379 1326 415 1330
rect 419 1326 439 1330
rect 443 1326 495 1330
rect 499 1326 527 1330
rect 531 1326 543 1330
rect 547 1326 591 1330
rect 595 1326 639 1330
rect 643 1326 687 1330
rect 691 1326 743 1330
rect 747 1326 751 1330
rect 755 1326 791 1330
rect 795 1326 839 1330
rect 843 1326 863 1330
rect 867 1326 887 1330
rect 891 1326 935 1330
rect 939 1326 967 1330
rect 971 1326 991 1330
rect 995 1326 1047 1330
rect 1051 1326 1063 1330
rect 1067 1326 1103 1330
rect 1107 1326 1151 1330
rect 1155 1326 1159 1330
rect 1163 1326 1215 1330
rect 1219 1326 1231 1330
rect 1235 1326 1271 1330
rect 1275 1326 1311 1330
rect 1315 1326 1327 1330
rect 1331 1326 1375 1330
rect 1379 1326 1383 1330
rect 1387 1326 1423 1330
rect 1427 1326 1455 1330
rect 1459 1326 1471 1330
rect 1475 1326 1527 1330
rect 1531 1326 1535 1330
rect 1539 1326 1583 1330
rect 1587 1326 1619 1330
rect 103 1325 1619 1326
rect 1625 1325 1626 1331
rect 84 1289 85 1295
rect 91 1294 1607 1295
rect 91 1290 111 1294
rect 115 1290 135 1294
rect 139 1290 183 1294
rect 187 1290 191 1294
rect 195 1290 247 1294
rect 251 1290 255 1294
rect 259 1290 311 1294
rect 315 1290 327 1294
rect 331 1290 375 1294
rect 379 1290 391 1294
rect 395 1290 439 1294
rect 443 1290 463 1294
rect 467 1290 495 1294
rect 499 1290 535 1294
rect 539 1290 543 1294
rect 547 1290 591 1294
rect 595 1290 599 1294
rect 603 1290 639 1294
rect 643 1290 663 1294
rect 667 1290 687 1294
rect 691 1290 727 1294
rect 731 1290 743 1294
rect 747 1290 791 1294
rect 795 1290 839 1294
rect 843 1290 855 1294
rect 859 1290 887 1294
rect 891 1290 927 1294
rect 931 1290 935 1294
rect 939 1290 991 1294
rect 995 1290 999 1294
rect 1003 1290 1047 1294
rect 1051 1290 1063 1294
rect 1067 1290 1103 1294
rect 1107 1290 1127 1294
rect 1131 1290 1159 1294
rect 1163 1290 1191 1294
rect 1195 1290 1215 1294
rect 1219 1290 1247 1294
rect 1251 1290 1271 1294
rect 1275 1290 1303 1294
rect 1307 1290 1327 1294
rect 1331 1290 1367 1294
rect 1371 1290 1375 1294
rect 1379 1290 1423 1294
rect 1427 1290 1431 1294
rect 1435 1290 1471 1294
rect 1475 1290 1527 1294
rect 1531 1290 1583 1294
rect 1587 1290 1607 1294
rect 91 1289 1607 1290
rect 1613 1289 1614 1295
rect 96 1253 97 1259
rect 103 1258 1619 1259
rect 103 1254 111 1258
rect 115 1254 135 1258
rect 139 1254 175 1258
rect 179 1254 191 1258
rect 195 1254 231 1258
rect 235 1254 255 1258
rect 259 1254 287 1258
rect 291 1254 327 1258
rect 331 1254 351 1258
rect 355 1254 391 1258
rect 395 1254 415 1258
rect 419 1254 463 1258
rect 467 1254 479 1258
rect 483 1254 535 1258
rect 539 1254 543 1258
rect 547 1254 599 1258
rect 603 1254 607 1258
rect 611 1254 663 1258
rect 667 1254 671 1258
rect 675 1254 727 1258
rect 731 1254 735 1258
rect 739 1254 791 1258
rect 795 1254 799 1258
rect 803 1254 855 1258
rect 859 1254 863 1258
rect 867 1254 927 1258
rect 931 1254 991 1258
rect 995 1254 999 1258
rect 1003 1254 1055 1258
rect 1059 1254 1063 1258
rect 1067 1254 1119 1258
rect 1123 1254 1127 1258
rect 1131 1254 1183 1258
rect 1187 1254 1191 1258
rect 1195 1254 1247 1258
rect 1251 1254 1303 1258
rect 1307 1254 1311 1258
rect 1315 1254 1367 1258
rect 1371 1254 1375 1258
rect 1379 1254 1431 1258
rect 1435 1254 1439 1258
rect 1443 1254 1503 1258
rect 1507 1254 1543 1258
rect 1547 1254 1583 1258
rect 1587 1254 1619 1258
rect 103 1253 1619 1254
rect 1625 1253 1626 1259
rect 84 1217 85 1223
rect 91 1222 1607 1223
rect 91 1218 111 1222
rect 115 1218 135 1222
rect 139 1218 143 1222
rect 147 1218 175 1222
rect 179 1218 215 1222
rect 219 1218 231 1222
rect 235 1218 263 1222
rect 267 1218 287 1222
rect 291 1218 311 1222
rect 315 1218 351 1222
rect 355 1218 359 1222
rect 363 1218 415 1222
rect 419 1218 471 1222
rect 475 1218 479 1222
rect 483 1218 527 1222
rect 531 1218 543 1222
rect 547 1218 583 1222
rect 587 1218 607 1222
rect 611 1218 639 1222
rect 643 1218 671 1222
rect 675 1218 687 1222
rect 691 1218 735 1222
rect 739 1218 783 1222
rect 787 1218 799 1222
rect 803 1218 831 1222
rect 835 1218 863 1222
rect 867 1218 879 1222
rect 883 1218 927 1222
rect 931 1218 935 1222
rect 939 1218 983 1222
rect 987 1218 991 1222
rect 995 1218 1039 1222
rect 1043 1218 1055 1222
rect 1059 1218 1095 1222
rect 1099 1218 1119 1222
rect 1123 1218 1159 1222
rect 1163 1218 1183 1222
rect 1187 1218 1231 1222
rect 1235 1218 1247 1222
rect 1251 1218 1303 1222
rect 1307 1218 1311 1222
rect 1315 1218 1375 1222
rect 1379 1218 1383 1222
rect 1387 1218 1439 1222
rect 1443 1218 1471 1222
rect 1475 1218 1503 1222
rect 1507 1218 1543 1222
rect 1547 1218 1583 1222
rect 1587 1218 1607 1222
rect 91 1217 1607 1218
rect 1613 1217 1614 1223
rect 96 1181 97 1187
rect 103 1186 1619 1187
rect 103 1182 111 1186
rect 115 1182 143 1186
rect 147 1182 175 1186
rect 179 1182 215 1186
rect 219 1182 255 1186
rect 259 1182 263 1186
rect 267 1182 303 1186
rect 307 1182 311 1186
rect 315 1182 359 1186
rect 363 1182 415 1186
rect 419 1182 471 1186
rect 475 1182 527 1186
rect 531 1182 583 1186
rect 587 1182 591 1186
rect 595 1182 639 1186
rect 643 1182 655 1186
rect 659 1182 687 1186
rect 691 1182 719 1186
rect 723 1182 735 1186
rect 739 1182 783 1186
rect 787 1182 791 1186
rect 795 1182 831 1186
rect 835 1182 855 1186
rect 859 1182 879 1186
rect 883 1182 919 1186
rect 923 1182 935 1186
rect 939 1182 983 1186
rect 987 1182 1039 1186
rect 1043 1182 1095 1186
rect 1099 1182 1103 1186
rect 1107 1182 1159 1186
rect 1163 1182 1167 1186
rect 1171 1182 1231 1186
rect 1235 1182 1239 1186
rect 1243 1182 1303 1186
rect 1307 1182 1311 1186
rect 1315 1182 1383 1186
rect 1387 1182 1391 1186
rect 1395 1182 1471 1186
rect 1475 1182 1479 1186
rect 1483 1182 1543 1186
rect 1547 1182 1583 1186
rect 1587 1182 1619 1186
rect 103 1181 1619 1182
rect 1625 1181 1626 1187
rect 84 1145 85 1151
rect 91 1150 1607 1151
rect 91 1146 111 1150
rect 115 1146 135 1150
rect 139 1146 143 1150
rect 147 1146 167 1150
rect 171 1146 175 1150
rect 179 1146 199 1150
rect 203 1146 215 1150
rect 219 1146 231 1150
rect 235 1146 255 1150
rect 259 1146 263 1150
rect 267 1146 295 1150
rect 299 1146 303 1150
rect 307 1146 327 1150
rect 331 1146 359 1150
rect 363 1146 391 1150
rect 395 1146 415 1150
rect 419 1146 447 1150
rect 451 1146 471 1150
rect 475 1146 503 1150
rect 507 1146 527 1150
rect 531 1146 559 1150
rect 563 1146 591 1150
rect 595 1146 615 1150
rect 619 1146 655 1150
rect 659 1146 671 1150
rect 675 1146 719 1150
rect 723 1146 727 1150
rect 731 1146 783 1150
rect 787 1146 791 1150
rect 795 1146 839 1150
rect 843 1146 855 1150
rect 859 1146 895 1150
rect 899 1146 919 1150
rect 923 1146 951 1150
rect 955 1146 983 1150
rect 987 1146 1007 1150
rect 1011 1146 1039 1150
rect 1043 1146 1063 1150
rect 1067 1146 1103 1150
rect 1107 1146 1127 1150
rect 1131 1146 1167 1150
rect 1171 1146 1191 1150
rect 1195 1146 1239 1150
rect 1243 1146 1255 1150
rect 1259 1146 1311 1150
rect 1315 1146 1327 1150
rect 1331 1146 1391 1150
rect 1395 1146 1399 1150
rect 1403 1146 1479 1150
rect 1483 1146 1543 1150
rect 1547 1146 1583 1150
rect 1587 1146 1607 1150
rect 91 1145 1607 1146
rect 1613 1145 1614 1151
rect 96 1109 97 1115
rect 103 1114 1619 1115
rect 103 1110 111 1114
rect 115 1110 135 1114
rect 139 1110 151 1114
rect 155 1110 167 1114
rect 171 1110 183 1114
rect 187 1110 199 1114
rect 203 1110 223 1114
rect 227 1110 231 1114
rect 235 1110 263 1114
rect 267 1110 271 1114
rect 275 1110 295 1114
rect 299 1110 327 1114
rect 331 1110 359 1114
rect 363 1110 383 1114
rect 387 1110 391 1114
rect 395 1110 439 1114
rect 443 1110 447 1114
rect 451 1110 503 1114
rect 507 1110 559 1114
rect 563 1110 567 1114
rect 571 1110 615 1114
rect 619 1110 639 1114
rect 643 1110 671 1114
rect 675 1110 711 1114
rect 715 1110 727 1114
rect 731 1110 783 1114
rect 787 1110 839 1114
rect 843 1110 855 1114
rect 859 1110 895 1114
rect 899 1110 919 1114
rect 923 1110 951 1114
rect 955 1110 983 1114
rect 987 1110 1007 1114
rect 1011 1110 1039 1114
rect 1043 1110 1063 1114
rect 1067 1110 1095 1114
rect 1099 1110 1127 1114
rect 1131 1110 1151 1114
rect 1155 1110 1191 1114
rect 1195 1110 1207 1114
rect 1211 1110 1255 1114
rect 1259 1110 1263 1114
rect 1267 1110 1319 1114
rect 1323 1110 1327 1114
rect 1331 1110 1375 1114
rect 1379 1110 1399 1114
rect 1403 1110 1439 1114
rect 1443 1110 1479 1114
rect 1483 1110 1503 1114
rect 1507 1110 1543 1114
rect 1547 1110 1583 1114
rect 1587 1110 1619 1114
rect 103 1109 1619 1110
rect 1625 1109 1626 1115
rect 166 1100 172 1101
rect 310 1100 316 1101
rect 166 1096 167 1100
rect 171 1096 311 1100
rect 315 1096 316 1100
rect 166 1095 172 1096
rect 310 1095 316 1096
rect 84 1065 85 1071
rect 91 1070 1607 1071
rect 91 1066 111 1070
rect 115 1066 151 1070
rect 155 1066 183 1070
rect 187 1066 223 1070
rect 227 1066 271 1070
rect 275 1066 327 1070
rect 331 1066 383 1070
rect 387 1066 439 1070
rect 443 1066 447 1070
rect 451 1066 487 1070
rect 491 1066 503 1070
rect 507 1066 543 1070
rect 547 1066 567 1070
rect 571 1066 599 1070
rect 603 1066 639 1070
rect 643 1066 663 1070
rect 667 1066 711 1070
rect 715 1066 727 1070
rect 731 1066 783 1070
rect 787 1066 791 1070
rect 795 1066 855 1070
rect 859 1066 863 1070
rect 867 1066 919 1070
rect 923 1066 935 1070
rect 939 1066 983 1070
rect 987 1066 1007 1070
rect 1011 1066 1039 1070
rect 1043 1066 1079 1070
rect 1083 1066 1095 1070
rect 1099 1066 1151 1070
rect 1155 1066 1207 1070
rect 1211 1066 1215 1070
rect 1219 1066 1263 1070
rect 1267 1066 1279 1070
rect 1283 1066 1319 1070
rect 1323 1066 1335 1070
rect 1339 1066 1375 1070
rect 1379 1066 1391 1070
rect 1395 1066 1439 1070
rect 1443 1066 1447 1070
rect 1451 1066 1503 1070
rect 1507 1066 1543 1070
rect 1547 1066 1583 1070
rect 1587 1066 1607 1070
rect 91 1065 1607 1066
rect 1613 1065 1614 1071
rect 96 1025 97 1031
rect 103 1030 1619 1031
rect 103 1026 111 1030
rect 115 1026 447 1030
rect 451 1026 487 1030
rect 491 1026 511 1030
rect 515 1026 543 1030
rect 547 1026 575 1030
rect 579 1026 599 1030
rect 603 1026 615 1030
rect 619 1026 663 1030
rect 667 1026 711 1030
rect 715 1026 727 1030
rect 731 1026 775 1030
rect 779 1026 791 1030
rect 795 1026 847 1030
rect 851 1026 863 1030
rect 867 1026 927 1030
rect 931 1026 935 1030
rect 939 1026 1007 1030
rect 1011 1026 1079 1030
rect 1083 1026 1087 1030
rect 1091 1026 1151 1030
rect 1155 1026 1167 1030
rect 1171 1026 1215 1030
rect 1219 1026 1239 1030
rect 1243 1026 1279 1030
rect 1283 1026 1303 1030
rect 1307 1026 1335 1030
rect 1339 1026 1359 1030
rect 1363 1026 1391 1030
rect 1395 1026 1407 1030
rect 1411 1026 1447 1030
rect 1451 1026 1455 1030
rect 1459 1026 1503 1030
rect 1507 1026 1511 1030
rect 1515 1026 1543 1030
rect 1547 1026 1583 1030
rect 1587 1026 1619 1030
rect 103 1025 1619 1026
rect 1625 1025 1626 1031
rect 84 981 85 987
rect 91 986 1607 987
rect 91 982 111 986
rect 115 982 159 986
rect 163 982 199 986
rect 203 982 255 986
rect 259 982 311 986
rect 315 982 375 986
rect 379 982 439 986
rect 443 982 503 986
rect 507 982 511 986
rect 515 982 543 986
rect 547 982 559 986
rect 563 982 575 986
rect 579 982 615 986
rect 619 982 663 986
rect 667 982 703 986
rect 707 982 711 986
rect 715 982 735 986
rect 739 982 775 986
rect 779 982 831 986
rect 835 982 847 986
rect 851 982 895 986
rect 899 982 927 986
rect 931 982 967 986
rect 971 982 1007 986
rect 1011 982 1047 986
rect 1051 982 1087 986
rect 1091 982 1127 986
rect 1131 982 1167 986
rect 1171 982 1199 986
rect 1203 982 1239 986
rect 1243 982 1271 986
rect 1275 982 1303 986
rect 1307 982 1343 986
rect 1347 982 1359 986
rect 1363 982 1407 986
rect 1411 982 1415 986
rect 1419 982 1455 986
rect 1459 982 1487 986
rect 1491 982 1511 986
rect 1515 982 1543 986
rect 1547 982 1583 986
rect 1587 982 1607 986
rect 91 981 1607 982
rect 1613 981 1614 987
rect 522 972 528 973
rect 586 972 592 973
rect 522 968 523 972
rect 527 968 587 972
rect 591 968 592 972
rect 522 967 528 968
rect 586 967 592 968
rect 96 945 97 951
rect 103 950 1619 951
rect 103 946 111 950
rect 115 946 151 950
rect 155 946 159 950
rect 163 946 191 950
rect 195 946 199 950
rect 203 946 247 950
rect 251 946 255 950
rect 259 946 303 950
rect 307 946 311 950
rect 315 946 367 950
rect 371 946 375 950
rect 379 946 431 950
rect 435 946 439 950
rect 443 946 495 950
rect 499 946 503 950
rect 507 946 559 950
rect 563 946 615 950
rect 619 946 663 950
rect 667 946 671 950
rect 675 946 703 950
rect 707 946 719 950
rect 723 946 735 950
rect 739 946 767 950
rect 771 946 775 950
rect 779 946 815 950
rect 819 946 831 950
rect 835 946 871 950
rect 875 946 895 950
rect 899 946 935 950
rect 939 946 967 950
rect 971 946 1007 950
rect 1011 946 1047 950
rect 1051 946 1079 950
rect 1083 946 1127 950
rect 1131 946 1143 950
rect 1147 946 1199 950
rect 1203 946 1207 950
rect 1211 946 1271 950
rect 1275 946 1327 950
rect 1331 946 1343 950
rect 1347 946 1375 950
rect 1379 946 1415 950
rect 1419 946 1423 950
rect 1427 946 1471 950
rect 1475 946 1487 950
rect 1491 946 1511 950
rect 1515 946 1543 950
rect 1547 946 1583 950
rect 1587 946 1619 950
rect 103 945 1619 946
rect 1625 945 1626 951
rect 84 905 85 911
rect 91 910 1607 911
rect 91 906 111 910
rect 115 906 135 910
rect 139 906 151 910
rect 155 906 167 910
rect 171 906 191 910
rect 195 906 223 910
rect 227 906 247 910
rect 251 906 279 910
rect 283 906 303 910
rect 307 906 335 910
rect 339 906 367 910
rect 371 906 391 910
rect 395 906 431 910
rect 435 906 447 910
rect 451 906 495 910
rect 499 906 503 910
rect 507 906 559 910
rect 563 906 615 910
rect 619 906 623 910
rect 627 906 671 910
rect 675 906 695 910
rect 699 906 719 910
rect 723 906 759 910
rect 763 906 767 910
rect 771 906 815 910
rect 819 906 823 910
rect 827 906 871 910
rect 875 906 887 910
rect 891 906 935 910
rect 939 906 951 910
rect 955 906 1007 910
rect 1011 906 1015 910
rect 1019 906 1079 910
rect 1083 906 1135 910
rect 1139 906 1143 910
rect 1147 906 1191 910
rect 1195 906 1207 910
rect 1211 906 1247 910
rect 1251 906 1271 910
rect 1275 906 1303 910
rect 1307 906 1327 910
rect 1331 906 1359 910
rect 1363 906 1375 910
rect 1379 906 1407 910
rect 1411 906 1423 910
rect 1427 906 1455 910
rect 1459 906 1471 910
rect 1475 906 1511 910
rect 1515 906 1543 910
rect 1547 906 1583 910
rect 1587 906 1607 910
rect 91 905 1607 906
rect 1613 905 1614 911
rect 96 869 97 875
rect 103 874 1619 875
rect 103 870 111 874
rect 115 870 135 874
rect 139 870 167 874
rect 171 870 207 874
rect 211 870 223 874
rect 227 870 255 874
rect 259 870 279 874
rect 283 870 303 874
rect 307 870 335 874
rect 339 870 343 874
rect 347 870 383 874
rect 387 870 391 874
rect 395 870 439 874
rect 443 870 447 874
rect 451 870 503 874
rect 507 870 511 874
rect 515 870 559 874
rect 563 870 591 874
rect 595 870 623 874
rect 627 870 679 874
rect 683 870 695 874
rect 699 870 759 874
rect 763 870 767 874
rect 771 870 823 874
rect 827 870 847 874
rect 851 870 887 874
rect 891 870 919 874
rect 923 870 951 874
rect 955 870 983 874
rect 987 870 1015 874
rect 1019 870 1039 874
rect 1043 870 1079 874
rect 1083 870 1095 874
rect 1099 870 1135 874
rect 1139 870 1151 874
rect 1155 870 1191 874
rect 1195 870 1207 874
rect 1211 870 1247 874
rect 1251 870 1263 874
rect 1267 870 1303 874
rect 1307 870 1327 874
rect 1331 870 1359 874
rect 1363 870 1399 874
rect 1403 870 1407 874
rect 1411 870 1455 874
rect 1459 870 1479 874
rect 1483 870 1511 874
rect 1515 870 1543 874
rect 1547 870 1583 874
rect 1587 870 1619 874
rect 103 869 1619 870
rect 1625 869 1626 875
rect 84 829 85 835
rect 91 834 1607 835
rect 91 830 111 834
rect 115 830 135 834
rect 139 830 167 834
rect 171 830 207 834
rect 211 830 223 834
rect 227 830 255 834
rect 259 830 287 834
rect 291 830 303 834
rect 307 830 343 834
rect 347 830 351 834
rect 355 830 383 834
rect 387 830 423 834
rect 427 830 439 834
rect 443 830 495 834
rect 499 830 511 834
rect 515 830 567 834
rect 571 830 591 834
rect 595 830 639 834
rect 643 830 679 834
rect 683 830 719 834
rect 723 830 767 834
rect 771 830 791 834
rect 795 830 847 834
rect 851 830 863 834
rect 867 830 919 834
rect 923 830 935 834
rect 939 830 983 834
rect 987 830 999 834
rect 1003 830 1039 834
rect 1043 830 1055 834
rect 1059 830 1095 834
rect 1099 830 1103 834
rect 1107 830 1143 834
rect 1147 830 1151 834
rect 1155 830 1183 834
rect 1187 830 1207 834
rect 1211 830 1231 834
rect 1235 830 1263 834
rect 1267 830 1279 834
rect 1283 830 1327 834
rect 1331 830 1399 834
rect 1403 830 1479 834
rect 1483 830 1543 834
rect 1547 830 1583 834
rect 1587 830 1607 834
rect 91 829 1607 830
rect 1613 829 1614 835
rect 96 793 97 799
rect 103 798 1619 799
rect 103 794 111 798
rect 115 794 135 798
rect 139 794 167 798
rect 171 794 199 798
rect 203 794 223 798
rect 227 794 247 798
rect 251 794 287 798
rect 291 794 303 798
rect 307 794 351 798
rect 355 794 359 798
rect 363 794 423 798
rect 427 794 487 798
rect 491 794 495 798
rect 499 794 551 798
rect 555 794 567 798
rect 571 794 607 798
rect 611 794 639 798
rect 643 794 671 798
rect 675 794 719 798
rect 723 794 735 798
rect 739 794 791 798
rect 795 794 799 798
rect 803 794 863 798
rect 867 794 871 798
rect 875 794 935 798
rect 939 794 999 798
rect 1003 794 1055 798
rect 1059 794 1063 798
rect 1067 794 1103 798
rect 1107 794 1127 798
rect 1131 794 1143 798
rect 1147 794 1183 798
rect 1187 794 1191 798
rect 1195 794 1231 798
rect 1235 794 1255 798
rect 1259 794 1279 798
rect 1283 794 1319 798
rect 1323 794 1327 798
rect 1331 794 1383 798
rect 1387 794 1583 798
rect 1587 794 1619 798
rect 103 793 1619 794
rect 1625 793 1626 799
rect 84 757 85 763
rect 91 762 1607 763
rect 91 758 111 762
rect 115 758 135 762
rect 139 758 167 762
rect 171 758 199 762
rect 203 758 247 762
rect 251 758 255 762
rect 259 758 303 762
rect 307 758 319 762
rect 323 758 359 762
rect 363 758 391 762
rect 395 758 423 762
rect 427 758 463 762
rect 467 758 487 762
rect 491 758 543 762
rect 547 758 551 762
rect 555 758 607 762
rect 611 758 623 762
rect 627 758 671 762
rect 675 758 703 762
rect 707 758 735 762
rect 739 758 775 762
rect 779 758 799 762
rect 803 758 847 762
rect 851 758 871 762
rect 875 758 919 762
rect 923 758 935 762
rect 939 758 991 762
rect 995 758 999 762
rect 1003 758 1063 762
rect 1067 758 1127 762
rect 1131 758 1135 762
rect 1139 758 1191 762
rect 1195 758 1207 762
rect 1211 758 1255 762
rect 1259 758 1271 762
rect 1275 758 1319 762
rect 1323 758 1327 762
rect 1331 758 1375 762
rect 1379 758 1383 762
rect 1387 758 1423 762
rect 1427 758 1471 762
rect 1475 758 1511 762
rect 1515 758 1543 762
rect 1547 758 1583 762
rect 1587 758 1607 762
rect 91 757 1607 758
rect 1613 757 1614 763
rect 96 721 97 727
rect 103 726 1619 727
rect 103 722 111 726
rect 115 722 135 726
rect 139 722 167 726
rect 171 722 199 726
rect 203 722 207 726
rect 211 722 255 726
rect 259 722 311 726
rect 315 722 319 726
rect 323 722 367 726
rect 371 722 391 726
rect 395 722 423 726
rect 427 722 463 726
rect 467 722 479 726
rect 483 722 543 726
rect 547 722 615 726
rect 619 722 623 726
rect 627 722 687 726
rect 691 722 703 726
rect 707 722 759 726
rect 763 722 775 726
rect 779 722 839 726
rect 843 722 847 726
rect 851 722 919 726
rect 923 722 991 726
rect 995 722 1007 726
rect 1011 722 1063 726
rect 1067 722 1087 726
rect 1091 722 1135 726
rect 1139 722 1167 726
rect 1171 722 1207 726
rect 1211 722 1239 726
rect 1243 722 1271 726
rect 1275 722 1303 726
rect 1307 722 1327 726
rect 1331 722 1359 726
rect 1363 722 1375 726
rect 1379 722 1407 726
rect 1411 722 1423 726
rect 1427 722 1455 726
rect 1459 722 1471 726
rect 1475 722 1511 726
rect 1515 722 1543 726
rect 1547 722 1583 726
rect 1587 722 1619 726
rect 103 721 1619 722
rect 1625 721 1626 727
rect 84 685 85 691
rect 91 690 1607 691
rect 91 686 111 690
rect 115 686 135 690
rect 139 686 159 690
rect 163 686 167 690
rect 171 686 207 690
rect 211 686 255 690
rect 259 686 303 690
rect 307 686 311 690
rect 315 686 359 690
rect 363 686 367 690
rect 371 686 415 690
rect 419 686 423 690
rect 427 686 471 690
rect 475 686 479 690
rect 483 686 527 690
rect 531 686 543 690
rect 547 686 583 690
rect 587 686 615 690
rect 619 686 639 690
rect 643 686 687 690
rect 691 686 695 690
rect 699 686 759 690
rect 763 686 823 690
rect 827 686 839 690
rect 843 686 887 690
rect 891 686 919 690
rect 923 686 951 690
rect 955 686 1007 690
rect 1011 686 1015 690
rect 1019 686 1079 690
rect 1083 686 1087 690
rect 1091 686 1135 690
rect 1139 686 1167 690
rect 1171 686 1191 690
rect 1195 686 1239 690
rect 1243 686 1247 690
rect 1251 686 1303 690
rect 1307 686 1359 690
rect 1363 686 1407 690
rect 1411 686 1455 690
rect 1459 686 1511 690
rect 1515 686 1543 690
rect 1547 686 1583 690
rect 1587 686 1607 690
rect 91 685 1607 686
rect 1613 685 1614 691
rect 96 645 97 651
rect 103 650 1619 651
rect 103 646 111 650
rect 115 646 159 650
rect 163 646 167 650
rect 171 646 207 650
rect 211 646 215 650
rect 219 646 255 650
rect 259 646 271 650
rect 275 646 303 650
rect 307 646 327 650
rect 331 646 359 650
rect 363 646 383 650
rect 387 646 415 650
rect 419 646 431 650
rect 435 646 471 650
rect 475 646 487 650
rect 491 646 527 650
rect 531 646 535 650
rect 539 646 583 650
rect 587 646 591 650
rect 595 646 639 650
rect 643 646 647 650
rect 651 646 695 650
rect 699 646 703 650
rect 707 646 759 650
rect 763 646 823 650
rect 827 646 887 650
rect 891 646 943 650
rect 947 646 951 650
rect 955 646 999 650
rect 1003 646 1015 650
rect 1019 646 1055 650
rect 1059 646 1079 650
rect 1083 646 1111 650
rect 1115 646 1135 650
rect 1139 646 1167 650
rect 1171 646 1191 650
rect 1195 646 1215 650
rect 1219 646 1247 650
rect 1251 646 1271 650
rect 1275 646 1303 650
rect 1307 646 1327 650
rect 1331 646 1359 650
rect 1363 646 1383 650
rect 1387 646 1439 650
rect 1443 646 1503 650
rect 1507 646 1543 650
rect 1547 646 1583 650
rect 1587 646 1619 650
rect 103 645 1619 646
rect 1625 645 1626 651
rect 84 609 85 615
rect 91 614 1607 615
rect 91 610 111 614
rect 115 610 167 614
rect 171 610 215 614
rect 219 610 223 614
rect 227 610 255 614
rect 259 610 271 614
rect 275 610 287 614
rect 291 610 319 614
rect 323 610 327 614
rect 331 610 351 614
rect 355 610 383 614
rect 387 610 423 614
rect 427 610 431 614
rect 435 610 463 614
rect 467 610 487 614
rect 491 610 519 614
rect 523 610 535 614
rect 539 610 583 614
rect 587 610 591 614
rect 595 610 647 614
rect 651 610 703 614
rect 707 610 719 614
rect 723 610 759 614
rect 763 610 799 614
rect 803 610 823 614
rect 827 610 887 614
rect 891 610 943 614
rect 947 610 975 614
rect 979 610 999 614
rect 1003 610 1055 614
rect 1059 610 1063 614
rect 1067 610 1111 614
rect 1115 610 1143 614
rect 1147 610 1167 614
rect 1171 610 1215 614
rect 1219 610 1271 614
rect 1275 610 1287 614
rect 1291 610 1327 614
rect 1331 610 1351 614
rect 1355 610 1383 614
rect 1387 610 1407 614
rect 1411 610 1439 614
rect 1443 610 1455 614
rect 1459 610 1503 614
rect 1507 610 1511 614
rect 1515 610 1543 614
rect 1547 610 1583 614
rect 1587 610 1607 614
rect 91 609 1607 610
rect 1613 609 1614 615
rect 96 573 97 579
rect 103 578 1619 579
rect 103 574 111 578
rect 115 574 191 578
rect 195 574 223 578
rect 227 574 255 578
rect 259 574 287 578
rect 291 574 319 578
rect 323 574 327 578
rect 331 574 351 578
rect 355 574 383 578
rect 387 574 399 578
rect 403 574 423 578
rect 427 574 463 578
rect 467 574 471 578
rect 475 574 519 578
rect 523 574 535 578
rect 539 574 583 578
rect 587 574 599 578
rect 603 574 647 578
rect 651 574 663 578
rect 667 574 719 578
rect 723 574 727 578
rect 731 574 783 578
rect 787 574 799 578
rect 803 574 839 578
rect 843 574 887 578
rect 891 574 903 578
rect 907 574 967 578
rect 971 574 975 578
rect 979 574 1039 578
rect 1043 574 1063 578
rect 1067 574 1103 578
rect 1107 574 1143 578
rect 1147 574 1167 578
rect 1171 574 1215 578
rect 1219 574 1231 578
rect 1235 574 1287 578
rect 1291 574 1335 578
rect 1339 574 1351 578
rect 1355 574 1383 578
rect 1387 574 1407 578
rect 1411 574 1423 578
rect 1427 574 1455 578
rect 1459 574 1471 578
rect 1475 574 1511 578
rect 1515 574 1543 578
rect 1547 574 1583 578
rect 1587 574 1619 578
rect 103 573 1619 574
rect 1625 573 1626 579
rect 84 537 85 543
rect 91 542 1607 543
rect 91 538 111 542
rect 115 538 135 542
rect 139 538 175 542
rect 179 538 191 542
rect 195 538 231 542
rect 235 538 255 542
rect 259 538 295 542
rect 299 538 327 542
rect 331 538 359 542
rect 363 538 399 542
rect 403 538 423 542
rect 427 538 471 542
rect 475 538 479 542
rect 483 538 535 542
rect 539 538 543 542
rect 547 538 599 542
rect 603 538 655 542
rect 659 538 663 542
rect 667 538 711 542
rect 715 538 727 542
rect 731 538 767 542
rect 771 538 783 542
rect 787 538 831 542
rect 835 538 839 542
rect 843 538 895 542
rect 899 538 903 542
rect 907 538 967 542
rect 971 538 1031 542
rect 1035 538 1039 542
rect 1043 538 1095 542
rect 1099 538 1103 542
rect 1107 538 1167 542
rect 1171 538 1231 542
rect 1235 538 1239 542
rect 1243 538 1287 542
rect 1291 538 1311 542
rect 1315 538 1335 542
rect 1339 538 1383 542
rect 1387 538 1391 542
rect 1395 538 1423 542
rect 1427 538 1471 542
rect 1475 538 1479 542
rect 1483 538 1511 542
rect 1515 538 1543 542
rect 1547 538 1583 542
rect 1587 538 1607 542
rect 91 537 1607 538
rect 1613 537 1614 543
rect 96 501 97 507
rect 103 506 1619 507
rect 103 502 111 506
rect 115 502 135 506
rect 139 502 167 506
rect 171 502 175 506
rect 179 502 199 506
rect 203 502 231 506
rect 235 502 247 506
rect 251 502 295 506
rect 299 502 343 506
rect 347 502 359 506
rect 363 502 399 506
rect 403 502 423 506
rect 427 502 455 506
rect 459 502 479 506
rect 483 502 511 506
rect 515 502 543 506
rect 547 502 567 506
rect 571 502 599 506
rect 603 502 623 506
rect 627 502 655 506
rect 659 502 679 506
rect 683 502 711 506
rect 715 502 743 506
rect 747 502 767 506
rect 771 502 815 506
rect 819 502 831 506
rect 835 502 887 506
rect 891 502 895 506
rect 899 502 959 506
rect 963 502 967 506
rect 971 502 1031 506
rect 1035 502 1039 506
rect 1043 502 1095 506
rect 1099 502 1127 506
rect 1131 502 1167 506
rect 1171 502 1223 506
rect 1227 502 1239 506
rect 1243 502 1311 506
rect 1315 502 1327 506
rect 1331 502 1391 506
rect 1395 502 1439 506
rect 1443 502 1479 506
rect 1483 502 1543 506
rect 1547 502 1583 506
rect 1587 502 1619 506
rect 103 501 1619 502
rect 1625 501 1626 507
rect 84 465 85 471
rect 91 470 1607 471
rect 91 466 111 470
rect 115 466 135 470
rect 139 466 167 470
rect 171 466 199 470
rect 203 466 247 470
rect 251 466 255 470
rect 259 466 295 470
rect 299 466 311 470
rect 315 466 343 470
rect 347 466 367 470
rect 371 466 399 470
rect 403 466 423 470
rect 427 466 455 470
rect 459 466 479 470
rect 483 466 511 470
rect 515 466 535 470
rect 539 466 567 470
rect 571 466 599 470
rect 603 466 623 470
rect 627 466 663 470
rect 667 466 679 470
rect 683 466 735 470
rect 739 466 743 470
rect 747 466 807 470
rect 811 466 815 470
rect 819 466 871 470
rect 875 466 887 470
rect 891 466 935 470
rect 939 466 959 470
rect 963 466 991 470
rect 995 466 1039 470
rect 1043 466 1047 470
rect 1051 466 1095 470
rect 1099 466 1127 470
rect 1131 466 1143 470
rect 1147 466 1199 470
rect 1203 466 1223 470
rect 1227 466 1263 470
rect 1267 466 1327 470
rect 1331 466 1399 470
rect 1403 466 1439 470
rect 1443 466 1479 470
rect 1483 466 1543 470
rect 1547 466 1583 470
rect 1587 466 1607 470
rect 91 465 1607 466
rect 1613 465 1614 471
rect 96 425 97 431
rect 103 430 1619 431
rect 103 426 111 430
rect 115 426 135 430
rect 139 426 167 430
rect 171 426 199 430
rect 203 426 231 430
rect 235 426 255 430
rect 259 426 295 430
rect 299 426 311 430
rect 315 426 359 430
rect 363 426 367 430
rect 371 426 423 430
rect 427 426 479 430
rect 483 426 487 430
rect 491 426 535 430
rect 539 426 543 430
rect 547 426 591 430
rect 595 426 599 430
rect 603 426 639 430
rect 643 426 663 430
rect 667 426 679 430
rect 683 426 719 430
rect 723 426 735 430
rect 739 426 759 430
rect 763 426 807 430
rect 811 426 863 430
rect 867 426 871 430
rect 875 426 919 430
rect 923 426 935 430
rect 939 426 975 430
rect 979 426 991 430
rect 995 426 1031 430
rect 1035 426 1047 430
rect 1051 426 1087 430
rect 1091 426 1095 430
rect 1099 426 1143 430
rect 1147 426 1151 430
rect 1155 426 1199 430
rect 1203 426 1223 430
rect 1227 426 1263 430
rect 1267 426 1303 430
rect 1307 426 1327 430
rect 1331 426 1383 430
rect 1387 426 1399 430
rect 1403 426 1471 430
rect 1475 426 1479 430
rect 1483 426 1543 430
rect 1547 426 1583 430
rect 1587 426 1619 430
rect 103 425 1619 426
rect 1625 425 1626 431
rect 84 389 85 395
rect 91 394 1607 395
rect 91 390 111 394
rect 115 390 135 394
rect 139 390 167 394
rect 171 390 207 394
rect 211 390 231 394
rect 235 390 295 394
rect 299 390 359 394
rect 363 390 383 394
rect 387 390 423 394
rect 427 390 463 394
rect 467 390 487 394
rect 491 390 535 394
rect 539 390 543 394
rect 547 390 591 394
rect 595 390 599 394
rect 603 390 639 394
rect 643 390 655 394
rect 659 390 679 394
rect 683 390 703 394
rect 707 390 719 394
rect 723 390 751 394
rect 755 390 759 394
rect 763 390 807 394
rect 811 390 863 394
rect 867 390 919 394
rect 923 390 975 394
rect 979 390 983 394
rect 987 390 1031 394
rect 1035 390 1055 394
rect 1059 390 1087 394
rect 1091 390 1127 394
rect 1131 390 1151 394
rect 1155 390 1199 394
rect 1203 390 1223 394
rect 1227 390 1271 394
rect 1275 390 1303 394
rect 1307 390 1343 394
rect 1347 390 1383 394
rect 1387 390 1415 394
rect 1419 390 1471 394
rect 1475 390 1487 394
rect 1491 390 1543 394
rect 1547 390 1583 394
rect 1587 390 1607 394
rect 91 389 1607 390
rect 1613 389 1614 395
rect 96 353 97 359
rect 103 358 1619 359
rect 103 354 111 358
rect 115 354 135 358
rect 139 354 175 358
rect 179 354 207 358
rect 211 354 223 358
rect 227 354 279 358
rect 283 354 295 358
rect 299 354 335 358
rect 339 354 383 358
rect 387 354 391 358
rect 395 354 447 358
rect 451 354 463 358
rect 467 354 503 358
rect 507 354 535 358
rect 539 354 567 358
rect 571 354 599 358
rect 603 354 631 358
rect 635 354 655 358
rect 659 354 687 358
rect 691 354 703 358
rect 707 354 751 358
rect 755 354 807 358
rect 811 354 815 358
rect 819 354 863 358
rect 867 354 879 358
rect 883 354 919 358
rect 923 354 951 358
rect 955 354 983 358
rect 987 354 1031 358
rect 1035 354 1055 358
rect 1059 354 1103 358
rect 1107 354 1127 358
rect 1131 354 1175 358
rect 1179 354 1199 358
rect 1203 354 1247 358
rect 1251 354 1271 358
rect 1275 354 1327 358
rect 1331 354 1343 358
rect 1347 354 1407 358
rect 1411 354 1415 358
rect 1419 354 1487 358
rect 1491 354 1543 358
rect 1547 354 1583 358
rect 1587 354 1619 358
rect 103 353 1619 354
rect 1625 353 1626 359
rect 84 317 85 323
rect 91 322 1607 323
rect 91 318 111 322
rect 115 318 135 322
rect 139 318 175 322
rect 179 318 191 322
rect 195 318 223 322
rect 227 318 255 322
rect 259 318 279 322
rect 283 318 295 322
rect 299 318 335 322
rect 339 318 367 322
rect 371 318 391 322
rect 395 318 407 322
rect 411 318 447 322
rect 451 318 455 322
rect 459 318 503 322
rect 507 318 519 322
rect 523 318 567 322
rect 571 318 591 322
rect 595 318 631 322
rect 635 318 663 322
rect 667 318 687 322
rect 691 318 735 322
rect 739 318 751 322
rect 755 318 807 322
rect 811 318 815 322
rect 819 318 879 322
rect 883 318 951 322
rect 955 318 1023 322
rect 1027 318 1031 322
rect 1035 318 1095 322
rect 1099 318 1103 322
rect 1107 318 1167 322
rect 1171 318 1175 322
rect 1179 318 1231 322
rect 1235 318 1247 322
rect 1251 318 1295 322
rect 1299 318 1327 322
rect 1331 318 1351 322
rect 1355 318 1399 322
rect 1403 318 1407 322
rect 1411 318 1455 322
rect 1459 318 1487 322
rect 1491 318 1511 322
rect 1515 318 1543 322
rect 1547 318 1583 322
rect 1587 318 1607 322
rect 91 317 1607 318
rect 1613 317 1614 323
rect 96 277 97 283
rect 103 282 1619 283
rect 103 278 111 282
rect 115 278 151 282
rect 155 278 183 282
rect 187 278 191 282
rect 195 278 215 282
rect 219 278 223 282
rect 227 278 247 282
rect 251 278 255 282
rect 259 278 279 282
rect 283 278 295 282
rect 299 278 311 282
rect 315 278 335 282
rect 339 278 351 282
rect 355 278 367 282
rect 371 278 407 282
rect 411 278 455 282
rect 459 278 479 282
rect 483 278 519 282
rect 523 278 559 282
rect 563 278 591 282
rect 595 278 647 282
rect 651 278 663 282
rect 667 278 735 282
rect 739 278 807 282
rect 811 278 823 282
rect 827 278 879 282
rect 883 278 903 282
rect 907 278 951 282
rect 955 278 983 282
rect 987 278 1023 282
rect 1027 278 1055 282
rect 1059 278 1095 282
rect 1099 278 1119 282
rect 1123 278 1167 282
rect 1171 278 1175 282
rect 1179 278 1223 282
rect 1227 278 1231 282
rect 1235 278 1263 282
rect 1267 278 1295 282
rect 1299 278 1303 282
rect 1307 278 1351 282
rect 1355 278 1399 282
rect 1403 278 1447 282
rect 1451 278 1455 282
rect 1459 278 1503 282
rect 1507 278 1511 282
rect 1515 278 1543 282
rect 1547 278 1583 282
rect 1587 278 1619 282
rect 103 277 1619 278
rect 1625 277 1626 283
rect 84 241 85 247
rect 91 246 1607 247
rect 91 242 111 246
rect 115 242 135 246
rect 139 242 151 246
rect 155 242 167 246
rect 171 242 183 246
rect 187 242 207 246
rect 211 242 215 246
rect 219 242 247 246
rect 251 242 255 246
rect 259 242 279 246
rect 283 242 303 246
rect 307 242 311 246
rect 315 242 343 246
rect 347 242 351 246
rect 355 242 383 246
rect 387 242 407 246
rect 411 242 439 246
rect 443 242 479 246
rect 483 242 511 246
rect 515 242 559 246
rect 563 242 591 246
rect 595 242 647 246
rect 651 242 679 246
rect 683 242 735 246
rect 739 242 767 246
rect 771 242 823 246
rect 827 242 847 246
rect 851 242 903 246
rect 907 242 919 246
rect 923 242 983 246
rect 987 242 1047 246
rect 1051 242 1055 246
rect 1059 242 1103 246
rect 1107 242 1119 246
rect 1123 242 1159 246
rect 1163 242 1175 246
rect 1179 242 1215 246
rect 1219 242 1223 246
rect 1227 242 1263 246
rect 1267 242 1271 246
rect 1275 242 1303 246
rect 1307 242 1327 246
rect 1331 242 1351 246
rect 1355 242 1383 246
rect 1387 242 1399 246
rect 1403 242 1439 246
rect 1443 242 1447 246
rect 1451 242 1503 246
rect 1507 242 1543 246
rect 1547 242 1583 246
rect 1587 242 1607 246
rect 91 241 1607 242
rect 1613 241 1614 247
rect 96 201 97 207
rect 103 206 1619 207
rect 103 202 111 206
rect 115 202 135 206
rect 139 202 167 206
rect 171 202 207 206
rect 211 202 215 206
rect 219 202 255 206
rect 259 202 263 206
rect 267 202 303 206
rect 307 202 311 206
rect 315 202 343 206
rect 347 202 359 206
rect 363 202 383 206
rect 387 202 415 206
rect 419 202 439 206
rect 443 202 471 206
rect 475 202 511 206
rect 515 202 535 206
rect 539 202 591 206
rect 595 202 607 206
rect 611 202 679 206
rect 683 202 751 206
rect 755 202 767 206
rect 771 202 815 206
rect 819 202 847 206
rect 851 202 879 206
rect 883 202 919 206
rect 923 202 943 206
rect 947 202 983 206
rect 987 202 1007 206
rect 1011 202 1047 206
rect 1051 202 1063 206
rect 1067 202 1103 206
rect 1107 202 1119 206
rect 1123 202 1159 206
rect 1163 202 1175 206
rect 1179 202 1215 206
rect 1219 202 1231 206
rect 1235 202 1271 206
rect 1275 202 1287 206
rect 1291 202 1327 206
rect 1331 202 1343 206
rect 1347 202 1383 206
rect 1387 202 1399 206
rect 1403 202 1439 206
rect 1443 202 1455 206
rect 1459 202 1503 206
rect 1507 202 1511 206
rect 1515 202 1543 206
rect 1547 202 1583 206
rect 1587 202 1619 206
rect 103 201 1619 202
rect 1625 201 1626 207
rect 84 165 85 171
rect 91 170 1607 171
rect 91 166 111 170
rect 115 166 135 170
rect 139 166 143 170
rect 147 166 167 170
rect 171 166 191 170
rect 195 166 215 170
rect 219 166 239 170
rect 243 166 263 170
rect 267 166 295 170
rect 299 166 311 170
rect 315 166 351 170
rect 355 166 359 170
rect 363 166 407 170
rect 411 166 415 170
rect 419 166 463 170
rect 467 166 471 170
rect 475 166 519 170
rect 523 166 535 170
rect 539 166 575 170
rect 579 166 607 170
rect 611 166 631 170
rect 635 166 679 170
rect 683 166 687 170
rect 691 166 743 170
rect 747 166 751 170
rect 755 166 799 170
rect 803 166 815 170
rect 819 166 855 170
rect 859 166 879 170
rect 883 166 911 170
rect 915 166 943 170
rect 947 166 975 170
rect 979 166 1007 170
rect 1011 166 1039 170
rect 1043 166 1063 170
rect 1067 166 1095 170
rect 1099 166 1119 170
rect 1123 166 1151 170
rect 1155 166 1175 170
rect 1179 166 1207 170
rect 1211 166 1231 170
rect 1235 166 1255 170
rect 1259 166 1287 170
rect 1291 166 1303 170
rect 1307 166 1343 170
rect 1347 166 1351 170
rect 1355 166 1399 170
rect 1403 166 1455 170
rect 1459 166 1511 170
rect 1515 166 1543 170
rect 1547 166 1583 170
rect 1587 166 1607 170
rect 91 165 1607 166
rect 1613 165 1614 171
rect 96 117 97 123
rect 103 122 1619 123
rect 103 118 111 122
rect 115 118 135 122
rect 139 118 143 122
rect 147 118 167 122
rect 171 118 191 122
rect 195 118 199 122
rect 203 118 231 122
rect 235 118 239 122
rect 243 118 263 122
rect 267 118 295 122
rect 299 118 327 122
rect 331 118 351 122
rect 355 118 359 122
rect 363 118 391 122
rect 395 118 407 122
rect 411 118 423 122
rect 427 118 455 122
rect 459 118 463 122
rect 467 118 487 122
rect 491 118 519 122
rect 523 118 551 122
rect 555 118 575 122
rect 579 118 583 122
rect 587 118 615 122
rect 619 118 631 122
rect 635 118 647 122
rect 651 118 679 122
rect 683 118 687 122
rect 691 118 711 122
rect 715 118 743 122
rect 747 118 775 122
rect 779 118 799 122
rect 803 118 807 122
rect 811 118 839 122
rect 843 118 855 122
rect 859 118 871 122
rect 875 118 903 122
rect 907 118 911 122
rect 915 118 943 122
rect 947 118 975 122
rect 979 118 983 122
rect 987 118 1031 122
rect 1035 118 1039 122
rect 1043 118 1079 122
rect 1083 118 1095 122
rect 1099 118 1127 122
rect 1131 118 1151 122
rect 1155 118 1175 122
rect 1179 118 1207 122
rect 1211 118 1223 122
rect 1227 118 1255 122
rect 1259 118 1263 122
rect 1267 118 1303 122
rect 1307 118 1343 122
rect 1347 118 1351 122
rect 1355 118 1383 122
rect 1387 118 1399 122
rect 1403 118 1423 122
rect 1427 118 1455 122
rect 1459 118 1471 122
rect 1475 118 1511 122
rect 1515 118 1543 122
rect 1547 118 1583 122
rect 1587 118 1619 122
rect 103 117 1619 118
rect 1625 117 1626 123
rect 84 81 85 87
rect 91 86 1607 87
rect 91 82 111 86
rect 115 82 135 86
rect 139 82 167 86
rect 171 82 199 86
rect 203 82 231 86
rect 235 82 263 86
rect 267 82 295 86
rect 299 82 327 86
rect 331 82 359 86
rect 363 82 391 86
rect 395 82 423 86
rect 427 82 455 86
rect 459 82 487 86
rect 491 82 519 86
rect 523 82 551 86
rect 555 82 583 86
rect 587 82 615 86
rect 619 82 647 86
rect 651 82 679 86
rect 683 82 711 86
rect 715 82 743 86
rect 747 82 775 86
rect 779 82 807 86
rect 811 82 839 86
rect 843 82 871 86
rect 875 82 903 86
rect 907 82 943 86
rect 947 82 983 86
rect 987 82 1031 86
rect 1035 82 1079 86
rect 1083 82 1127 86
rect 1131 82 1175 86
rect 1179 82 1223 86
rect 1227 82 1263 86
rect 1267 82 1303 86
rect 1307 82 1343 86
rect 1347 82 1383 86
rect 1387 82 1423 86
rect 1427 82 1471 86
rect 1475 82 1511 86
rect 1515 82 1543 86
rect 1547 82 1583 86
rect 1587 82 1607 86
rect 91 81 1607 82
rect 1613 81 1614 87
<< m5c >>
rect 85 1649 91 1655
rect 1607 1649 1613 1655
rect 97 1613 103 1619
rect 1619 1613 1625 1619
rect 85 1577 91 1583
rect 1607 1577 1613 1583
rect 97 1541 103 1547
rect 1619 1541 1625 1547
rect 85 1505 91 1511
rect 1607 1505 1613 1511
rect 97 1469 103 1475
rect 1619 1469 1625 1475
rect 85 1433 91 1439
rect 1607 1433 1613 1439
rect 97 1397 103 1403
rect 1619 1397 1625 1403
rect 85 1361 91 1367
rect 1607 1361 1613 1367
rect 97 1325 103 1331
rect 1619 1325 1625 1331
rect 85 1289 91 1295
rect 1607 1289 1613 1295
rect 97 1253 103 1259
rect 1619 1253 1625 1259
rect 85 1217 91 1223
rect 1607 1217 1613 1223
rect 97 1181 103 1187
rect 1619 1181 1625 1187
rect 85 1145 91 1151
rect 1607 1145 1613 1151
rect 97 1109 103 1115
rect 1619 1109 1625 1115
rect 85 1065 91 1071
rect 1607 1065 1613 1071
rect 97 1025 103 1031
rect 1619 1025 1625 1031
rect 85 981 91 987
rect 1607 981 1613 987
rect 97 945 103 951
rect 1619 945 1625 951
rect 85 905 91 911
rect 1607 905 1613 911
rect 97 869 103 875
rect 1619 869 1625 875
rect 85 829 91 835
rect 1607 829 1613 835
rect 97 793 103 799
rect 1619 793 1625 799
rect 85 757 91 763
rect 1607 757 1613 763
rect 97 721 103 727
rect 1619 721 1625 727
rect 85 685 91 691
rect 1607 685 1613 691
rect 97 645 103 651
rect 1619 645 1625 651
rect 85 609 91 615
rect 1607 609 1613 615
rect 97 573 103 579
rect 1619 573 1625 579
rect 85 537 91 543
rect 1607 537 1613 543
rect 97 501 103 507
rect 1619 501 1625 507
rect 85 465 91 471
rect 1607 465 1613 471
rect 97 425 103 431
rect 1619 425 1625 431
rect 85 389 91 395
rect 1607 389 1613 395
rect 97 353 103 359
rect 1619 353 1625 359
rect 85 317 91 323
rect 1607 317 1613 323
rect 97 277 103 283
rect 1619 277 1625 283
rect 85 241 91 247
rect 1607 241 1613 247
rect 97 201 103 207
rect 1619 201 1625 207
rect 85 165 91 171
rect 1607 165 1613 171
rect 97 117 103 123
rect 1619 117 1625 123
rect 85 81 91 87
rect 1607 81 1613 87
<< m5 >>
rect 84 1655 92 1656
rect 84 1649 85 1655
rect 91 1649 92 1655
rect 84 1583 92 1649
rect 84 1577 85 1583
rect 91 1577 92 1583
rect 84 1511 92 1577
rect 84 1505 85 1511
rect 91 1505 92 1511
rect 84 1439 92 1505
rect 84 1433 85 1439
rect 91 1433 92 1439
rect 84 1367 92 1433
rect 84 1361 85 1367
rect 91 1361 92 1367
rect 84 1295 92 1361
rect 84 1289 85 1295
rect 91 1289 92 1295
rect 84 1223 92 1289
rect 84 1217 85 1223
rect 91 1217 92 1223
rect 84 1151 92 1217
rect 84 1145 85 1151
rect 91 1145 92 1151
rect 84 1071 92 1145
rect 84 1065 85 1071
rect 91 1065 92 1071
rect 84 987 92 1065
rect 84 981 85 987
rect 91 981 92 987
rect 84 911 92 981
rect 84 905 85 911
rect 91 905 92 911
rect 84 835 92 905
rect 84 829 85 835
rect 91 829 92 835
rect 84 763 92 829
rect 84 757 85 763
rect 91 757 92 763
rect 84 691 92 757
rect 84 685 85 691
rect 91 685 92 691
rect 84 615 92 685
rect 84 609 85 615
rect 91 609 92 615
rect 84 543 92 609
rect 84 537 85 543
rect 91 537 92 543
rect 84 471 92 537
rect 84 465 85 471
rect 91 465 92 471
rect 84 395 92 465
rect 84 389 85 395
rect 91 389 92 395
rect 84 323 92 389
rect 84 317 85 323
rect 91 317 92 323
rect 84 247 92 317
rect 84 241 85 247
rect 91 241 92 247
rect 84 171 92 241
rect 84 165 85 171
rect 91 165 92 171
rect 84 87 92 165
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 1619 104 1656
rect 96 1613 97 1619
rect 103 1613 104 1619
rect 96 1547 104 1613
rect 96 1541 97 1547
rect 103 1541 104 1547
rect 96 1475 104 1541
rect 96 1469 97 1475
rect 103 1469 104 1475
rect 96 1403 104 1469
rect 96 1397 97 1403
rect 103 1397 104 1403
rect 96 1331 104 1397
rect 96 1325 97 1331
rect 103 1325 104 1331
rect 96 1259 104 1325
rect 96 1253 97 1259
rect 103 1253 104 1259
rect 96 1187 104 1253
rect 96 1181 97 1187
rect 103 1181 104 1187
rect 96 1115 104 1181
rect 96 1109 97 1115
rect 103 1109 104 1115
rect 96 1031 104 1109
rect 96 1025 97 1031
rect 103 1025 104 1031
rect 96 951 104 1025
rect 96 945 97 951
rect 103 945 104 951
rect 96 875 104 945
rect 96 869 97 875
rect 103 869 104 875
rect 96 799 104 869
rect 96 793 97 799
rect 103 793 104 799
rect 96 727 104 793
rect 96 721 97 727
rect 103 721 104 727
rect 96 651 104 721
rect 96 645 97 651
rect 103 645 104 651
rect 96 579 104 645
rect 96 573 97 579
rect 103 573 104 579
rect 96 507 104 573
rect 96 501 97 507
rect 103 501 104 507
rect 96 431 104 501
rect 96 425 97 431
rect 103 425 104 431
rect 96 359 104 425
rect 96 353 97 359
rect 103 353 104 359
rect 96 283 104 353
rect 96 277 97 283
rect 103 277 104 283
rect 96 207 104 277
rect 96 201 97 207
rect 103 201 104 207
rect 96 123 104 201
rect 96 117 97 123
rect 103 117 104 123
rect 96 72 104 117
rect 1606 1655 1614 1656
rect 1606 1649 1607 1655
rect 1613 1649 1614 1655
rect 1606 1583 1614 1649
rect 1606 1577 1607 1583
rect 1613 1577 1614 1583
rect 1606 1511 1614 1577
rect 1606 1505 1607 1511
rect 1613 1505 1614 1511
rect 1606 1439 1614 1505
rect 1606 1433 1607 1439
rect 1613 1433 1614 1439
rect 1606 1367 1614 1433
rect 1606 1361 1607 1367
rect 1613 1361 1614 1367
rect 1606 1295 1614 1361
rect 1606 1289 1607 1295
rect 1613 1289 1614 1295
rect 1606 1223 1614 1289
rect 1606 1217 1607 1223
rect 1613 1217 1614 1223
rect 1606 1151 1614 1217
rect 1606 1145 1607 1151
rect 1613 1145 1614 1151
rect 1606 1071 1614 1145
rect 1606 1065 1607 1071
rect 1613 1065 1614 1071
rect 1606 987 1614 1065
rect 1606 981 1607 987
rect 1613 981 1614 987
rect 1606 911 1614 981
rect 1606 905 1607 911
rect 1613 905 1614 911
rect 1606 835 1614 905
rect 1606 829 1607 835
rect 1613 829 1614 835
rect 1606 763 1614 829
rect 1606 757 1607 763
rect 1613 757 1614 763
rect 1606 691 1614 757
rect 1606 685 1607 691
rect 1613 685 1614 691
rect 1606 615 1614 685
rect 1606 609 1607 615
rect 1613 609 1614 615
rect 1606 543 1614 609
rect 1606 537 1607 543
rect 1613 537 1614 543
rect 1606 471 1614 537
rect 1606 465 1607 471
rect 1613 465 1614 471
rect 1606 395 1614 465
rect 1606 389 1607 395
rect 1613 389 1614 395
rect 1606 323 1614 389
rect 1606 317 1607 323
rect 1613 317 1614 323
rect 1606 247 1614 317
rect 1606 241 1607 247
rect 1613 241 1614 247
rect 1606 171 1614 241
rect 1606 165 1607 171
rect 1613 165 1614 171
rect 1606 87 1614 165
rect 1606 81 1607 87
rect 1613 81 1614 87
rect 1606 72 1614 81
rect 1618 1619 1626 1656
rect 1618 1613 1619 1619
rect 1625 1613 1626 1619
rect 1618 1547 1626 1613
rect 1618 1541 1619 1547
rect 1625 1541 1626 1547
rect 1618 1475 1626 1541
rect 1618 1469 1619 1475
rect 1625 1469 1626 1475
rect 1618 1403 1626 1469
rect 1618 1397 1619 1403
rect 1625 1397 1626 1403
rect 1618 1331 1626 1397
rect 1618 1325 1619 1331
rect 1625 1325 1626 1331
rect 1618 1259 1626 1325
rect 1618 1253 1619 1259
rect 1625 1253 1626 1259
rect 1618 1187 1626 1253
rect 1618 1181 1619 1187
rect 1625 1181 1626 1187
rect 1618 1115 1626 1181
rect 1618 1109 1619 1115
rect 1625 1109 1626 1115
rect 1618 1031 1626 1109
rect 1618 1025 1619 1031
rect 1625 1025 1626 1031
rect 1618 951 1626 1025
rect 1618 945 1619 951
rect 1625 945 1626 951
rect 1618 875 1626 945
rect 1618 869 1619 875
rect 1625 869 1626 875
rect 1618 799 1626 869
rect 1618 793 1619 799
rect 1625 793 1626 799
rect 1618 727 1626 793
rect 1618 721 1619 727
rect 1625 721 1626 727
rect 1618 651 1626 721
rect 1618 645 1619 651
rect 1625 645 1626 651
rect 1618 579 1626 645
rect 1618 573 1619 579
rect 1625 573 1626 579
rect 1618 507 1626 573
rect 1618 501 1619 507
rect 1625 501 1626 507
rect 1618 431 1626 501
rect 1618 425 1619 431
rect 1625 425 1626 431
rect 1618 359 1626 425
rect 1618 353 1619 359
rect 1625 353 1626 359
rect 1618 283 1626 353
rect 1618 277 1619 283
rect 1625 277 1626 283
rect 1618 207 1626 277
rect 1618 201 1619 207
rect 1625 201 1626 207
rect 1618 123 1626 201
rect 1618 117 1619 123
rect 1625 117 1626 123
rect 1618 72 1626 117
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__83
timestamp 1731220378
transform 1 0 1576 0 -1 1648
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220378
transform 1 0 104 0 -1 1648
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220378
transform 1 0 1576 0 1 1584
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220378
transform 1 0 104 0 1 1584
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220378
transform 1 0 1576 0 -1 1576
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220378
transform 1 0 104 0 -1 1576
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220378
transform 1 0 1576 0 1 1512
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220378
transform 1 0 104 0 1 1512
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220378
transform 1 0 1576 0 -1 1504
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220378
transform 1 0 104 0 -1 1504
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220378
transform 1 0 1576 0 1 1440
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220378
transform 1 0 104 0 1 1440
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220378
transform 1 0 1576 0 -1 1432
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220378
transform 1 0 104 0 -1 1432
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220378
transform 1 0 1576 0 1 1368
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220378
transform 1 0 104 0 1 1368
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220378
transform 1 0 1576 0 -1 1360
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220378
transform 1 0 104 0 -1 1360
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220378
transform 1 0 1576 0 1 1296
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220378
transform 1 0 104 0 1 1296
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220378
transform 1 0 1576 0 -1 1288
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220378
transform 1 0 104 0 -1 1288
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220378
transform 1 0 1576 0 1 1224
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220378
transform 1 0 104 0 1 1224
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220378
transform 1 0 1576 0 -1 1216
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220378
transform 1 0 104 0 -1 1216
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220378
transform 1 0 1576 0 1 1152
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220378
transform 1 0 104 0 1 1152
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220378
transform 1 0 1576 0 -1 1144
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220378
transform 1 0 104 0 -1 1144
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220378
transform 1 0 1576 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220378
transform 1 0 104 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220378
transform 1 0 1576 0 -1 1064
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220378
transform 1 0 104 0 -1 1064
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220378
transform 1 0 1576 0 1 996
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220378
transform 1 0 104 0 1 996
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220378
transform 1 0 1576 0 -1 980
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220378
transform 1 0 104 0 -1 980
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220378
transform 1 0 1576 0 1 916
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220378
transform 1 0 104 0 1 916
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220378
transform 1 0 1576 0 -1 904
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220378
transform 1 0 104 0 -1 904
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220378
transform 1 0 1576 0 1 840
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220378
transform 1 0 104 0 1 840
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220378
transform 1 0 1576 0 -1 828
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220378
transform 1 0 104 0 -1 828
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220378
transform 1 0 1576 0 1 764
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220378
transform 1 0 104 0 1 764
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220378
transform 1 0 1576 0 -1 756
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220378
transform 1 0 104 0 -1 756
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220378
transform 1 0 1576 0 1 692
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220378
transform 1 0 104 0 1 692
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220378
transform 1 0 1576 0 -1 684
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220378
transform 1 0 104 0 -1 684
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220378
transform 1 0 1576 0 1 616
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220378
transform 1 0 104 0 1 616
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220378
transform 1 0 1576 0 -1 608
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220378
transform 1 0 104 0 -1 608
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220378
transform 1 0 1576 0 1 544
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220378
transform 1 0 104 0 1 544
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220378
transform 1 0 1576 0 -1 536
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220378
transform 1 0 104 0 -1 536
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220378
transform 1 0 1576 0 1 472
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220378
transform 1 0 104 0 1 472
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220378
transform 1 0 1576 0 -1 464
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220378
transform 1 0 104 0 -1 464
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220378
transform 1 0 1576 0 1 396
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220378
transform 1 0 104 0 1 396
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220378
transform 1 0 1576 0 -1 388
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220378
transform 1 0 104 0 -1 388
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220378
transform 1 0 1576 0 1 324
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220378
transform 1 0 104 0 1 324
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220378
transform 1 0 1576 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220378
transform 1 0 104 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220378
transform 1 0 1576 0 1 248
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220378
transform 1 0 104 0 1 248
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220378
transform 1 0 1576 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220378
transform 1 0 104 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220378
transform 1 0 1576 0 1 172
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220378
transform 1 0 104 0 1 172
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220378
transform 1 0 1576 0 -1 164
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220378
transform 1 0 104 0 -1 164
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220378
transform 1 0 1576 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220378
transform 1 0 104 0 1 88
box 7 3 12 24
use _0_0cell_0_0ginvx0  tst_5999_6
timestamp 1731220378
transform 1 0 1504 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5998_6
timestamp 1731220378
transform 1 0 1536 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5997_6
timestamp 1731220378
transform 1 0 1536 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5996_6
timestamp 1731220378
transform 1 0 1504 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5995_6
timestamp 1731220378
transform 1 0 1504 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5994_6
timestamp 1731220378
transform 1 0 1536 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5993_6
timestamp 1731220378
transform 1 0 1536 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5992_6
timestamp 1731220378
transform 1 0 1536 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5991_6
timestamp 1731220378
transform 1 0 1536 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5990_6
timestamp 1731220378
transform 1 0 1504 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5989_6
timestamp 1731220378
transform 1 0 1536 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5988_6
timestamp 1731220378
transform 1 0 1536 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5987_6
timestamp 1731220378
transform 1 0 1536 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5986_6
timestamp 1731220378
transform 1 0 1536 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5985_6
timestamp 1731220378
transform 1 0 1536 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5984_6
timestamp 1731220378
transform 1 0 1536 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5983_6
timestamp 1731220378
transform 1 0 1536 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5982_6
timestamp 1731220378
transform 1 0 1536 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5981_6
timestamp 1731220378
transform 1 0 1496 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5980_6
timestamp 1731220378
transform 1 0 1504 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5979_6
timestamp 1731220378
transform 1 0 1504 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5978_6
timestamp 1731220378
transform 1 0 1536 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5977_6
timestamp 1731220378
transform 1 0 1472 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5976_6
timestamp 1731220378
transform 1 0 1464 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5975_6
timestamp 1731220378
transform 1 0 1480 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5974_6
timestamp 1731220378
transform 1 0 1408 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5973_6
timestamp 1731220378
transform 1 0 1400 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5972_6
timestamp 1731220378
transform 1 0 1480 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5971_6
timestamp 1731220378
transform 1 0 1448 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5970_6
timestamp 1731220378
transform 1 0 1392 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5969_6
timestamp 1731220378
transform 1 0 1344 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5968_6
timestamp 1731220378
transform 1 0 1392 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5967_6
timestamp 1731220378
transform 1 0 1440 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5966_6
timestamp 1731220378
transform 1 0 1496 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5965_6
timestamp 1731220378
transform 1 0 1496 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5964_6
timestamp 1731220378
transform 1 0 1432 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5963_6
timestamp 1731220378
transform 1 0 1376 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5962_6
timestamp 1731220378
transform 1 0 1448 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5961_6
timestamp 1731220378
transform 1 0 1392 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5960_6
timestamp 1731220378
transform 1 0 1336 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5959_6
timestamp 1731220378
transform 1 0 1344 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5958_6
timestamp 1731220378
transform 1 0 1392 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5957_6
timestamp 1731220378
transform 1 0 1448 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5956_6
timestamp 1731220378
transform 1 0 1464 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5955_6
timestamp 1731220378
transform 1 0 1416 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5954_6
timestamp 1731220378
transform 1 0 1376 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5953_6
timestamp 1731220378
transform 1 0 1336 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5952_6
timestamp 1731220378
transform 1 0 1296 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5951_6
timestamp 1731220378
transform 1 0 1256 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5950_6
timestamp 1731220378
transform 1 0 1216 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5949_6
timestamp 1731220378
transform 1 0 1168 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5948_6
timestamp 1731220378
transform 1 0 1296 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5947_6
timestamp 1731220378
transform 1 0 1248 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5946_6
timestamp 1731220378
transform 1 0 1200 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5945_6
timestamp 1731220378
transform 1 0 1144 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5944_6
timestamp 1731220378
transform 1 0 1168 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5943_6
timestamp 1731220378
transform 1 0 1280 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5942_6
timestamp 1731220378
transform 1 0 1224 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5941_6
timestamp 1731220378
transform 1 0 1208 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5940_6
timestamp 1731220378
transform 1 0 1264 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5939_6
timestamp 1731220378
transform 1 0 1320 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5938_6
timestamp 1731220378
transform 1 0 1344 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5937_6
timestamp 1731220378
transform 1 0 1296 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5936_6
timestamp 1731220378
transform 1 0 1256 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5935_6
timestamp 1731220378
transform 1 0 1216 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5934_6
timestamp 1731220378
transform 1 0 1288 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5933_6
timestamp 1731220378
transform 1 0 1224 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5932_6
timestamp 1731220378
transform 1 0 1168 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5931_6
timestamp 1731220378
transform 1 0 1240 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5930_6
timestamp 1731220378
transform 1 0 1320 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5929_6
timestamp 1731220378
transform 1 0 1336 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5928_6
timestamp 1731220378
transform 1 0 1264 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5927_6
timestamp 1731220378
transform 1 0 1192 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5926_6
timestamp 1731220378
transform 1 0 1120 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5925_6
timestamp 1731220378
transform 1 0 1376 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5924_6
timestamp 1731220378
transform 1 0 1296 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5923_6
timestamp 1731220378
transform 1 0 1216 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5922_6
timestamp 1731220378
transform 1 0 1144 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5921_6
timestamp 1731220378
transform 1 0 1080 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5920_6
timestamp 1731220378
transform 1 0 1024 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5919_6
timestamp 1731220378
transform 1 0 984 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5918_6
timestamp 1731220378
transform 1 0 928 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5917_6
timestamp 1731220378
transform 1 0 1040 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5916_6
timestamp 1731220378
transform 1 0 1088 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5915_6
timestamp 1731220378
transform 1 0 1136 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5914_6
timestamp 1731220378
transform 1 0 1192 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5913_6
timestamp 1731220378
transform 1 0 1392 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5912_6
timestamp 1731220378
transform 1 0 1320 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5911_6
timestamp 1731220378
transform 1 0 1256 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5910_6
timestamp 1731220378
transform 1 0 1216 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5909_6
timestamp 1731220378
transform 1 0 1120 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5908_6
timestamp 1731220378
transform 1 0 1320 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5907_6
timestamp 1731220378
transform 1 0 1432 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5906_6
timestamp 1731220378
transform 1 0 1472 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5905_6
timestamp 1731220378
transform 1 0 1384 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5904_6
timestamp 1731220378
transform 1 0 1304 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5903_6
timestamp 1731220378
transform 1 0 1232 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5902_6
timestamp 1731220378
transform 1 0 1160 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5901_6
timestamp 1731220378
transform 1 0 1224 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5900_6
timestamp 1731220378
transform 1 0 1280 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5899_6
timestamp 1731220378
transform 1 0 1328 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5898_6
timestamp 1731220378
transform 1 0 1376 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5897_6
timestamp 1731220378
transform 1 0 1416 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5896_6
timestamp 1731220378
transform 1 0 1464 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5895_6
timestamp 1731220378
transform 1 0 1448 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5894_6
timestamp 1731220378
transform 1 0 1400 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5893_6
timestamp 1731220378
transform 1 0 1344 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5892_6
timestamp 1731220378
transform 1 0 1280 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5891_6
timestamp 1731220378
transform 1 0 1208 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5890_6
timestamp 1731220378
transform 1 0 1432 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5889_6
timestamp 1731220378
transform 1 0 1376 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5888_6
timestamp 1731220378
transform 1 0 1320 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5887_6
timestamp 1731220378
transform 1 0 1264 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5886_6
timestamp 1731220378
transform 1 0 1208 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5885_6
timestamp 1731220378
transform 1 0 1160 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5884_6
timestamp 1731220378
transform 1 0 1128 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5883_6
timestamp 1731220378
transform 1 0 1184 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5882_6
timestamp 1731220378
transform 1 0 1240 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5881_6
timestamp 1731220378
transform 1 0 1296 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5880_6
timestamp 1731220378
transform 1 0 1352 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5879_6
timestamp 1731220378
transform 1 0 1296 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5878_6
timestamp 1731220378
transform 1 0 1232 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5877_6
timestamp 1731220378
transform 1 0 1352 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5876_6
timestamp 1731220378
transform 1 0 1400 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5875_6
timestamp 1731220378
transform 1 0 1448 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5874_6
timestamp 1731220378
transform 1 0 1504 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5873_6
timestamp 1731220378
transform 1 0 1536 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5872_6
timestamp 1731220378
transform 1 0 1536 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5871_6
timestamp 1731220378
transform 1 0 1504 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5870_6
timestamp 1731220378
transform 1 0 1464 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5869_6
timestamp 1731220378
transform 1 0 1416 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5868_6
timestamp 1731220378
transform 1 0 1368 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5867_6
timestamp 1731220378
transform 1 0 1320 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5866_6
timestamp 1731220378
transform 1 0 1264 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5865_6
timestamp 1731220378
transform 1 0 1376 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5864_6
timestamp 1731220378
transform 1 0 1312 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5863_6
timestamp 1731220378
transform 1 0 1248 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5862_6
timestamp 1731220378
transform 1 0 1184 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5861_6
timestamp 1731220378
transform 1 0 1320 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5860_6
timestamp 1731220378
transform 1 0 1272 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5859_6
timestamp 1731220378
transform 1 0 1224 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5858_6
timestamp 1731220378
transform 1 0 1176 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5857_6
timestamp 1731220378
transform 1 0 1136 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5856_6
timestamp 1731220378
transform 1 0 1096 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5855_6
timestamp 1731220378
transform 1 0 1144 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5854_6
timestamp 1731220378
transform 1 0 1200 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5853_6
timestamp 1731220378
transform 1 0 1392 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5852_6
timestamp 1731220378
transform 1 0 1320 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5851_6
timestamp 1731220378
transform 1 0 1256 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5850_6
timestamp 1731220378
transform 1 0 1240 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5849_6
timestamp 1731220378
transform 1 0 1184 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5848_6
timestamp 1731220378
transform 1 0 1296 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5847_6
timestamp 1731220378
transform 1 0 1352 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5846_6
timestamp 1731220378
transform 1 0 1320 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5845_6
timestamp 1731220378
transform 1 0 1264 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5844_6
timestamp 1731220378
transform 1 0 1200 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5843_6
timestamp 1731220378
transform 1 0 1192 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5842_6
timestamp 1731220378
transform 1 0 1264 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5841_6
timestamp 1731220378
transform 1 0 1336 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5840_6
timestamp 1731220378
transform 1 0 1408 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5839_6
timestamp 1731220378
transform 1 0 1480 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5838_6
timestamp 1731220378
transform 1 0 1464 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5837_6
timestamp 1731220378
transform 1 0 1416 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5836_6
timestamp 1731220378
transform 1 0 1368 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5835_6
timestamp 1731220378
transform 1 0 1400 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5834_6
timestamp 1731220378
transform 1 0 1448 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5833_6
timestamp 1731220378
transform 1 0 1472 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5832_6
timestamp 1731220378
transform 1 0 1536 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5831_6
timestamp 1731220378
transform 1 0 1536 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5830_6
timestamp 1731220378
transform 1 0 1504 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5829_6
timestamp 1731220378
transform 1 0 1504 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5828_6
timestamp 1731220378
transform 1 0 1536 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5827_6
timestamp 1731220378
transform 1 0 1536 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5826_6
timestamp 1731220378
transform 1 0 1536 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5825_6
timestamp 1731220378
transform 1 0 1504 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5824_6
timestamp 1731220378
transform 1 0 1536 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5823_6
timestamp 1731220378
transform 1 0 1536 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5822_6
timestamp 1731220378
transform 1 0 1536 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5821_6
timestamp 1731220378
transform 1 0 1536 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5820_6
timestamp 1731220378
transform 1 0 1536 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5819_6
timestamp 1731220378
transform 1 0 1536 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5818_6
timestamp 1731220378
transform 1 0 1496 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5817_6
timestamp 1731220378
transform 1 0 1432 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5816_6
timestamp 1731220378
transform 1 0 1464 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5815_6
timestamp 1731220378
transform 1 0 1472 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5814_6
timestamp 1731220378
transform 1 0 1472 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5813_6
timestamp 1731220378
transform 1 0 1496 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5812_6
timestamp 1731220378
transform 1 0 1432 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5811_6
timestamp 1731220378
transform 1 0 1384 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5810_6
timestamp 1731220378
transform 1 0 1440 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5809_6
timestamp 1731220378
transform 1 0 1496 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5808_6
timestamp 1731220378
transform 1 0 1448 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5807_6
timestamp 1731220378
transform 1 0 1400 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5806_6
timestamp 1731220378
transform 1 0 1352 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5805_6
timestamp 1731220378
transform 1 0 1296 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5804_6
timestamp 1731220378
transform 1 0 1232 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5803_6
timestamp 1731220378
transform 1 0 1160 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5802_6
timestamp 1731220378
transform 1 0 1208 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5801_6
timestamp 1731220378
transform 1 0 1272 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5800_6
timestamp 1731220378
transform 1 0 1328 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5799_6
timestamp 1731220378
transform 1 0 1368 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5798_6
timestamp 1731220378
transform 1 0 1312 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5797_6
timestamp 1731220378
transform 1 0 1256 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5796_6
timestamp 1731220378
transform 1 0 1200 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5795_6
timestamp 1731220378
transform 1 0 1392 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5794_6
timestamp 1731220378
transform 1 0 1320 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5793_6
timestamp 1731220378
transform 1 0 1248 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5792_6
timestamp 1731220378
transform 1 0 1184 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5791_6
timestamp 1731220378
transform 1 0 1120 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5790_6
timestamp 1731220378
transform 1 0 1384 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5789_6
timestamp 1731220378
transform 1 0 1304 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5788_6
timestamp 1731220378
transform 1 0 1232 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5787_6
timestamp 1731220378
transform 1 0 1160 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5786_6
timestamp 1731220378
transform 1 0 1096 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5785_6
timestamp 1731220378
transform 1 0 1032 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5784_6
timestamp 1731220378
transform 1 0 1088 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5783_6
timestamp 1731220378
transform 1 0 1152 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5782_6
timestamp 1731220378
transform 1 0 1224 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5781_6
timestamp 1731220378
transform 1 0 1376 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5780_6
timestamp 1731220378
transform 1 0 1296 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5779_6
timestamp 1731220378
transform 1 0 1240 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5778_6
timestamp 1731220378
transform 1 0 1176 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5777_6
timestamp 1731220378
transform 1 0 1112 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5776_6
timestamp 1731220378
transform 1 0 1368 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5775_6
timestamp 1731220378
transform 1 0 1304 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5774_6
timestamp 1731220378
transform 1 0 1240 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5773_6
timestamp 1731220378
transform 1 0 1184 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5772_6
timestamp 1731220378
transform 1 0 1296 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5771_6
timestamp 1731220378
transform 1 0 1424 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5770_6
timestamp 1731220378
transform 1 0 1360 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5769_6
timestamp 1731220378
transform 1 0 1320 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5768_6
timestamp 1731220378
transform 1 0 1264 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5767_6
timestamp 1731220378
transform 1 0 1368 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5766_6
timestamp 1731220378
transform 1 0 1520 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5765_6
timestamp 1731220378
transform 1 0 1464 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5764_6
timestamp 1731220378
transform 1 0 1416 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5763_6
timestamp 1731220378
transform 1 0 1376 0 -1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5762_6
timestamp 1731220378
transform 1 0 1304 0 -1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5761_6
timestamp 1731220378
transform 1 0 1528 0 -1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5760_6
timestamp 1731220378
transform 1 0 1448 0 -1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5759_6
timestamp 1731220378
transform 1 0 1408 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5758_6
timestamp 1731220378
transform 1 0 1344 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5757_6
timestamp 1731220378
transform 1 0 1536 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5756_6
timestamp 1731220378
transform 1 0 1472 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5755_6
timestamp 1731220378
transform 1 0 1448 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5754_6
timestamp 1731220378
transform 1 0 1392 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5753_6
timestamp 1731220378
transform 1 0 1336 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5752_6
timestamp 1731220378
transform 1 0 1536 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5751_6
timestamp 1731220378
transform 1 0 1504 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5750_6
timestamp 1731220378
transform 1 0 1472 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5749_6
timestamp 1731220378
transform 1 0 1536 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5748_6
timestamp 1731220378
transform 1 0 1536 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5747_6
timestamp 1731220378
transform 1 0 1488 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5746_6
timestamp 1731220378
transform 1 0 1488 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5745_6
timestamp 1731220378
transform 1 0 1536 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5744_6
timestamp 1731220378
transform 1 0 1536 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5743_6
timestamp 1731220378
transform 1 0 1472 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5742_6
timestamp 1731220378
transform 1 0 1536 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5741_6
timestamp 1731220378
transform 1 0 1504 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5740_6
timestamp 1731220378
transform 1 0 1472 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5739_6
timestamp 1731220378
transform 1 0 1440 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5738_6
timestamp 1731220378
transform 1 0 1400 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5737_6
timestamp 1731220378
transform 1 0 1360 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5736_6
timestamp 1731220378
transform 1 0 1320 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5735_6
timestamp 1731220378
transform 1 0 1280 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5734_6
timestamp 1731220378
transform 1 0 1232 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5733_6
timestamp 1731220378
transform 1 0 1184 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5732_6
timestamp 1731220378
transform 1 0 1152 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5731_6
timestamp 1731220378
transform 1 0 1232 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5730_6
timestamp 1731220378
transform 1 0 1392 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5729_6
timestamp 1731220378
transform 1 0 1312 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5728_6
timestamp 1731220378
transform 1 0 1288 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5727_6
timestamp 1731220378
transform 1 0 1224 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5726_6
timestamp 1731220378
transform 1 0 1160 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5725_6
timestamp 1731220378
transform 1 0 1352 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5724_6
timestamp 1731220378
transform 1 0 1416 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5723_6
timestamp 1731220378
transform 1 0 1416 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5722_6
timestamp 1731220378
transform 1 0 1344 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5721_6
timestamp 1731220378
transform 1 0 1272 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5720_6
timestamp 1731220378
transform 1 0 1208 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5719_6
timestamp 1731220378
transform 1 0 1144 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5718_6
timestamp 1731220378
transform 1 0 1392 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5717_6
timestamp 1731220378
transform 1 0 1312 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5716_6
timestamp 1731220378
transform 1 0 1232 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5715_6
timestamp 1731220378
transform 1 0 1152 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5714_6
timestamp 1731220378
transform 1 0 1152 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5713_6
timestamp 1731220378
transform 1 0 1216 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5712_6
timestamp 1731220378
transform 1 0 1280 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5711_6
timestamp 1731220378
transform 1 0 1288 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5710_6
timestamp 1731220378
transform 1 0 1232 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5709_6
timestamp 1731220378
transform 1 0 1168 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5708_6
timestamp 1731220378
transform 1 0 1144 0 -1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5707_6
timestamp 1731220378
transform 1 0 1056 0 -1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5706_6
timestamp 1731220378
transform 1 0 1224 0 -1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5705_6
timestamp 1731220378
transform 1 0 1208 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5704_6
timestamp 1731220378
transform 1 0 1152 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5703_6
timestamp 1731220378
transform 1 0 1096 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5702_6
timestamp 1731220378
transform 1 0 1040 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5701_6
timestamp 1731220378
transform 1 0 992 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5700_6
timestamp 1731220378
transform 1 0 1120 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5699_6
timestamp 1731220378
transform 1 0 1056 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5698_6
timestamp 1731220378
transform 1 0 1048 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5697_6
timestamp 1731220378
transform 1 0 984 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5696_6
timestamp 1731220378
transform 1 0 1032 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5695_6
timestamp 1731220378
transform 1 0 872 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5694_6
timestamp 1731220378
transform 1 0 824 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5693_6
timestamp 1731220378
transform 1 0 776 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5692_6
timestamp 1731220378
transform 1 0 728 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5691_6
timestamp 1731220378
transform 1 0 680 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5690_6
timestamp 1731220378
transform 1 0 664 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5689_6
timestamp 1731220378
transform 1 0 728 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5688_6
timestamp 1731220378
transform 1 0 792 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5687_6
timestamp 1731220378
transform 1 0 720 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5686_6
timestamp 1731220378
transform 1 0 656 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5685_6
timestamp 1731220378
transform 1 0 784 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5684_6
timestamp 1731220378
transform 1 0 832 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5683_6
timestamp 1731220378
transform 1 0 784 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5682_6
timestamp 1731220378
transform 1 0 736 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5681_6
timestamp 1731220378
transform 1 0 680 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5680_6
timestamp 1731220378
transform 1 0 632 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5679_6
timestamp 1731220378
transform 1 0 584 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5678_6
timestamp 1731220378
transform 1 0 536 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5677_6
timestamp 1731220378
transform 1 0 488 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5676_6
timestamp 1731220378
transform 1 0 432 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5675_6
timestamp 1731220378
transform 1 0 456 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5674_6
timestamp 1731220378
transform 1 0 528 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5673_6
timestamp 1731220378
transform 1 0 592 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5672_6
timestamp 1731220378
transform 1 0 600 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5671_6
timestamp 1731220378
transform 1 0 536 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5670_6
timestamp 1731220378
transform 1 0 472 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5669_6
timestamp 1731220378
transform 1 0 408 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5668_6
timestamp 1731220378
transform 1 0 408 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5667_6
timestamp 1731220378
transform 1 0 464 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5666_6
timestamp 1731220378
transform 1 0 520 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5665_6
timestamp 1731220378
transform 1 0 576 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5664_6
timestamp 1731220378
transform 1 0 632 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5663_6
timestamp 1731220378
transform 1 0 584 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5662_6
timestamp 1731220378
transform 1 0 520 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5661_6
timestamp 1731220378
transform 1 0 464 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5660_6
timestamp 1731220378
transform 1 0 648 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5659_6
timestamp 1731220378
transform 1 0 712 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5658_6
timestamp 1731220378
transform 1 0 784 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5657_6
timestamp 1731220378
transform 1 0 776 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5656_6
timestamp 1731220378
transform 1 0 720 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5655_6
timestamp 1731220378
transform 1 0 664 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5654_6
timestamp 1731220378
transform 1 0 608 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5653_6
timestamp 1731220378
transform 1 0 552 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5652_6
timestamp 1731220378
transform 1 0 776 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5651_6
timestamp 1731220378
transform 1 0 704 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5650_6
timestamp 1731220378
transform 1 0 632 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5649_6
timestamp 1731220378
transform 1 0 560 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5648_6
timestamp 1731220378
transform 1 0 496 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5647_6
timestamp 1731220378
transform 1 0 432 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5646_6
timestamp 1731220378
transform 1 0 720 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5645_6
timestamp 1731220378
transform 1 0 656 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5644_6
timestamp 1731220378
transform 1 0 592 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5643_6
timestamp 1731220378
transform 1 0 536 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5642_6
timestamp 1731220378
transform 1 0 480 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5641_6
timestamp 1731220378
transform 1 0 440 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5640_6
timestamp 1731220378
transform 1 0 504 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5639_6
timestamp 1731220378
transform 1 0 536 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5638_6
timestamp 1731220378
transform 1 0 568 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5637_6
timestamp 1731220378
transform 1 0 704 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5636_6
timestamp 1731220378
transform 1 0 656 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5635_6
timestamp 1731220378
transform 1 0 608 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5634_6
timestamp 1731220378
transform 1 0 552 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5633_6
timestamp 1731220378
transform 1 0 496 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5632_6
timestamp 1731220378
transform 1 0 608 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5631_6
timestamp 1731220378
transform 1 0 656 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5630_6
timestamp 1731220378
transform 1 0 696 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5629_6
timestamp 1731220378
transform 1 0 728 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5628_6
timestamp 1731220378
transform 1 0 760 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5627_6
timestamp 1731220378
transform 1 0 712 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5626_6
timestamp 1731220378
transform 1 0 664 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5625_6
timestamp 1731220378
transform 1 0 608 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5624_6
timestamp 1731220378
transform 1 0 552 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5623_6
timestamp 1731220378
transform 1 0 488 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5622_6
timestamp 1731220378
transform 1 0 752 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5621_6
timestamp 1731220378
transform 1 0 688 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5620_6
timestamp 1731220378
transform 1 0 616 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5619_6
timestamp 1731220378
transform 1 0 552 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5618_6
timestamp 1731220378
transform 1 0 496 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5617_6
timestamp 1731220378
transform 1 0 440 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5616_6
timestamp 1731220378
transform 1 0 760 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5615_6
timestamp 1731220378
transform 1 0 672 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5614_6
timestamp 1731220378
transform 1 0 584 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5613_6
timestamp 1731220378
transform 1 0 504 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5612_6
timestamp 1731220378
transform 1 0 432 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5611_6
timestamp 1731220378
transform 1 0 376 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5610_6
timestamp 1731220378
transform 1 0 416 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5609_6
timestamp 1731220378
transform 1 0 488 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5608_6
timestamp 1731220378
transform 1 0 456 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5607_6
timestamp 1731220378
transform 1 0 416 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5606_6
timestamp 1731220378
transform 1 0 408 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5605_6
timestamp 1731220378
transform 1 0 376 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5604_6
timestamp 1731220378
transform 1 0 320 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5603_6
timestamp 1731220378
transform 1 0 312 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5602_6
timestamp 1731220378
transform 1 0 344 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5601_6
timestamp 1731220378
transform 1 0 376 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5600_6
timestamp 1731220378
transform 1 0 392 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5599_6
timestamp 1731220378
transform 1 0 464 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5598_6
timestamp 1731220378
transform 1 0 416 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5597_6
timestamp 1731220378
transform 1 0 352 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5596_6
timestamp 1731220378
transform 1 0 336 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5595_6
timestamp 1731220378
transform 1 0 288 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5594_6
timestamp 1731220378
transform 1 0 304 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5593_6
timestamp 1731220378
transform 1 0 360 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5592_6
timestamp 1731220378
transform 1 0 352 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5591_6
timestamp 1731220378
transform 1 0 416 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5590_6
timestamp 1731220378
transform 1 0 456 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5589_6
timestamp 1731220378
transform 1 0 376 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5588_6
timestamp 1731220378
transform 1 0 288 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5587_6
timestamp 1731220378
transform 1 0 328 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5586_6
timestamp 1731220378
transform 1 0 384 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5585_6
timestamp 1731220378
transform 1 0 360 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5584_6
timestamp 1731220378
transform 1 0 328 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5583_6
timestamp 1731220378
transform 1 0 304 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5582_6
timestamp 1731220378
transform 1 0 272 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5581_6
timestamp 1731220378
transform 1 0 240 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5580_6
timestamp 1731220378
transform 1 0 248 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5579_6
timestamp 1731220378
transform 1 0 296 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5578_6
timestamp 1731220378
transform 1 0 336 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5577_6
timestamp 1731220378
transform 1 0 352 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5576_6
timestamp 1731220378
transform 1 0 304 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5575_6
timestamp 1731220378
transform 1 0 288 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5574_6
timestamp 1731220378
transform 1 0 344 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5573_6
timestamp 1731220378
transform 1 0 400 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5572_6
timestamp 1731220378
transform 1 0 416 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5571_6
timestamp 1731220378
transform 1 0 384 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5570_6
timestamp 1731220378
transform 1 0 352 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5569_6
timestamp 1731220378
transform 1 0 320 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5568_6
timestamp 1731220378
transform 1 0 288 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5567_6
timestamp 1731220378
transform 1 0 256 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5566_6
timestamp 1731220378
transform 1 0 224 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5565_6
timestamp 1731220378
transform 1 0 192 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5564_6
timestamp 1731220378
transform 1 0 160 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5563_6
timestamp 1731220378
transform 1 0 128 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5562_6
timestamp 1731220378
transform 1 0 136 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5561_6
timestamp 1731220378
transform 1 0 184 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5560_6
timestamp 1731220378
transform 1 0 232 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5559_6
timestamp 1731220378
transform 1 0 256 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5558_6
timestamp 1731220378
transform 1 0 208 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5557_6
timestamp 1731220378
transform 1 0 160 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5556_6
timestamp 1731220378
transform 1 0 128 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5555_6
timestamp 1731220378
transform 1 0 128 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5554_6
timestamp 1731220378
transform 1 0 160 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5553_6
timestamp 1731220378
transform 1 0 200 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5552_6
timestamp 1731220378
transform 1 0 208 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5551_6
timestamp 1731220378
transform 1 0 176 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5550_6
timestamp 1731220378
transform 1 0 144 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5549_6
timestamp 1731220378
transform 1 0 184 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5548_6
timestamp 1731220378
transform 1 0 216 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5547_6
timestamp 1731220378
transform 1 0 248 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5546_6
timestamp 1731220378
transform 1 0 288 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5545_6
timestamp 1731220378
transform 1 0 272 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5544_6
timestamp 1731220378
transform 1 0 216 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5543_6
timestamp 1731220378
transform 1 0 168 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5542_6
timestamp 1731220378
transform 1 0 128 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5541_6
timestamp 1731220378
transform 1 0 128 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5540_6
timestamp 1731220378
transform 1 0 200 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5539_6
timestamp 1731220378
transform 1 0 288 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5538_6
timestamp 1731220378
transform 1 0 224 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5537_6
timestamp 1731220378
transform 1 0 160 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5536_6
timestamp 1731220378
transform 1 0 128 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5535_6
timestamp 1731220378
transform 1 0 128 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5534_6
timestamp 1731220378
transform 1 0 160 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5533_6
timestamp 1731220378
transform 1 0 192 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5532_6
timestamp 1731220378
transform 1 0 248 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5531_6
timestamp 1731220378
transform 1 0 240 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5530_6
timestamp 1731220378
transform 1 0 192 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5529_6
timestamp 1731220378
transform 1 0 160 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5528_6
timestamp 1731220378
transform 1 0 128 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5527_6
timestamp 1731220378
transform 1 0 128 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5526_6
timestamp 1731220378
transform 1 0 168 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5525_6
timestamp 1731220378
transform 1 0 224 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5524_6
timestamp 1731220378
transform 1 0 288 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5523_6
timestamp 1731220378
transform 1 0 320 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5522_6
timestamp 1731220378
transform 1 0 248 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5521_6
timestamp 1731220378
transform 1 0 184 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5520_6
timestamp 1731220378
transform 1 0 216 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5519_6
timestamp 1731220378
transform 1 0 248 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5518_6
timestamp 1731220378
transform 1 0 280 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5517_6
timestamp 1731220378
transform 1 0 264 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5516_6
timestamp 1731220378
transform 1 0 208 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5515_6
timestamp 1731220378
transform 1 0 160 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5514_6
timestamp 1731220378
transform 1 0 152 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5513_6
timestamp 1731220378
transform 1 0 200 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5512_6
timestamp 1731220378
transform 1 0 200 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5511_6
timestamp 1731220378
transform 1 0 160 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5510_6
timestamp 1731220378
transform 1 0 128 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5509_6
timestamp 1731220378
transform 1 0 128 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5508_6
timestamp 1731220378
transform 1 0 160 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5507_6
timestamp 1731220378
transform 1 0 192 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5506_6
timestamp 1731220378
transform 1 0 160 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5505_6
timestamp 1731220378
transform 1 0 128 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5504_6
timestamp 1731220378
transform 1 0 128 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5503_6
timestamp 1731220378
transform 1 0 160 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5502_6
timestamp 1731220378
transform 1 0 200 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5501_6
timestamp 1731220378
transform 1 0 160 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5500_6
timestamp 1731220378
transform 1 0 128 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5499_6
timestamp 1731220378
transform 1 0 128 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5498_6
timestamp 1731220378
transform 1 0 160 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5497_6
timestamp 1731220378
transform 1 0 216 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5496_6
timestamp 1731220378
transform 1 0 240 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5495_6
timestamp 1731220378
transform 1 0 184 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5494_6
timestamp 1731220378
transform 1 0 144 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5493_6
timestamp 1731220378
transform 1 0 152 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5492_6
timestamp 1731220378
transform 1 0 192 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5491_6
timestamp 1731220378
transform 1 0 248 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5490_6
timestamp 1731220378
transform 1 0 304 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5489_6
timestamp 1731220378
transform 1 0 368 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5488_6
timestamp 1731220378
transform 1 0 432 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5487_6
timestamp 1731220378
transform 1 0 424 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5486_6
timestamp 1731220378
transform 1 0 360 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5485_6
timestamp 1731220378
transform 1 0 296 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5484_6
timestamp 1731220378
transform 1 0 272 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5483_6
timestamp 1731220378
transform 1 0 328 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5482_6
timestamp 1731220378
transform 1 0 384 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5481_6
timestamp 1731220378
transform 1 0 336 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5480_6
timestamp 1731220378
transform 1 0 296 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5479_6
timestamp 1731220378
transform 1 0 248 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5478_6
timestamp 1731220378
transform 1 0 216 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5477_6
timestamp 1731220378
transform 1 0 280 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5476_6
timestamp 1731220378
transform 1 0 344 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5475_6
timestamp 1731220378
transform 1 0 352 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5474_6
timestamp 1731220378
transform 1 0 296 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5473_6
timestamp 1731220378
transform 1 0 240 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5472_6
timestamp 1731220378
transform 1 0 192 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5471_6
timestamp 1731220378
transform 1 0 248 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5470_6
timestamp 1731220378
transform 1 0 312 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5469_6
timestamp 1731220378
transform 1 0 384 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5468_6
timestamp 1731220378
transform 1 0 360 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5467_6
timestamp 1731220378
transform 1 0 304 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5466_6
timestamp 1731220378
transform 1 0 248 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5465_6
timestamp 1731220378
transform 1 0 248 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5464_6
timestamp 1731220378
transform 1 0 296 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5463_6
timestamp 1731220378
transform 1 0 352 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5462_6
timestamp 1731220378
transform 1 0 464 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5461_6
timestamp 1731220378
transform 1 0 424 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5460_6
timestamp 1731220378
transform 1 0 416 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5459_6
timestamp 1731220378
transform 1 0 456 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5458_6
timestamp 1731220378
transform 1 0 512 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5457_6
timestamp 1731220378
transform 1 0 640 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5456_6
timestamp 1731220378
transform 1 0 576 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5455_6
timestamp 1731220378
transform 1 0 528 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5454_6
timestamp 1731220378
transform 1 0 480 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5453_6
timestamp 1731220378
transform 1 0 520 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5452_6
timestamp 1731220378
transform 1 0 472 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5451_6
timestamp 1731220378
transform 1 0 536 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5450_6
timestamp 1731220378
transform 1 0 536 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5449_6
timestamp 1731220378
transform 1 0 480 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5448_6
timestamp 1731220378
transform 1 0 416 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5447_6
timestamp 1731220378
transform 1 0 560 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5446_6
timestamp 1731220378
transform 1 0 632 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5445_6
timestamp 1731220378
transform 1 0 664 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5444_6
timestamp 1731220378
transform 1 0 600 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5443_6
timestamp 1731220378
transform 1 0 544 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5442_6
timestamp 1731220378
transform 1 0 616 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5441_6
timestamp 1731220378
transform 1 0 608 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5440_6
timestamp 1731220378
transform 1 0 680 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5439_6
timestamp 1731220378
transform 1 0 632 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5438_6
timestamp 1731220378
transform 1 0 576 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5437_6
timestamp 1731220378
transform 1 0 584 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5436_6
timestamp 1731220378
transform 1 0 640 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5435_6
timestamp 1731220378
transform 1 0 696 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5434_6
timestamp 1731220378
transform 1 0 752 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5433_6
timestamp 1731220378
transform 1 0 752 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5432_6
timestamp 1731220378
transform 1 0 688 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5431_6
timestamp 1731220378
transform 1 0 752 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5430_6
timestamp 1731220378
transform 1 0 696 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5429_6
timestamp 1731220378
transform 1 0 768 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5428_6
timestamp 1731220378
transform 1 0 792 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5427_6
timestamp 1731220378
transform 1 0 728 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5426_6
timestamp 1731220378
transform 1 0 712 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5425_6
timestamp 1731220378
transform 1 0 784 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5424_6
timestamp 1731220378
transform 1 0 856 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5423_6
timestamp 1731220378
transform 1 0 928 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5422_6
timestamp 1731220378
transform 1 0 992 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5421_6
timestamp 1731220378
transform 1 0 928 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5420_6
timestamp 1731220378
transform 1 0 864 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5419_6
timestamp 1731220378
transform 1 0 840 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5418_6
timestamp 1731220378
transform 1 0 912 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5417_6
timestamp 1731220378
transform 1 0 984 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5416_6
timestamp 1731220378
transform 1 0 1000 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5415_6
timestamp 1731220378
transform 1 0 912 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5414_6
timestamp 1731220378
transform 1 0 832 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5413_6
timestamp 1731220378
transform 1 0 816 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5412_6
timestamp 1731220378
transform 1 0 880 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5411_6
timestamp 1731220378
transform 1 0 944 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5410_6
timestamp 1731220378
transform 1 0 880 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5409_6
timestamp 1731220378
transform 1 0 816 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5408_6
timestamp 1731220378
transform 1 0 792 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5407_6
timestamp 1731220378
transform 1 0 712 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5406_6
timestamp 1731220378
transform 1 0 880 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5405_6
timestamp 1731220378
transform 1 0 832 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5404_6
timestamp 1731220378
transform 1 0 776 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5403_6
timestamp 1731220378
transform 1 0 720 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5402_6
timestamp 1731220378
transform 1 0 656 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5401_6
timestamp 1731220378
transform 1 0 592 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5400_6
timestamp 1731220378
transform 1 0 528 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5399_6
timestamp 1731220378
transform 1 0 760 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5398_6
timestamp 1731220378
transform 1 0 704 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5397_6
timestamp 1731220378
transform 1 0 648 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5396_6
timestamp 1731220378
transform 1 0 592 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5395_6
timestamp 1731220378
transform 1 0 536 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5394_6
timestamp 1731220378
transform 1 0 472 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5393_6
timestamp 1731220378
transform 1 0 672 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5392_6
timestamp 1731220378
transform 1 0 616 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5391_6
timestamp 1731220378
transform 1 0 560 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5390_6
timestamp 1731220378
transform 1 0 504 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5389_6
timestamp 1731220378
transform 1 0 448 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5388_6
timestamp 1731220378
transform 1 0 392 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5387_6
timestamp 1731220378
transform 1 0 416 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5386_6
timestamp 1731220378
transform 1 0 472 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5385_6
timestamp 1731220378
transform 1 0 528 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5384_6
timestamp 1731220378
transform 1 0 728 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5383_6
timestamp 1731220378
transform 1 0 656 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5382_6
timestamp 1731220378
transform 1 0 592 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5381_6
timestamp 1731220378
transform 1 0 536 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5380_6
timestamp 1731220378
transform 1 0 480 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5379_6
timestamp 1731220378
transform 1 0 584 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5378_6
timestamp 1731220378
transform 1 0 632 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5377_6
timestamp 1731220378
transform 1 0 672 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5376_6
timestamp 1731220378
transform 1 0 712 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5375_6
timestamp 1731220378
transform 1 0 744 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5374_6
timestamp 1731220378
transform 1 0 696 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5373_6
timestamp 1731220378
transform 1 0 648 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5372_6
timestamp 1731220378
transform 1 0 592 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5371_6
timestamp 1731220378
transform 1 0 528 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5370_6
timestamp 1731220378
transform 1 0 744 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5369_6
timestamp 1731220378
transform 1 0 680 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5368_6
timestamp 1731220378
transform 1 0 624 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5367_6
timestamp 1731220378
transform 1 0 560 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5366_6
timestamp 1731220378
transform 1 0 496 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5365_6
timestamp 1731220378
transform 1 0 440 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5364_6
timestamp 1731220378
transform 1 0 728 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5363_6
timestamp 1731220378
transform 1 0 656 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5362_6
timestamp 1731220378
transform 1 0 584 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5361_6
timestamp 1731220378
transform 1 0 512 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5360_6
timestamp 1731220378
transform 1 0 448 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5359_6
timestamp 1731220378
transform 1 0 400 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5358_6
timestamp 1731220378
transform 1 0 728 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5357_6
timestamp 1731220378
transform 1 0 640 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5356_6
timestamp 1731220378
transform 1 0 552 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5355_6
timestamp 1731220378
transform 1 0 472 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5354_6
timestamp 1731220378
transform 1 0 400 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5353_6
timestamp 1731220378
transform 1 0 344 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5352_6
timestamp 1731220378
transform 1 0 376 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5351_6
timestamp 1731220378
transform 1 0 432 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5350_6
timestamp 1731220378
transform 1 0 504 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5349_6
timestamp 1731220378
transform 1 0 760 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5348_6
timestamp 1731220378
transform 1 0 672 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5347_6
timestamp 1731220378
transform 1 0 584 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5346_6
timestamp 1731220378
transform 1 0 528 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5345_6
timestamp 1731220378
transform 1 0 464 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5344_6
timestamp 1731220378
transform 1 0 408 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5343_6
timestamp 1731220378
transform 1 0 744 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5342_6
timestamp 1731220378
transform 1 0 672 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5341_6
timestamp 1731220378
transform 1 0 600 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5340_6
timestamp 1731220378
transform 1 0 568 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5339_6
timestamp 1731220378
transform 1 0 512 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5338_6
timestamp 1731220378
transform 1 0 456 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5337_6
timestamp 1731220378
transform 1 0 736 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5336_6
timestamp 1731220378
transform 1 0 680 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5335_6
timestamp 1731220378
transform 1 0 624 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5334_6
timestamp 1731220378
transform 1 0 512 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5333_6
timestamp 1731220378
transform 1 0 480 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5332_6
timestamp 1731220378
transform 1 0 448 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5331_6
timestamp 1731220378
transform 1 0 544 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5330_6
timestamp 1731220378
transform 1 0 576 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5329_6
timestamp 1731220378
transform 1 0 608 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5328_6
timestamp 1731220378
transform 1 0 640 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5327_6
timestamp 1731220378
transform 1 0 672 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5326_6
timestamp 1731220378
transform 1 0 704 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5325_6
timestamp 1731220378
transform 1 0 736 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5324_6
timestamp 1731220378
transform 1 0 768 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5323_6
timestamp 1731220378
transform 1 0 800 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5322_6
timestamp 1731220378
transform 1 0 832 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5321_6
timestamp 1731220378
transform 1 0 864 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5320_6
timestamp 1731220378
transform 1 0 896 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5319_6
timestamp 1731220378
transform 1 0 936 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5318_6
timestamp 1731220378
transform 1 0 976 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5317_6
timestamp 1731220378
transform 1 0 1120 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5316_6
timestamp 1731220378
transform 1 0 1072 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5315_6
timestamp 1731220378
transform 1 0 1024 0 1 84
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5314_6
timestamp 1731220378
transform 1 0 904 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5313_6
timestamp 1731220378
transform 1 0 848 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5312_6
timestamp 1731220378
transform 1 0 792 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5311_6
timestamp 1731220378
transform 1 0 1088 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5310_6
timestamp 1731220378
transform 1 0 1032 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5309_6
timestamp 1731220378
transform 1 0 968 0 -1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5308_6
timestamp 1731220378
transform 1 0 936 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5307_6
timestamp 1731220378
transform 1 0 872 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5306_6
timestamp 1731220378
transform 1 0 808 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5305_6
timestamp 1731220378
transform 1 0 1112 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5304_6
timestamp 1731220378
transform 1 0 1056 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5303_6
timestamp 1731220378
transform 1 0 1000 0 1 168
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5302_6
timestamp 1731220378
transform 1 0 976 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5301_6
timestamp 1731220378
transform 1 0 912 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5300_6
timestamp 1731220378
transform 1 0 840 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5299_6
timestamp 1731220378
transform 1 0 1040 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5298_6
timestamp 1731220378
transform 1 0 1096 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5297_6
timestamp 1731220378
transform 1 0 1152 0 -1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5296_6
timestamp 1731220378
transform 1 0 1168 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5295_6
timestamp 1731220378
transform 1 0 1112 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5294_6
timestamp 1731220378
transform 1 0 1048 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5293_6
timestamp 1731220378
transform 1 0 976 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5292_6
timestamp 1731220378
transform 1 0 896 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5291_6
timestamp 1731220378
transform 1 0 816 0 1 244
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5290_6
timestamp 1731220378
transform 1 0 1160 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5289_6
timestamp 1731220378
transform 1 0 1088 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5288_6
timestamp 1731220378
transform 1 0 1016 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5287_6
timestamp 1731220378
transform 1 0 944 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5286_6
timestamp 1731220378
transform 1 0 872 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5285_6
timestamp 1731220378
transform 1 0 800 0 -1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5284_6
timestamp 1731220378
transform 1 0 1096 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5283_6
timestamp 1731220378
transform 1 0 1024 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5282_6
timestamp 1731220378
transform 1 0 944 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5281_6
timestamp 1731220378
transform 1 0 872 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5280_6
timestamp 1731220378
transform 1 0 808 0 1 320
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5279_6
timestamp 1731220378
transform 1 0 1048 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5278_6
timestamp 1731220378
transform 1 0 976 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5277_6
timestamp 1731220378
transform 1 0 912 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5276_6
timestamp 1731220378
transform 1 0 856 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5275_6
timestamp 1731220378
transform 1 0 800 0 -1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5274_6
timestamp 1731220378
transform 1 0 968 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5273_6
timestamp 1731220378
transform 1 0 912 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5272_6
timestamp 1731220378
transform 1 0 856 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5271_6
timestamp 1731220378
transform 1 0 800 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5270_6
timestamp 1731220378
transform 1 0 752 0 1 392
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5269_6
timestamp 1731220378
transform 1 0 800 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5268_6
timestamp 1731220378
transform 1 0 864 0 -1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5267_6
timestamp 1731220378
transform 1 0 1032 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5266_6
timestamp 1731220378
transform 1 0 952 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5265_6
timestamp 1731220378
transform 1 0 880 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5264_6
timestamp 1731220378
transform 1 0 808 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5263_6
timestamp 1731220378
transform 1 0 736 0 1 468
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5262_6
timestamp 1731220378
transform 1 0 824 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5261_6
timestamp 1731220378
transform 1 0 888 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5260_6
timestamp 1731220378
transform 1 0 1088 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5259_6
timestamp 1731220378
transform 1 0 1024 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5258_6
timestamp 1731220378
transform 1 0 960 0 -1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5257_6
timestamp 1731220378
transform 1 0 896 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5256_6
timestamp 1731220378
transform 1 0 960 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5255_6
timestamp 1731220378
transform 1 0 1032 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5254_6
timestamp 1731220378
transform 1 0 1096 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5253_6
timestamp 1731220378
transform 1 0 1160 0 1 540
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5252_6
timestamp 1731220378
transform 1 0 1136 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5251_6
timestamp 1731220378
transform 1 0 1056 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5250_6
timestamp 1731220378
transform 1 0 968 0 -1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5249_6
timestamp 1731220378
transform 1 0 936 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5248_6
timestamp 1731220378
transform 1 0 992 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5247_6
timestamp 1731220378
transform 1 0 1048 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5246_6
timestamp 1731220378
transform 1 0 1104 0 1 612
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5245_6
timestamp 1731220378
transform 1 0 1072 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5244_6
timestamp 1731220378
transform 1 0 1008 0 -1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5243_6
timestamp 1731220378
transform 1 0 1080 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5242_6
timestamp 1731220378
transform 1 0 1160 0 1 688
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5241_6
timestamp 1731220378
transform 1 0 1200 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5240_6
timestamp 1731220378
transform 1 0 1128 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5239_6
timestamp 1731220378
transform 1 0 1056 0 -1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5238_6
timestamp 1731220378
transform 1 0 1056 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5237_6
timestamp 1731220378
transform 1 0 1120 0 1 760
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5236_6
timestamp 1731220378
transform 1 0 1048 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5235_6
timestamp 1731220378
transform 1 0 992 0 -1 832
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5234_6
timestamp 1731220378
transform 1 0 1088 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5233_6
timestamp 1731220378
transform 1 0 1032 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5232_6
timestamp 1731220378
transform 1 0 976 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5231_6
timestamp 1731220378
transform 1 0 912 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5230_6
timestamp 1731220378
transform 1 0 840 0 1 836
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5229_6
timestamp 1731220378
transform 1 0 1128 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5228_6
timestamp 1731220378
transform 1 0 1072 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5227_6
timestamp 1731220378
transform 1 0 1008 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5226_6
timestamp 1731220378
transform 1 0 944 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5225_6
timestamp 1731220378
transform 1 0 880 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5224_6
timestamp 1731220378
transform 1 0 816 0 -1 908
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5223_6
timestamp 1731220378
transform 1 0 1136 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5222_6
timestamp 1731220378
transform 1 0 1072 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5221_6
timestamp 1731220378
transform 1 0 1000 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5220_6
timestamp 1731220378
transform 1 0 928 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5219_6
timestamp 1731220378
transform 1 0 864 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5218_6
timestamp 1731220378
transform 1 0 808 0 1 912
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5217_6
timestamp 1731220378
transform 1 0 1120 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5216_6
timestamp 1731220378
transform 1 0 1040 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5215_6
timestamp 1731220378
transform 1 0 960 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5214_6
timestamp 1731220378
transform 1 0 888 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5213_6
timestamp 1731220378
transform 1 0 824 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5212_6
timestamp 1731220378
transform 1 0 768 0 -1 984
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5211_6
timestamp 1731220378
transform 1 0 768 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5210_6
timestamp 1731220378
transform 1 0 840 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5209_6
timestamp 1731220378
transform 1 0 920 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5208_6
timestamp 1731220378
transform 1 0 1080 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5207_6
timestamp 1731220378
transform 1 0 1000 0 1 992
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5206_6
timestamp 1731220378
transform 1 0 928 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5205_6
timestamp 1731220378
transform 1 0 856 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5204_6
timestamp 1731220378
transform 1 0 784 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5203_6
timestamp 1731220378
transform 1 0 1000 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5202_6
timestamp 1731220378
transform 1 0 1072 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5201_6
timestamp 1731220378
transform 1 0 1144 0 -1 1068
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5200_6
timestamp 1731220378
transform 1 0 1144 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5199_6
timestamp 1731220378
transform 1 0 1088 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5198_6
timestamp 1731220378
transform 1 0 1032 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5197_6
timestamp 1731220378
transform 1 0 976 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5196_6
timestamp 1731220378
transform 1 0 912 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5195_6
timestamp 1731220378
transform 1 0 848 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5194_6
timestamp 1731220378
transform 1 0 1056 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5193_6
timestamp 1731220378
transform 1 0 1000 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5192_6
timestamp 1731220378
transform 1 0 944 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5191_6
timestamp 1731220378
transform 1 0 888 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5190_6
timestamp 1731220378
transform 1 0 832 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5189_6
timestamp 1731220378
transform 1 0 848 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5188_6
timestamp 1731220378
transform 1 0 912 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5187_6
timestamp 1731220378
transform 1 0 976 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5186_6
timestamp 1731220378
transform 1 0 976 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5185_6
timestamp 1731220378
transform 1 0 928 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5184_6
timestamp 1731220378
transform 1 0 920 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5183_6
timestamp 1731220378
transform 1 0 856 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5182_6
timestamp 1731220378
transform 1 0 848 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5181_6
timestamp 1731220378
transform 1 0 920 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5180_6
timestamp 1731220378
transform 1 0 984 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5179_6
timestamp 1731220378
transform 1 0 928 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5178_6
timestamp 1731220378
transform 1 0 880 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5177_6
timestamp 1731220378
transform 1 0 856 0 -1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5176_6
timestamp 1731220378
transform 1 0 744 0 -1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5175_6
timestamp 1731220378
transform 1 0 960 0 -1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5174_6
timestamp 1731220378
transform 1 0 1104 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5173_6
timestamp 1731220378
transform 1 0 1048 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5172_6
timestamp 1731220378
transform 1 0 992 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5171_6
timestamp 1731220378
transform 1 0 944 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5170_6
timestamp 1731220378
transform 1 0 888 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5169_6
timestamp 1731220378
transform 1 0 1088 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5168_6
timestamp 1731220378
transform 1 0 1016 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5167_6
timestamp 1731220378
transform 1 0 944 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5166_6
timestamp 1731220378
transform 1 0 872 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5165_6
timestamp 1731220378
transform 1 0 1080 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5164_6
timestamp 1731220378
transform 1 0 1008 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5163_6
timestamp 1731220378
transform 1 0 936 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5162_6
timestamp 1731220378
transform 1 0 872 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5161_6
timestamp 1731220378
transform 1 0 928 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5160_6
timestamp 1731220378
transform 1 0 1000 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5159_6
timestamp 1731220378
transform 1 0 1072 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5158_6
timestamp 1731220378
transform 1 0 1096 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5157_6
timestamp 1731220378
transform 1 0 1032 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5156_6
timestamp 1731220378
transform 1 0 960 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5155_6
timestamp 1731220378
transform 1 0 1008 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5154_6
timestamp 1731220378
transform 1 0 1080 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5153_6
timestamp 1731220378
transform 1 0 1136 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5152_6
timestamp 1731220378
transform 1 0 1088 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5151_6
timestamp 1731220378
transform 1 0 1040 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5150_6
timestamp 1731220378
transform 1 0 984 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5149_6
timestamp 1731220378
transform 1 0 928 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5148_6
timestamp 1731220378
transform 1 0 880 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5147_6
timestamp 1731220378
transform 1 0 832 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5146_6
timestamp 1731220378
transform 1 0 784 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5145_6
timestamp 1731220378
transform 1 0 848 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5144_6
timestamp 1731220378
transform 1 0 928 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5143_6
timestamp 1731220378
transform 1 0 888 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5142_6
timestamp 1731220378
transform 1 0 816 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5141_6
timestamp 1731220378
transform 1 0 752 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5140_6
timestamp 1731220378
transform 1 0 712 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5139_6
timestamp 1731220378
transform 1 0 776 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5138_6
timestamp 1731220378
transform 1 0 848 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5137_6
timestamp 1731220378
transform 1 0 808 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5136_6
timestamp 1731220378
transform 1 0 744 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5135_6
timestamp 1731220378
transform 1 0 680 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5134_6
timestamp 1731220378
transform 1 0 672 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5133_6
timestamp 1731220378
transform 1 0 736 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5132_6
timestamp 1731220378
transform 1 0 808 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5131_6
timestamp 1731220378
transform 1 0 832 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5130_6
timestamp 1731220378
transform 1 0 768 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5129_6
timestamp 1731220378
transform 1 0 704 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5128_6
timestamp 1731220378
transform 1 0 640 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5127_6
timestamp 1731220378
transform 1 0 576 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5126_6
timestamp 1731220378
transform 1 0 512 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5125_6
timestamp 1731220378
transform 1 0 448 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5124_6
timestamp 1731220378
transform 1 0 464 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5123_6
timestamp 1731220378
transform 1 0 536 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5122_6
timestamp 1731220378
transform 1 0 608 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5121_6
timestamp 1731220378
transform 1 0 624 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5120_6
timestamp 1731220378
transform 1 0 568 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5119_6
timestamp 1731220378
transform 1 0 504 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5118_6
timestamp 1731220378
transform 1 0 448 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5117_6
timestamp 1731220378
transform 1 0 648 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5116_6
timestamp 1731220378
transform 1 0 584 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5115_6
timestamp 1731220378
transform 1 0 520 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5114_6
timestamp 1731220378
transform 1 0 456 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5113_6
timestamp 1731220378
transform 1 0 400 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5112_6
timestamp 1731220378
transform 1 0 464 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5111_6
timestamp 1731220378
transform 1 0 520 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5110_6
timestamp 1731220378
transform 1 0 576 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5109_6
timestamp 1731220378
transform 1 0 632 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5108_6
timestamp 1731220378
transform 1 0 688 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5107_6
timestamp 1731220378
transform 1 0 768 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5106_6
timestamp 1731220378
transform 1 0 696 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5105_6
timestamp 1731220378
transform 1 0 632 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5104_6
timestamp 1731220378
transform 1 0 576 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5103_6
timestamp 1731220378
transform 1 0 736 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5102_6
timestamp 1731220378
transform 1 0 688 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5101_6
timestamp 1731220378
transform 1 0 640 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_5100_6
timestamp 1731220378
transform 1 0 592 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_599_6
timestamp 1731220378
transform 1 0 544 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_598_6
timestamp 1731220378
transform 1 0 496 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_597_6
timestamp 1731220378
transform 1 0 448 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_596_6
timestamp 1731220378
transform 1 0 400 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_595_6
timestamp 1731220378
transform 1 0 344 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_594_6
timestamp 1731220378
transform 1 0 528 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_593_6
timestamp 1731220378
transform 1 0 480 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_592_6
timestamp 1731220378
transform 1 0 432 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_591_6
timestamp 1731220378
transform 1 0 384 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_590_6
timestamp 1731220378
transform 1 0 336 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_589_6
timestamp 1731220378
transform 1 0 288 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_588_6
timestamp 1731220378
transform 1 0 248 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_587_6
timestamp 1731220378
transform 1 0 304 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_586_6
timestamp 1731220378
transform 1 0 408 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_585_6
timestamp 1731220378
transform 1 0 352 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_584_6
timestamp 1731220378
transform 1 0 344 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_583_6
timestamp 1731220378
transform 1 0 296 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_582_6
timestamp 1731220378
transform 1 0 248 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_581_6
timestamp 1731220378
transform 1 0 392 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_580_6
timestamp 1731220378
transform 1 0 336 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_579_6
timestamp 1731220378
transform 1 0 280 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_578_6
timestamp 1731220378
transform 1 0 224 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_577_6
timestamp 1731220378
transform 1 0 392 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_576_6
timestamp 1731220378
transform 1 0 320 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_575_6
timestamp 1731220378
transform 1 0 248 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_574_6
timestamp 1731220378
transform 1 0 240 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_573_6
timestamp 1731220378
transform 1 0 312 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_572_6
timestamp 1731220378
transform 1 0 384 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_571_6
timestamp 1731220378
transform 1 0 632 0 -1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_570_6
timestamp 1731220378
transform 1 0 520 0 -1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_569_6
timestamp 1731220378
transform 1 0 408 0 -1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_568_6
timestamp 1731220378
transform 1 0 296 0 -1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_567_6
timestamp 1731220378
transform 1 0 240 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_566_6
timestamp 1731220378
transform 1 0 304 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_565_6
timestamp 1731220378
transform 1 0 368 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_564_6
timestamp 1731220378
transform 1 0 384 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_563_6
timestamp 1731220378
transform 1 0 320 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_562_6
timestamp 1731220378
transform 1 0 248 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_561_6
timestamp 1731220378
transform 1 0 280 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_560_6
timestamp 1731220378
transform 1 0 344 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_559_6
timestamp 1731220378
transform 1 0 304 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_558_6
timestamp 1731220378
transform 1 0 256 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_557_6
timestamp 1731220378
transform 1 0 352 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_556_6
timestamp 1731220378
transform 1 0 408 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_555_6
timestamp 1731220378
transform 1 0 352 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_554_6
timestamp 1731220378
transform 1 0 296 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_553_6
timestamp 1731220378
transform 1 0 248 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_552_6
timestamp 1731220378
transform 1 0 496 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_551_6
timestamp 1731220378
transform 1 0 440 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_550_6
timestamp 1731220378
transform 1 0 384 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_549_6
timestamp 1731220378
transform 1 0 352 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_548_6
timestamp 1731220378
transform 1 0 320 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_547_6
timestamp 1731220378
transform 1 0 376 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_546_6
timestamp 1731220378
transform 1 0 320 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_545_6
timestamp 1731220378
transform 1 0 264 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_544_6
timestamp 1731220378
transform 1 0 216 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_543_6
timestamp 1731220378
transform 1 0 176 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_542_6
timestamp 1731220378
transform 1 0 144 0 1 1076
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_541_6
timestamp 1731220378
transform 1 0 288 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_540_6
timestamp 1731220378
transform 1 0 256 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_539_6
timestamp 1731220378
transform 1 0 224 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_538_6
timestamp 1731220378
transform 1 0 192 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_537_6
timestamp 1731220378
transform 1 0 160 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_536_6
timestamp 1731220378
transform 1 0 128 0 -1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_535_6
timestamp 1731220378
transform 1 0 136 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_534_6
timestamp 1731220378
transform 1 0 168 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_533_6
timestamp 1731220378
transform 1 0 208 0 1 1148
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_532_6
timestamp 1731220378
transform 1 0 208 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_531_6
timestamp 1731220378
transform 1 0 168 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_530_6
timestamp 1731220378
transform 1 0 136 0 -1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_529_6
timestamp 1731220378
transform 1 0 128 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_528_6
timestamp 1731220378
transform 1 0 168 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_527_6
timestamp 1731220378
transform 1 0 224 0 1 1220
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_526_6
timestamp 1731220378
transform 1 0 184 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_525_6
timestamp 1731220378
transform 1 0 128 0 -1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_524_6
timestamp 1731220378
transform 1 0 128 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_523_6
timestamp 1731220378
transform 1 0 176 0 1 1292
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_522_6
timestamp 1731220378
transform 1 0 208 0 -1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_521_6
timestamp 1731220378
transform 1 0 160 0 -1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_520_6
timestamp 1731220378
transform 1 0 128 0 -1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_519_6
timestamp 1731220378
transform 1 0 128 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_518_6
timestamp 1731220378
transform 1 0 168 0 1 1364
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_517_6
timestamp 1731220378
transform 1 0 176 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_516_6
timestamp 1731220378
transform 1 0 128 0 -1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_515_6
timestamp 1731220378
transform 1 0 128 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_514_6
timestamp 1731220378
transform 1 0 176 0 1 1436
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_513_6
timestamp 1731220378
transform 1 0 200 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_512_6
timestamp 1731220378
transform 1 0 152 0 -1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_511_6
timestamp 1731220378
transform 1 0 152 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_510_6
timestamp 1731220378
transform 1 0 200 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_59_6
timestamp 1731220378
transform 1 0 248 0 1 1508
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_58_6
timestamp 1731220378
transform 1 0 208 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_57_6
timestamp 1731220378
transform 1 0 168 0 -1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_56_6
timestamp 1731220378
transform 1 0 288 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_55_6
timestamp 1731220378
transform 1 0 232 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_54_6
timestamp 1731220378
transform 1 0 168 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_53_6
timestamp 1731220378
transform 1 0 128 0 1 1580
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_52_6
timestamp 1731220378
transform 1 0 128 0 -1 1652
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_51_6
timestamp 1731220378
transform 1 0 160 0 -1 1652
box 8 6 28 32
use _0_0cell_0_0ginvx0  tst_50_6
timestamp 1731220378
transform 1 0 192 0 -1 1652
box 8 6 28 32
<< end >>
