magic
tech sky130l
timestamp 1731220306
<< checkpaint >>
rect -28 76 40 80
rect -28 60 64 76
rect -28 12 80 60
rect -27 6 80 12
rect -24 -8 80 6
rect -24 -21 73 -8
rect -24 -26 66 -21
rect -24 -28 61 -26
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 11 20 12
rect 15 8 16 11
rect 19 8 20 11
rect 15 6 20 8
rect 22 10 27 12
rect 22 7 23 10
rect 26 7 27 10
rect 22 6 27 7
rect 29 11 34 12
rect 29 8 30 11
rect 33 8 34 11
rect 29 6 34 8
<< ndc >>
rect 9 7 12 10
rect 16 8 19 11
rect 23 7 26 10
rect 30 8 33 11
<< ntransistor >>
rect 13 6 15 12
rect 20 6 22 12
rect 27 6 29 12
<< pdiffusion >>
rect 8 23 13 34
rect 8 20 9 23
rect 12 20 13 23
rect 8 19 13 20
rect 15 19 20 34
rect 22 27 26 34
rect 22 26 27 27
rect 22 23 23 26
rect 26 23 27 26
rect 22 19 27 23
rect 29 23 34 27
rect 29 20 30 23
rect 33 20 34 23
rect 29 19 34 20
<< pdc >>
rect 9 20 12 23
rect 23 23 26 26
rect 30 20 33 23
<< ptransistor >>
rect 13 19 15 34
rect 20 19 22 34
rect 27 19 29 27
<< polysilicon >>
rect 10 41 15 42
rect 10 38 11 41
rect 14 38 15 41
rect 10 37 15 38
rect 13 34 15 37
rect 20 41 25 42
rect 20 38 21 41
rect 24 38 25 41
rect 20 37 25 38
rect 20 34 22 37
rect 27 27 29 29
rect 13 12 15 19
rect 20 12 22 19
rect 27 16 29 19
rect 27 15 41 16
rect 27 14 37 15
rect 27 12 29 14
rect 36 12 37 14
rect 40 12 41 15
rect 36 11 41 12
rect 13 4 15 6
rect 20 4 22 6
rect 27 4 29 6
<< pc >>
rect 11 38 14 41
rect 21 38 24 41
rect 37 12 40 15
<< m1 >>
rect 4 44 8 48
rect 5 41 8 44
rect 28 41 32 44
rect 5 38 11 41
rect 14 38 15 41
rect 20 38 21 41
rect 24 40 32 41
rect 24 38 31 40
rect 44 27 48 28
rect 23 26 26 27
rect 9 23 12 24
rect 23 22 26 23
rect 30 24 48 27
rect 30 23 33 24
rect 9 17 12 20
rect 9 13 12 14
rect 16 17 19 18
rect 16 11 19 14
rect 30 11 33 20
rect 37 15 40 16
rect 37 11 40 12
rect 8 7 9 10
rect 12 7 13 10
rect 16 7 19 8
rect 23 10 26 11
rect 30 7 33 8
rect 8 4 13 7
rect 23 6 26 7
<< m2c >>
rect 23 23 26 26
rect 9 14 12 17
rect 16 14 19 17
rect 37 12 40 15
rect 9 7 12 10
rect 23 7 26 10
<< m2 >>
rect 22 26 27 27
rect 22 23 23 26
rect 26 23 27 26
rect 22 22 27 23
rect 8 17 13 18
rect 15 17 20 18
rect 8 14 9 17
rect 12 15 16 17
rect 12 14 13 15
rect 8 13 13 14
rect 15 14 16 15
rect 19 16 20 17
rect 19 15 41 16
rect 19 14 37 15
rect 15 13 20 14
rect 36 12 37 14
rect 40 12 41 15
rect 36 11 41 12
rect 8 10 27 11
rect 8 7 9 10
rect 12 7 23 10
rect 26 7 27 10
rect 8 6 27 7
<< labels >>
rlabel space 0 0 56 52 6 prboundary
rlabel ndiffusion 34 9 34 9 3 Y
rlabel pdiffusion 34 21 34 21 3 Y
rlabel ndiffusion 30 7 30 7 3 Y
rlabel ndiffusion 30 9 30 9 3 Y
rlabel ndiffusion 30 12 30 12 3 Y
rlabel pdiffusion 30 20 30 20 3 Y
rlabel pdiffusion 30 21 30 21 3 Y
rlabel pdiffusion 30 24 30 24 3 Y
rlabel polysilicon 28 28 28 28 3 _Y
rlabel polysilicon 28 5 28 5 3 _Y
rlabel ntransistor 28 7 28 7 3 _Y
rlabel polysilicon 28 13 28 13 3 _Y
rlabel polysilicon 28 15 28 15 3 _Y
rlabel polysilicon 28 16 28 16 3 _Y
rlabel polysilicon 28 17 28 17 3 _Y
rlabel ptransistor 28 20 28 20 3 _Y
rlabel ndiffusion 23 7 23 7 3 GND
rlabel ndiffusion 23 8 23 8 3 GND
rlabel ndiffusion 23 11 23 11 3 GND
rlabel ndiffusion 20 9 20 9 3 _Y
rlabel pdiffusion 23 20 23 20 3 Vdd
rlabel pdiffusion 23 28 23 28 3 Vdd
rlabel polysilicon 21 35 21 35 3 A
rlabel polysilicon 21 38 21 38 3 A
rlabel polysilicon 21 42 21 42 3 A
rlabel polysilicon 21 5 21 5 3 A
rlabel ntransistor 21 7 21 7 3 A
rlabel polysilicon 21 13 21 13 3 A
rlabel ptransistor 21 20 21 20 3 A
rlabel ndiffusion 16 7 16 7 3 _Y
rlabel ndiffusion 16 9 16 9 3 _Y
rlabel ndiffusion 16 12 16 12 3 _Y
rlabel pdiffusion 13 21 13 21 3 _Y
rlabel polysilicon 14 35 14 35 3 B
rlabel polysilicon 14 5 14 5 3 B
rlabel ntransistor 14 7 14 7 3 B
rlabel polysilicon 14 13 14 13 3 B
rlabel ptransistor 14 20 14 20 3 B
rlabel polysilicon 11 38 11 38 3 B
rlabel polysilicon 11 39 11 39 3 B
rlabel polysilicon 11 42 11 42 3 B
rlabel pdiffusion 9 20 9 20 3 _Y
rlabel pdiffusion 9 21 9 21 3 _Y
rlabel pdiffusion 9 24 9 24 3 _Y
rlabel m1 45 28 45 28 3 Y
port 1 e
rlabel m1 38 12 38 12 3 _Y
rlabel m1 38 16 38 16 3 _Y
rlabel m1 29 42 29 42 3 A
port 2 e
rlabel ndc 31 9 31 9 3 Y
port 1 e
rlabel m1 31 12 31 12 3 Y
port 1 e
rlabel pdc 31 21 31 21 3 Y
port 1 e
rlabel m1 31 24 31 24 3 Y
port 1 e
rlabel m1 31 25 31 25 3 Y
port 1 e
rlabel m1 31 8 31 8 3 Y
port 1 e
rlabel m1 24 11 24 11 3 GND
rlabel m1 24 23 24 23 3 Vdd
rlabel m1 24 27 24 27 3 Vdd
rlabel m1 25 39 25 39 3 A
port 2 e
rlabel m1 25 41 25 41 3 A
port 2 e
rlabel pc 22 39 22 39 3 A
port 2 e
rlabel m1 21 39 21 39 3 A
port 2 e
rlabel m1 17 8 17 8 3 _Y
rlabel ndc 17 9 17 9 3 _Y
rlabel m1 17 12 17 12 3 _Y
rlabel m1 17 18 17 18 3 _Y
rlabel m1 24 7 24 7 3 GND
rlabel m1 10 14 10 14 3 _Y
rlabel m1 10 18 10 18 3 _Y
rlabel pdc 10 21 10 21 3 _Y
rlabel m1 10 24 10 24 3 _Y
rlabel m1 15 39 15 39 3 B
port 3 e
rlabel m1 9 5 9 5 3 GND
rlabel pc 12 39 12 39 3 B
port 3 e
rlabel m1 6 39 6 39 3 B
port 3 e
rlabel m1 6 42 6 42 3 B
port 3 e
rlabel m1 5 45 5 45 3 B
port 3 e
rlabel m2 20 15 20 15 3 _Y
rlabel m2 20 16 20 16 3 _Y
rlabel m2 20 17 20 17 3 _Y
rlabel m2 27 24 27 24 3 Vdd
rlabel m2c 17 15 17 15 3 _Y
rlabel m2c 24 24 24 24 3 Vdd
rlabel m2 27 8 27 8 3 GND
rlabel m2 41 13 41 13 3 _Y
rlabel m2 16 15 16 15 3 _Y
rlabel m2 23 23 23 23 3 Vdd
rlabel m2 23 24 23 24 3 Vdd
rlabel m2 23 27 23 27 3 Vdd
rlabel m2c 24 8 24 8 3 GND
rlabel m2c 38 13 38 13 3 _Y
rlabel m2 13 8 13 8 3 GND
rlabel m2 37 12 37 12 3 _Y
rlabel m2 37 13 37 13 3 _Y
rlabel m2 16 14 16 14 3 _Y
rlabel m2 13 15 13 15 3 _Y
rlabel m2 13 16 13 16 3 _Y
rlabel m2 16 18 16 18 3 _Y
rlabel m2c 10 8 10 8 3 GND
rlabel m2c 10 15 10 15 3 _Y
rlabel m2 9 7 9 7 3 GND
rlabel m2 9 8 9 8 3 GND
rlabel m2 9 11 9 11 3 GND
rlabel m2 9 14 9 14 3 _Y
rlabel m2 9 15 9 15 3 _Y
rlabel m2 9 18 9 18 3 _Y
<< end >>
