magic
tech sky130l
timestamp 1730767052
<< m1 >>
rect 1104 483 1108 543
<< m2c >>
rect 608 1511 612 1515
rect 696 1511 700 1515
rect 784 1511 788 1515
rect 872 1511 876 1515
rect 960 1511 964 1515
rect 111 1497 115 1501
rect 1567 1497 1571 1501
rect 111 1479 115 1483
rect 1567 1479 1571 1483
rect 111 1445 115 1449
rect 1567 1445 1571 1449
rect 656 1439 660 1443
rect 816 1439 820 1443
rect 1160 1439 1164 1443
rect 111 1427 115 1431
rect 1567 1427 1571 1431
rect 536 1411 540 1415
rect 680 1411 684 1415
rect 840 1411 844 1415
rect 1008 1411 1012 1415
rect 1184 1411 1188 1415
rect 1536 1411 1540 1415
rect 488 1383 492 1387
rect 728 1379 732 1383
rect 976 1379 980 1383
rect 1232 1379 1236 1383
rect 1496 1381 1500 1385
rect 111 1365 115 1369
rect 1567 1365 1571 1369
rect 111 1347 115 1351
rect 1567 1347 1571 1351
rect 111 1301 115 1305
rect 1567 1301 1571 1305
rect 768 1295 772 1299
rect 1504 1295 1508 1299
rect 111 1283 115 1287
rect 1567 1283 1571 1287
rect 552 1267 556 1271
rect 792 1267 796 1271
rect 1032 1267 1036 1271
rect 1280 1267 1284 1271
rect 1528 1267 1532 1271
rect 600 1231 604 1235
rect 1464 1231 1468 1235
rect 808 1227 812 1231
rect 1024 1227 1028 1231
rect 1240 1227 1244 1231
rect 111 1213 115 1217
rect 1567 1213 1571 1217
rect 111 1195 115 1199
rect 1567 1195 1571 1199
rect 111 1145 115 1149
rect 1567 1145 1571 1149
rect 872 1139 876 1143
rect 1056 1139 1060 1143
rect 111 1127 115 1131
rect 1567 1127 1571 1131
rect 720 1111 724 1115
rect 896 1111 900 1115
rect 1080 1111 1084 1115
rect 1272 1111 1276 1115
rect 1464 1111 1468 1115
rect 728 1075 732 1079
rect 1488 1075 1492 1079
rect 912 1071 916 1075
rect 1096 1071 1100 1075
rect 1288 1071 1292 1075
rect 111 1057 115 1061
rect 1567 1057 1571 1061
rect 111 1039 115 1043
rect 1567 1039 1571 1043
rect 111 989 115 993
rect 1567 989 1571 993
rect 800 983 804 987
rect 111 971 115 975
rect 1567 971 1571 975
rect 616 955 620 959
rect 824 955 828 959
rect 1040 955 1044 959
rect 1264 955 1268 959
rect 1496 955 1500 959
rect 464 919 468 923
rect 728 919 732 923
rect 992 919 996 923
rect 1536 919 1540 923
rect 1264 915 1268 919
rect 111 901 115 905
rect 1567 901 1571 905
rect 111 883 115 887
rect 1567 883 1571 887
rect 111 837 115 841
rect 1567 837 1571 841
rect 576 831 580 835
rect 864 831 868 835
rect 111 819 115 823
rect 1567 819 1571 823
rect 320 803 324 807
rect 600 803 604 807
rect 888 803 892 807
rect 1176 803 1180 807
rect 1472 803 1476 807
rect 264 767 268 771
rect 1464 767 1468 771
rect 552 763 556 767
rect 848 763 852 767
rect 1152 763 1156 767
rect 111 749 115 753
rect 1567 749 1571 753
rect 111 731 115 735
rect 1567 731 1571 735
rect 111 689 115 693
rect 1567 689 1571 693
rect 111 671 115 675
rect 1567 671 1571 675
rect 320 655 324 659
rect 592 655 596 659
rect 880 655 884 659
rect 1176 655 1180 659
rect 1472 655 1476 659
rect 824 627 828 631
rect 1040 627 1044 631
rect 1480 627 1484 631
rect 616 623 620 627
rect 1256 623 1260 627
rect 111 609 115 613
rect 1567 609 1571 613
rect 111 591 115 595
rect 1567 591 1571 595
rect 111 549 115 553
rect 1567 549 1571 553
rect 1104 543 1108 547
rect 1152 543 1156 547
rect 111 531 115 535
rect 792 515 796 519
rect 912 515 916 519
rect 1040 515 1044 519
rect 1567 531 1571 535
rect 1176 515 1180 519
rect 1320 515 1324 519
rect 1472 515 1476 519
rect 1096 479 1100 483
rect 1104 479 1108 483
rect 1536 479 1540 483
rect 832 475 836 479
rect 920 475 924 479
rect 1008 475 1012 479
rect 1184 475 1188 479
rect 1272 475 1276 479
rect 1360 475 1364 479
rect 1448 475 1452 479
rect 111 461 115 465
rect 1567 461 1571 465
rect 111 443 115 447
rect 1567 443 1571 447
rect 111 393 115 397
rect 1567 393 1571 397
rect 752 387 756 391
rect 840 387 844 391
rect 111 375 115 379
rect 1567 375 1571 379
rect 688 359 692 363
rect 776 359 780 363
rect 864 359 868 363
rect 952 359 956 363
rect 728 319 732 323
rect 464 315 468 319
rect 552 315 556 319
rect 640 315 644 319
rect 111 301 115 305
rect 1567 301 1571 305
rect 111 283 115 287
rect 1567 283 1571 287
rect 111 229 115 233
rect 1567 229 1571 233
rect 344 223 348 227
rect 432 223 436 227
rect 520 223 524 227
rect 111 211 115 215
rect 1567 211 1571 215
rect 280 195 284 199
rect 368 195 372 199
rect 456 195 460 199
rect 544 195 548 199
rect 640 139 644 143
rect 200 135 204 139
rect 288 135 292 139
rect 376 135 380 139
rect 464 135 468 139
rect 552 135 556 139
rect 111 121 115 125
rect 1567 121 1571 125
rect 111 103 115 107
rect 1567 103 1571 107
<< m2 >>
rect 542 1518 548 1519
rect 542 1514 543 1518
rect 547 1514 548 1518
rect 630 1518 636 1519
rect 542 1513 548 1514
rect 607 1515 613 1516
rect 607 1511 608 1515
rect 612 1514 613 1515
rect 630 1514 631 1518
rect 635 1514 636 1518
rect 718 1518 724 1519
rect 612 1512 626 1514
rect 630 1513 636 1514
rect 695 1515 701 1516
rect 612 1511 613 1512
rect 607 1510 613 1511
rect 624 1506 626 1512
rect 695 1511 696 1515
rect 700 1514 701 1515
rect 718 1514 719 1518
rect 723 1514 724 1518
rect 806 1518 812 1519
rect 700 1512 714 1514
rect 718 1513 724 1514
rect 783 1515 789 1516
rect 700 1511 701 1512
rect 695 1510 701 1511
rect 646 1507 652 1508
rect 646 1506 647 1507
rect 624 1504 647 1506
rect 646 1503 647 1504
rect 651 1503 652 1507
rect 712 1506 714 1512
rect 783 1511 784 1515
rect 788 1514 789 1515
rect 806 1514 807 1518
rect 811 1514 812 1518
rect 894 1518 900 1519
rect 788 1512 802 1514
rect 806 1513 812 1514
rect 871 1515 877 1516
rect 788 1511 789 1512
rect 783 1510 789 1511
rect 734 1507 740 1508
rect 734 1506 735 1507
rect 712 1504 735 1506
rect 646 1502 652 1503
rect 734 1503 735 1504
rect 739 1503 740 1507
rect 800 1506 802 1512
rect 871 1511 872 1515
rect 876 1514 877 1515
rect 886 1515 892 1516
rect 886 1514 887 1515
rect 876 1512 887 1514
rect 876 1511 877 1512
rect 871 1510 877 1511
rect 886 1511 887 1512
rect 891 1511 892 1515
rect 894 1514 895 1518
rect 899 1514 900 1518
rect 894 1513 900 1514
rect 959 1515 965 1516
rect 886 1510 892 1511
rect 959 1511 960 1515
rect 964 1514 965 1515
rect 974 1515 980 1516
rect 974 1514 975 1515
rect 964 1512 975 1514
rect 964 1511 965 1512
rect 959 1510 965 1511
rect 974 1511 975 1512
rect 979 1511 980 1515
rect 974 1510 980 1511
rect 822 1507 828 1508
rect 822 1506 823 1507
rect 800 1504 823 1506
rect 734 1502 740 1503
rect 822 1503 823 1504
rect 827 1503 828 1507
rect 822 1502 828 1503
rect 110 1501 116 1502
rect 110 1497 111 1501
rect 115 1497 116 1501
rect 110 1496 116 1497
rect 1566 1501 1572 1502
rect 1566 1497 1567 1501
rect 1571 1497 1572 1501
rect 1566 1496 1572 1497
rect 886 1487 892 1488
rect 110 1483 116 1484
rect 110 1479 111 1483
rect 115 1479 116 1483
rect 886 1483 887 1487
rect 891 1486 892 1487
rect 891 1484 962 1486
rect 891 1483 892 1484
rect 886 1482 892 1483
rect 110 1478 116 1479
rect 960 1473 962 1484
rect 1566 1483 1572 1484
rect 1566 1479 1567 1483
rect 1571 1479 1572 1483
rect 1566 1478 1572 1479
rect 542 1472 548 1473
rect 630 1472 636 1473
rect 718 1472 724 1473
rect 806 1472 812 1473
rect 894 1472 900 1473
rect 542 1468 543 1472
rect 547 1468 548 1472
rect 622 1471 628 1472
rect 622 1470 623 1471
rect 613 1468 623 1470
rect 542 1467 548 1468
rect 622 1467 623 1468
rect 627 1467 628 1471
rect 630 1468 631 1472
rect 635 1468 636 1472
rect 630 1467 636 1468
rect 646 1471 652 1472
rect 646 1467 647 1471
rect 651 1470 652 1471
rect 651 1468 665 1470
rect 718 1468 719 1472
rect 723 1468 724 1472
rect 651 1467 652 1468
rect 718 1467 724 1468
rect 734 1471 740 1472
rect 734 1467 735 1471
rect 739 1470 740 1471
rect 739 1468 753 1470
rect 806 1468 807 1472
rect 811 1468 812 1472
rect 739 1467 740 1468
rect 806 1467 812 1468
rect 822 1471 828 1472
rect 822 1467 823 1471
rect 827 1470 828 1471
rect 827 1468 841 1470
rect 894 1468 895 1472
rect 899 1468 900 1472
rect 827 1467 828 1468
rect 894 1467 900 1468
rect 622 1466 628 1467
rect 646 1466 652 1467
rect 734 1466 740 1467
rect 822 1466 828 1467
rect 470 1460 476 1461
rect 614 1460 620 1461
rect 470 1456 471 1460
rect 475 1456 476 1460
rect 470 1455 476 1456
rect 502 1459 508 1460
rect 502 1455 503 1459
rect 507 1455 508 1459
rect 614 1456 615 1460
rect 619 1456 620 1460
rect 614 1455 620 1456
rect 774 1460 780 1461
rect 774 1456 775 1460
rect 779 1456 780 1460
rect 774 1455 780 1456
rect 942 1460 948 1461
rect 1118 1460 1124 1461
rect 942 1456 943 1460
rect 947 1456 948 1460
rect 942 1455 948 1456
rect 974 1459 980 1460
rect 974 1455 975 1459
rect 979 1455 980 1459
rect 1118 1456 1119 1460
rect 1123 1456 1124 1460
rect 1118 1455 1124 1456
rect 1302 1460 1308 1461
rect 1470 1460 1476 1461
rect 1302 1456 1303 1460
rect 1307 1456 1308 1460
rect 1434 1459 1440 1460
rect 1434 1458 1435 1459
rect 1373 1456 1435 1458
rect 1302 1455 1308 1456
rect 1434 1455 1435 1456
rect 1439 1455 1440 1459
rect 1470 1456 1471 1460
rect 1475 1456 1476 1460
rect 1470 1455 1476 1456
rect 1494 1459 1500 1460
rect 1494 1455 1495 1459
rect 1499 1458 1500 1459
rect 1499 1456 1505 1458
rect 1499 1455 1500 1456
rect 502 1454 508 1455
rect 974 1454 980 1455
rect 1434 1454 1440 1455
rect 1494 1454 1500 1455
rect 110 1449 116 1450
rect 110 1445 111 1449
rect 115 1445 116 1449
rect 110 1444 116 1445
rect 1566 1449 1572 1450
rect 1566 1445 1567 1449
rect 1571 1445 1572 1449
rect 1566 1444 1572 1445
rect 538 1443 544 1444
rect 538 1439 539 1443
rect 543 1442 544 1443
rect 655 1443 661 1444
rect 655 1442 656 1443
rect 543 1440 656 1442
rect 543 1439 544 1440
rect 538 1438 544 1439
rect 655 1439 656 1440
rect 660 1439 661 1443
rect 655 1438 661 1439
rect 682 1443 688 1444
rect 682 1439 683 1443
rect 687 1442 688 1443
rect 815 1443 821 1444
rect 815 1442 816 1443
rect 687 1440 816 1442
rect 687 1439 688 1440
rect 682 1438 688 1439
rect 815 1439 816 1440
rect 820 1439 821 1443
rect 815 1438 821 1439
rect 1010 1443 1016 1444
rect 1010 1439 1011 1443
rect 1015 1442 1016 1443
rect 1159 1443 1165 1444
rect 1159 1442 1160 1443
rect 1015 1440 1160 1442
rect 1015 1439 1016 1440
rect 1010 1438 1016 1439
rect 1159 1439 1160 1440
rect 1164 1439 1165 1443
rect 1159 1438 1165 1439
rect 110 1431 116 1432
rect 110 1427 111 1431
rect 115 1427 116 1431
rect 110 1426 116 1427
rect 1566 1431 1572 1432
rect 1566 1427 1567 1431
rect 1571 1427 1572 1431
rect 1566 1426 1572 1427
rect 1434 1423 1440 1424
rect 1434 1419 1435 1423
rect 1439 1422 1440 1423
rect 1439 1420 1498 1422
rect 1439 1419 1440 1420
rect 1434 1418 1440 1419
rect 535 1415 544 1416
rect 679 1415 688 1416
rect 839 1415 845 1416
rect 1007 1415 1016 1416
rect 1183 1415 1189 1416
rect 470 1414 476 1415
rect 470 1410 471 1414
rect 475 1410 476 1414
rect 535 1411 536 1415
rect 543 1411 544 1415
rect 535 1410 544 1411
rect 614 1414 620 1415
rect 614 1410 615 1414
rect 619 1410 620 1414
rect 679 1411 680 1415
rect 687 1411 688 1415
rect 679 1410 688 1411
rect 774 1414 780 1415
rect 839 1414 840 1415
rect 774 1410 775 1414
rect 779 1410 780 1414
rect 470 1409 476 1410
rect 614 1409 620 1410
rect 774 1409 780 1410
rect 800 1412 840 1414
rect 622 1407 628 1408
rect 622 1403 623 1407
rect 627 1406 628 1407
rect 800 1406 802 1412
rect 839 1411 840 1412
rect 844 1411 845 1415
rect 839 1410 845 1411
rect 942 1414 948 1415
rect 942 1410 943 1414
rect 947 1410 948 1414
rect 1007 1411 1008 1415
rect 1015 1411 1016 1415
rect 1007 1410 1016 1411
rect 1118 1414 1124 1415
rect 1118 1410 1119 1414
rect 1123 1410 1124 1414
rect 1183 1411 1184 1415
rect 1188 1414 1189 1415
rect 1198 1415 1204 1416
rect 1198 1414 1199 1415
rect 1188 1412 1199 1414
rect 1188 1411 1189 1412
rect 1183 1410 1189 1411
rect 1198 1411 1199 1412
rect 1203 1411 1204 1415
rect 1198 1410 1204 1411
rect 1302 1414 1308 1415
rect 1302 1410 1303 1414
rect 1307 1410 1308 1414
rect 942 1409 948 1410
rect 1118 1409 1124 1410
rect 1302 1409 1308 1410
rect 1470 1414 1476 1415
rect 1470 1410 1471 1414
rect 1475 1410 1476 1414
rect 1496 1414 1498 1420
rect 1535 1415 1541 1416
rect 1535 1414 1536 1415
rect 1496 1412 1536 1414
rect 1535 1411 1536 1412
rect 1540 1411 1541 1415
rect 1535 1410 1541 1411
rect 1470 1409 1476 1410
rect 627 1404 802 1406
rect 627 1403 628 1404
rect 622 1402 628 1403
rect 487 1387 493 1388
rect 422 1386 428 1387
rect 422 1382 423 1386
rect 427 1382 428 1386
rect 487 1383 488 1387
rect 492 1386 493 1387
rect 502 1387 508 1388
rect 1494 1387 1500 1388
rect 502 1386 503 1387
rect 492 1384 503 1386
rect 492 1383 493 1384
rect 487 1382 493 1383
rect 502 1383 503 1384
rect 507 1383 508 1387
rect 502 1382 508 1383
rect 662 1386 668 1387
rect 662 1382 663 1386
rect 667 1382 668 1386
rect 910 1386 916 1387
rect 727 1383 733 1384
rect 727 1382 728 1383
rect 422 1381 428 1382
rect 662 1381 668 1382
rect 688 1380 728 1382
rect 590 1375 596 1376
rect 590 1371 591 1375
rect 595 1374 596 1375
rect 688 1374 690 1380
rect 727 1379 728 1380
rect 732 1379 733 1383
rect 910 1382 911 1386
rect 915 1382 916 1386
rect 1166 1386 1172 1387
rect 910 1381 916 1382
rect 975 1383 984 1384
rect 727 1378 733 1379
rect 975 1379 976 1383
rect 983 1379 984 1383
rect 1166 1382 1167 1386
rect 1171 1382 1172 1386
rect 1430 1386 1436 1387
rect 1166 1381 1172 1382
rect 1206 1383 1212 1384
rect 975 1378 984 1379
rect 1206 1379 1207 1383
rect 1211 1382 1212 1383
rect 1231 1383 1237 1384
rect 1231 1382 1232 1383
rect 1211 1380 1232 1382
rect 1211 1379 1212 1380
rect 1206 1378 1212 1379
rect 1231 1379 1232 1380
rect 1236 1379 1237 1383
rect 1430 1382 1431 1386
rect 1435 1382 1436 1386
rect 1494 1383 1495 1387
rect 1499 1386 1500 1387
rect 1499 1385 1501 1386
rect 1494 1382 1496 1383
rect 1430 1381 1436 1382
rect 1495 1381 1496 1382
rect 1500 1381 1501 1385
rect 1495 1380 1501 1381
rect 1231 1378 1237 1379
rect 595 1372 690 1374
rect 595 1371 596 1372
rect 590 1370 596 1371
rect 110 1369 116 1370
rect 110 1365 111 1369
rect 115 1365 116 1369
rect 110 1364 116 1365
rect 1566 1369 1572 1370
rect 1566 1365 1567 1369
rect 1571 1365 1572 1369
rect 1566 1364 1572 1365
rect 730 1359 736 1360
rect 730 1355 731 1359
rect 735 1358 736 1359
rect 978 1359 984 1360
rect 978 1358 979 1359
rect 735 1356 979 1358
rect 735 1355 736 1356
rect 730 1354 736 1355
rect 978 1355 979 1356
rect 983 1355 984 1359
rect 978 1354 984 1355
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 110 1346 116 1347
rect 1566 1351 1572 1352
rect 1566 1347 1567 1351
rect 1571 1347 1572 1351
rect 1566 1346 1572 1347
rect 730 1343 736 1344
rect 422 1340 428 1341
rect 662 1340 668 1341
rect 422 1336 423 1340
rect 427 1336 428 1340
rect 590 1339 596 1340
rect 590 1338 591 1339
rect 493 1336 591 1338
rect 422 1335 428 1336
rect 590 1335 591 1336
rect 595 1335 596 1339
rect 662 1336 663 1340
rect 667 1336 668 1340
rect 730 1339 731 1343
rect 735 1339 736 1343
rect 730 1338 736 1339
rect 910 1340 916 1341
rect 662 1335 668 1336
rect 910 1336 911 1340
rect 915 1336 916 1340
rect 1166 1340 1172 1341
rect 1430 1340 1436 1341
rect 910 1335 916 1336
rect 590 1334 596 1335
rect 854 1331 860 1332
rect 854 1327 855 1331
rect 859 1330 860 1331
rect 944 1330 946 1337
rect 1166 1336 1167 1340
rect 1171 1336 1172 1340
rect 1166 1335 1172 1336
rect 1198 1339 1204 1340
rect 1198 1335 1199 1339
rect 1203 1335 1204 1339
rect 1430 1336 1431 1340
rect 1435 1336 1436 1340
rect 1430 1335 1436 1336
rect 1498 1339 1504 1340
rect 1498 1335 1499 1339
rect 1503 1335 1504 1339
rect 1198 1334 1204 1335
rect 1498 1334 1504 1335
rect 859 1328 946 1330
rect 859 1327 860 1328
rect 854 1326 860 1327
rect 486 1316 492 1317
rect 726 1316 732 1317
rect 486 1312 487 1316
rect 491 1312 492 1316
rect 562 1315 568 1316
rect 562 1314 563 1315
rect 557 1312 563 1314
rect 486 1311 492 1312
rect 562 1311 563 1312
rect 567 1311 568 1315
rect 726 1312 727 1316
rect 731 1312 732 1316
rect 726 1311 732 1312
rect 966 1316 972 1317
rect 1214 1316 1220 1317
rect 1462 1316 1468 1317
rect 966 1312 967 1316
rect 971 1312 972 1316
rect 1206 1315 1212 1316
rect 1206 1314 1207 1315
rect 1037 1312 1207 1314
rect 966 1311 972 1312
rect 1206 1311 1207 1312
rect 1211 1311 1212 1315
rect 1214 1312 1215 1316
rect 1219 1312 1220 1316
rect 1422 1315 1428 1316
rect 1422 1314 1423 1315
rect 1285 1312 1423 1314
rect 1214 1311 1220 1312
rect 1422 1311 1423 1312
rect 1427 1311 1428 1315
rect 1462 1312 1463 1316
rect 1467 1312 1468 1316
rect 1462 1311 1468 1312
rect 562 1310 568 1311
rect 1206 1310 1212 1311
rect 1422 1310 1428 1311
rect 110 1305 116 1306
rect 110 1301 111 1305
rect 115 1301 116 1305
rect 110 1300 116 1301
rect 1566 1305 1572 1306
rect 1566 1301 1567 1305
rect 1571 1301 1572 1305
rect 1566 1300 1572 1301
rect 554 1299 560 1300
rect 554 1295 555 1299
rect 559 1298 560 1299
rect 767 1299 773 1300
rect 767 1298 768 1299
rect 559 1296 768 1298
rect 559 1295 560 1296
rect 554 1294 560 1295
rect 767 1295 768 1296
rect 772 1295 773 1299
rect 767 1294 773 1295
rect 1282 1299 1288 1300
rect 1282 1295 1283 1299
rect 1287 1298 1288 1299
rect 1503 1299 1509 1300
rect 1503 1298 1504 1299
rect 1287 1296 1504 1298
rect 1287 1295 1288 1296
rect 1282 1294 1288 1295
rect 1503 1295 1504 1296
rect 1508 1295 1509 1299
rect 1503 1294 1509 1295
rect 110 1287 116 1288
rect 110 1283 111 1287
rect 115 1283 116 1287
rect 110 1282 116 1283
rect 1566 1287 1572 1288
rect 1566 1283 1567 1287
rect 1571 1283 1572 1287
rect 1566 1282 1572 1283
rect 551 1271 560 1272
rect 791 1271 797 1272
rect 486 1270 492 1271
rect 486 1266 487 1270
rect 491 1266 492 1270
rect 551 1267 552 1271
rect 559 1267 560 1271
rect 551 1266 560 1267
rect 726 1270 732 1271
rect 726 1266 727 1270
rect 731 1266 732 1270
rect 791 1267 792 1271
rect 796 1270 797 1271
rect 854 1271 860 1272
rect 1031 1271 1037 1272
rect 854 1270 855 1271
rect 796 1268 855 1270
rect 796 1267 797 1268
rect 791 1266 797 1267
rect 854 1267 855 1268
rect 859 1267 860 1271
rect 854 1266 860 1267
rect 966 1270 972 1271
rect 966 1266 967 1270
rect 971 1266 972 1270
rect 1031 1267 1032 1271
rect 1036 1270 1037 1271
rect 1206 1271 1212 1272
rect 1279 1271 1288 1272
rect 1498 1271 1504 1272
rect 1206 1270 1207 1271
rect 1036 1268 1207 1270
rect 1036 1267 1037 1268
rect 1031 1266 1037 1267
rect 1206 1267 1207 1268
rect 1211 1267 1212 1271
rect 1206 1266 1212 1267
rect 1214 1270 1220 1271
rect 1214 1266 1215 1270
rect 1219 1266 1220 1270
rect 1279 1267 1280 1271
rect 1287 1267 1288 1271
rect 1279 1266 1288 1267
rect 1462 1270 1468 1271
rect 1462 1266 1463 1270
rect 1467 1266 1468 1270
rect 1498 1267 1499 1271
rect 1503 1270 1504 1271
rect 1527 1271 1533 1272
rect 1527 1270 1528 1271
rect 1503 1268 1528 1270
rect 1503 1267 1504 1268
rect 1498 1266 1504 1267
rect 1527 1267 1528 1268
rect 1532 1267 1533 1271
rect 1527 1266 1533 1267
rect 486 1265 492 1266
rect 726 1265 732 1266
rect 966 1265 972 1266
rect 1214 1265 1220 1266
rect 1462 1265 1468 1266
rect 562 1235 568 1236
rect 534 1234 540 1235
rect 534 1230 535 1234
rect 539 1230 540 1234
rect 562 1231 563 1235
rect 567 1234 568 1235
rect 599 1235 605 1236
rect 1422 1235 1428 1236
rect 599 1234 600 1235
rect 567 1232 600 1234
rect 567 1231 568 1232
rect 562 1230 568 1231
rect 599 1231 600 1232
rect 604 1231 605 1235
rect 599 1230 605 1231
rect 742 1234 748 1235
rect 742 1230 743 1234
rect 747 1230 748 1234
rect 958 1234 964 1235
rect 807 1231 813 1232
rect 807 1230 808 1231
rect 534 1229 540 1230
rect 742 1229 748 1230
rect 768 1228 808 1230
rect 686 1223 692 1224
rect 686 1219 687 1223
rect 691 1222 692 1223
rect 768 1222 770 1228
rect 807 1227 808 1228
rect 812 1227 813 1231
rect 958 1230 959 1234
rect 963 1230 964 1234
rect 1174 1234 1180 1235
rect 958 1229 964 1230
rect 982 1231 988 1232
rect 807 1226 813 1227
rect 982 1227 983 1231
rect 987 1230 988 1231
rect 1023 1231 1029 1232
rect 1023 1230 1024 1231
rect 987 1228 1024 1230
rect 987 1227 988 1228
rect 982 1226 988 1227
rect 1023 1227 1024 1228
rect 1028 1227 1029 1231
rect 1174 1230 1175 1234
rect 1179 1230 1180 1234
rect 1398 1234 1404 1235
rect 1174 1229 1180 1230
rect 1238 1231 1245 1232
rect 1023 1226 1029 1227
rect 1238 1227 1239 1231
rect 1244 1227 1245 1231
rect 1398 1230 1399 1234
rect 1403 1230 1404 1234
rect 1422 1231 1423 1235
rect 1427 1234 1428 1235
rect 1463 1235 1469 1236
rect 1463 1234 1464 1235
rect 1427 1232 1464 1234
rect 1427 1231 1428 1232
rect 1422 1230 1428 1231
rect 1463 1231 1464 1232
rect 1468 1231 1469 1235
rect 1463 1230 1469 1231
rect 1398 1229 1404 1230
rect 1238 1226 1245 1227
rect 691 1220 770 1222
rect 691 1219 692 1220
rect 686 1218 692 1219
rect 110 1217 116 1218
rect 110 1213 111 1217
rect 115 1213 116 1217
rect 110 1212 116 1213
rect 1566 1217 1572 1218
rect 1566 1213 1567 1217
rect 1571 1213 1572 1217
rect 1566 1212 1572 1213
rect 110 1199 116 1200
rect 110 1195 111 1199
rect 115 1195 116 1199
rect 110 1194 116 1195
rect 1566 1199 1572 1200
rect 1566 1195 1567 1199
rect 1571 1195 1572 1199
rect 1566 1194 1572 1195
rect 534 1188 540 1189
rect 742 1188 748 1189
rect 534 1184 535 1188
rect 539 1184 540 1188
rect 686 1187 692 1188
rect 686 1186 687 1187
rect 605 1184 687 1186
rect 534 1183 540 1184
rect 686 1183 687 1184
rect 691 1183 692 1187
rect 742 1184 743 1188
rect 747 1184 748 1188
rect 958 1188 964 1189
rect 1174 1188 1180 1189
rect 1398 1188 1404 1189
rect 813 1184 850 1186
rect 742 1183 748 1184
rect 686 1182 692 1183
rect 848 1178 850 1184
rect 958 1184 959 1188
rect 963 1184 964 1188
rect 1038 1187 1044 1188
rect 1038 1186 1039 1187
rect 1029 1184 1039 1186
rect 958 1183 964 1184
rect 1038 1183 1039 1184
rect 1043 1183 1044 1187
rect 1174 1184 1175 1188
rect 1179 1184 1180 1188
rect 1174 1183 1180 1184
rect 1206 1187 1212 1188
rect 1206 1183 1207 1187
rect 1211 1183 1212 1187
rect 1398 1184 1399 1188
rect 1403 1184 1404 1188
rect 1398 1183 1404 1184
rect 1462 1187 1468 1188
rect 1462 1183 1463 1187
rect 1467 1183 1468 1187
rect 1038 1182 1044 1183
rect 1206 1182 1212 1183
rect 1462 1182 1468 1183
rect 982 1179 988 1180
rect 982 1178 983 1179
rect 848 1176 983 1178
rect 982 1175 983 1176
rect 987 1175 988 1179
rect 982 1174 988 1175
rect 654 1160 660 1161
rect 830 1160 836 1161
rect 654 1156 655 1160
rect 659 1156 660 1160
rect 730 1159 736 1160
rect 730 1158 731 1159
rect 725 1156 731 1158
rect 654 1155 660 1156
rect 730 1155 731 1156
rect 735 1155 736 1159
rect 830 1156 831 1160
rect 835 1156 836 1160
rect 830 1155 836 1156
rect 1014 1160 1020 1161
rect 1014 1156 1015 1160
rect 1019 1156 1020 1160
rect 1014 1155 1020 1156
rect 1206 1160 1212 1161
rect 1398 1160 1404 1161
rect 1206 1156 1207 1160
rect 1211 1156 1212 1160
rect 1206 1155 1212 1156
rect 1238 1159 1244 1160
rect 1238 1155 1239 1159
rect 1243 1155 1244 1159
rect 1398 1156 1399 1160
rect 1403 1156 1404 1160
rect 1474 1159 1480 1160
rect 1474 1158 1475 1159
rect 1469 1156 1475 1158
rect 1398 1155 1404 1156
rect 1474 1155 1475 1156
rect 1479 1155 1480 1159
rect 730 1154 736 1155
rect 1238 1154 1244 1155
rect 1474 1154 1480 1155
rect 110 1149 116 1150
rect 110 1145 111 1149
rect 115 1145 116 1149
rect 110 1144 116 1145
rect 1566 1149 1572 1150
rect 1566 1145 1567 1149
rect 1571 1145 1572 1149
rect 1566 1144 1572 1145
rect 722 1143 728 1144
rect 722 1139 723 1143
rect 727 1142 728 1143
rect 871 1143 877 1144
rect 871 1142 872 1143
rect 727 1140 872 1142
rect 727 1139 728 1140
rect 722 1138 728 1139
rect 871 1139 872 1140
rect 876 1139 877 1143
rect 871 1138 877 1139
rect 954 1143 960 1144
rect 954 1139 955 1143
rect 959 1142 960 1143
rect 1055 1143 1061 1144
rect 1055 1142 1056 1143
rect 959 1140 1056 1142
rect 959 1139 960 1140
rect 954 1138 960 1139
rect 1055 1139 1056 1140
rect 1060 1139 1061 1143
rect 1055 1138 1061 1139
rect 110 1131 116 1132
rect 110 1127 111 1131
rect 115 1127 116 1131
rect 110 1126 116 1127
rect 1566 1131 1572 1132
rect 1566 1127 1567 1131
rect 1571 1127 1572 1131
rect 1566 1126 1572 1127
rect 719 1115 728 1116
rect 895 1115 901 1116
rect 654 1114 660 1115
rect 654 1110 655 1114
rect 659 1110 660 1114
rect 719 1111 720 1115
rect 727 1111 728 1115
rect 719 1110 728 1111
rect 830 1114 836 1115
rect 830 1110 831 1114
rect 835 1110 836 1114
rect 895 1111 896 1115
rect 900 1114 901 1115
rect 954 1115 960 1116
rect 1038 1115 1044 1116
rect 954 1114 955 1115
rect 900 1112 955 1114
rect 900 1111 901 1112
rect 895 1110 901 1111
rect 954 1111 955 1112
rect 959 1111 960 1115
rect 954 1110 960 1111
rect 1014 1114 1020 1115
rect 1014 1110 1015 1114
rect 1019 1110 1020 1114
rect 1038 1111 1039 1115
rect 1043 1114 1044 1115
rect 1079 1115 1085 1116
rect 1270 1115 1277 1116
rect 1462 1115 1469 1116
rect 1079 1114 1080 1115
rect 1043 1112 1080 1114
rect 1043 1111 1044 1112
rect 1038 1110 1044 1111
rect 1079 1111 1080 1112
rect 1084 1111 1085 1115
rect 1079 1110 1085 1111
rect 1206 1114 1212 1115
rect 1206 1110 1207 1114
rect 1211 1110 1212 1114
rect 1270 1111 1271 1115
rect 1276 1111 1277 1115
rect 1270 1110 1277 1111
rect 1398 1114 1404 1115
rect 1398 1110 1399 1114
rect 1403 1110 1404 1114
rect 1462 1111 1463 1115
rect 1468 1111 1469 1115
rect 1462 1110 1469 1111
rect 654 1109 660 1110
rect 830 1109 836 1110
rect 1014 1109 1020 1110
rect 1206 1109 1212 1110
rect 1398 1109 1404 1110
rect 727 1079 736 1080
rect 1474 1079 1480 1080
rect 662 1078 668 1079
rect 662 1074 663 1078
rect 667 1074 668 1078
rect 727 1075 728 1079
rect 735 1075 736 1079
rect 727 1074 736 1075
rect 846 1078 852 1079
rect 846 1074 847 1078
rect 851 1074 852 1078
rect 1030 1078 1036 1079
rect 911 1075 917 1076
rect 911 1074 912 1075
rect 662 1073 668 1074
rect 846 1073 852 1074
rect 872 1072 912 1074
rect 802 1067 808 1068
rect 802 1063 803 1067
rect 807 1066 808 1067
rect 872 1066 874 1072
rect 911 1071 912 1072
rect 916 1071 917 1075
rect 1030 1074 1031 1078
rect 1035 1074 1036 1078
rect 1222 1078 1228 1079
rect 1030 1073 1036 1074
rect 1095 1075 1104 1076
rect 911 1070 917 1071
rect 1095 1071 1096 1075
rect 1103 1071 1104 1075
rect 1222 1074 1223 1078
rect 1227 1074 1228 1078
rect 1422 1078 1428 1079
rect 1222 1073 1228 1074
rect 1286 1075 1293 1076
rect 1095 1070 1104 1071
rect 1286 1071 1287 1075
rect 1292 1071 1293 1075
rect 1422 1074 1423 1078
rect 1427 1074 1428 1078
rect 1474 1075 1475 1079
rect 1479 1078 1480 1079
rect 1487 1079 1493 1080
rect 1487 1078 1488 1079
rect 1479 1076 1488 1078
rect 1479 1075 1480 1076
rect 1474 1074 1480 1075
rect 1487 1075 1488 1076
rect 1492 1075 1493 1079
rect 1487 1074 1493 1075
rect 1422 1073 1428 1074
rect 1286 1070 1293 1071
rect 807 1064 874 1066
rect 807 1063 808 1064
rect 802 1062 808 1063
rect 110 1061 116 1062
rect 110 1057 111 1061
rect 115 1057 116 1061
rect 110 1056 116 1057
rect 1566 1061 1572 1062
rect 1566 1057 1567 1061
rect 1571 1057 1572 1061
rect 1566 1056 1572 1057
rect 914 1051 920 1052
rect 914 1047 915 1051
rect 919 1050 920 1051
rect 1098 1051 1104 1052
rect 1098 1050 1099 1051
rect 919 1048 1099 1050
rect 919 1047 920 1048
rect 914 1046 920 1047
rect 1098 1047 1099 1048
rect 1103 1047 1104 1051
rect 1098 1046 1104 1047
rect 110 1043 116 1044
rect 110 1039 111 1043
rect 115 1039 116 1043
rect 110 1038 116 1039
rect 1566 1043 1572 1044
rect 1566 1039 1567 1043
rect 1571 1039 1572 1043
rect 1566 1038 1572 1039
rect 914 1035 920 1036
rect 662 1032 668 1033
rect 846 1032 852 1033
rect 662 1028 663 1032
rect 667 1028 668 1032
rect 802 1031 808 1032
rect 802 1030 803 1031
rect 733 1028 803 1030
rect 662 1027 668 1028
rect 802 1027 803 1028
rect 807 1027 808 1031
rect 846 1028 847 1032
rect 851 1028 852 1032
rect 914 1031 915 1035
rect 919 1031 920 1035
rect 914 1030 920 1031
rect 1030 1032 1036 1033
rect 1222 1032 1228 1033
rect 1422 1032 1428 1033
rect 846 1027 852 1028
rect 1030 1028 1031 1032
rect 1035 1028 1036 1032
rect 1030 1027 1036 1028
rect 1062 1031 1068 1032
rect 1062 1027 1063 1031
rect 1067 1027 1068 1031
rect 1222 1028 1223 1032
rect 1227 1028 1228 1032
rect 1222 1027 1228 1028
rect 1270 1031 1276 1032
rect 1270 1027 1271 1031
rect 1275 1027 1276 1031
rect 1422 1028 1423 1032
rect 1427 1028 1428 1032
rect 1422 1027 1428 1028
rect 1490 1031 1496 1032
rect 1490 1027 1491 1031
rect 1495 1027 1496 1031
rect 802 1026 808 1027
rect 1062 1026 1068 1027
rect 1270 1026 1276 1027
rect 1490 1026 1496 1027
rect 550 1004 556 1005
rect 758 1004 764 1005
rect 550 1000 551 1004
rect 555 1000 556 1004
rect 550 999 556 1000
rect 582 1003 588 1004
rect 582 999 583 1003
rect 587 999 588 1003
rect 758 1000 759 1004
rect 763 1000 764 1004
rect 758 999 764 1000
rect 974 1004 980 1005
rect 1198 1004 1204 1005
rect 1430 1004 1436 1005
rect 974 1000 975 1004
rect 979 1000 980 1004
rect 974 999 980 1000
rect 1006 1003 1012 1004
rect 1006 999 1007 1003
rect 1011 999 1012 1003
rect 1198 1000 1199 1004
rect 1203 1000 1204 1004
rect 1286 1003 1292 1004
rect 1286 1002 1287 1003
rect 1269 1000 1287 1002
rect 1198 999 1204 1000
rect 1286 999 1287 1000
rect 1291 999 1292 1003
rect 1430 1000 1431 1004
rect 1435 1000 1436 1004
rect 1430 999 1436 1000
rect 1498 1003 1504 1004
rect 1498 999 1499 1003
rect 1503 999 1504 1003
rect 582 998 588 999
rect 1006 998 1012 999
rect 1286 998 1292 999
rect 1498 998 1504 999
rect 110 993 116 994
rect 110 989 111 993
rect 115 989 116 993
rect 110 988 116 989
rect 1566 993 1572 994
rect 1566 989 1567 993
rect 1571 989 1572 993
rect 1566 988 1572 989
rect 618 987 624 988
rect 618 983 619 987
rect 623 986 624 987
rect 799 987 805 988
rect 799 986 800 987
rect 623 984 800 986
rect 623 983 624 984
rect 618 982 624 983
rect 799 983 800 984
rect 804 983 805 987
rect 799 982 805 983
rect 110 975 116 976
rect 110 971 111 975
rect 115 971 116 975
rect 110 970 116 971
rect 1566 975 1572 976
rect 1566 971 1567 975
rect 1571 971 1572 975
rect 1566 970 1572 971
rect 615 959 624 960
rect 823 959 829 960
rect 1039 959 1045 960
rect 550 958 556 959
rect 550 954 551 958
rect 555 954 556 958
rect 615 955 616 959
rect 623 955 624 959
rect 615 954 624 955
rect 758 958 764 959
rect 758 954 759 958
rect 763 954 764 958
rect 823 955 824 959
rect 828 958 829 959
rect 974 958 980 959
rect 828 956 874 958
rect 828 955 829 956
rect 823 954 829 955
rect 550 953 556 954
rect 758 953 764 954
rect 872 950 874 956
rect 974 954 975 958
rect 979 954 980 958
rect 1039 955 1040 959
rect 1044 958 1045 959
rect 1062 959 1068 960
rect 1263 959 1272 960
rect 1490 959 1501 960
rect 1062 958 1063 959
rect 1044 956 1063 958
rect 1044 955 1045 956
rect 1039 954 1045 955
rect 1062 955 1063 956
rect 1067 955 1068 959
rect 1062 954 1068 955
rect 1198 958 1204 959
rect 1198 954 1199 958
rect 1203 954 1204 958
rect 1263 955 1264 959
rect 1271 955 1272 959
rect 1263 954 1272 955
rect 1430 958 1436 959
rect 1430 954 1431 958
rect 1435 954 1436 958
rect 1490 955 1491 959
rect 1495 955 1496 959
rect 1500 955 1501 959
rect 1490 954 1501 955
rect 974 953 980 954
rect 1198 953 1204 954
rect 1430 953 1436 954
rect 1006 951 1012 952
rect 1006 950 1007 951
rect 872 948 1007 950
rect 1006 947 1007 948
rect 1011 947 1012 951
rect 1006 946 1012 947
rect 614 931 620 932
rect 614 927 615 931
rect 619 930 620 931
rect 854 931 860 932
rect 619 928 690 930
rect 619 927 620 928
rect 614 926 620 927
rect 463 923 469 924
rect 398 922 404 923
rect 398 918 399 922
rect 403 918 404 922
rect 463 919 464 923
rect 468 922 469 923
rect 582 923 588 924
rect 582 922 583 923
rect 468 920 583 922
rect 468 919 469 920
rect 463 918 469 919
rect 582 919 583 920
rect 587 919 588 923
rect 582 918 588 919
rect 662 922 668 923
rect 662 918 663 922
rect 667 918 668 922
rect 688 922 690 928
rect 854 927 855 931
rect 859 930 860 931
rect 859 928 958 930
rect 859 927 860 928
rect 854 926 860 927
rect 727 923 733 924
rect 727 922 728 923
rect 688 920 728 922
rect 727 919 728 920
rect 732 919 733 923
rect 727 918 733 919
rect 926 922 932 923
rect 926 918 927 922
rect 931 918 932 922
rect 956 922 958 928
rect 991 923 997 924
rect 1498 923 1504 924
rect 991 922 992 923
rect 956 920 992 922
rect 991 919 992 920
rect 996 919 997 923
rect 991 918 997 919
rect 1198 922 1204 923
rect 1198 918 1199 922
rect 1203 918 1204 922
rect 1470 922 1476 923
rect 398 917 404 918
rect 662 917 668 918
rect 926 917 932 918
rect 1198 917 1204 918
rect 1263 919 1269 920
rect 1263 915 1264 919
rect 1268 918 1269 919
rect 1334 919 1340 920
rect 1334 918 1335 919
rect 1268 916 1335 918
rect 1268 915 1269 916
rect 1263 914 1269 915
rect 1334 915 1335 916
rect 1339 915 1340 919
rect 1470 918 1471 922
rect 1475 918 1476 922
rect 1498 919 1499 923
rect 1503 922 1504 923
rect 1535 923 1541 924
rect 1535 922 1536 923
rect 1503 920 1536 922
rect 1503 919 1504 920
rect 1498 918 1504 919
rect 1535 919 1536 920
rect 1540 919 1541 923
rect 1535 918 1541 919
rect 1470 917 1476 918
rect 1334 914 1340 915
rect 110 905 116 906
rect 110 901 111 905
rect 115 901 116 905
rect 110 900 116 901
rect 1566 905 1572 906
rect 1566 901 1567 905
rect 1571 901 1572 905
rect 1566 900 1572 901
rect 110 887 116 888
rect 110 883 111 887
rect 115 883 116 887
rect 110 882 116 883
rect 1566 887 1572 888
rect 1566 883 1567 887
rect 1571 883 1572 887
rect 1566 882 1572 883
rect 398 876 404 877
rect 662 876 668 877
rect 926 876 932 877
rect 1198 876 1204 877
rect 1470 876 1476 877
rect 398 872 399 876
rect 403 872 404 876
rect 614 875 620 876
rect 614 874 615 875
rect 469 872 615 874
rect 398 871 404 872
rect 614 871 615 872
rect 619 871 620 875
rect 662 872 663 876
rect 667 872 668 876
rect 854 875 860 876
rect 854 874 855 875
rect 733 872 855 874
rect 662 871 668 872
rect 854 871 855 872
rect 859 871 860 875
rect 926 872 927 876
rect 931 872 932 876
rect 926 871 932 872
rect 958 875 964 876
rect 958 871 959 875
rect 963 871 964 875
rect 1198 872 1199 876
rect 1203 872 1204 876
rect 1430 875 1436 876
rect 1430 874 1431 875
rect 1269 872 1431 874
rect 1198 871 1204 872
rect 1430 871 1431 872
rect 1435 871 1436 875
rect 1470 872 1471 876
rect 1475 872 1476 876
rect 1470 871 1476 872
rect 614 870 620 871
rect 854 870 860 871
rect 958 870 964 871
rect 1430 870 1436 871
rect 1334 867 1340 868
rect 1334 863 1335 867
rect 1339 866 1340 867
rect 1504 866 1506 873
rect 1339 864 1506 866
rect 1339 863 1340 864
rect 1334 862 1340 863
rect 254 852 260 853
rect 534 852 540 853
rect 254 848 255 852
rect 259 848 260 852
rect 254 847 260 848
rect 286 851 292 852
rect 286 847 287 851
rect 291 847 292 851
rect 534 848 535 852
rect 539 848 540 852
rect 534 847 540 848
rect 822 852 828 853
rect 822 848 823 852
rect 827 848 828 852
rect 822 847 828 848
rect 1110 852 1116 853
rect 1406 852 1412 853
rect 1110 848 1111 852
rect 1115 848 1116 852
rect 1266 851 1272 852
rect 1266 850 1267 851
rect 1181 848 1267 850
rect 1110 847 1116 848
rect 1266 847 1267 848
rect 1271 847 1272 851
rect 1406 848 1407 852
rect 1411 848 1412 852
rect 1406 847 1412 848
rect 1462 851 1468 852
rect 1462 847 1463 851
rect 1467 847 1468 851
rect 286 846 292 847
rect 1266 846 1272 847
rect 1462 846 1468 847
rect 110 841 116 842
rect 110 837 111 841
rect 115 837 116 841
rect 110 836 116 837
rect 1566 841 1572 842
rect 1566 837 1567 841
rect 1571 837 1572 841
rect 1566 836 1572 837
rect 322 835 328 836
rect 322 831 323 835
rect 327 834 328 835
rect 575 835 581 836
rect 575 834 576 835
rect 327 832 576 834
rect 327 831 328 832
rect 322 830 328 831
rect 575 831 576 832
rect 580 831 581 835
rect 575 830 581 831
rect 602 835 608 836
rect 602 831 603 835
rect 607 834 608 835
rect 863 835 869 836
rect 863 834 864 835
rect 607 832 864 834
rect 607 831 608 832
rect 602 830 608 831
rect 863 831 864 832
rect 868 831 869 835
rect 863 830 869 831
rect 110 823 116 824
rect 110 819 111 823
rect 115 819 116 823
rect 110 818 116 819
rect 1566 823 1572 824
rect 1566 819 1567 823
rect 1571 819 1572 823
rect 1566 818 1572 819
rect 319 807 328 808
rect 599 807 608 808
rect 887 807 893 808
rect 254 806 260 807
rect 254 802 255 806
rect 259 802 260 806
rect 319 803 320 807
rect 327 803 328 807
rect 319 802 328 803
rect 534 806 540 807
rect 534 802 535 806
rect 539 802 540 806
rect 599 803 600 807
rect 607 803 608 807
rect 599 802 608 803
rect 822 806 828 807
rect 822 802 823 806
rect 827 802 828 806
rect 887 803 888 807
rect 892 806 893 807
rect 958 807 964 808
rect 1154 807 1160 808
rect 958 806 959 807
rect 892 804 959 806
rect 892 803 893 804
rect 887 802 893 803
rect 958 803 959 804
rect 963 803 964 807
rect 958 802 964 803
rect 1110 806 1116 807
rect 1110 802 1111 806
rect 1115 802 1116 806
rect 1154 803 1155 807
rect 1159 806 1160 807
rect 1175 807 1181 808
rect 1430 807 1436 808
rect 1175 806 1176 807
rect 1159 804 1176 806
rect 1159 803 1160 804
rect 1154 802 1160 803
rect 1175 803 1176 804
rect 1180 803 1181 807
rect 1175 802 1181 803
rect 1406 806 1412 807
rect 1406 802 1407 806
rect 1411 802 1412 806
rect 1430 803 1431 807
rect 1435 806 1436 807
rect 1471 807 1477 808
rect 1471 806 1472 807
rect 1435 804 1472 806
rect 1435 803 1436 804
rect 1430 802 1436 803
rect 1471 803 1472 804
rect 1476 803 1477 807
rect 1471 802 1477 803
rect 254 801 260 802
rect 534 801 540 802
rect 822 801 828 802
rect 1110 801 1116 802
rect 1406 801 1412 802
rect 263 771 269 772
rect 198 770 204 771
rect 198 766 199 770
rect 203 766 204 770
rect 263 767 264 771
rect 268 770 269 771
rect 286 771 292 772
rect 1462 771 1469 772
rect 286 770 287 771
rect 268 768 287 770
rect 268 767 269 768
rect 263 766 269 767
rect 286 767 287 768
rect 291 767 292 771
rect 286 766 292 767
rect 486 770 492 771
rect 486 766 487 770
rect 491 766 492 770
rect 782 770 788 771
rect 198 765 204 766
rect 486 765 492 766
rect 551 767 557 768
rect 551 763 552 767
rect 556 766 557 767
rect 782 766 783 770
rect 787 766 788 770
rect 1086 770 1092 771
rect 556 764 686 766
rect 782 765 788 766
rect 847 767 856 768
rect 556 763 557 764
rect 551 762 557 763
rect 684 758 686 764
rect 847 763 848 767
rect 855 763 856 767
rect 1086 766 1087 770
rect 1091 766 1092 770
rect 1398 770 1404 771
rect 1086 765 1092 766
rect 1151 767 1157 768
rect 847 762 856 763
rect 1151 763 1152 767
rect 1156 766 1157 767
rect 1222 767 1228 768
rect 1222 766 1223 767
rect 1156 764 1223 766
rect 1156 763 1157 764
rect 1151 762 1157 763
rect 1222 763 1223 764
rect 1227 763 1228 767
rect 1398 766 1399 770
rect 1403 766 1404 770
rect 1462 767 1463 771
rect 1468 767 1469 771
rect 1462 766 1469 767
rect 1398 765 1404 766
rect 1222 762 1228 763
rect 798 759 804 760
rect 798 758 799 759
rect 684 756 799 758
rect 798 755 799 756
rect 803 755 804 759
rect 798 754 804 755
rect 110 753 116 754
rect 110 749 111 753
rect 115 749 116 753
rect 110 748 116 749
rect 1566 753 1572 754
rect 1566 749 1567 753
rect 1571 749 1572 753
rect 1566 748 1572 749
rect 850 739 856 740
rect 850 738 851 739
rect 264 736 851 738
rect 110 735 116 736
rect 110 731 111 735
rect 115 731 116 735
rect 110 730 116 731
rect 264 725 266 736
rect 850 735 851 736
rect 855 735 856 739
rect 850 734 856 735
rect 1566 735 1572 736
rect 1566 731 1567 735
rect 1571 731 1572 735
rect 1566 730 1572 731
rect 1154 727 1160 728
rect 198 724 204 725
rect 198 720 199 724
rect 203 720 204 724
rect 198 719 204 720
rect 486 724 492 725
rect 782 724 788 725
rect 1086 724 1092 725
rect 486 720 487 724
rect 491 720 492 724
rect 486 719 492 720
rect 518 723 524 724
rect 518 719 519 723
rect 523 719 524 723
rect 782 720 783 724
rect 787 720 788 724
rect 782 719 788 720
rect 798 723 804 724
rect 798 719 799 723
rect 803 722 804 723
rect 803 720 817 722
rect 1086 720 1087 724
rect 1091 720 1092 724
rect 1154 723 1155 727
rect 1159 723 1160 727
rect 1154 722 1160 723
rect 1398 724 1404 725
rect 803 719 804 720
rect 1086 719 1092 720
rect 1398 720 1399 724
rect 1403 720 1404 724
rect 1398 719 1404 720
rect 1466 723 1472 724
rect 1466 719 1467 723
rect 1471 719 1472 723
rect 518 718 524 719
rect 798 718 804 719
rect 1466 718 1472 719
rect 254 704 260 705
rect 526 704 532 705
rect 814 704 820 705
rect 1110 704 1116 705
rect 1406 704 1412 705
rect 254 700 255 704
rect 259 700 260 704
rect 438 703 444 704
rect 438 702 439 703
rect 325 700 439 702
rect 254 699 260 700
rect 438 699 439 700
rect 443 699 444 703
rect 526 700 527 704
rect 531 700 532 704
rect 798 703 804 704
rect 798 702 799 703
rect 597 700 799 702
rect 526 699 532 700
rect 798 699 799 700
rect 803 699 804 703
rect 814 700 815 704
rect 819 700 820 704
rect 1098 703 1104 704
rect 1098 702 1099 703
rect 885 700 1099 702
rect 814 699 820 700
rect 1098 699 1099 700
rect 1103 699 1104 703
rect 1110 700 1111 704
rect 1115 700 1116 704
rect 1110 699 1116 700
rect 1142 703 1148 704
rect 1142 699 1143 703
rect 1147 699 1148 703
rect 1406 700 1407 704
rect 1411 700 1412 704
rect 1406 699 1412 700
rect 1474 703 1480 704
rect 1474 699 1475 703
rect 1479 699 1480 703
rect 438 698 444 699
rect 798 698 804 699
rect 1098 698 1104 699
rect 1142 698 1148 699
rect 1474 698 1480 699
rect 110 693 116 694
rect 110 689 111 693
rect 115 689 116 693
rect 110 688 116 689
rect 1566 693 1572 694
rect 1566 689 1567 693
rect 1571 689 1572 693
rect 1566 688 1572 689
rect 110 675 116 676
rect 110 671 111 675
rect 115 671 116 675
rect 110 670 116 671
rect 1566 675 1572 676
rect 1566 671 1567 675
rect 1571 671 1572 675
rect 1566 670 1572 671
rect 438 667 444 668
rect 438 663 439 667
rect 443 666 444 667
rect 798 667 804 668
rect 443 664 554 666
rect 443 663 444 664
rect 438 662 444 663
rect 319 659 325 660
rect 254 658 260 659
rect 254 654 255 658
rect 259 654 260 658
rect 319 655 320 659
rect 324 658 325 659
rect 518 659 524 660
rect 518 658 519 659
rect 324 656 519 658
rect 324 655 325 656
rect 319 654 325 655
rect 518 655 519 656
rect 523 655 524 659
rect 518 654 524 655
rect 526 658 532 659
rect 526 654 527 658
rect 531 654 532 658
rect 552 658 554 664
rect 798 663 799 667
rect 803 666 804 667
rect 1098 667 1104 668
rect 803 664 842 666
rect 803 663 804 664
rect 798 662 804 663
rect 591 659 597 660
rect 591 658 592 659
rect 552 656 592 658
rect 591 655 592 656
rect 596 655 597 659
rect 591 654 597 655
rect 814 658 820 659
rect 814 654 815 658
rect 819 654 820 658
rect 840 658 842 664
rect 1098 663 1099 667
rect 1103 666 1104 667
rect 1103 664 1138 666
rect 1103 663 1104 664
rect 1098 662 1104 663
rect 879 659 885 660
rect 879 658 880 659
rect 840 656 880 658
rect 879 655 880 656
rect 884 655 885 659
rect 879 654 885 655
rect 1110 658 1116 659
rect 1110 654 1111 658
rect 1115 654 1116 658
rect 1136 658 1138 664
rect 1175 659 1181 660
rect 1466 659 1477 660
rect 1175 658 1176 659
rect 1136 656 1176 658
rect 1175 655 1176 656
rect 1180 655 1181 659
rect 1175 654 1181 655
rect 1406 658 1412 659
rect 1406 654 1407 658
rect 1411 654 1412 658
rect 1466 655 1467 659
rect 1471 655 1472 659
rect 1476 655 1477 659
rect 1466 654 1477 655
rect 254 653 260 654
rect 526 653 532 654
rect 814 653 820 654
rect 1110 653 1116 654
rect 1406 653 1412 654
rect 1006 639 1012 640
rect 1006 638 1007 639
rect 872 636 1007 638
rect 823 631 829 632
rect 550 630 556 631
rect 550 626 551 630
rect 555 626 556 630
rect 758 630 764 631
rect 550 625 556 626
rect 615 627 621 628
rect 615 623 616 627
rect 620 626 621 627
rect 758 626 759 630
rect 763 626 764 630
rect 823 627 824 631
rect 828 630 829 631
rect 872 630 874 636
rect 1006 635 1007 636
rect 1011 635 1012 639
rect 1006 634 1012 635
rect 1039 631 1045 632
rect 828 628 874 630
rect 974 630 980 631
rect 828 627 829 628
rect 823 626 829 627
rect 974 626 975 630
rect 979 626 980 630
rect 1039 627 1040 631
rect 1044 630 1045 631
rect 1142 631 1148 632
rect 1474 631 1485 632
rect 1142 630 1143 631
rect 1044 628 1143 630
rect 1044 627 1045 628
rect 1039 626 1045 627
rect 1142 627 1143 628
rect 1147 627 1148 631
rect 1142 626 1148 627
rect 1190 630 1196 631
rect 1190 626 1191 630
rect 1195 626 1196 630
rect 1414 630 1420 631
rect 620 624 706 626
rect 758 625 764 626
rect 974 625 980 626
rect 1190 625 1196 626
rect 1255 627 1261 628
rect 620 623 621 624
rect 615 622 621 623
rect 704 618 706 624
rect 1255 623 1256 627
rect 1260 626 1261 627
rect 1286 627 1292 628
rect 1286 626 1287 627
rect 1260 624 1287 626
rect 1260 623 1261 624
rect 1255 622 1261 623
rect 1286 623 1287 624
rect 1291 623 1292 627
rect 1414 626 1415 630
rect 1419 626 1420 630
rect 1474 627 1475 631
rect 1479 627 1480 631
rect 1484 627 1485 631
rect 1474 626 1485 627
rect 1414 625 1420 626
rect 1286 622 1292 623
rect 774 619 780 620
rect 774 618 775 619
rect 704 616 775 618
rect 774 615 775 616
rect 779 615 780 619
rect 774 614 780 615
rect 110 613 116 614
rect 110 609 111 613
rect 115 609 116 613
rect 110 608 116 609
rect 1566 613 1572 614
rect 1566 609 1567 613
rect 1571 609 1572 613
rect 1566 608 1572 609
rect 110 595 116 596
rect 110 591 111 595
rect 115 591 116 595
rect 110 590 116 591
rect 1566 595 1572 596
rect 1566 591 1567 595
rect 1571 591 1572 595
rect 1566 590 1572 591
rect 550 584 556 585
rect 758 584 764 585
rect 974 584 980 585
rect 1190 584 1196 585
rect 1414 584 1420 585
rect 550 580 551 584
rect 555 580 556 584
rect 750 583 756 584
rect 750 582 751 583
rect 621 580 751 582
rect 550 579 556 580
rect 750 579 751 580
rect 755 579 756 583
rect 758 580 759 584
rect 763 580 764 584
rect 758 579 764 580
rect 774 583 780 584
rect 774 579 775 583
rect 779 582 780 583
rect 779 580 793 582
rect 974 580 975 584
rect 979 580 980 584
rect 779 579 780 580
rect 974 579 980 580
rect 1006 583 1012 584
rect 1006 579 1007 583
rect 1011 579 1012 583
rect 1190 580 1191 584
rect 1195 580 1196 584
rect 1190 579 1196 580
rect 1222 583 1228 584
rect 1222 579 1223 583
rect 1227 579 1228 583
rect 1414 580 1415 584
rect 1419 580 1420 584
rect 1414 579 1420 580
rect 1470 583 1476 584
rect 1470 579 1471 583
rect 1475 579 1476 583
rect 750 578 756 579
rect 774 578 780 579
rect 1006 578 1012 579
rect 1222 578 1228 579
rect 1470 578 1476 579
rect 726 564 732 565
rect 846 564 852 565
rect 974 564 980 565
rect 1110 564 1116 565
rect 726 560 727 564
rect 731 560 732 564
rect 834 563 840 564
rect 834 562 835 563
rect 797 560 835 562
rect 726 559 732 560
rect 834 559 835 560
rect 839 559 840 563
rect 846 560 847 564
rect 851 560 852 564
rect 846 559 852 560
rect 914 563 920 564
rect 914 559 915 563
rect 919 559 920 563
rect 974 560 975 564
rect 979 560 980 564
rect 1090 563 1096 564
rect 1090 562 1091 563
rect 1045 560 1091 562
rect 974 559 980 560
rect 1090 559 1091 560
rect 1095 559 1096 563
rect 1110 560 1111 564
rect 1115 560 1116 564
rect 1110 559 1116 560
rect 1254 564 1260 565
rect 1406 564 1412 565
rect 1254 560 1255 564
rect 1259 560 1260 564
rect 1254 559 1260 560
rect 1286 563 1292 564
rect 1286 559 1287 563
rect 1291 559 1292 563
rect 1406 560 1407 564
rect 1411 560 1412 564
rect 1494 563 1500 564
rect 1494 562 1495 563
rect 1477 560 1495 562
rect 1406 559 1412 560
rect 1494 559 1495 560
rect 1499 559 1500 563
rect 834 558 840 559
rect 914 558 920 559
rect 1090 558 1096 559
rect 1286 558 1292 559
rect 1494 558 1500 559
rect 110 553 116 554
rect 110 549 111 553
rect 115 549 116 553
rect 110 548 116 549
rect 1566 553 1572 554
rect 1566 549 1567 553
rect 1571 549 1572 553
rect 1566 548 1572 549
rect 1103 547 1109 548
rect 1103 543 1104 547
rect 1108 546 1109 547
rect 1151 547 1157 548
rect 1151 546 1152 547
rect 1108 544 1152 546
rect 1108 543 1109 544
rect 1103 542 1109 543
rect 1151 543 1152 544
rect 1156 543 1157 547
rect 1151 542 1157 543
rect 110 535 116 536
rect 110 531 111 535
rect 115 531 116 535
rect 110 530 116 531
rect 1566 535 1572 536
rect 1566 531 1567 535
rect 1571 531 1572 535
rect 1566 530 1572 531
rect 834 527 840 528
rect 834 523 835 527
rect 839 526 840 527
rect 1090 527 1096 528
rect 839 524 874 526
rect 839 523 840 524
rect 834 522 840 523
rect 750 519 756 520
rect 726 518 732 519
rect 726 514 727 518
rect 731 514 732 518
rect 750 515 751 519
rect 755 518 756 519
rect 791 519 797 520
rect 791 518 792 519
rect 755 516 792 518
rect 755 515 756 516
rect 750 514 756 515
rect 791 515 792 516
rect 796 515 797 519
rect 791 514 797 515
rect 846 518 852 519
rect 846 514 847 518
rect 851 514 852 518
rect 872 518 874 524
rect 1090 523 1091 527
rect 1095 526 1096 527
rect 1095 524 1138 526
rect 1095 523 1096 524
rect 1090 522 1096 523
rect 911 519 917 520
rect 1039 519 1045 520
rect 911 518 912 519
rect 872 516 912 518
rect 911 515 912 516
rect 916 515 917 519
rect 911 514 917 515
rect 974 518 980 519
rect 1039 518 1040 519
rect 974 514 975 518
rect 979 514 980 518
rect 726 513 732 514
rect 846 513 852 514
rect 974 513 980 514
rect 1000 516 1040 518
rect 914 511 920 512
rect 914 507 915 511
rect 919 510 920 511
rect 1000 510 1002 516
rect 1039 515 1040 516
rect 1044 515 1045 519
rect 1039 514 1045 515
rect 1110 518 1116 519
rect 1110 514 1111 518
rect 1115 514 1116 518
rect 1136 518 1138 524
rect 1175 519 1181 520
rect 1319 519 1325 520
rect 1470 519 1477 520
rect 1175 518 1176 519
rect 1136 516 1176 518
rect 1175 515 1176 516
rect 1180 515 1181 519
rect 1175 514 1181 515
rect 1254 518 1260 519
rect 1319 518 1320 519
rect 1254 514 1255 518
rect 1259 514 1260 518
rect 1110 513 1116 514
rect 1254 513 1260 514
rect 1280 516 1320 518
rect 919 508 1002 510
rect 1186 511 1192 512
rect 919 507 920 508
rect 914 506 920 507
rect 1186 507 1187 511
rect 1191 510 1192 511
rect 1280 510 1282 516
rect 1319 515 1320 516
rect 1324 515 1325 519
rect 1319 514 1325 515
rect 1406 518 1412 519
rect 1406 514 1407 518
rect 1411 514 1412 518
rect 1470 515 1471 519
rect 1476 515 1477 519
rect 1470 514 1477 515
rect 1406 513 1412 514
rect 1191 508 1282 510
rect 1191 507 1192 508
rect 1186 506 1192 507
rect 1095 483 1101 484
rect 766 482 772 483
rect 766 478 767 482
rect 771 478 772 482
rect 854 482 860 483
rect 766 477 772 478
rect 831 479 837 480
rect 831 475 832 479
rect 836 478 837 479
rect 854 478 855 482
rect 859 478 860 482
rect 942 482 948 483
rect 836 476 850 478
rect 854 477 860 478
rect 919 479 925 480
rect 836 475 837 476
rect 831 474 837 475
rect 848 470 850 476
rect 919 475 920 479
rect 924 478 925 479
rect 942 478 943 482
rect 947 478 948 482
rect 1030 482 1036 483
rect 924 476 938 478
rect 942 477 948 478
rect 1007 479 1013 480
rect 924 475 925 476
rect 919 474 925 475
rect 870 471 876 472
rect 870 470 871 471
rect 848 468 871 470
rect 870 467 871 468
rect 875 467 876 471
rect 936 470 938 476
rect 1007 475 1008 479
rect 1012 478 1013 479
rect 1030 478 1031 482
rect 1035 478 1036 482
rect 1095 479 1096 483
rect 1100 482 1101 483
rect 1103 483 1109 484
rect 1494 483 1500 484
rect 1103 482 1104 483
rect 1100 480 1104 482
rect 1100 479 1101 480
rect 1095 478 1101 479
rect 1103 479 1104 480
rect 1108 479 1109 483
rect 1103 478 1109 479
rect 1118 482 1124 483
rect 1118 478 1119 482
rect 1123 478 1124 482
rect 1206 482 1212 483
rect 1012 476 1026 478
rect 1030 477 1036 478
rect 1118 477 1124 478
rect 1183 479 1189 480
rect 1012 475 1013 476
rect 1007 474 1013 475
rect 958 471 964 472
rect 958 470 959 471
rect 936 468 959 470
rect 870 466 876 467
rect 958 467 959 468
rect 963 467 964 471
rect 1024 470 1026 476
rect 1183 475 1184 479
rect 1188 478 1189 479
rect 1206 478 1207 482
rect 1211 478 1212 482
rect 1294 482 1300 483
rect 1188 476 1202 478
rect 1206 477 1212 478
rect 1271 479 1277 480
rect 1188 475 1189 476
rect 1183 474 1189 475
rect 1046 471 1052 472
rect 1046 470 1047 471
rect 1024 468 1047 470
rect 958 466 964 467
rect 1046 467 1047 468
rect 1051 467 1052 471
rect 1200 470 1202 476
rect 1271 475 1272 479
rect 1276 478 1277 479
rect 1294 478 1295 482
rect 1299 478 1300 482
rect 1382 482 1388 483
rect 1276 476 1290 478
rect 1294 477 1300 478
rect 1359 479 1365 480
rect 1276 475 1277 476
rect 1271 474 1277 475
rect 1222 471 1228 472
rect 1222 470 1223 471
rect 1200 468 1223 470
rect 1046 466 1052 467
rect 1222 467 1223 468
rect 1227 467 1228 471
rect 1288 470 1290 476
rect 1359 475 1360 479
rect 1364 478 1365 479
rect 1382 478 1383 482
rect 1387 478 1388 482
rect 1470 482 1476 483
rect 1364 476 1378 478
rect 1382 477 1388 478
rect 1447 479 1453 480
rect 1364 475 1365 476
rect 1359 474 1365 475
rect 1310 471 1316 472
rect 1310 470 1311 471
rect 1288 468 1311 470
rect 1222 466 1228 467
rect 1310 467 1311 468
rect 1315 467 1316 471
rect 1376 470 1378 476
rect 1447 475 1448 479
rect 1452 478 1453 479
rect 1470 478 1471 482
rect 1475 478 1476 482
rect 1494 479 1495 483
rect 1499 482 1500 483
rect 1535 483 1541 484
rect 1535 482 1536 483
rect 1499 480 1536 482
rect 1499 479 1500 480
rect 1494 478 1500 479
rect 1535 479 1536 480
rect 1540 479 1541 483
rect 1535 478 1541 479
rect 1452 476 1466 478
rect 1470 477 1476 478
rect 1452 475 1453 476
rect 1447 474 1453 475
rect 1398 471 1404 472
rect 1398 470 1399 471
rect 1376 468 1399 470
rect 1310 466 1316 467
rect 1398 467 1399 468
rect 1403 467 1404 471
rect 1464 470 1466 476
rect 1486 471 1492 472
rect 1486 470 1487 471
rect 1464 468 1487 470
rect 1398 466 1404 467
rect 1486 467 1487 468
rect 1491 467 1492 471
rect 1486 466 1492 467
rect 110 465 116 466
rect 110 461 111 465
rect 115 461 116 465
rect 110 460 116 461
rect 1566 465 1572 466
rect 1566 461 1567 465
rect 1571 461 1572 465
rect 1566 460 1572 461
rect 934 451 940 452
rect 934 450 935 451
rect 832 448 935 450
rect 110 447 116 448
rect 110 443 111 447
rect 115 443 116 447
rect 110 442 116 443
rect 832 437 834 448
rect 934 447 935 448
rect 939 447 940 451
rect 934 446 940 447
rect 1566 447 1572 448
rect 1566 443 1567 447
rect 1571 443 1572 447
rect 1566 442 1572 443
rect 1186 439 1192 440
rect 766 436 772 437
rect 766 432 767 436
rect 771 432 772 436
rect 766 431 772 432
rect 854 436 860 437
rect 942 436 948 437
rect 1030 436 1036 437
rect 1118 436 1124 437
rect 854 432 855 436
rect 859 432 860 436
rect 854 431 860 432
rect 870 435 876 436
rect 870 431 871 435
rect 875 434 876 435
rect 875 432 889 434
rect 942 432 943 436
rect 947 432 948 436
rect 875 431 876 432
rect 942 431 948 432
rect 958 435 964 436
rect 958 431 959 435
rect 963 434 964 435
rect 963 432 977 434
rect 1030 432 1031 436
rect 1035 432 1036 436
rect 963 431 964 432
rect 1030 431 1036 432
rect 1046 435 1052 436
rect 1046 431 1047 435
rect 1051 434 1052 435
rect 1051 432 1065 434
rect 1118 432 1119 436
rect 1123 432 1124 436
rect 1186 435 1187 439
rect 1191 435 1192 439
rect 1186 434 1192 435
rect 1206 436 1212 437
rect 1294 436 1300 437
rect 1382 436 1388 437
rect 1470 436 1476 437
rect 1051 431 1052 432
rect 1118 431 1124 432
rect 1206 432 1207 436
rect 1211 432 1212 436
rect 1206 431 1212 432
rect 1222 435 1228 436
rect 1222 431 1223 435
rect 1227 434 1228 435
rect 1227 432 1241 434
rect 1294 432 1295 436
rect 1299 432 1300 436
rect 1227 431 1228 432
rect 1294 431 1300 432
rect 1310 435 1316 436
rect 1310 431 1311 435
rect 1315 434 1316 435
rect 1315 432 1329 434
rect 1382 432 1383 436
rect 1387 432 1388 436
rect 1315 431 1316 432
rect 1382 431 1388 432
rect 1398 435 1404 436
rect 1398 431 1399 435
rect 1403 434 1404 435
rect 1403 432 1417 434
rect 1470 432 1471 436
rect 1475 432 1476 436
rect 1403 431 1404 432
rect 1470 431 1476 432
rect 1486 435 1492 436
rect 1486 431 1487 435
rect 1491 434 1492 435
rect 1491 432 1505 434
rect 1491 431 1492 432
rect 870 430 876 431
rect 958 430 964 431
rect 1046 430 1052 431
rect 1222 430 1228 431
rect 1310 430 1316 431
rect 1398 430 1404 431
rect 1486 430 1492 431
rect 622 408 628 409
rect 710 408 716 409
rect 622 404 623 408
rect 627 404 628 408
rect 698 407 704 408
rect 698 406 699 407
rect 693 404 699 406
rect 622 403 628 404
rect 698 403 699 404
rect 703 403 704 407
rect 710 404 711 408
rect 715 404 716 408
rect 710 403 716 404
rect 798 408 804 409
rect 798 404 799 408
rect 803 404 804 408
rect 798 403 804 404
rect 886 408 892 409
rect 886 404 887 408
rect 891 404 892 408
rect 886 403 892 404
rect 918 407 924 408
rect 918 403 919 407
rect 923 403 924 407
rect 698 402 704 403
rect 918 402 924 403
rect 110 397 116 398
rect 110 393 111 397
rect 115 393 116 397
rect 110 392 116 393
rect 1566 397 1572 398
rect 1566 393 1567 397
rect 1571 393 1572 397
rect 1566 392 1572 393
rect 690 391 696 392
rect 690 387 691 391
rect 695 390 696 391
rect 751 391 757 392
rect 751 390 752 391
rect 695 388 752 390
rect 695 387 696 388
rect 690 386 696 387
rect 751 387 752 388
rect 756 387 757 391
rect 751 386 757 387
rect 778 391 784 392
rect 778 387 779 391
rect 783 390 784 391
rect 839 391 845 392
rect 839 390 840 391
rect 783 388 840 390
rect 783 387 784 388
rect 778 386 784 387
rect 839 387 840 388
rect 844 387 845 391
rect 839 386 845 387
rect 110 379 116 380
rect 110 375 111 379
rect 115 375 116 379
rect 110 374 116 375
rect 1566 379 1572 380
rect 1566 375 1567 379
rect 1571 375 1572 379
rect 1566 374 1572 375
rect 687 363 696 364
rect 775 363 784 364
rect 863 363 869 364
rect 934 363 940 364
rect 622 362 628 363
rect 622 358 623 362
rect 627 358 628 362
rect 687 359 688 363
rect 695 359 696 363
rect 687 358 696 359
rect 710 362 716 363
rect 710 358 711 362
rect 715 358 716 362
rect 775 359 776 363
rect 783 359 784 363
rect 775 358 784 359
rect 798 362 804 363
rect 798 358 799 362
rect 803 358 804 362
rect 863 359 864 363
rect 868 362 869 363
rect 886 362 892 363
rect 868 360 882 362
rect 868 359 869 360
rect 863 358 869 359
rect 622 357 628 358
rect 710 357 716 358
rect 798 357 804 358
rect 880 354 882 360
rect 886 358 887 362
rect 891 358 892 362
rect 934 359 935 363
rect 939 362 940 363
rect 951 363 957 364
rect 951 362 952 363
rect 939 360 952 362
rect 939 359 940 360
rect 934 358 940 359
rect 951 359 952 360
rect 956 359 957 363
rect 951 358 957 359
rect 886 357 892 358
rect 918 355 924 356
rect 918 354 919 355
rect 880 352 919 354
rect 918 351 919 352
rect 923 351 924 355
rect 918 350 924 351
rect 698 323 704 324
rect 398 322 404 323
rect 398 318 399 322
rect 403 318 404 322
rect 486 322 492 323
rect 398 317 404 318
rect 463 319 469 320
rect 463 315 464 319
rect 468 318 469 319
rect 486 318 487 322
rect 491 318 492 322
rect 574 322 580 323
rect 468 316 482 318
rect 486 317 492 318
rect 551 319 557 320
rect 468 315 469 316
rect 463 314 469 315
rect 480 310 482 316
rect 551 315 552 319
rect 556 318 557 319
rect 574 318 575 322
rect 579 318 580 322
rect 662 322 668 323
rect 556 316 570 318
rect 574 317 580 318
rect 639 319 645 320
rect 556 315 557 316
rect 551 314 557 315
rect 502 311 508 312
rect 502 310 503 311
rect 480 308 503 310
rect 502 307 503 308
rect 507 307 508 311
rect 568 310 570 316
rect 639 315 640 319
rect 644 318 645 319
rect 662 318 663 322
rect 667 318 668 322
rect 698 319 699 323
rect 703 322 704 323
rect 727 323 733 324
rect 727 322 728 323
rect 703 320 728 322
rect 703 319 704 320
rect 698 318 704 319
rect 727 319 728 320
rect 732 319 733 323
rect 727 318 733 319
rect 644 316 658 318
rect 662 317 668 318
rect 644 315 645 316
rect 639 314 645 315
rect 590 311 596 312
rect 590 310 591 311
rect 568 308 591 310
rect 502 306 508 307
rect 590 307 591 308
rect 595 307 596 311
rect 656 310 658 316
rect 678 311 684 312
rect 678 310 679 311
rect 656 308 679 310
rect 590 306 596 307
rect 678 307 679 308
rect 683 307 684 311
rect 678 306 684 307
rect 110 305 116 306
rect 110 301 111 305
rect 115 301 116 305
rect 110 300 116 301
rect 1566 305 1572 306
rect 1566 301 1567 305
rect 1571 301 1572 305
rect 1566 300 1572 301
rect 110 287 116 288
rect 110 283 111 287
rect 115 283 116 287
rect 110 282 116 283
rect 1566 287 1572 288
rect 1566 283 1567 287
rect 1571 283 1572 287
rect 1566 282 1572 283
rect 398 276 404 277
rect 486 276 492 277
rect 574 276 580 277
rect 662 276 668 277
rect 398 272 399 276
rect 403 272 404 276
rect 398 271 404 272
rect 466 275 472 276
rect 466 271 467 275
rect 471 271 472 275
rect 486 272 487 276
rect 491 272 492 276
rect 486 271 492 272
rect 502 275 508 276
rect 502 271 503 275
rect 507 274 508 275
rect 507 272 521 274
rect 574 272 575 276
rect 579 272 580 276
rect 507 271 508 272
rect 574 271 580 272
rect 590 275 596 276
rect 590 271 591 275
rect 595 274 596 275
rect 595 272 609 274
rect 662 272 663 276
rect 667 272 668 276
rect 595 271 596 272
rect 662 271 668 272
rect 678 275 684 276
rect 678 271 679 275
rect 683 274 684 275
rect 683 272 697 274
rect 683 271 684 272
rect 466 270 472 271
rect 502 270 508 271
rect 590 270 596 271
rect 678 270 684 271
rect 214 244 220 245
rect 302 244 308 245
rect 214 240 215 244
rect 219 240 220 244
rect 214 239 220 240
rect 274 243 280 244
rect 274 239 275 243
rect 279 239 280 243
rect 302 240 303 244
rect 307 240 308 244
rect 302 239 308 240
rect 390 244 396 245
rect 390 240 391 244
rect 395 240 396 244
rect 390 239 396 240
rect 478 244 484 245
rect 478 240 479 244
rect 483 240 484 244
rect 478 239 484 240
rect 274 238 280 239
rect 110 233 116 234
rect 110 229 111 233
rect 115 229 116 233
rect 110 228 116 229
rect 1566 233 1572 234
rect 1566 229 1567 233
rect 1571 229 1572 233
rect 1566 228 1572 229
rect 282 227 288 228
rect 282 223 283 227
rect 287 226 288 227
rect 343 227 349 228
rect 343 226 344 227
rect 287 224 344 226
rect 287 223 288 224
rect 282 222 288 223
rect 343 223 344 224
rect 348 223 349 227
rect 343 222 349 223
rect 370 227 376 228
rect 370 223 371 227
rect 375 226 376 227
rect 431 227 437 228
rect 431 226 432 227
rect 375 224 432 226
rect 375 223 376 224
rect 370 222 376 223
rect 431 223 432 224
rect 436 223 437 227
rect 431 222 437 223
rect 458 227 464 228
rect 458 223 459 227
rect 463 226 464 227
rect 519 227 525 228
rect 519 226 520 227
rect 463 224 520 226
rect 463 223 464 224
rect 458 222 464 223
rect 519 223 520 224
rect 524 223 525 227
rect 519 222 525 223
rect 110 215 116 216
rect 110 211 111 215
rect 115 211 116 215
rect 110 210 116 211
rect 1566 215 1572 216
rect 1566 211 1567 215
rect 1571 211 1572 215
rect 1566 210 1572 211
rect 466 207 472 208
rect 466 203 467 207
rect 471 206 472 207
rect 471 204 506 206
rect 471 203 472 204
rect 466 202 472 203
rect 279 199 288 200
rect 367 199 376 200
rect 455 199 464 200
rect 214 198 220 199
rect 214 194 215 198
rect 219 194 220 198
rect 279 195 280 199
rect 287 195 288 199
rect 279 194 288 195
rect 302 198 308 199
rect 302 194 303 198
rect 307 194 308 198
rect 367 195 368 199
rect 375 195 376 199
rect 367 194 376 195
rect 390 198 396 199
rect 390 194 391 198
rect 395 194 396 198
rect 455 195 456 199
rect 463 195 464 199
rect 455 194 464 195
rect 478 198 484 199
rect 478 194 479 198
rect 483 194 484 198
rect 504 198 506 204
rect 543 199 549 200
rect 543 198 544 199
rect 504 196 544 198
rect 543 195 544 196
rect 548 195 549 199
rect 543 194 549 195
rect 214 193 220 194
rect 302 193 308 194
rect 390 193 396 194
rect 478 193 484 194
rect 598 143 604 144
rect 134 142 140 143
rect 134 138 135 142
rect 139 138 140 142
rect 222 142 228 143
rect 134 137 140 138
rect 199 139 205 140
rect 199 135 200 139
rect 204 138 205 139
rect 222 138 223 142
rect 227 138 228 142
rect 310 142 316 143
rect 204 136 218 138
rect 222 137 228 138
rect 287 139 293 140
rect 204 135 205 136
rect 199 134 205 135
rect 216 130 218 136
rect 287 135 288 139
rect 292 138 293 139
rect 310 138 311 142
rect 315 138 316 142
rect 398 142 404 143
rect 292 136 306 138
rect 310 137 316 138
rect 375 139 381 140
rect 292 135 293 136
rect 287 134 293 135
rect 238 131 244 132
rect 238 130 239 131
rect 216 128 239 130
rect 238 127 239 128
rect 243 127 244 131
rect 304 130 306 136
rect 375 135 376 139
rect 380 138 381 139
rect 398 138 399 142
rect 403 138 404 142
rect 486 142 492 143
rect 380 136 394 138
rect 398 137 404 138
rect 463 139 469 140
rect 380 135 381 136
rect 375 134 381 135
rect 326 131 332 132
rect 326 130 327 131
rect 304 128 327 130
rect 238 126 244 127
rect 326 127 327 128
rect 331 127 332 131
rect 392 130 394 136
rect 463 135 464 139
rect 468 138 469 139
rect 486 138 487 142
rect 491 138 492 142
rect 574 142 580 143
rect 468 136 482 138
rect 486 137 492 138
rect 551 139 557 140
rect 468 135 469 136
rect 463 134 469 135
rect 414 131 420 132
rect 414 130 415 131
rect 392 128 415 130
rect 326 126 332 127
rect 414 127 415 128
rect 419 127 420 131
rect 480 130 482 136
rect 551 135 552 139
rect 556 138 557 139
rect 574 138 575 142
rect 579 138 580 142
rect 598 139 599 143
rect 603 142 604 143
rect 639 143 645 144
rect 639 142 640 143
rect 603 140 640 142
rect 603 139 604 140
rect 598 138 604 139
rect 639 139 640 140
rect 644 139 645 143
rect 639 138 645 139
rect 556 136 570 138
rect 574 137 580 138
rect 556 135 557 136
rect 551 134 557 135
rect 502 131 508 132
rect 502 130 503 131
rect 480 128 503 130
rect 414 126 420 127
rect 502 127 503 128
rect 507 127 508 131
rect 568 130 570 136
rect 590 131 596 132
rect 590 130 591 131
rect 568 128 591 130
rect 502 126 508 127
rect 590 127 591 128
rect 595 127 596 131
rect 590 126 596 127
rect 110 125 116 126
rect 110 121 111 125
rect 115 121 116 125
rect 110 120 116 121
rect 1566 125 1572 126
rect 1566 121 1567 125
rect 1571 121 1572 125
rect 1566 120 1572 121
rect 110 107 116 108
rect 110 103 111 107
rect 115 103 116 107
rect 110 102 116 103
rect 1566 107 1572 108
rect 1566 103 1567 107
rect 1571 103 1572 107
rect 1566 102 1572 103
rect 134 96 140 97
rect 134 92 135 96
rect 139 92 140 96
rect 134 91 140 92
rect 222 96 228 97
rect 310 96 316 97
rect 398 96 404 97
rect 486 96 492 97
rect 574 96 580 97
rect 222 92 223 96
rect 227 92 228 96
rect 222 91 228 92
rect 238 95 244 96
rect 238 91 239 95
rect 243 94 244 95
rect 243 92 257 94
rect 310 92 311 96
rect 315 92 316 96
rect 243 91 244 92
rect 310 91 316 92
rect 326 95 332 96
rect 326 91 327 95
rect 331 94 332 95
rect 331 92 345 94
rect 398 92 399 96
rect 403 92 404 96
rect 331 91 332 92
rect 398 91 404 92
rect 414 95 420 96
rect 414 91 415 95
rect 419 94 420 95
rect 419 92 433 94
rect 486 92 487 96
rect 491 92 492 96
rect 419 91 420 92
rect 486 91 492 92
rect 502 95 508 96
rect 502 91 503 95
rect 507 94 508 95
rect 507 92 521 94
rect 574 92 575 96
rect 579 92 580 96
rect 507 91 508 92
rect 574 91 580 92
rect 590 95 596 96
rect 590 91 591 95
rect 595 94 596 95
rect 595 92 609 94
rect 595 91 596 92
rect 238 90 244 91
rect 326 90 332 91
rect 414 90 420 91
rect 502 90 508 91
rect 590 90 596 91
<< m3c >>
rect 543 1514 547 1518
rect 631 1514 635 1518
rect 719 1514 723 1518
rect 647 1503 651 1507
rect 807 1514 811 1518
rect 735 1503 739 1507
rect 887 1511 891 1515
rect 895 1514 899 1518
rect 975 1511 979 1515
rect 823 1503 827 1507
rect 111 1497 115 1501
rect 1567 1497 1571 1501
rect 111 1479 115 1483
rect 887 1483 891 1487
rect 1567 1479 1571 1483
rect 543 1468 547 1472
rect 623 1467 627 1471
rect 631 1468 635 1472
rect 647 1467 651 1471
rect 719 1468 723 1472
rect 735 1467 739 1471
rect 807 1468 811 1472
rect 823 1467 827 1471
rect 895 1468 899 1472
rect 471 1456 475 1460
rect 503 1455 507 1459
rect 615 1456 619 1460
rect 775 1456 779 1460
rect 943 1456 947 1460
rect 975 1455 979 1459
rect 1119 1456 1123 1460
rect 1303 1456 1307 1460
rect 1435 1455 1439 1459
rect 1471 1456 1475 1460
rect 1495 1455 1499 1459
rect 111 1445 115 1449
rect 1567 1445 1571 1449
rect 539 1439 543 1443
rect 683 1439 687 1443
rect 1011 1439 1015 1443
rect 111 1427 115 1431
rect 1567 1427 1571 1431
rect 1435 1419 1439 1423
rect 471 1410 475 1414
rect 539 1411 540 1415
rect 540 1411 543 1415
rect 615 1410 619 1414
rect 683 1411 684 1415
rect 684 1411 687 1415
rect 775 1410 779 1414
rect 623 1403 627 1407
rect 943 1410 947 1414
rect 1011 1411 1012 1415
rect 1012 1411 1015 1415
rect 1119 1410 1123 1414
rect 1199 1411 1203 1415
rect 1303 1410 1307 1414
rect 1471 1410 1475 1414
rect 423 1382 427 1386
rect 503 1383 507 1387
rect 663 1382 667 1386
rect 591 1371 595 1375
rect 911 1382 915 1386
rect 979 1379 980 1383
rect 980 1379 983 1383
rect 1167 1382 1171 1386
rect 1207 1379 1211 1383
rect 1431 1382 1435 1386
rect 1495 1385 1499 1387
rect 1495 1383 1496 1385
rect 1496 1383 1499 1385
rect 111 1365 115 1369
rect 1567 1365 1571 1369
rect 731 1355 735 1359
rect 979 1355 983 1359
rect 111 1347 115 1351
rect 1567 1347 1571 1351
rect 423 1336 427 1340
rect 591 1335 595 1339
rect 663 1336 667 1340
rect 731 1339 735 1343
rect 911 1336 915 1340
rect 855 1327 859 1331
rect 1167 1336 1171 1340
rect 1199 1335 1203 1339
rect 1431 1336 1435 1340
rect 1499 1335 1503 1339
rect 487 1312 491 1316
rect 563 1311 567 1315
rect 727 1312 731 1316
rect 967 1312 971 1316
rect 1207 1311 1211 1315
rect 1215 1312 1219 1316
rect 1423 1311 1427 1315
rect 1463 1312 1467 1316
rect 111 1301 115 1305
rect 1567 1301 1571 1305
rect 555 1295 559 1299
rect 1283 1295 1287 1299
rect 111 1283 115 1287
rect 1567 1283 1571 1287
rect 487 1266 491 1270
rect 555 1267 556 1271
rect 556 1267 559 1271
rect 727 1266 731 1270
rect 855 1267 859 1271
rect 967 1266 971 1270
rect 1207 1267 1211 1271
rect 1215 1266 1219 1270
rect 1283 1267 1284 1271
rect 1284 1267 1287 1271
rect 1463 1266 1467 1270
rect 1499 1267 1503 1271
rect 535 1230 539 1234
rect 563 1231 567 1235
rect 743 1230 747 1234
rect 687 1219 691 1223
rect 959 1230 963 1234
rect 983 1227 987 1231
rect 1175 1230 1179 1234
rect 1239 1227 1240 1231
rect 1240 1227 1243 1231
rect 1399 1230 1403 1234
rect 1423 1231 1427 1235
rect 111 1213 115 1217
rect 1567 1213 1571 1217
rect 111 1195 115 1199
rect 1567 1195 1571 1199
rect 535 1184 539 1188
rect 687 1183 691 1187
rect 743 1184 747 1188
rect 959 1184 963 1188
rect 1039 1183 1043 1187
rect 1175 1184 1179 1188
rect 1207 1183 1211 1187
rect 1399 1184 1403 1188
rect 1463 1183 1467 1187
rect 983 1175 987 1179
rect 655 1156 659 1160
rect 731 1155 735 1159
rect 831 1156 835 1160
rect 1015 1156 1019 1160
rect 1207 1156 1211 1160
rect 1239 1155 1243 1159
rect 1399 1156 1403 1160
rect 1475 1155 1479 1159
rect 111 1145 115 1149
rect 1567 1145 1571 1149
rect 723 1139 727 1143
rect 955 1139 959 1143
rect 111 1127 115 1131
rect 1567 1127 1571 1131
rect 655 1110 659 1114
rect 723 1111 724 1115
rect 724 1111 727 1115
rect 831 1110 835 1114
rect 955 1111 959 1115
rect 1015 1110 1019 1114
rect 1039 1111 1043 1115
rect 1207 1110 1211 1114
rect 1271 1111 1272 1115
rect 1272 1111 1275 1115
rect 1399 1110 1403 1114
rect 1463 1111 1464 1115
rect 1464 1111 1467 1115
rect 663 1074 667 1078
rect 731 1075 732 1079
rect 732 1075 735 1079
rect 847 1074 851 1078
rect 803 1063 807 1067
rect 1031 1074 1035 1078
rect 1099 1071 1100 1075
rect 1100 1071 1103 1075
rect 1223 1074 1227 1078
rect 1287 1071 1288 1075
rect 1288 1071 1291 1075
rect 1423 1074 1427 1078
rect 1475 1075 1479 1079
rect 111 1057 115 1061
rect 1567 1057 1571 1061
rect 915 1047 919 1051
rect 1099 1047 1103 1051
rect 111 1039 115 1043
rect 1567 1039 1571 1043
rect 663 1028 667 1032
rect 803 1027 807 1031
rect 847 1028 851 1032
rect 915 1031 919 1035
rect 1031 1028 1035 1032
rect 1063 1027 1067 1031
rect 1223 1028 1227 1032
rect 1271 1027 1275 1031
rect 1423 1028 1427 1032
rect 1491 1027 1495 1031
rect 551 1000 555 1004
rect 583 999 587 1003
rect 759 1000 763 1004
rect 975 1000 979 1004
rect 1007 999 1011 1003
rect 1199 1000 1203 1004
rect 1287 999 1291 1003
rect 1431 1000 1435 1004
rect 1499 999 1503 1003
rect 111 989 115 993
rect 1567 989 1571 993
rect 619 983 623 987
rect 111 971 115 975
rect 1567 971 1571 975
rect 551 954 555 958
rect 619 955 620 959
rect 620 955 623 959
rect 759 954 763 958
rect 975 954 979 958
rect 1063 955 1067 959
rect 1199 954 1203 958
rect 1267 955 1268 959
rect 1268 955 1271 959
rect 1431 954 1435 958
rect 1491 955 1495 959
rect 1007 947 1011 951
rect 615 927 619 931
rect 399 918 403 922
rect 583 919 587 923
rect 663 918 667 922
rect 855 927 859 931
rect 927 918 931 922
rect 1199 918 1203 922
rect 1335 915 1339 919
rect 1471 918 1475 922
rect 1499 919 1503 923
rect 111 901 115 905
rect 1567 901 1571 905
rect 111 883 115 887
rect 1567 883 1571 887
rect 399 872 403 876
rect 615 871 619 875
rect 663 872 667 876
rect 855 871 859 875
rect 927 872 931 876
rect 959 871 963 875
rect 1199 872 1203 876
rect 1431 871 1435 875
rect 1471 872 1475 876
rect 1335 863 1339 867
rect 255 848 259 852
rect 287 847 291 851
rect 535 848 539 852
rect 823 848 827 852
rect 1111 848 1115 852
rect 1267 847 1271 851
rect 1407 848 1411 852
rect 1463 847 1467 851
rect 111 837 115 841
rect 1567 837 1571 841
rect 323 831 327 835
rect 603 831 607 835
rect 111 819 115 823
rect 1567 819 1571 823
rect 255 802 259 806
rect 323 803 324 807
rect 324 803 327 807
rect 535 802 539 806
rect 603 803 604 807
rect 604 803 607 807
rect 823 802 827 806
rect 959 803 963 807
rect 1111 802 1115 806
rect 1155 803 1159 807
rect 1407 802 1411 806
rect 1431 803 1435 807
rect 199 766 203 770
rect 287 767 291 771
rect 487 766 491 770
rect 783 766 787 770
rect 851 763 852 767
rect 852 763 855 767
rect 1087 766 1091 770
rect 1223 763 1227 767
rect 1399 766 1403 770
rect 1463 767 1464 771
rect 1464 767 1467 771
rect 799 755 803 759
rect 111 749 115 753
rect 1567 749 1571 753
rect 111 731 115 735
rect 851 735 855 739
rect 1567 731 1571 735
rect 199 720 203 724
rect 487 720 491 724
rect 519 719 523 723
rect 783 720 787 724
rect 799 719 803 723
rect 1087 720 1091 724
rect 1155 723 1159 727
rect 1399 720 1403 724
rect 1467 719 1471 723
rect 255 700 259 704
rect 439 699 443 703
rect 527 700 531 704
rect 799 699 803 703
rect 815 700 819 704
rect 1099 699 1103 703
rect 1111 700 1115 704
rect 1143 699 1147 703
rect 1407 700 1411 704
rect 1475 699 1479 703
rect 111 689 115 693
rect 1567 689 1571 693
rect 111 671 115 675
rect 1567 671 1571 675
rect 439 663 443 667
rect 255 654 259 658
rect 519 655 523 659
rect 527 654 531 658
rect 799 663 803 667
rect 815 654 819 658
rect 1099 663 1103 667
rect 1111 654 1115 658
rect 1407 654 1411 658
rect 1467 655 1471 659
rect 551 626 555 630
rect 759 626 763 630
rect 1007 635 1011 639
rect 975 626 979 630
rect 1143 627 1147 631
rect 1191 626 1195 630
rect 1287 623 1291 627
rect 1415 626 1419 630
rect 1475 627 1479 631
rect 775 615 779 619
rect 111 609 115 613
rect 1567 609 1571 613
rect 111 591 115 595
rect 1567 591 1571 595
rect 551 580 555 584
rect 751 579 755 583
rect 759 580 763 584
rect 775 579 779 583
rect 975 580 979 584
rect 1007 579 1011 583
rect 1191 580 1195 584
rect 1223 579 1227 583
rect 1415 580 1419 584
rect 1471 579 1475 583
rect 727 560 731 564
rect 835 559 839 563
rect 847 560 851 564
rect 915 559 919 563
rect 975 560 979 564
rect 1091 559 1095 563
rect 1111 560 1115 564
rect 1255 560 1259 564
rect 1287 559 1291 563
rect 1407 560 1411 564
rect 1495 559 1499 563
rect 111 549 115 553
rect 1567 549 1571 553
rect 111 531 115 535
rect 1567 531 1571 535
rect 835 523 839 527
rect 727 514 731 518
rect 751 515 755 519
rect 847 514 851 518
rect 1091 523 1095 527
rect 975 514 979 518
rect 915 507 919 511
rect 1111 514 1115 518
rect 1255 514 1259 518
rect 1187 507 1191 511
rect 1407 514 1411 518
rect 1471 515 1472 519
rect 1472 515 1475 519
rect 767 478 771 482
rect 855 478 859 482
rect 943 478 947 482
rect 871 467 875 471
rect 1031 478 1035 482
rect 1119 478 1123 482
rect 959 467 963 471
rect 1207 478 1211 482
rect 1047 467 1051 471
rect 1295 478 1299 482
rect 1223 467 1227 471
rect 1383 478 1387 482
rect 1311 467 1315 471
rect 1471 478 1475 482
rect 1495 479 1499 483
rect 1399 467 1403 471
rect 1487 467 1491 471
rect 111 461 115 465
rect 1567 461 1571 465
rect 111 443 115 447
rect 935 447 939 451
rect 1567 443 1571 447
rect 767 432 771 436
rect 855 432 859 436
rect 871 431 875 435
rect 943 432 947 436
rect 959 431 963 435
rect 1031 432 1035 436
rect 1047 431 1051 435
rect 1119 432 1123 436
rect 1187 435 1191 439
rect 1207 432 1211 436
rect 1223 431 1227 435
rect 1295 432 1299 436
rect 1311 431 1315 435
rect 1383 432 1387 436
rect 1399 431 1403 435
rect 1471 432 1475 436
rect 1487 431 1491 435
rect 623 404 627 408
rect 699 403 703 407
rect 711 404 715 408
rect 799 404 803 408
rect 887 404 891 408
rect 919 403 923 407
rect 111 393 115 397
rect 1567 393 1571 397
rect 691 387 695 391
rect 779 387 783 391
rect 111 375 115 379
rect 1567 375 1571 379
rect 623 358 627 362
rect 691 359 692 363
rect 692 359 695 363
rect 711 358 715 362
rect 779 359 780 363
rect 780 359 783 363
rect 799 358 803 362
rect 887 358 891 362
rect 935 359 939 363
rect 919 351 923 355
rect 399 318 403 322
rect 487 318 491 322
rect 575 318 579 322
rect 503 307 507 311
rect 663 318 667 322
rect 699 319 703 323
rect 591 307 595 311
rect 679 307 683 311
rect 111 301 115 305
rect 1567 301 1571 305
rect 111 283 115 287
rect 1567 283 1571 287
rect 399 272 403 276
rect 467 271 471 275
rect 487 272 491 276
rect 503 271 507 275
rect 575 272 579 276
rect 591 271 595 275
rect 663 272 667 276
rect 679 271 683 275
rect 215 240 219 244
rect 275 239 279 243
rect 303 240 307 244
rect 391 240 395 244
rect 479 240 483 244
rect 111 229 115 233
rect 1567 229 1571 233
rect 283 223 287 227
rect 371 223 375 227
rect 459 223 463 227
rect 111 211 115 215
rect 1567 211 1571 215
rect 467 203 471 207
rect 215 194 219 198
rect 283 195 284 199
rect 284 195 287 199
rect 303 194 307 198
rect 371 195 372 199
rect 372 195 375 199
rect 391 194 395 198
rect 459 195 460 199
rect 460 195 463 199
rect 479 194 483 198
rect 135 138 139 142
rect 223 138 227 142
rect 311 138 315 142
rect 239 127 243 131
rect 399 138 403 142
rect 327 127 331 131
rect 487 138 491 142
rect 415 127 419 131
rect 575 138 579 142
rect 599 139 603 143
rect 503 127 507 131
rect 591 127 595 131
rect 111 121 115 125
rect 1567 121 1571 125
rect 111 103 115 107
rect 1567 103 1571 107
rect 135 92 139 96
rect 223 92 227 96
rect 239 91 243 95
rect 311 92 315 96
rect 327 91 331 95
rect 399 92 403 96
rect 415 91 419 95
rect 487 92 491 96
rect 503 91 507 95
rect 575 92 579 96
rect 591 91 595 95
<< m3 >>
rect 111 1530 115 1531
rect 111 1525 115 1526
rect 543 1530 547 1531
rect 543 1525 547 1526
rect 631 1530 635 1531
rect 631 1525 635 1526
rect 719 1530 723 1531
rect 719 1525 723 1526
rect 807 1530 811 1531
rect 807 1525 811 1526
rect 895 1530 899 1531
rect 895 1525 899 1526
rect 1567 1530 1571 1531
rect 1567 1525 1571 1526
rect 112 1502 114 1525
rect 544 1519 546 1525
rect 632 1519 634 1525
rect 720 1519 722 1525
rect 808 1519 810 1525
rect 896 1519 898 1525
rect 542 1518 548 1519
rect 542 1514 543 1518
rect 547 1514 548 1518
rect 542 1513 548 1514
rect 630 1518 636 1519
rect 630 1514 631 1518
rect 635 1514 636 1518
rect 630 1513 636 1514
rect 718 1518 724 1519
rect 718 1514 719 1518
rect 723 1514 724 1518
rect 718 1513 724 1514
rect 806 1518 812 1519
rect 806 1514 807 1518
rect 811 1514 812 1518
rect 894 1518 900 1519
rect 806 1513 812 1514
rect 886 1515 892 1516
rect 886 1511 887 1515
rect 891 1511 892 1515
rect 894 1514 895 1518
rect 899 1514 900 1518
rect 894 1513 900 1514
rect 974 1515 980 1516
rect 886 1510 892 1511
rect 974 1511 975 1515
rect 979 1511 980 1515
rect 974 1510 980 1511
rect 646 1507 652 1508
rect 646 1503 647 1507
rect 651 1503 652 1507
rect 646 1502 652 1503
rect 734 1507 740 1508
rect 734 1503 735 1507
rect 739 1503 740 1507
rect 734 1502 740 1503
rect 822 1507 828 1508
rect 822 1503 823 1507
rect 827 1503 828 1507
rect 822 1502 828 1503
rect 110 1501 116 1502
rect 110 1497 111 1501
rect 115 1497 116 1501
rect 110 1496 116 1497
rect 110 1483 116 1484
rect 110 1479 111 1483
rect 115 1479 116 1483
rect 110 1478 116 1479
rect 112 1467 114 1478
rect 542 1472 548 1473
rect 630 1472 636 1473
rect 648 1472 650 1502
rect 718 1472 724 1473
rect 736 1472 738 1502
rect 806 1472 812 1473
rect 824 1472 826 1502
rect 888 1488 890 1510
rect 886 1487 892 1488
rect 886 1483 887 1487
rect 891 1483 892 1487
rect 886 1482 892 1483
rect 894 1472 900 1473
rect 542 1468 543 1472
rect 547 1468 548 1472
rect 542 1467 548 1468
rect 622 1471 628 1472
rect 622 1467 623 1471
rect 627 1467 628 1471
rect 630 1468 631 1472
rect 635 1468 636 1472
rect 630 1467 636 1468
rect 646 1471 652 1472
rect 646 1467 647 1471
rect 651 1467 652 1471
rect 718 1468 719 1472
rect 723 1468 724 1472
rect 718 1467 724 1468
rect 734 1471 740 1472
rect 734 1467 735 1471
rect 739 1467 740 1471
rect 806 1468 807 1472
rect 811 1468 812 1472
rect 806 1467 812 1468
rect 822 1471 828 1472
rect 822 1467 823 1471
rect 827 1467 828 1471
rect 894 1468 895 1472
rect 899 1468 900 1472
rect 894 1467 900 1468
rect 111 1466 115 1467
rect 111 1461 115 1462
rect 471 1466 475 1467
rect 471 1461 475 1462
rect 543 1466 547 1467
rect 543 1461 547 1462
rect 615 1466 619 1467
rect 622 1466 628 1467
rect 631 1466 635 1467
rect 646 1466 652 1467
rect 719 1466 723 1467
rect 734 1466 740 1467
rect 775 1466 779 1467
rect 615 1461 619 1462
rect 112 1450 114 1461
rect 470 1460 476 1461
rect 614 1460 620 1461
rect 470 1456 471 1460
rect 475 1456 476 1460
rect 470 1455 476 1456
rect 502 1459 508 1460
rect 502 1455 503 1459
rect 507 1455 508 1459
rect 614 1456 615 1460
rect 619 1456 620 1460
rect 614 1455 620 1456
rect 502 1454 508 1455
rect 110 1449 116 1450
rect 110 1445 111 1449
rect 115 1445 116 1449
rect 110 1444 116 1445
rect 110 1431 116 1432
rect 110 1427 111 1431
rect 115 1427 116 1431
rect 110 1426 116 1427
rect 112 1399 114 1426
rect 470 1414 476 1415
rect 470 1410 471 1414
rect 475 1410 476 1414
rect 470 1409 476 1410
rect 472 1399 474 1409
rect 111 1398 115 1399
rect 111 1393 115 1394
rect 423 1398 427 1399
rect 423 1393 427 1394
rect 471 1398 475 1399
rect 471 1393 475 1394
rect 112 1370 114 1393
rect 424 1387 426 1393
rect 504 1388 506 1454
rect 538 1443 544 1444
rect 538 1439 539 1443
rect 543 1439 544 1443
rect 538 1438 544 1439
rect 540 1416 542 1438
rect 538 1415 544 1416
rect 538 1411 539 1415
rect 543 1411 544 1415
rect 538 1410 544 1411
rect 614 1414 620 1415
rect 614 1410 615 1414
rect 619 1410 620 1414
rect 614 1409 620 1410
rect 616 1399 618 1409
rect 624 1408 626 1466
rect 631 1461 635 1462
rect 719 1461 723 1462
rect 775 1461 779 1462
rect 807 1466 811 1467
rect 822 1466 828 1467
rect 895 1466 899 1467
rect 807 1461 811 1462
rect 895 1461 899 1462
rect 943 1466 947 1467
rect 943 1461 947 1462
rect 774 1460 780 1461
rect 774 1456 775 1460
rect 779 1456 780 1460
rect 774 1455 780 1456
rect 942 1460 948 1461
rect 976 1460 978 1510
rect 1568 1502 1570 1525
rect 1566 1501 1572 1502
rect 1566 1497 1567 1501
rect 1571 1497 1572 1501
rect 1566 1496 1572 1497
rect 1566 1483 1572 1484
rect 1566 1479 1567 1483
rect 1571 1479 1572 1483
rect 1566 1478 1572 1479
rect 1568 1467 1570 1478
rect 1119 1466 1123 1467
rect 1119 1461 1123 1462
rect 1303 1466 1307 1467
rect 1303 1461 1307 1462
rect 1471 1466 1475 1467
rect 1471 1461 1475 1462
rect 1567 1466 1571 1467
rect 1567 1461 1571 1462
rect 1118 1460 1124 1461
rect 942 1456 943 1460
rect 947 1456 948 1460
rect 942 1455 948 1456
rect 974 1459 980 1460
rect 974 1455 975 1459
rect 979 1455 980 1459
rect 1118 1456 1119 1460
rect 1123 1456 1124 1460
rect 1118 1455 1124 1456
rect 1302 1460 1308 1461
rect 1470 1460 1476 1461
rect 1302 1456 1303 1460
rect 1307 1456 1308 1460
rect 1302 1455 1308 1456
rect 1434 1459 1440 1460
rect 1434 1455 1435 1459
rect 1439 1455 1440 1459
rect 1470 1456 1471 1460
rect 1475 1456 1476 1460
rect 1470 1455 1476 1456
rect 1494 1459 1500 1460
rect 1494 1455 1495 1459
rect 1499 1455 1500 1459
rect 974 1454 980 1455
rect 1434 1454 1440 1455
rect 1494 1454 1500 1455
rect 682 1443 688 1444
rect 682 1439 683 1443
rect 687 1439 688 1443
rect 682 1438 688 1439
rect 1010 1443 1016 1444
rect 1010 1439 1011 1443
rect 1015 1439 1016 1443
rect 1010 1438 1016 1439
rect 684 1416 686 1438
rect 1012 1416 1014 1438
rect 1436 1424 1438 1454
rect 1434 1423 1440 1424
rect 1434 1419 1435 1423
rect 1439 1419 1440 1423
rect 1434 1418 1440 1419
rect 682 1415 688 1416
rect 1010 1415 1016 1416
rect 1198 1415 1204 1416
rect 682 1411 683 1415
rect 687 1411 688 1415
rect 682 1410 688 1411
rect 774 1414 780 1415
rect 774 1410 775 1414
rect 779 1410 780 1414
rect 774 1409 780 1410
rect 942 1414 948 1415
rect 942 1410 943 1414
rect 947 1410 948 1414
rect 1010 1411 1011 1415
rect 1015 1411 1016 1415
rect 1010 1410 1016 1411
rect 1118 1414 1124 1415
rect 1118 1410 1119 1414
rect 1123 1410 1124 1414
rect 1198 1411 1199 1415
rect 1203 1411 1204 1415
rect 1198 1410 1204 1411
rect 1302 1414 1308 1415
rect 1302 1410 1303 1414
rect 1307 1410 1308 1414
rect 942 1409 948 1410
rect 1118 1409 1124 1410
rect 622 1407 628 1408
rect 622 1403 623 1407
rect 627 1403 628 1407
rect 622 1402 628 1403
rect 776 1399 778 1409
rect 944 1399 946 1409
rect 1120 1399 1122 1409
rect 615 1398 619 1399
rect 615 1393 619 1394
rect 663 1398 667 1399
rect 663 1393 667 1394
rect 775 1398 779 1399
rect 775 1393 779 1394
rect 911 1398 915 1399
rect 911 1393 915 1394
rect 943 1398 947 1399
rect 943 1393 947 1394
rect 1119 1398 1123 1399
rect 1119 1393 1123 1394
rect 1167 1398 1171 1399
rect 1167 1393 1171 1394
rect 502 1387 508 1388
rect 664 1387 666 1393
rect 912 1387 914 1393
rect 1168 1387 1170 1393
rect 422 1386 428 1387
rect 422 1382 423 1386
rect 427 1382 428 1386
rect 502 1383 503 1387
rect 507 1383 508 1387
rect 502 1382 508 1383
rect 662 1386 668 1387
rect 662 1382 663 1386
rect 667 1382 668 1386
rect 422 1381 428 1382
rect 662 1381 668 1382
rect 910 1386 916 1387
rect 910 1382 911 1386
rect 915 1382 916 1386
rect 1166 1386 1172 1387
rect 910 1381 916 1382
rect 978 1383 984 1384
rect 978 1379 979 1383
rect 983 1379 984 1383
rect 1166 1382 1167 1386
rect 1171 1382 1172 1386
rect 1166 1381 1172 1382
rect 978 1378 984 1379
rect 590 1375 596 1376
rect 590 1371 591 1375
rect 595 1371 596 1375
rect 590 1370 596 1371
rect 110 1369 116 1370
rect 110 1365 111 1369
rect 115 1365 116 1369
rect 110 1364 116 1365
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 110 1346 116 1347
rect 112 1323 114 1346
rect 422 1340 428 1341
rect 592 1340 594 1370
rect 980 1360 982 1378
rect 730 1359 736 1360
rect 730 1355 731 1359
rect 735 1355 736 1359
rect 730 1354 736 1355
rect 978 1359 984 1360
rect 978 1355 979 1359
rect 983 1355 984 1359
rect 978 1354 984 1355
rect 732 1344 734 1354
rect 730 1343 736 1344
rect 662 1340 668 1341
rect 422 1336 423 1340
rect 427 1336 428 1340
rect 422 1335 428 1336
rect 590 1339 596 1340
rect 590 1335 591 1339
rect 595 1335 596 1339
rect 662 1336 663 1340
rect 667 1336 668 1340
rect 730 1339 731 1343
rect 735 1339 736 1343
rect 730 1338 736 1339
rect 910 1340 916 1341
rect 662 1335 668 1336
rect 910 1336 911 1340
rect 915 1336 916 1340
rect 910 1335 916 1336
rect 1166 1340 1172 1341
rect 1200 1340 1202 1410
rect 1302 1409 1308 1410
rect 1470 1414 1476 1415
rect 1470 1410 1471 1414
rect 1475 1410 1476 1414
rect 1470 1409 1476 1410
rect 1304 1399 1306 1409
rect 1472 1399 1474 1409
rect 1303 1398 1307 1399
rect 1303 1393 1307 1394
rect 1431 1398 1435 1399
rect 1431 1393 1435 1394
rect 1471 1398 1475 1399
rect 1471 1393 1475 1394
rect 1432 1387 1434 1393
rect 1496 1388 1498 1454
rect 1568 1450 1570 1461
rect 1566 1449 1572 1450
rect 1566 1445 1567 1449
rect 1571 1445 1572 1449
rect 1566 1444 1572 1445
rect 1566 1431 1572 1432
rect 1566 1427 1567 1431
rect 1571 1427 1572 1431
rect 1566 1426 1572 1427
rect 1568 1399 1570 1426
rect 1567 1398 1571 1399
rect 1567 1393 1571 1394
rect 1494 1387 1500 1388
rect 1430 1386 1436 1387
rect 1206 1383 1212 1384
rect 1206 1379 1207 1383
rect 1211 1379 1212 1383
rect 1430 1382 1431 1386
rect 1435 1382 1436 1386
rect 1494 1383 1495 1387
rect 1499 1383 1500 1387
rect 1494 1382 1500 1383
rect 1430 1381 1436 1382
rect 1206 1378 1212 1379
rect 1166 1336 1167 1340
rect 1171 1336 1172 1340
rect 1166 1335 1172 1336
rect 1198 1339 1204 1340
rect 1198 1335 1199 1339
rect 1203 1335 1204 1339
rect 424 1323 426 1335
rect 590 1334 596 1335
rect 664 1323 666 1335
rect 854 1331 860 1332
rect 854 1327 855 1331
rect 859 1327 860 1331
rect 854 1326 860 1327
rect 111 1322 115 1323
rect 111 1317 115 1318
rect 423 1322 427 1323
rect 423 1317 427 1318
rect 487 1322 491 1323
rect 487 1317 491 1318
rect 663 1322 667 1323
rect 663 1317 667 1318
rect 727 1322 731 1323
rect 727 1317 731 1318
rect 112 1306 114 1317
rect 486 1316 492 1317
rect 726 1316 732 1317
rect 486 1312 487 1316
rect 491 1312 492 1316
rect 486 1311 492 1312
rect 562 1315 568 1316
rect 562 1311 563 1315
rect 567 1311 568 1315
rect 726 1312 727 1316
rect 731 1312 732 1316
rect 726 1311 732 1312
rect 562 1310 568 1311
rect 110 1305 116 1306
rect 110 1301 111 1305
rect 115 1301 116 1305
rect 110 1300 116 1301
rect 554 1299 560 1300
rect 554 1295 555 1299
rect 559 1295 560 1299
rect 554 1294 560 1295
rect 110 1287 116 1288
rect 110 1283 111 1287
rect 115 1283 116 1287
rect 110 1282 116 1283
rect 112 1247 114 1282
rect 556 1272 558 1294
rect 554 1271 560 1272
rect 486 1270 492 1271
rect 486 1266 487 1270
rect 491 1266 492 1270
rect 554 1267 555 1271
rect 559 1267 560 1271
rect 554 1266 560 1267
rect 486 1265 492 1266
rect 488 1247 490 1265
rect 111 1246 115 1247
rect 111 1241 115 1242
rect 487 1246 491 1247
rect 487 1241 491 1242
rect 535 1246 539 1247
rect 535 1241 539 1242
rect 112 1218 114 1241
rect 536 1235 538 1241
rect 564 1236 566 1310
rect 856 1272 858 1326
rect 912 1323 914 1335
rect 1168 1323 1170 1335
rect 1198 1334 1204 1335
rect 911 1322 915 1323
rect 911 1317 915 1318
rect 967 1322 971 1323
rect 967 1317 971 1318
rect 1167 1322 1171 1323
rect 1167 1317 1171 1318
rect 966 1316 972 1317
rect 1208 1316 1210 1378
rect 1568 1370 1570 1393
rect 1566 1369 1572 1370
rect 1566 1365 1567 1369
rect 1571 1365 1572 1369
rect 1566 1364 1572 1365
rect 1566 1351 1572 1352
rect 1566 1347 1567 1351
rect 1571 1347 1572 1351
rect 1566 1346 1572 1347
rect 1430 1340 1436 1341
rect 1430 1336 1431 1340
rect 1435 1336 1436 1340
rect 1430 1335 1436 1336
rect 1498 1339 1504 1340
rect 1498 1335 1499 1339
rect 1503 1335 1504 1339
rect 1432 1323 1434 1335
rect 1498 1334 1504 1335
rect 1215 1322 1219 1323
rect 1215 1317 1219 1318
rect 1431 1322 1435 1323
rect 1431 1317 1435 1318
rect 1463 1322 1467 1323
rect 1463 1317 1467 1318
rect 1214 1316 1220 1317
rect 1462 1316 1468 1317
rect 966 1312 967 1316
rect 971 1312 972 1316
rect 966 1311 972 1312
rect 1206 1315 1212 1316
rect 1206 1311 1207 1315
rect 1211 1311 1212 1315
rect 1214 1312 1215 1316
rect 1219 1312 1220 1316
rect 1214 1311 1220 1312
rect 1422 1315 1428 1316
rect 1422 1311 1423 1315
rect 1427 1311 1428 1315
rect 1462 1312 1463 1316
rect 1467 1312 1468 1316
rect 1462 1311 1468 1312
rect 1206 1310 1212 1311
rect 1422 1310 1428 1311
rect 1282 1299 1288 1300
rect 1282 1295 1283 1299
rect 1287 1295 1288 1299
rect 1282 1294 1288 1295
rect 1284 1272 1286 1294
rect 854 1271 860 1272
rect 1206 1271 1212 1272
rect 1282 1271 1288 1272
rect 726 1270 732 1271
rect 726 1266 727 1270
rect 731 1266 732 1270
rect 854 1267 855 1271
rect 859 1267 860 1271
rect 854 1266 860 1267
rect 966 1270 972 1271
rect 966 1266 967 1270
rect 971 1266 972 1270
rect 1206 1267 1207 1271
rect 1211 1267 1212 1271
rect 1206 1266 1212 1267
rect 1214 1270 1220 1271
rect 1214 1266 1215 1270
rect 1219 1266 1220 1270
rect 1282 1267 1283 1271
rect 1287 1267 1288 1271
rect 1282 1266 1288 1267
rect 726 1265 732 1266
rect 966 1265 972 1266
rect 728 1247 730 1265
rect 968 1247 970 1265
rect 727 1246 731 1247
rect 727 1241 731 1242
rect 743 1246 747 1247
rect 743 1241 747 1242
rect 959 1246 963 1247
rect 959 1241 963 1242
rect 967 1246 971 1247
rect 967 1241 971 1242
rect 1175 1246 1179 1247
rect 1175 1241 1179 1242
rect 562 1235 568 1236
rect 744 1235 746 1241
rect 960 1235 962 1241
rect 1176 1235 1178 1241
rect 534 1234 540 1235
rect 534 1230 535 1234
rect 539 1230 540 1234
rect 562 1231 563 1235
rect 567 1231 568 1235
rect 562 1230 568 1231
rect 742 1234 748 1235
rect 742 1230 743 1234
rect 747 1230 748 1234
rect 534 1229 540 1230
rect 742 1229 748 1230
rect 958 1234 964 1235
rect 958 1230 959 1234
rect 963 1230 964 1234
rect 1174 1234 1180 1235
rect 958 1229 964 1230
rect 982 1231 988 1232
rect 982 1227 983 1231
rect 987 1227 988 1231
rect 1174 1230 1175 1234
rect 1179 1230 1180 1234
rect 1174 1229 1180 1230
rect 982 1226 988 1227
rect 686 1223 692 1224
rect 686 1219 687 1223
rect 691 1219 692 1223
rect 686 1218 692 1219
rect 110 1217 116 1218
rect 110 1213 111 1217
rect 115 1213 116 1217
rect 110 1212 116 1213
rect 110 1199 116 1200
rect 110 1195 111 1199
rect 115 1195 116 1199
rect 110 1194 116 1195
rect 112 1167 114 1194
rect 534 1188 540 1189
rect 688 1188 690 1218
rect 742 1188 748 1189
rect 534 1184 535 1188
rect 539 1184 540 1188
rect 534 1183 540 1184
rect 686 1187 692 1188
rect 686 1183 687 1187
rect 691 1183 692 1187
rect 742 1184 743 1188
rect 747 1184 748 1188
rect 742 1183 748 1184
rect 958 1188 964 1189
rect 958 1184 959 1188
rect 963 1184 964 1188
rect 958 1183 964 1184
rect 536 1167 538 1183
rect 686 1182 692 1183
rect 744 1167 746 1183
rect 960 1167 962 1183
rect 984 1180 986 1226
rect 1174 1188 1180 1189
rect 1208 1188 1210 1266
rect 1214 1265 1220 1266
rect 1216 1247 1218 1265
rect 1215 1246 1219 1247
rect 1215 1241 1219 1242
rect 1399 1246 1403 1247
rect 1399 1241 1403 1242
rect 1400 1235 1402 1241
rect 1424 1236 1426 1310
rect 1500 1272 1502 1334
rect 1568 1323 1570 1346
rect 1567 1322 1571 1323
rect 1567 1317 1571 1318
rect 1568 1306 1570 1317
rect 1566 1305 1572 1306
rect 1566 1301 1567 1305
rect 1571 1301 1572 1305
rect 1566 1300 1572 1301
rect 1566 1287 1572 1288
rect 1566 1283 1567 1287
rect 1571 1283 1572 1287
rect 1566 1282 1572 1283
rect 1498 1271 1504 1272
rect 1462 1270 1468 1271
rect 1462 1266 1463 1270
rect 1467 1266 1468 1270
rect 1498 1267 1499 1271
rect 1503 1267 1504 1271
rect 1498 1266 1504 1267
rect 1462 1265 1468 1266
rect 1464 1247 1466 1265
rect 1568 1247 1570 1282
rect 1463 1246 1467 1247
rect 1463 1241 1467 1242
rect 1567 1246 1571 1247
rect 1567 1241 1571 1242
rect 1422 1235 1428 1236
rect 1398 1234 1404 1235
rect 1238 1231 1244 1232
rect 1238 1227 1239 1231
rect 1243 1227 1244 1231
rect 1398 1230 1399 1234
rect 1403 1230 1404 1234
rect 1422 1231 1423 1235
rect 1427 1231 1428 1235
rect 1422 1230 1428 1231
rect 1398 1229 1404 1230
rect 1238 1226 1244 1227
rect 1038 1187 1044 1188
rect 1038 1183 1039 1187
rect 1043 1183 1044 1187
rect 1174 1184 1175 1188
rect 1179 1184 1180 1188
rect 1174 1183 1180 1184
rect 1206 1187 1212 1188
rect 1206 1183 1207 1187
rect 1211 1183 1212 1187
rect 1038 1182 1044 1183
rect 982 1179 988 1180
rect 982 1175 983 1179
rect 987 1175 988 1179
rect 982 1174 988 1175
rect 111 1166 115 1167
rect 111 1161 115 1162
rect 535 1166 539 1167
rect 535 1161 539 1162
rect 655 1166 659 1167
rect 655 1161 659 1162
rect 743 1166 747 1167
rect 743 1161 747 1162
rect 831 1166 835 1167
rect 831 1161 835 1162
rect 959 1166 963 1167
rect 959 1161 963 1162
rect 1015 1166 1019 1167
rect 1015 1161 1019 1162
rect 112 1150 114 1161
rect 654 1160 660 1161
rect 830 1160 836 1161
rect 654 1156 655 1160
rect 659 1156 660 1160
rect 654 1155 660 1156
rect 730 1159 736 1160
rect 730 1155 731 1159
rect 735 1155 736 1159
rect 830 1156 831 1160
rect 835 1156 836 1160
rect 830 1155 836 1156
rect 1014 1160 1020 1161
rect 1014 1156 1015 1160
rect 1019 1156 1020 1160
rect 1014 1155 1020 1156
rect 730 1154 736 1155
rect 110 1149 116 1150
rect 110 1145 111 1149
rect 115 1145 116 1149
rect 110 1144 116 1145
rect 722 1143 728 1144
rect 722 1139 723 1143
rect 727 1139 728 1143
rect 722 1138 728 1139
rect 110 1131 116 1132
rect 110 1127 111 1131
rect 115 1127 116 1131
rect 110 1126 116 1127
rect 112 1091 114 1126
rect 724 1116 726 1138
rect 722 1115 728 1116
rect 654 1114 660 1115
rect 654 1110 655 1114
rect 659 1110 660 1114
rect 722 1111 723 1115
rect 727 1111 728 1115
rect 722 1110 728 1111
rect 654 1109 660 1110
rect 656 1091 658 1109
rect 111 1090 115 1091
rect 111 1085 115 1086
rect 655 1090 659 1091
rect 655 1085 659 1086
rect 663 1090 667 1091
rect 663 1085 667 1086
rect 112 1062 114 1085
rect 664 1079 666 1085
rect 732 1080 734 1154
rect 954 1143 960 1144
rect 954 1139 955 1143
rect 959 1139 960 1143
rect 954 1138 960 1139
rect 956 1116 958 1138
rect 1040 1116 1042 1182
rect 1176 1167 1178 1183
rect 1206 1182 1212 1183
rect 1175 1166 1179 1167
rect 1175 1161 1179 1162
rect 1207 1166 1211 1167
rect 1207 1161 1211 1162
rect 1206 1160 1212 1161
rect 1240 1160 1242 1226
rect 1568 1218 1570 1241
rect 1566 1217 1572 1218
rect 1566 1213 1567 1217
rect 1571 1213 1572 1217
rect 1566 1212 1572 1213
rect 1566 1199 1572 1200
rect 1566 1195 1567 1199
rect 1571 1195 1572 1199
rect 1566 1194 1572 1195
rect 1398 1188 1404 1189
rect 1398 1184 1399 1188
rect 1403 1184 1404 1188
rect 1398 1183 1404 1184
rect 1462 1187 1468 1188
rect 1462 1183 1463 1187
rect 1467 1183 1468 1187
rect 1400 1167 1402 1183
rect 1462 1182 1468 1183
rect 1399 1166 1403 1167
rect 1399 1161 1403 1162
rect 1398 1160 1404 1161
rect 1206 1156 1207 1160
rect 1211 1156 1212 1160
rect 1206 1155 1212 1156
rect 1238 1159 1244 1160
rect 1238 1155 1239 1159
rect 1243 1155 1244 1159
rect 1398 1156 1399 1160
rect 1403 1156 1404 1160
rect 1398 1155 1404 1156
rect 1238 1154 1244 1155
rect 1464 1116 1466 1182
rect 1568 1167 1570 1194
rect 1567 1166 1571 1167
rect 1567 1161 1571 1162
rect 1474 1159 1480 1160
rect 1474 1155 1475 1159
rect 1479 1155 1480 1159
rect 1474 1154 1480 1155
rect 954 1115 960 1116
rect 1038 1115 1044 1116
rect 1270 1115 1276 1116
rect 1462 1115 1468 1116
rect 830 1114 836 1115
rect 830 1110 831 1114
rect 835 1110 836 1114
rect 954 1111 955 1115
rect 959 1111 960 1115
rect 954 1110 960 1111
rect 1014 1114 1020 1115
rect 1014 1110 1015 1114
rect 1019 1110 1020 1114
rect 1038 1111 1039 1115
rect 1043 1111 1044 1115
rect 1038 1110 1044 1111
rect 1206 1114 1212 1115
rect 1206 1110 1207 1114
rect 1211 1110 1212 1114
rect 1270 1111 1271 1115
rect 1275 1111 1276 1115
rect 1270 1110 1276 1111
rect 1398 1114 1404 1115
rect 1398 1110 1399 1114
rect 1403 1110 1404 1114
rect 1462 1111 1463 1115
rect 1467 1111 1468 1115
rect 1462 1110 1468 1111
rect 830 1109 836 1110
rect 1014 1109 1020 1110
rect 1206 1109 1212 1110
rect 832 1091 834 1109
rect 1016 1091 1018 1109
rect 1208 1091 1210 1109
rect 831 1090 835 1091
rect 831 1085 835 1086
rect 847 1090 851 1091
rect 847 1085 851 1086
rect 1015 1090 1019 1091
rect 1015 1085 1019 1086
rect 1031 1090 1035 1091
rect 1031 1085 1035 1086
rect 1207 1090 1211 1091
rect 1207 1085 1211 1086
rect 1223 1090 1227 1091
rect 1223 1085 1227 1086
rect 730 1079 736 1080
rect 848 1079 850 1085
rect 1032 1079 1034 1085
rect 1224 1079 1226 1085
rect 662 1078 668 1079
rect 662 1074 663 1078
rect 667 1074 668 1078
rect 730 1075 731 1079
rect 735 1075 736 1079
rect 730 1074 736 1075
rect 846 1078 852 1079
rect 846 1074 847 1078
rect 851 1074 852 1078
rect 662 1073 668 1074
rect 846 1073 852 1074
rect 1030 1078 1036 1079
rect 1030 1074 1031 1078
rect 1035 1074 1036 1078
rect 1222 1078 1228 1079
rect 1030 1073 1036 1074
rect 1098 1075 1104 1076
rect 1098 1071 1099 1075
rect 1103 1071 1104 1075
rect 1222 1074 1223 1078
rect 1227 1074 1228 1078
rect 1222 1073 1228 1074
rect 1098 1070 1104 1071
rect 802 1067 808 1068
rect 802 1063 803 1067
rect 807 1063 808 1067
rect 802 1062 808 1063
rect 110 1061 116 1062
rect 110 1057 111 1061
rect 115 1057 116 1061
rect 110 1056 116 1057
rect 110 1043 116 1044
rect 110 1039 111 1043
rect 115 1039 116 1043
rect 110 1038 116 1039
rect 112 1011 114 1038
rect 662 1032 668 1033
rect 804 1032 806 1062
rect 1100 1052 1102 1070
rect 914 1051 920 1052
rect 914 1047 915 1051
rect 919 1047 920 1051
rect 914 1046 920 1047
rect 1098 1051 1104 1052
rect 1098 1047 1099 1051
rect 1103 1047 1104 1051
rect 1098 1046 1104 1047
rect 916 1036 918 1046
rect 914 1035 920 1036
rect 846 1032 852 1033
rect 662 1028 663 1032
rect 667 1028 668 1032
rect 662 1027 668 1028
rect 802 1031 808 1032
rect 802 1027 803 1031
rect 807 1027 808 1031
rect 846 1028 847 1032
rect 851 1028 852 1032
rect 914 1031 915 1035
rect 919 1031 920 1035
rect 914 1030 920 1031
rect 1030 1032 1036 1033
rect 1222 1032 1228 1033
rect 1272 1032 1274 1110
rect 1398 1109 1404 1110
rect 1400 1091 1402 1109
rect 1399 1090 1403 1091
rect 1399 1085 1403 1086
rect 1423 1090 1427 1091
rect 1423 1085 1427 1086
rect 1424 1079 1426 1085
rect 1476 1080 1478 1154
rect 1568 1150 1570 1161
rect 1566 1149 1572 1150
rect 1566 1145 1567 1149
rect 1571 1145 1572 1149
rect 1566 1144 1572 1145
rect 1566 1131 1572 1132
rect 1566 1127 1567 1131
rect 1571 1127 1572 1131
rect 1566 1126 1572 1127
rect 1568 1091 1570 1126
rect 1567 1090 1571 1091
rect 1567 1085 1571 1086
rect 1474 1079 1480 1080
rect 1422 1078 1428 1079
rect 1286 1075 1292 1076
rect 1286 1071 1287 1075
rect 1291 1071 1292 1075
rect 1422 1074 1423 1078
rect 1427 1074 1428 1078
rect 1474 1075 1475 1079
rect 1479 1075 1480 1079
rect 1474 1074 1480 1075
rect 1422 1073 1428 1074
rect 1286 1070 1292 1071
rect 846 1027 852 1028
rect 1030 1028 1031 1032
rect 1035 1028 1036 1032
rect 1030 1027 1036 1028
rect 1062 1031 1068 1032
rect 1062 1027 1063 1031
rect 1067 1027 1068 1031
rect 1222 1028 1223 1032
rect 1227 1028 1228 1032
rect 1222 1027 1228 1028
rect 1270 1031 1276 1032
rect 1270 1027 1271 1031
rect 1275 1027 1276 1031
rect 664 1011 666 1027
rect 802 1026 808 1027
rect 848 1011 850 1027
rect 1032 1011 1034 1027
rect 1062 1026 1068 1027
rect 111 1010 115 1011
rect 111 1005 115 1006
rect 551 1010 555 1011
rect 551 1005 555 1006
rect 663 1010 667 1011
rect 663 1005 667 1006
rect 759 1010 763 1011
rect 759 1005 763 1006
rect 847 1010 851 1011
rect 847 1005 851 1006
rect 975 1010 979 1011
rect 975 1005 979 1006
rect 1031 1010 1035 1011
rect 1031 1005 1035 1006
rect 112 994 114 1005
rect 550 1004 556 1005
rect 758 1004 764 1005
rect 550 1000 551 1004
rect 555 1000 556 1004
rect 550 999 556 1000
rect 582 1003 588 1004
rect 582 999 583 1003
rect 587 999 588 1003
rect 758 1000 759 1004
rect 763 1000 764 1004
rect 758 999 764 1000
rect 974 1004 980 1005
rect 974 1000 975 1004
rect 979 1000 980 1004
rect 974 999 980 1000
rect 1006 1003 1012 1004
rect 1006 999 1007 1003
rect 1011 999 1012 1003
rect 582 998 588 999
rect 1006 998 1012 999
rect 110 993 116 994
rect 110 989 111 993
rect 115 989 116 993
rect 110 988 116 989
rect 110 975 116 976
rect 110 971 111 975
rect 115 971 116 975
rect 110 970 116 971
rect 112 935 114 970
rect 550 958 556 959
rect 550 954 551 958
rect 555 954 556 958
rect 550 953 556 954
rect 552 935 554 953
rect 111 934 115 935
rect 111 929 115 930
rect 399 934 403 935
rect 399 929 403 930
rect 551 934 555 935
rect 551 929 555 930
rect 112 906 114 929
rect 400 923 402 929
rect 584 924 586 998
rect 618 987 624 988
rect 618 983 619 987
rect 623 983 624 987
rect 618 982 624 983
rect 620 960 622 982
rect 618 959 624 960
rect 618 955 619 959
rect 623 955 624 959
rect 618 954 624 955
rect 758 958 764 959
rect 758 954 759 958
rect 763 954 764 958
rect 758 953 764 954
rect 974 958 980 959
rect 974 954 975 958
rect 979 954 980 958
rect 974 953 980 954
rect 760 935 762 953
rect 976 935 978 953
rect 1008 952 1010 998
rect 1064 960 1066 1026
rect 1224 1011 1226 1027
rect 1270 1026 1276 1027
rect 1199 1010 1203 1011
rect 1199 1005 1203 1006
rect 1223 1010 1227 1011
rect 1223 1005 1227 1006
rect 1198 1004 1204 1005
rect 1288 1004 1290 1070
rect 1568 1062 1570 1085
rect 1566 1061 1572 1062
rect 1566 1057 1567 1061
rect 1571 1057 1572 1061
rect 1566 1056 1572 1057
rect 1566 1043 1572 1044
rect 1566 1039 1567 1043
rect 1571 1039 1572 1043
rect 1566 1038 1572 1039
rect 1422 1032 1428 1033
rect 1422 1028 1423 1032
rect 1427 1028 1428 1032
rect 1422 1027 1428 1028
rect 1490 1031 1496 1032
rect 1490 1027 1491 1031
rect 1495 1027 1496 1031
rect 1424 1011 1426 1027
rect 1490 1026 1496 1027
rect 1423 1010 1427 1011
rect 1423 1005 1427 1006
rect 1431 1010 1435 1011
rect 1431 1005 1435 1006
rect 1430 1004 1436 1005
rect 1198 1000 1199 1004
rect 1203 1000 1204 1004
rect 1198 999 1204 1000
rect 1286 1003 1292 1004
rect 1286 999 1287 1003
rect 1291 999 1292 1003
rect 1430 1000 1431 1004
rect 1435 1000 1436 1004
rect 1430 999 1436 1000
rect 1286 998 1292 999
rect 1492 960 1494 1026
rect 1568 1011 1570 1038
rect 1567 1010 1571 1011
rect 1567 1005 1571 1006
rect 1498 1003 1504 1004
rect 1498 999 1499 1003
rect 1503 999 1504 1003
rect 1498 998 1504 999
rect 1062 959 1068 960
rect 1266 959 1272 960
rect 1490 959 1496 960
rect 1062 955 1063 959
rect 1067 955 1068 959
rect 1062 954 1068 955
rect 1198 958 1204 959
rect 1198 954 1199 958
rect 1203 954 1204 958
rect 1266 955 1267 959
rect 1271 955 1272 959
rect 1266 954 1272 955
rect 1430 958 1436 959
rect 1430 954 1431 958
rect 1435 954 1436 958
rect 1490 955 1491 959
rect 1495 955 1496 959
rect 1490 954 1496 955
rect 1198 953 1204 954
rect 1006 951 1012 952
rect 1006 947 1007 951
rect 1011 947 1012 951
rect 1006 946 1012 947
rect 1200 935 1202 953
rect 663 934 667 935
rect 614 931 620 932
rect 614 927 615 931
rect 619 927 620 931
rect 663 929 667 930
rect 759 934 763 935
rect 927 934 931 935
rect 759 929 763 930
rect 854 931 860 932
rect 614 926 620 927
rect 582 923 588 924
rect 398 922 404 923
rect 398 918 399 922
rect 403 918 404 922
rect 582 919 583 923
rect 587 919 588 923
rect 582 918 588 919
rect 398 917 404 918
rect 110 905 116 906
rect 110 901 111 905
rect 115 901 116 905
rect 110 900 116 901
rect 110 887 116 888
rect 110 883 111 887
rect 115 883 116 887
rect 110 882 116 883
rect 112 859 114 882
rect 398 876 404 877
rect 616 876 618 926
rect 664 923 666 929
rect 854 927 855 931
rect 859 927 860 931
rect 927 929 931 930
rect 975 934 979 935
rect 975 929 979 930
rect 1199 934 1203 935
rect 1199 929 1203 930
rect 854 926 860 927
rect 662 922 668 923
rect 662 918 663 922
rect 667 918 668 922
rect 662 917 668 918
rect 662 876 668 877
rect 856 876 858 926
rect 928 923 930 929
rect 1200 923 1202 929
rect 926 922 932 923
rect 926 918 927 922
rect 931 918 932 922
rect 926 917 932 918
rect 1198 922 1204 923
rect 1198 918 1199 922
rect 1203 918 1204 922
rect 1198 917 1204 918
rect 926 876 932 877
rect 1198 876 1204 877
rect 398 872 399 876
rect 403 872 404 876
rect 398 871 404 872
rect 614 875 620 876
rect 614 871 615 875
rect 619 871 620 875
rect 662 872 663 876
rect 667 872 668 876
rect 662 871 668 872
rect 854 875 860 876
rect 854 871 855 875
rect 859 871 860 875
rect 926 872 927 876
rect 931 872 932 876
rect 926 871 932 872
rect 958 875 964 876
rect 958 871 959 875
rect 963 871 964 875
rect 1198 872 1199 876
rect 1203 872 1204 876
rect 1198 871 1204 872
rect 400 859 402 871
rect 614 870 620 871
rect 664 859 666 871
rect 854 870 860 871
rect 928 859 930 871
rect 958 870 964 871
rect 111 858 115 859
rect 111 853 115 854
rect 255 858 259 859
rect 255 853 259 854
rect 399 858 403 859
rect 399 853 403 854
rect 535 858 539 859
rect 535 853 539 854
rect 663 858 667 859
rect 663 853 667 854
rect 823 858 827 859
rect 823 853 827 854
rect 927 858 931 859
rect 927 853 931 854
rect 112 842 114 853
rect 254 852 260 853
rect 534 852 540 853
rect 254 848 255 852
rect 259 848 260 852
rect 254 847 260 848
rect 286 851 292 852
rect 286 847 287 851
rect 291 847 292 851
rect 534 848 535 852
rect 539 848 540 852
rect 534 847 540 848
rect 822 852 828 853
rect 822 848 823 852
rect 827 848 828 852
rect 822 847 828 848
rect 286 846 292 847
rect 110 841 116 842
rect 110 837 111 841
rect 115 837 116 841
rect 110 836 116 837
rect 110 823 116 824
rect 110 819 111 823
rect 115 819 116 823
rect 110 818 116 819
rect 112 783 114 818
rect 254 806 260 807
rect 254 802 255 806
rect 259 802 260 806
rect 254 801 260 802
rect 256 783 258 801
rect 111 782 115 783
rect 111 777 115 778
rect 199 782 203 783
rect 199 777 203 778
rect 255 782 259 783
rect 255 777 259 778
rect 112 754 114 777
rect 200 771 202 777
rect 288 772 290 846
rect 322 835 328 836
rect 322 831 323 835
rect 327 831 328 835
rect 322 830 328 831
rect 602 835 608 836
rect 602 831 603 835
rect 607 831 608 835
rect 602 830 608 831
rect 324 808 326 830
rect 604 808 606 830
rect 960 808 962 870
rect 1200 859 1202 871
rect 1111 858 1115 859
rect 1111 853 1115 854
rect 1199 858 1203 859
rect 1199 853 1203 854
rect 1110 852 1116 853
rect 1268 852 1270 954
rect 1430 953 1436 954
rect 1432 935 1434 953
rect 1431 934 1435 935
rect 1431 929 1435 930
rect 1471 934 1475 935
rect 1471 929 1475 930
rect 1472 923 1474 929
rect 1500 924 1502 998
rect 1568 994 1570 1005
rect 1566 993 1572 994
rect 1566 989 1567 993
rect 1571 989 1572 993
rect 1566 988 1572 989
rect 1566 975 1572 976
rect 1566 971 1567 975
rect 1571 971 1572 975
rect 1566 970 1572 971
rect 1568 935 1570 970
rect 1567 934 1571 935
rect 1567 929 1571 930
rect 1498 923 1504 924
rect 1470 922 1476 923
rect 1334 919 1340 920
rect 1334 915 1335 919
rect 1339 915 1340 919
rect 1470 918 1471 922
rect 1475 918 1476 922
rect 1498 919 1499 923
rect 1503 919 1504 923
rect 1498 918 1504 919
rect 1470 917 1476 918
rect 1334 914 1340 915
rect 1336 868 1338 914
rect 1568 906 1570 929
rect 1566 905 1572 906
rect 1566 901 1567 905
rect 1571 901 1572 905
rect 1566 900 1572 901
rect 1566 887 1572 888
rect 1566 883 1567 887
rect 1571 883 1572 887
rect 1566 882 1572 883
rect 1470 876 1476 877
rect 1430 875 1436 876
rect 1430 871 1431 875
rect 1435 871 1436 875
rect 1470 872 1471 876
rect 1475 872 1476 876
rect 1470 871 1476 872
rect 1430 870 1436 871
rect 1334 867 1340 868
rect 1334 863 1335 867
rect 1339 863 1340 867
rect 1334 862 1340 863
rect 1407 858 1411 859
rect 1407 853 1411 854
rect 1406 852 1412 853
rect 1110 848 1111 852
rect 1115 848 1116 852
rect 1110 847 1116 848
rect 1266 851 1272 852
rect 1266 847 1267 851
rect 1271 847 1272 851
rect 1406 848 1407 852
rect 1411 848 1412 852
rect 1406 847 1412 848
rect 1266 846 1272 847
rect 1432 808 1434 870
rect 1472 859 1474 871
rect 1568 859 1570 882
rect 1471 858 1475 859
rect 1471 853 1475 854
rect 1567 858 1571 859
rect 1567 853 1571 854
rect 1462 851 1468 852
rect 1462 847 1463 851
rect 1467 847 1468 851
rect 1462 846 1468 847
rect 322 807 328 808
rect 602 807 608 808
rect 958 807 964 808
rect 1154 807 1160 808
rect 1430 807 1436 808
rect 322 803 323 807
rect 327 803 328 807
rect 322 802 328 803
rect 534 806 540 807
rect 534 802 535 806
rect 539 802 540 806
rect 602 803 603 807
rect 607 803 608 807
rect 602 802 608 803
rect 822 806 828 807
rect 822 802 823 806
rect 827 802 828 806
rect 958 803 959 807
rect 963 803 964 807
rect 958 802 964 803
rect 1110 806 1116 807
rect 1110 802 1111 806
rect 1115 802 1116 806
rect 1154 803 1155 807
rect 1159 803 1160 807
rect 1154 802 1160 803
rect 1406 806 1412 807
rect 1406 802 1407 806
rect 1411 802 1412 806
rect 1430 803 1431 807
rect 1435 803 1436 807
rect 1430 802 1436 803
rect 534 801 540 802
rect 822 801 828 802
rect 1110 801 1116 802
rect 536 783 538 801
rect 824 783 826 801
rect 1112 783 1114 801
rect 487 782 491 783
rect 487 777 491 778
rect 535 782 539 783
rect 535 777 539 778
rect 783 782 787 783
rect 783 777 787 778
rect 823 782 827 783
rect 823 777 827 778
rect 1087 782 1091 783
rect 1087 777 1091 778
rect 1111 782 1115 783
rect 1111 777 1115 778
rect 286 771 292 772
rect 488 771 490 777
rect 784 771 786 777
rect 1088 771 1090 777
rect 198 770 204 771
rect 198 766 199 770
rect 203 766 204 770
rect 286 767 287 771
rect 291 767 292 771
rect 286 766 292 767
rect 486 770 492 771
rect 486 766 487 770
rect 491 766 492 770
rect 198 765 204 766
rect 486 765 492 766
rect 782 770 788 771
rect 782 766 783 770
rect 787 766 788 770
rect 1086 770 1092 771
rect 782 765 788 766
rect 850 767 856 768
rect 850 763 851 767
rect 855 763 856 767
rect 1086 766 1087 770
rect 1091 766 1092 770
rect 1086 765 1092 766
rect 850 762 856 763
rect 798 759 804 760
rect 798 755 799 759
rect 803 755 804 759
rect 798 754 804 755
rect 110 753 116 754
rect 110 749 111 753
rect 115 749 116 753
rect 110 748 116 749
rect 110 735 116 736
rect 110 731 111 735
rect 115 731 116 735
rect 110 730 116 731
rect 112 711 114 730
rect 198 724 204 725
rect 198 720 199 724
rect 203 720 204 724
rect 198 719 204 720
rect 486 724 492 725
rect 782 724 788 725
rect 800 724 802 754
rect 852 740 854 762
rect 850 739 856 740
rect 850 735 851 739
rect 855 735 856 739
rect 850 734 856 735
rect 1156 728 1158 802
rect 1406 801 1412 802
rect 1408 783 1410 801
rect 1399 782 1403 783
rect 1399 777 1403 778
rect 1407 782 1411 783
rect 1407 777 1411 778
rect 1400 771 1402 777
rect 1464 772 1466 846
rect 1568 842 1570 853
rect 1566 841 1572 842
rect 1566 837 1567 841
rect 1571 837 1572 841
rect 1566 836 1572 837
rect 1566 823 1572 824
rect 1566 819 1567 823
rect 1571 819 1572 823
rect 1566 818 1572 819
rect 1568 783 1570 818
rect 1567 782 1571 783
rect 1567 777 1571 778
rect 1462 771 1468 772
rect 1398 770 1404 771
rect 1222 767 1228 768
rect 1222 763 1223 767
rect 1227 763 1228 767
rect 1398 766 1399 770
rect 1403 766 1404 770
rect 1462 767 1463 771
rect 1467 767 1468 771
rect 1462 766 1468 767
rect 1398 765 1404 766
rect 1222 762 1228 763
rect 1154 727 1160 728
rect 1086 724 1092 725
rect 486 720 487 724
rect 491 720 492 724
rect 486 719 492 720
rect 518 723 524 724
rect 518 719 519 723
rect 523 719 524 723
rect 782 720 783 724
rect 787 720 788 724
rect 782 719 788 720
rect 798 723 804 724
rect 798 719 799 723
rect 803 719 804 723
rect 1086 720 1087 724
rect 1091 720 1092 724
rect 1154 723 1155 727
rect 1159 723 1160 727
rect 1154 722 1160 723
rect 1086 719 1092 720
rect 200 711 202 719
rect 488 711 490 719
rect 518 718 524 719
rect 111 710 115 711
rect 111 705 115 706
rect 199 710 203 711
rect 199 705 203 706
rect 255 710 259 711
rect 255 705 259 706
rect 487 710 491 711
rect 487 705 491 706
rect 112 694 114 705
rect 254 704 260 705
rect 254 700 255 704
rect 259 700 260 704
rect 254 699 260 700
rect 438 703 444 704
rect 438 699 439 703
rect 443 699 444 703
rect 438 698 444 699
rect 110 693 116 694
rect 110 689 111 693
rect 115 689 116 693
rect 110 688 116 689
rect 110 675 116 676
rect 110 671 111 675
rect 115 671 116 675
rect 110 670 116 671
rect 112 643 114 670
rect 440 668 442 698
rect 438 667 444 668
rect 438 663 439 667
rect 443 663 444 667
rect 438 662 444 663
rect 520 660 522 718
rect 784 711 786 719
rect 798 718 804 719
rect 1088 711 1090 719
rect 527 710 531 711
rect 527 705 531 706
rect 783 710 787 711
rect 783 705 787 706
rect 815 710 819 711
rect 815 705 819 706
rect 1087 710 1091 711
rect 1087 705 1091 706
rect 1111 710 1115 711
rect 1111 705 1115 706
rect 526 704 532 705
rect 814 704 820 705
rect 1110 704 1116 705
rect 526 700 527 704
rect 531 700 532 704
rect 526 699 532 700
rect 798 703 804 704
rect 798 699 799 703
rect 803 699 804 703
rect 814 700 815 704
rect 819 700 820 704
rect 814 699 820 700
rect 1098 703 1104 704
rect 1098 699 1099 703
rect 1103 699 1104 703
rect 1110 700 1111 704
rect 1115 700 1116 704
rect 1110 699 1116 700
rect 1142 703 1148 704
rect 1142 699 1143 703
rect 1147 699 1148 703
rect 798 698 804 699
rect 1098 698 1104 699
rect 1142 698 1148 699
rect 800 668 802 698
rect 1100 668 1102 698
rect 798 667 804 668
rect 798 663 799 667
rect 803 663 804 667
rect 798 662 804 663
rect 1098 667 1104 668
rect 1098 663 1099 667
rect 1103 663 1104 667
rect 1098 662 1104 663
rect 518 659 524 660
rect 254 658 260 659
rect 254 654 255 658
rect 259 654 260 658
rect 518 655 519 659
rect 523 655 524 659
rect 518 654 524 655
rect 526 658 532 659
rect 526 654 527 658
rect 531 654 532 658
rect 254 653 260 654
rect 526 653 532 654
rect 814 658 820 659
rect 814 654 815 658
rect 819 654 820 658
rect 814 653 820 654
rect 1110 658 1116 659
rect 1110 654 1111 658
rect 1115 654 1116 658
rect 1110 653 1116 654
rect 256 643 258 653
rect 528 643 530 653
rect 816 643 818 653
rect 1112 643 1114 653
rect 111 642 115 643
rect 111 637 115 638
rect 255 642 259 643
rect 255 637 259 638
rect 527 642 531 643
rect 527 637 531 638
rect 551 642 555 643
rect 551 637 555 638
rect 759 642 763 643
rect 759 637 763 638
rect 815 642 819 643
rect 815 637 819 638
rect 975 642 979 643
rect 1111 642 1115 643
rect 975 637 979 638
rect 1006 639 1012 640
rect 112 614 114 637
rect 552 631 554 637
rect 760 631 762 637
rect 976 631 978 637
rect 1006 635 1007 639
rect 1011 635 1012 639
rect 1111 637 1115 638
rect 1006 634 1012 635
rect 550 630 556 631
rect 550 626 551 630
rect 555 626 556 630
rect 550 625 556 626
rect 758 630 764 631
rect 758 626 759 630
rect 763 626 764 630
rect 758 625 764 626
rect 974 630 980 631
rect 974 626 975 630
rect 979 626 980 630
rect 974 625 980 626
rect 774 619 780 620
rect 774 615 775 619
rect 779 615 780 619
rect 774 614 780 615
rect 110 613 116 614
rect 110 609 111 613
rect 115 609 116 613
rect 110 608 116 609
rect 110 595 116 596
rect 110 591 111 595
rect 115 591 116 595
rect 110 590 116 591
rect 112 571 114 590
rect 550 584 556 585
rect 758 584 764 585
rect 776 584 778 614
rect 974 584 980 585
rect 1008 584 1010 634
rect 1144 632 1146 698
rect 1191 642 1195 643
rect 1191 637 1195 638
rect 1142 631 1148 632
rect 1192 631 1194 637
rect 1142 627 1143 631
rect 1147 627 1148 631
rect 1142 626 1148 627
rect 1190 630 1196 631
rect 1190 626 1191 630
rect 1195 626 1196 630
rect 1190 625 1196 626
rect 1190 584 1196 585
rect 1224 584 1226 762
rect 1568 754 1570 777
rect 1566 753 1572 754
rect 1566 749 1567 753
rect 1571 749 1572 753
rect 1566 748 1572 749
rect 1566 735 1572 736
rect 1566 731 1567 735
rect 1571 731 1572 735
rect 1566 730 1572 731
rect 1398 724 1404 725
rect 1398 720 1399 724
rect 1403 720 1404 724
rect 1398 719 1404 720
rect 1466 723 1472 724
rect 1466 719 1467 723
rect 1471 719 1472 723
rect 1400 711 1402 719
rect 1466 718 1472 719
rect 1399 710 1403 711
rect 1399 705 1403 706
rect 1407 710 1411 711
rect 1407 705 1411 706
rect 1406 704 1412 705
rect 1406 700 1407 704
rect 1411 700 1412 704
rect 1406 699 1412 700
rect 1468 660 1470 718
rect 1568 711 1570 730
rect 1567 710 1571 711
rect 1567 705 1571 706
rect 1474 703 1480 704
rect 1474 699 1475 703
rect 1479 699 1480 703
rect 1474 698 1480 699
rect 1466 659 1472 660
rect 1406 658 1412 659
rect 1406 654 1407 658
rect 1411 654 1412 658
rect 1466 655 1467 659
rect 1471 655 1472 659
rect 1466 654 1472 655
rect 1406 653 1412 654
rect 1408 643 1410 653
rect 1407 642 1411 643
rect 1407 637 1411 638
rect 1415 642 1419 643
rect 1415 637 1419 638
rect 1416 631 1418 637
rect 1476 632 1478 698
rect 1568 694 1570 705
rect 1566 693 1572 694
rect 1566 689 1567 693
rect 1571 689 1572 693
rect 1566 688 1572 689
rect 1566 675 1572 676
rect 1566 671 1567 675
rect 1571 671 1572 675
rect 1566 670 1572 671
rect 1568 643 1570 670
rect 1567 642 1571 643
rect 1567 637 1571 638
rect 1474 631 1480 632
rect 1414 630 1420 631
rect 1286 627 1292 628
rect 1286 623 1287 627
rect 1291 623 1292 627
rect 1414 626 1415 630
rect 1419 626 1420 630
rect 1474 627 1475 631
rect 1479 627 1480 631
rect 1474 626 1480 627
rect 1414 625 1420 626
rect 1286 622 1292 623
rect 550 580 551 584
rect 555 580 556 584
rect 550 579 556 580
rect 750 583 756 584
rect 750 579 751 583
rect 755 579 756 583
rect 758 580 759 584
rect 763 580 764 584
rect 758 579 764 580
rect 774 583 780 584
rect 774 579 775 583
rect 779 579 780 583
rect 974 580 975 584
rect 979 580 980 584
rect 974 579 980 580
rect 1006 583 1012 584
rect 1006 579 1007 583
rect 1011 579 1012 583
rect 1190 580 1191 584
rect 1195 580 1196 584
rect 1190 579 1196 580
rect 1222 583 1228 584
rect 1222 579 1223 583
rect 1227 579 1228 583
rect 552 571 554 579
rect 750 578 756 579
rect 111 570 115 571
rect 111 565 115 566
rect 551 570 555 571
rect 551 565 555 566
rect 727 570 731 571
rect 727 565 731 566
rect 112 554 114 565
rect 726 564 732 565
rect 726 560 727 564
rect 731 560 732 564
rect 726 559 732 560
rect 110 553 116 554
rect 110 549 111 553
rect 115 549 116 553
rect 110 548 116 549
rect 110 535 116 536
rect 110 531 111 535
rect 115 531 116 535
rect 110 530 116 531
rect 112 495 114 530
rect 752 520 754 578
rect 760 571 762 579
rect 774 578 780 579
rect 976 571 978 579
rect 1006 578 1012 579
rect 1192 571 1194 579
rect 1222 578 1228 579
rect 759 570 763 571
rect 759 565 763 566
rect 847 570 851 571
rect 847 565 851 566
rect 975 570 979 571
rect 975 565 979 566
rect 1111 570 1115 571
rect 1111 565 1115 566
rect 1191 570 1195 571
rect 1191 565 1195 566
rect 1255 570 1259 571
rect 1255 565 1259 566
rect 846 564 852 565
rect 974 564 980 565
rect 1110 564 1116 565
rect 834 563 840 564
rect 834 559 835 563
rect 839 559 840 563
rect 846 560 847 564
rect 851 560 852 564
rect 846 559 852 560
rect 914 563 920 564
rect 914 559 915 563
rect 919 559 920 563
rect 974 560 975 564
rect 979 560 980 564
rect 974 559 980 560
rect 1090 563 1096 564
rect 1090 559 1091 563
rect 1095 559 1096 563
rect 1110 560 1111 564
rect 1115 560 1116 564
rect 1110 559 1116 560
rect 1254 564 1260 565
rect 1288 564 1290 622
rect 1568 614 1570 637
rect 1566 613 1572 614
rect 1566 609 1567 613
rect 1571 609 1572 613
rect 1566 608 1572 609
rect 1566 595 1572 596
rect 1566 591 1567 595
rect 1571 591 1572 595
rect 1566 590 1572 591
rect 1414 584 1420 585
rect 1414 580 1415 584
rect 1419 580 1420 584
rect 1414 579 1420 580
rect 1470 583 1476 584
rect 1470 579 1471 583
rect 1475 579 1476 583
rect 1416 571 1418 579
rect 1470 578 1476 579
rect 1407 570 1411 571
rect 1407 565 1411 566
rect 1415 570 1419 571
rect 1415 565 1419 566
rect 1406 564 1412 565
rect 1254 560 1255 564
rect 1259 560 1260 564
rect 1254 559 1260 560
rect 1286 563 1292 564
rect 1286 559 1287 563
rect 1291 559 1292 563
rect 1406 560 1407 564
rect 1411 560 1412 564
rect 1406 559 1412 560
rect 834 558 840 559
rect 914 558 920 559
rect 1090 558 1096 559
rect 1286 558 1292 559
rect 836 528 838 558
rect 834 527 840 528
rect 834 523 835 527
rect 839 523 840 527
rect 834 522 840 523
rect 750 519 756 520
rect 726 518 732 519
rect 726 514 727 518
rect 731 514 732 518
rect 750 515 751 519
rect 755 515 756 519
rect 750 514 756 515
rect 846 518 852 519
rect 846 514 847 518
rect 851 514 852 518
rect 726 513 732 514
rect 846 513 852 514
rect 728 495 730 513
rect 848 495 850 513
rect 916 512 918 558
rect 1092 528 1094 558
rect 1090 527 1096 528
rect 1090 523 1091 527
rect 1095 523 1096 527
rect 1090 522 1096 523
rect 1472 520 1474 578
rect 1568 571 1570 590
rect 1567 570 1571 571
rect 1567 565 1571 566
rect 1494 563 1500 564
rect 1494 559 1495 563
rect 1499 559 1500 563
rect 1494 558 1500 559
rect 1470 519 1476 520
rect 974 518 980 519
rect 974 514 975 518
rect 979 514 980 518
rect 974 513 980 514
rect 1110 518 1116 519
rect 1110 514 1111 518
rect 1115 514 1116 518
rect 1110 513 1116 514
rect 1254 518 1260 519
rect 1254 514 1255 518
rect 1259 514 1260 518
rect 1254 513 1260 514
rect 1406 518 1412 519
rect 1406 514 1407 518
rect 1411 514 1412 518
rect 1470 515 1471 519
rect 1475 515 1476 519
rect 1470 514 1476 515
rect 1406 513 1412 514
rect 914 511 920 512
rect 914 507 915 511
rect 919 507 920 511
rect 914 506 920 507
rect 976 495 978 513
rect 1112 495 1114 513
rect 1186 511 1192 512
rect 1186 507 1187 511
rect 1191 507 1192 511
rect 1186 506 1192 507
rect 111 494 115 495
rect 111 489 115 490
rect 727 494 731 495
rect 727 489 731 490
rect 767 494 771 495
rect 767 489 771 490
rect 847 494 851 495
rect 847 489 851 490
rect 855 494 859 495
rect 855 489 859 490
rect 943 494 947 495
rect 943 489 947 490
rect 975 494 979 495
rect 975 489 979 490
rect 1031 494 1035 495
rect 1031 489 1035 490
rect 1111 494 1115 495
rect 1111 489 1115 490
rect 1119 494 1123 495
rect 1119 489 1123 490
rect 112 466 114 489
rect 768 483 770 489
rect 856 483 858 489
rect 944 483 946 489
rect 1032 483 1034 489
rect 1120 483 1122 489
rect 766 482 772 483
rect 766 478 767 482
rect 771 478 772 482
rect 766 477 772 478
rect 854 482 860 483
rect 854 478 855 482
rect 859 478 860 482
rect 854 477 860 478
rect 942 482 948 483
rect 942 478 943 482
rect 947 478 948 482
rect 942 477 948 478
rect 1030 482 1036 483
rect 1030 478 1031 482
rect 1035 478 1036 482
rect 1030 477 1036 478
rect 1118 482 1124 483
rect 1118 478 1119 482
rect 1123 478 1124 482
rect 1118 477 1124 478
rect 870 471 876 472
rect 870 467 871 471
rect 875 467 876 471
rect 870 466 876 467
rect 958 471 964 472
rect 958 467 959 471
rect 963 467 964 471
rect 958 466 964 467
rect 1046 471 1052 472
rect 1046 467 1047 471
rect 1051 467 1052 471
rect 1046 466 1052 467
rect 110 465 116 466
rect 110 461 111 465
rect 115 461 116 465
rect 110 460 116 461
rect 110 447 116 448
rect 110 443 111 447
rect 115 443 116 447
rect 110 442 116 443
rect 112 415 114 442
rect 766 436 772 437
rect 766 432 767 436
rect 771 432 772 436
rect 766 431 772 432
rect 854 436 860 437
rect 872 436 874 466
rect 934 451 940 452
rect 934 447 935 451
rect 939 447 940 451
rect 934 446 940 447
rect 854 432 855 436
rect 859 432 860 436
rect 854 431 860 432
rect 870 435 876 436
rect 870 431 871 435
rect 875 431 876 435
rect 768 415 770 431
rect 856 415 858 431
rect 870 430 876 431
rect 111 414 115 415
rect 111 409 115 410
rect 623 414 627 415
rect 623 409 627 410
rect 711 414 715 415
rect 711 409 715 410
rect 767 414 771 415
rect 767 409 771 410
rect 799 414 803 415
rect 799 409 803 410
rect 855 414 859 415
rect 855 409 859 410
rect 887 414 891 415
rect 887 409 891 410
rect 112 398 114 409
rect 622 408 628 409
rect 710 408 716 409
rect 622 404 623 408
rect 627 404 628 408
rect 622 403 628 404
rect 698 407 704 408
rect 698 403 699 407
rect 703 403 704 407
rect 710 404 711 408
rect 715 404 716 408
rect 710 403 716 404
rect 798 408 804 409
rect 798 404 799 408
rect 803 404 804 408
rect 798 403 804 404
rect 886 408 892 409
rect 886 404 887 408
rect 891 404 892 408
rect 886 403 892 404
rect 918 407 924 408
rect 918 403 919 407
rect 923 403 924 407
rect 698 402 704 403
rect 918 402 924 403
rect 110 397 116 398
rect 110 393 111 397
rect 115 393 116 397
rect 110 392 116 393
rect 690 391 696 392
rect 690 387 691 391
rect 695 387 696 391
rect 690 386 696 387
rect 110 379 116 380
rect 110 375 111 379
rect 115 375 116 379
rect 110 374 116 375
rect 112 335 114 374
rect 692 364 694 386
rect 690 363 696 364
rect 622 362 628 363
rect 622 358 623 362
rect 627 358 628 362
rect 690 359 691 363
rect 695 359 696 363
rect 690 358 696 359
rect 622 357 628 358
rect 624 335 626 357
rect 111 334 115 335
rect 111 329 115 330
rect 399 334 403 335
rect 399 329 403 330
rect 487 334 491 335
rect 487 329 491 330
rect 575 334 579 335
rect 575 329 579 330
rect 623 334 627 335
rect 623 329 627 330
rect 663 334 667 335
rect 663 329 667 330
rect 112 306 114 329
rect 400 323 402 329
rect 488 323 490 329
rect 576 323 578 329
rect 664 323 666 329
rect 700 324 702 402
rect 778 391 784 392
rect 778 387 779 391
rect 783 387 784 391
rect 778 386 784 387
rect 780 364 782 386
rect 778 363 784 364
rect 710 362 716 363
rect 710 358 711 362
rect 715 358 716 362
rect 778 359 779 363
rect 783 359 784 363
rect 778 358 784 359
rect 798 362 804 363
rect 798 358 799 362
rect 803 358 804 362
rect 710 357 716 358
rect 798 357 804 358
rect 886 362 892 363
rect 886 358 887 362
rect 891 358 892 362
rect 886 357 892 358
rect 712 335 714 357
rect 800 335 802 357
rect 888 335 890 357
rect 920 356 922 402
rect 936 364 938 446
rect 942 436 948 437
rect 960 436 962 466
rect 1030 436 1036 437
rect 1048 436 1050 466
rect 1188 440 1190 506
rect 1256 495 1258 513
rect 1408 495 1410 513
rect 1207 494 1211 495
rect 1207 489 1211 490
rect 1255 494 1259 495
rect 1255 489 1259 490
rect 1295 494 1299 495
rect 1295 489 1299 490
rect 1383 494 1387 495
rect 1383 489 1387 490
rect 1407 494 1411 495
rect 1407 489 1411 490
rect 1471 494 1475 495
rect 1471 489 1475 490
rect 1208 483 1210 489
rect 1296 483 1298 489
rect 1384 483 1386 489
rect 1472 483 1474 489
rect 1496 484 1498 558
rect 1568 554 1570 565
rect 1566 553 1572 554
rect 1566 549 1567 553
rect 1571 549 1572 553
rect 1566 548 1572 549
rect 1566 535 1572 536
rect 1566 531 1567 535
rect 1571 531 1572 535
rect 1566 530 1572 531
rect 1568 495 1570 530
rect 1567 494 1571 495
rect 1567 489 1571 490
rect 1494 483 1500 484
rect 1206 482 1212 483
rect 1206 478 1207 482
rect 1211 478 1212 482
rect 1206 477 1212 478
rect 1294 482 1300 483
rect 1294 478 1295 482
rect 1299 478 1300 482
rect 1294 477 1300 478
rect 1382 482 1388 483
rect 1382 478 1383 482
rect 1387 478 1388 482
rect 1382 477 1388 478
rect 1470 482 1476 483
rect 1470 478 1471 482
rect 1475 478 1476 482
rect 1494 479 1495 483
rect 1499 479 1500 483
rect 1494 478 1500 479
rect 1470 477 1476 478
rect 1222 471 1228 472
rect 1222 467 1223 471
rect 1227 467 1228 471
rect 1222 466 1228 467
rect 1310 471 1316 472
rect 1310 467 1311 471
rect 1315 467 1316 471
rect 1310 466 1316 467
rect 1398 471 1404 472
rect 1398 467 1399 471
rect 1403 467 1404 471
rect 1398 466 1404 467
rect 1486 471 1492 472
rect 1486 467 1487 471
rect 1491 467 1492 471
rect 1486 466 1492 467
rect 1568 466 1570 489
rect 1186 439 1192 440
rect 1118 436 1124 437
rect 942 432 943 436
rect 947 432 948 436
rect 942 431 948 432
rect 958 435 964 436
rect 958 431 959 435
rect 963 431 964 435
rect 1030 432 1031 436
rect 1035 432 1036 436
rect 1030 431 1036 432
rect 1046 435 1052 436
rect 1046 431 1047 435
rect 1051 431 1052 435
rect 1118 432 1119 436
rect 1123 432 1124 436
rect 1186 435 1187 439
rect 1191 435 1192 439
rect 1186 434 1192 435
rect 1206 436 1212 437
rect 1224 436 1226 466
rect 1294 436 1300 437
rect 1312 436 1314 466
rect 1382 436 1388 437
rect 1400 436 1402 466
rect 1470 436 1476 437
rect 1488 436 1490 466
rect 1566 465 1572 466
rect 1566 461 1567 465
rect 1571 461 1572 465
rect 1566 460 1572 461
rect 1566 447 1572 448
rect 1566 443 1567 447
rect 1571 443 1572 447
rect 1566 442 1572 443
rect 1118 431 1124 432
rect 1206 432 1207 436
rect 1211 432 1212 436
rect 1206 431 1212 432
rect 1222 435 1228 436
rect 1222 431 1223 435
rect 1227 431 1228 435
rect 1294 432 1295 436
rect 1299 432 1300 436
rect 1294 431 1300 432
rect 1310 435 1316 436
rect 1310 431 1311 435
rect 1315 431 1316 435
rect 1382 432 1383 436
rect 1387 432 1388 436
rect 1382 431 1388 432
rect 1398 435 1404 436
rect 1398 431 1399 435
rect 1403 431 1404 435
rect 1470 432 1471 436
rect 1475 432 1476 436
rect 1470 431 1476 432
rect 1486 435 1492 436
rect 1486 431 1487 435
rect 1491 431 1492 435
rect 944 415 946 431
rect 958 430 964 431
rect 1032 415 1034 431
rect 1046 430 1052 431
rect 1120 415 1122 431
rect 1208 415 1210 431
rect 1222 430 1228 431
rect 1296 415 1298 431
rect 1310 430 1316 431
rect 1384 415 1386 431
rect 1398 430 1404 431
rect 1472 415 1474 431
rect 1486 430 1492 431
rect 1568 415 1570 442
rect 943 414 947 415
rect 943 409 947 410
rect 1031 414 1035 415
rect 1031 409 1035 410
rect 1119 414 1123 415
rect 1119 409 1123 410
rect 1207 414 1211 415
rect 1207 409 1211 410
rect 1295 414 1299 415
rect 1295 409 1299 410
rect 1383 414 1387 415
rect 1383 409 1387 410
rect 1471 414 1475 415
rect 1471 409 1475 410
rect 1567 414 1571 415
rect 1567 409 1571 410
rect 1568 398 1570 409
rect 1566 397 1572 398
rect 1566 393 1567 397
rect 1571 393 1572 397
rect 1566 392 1572 393
rect 1566 379 1572 380
rect 1566 375 1567 379
rect 1571 375 1572 379
rect 1566 374 1572 375
rect 934 363 940 364
rect 934 359 935 363
rect 939 359 940 363
rect 934 358 940 359
rect 918 355 924 356
rect 918 351 919 355
rect 923 351 924 355
rect 918 350 924 351
rect 1568 335 1570 374
rect 711 334 715 335
rect 711 329 715 330
rect 799 334 803 335
rect 799 329 803 330
rect 887 334 891 335
rect 887 329 891 330
rect 1567 334 1571 335
rect 1567 329 1571 330
rect 698 323 704 324
rect 398 322 404 323
rect 398 318 399 322
rect 403 318 404 322
rect 398 317 404 318
rect 486 322 492 323
rect 486 318 487 322
rect 491 318 492 322
rect 486 317 492 318
rect 574 322 580 323
rect 574 318 575 322
rect 579 318 580 322
rect 574 317 580 318
rect 662 322 668 323
rect 662 318 663 322
rect 667 318 668 322
rect 698 319 699 323
rect 703 319 704 323
rect 698 318 704 319
rect 662 317 668 318
rect 502 311 508 312
rect 502 307 503 311
rect 507 307 508 311
rect 502 306 508 307
rect 590 311 596 312
rect 590 307 591 311
rect 595 307 596 311
rect 590 306 596 307
rect 678 311 684 312
rect 678 307 679 311
rect 683 307 684 311
rect 678 306 684 307
rect 1568 306 1570 329
rect 110 305 116 306
rect 110 301 111 305
rect 115 301 116 305
rect 110 300 116 301
rect 110 287 116 288
rect 110 283 111 287
rect 115 283 116 287
rect 110 282 116 283
rect 112 251 114 282
rect 398 276 404 277
rect 486 276 492 277
rect 504 276 506 306
rect 574 276 580 277
rect 592 276 594 306
rect 662 276 668 277
rect 680 276 682 306
rect 1566 305 1572 306
rect 1566 301 1567 305
rect 1571 301 1572 305
rect 1566 300 1572 301
rect 1566 287 1572 288
rect 1566 283 1567 287
rect 1571 283 1572 287
rect 1566 282 1572 283
rect 398 272 399 276
rect 403 272 404 276
rect 398 271 404 272
rect 466 275 472 276
rect 466 271 467 275
rect 471 271 472 275
rect 486 272 487 276
rect 491 272 492 276
rect 486 271 492 272
rect 502 275 508 276
rect 502 271 503 275
rect 507 271 508 275
rect 574 272 575 276
rect 579 272 580 276
rect 574 271 580 272
rect 590 275 596 276
rect 590 271 591 275
rect 595 271 596 275
rect 662 272 663 276
rect 667 272 668 276
rect 662 271 668 272
rect 678 275 684 276
rect 678 271 679 275
rect 683 271 684 275
rect 400 251 402 271
rect 466 270 472 271
rect 111 250 115 251
rect 111 245 115 246
rect 215 250 219 251
rect 215 245 219 246
rect 303 250 307 251
rect 303 245 307 246
rect 391 250 395 251
rect 391 245 395 246
rect 399 250 403 251
rect 399 245 403 246
rect 112 234 114 245
rect 214 244 220 245
rect 302 244 308 245
rect 214 240 215 244
rect 219 240 220 244
rect 214 239 220 240
rect 274 243 280 244
rect 274 239 275 243
rect 279 239 280 243
rect 302 240 303 244
rect 307 240 308 244
rect 302 239 308 240
rect 390 244 396 245
rect 390 240 391 244
rect 395 240 396 244
rect 390 239 396 240
rect 274 238 280 239
rect 110 233 116 234
rect 110 229 111 233
rect 115 229 116 233
rect 110 228 116 229
rect 276 221 278 238
rect 282 227 288 228
rect 282 223 283 227
rect 287 223 288 227
rect 282 222 288 223
rect 370 227 376 228
rect 370 223 371 227
rect 375 223 376 227
rect 370 222 376 223
rect 458 227 464 228
rect 458 223 459 227
rect 463 223 464 227
rect 458 222 464 223
rect 275 220 279 221
rect 110 215 116 216
rect 275 215 279 216
rect 110 211 111 215
rect 115 211 116 215
rect 110 210 116 211
rect 112 155 114 210
rect 284 200 286 222
rect 372 200 374 222
rect 460 200 462 222
rect 468 208 470 270
rect 488 251 490 271
rect 502 270 508 271
rect 576 251 578 271
rect 590 270 596 271
rect 664 251 666 271
rect 678 270 684 271
rect 1568 251 1570 282
rect 479 250 483 251
rect 479 245 483 246
rect 487 250 491 251
rect 487 245 491 246
rect 575 250 579 251
rect 575 245 579 246
rect 663 250 667 251
rect 663 245 667 246
rect 1567 250 1571 251
rect 1567 245 1571 246
rect 478 244 484 245
rect 478 240 479 244
rect 483 240 484 244
rect 478 239 484 240
rect 1568 234 1570 245
rect 1566 233 1572 234
rect 1566 229 1567 233
rect 1571 229 1572 233
rect 1566 228 1572 229
rect 599 220 603 221
rect 599 215 603 216
rect 1566 215 1572 216
rect 466 207 472 208
rect 466 203 467 207
rect 471 203 472 207
rect 466 202 472 203
rect 282 199 288 200
rect 370 199 376 200
rect 458 199 464 200
rect 214 198 220 199
rect 214 194 215 198
rect 219 194 220 198
rect 282 195 283 199
rect 287 195 288 199
rect 282 194 288 195
rect 302 198 308 199
rect 302 194 303 198
rect 307 194 308 198
rect 370 195 371 199
rect 375 195 376 199
rect 370 194 376 195
rect 390 198 396 199
rect 390 194 391 198
rect 395 194 396 198
rect 458 195 459 199
rect 463 195 464 199
rect 458 194 464 195
rect 478 198 484 199
rect 478 194 479 198
rect 483 194 484 198
rect 214 193 220 194
rect 302 193 308 194
rect 390 193 396 194
rect 478 193 484 194
rect 216 155 218 193
rect 304 155 306 193
rect 392 155 394 193
rect 480 155 482 193
rect 111 154 115 155
rect 111 149 115 150
rect 135 154 139 155
rect 135 149 139 150
rect 215 154 219 155
rect 215 149 219 150
rect 223 154 227 155
rect 223 149 227 150
rect 303 154 307 155
rect 303 149 307 150
rect 311 154 315 155
rect 311 149 315 150
rect 391 154 395 155
rect 391 149 395 150
rect 399 154 403 155
rect 399 149 403 150
rect 479 154 483 155
rect 479 149 483 150
rect 487 154 491 155
rect 487 149 491 150
rect 575 154 579 155
rect 575 149 579 150
rect 112 126 114 149
rect 136 143 138 149
rect 224 143 226 149
rect 312 143 314 149
rect 400 143 402 149
rect 488 143 490 149
rect 576 143 578 149
rect 600 144 602 215
rect 1566 211 1567 215
rect 1571 211 1572 215
rect 1566 210 1572 211
rect 1568 155 1570 210
rect 1567 154 1571 155
rect 1567 149 1571 150
rect 598 143 604 144
rect 134 142 140 143
rect 134 138 135 142
rect 139 138 140 142
rect 134 137 140 138
rect 222 142 228 143
rect 222 138 223 142
rect 227 138 228 142
rect 222 137 228 138
rect 310 142 316 143
rect 310 138 311 142
rect 315 138 316 142
rect 310 137 316 138
rect 398 142 404 143
rect 398 138 399 142
rect 403 138 404 142
rect 398 137 404 138
rect 486 142 492 143
rect 486 138 487 142
rect 491 138 492 142
rect 486 137 492 138
rect 574 142 580 143
rect 574 138 575 142
rect 579 138 580 142
rect 598 139 599 143
rect 603 139 604 143
rect 598 138 604 139
rect 574 137 580 138
rect 238 131 244 132
rect 238 127 239 131
rect 243 127 244 131
rect 238 126 244 127
rect 326 131 332 132
rect 326 127 327 131
rect 331 127 332 131
rect 326 126 332 127
rect 414 131 420 132
rect 414 127 415 131
rect 419 127 420 131
rect 414 126 420 127
rect 502 131 508 132
rect 502 127 503 131
rect 507 127 508 131
rect 502 126 508 127
rect 590 131 596 132
rect 590 127 591 131
rect 595 127 596 131
rect 590 126 596 127
rect 1568 126 1570 149
rect 110 125 116 126
rect 110 121 111 125
rect 115 121 116 125
rect 110 120 116 121
rect 110 107 116 108
rect 110 103 111 107
rect 115 103 116 107
rect 110 102 116 103
rect 112 91 114 102
rect 134 96 140 97
rect 134 92 135 96
rect 139 92 140 96
rect 134 91 140 92
rect 222 96 228 97
rect 240 96 242 126
rect 310 96 316 97
rect 328 96 330 126
rect 398 96 404 97
rect 416 96 418 126
rect 486 96 492 97
rect 504 96 506 126
rect 574 96 580 97
rect 592 96 594 126
rect 1566 125 1572 126
rect 1566 121 1567 125
rect 1571 121 1572 125
rect 1566 120 1572 121
rect 1566 107 1572 108
rect 1566 103 1567 107
rect 1571 103 1572 107
rect 1566 102 1572 103
rect 222 92 223 96
rect 227 92 228 96
rect 222 91 228 92
rect 238 95 244 96
rect 238 91 239 95
rect 243 91 244 95
rect 310 92 311 96
rect 315 92 316 96
rect 310 91 316 92
rect 326 95 332 96
rect 326 91 327 95
rect 331 91 332 95
rect 398 92 399 96
rect 403 92 404 96
rect 398 91 404 92
rect 414 95 420 96
rect 414 91 415 95
rect 419 91 420 95
rect 486 92 487 96
rect 491 92 492 96
rect 486 91 492 92
rect 502 95 508 96
rect 502 91 503 95
rect 507 91 508 95
rect 574 92 575 96
rect 579 92 580 96
rect 574 91 580 92
rect 590 95 596 96
rect 590 91 591 95
rect 595 91 596 95
rect 1568 91 1570 102
rect 111 90 115 91
rect 111 85 115 86
rect 135 90 139 91
rect 135 85 139 86
rect 223 90 227 91
rect 238 90 244 91
rect 311 90 315 91
rect 326 90 332 91
rect 399 90 403 91
rect 414 90 420 91
rect 487 90 491 91
rect 502 90 508 91
rect 575 90 579 91
rect 590 90 596 91
rect 1567 90 1571 91
rect 223 85 227 86
rect 311 85 315 86
rect 399 85 403 86
rect 487 85 491 86
rect 575 85 579 86
rect 1567 85 1571 86
<< m4c >>
rect 111 1526 115 1530
rect 543 1526 547 1530
rect 631 1526 635 1530
rect 719 1526 723 1530
rect 807 1526 811 1530
rect 895 1526 899 1530
rect 1567 1526 1571 1530
rect 111 1462 115 1466
rect 471 1462 475 1466
rect 543 1462 547 1466
rect 615 1462 619 1466
rect 111 1394 115 1398
rect 423 1394 427 1398
rect 471 1394 475 1398
rect 631 1462 635 1466
rect 719 1462 723 1466
rect 775 1462 779 1466
rect 807 1462 811 1466
rect 895 1462 899 1466
rect 943 1462 947 1466
rect 1119 1462 1123 1466
rect 1303 1462 1307 1466
rect 1471 1462 1475 1466
rect 1567 1462 1571 1466
rect 615 1394 619 1398
rect 663 1394 667 1398
rect 775 1394 779 1398
rect 911 1394 915 1398
rect 943 1394 947 1398
rect 1119 1394 1123 1398
rect 1167 1394 1171 1398
rect 1303 1394 1307 1398
rect 1431 1394 1435 1398
rect 1471 1394 1475 1398
rect 1567 1394 1571 1398
rect 111 1318 115 1322
rect 423 1318 427 1322
rect 487 1318 491 1322
rect 663 1318 667 1322
rect 727 1318 731 1322
rect 111 1242 115 1246
rect 487 1242 491 1246
rect 535 1242 539 1246
rect 911 1318 915 1322
rect 967 1318 971 1322
rect 1167 1318 1171 1322
rect 1215 1318 1219 1322
rect 1431 1318 1435 1322
rect 1463 1318 1467 1322
rect 727 1242 731 1246
rect 743 1242 747 1246
rect 959 1242 963 1246
rect 967 1242 971 1246
rect 1175 1242 1179 1246
rect 1215 1242 1219 1246
rect 1399 1242 1403 1246
rect 1567 1318 1571 1322
rect 1463 1242 1467 1246
rect 1567 1242 1571 1246
rect 111 1162 115 1166
rect 535 1162 539 1166
rect 655 1162 659 1166
rect 743 1162 747 1166
rect 831 1162 835 1166
rect 959 1162 963 1166
rect 1015 1162 1019 1166
rect 111 1086 115 1090
rect 655 1086 659 1090
rect 663 1086 667 1090
rect 1175 1162 1179 1166
rect 1207 1162 1211 1166
rect 1399 1162 1403 1166
rect 1567 1162 1571 1166
rect 831 1086 835 1090
rect 847 1086 851 1090
rect 1015 1086 1019 1090
rect 1031 1086 1035 1090
rect 1207 1086 1211 1090
rect 1223 1086 1227 1090
rect 1399 1086 1403 1090
rect 1423 1086 1427 1090
rect 1567 1086 1571 1090
rect 111 1006 115 1010
rect 551 1006 555 1010
rect 663 1006 667 1010
rect 759 1006 763 1010
rect 847 1006 851 1010
rect 975 1006 979 1010
rect 1031 1006 1035 1010
rect 111 930 115 934
rect 399 930 403 934
rect 551 930 555 934
rect 1199 1006 1203 1010
rect 1223 1006 1227 1010
rect 1423 1006 1427 1010
rect 1431 1006 1435 1010
rect 1567 1006 1571 1010
rect 663 930 667 934
rect 759 930 763 934
rect 927 930 931 934
rect 975 930 979 934
rect 1199 930 1203 934
rect 111 854 115 858
rect 255 854 259 858
rect 399 854 403 858
rect 535 854 539 858
rect 663 854 667 858
rect 823 854 827 858
rect 927 854 931 858
rect 111 778 115 782
rect 199 778 203 782
rect 255 778 259 782
rect 1111 854 1115 858
rect 1199 854 1203 858
rect 1431 930 1435 934
rect 1471 930 1475 934
rect 1567 930 1571 934
rect 1407 854 1411 858
rect 1471 854 1475 858
rect 1567 854 1571 858
rect 487 778 491 782
rect 535 778 539 782
rect 783 778 787 782
rect 823 778 827 782
rect 1087 778 1091 782
rect 1111 778 1115 782
rect 1399 778 1403 782
rect 1407 778 1411 782
rect 1567 778 1571 782
rect 111 706 115 710
rect 199 706 203 710
rect 255 706 259 710
rect 487 706 491 710
rect 527 706 531 710
rect 783 706 787 710
rect 815 706 819 710
rect 1087 706 1091 710
rect 1111 706 1115 710
rect 111 638 115 642
rect 255 638 259 642
rect 527 638 531 642
rect 551 638 555 642
rect 759 638 763 642
rect 815 638 819 642
rect 975 638 979 642
rect 1111 638 1115 642
rect 1191 638 1195 642
rect 1399 706 1403 710
rect 1407 706 1411 710
rect 1567 706 1571 710
rect 1407 638 1411 642
rect 1415 638 1419 642
rect 1567 638 1571 642
rect 111 566 115 570
rect 551 566 555 570
rect 727 566 731 570
rect 759 566 763 570
rect 847 566 851 570
rect 975 566 979 570
rect 1111 566 1115 570
rect 1191 566 1195 570
rect 1255 566 1259 570
rect 1407 566 1411 570
rect 1415 566 1419 570
rect 1567 566 1571 570
rect 111 490 115 494
rect 727 490 731 494
rect 767 490 771 494
rect 847 490 851 494
rect 855 490 859 494
rect 943 490 947 494
rect 975 490 979 494
rect 1031 490 1035 494
rect 1111 490 1115 494
rect 1119 490 1123 494
rect 111 410 115 414
rect 623 410 627 414
rect 711 410 715 414
rect 767 410 771 414
rect 799 410 803 414
rect 855 410 859 414
rect 887 410 891 414
rect 111 330 115 334
rect 399 330 403 334
rect 487 330 491 334
rect 575 330 579 334
rect 623 330 627 334
rect 663 330 667 334
rect 1207 490 1211 494
rect 1255 490 1259 494
rect 1295 490 1299 494
rect 1383 490 1387 494
rect 1407 490 1411 494
rect 1471 490 1475 494
rect 1567 490 1571 494
rect 943 410 947 414
rect 1031 410 1035 414
rect 1119 410 1123 414
rect 1207 410 1211 414
rect 1295 410 1299 414
rect 1383 410 1387 414
rect 1471 410 1475 414
rect 1567 410 1571 414
rect 711 330 715 334
rect 799 330 803 334
rect 887 330 891 334
rect 1567 330 1571 334
rect 111 246 115 250
rect 215 246 219 250
rect 303 246 307 250
rect 391 246 395 250
rect 399 246 403 250
rect 275 216 279 220
rect 479 246 483 250
rect 487 246 491 250
rect 575 246 579 250
rect 663 246 667 250
rect 1567 246 1571 250
rect 599 216 603 220
rect 111 150 115 154
rect 135 150 139 154
rect 215 150 219 154
rect 223 150 227 154
rect 303 150 307 154
rect 311 150 315 154
rect 391 150 395 154
rect 399 150 403 154
rect 479 150 483 154
rect 487 150 491 154
rect 575 150 579 154
rect 1567 150 1571 154
rect 111 86 115 90
rect 135 86 139 90
rect 223 86 227 90
rect 311 86 315 90
rect 399 86 403 90
rect 487 86 491 90
rect 575 86 579 90
rect 1567 86 1571 90
<< m4 >>
rect 96 1525 97 1531
rect 103 1530 1603 1531
rect 103 1526 111 1530
rect 115 1526 543 1530
rect 547 1526 631 1530
rect 635 1526 719 1530
rect 723 1526 807 1530
rect 811 1526 895 1530
rect 899 1526 1567 1530
rect 1571 1526 1603 1530
rect 103 1525 1603 1526
rect 1609 1525 1610 1531
rect 84 1461 85 1467
rect 91 1466 1591 1467
rect 91 1462 111 1466
rect 115 1462 471 1466
rect 475 1462 543 1466
rect 547 1462 615 1466
rect 619 1462 631 1466
rect 635 1462 719 1466
rect 723 1462 775 1466
rect 779 1462 807 1466
rect 811 1462 895 1466
rect 899 1462 943 1466
rect 947 1462 1119 1466
rect 1123 1462 1303 1466
rect 1307 1462 1471 1466
rect 1475 1462 1567 1466
rect 1571 1462 1591 1466
rect 91 1461 1591 1462
rect 1597 1461 1598 1467
rect 96 1393 97 1399
rect 103 1398 1603 1399
rect 103 1394 111 1398
rect 115 1394 423 1398
rect 427 1394 471 1398
rect 475 1394 615 1398
rect 619 1394 663 1398
rect 667 1394 775 1398
rect 779 1394 911 1398
rect 915 1394 943 1398
rect 947 1394 1119 1398
rect 1123 1394 1167 1398
rect 1171 1394 1303 1398
rect 1307 1394 1431 1398
rect 1435 1394 1471 1398
rect 1475 1394 1567 1398
rect 1571 1394 1603 1398
rect 103 1393 1603 1394
rect 1609 1393 1610 1399
rect 84 1317 85 1323
rect 91 1322 1591 1323
rect 91 1318 111 1322
rect 115 1318 423 1322
rect 427 1318 487 1322
rect 491 1318 663 1322
rect 667 1318 727 1322
rect 731 1318 911 1322
rect 915 1318 967 1322
rect 971 1318 1167 1322
rect 1171 1318 1215 1322
rect 1219 1318 1431 1322
rect 1435 1318 1463 1322
rect 1467 1318 1567 1322
rect 1571 1318 1591 1322
rect 91 1317 1591 1318
rect 1597 1317 1598 1323
rect 96 1241 97 1247
rect 103 1246 1603 1247
rect 103 1242 111 1246
rect 115 1242 487 1246
rect 491 1242 535 1246
rect 539 1242 727 1246
rect 731 1242 743 1246
rect 747 1242 959 1246
rect 963 1242 967 1246
rect 971 1242 1175 1246
rect 1179 1242 1215 1246
rect 1219 1242 1399 1246
rect 1403 1242 1463 1246
rect 1467 1242 1567 1246
rect 1571 1242 1603 1246
rect 103 1241 1603 1242
rect 1609 1241 1610 1247
rect 84 1161 85 1167
rect 91 1166 1591 1167
rect 91 1162 111 1166
rect 115 1162 535 1166
rect 539 1162 655 1166
rect 659 1162 743 1166
rect 747 1162 831 1166
rect 835 1162 959 1166
rect 963 1162 1015 1166
rect 1019 1162 1175 1166
rect 1179 1162 1207 1166
rect 1211 1162 1399 1166
rect 1403 1162 1567 1166
rect 1571 1162 1591 1166
rect 91 1161 1591 1162
rect 1597 1161 1598 1167
rect 96 1085 97 1091
rect 103 1090 1603 1091
rect 103 1086 111 1090
rect 115 1086 655 1090
rect 659 1086 663 1090
rect 667 1086 831 1090
rect 835 1086 847 1090
rect 851 1086 1015 1090
rect 1019 1086 1031 1090
rect 1035 1086 1207 1090
rect 1211 1086 1223 1090
rect 1227 1086 1399 1090
rect 1403 1086 1423 1090
rect 1427 1086 1567 1090
rect 1571 1086 1603 1090
rect 103 1085 1603 1086
rect 1609 1085 1610 1091
rect 84 1005 85 1011
rect 91 1010 1591 1011
rect 91 1006 111 1010
rect 115 1006 551 1010
rect 555 1006 663 1010
rect 667 1006 759 1010
rect 763 1006 847 1010
rect 851 1006 975 1010
rect 979 1006 1031 1010
rect 1035 1006 1199 1010
rect 1203 1006 1223 1010
rect 1227 1006 1423 1010
rect 1427 1006 1431 1010
rect 1435 1006 1567 1010
rect 1571 1006 1591 1010
rect 91 1005 1591 1006
rect 1597 1005 1598 1011
rect 96 929 97 935
rect 103 934 1603 935
rect 103 930 111 934
rect 115 930 399 934
rect 403 930 551 934
rect 555 930 663 934
rect 667 930 759 934
rect 763 930 927 934
rect 931 930 975 934
rect 979 930 1199 934
rect 1203 930 1431 934
rect 1435 930 1471 934
rect 1475 930 1567 934
rect 1571 930 1603 934
rect 103 929 1603 930
rect 1609 929 1610 935
rect 84 853 85 859
rect 91 858 1591 859
rect 91 854 111 858
rect 115 854 255 858
rect 259 854 399 858
rect 403 854 535 858
rect 539 854 663 858
rect 667 854 823 858
rect 827 854 927 858
rect 931 854 1111 858
rect 1115 854 1199 858
rect 1203 854 1407 858
rect 1411 854 1471 858
rect 1475 854 1567 858
rect 1571 854 1591 858
rect 91 853 1591 854
rect 1597 853 1598 859
rect 96 777 97 783
rect 103 782 1603 783
rect 103 778 111 782
rect 115 778 199 782
rect 203 778 255 782
rect 259 778 487 782
rect 491 778 535 782
rect 539 778 783 782
rect 787 778 823 782
rect 827 778 1087 782
rect 1091 778 1111 782
rect 1115 778 1399 782
rect 1403 778 1407 782
rect 1411 778 1567 782
rect 1571 778 1603 782
rect 103 777 1603 778
rect 1609 777 1610 783
rect 84 705 85 711
rect 91 710 1591 711
rect 91 706 111 710
rect 115 706 199 710
rect 203 706 255 710
rect 259 706 487 710
rect 491 706 527 710
rect 531 706 783 710
rect 787 706 815 710
rect 819 706 1087 710
rect 1091 706 1111 710
rect 1115 706 1399 710
rect 1403 706 1407 710
rect 1411 706 1567 710
rect 1571 706 1591 710
rect 91 705 1591 706
rect 1597 705 1598 711
rect 96 637 97 643
rect 103 642 1603 643
rect 103 638 111 642
rect 115 638 255 642
rect 259 638 527 642
rect 531 638 551 642
rect 555 638 759 642
rect 763 638 815 642
rect 819 638 975 642
rect 979 638 1111 642
rect 1115 638 1191 642
rect 1195 638 1407 642
rect 1411 638 1415 642
rect 1419 638 1567 642
rect 1571 638 1603 642
rect 103 637 1603 638
rect 1609 637 1610 643
rect 84 565 85 571
rect 91 570 1591 571
rect 91 566 111 570
rect 115 566 551 570
rect 555 566 727 570
rect 731 566 759 570
rect 763 566 847 570
rect 851 566 975 570
rect 979 566 1111 570
rect 1115 566 1191 570
rect 1195 566 1255 570
rect 1259 566 1407 570
rect 1411 566 1415 570
rect 1419 566 1567 570
rect 1571 566 1591 570
rect 91 565 1591 566
rect 1597 565 1598 571
rect 96 489 97 495
rect 103 494 1603 495
rect 103 490 111 494
rect 115 490 727 494
rect 731 490 767 494
rect 771 490 847 494
rect 851 490 855 494
rect 859 490 943 494
rect 947 490 975 494
rect 979 490 1031 494
rect 1035 490 1111 494
rect 1115 490 1119 494
rect 1123 490 1207 494
rect 1211 490 1255 494
rect 1259 490 1295 494
rect 1299 490 1383 494
rect 1387 490 1407 494
rect 1411 490 1471 494
rect 1475 490 1567 494
rect 1571 490 1603 494
rect 103 489 1603 490
rect 1609 489 1610 495
rect 84 409 85 415
rect 91 414 1591 415
rect 91 410 111 414
rect 115 410 623 414
rect 627 410 711 414
rect 715 410 767 414
rect 771 410 799 414
rect 803 410 855 414
rect 859 410 887 414
rect 891 410 943 414
rect 947 410 1031 414
rect 1035 410 1119 414
rect 1123 410 1207 414
rect 1211 410 1295 414
rect 1299 410 1383 414
rect 1387 410 1471 414
rect 1475 410 1567 414
rect 1571 410 1591 414
rect 91 409 1591 410
rect 1597 409 1598 415
rect 96 329 97 335
rect 103 334 1603 335
rect 103 330 111 334
rect 115 330 399 334
rect 403 330 487 334
rect 491 330 575 334
rect 579 330 623 334
rect 627 330 663 334
rect 667 330 711 334
rect 715 330 799 334
rect 803 330 887 334
rect 891 330 1567 334
rect 1571 330 1603 334
rect 103 329 1603 330
rect 1609 329 1610 335
rect 84 245 85 251
rect 91 250 1591 251
rect 91 246 111 250
rect 115 246 215 250
rect 219 246 303 250
rect 307 246 391 250
rect 395 246 399 250
rect 403 246 479 250
rect 483 246 487 250
rect 491 246 575 250
rect 579 246 663 250
rect 667 246 1567 250
rect 1571 246 1591 250
rect 91 245 1591 246
rect 1597 245 1598 251
rect 274 220 280 221
rect 598 220 604 221
rect 274 216 275 220
rect 279 216 599 220
rect 603 216 604 220
rect 274 215 280 216
rect 598 215 604 216
rect 96 149 97 155
rect 103 154 1603 155
rect 103 150 111 154
rect 115 150 135 154
rect 139 150 215 154
rect 219 150 223 154
rect 227 150 303 154
rect 307 150 311 154
rect 315 150 391 154
rect 395 150 399 154
rect 403 150 479 154
rect 483 150 487 154
rect 491 150 575 154
rect 579 150 1567 154
rect 1571 150 1603 154
rect 103 149 1603 150
rect 1609 149 1610 155
rect 84 85 85 91
rect 91 90 1591 91
rect 91 86 111 90
rect 115 86 135 90
rect 139 86 223 90
rect 227 86 311 90
rect 315 86 399 90
rect 403 86 487 90
rect 491 86 575 90
rect 579 86 1567 90
rect 1571 86 1591 90
rect 91 85 1591 86
rect 1597 85 1598 91
<< m5c >>
rect 97 1525 103 1531
rect 1603 1525 1609 1531
rect 85 1461 91 1467
rect 1591 1461 1597 1467
rect 97 1393 103 1399
rect 1603 1393 1609 1399
rect 85 1317 91 1323
rect 1591 1317 1597 1323
rect 97 1241 103 1247
rect 1603 1241 1609 1247
rect 85 1161 91 1167
rect 1591 1161 1597 1167
rect 97 1085 103 1091
rect 1603 1085 1609 1091
rect 85 1005 91 1011
rect 1591 1005 1597 1011
rect 97 929 103 935
rect 1603 929 1609 935
rect 85 853 91 859
rect 1591 853 1597 859
rect 97 777 103 783
rect 1603 777 1609 783
rect 85 705 91 711
rect 1591 705 1597 711
rect 97 637 103 643
rect 1603 637 1609 643
rect 85 565 91 571
rect 1591 565 1597 571
rect 97 489 103 495
rect 1603 489 1609 495
rect 85 409 91 415
rect 1591 409 1597 415
rect 97 329 103 335
rect 1603 329 1609 335
rect 85 245 91 251
rect 1591 245 1597 251
rect 97 149 103 155
rect 1603 149 1609 155
rect 85 85 91 91
rect 1591 85 1597 91
<< m5 >>
rect 84 1467 92 1656
rect 84 1461 85 1467
rect 91 1461 92 1467
rect 84 1323 92 1461
rect 84 1317 85 1323
rect 91 1317 92 1323
rect 84 1167 92 1317
rect 84 1161 85 1167
rect 91 1161 92 1167
rect 84 1011 92 1161
rect 84 1005 85 1011
rect 91 1005 92 1011
rect 84 859 92 1005
rect 84 853 85 859
rect 91 853 92 859
rect 84 711 92 853
rect 84 705 85 711
rect 91 705 92 711
rect 84 571 92 705
rect 84 565 85 571
rect 91 565 92 571
rect 84 415 92 565
rect 84 409 85 415
rect 91 409 92 415
rect 84 251 92 409
rect 84 245 85 251
rect 91 245 92 251
rect 84 91 92 245
rect 84 85 85 91
rect 91 85 92 91
rect 84 72 92 85
rect 96 1531 104 1656
rect 96 1525 97 1531
rect 103 1525 104 1531
rect 96 1399 104 1525
rect 96 1393 97 1399
rect 103 1393 104 1399
rect 96 1247 104 1393
rect 96 1241 97 1247
rect 103 1241 104 1247
rect 96 1091 104 1241
rect 96 1085 97 1091
rect 103 1085 104 1091
rect 96 935 104 1085
rect 96 929 97 935
rect 103 929 104 935
rect 96 783 104 929
rect 96 777 97 783
rect 103 777 104 783
rect 96 643 104 777
rect 96 637 97 643
rect 103 637 104 643
rect 96 495 104 637
rect 96 489 97 495
rect 103 489 104 495
rect 96 335 104 489
rect 96 329 97 335
rect 103 329 104 335
rect 96 155 104 329
rect 96 149 97 155
rect 103 149 104 155
rect 96 72 104 149
rect 1590 1467 1598 1656
rect 1590 1461 1591 1467
rect 1597 1461 1598 1467
rect 1590 1323 1598 1461
rect 1590 1317 1591 1323
rect 1597 1317 1598 1323
rect 1590 1167 1598 1317
rect 1590 1161 1591 1167
rect 1597 1161 1598 1167
rect 1590 1011 1598 1161
rect 1590 1005 1591 1011
rect 1597 1005 1598 1011
rect 1590 859 1598 1005
rect 1590 853 1591 859
rect 1597 853 1598 859
rect 1590 711 1598 853
rect 1590 705 1591 711
rect 1597 705 1598 711
rect 1590 571 1598 705
rect 1590 565 1591 571
rect 1597 565 1598 571
rect 1590 415 1598 565
rect 1590 409 1591 415
rect 1597 409 1598 415
rect 1590 251 1598 409
rect 1590 245 1591 251
rect 1597 245 1598 251
rect 1590 91 1598 245
rect 1590 85 1591 91
rect 1597 85 1598 91
rect 1590 72 1598 85
rect 1602 1531 1610 1656
rect 1602 1525 1603 1531
rect 1609 1525 1610 1531
rect 1602 1399 1610 1525
rect 1602 1393 1603 1399
rect 1609 1393 1610 1399
rect 1602 1247 1610 1393
rect 1602 1241 1603 1247
rect 1609 1241 1610 1247
rect 1602 1091 1610 1241
rect 1602 1085 1603 1091
rect 1609 1085 1610 1091
rect 1602 935 1610 1085
rect 1602 929 1603 935
rect 1609 929 1610 935
rect 1602 783 1610 929
rect 1602 777 1603 783
rect 1609 777 1610 783
rect 1602 643 1610 777
rect 1602 637 1603 643
rect 1609 637 1610 643
rect 1602 495 1610 637
rect 1602 489 1603 495
rect 1609 489 1610 495
rect 1602 335 1610 489
rect 1602 329 1603 335
rect 1609 329 1610 335
rect 1602 155 1610 329
rect 1602 149 1603 155
rect 1609 149 1610 155
rect 1602 72 1610 149
use _0_0cell_0_0gcelem3x0  celem_599_6_acx0
timestamp 1730767052
transform 1 0 128 0 1 88
box 8 4 79 60
use welltap_svt  __well_tap__0
timestamp 1730767052
transform 1 0 104 0 1 100
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0cell_0_0gcelem3x0  celem_599_6_acx0
timestamp 1730767052
transform 1 0 128 0 1 88
box 8 4 79 60
use welltap_svt  __well_tap__0
timestamp 1730767052
transform 1 0 104 0 1 100
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0cell_0_0gcelem3x0  celem_598_6_acx0
timestamp 1730767052
transform 1 0 216 0 1 88
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_598_6_acx0
timestamp 1730767052
transform 1 0 216 0 1 88
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_597_6_acx0
timestamp 1730767052
transform 1 0 304 0 1 88
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_597_6_acx0
timestamp 1730767052
transform 1 0 304 0 1 88
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_596_6_acx0
timestamp 1730767052
transform 1 0 392 0 1 88
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_596_6_acx0
timestamp 1730767052
transform 1 0 392 0 1 88
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_595_6_acx0
timestamp 1730767052
transform 1 0 480 0 1 88
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_595_6_acx0
timestamp 1730767052
transform 1 0 480 0 1 88
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_594_6_acx0
timestamp 1730767052
transform 1 0 568 0 1 88
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_594_6_acx0
timestamp 1730767052
transform 1 0 568 0 1 88
box 8 4 79 60
use welltap_svt  __well_tap__1
timestamp 1730767052
transform 1 0 1560 0 1 100
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1730767052
transform 1 0 1560 0 1 100
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730767052
transform 1 0 104 0 -1 236
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730767052
transform 1 0 104 0 -1 236
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_593_6_acx0
timestamp 1730767052
transform 1 0 208 0 -1 248
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_593_6_acx0
timestamp 1730767052
transform 1 0 208 0 -1 248
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_592_6_acx0
timestamp 1730767052
transform 1 0 296 0 -1 248
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_592_6_acx0
timestamp 1730767052
transform 1 0 296 0 -1 248
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_591_6_acx0
timestamp 1730767052
transform 1 0 384 0 -1 248
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_591_6_acx0
timestamp 1730767052
transform 1 0 384 0 -1 248
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_590_6_acx0
timestamp 1730767052
transform 1 0 472 0 -1 248
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_590_6_acx0
timestamp 1730767052
transform 1 0 472 0 -1 248
box 8 4 79 60
use welltap_svt  __well_tap__3
timestamp 1730767052
transform 1 0 1560 0 -1 236
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730767052
transform 1 0 1560 0 -1 236
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730767052
transform 1 0 104 0 1 280
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730767052
transform 1 0 104 0 1 280
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_589_6_acx0
timestamp 1730767052
transform 1 0 392 0 1 268
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_589_6_acx0
timestamp 1730767052
transform 1 0 392 0 1 268
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_588_6_acx0
timestamp 1730767052
transform 1 0 480 0 1 268
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_588_6_acx0
timestamp 1730767052
transform 1 0 480 0 1 268
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_587_6_acx0
timestamp 1730767052
transform 1 0 568 0 1 268
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_587_6_acx0
timestamp 1730767052
transform 1 0 568 0 1 268
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_586_6_acx0
timestamp 1730767052
transform 1 0 656 0 1 268
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_586_6_acx0
timestamp 1730767052
transform 1 0 656 0 1 268
box 8 4 79 60
use welltap_svt  __well_tap__5
timestamp 1730767052
transform 1 0 1560 0 1 280
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730767052
transform 1 0 1560 0 1 280
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730767052
transform 1 0 104 0 -1 400
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730767052
transform 1 0 104 0 -1 400
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_585_6_acx0
timestamp 1730767052
transform 1 0 616 0 -1 412
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_585_6_acx0
timestamp 1730767052
transform 1 0 616 0 -1 412
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_584_6_acx0
timestamp 1730767052
transform 1 0 704 0 -1 412
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_584_6_acx0
timestamp 1730767052
transform 1 0 704 0 -1 412
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_583_6_acx0
timestamp 1730767052
transform 1 0 792 0 -1 412
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_583_6_acx0
timestamp 1730767052
transform 1 0 792 0 -1 412
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_582_6_acx0
timestamp 1730767052
transform 1 0 880 0 -1 412
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_582_6_acx0
timestamp 1730767052
transform 1 0 880 0 -1 412
box 8 4 79 60
use welltap_svt  __well_tap__7
timestamp 1730767052
transform 1 0 1560 0 -1 400
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1730767052
transform 1 0 1560 0 -1 400
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730767052
transform 1 0 104 0 1 440
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730767052
transform 1 0 104 0 1 440
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_581_6_acx0
timestamp 1730767052
transform 1 0 760 0 1 428
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_581_6_acx0
timestamp 1730767052
transform 1 0 760 0 1 428
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_580_6_acx0
timestamp 1730767052
transform 1 0 848 0 1 428
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_580_6_acx0
timestamp 1730767052
transform 1 0 848 0 1 428
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_579_6_acx0
timestamp 1730767052
transform 1 0 936 0 1 428
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_579_6_acx0
timestamp 1730767052
transform 1 0 936 0 1 428
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_578_6_acx0
timestamp 1730767052
transform 1 0 1024 0 1 428
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_578_6_acx0
timestamp 1730767052
transform 1 0 1024 0 1 428
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_520_6_acx0
timestamp 1730767052
transform 1 0 1112 0 1 428
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_520_6_acx0
timestamp 1730767052
transform 1 0 1112 0 1 428
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_519_6_acx0
timestamp 1730767052
transform 1 0 1200 0 1 428
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_519_6_acx0
timestamp 1730767052
transform 1 0 1200 0 1 428
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_518_6_acx0
timestamp 1730767052
transform 1 0 1288 0 1 428
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_518_6_acx0
timestamp 1730767052
transform 1 0 1288 0 1 428
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_517_6_acx0
timestamp 1730767052
transform 1 0 1376 0 1 428
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_517_6_acx0
timestamp 1730767052
transform 1 0 1376 0 1 428
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_516_6_acx0
timestamp 1730767052
transform 1 0 1464 0 1 428
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_516_6_acx0
timestamp 1730767052
transform 1 0 1464 0 1 428
box 8 4 79 60
use welltap_svt  __well_tap__9
timestamp 1730767052
transform 1 0 1560 0 1 440
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730767052
transform 1 0 1560 0 1 440
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730767052
transform 1 0 104 0 -1 556
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730767052
transform 1 0 104 0 1 588
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730767052
transform 1 0 104 0 -1 556
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730767052
transform 1 0 104 0 1 588
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_573_6_acx0
timestamp 1730767052
transform 1 0 544 0 1 576
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_573_6_acx0
timestamp 1730767052
transform 1 0 544 0 1 576
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_572_6_acx0
timestamp 1730767052
transform 1 0 752 0 1 576
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_574_6_acx0
timestamp 1730767052
transform 1 0 720 0 -1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_572_6_acx0
timestamp 1730767052
transform 1 0 752 0 1 576
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_574_6_acx0
timestamp 1730767052
transform 1 0 720 0 -1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_575_6_acx0
timestamp 1730767052
transform 1 0 840 0 -1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_575_6_acx0
timestamp 1730767052
transform 1 0 840 0 -1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_571_6_acx0
timestamp 1730767052
transform 1 0 968 0 1 576
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_576_6_acx0
timestamp 1730767052
transform 1 0 968 0 -1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_571_6_acx0
timestamp 1730767052
transform 1 0 968 0 1 576
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_576_6_acx0
timestamp 1730767052
transform 1 0 968 0 -1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_577_6_acx0
timestamp 1730767052
transform 1 0 1104 0 -1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_577_6_acx0
timestamp 1730767052
transform 1 0 1104 0 -1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_522_6_acx0
timestamp 1730767052
transform 1 0 1184 0 1 576
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_522_6_acx0
timestamp 1730767052
transform 1 0 1184 0 1 576
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_521_6_acx0
timestamp 1730767052
transform 1 0 1248 0 -1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_521_6_acx0
timestamp 1730767052
transform 1 0 1248 0 -1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_514_6_acx0
timestamp 1730767052
transform 1 0 1408 0 1 576
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_515_6_acx0
timestamp 1730767052
transform 1 0 1400 0 -1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_514_6_acx0
timestamp 1730767052
transform 1 0 1408 0 1 576
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_515_6_acx0
timestamp 1730767052
transform 1 0 1400 0 -1 568
box 8 4 79 60
use welltap_svt  __well_tap__11
timestamp 1730767052
transform 1 0 1560 0 -1 556
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730767052
transform 1 0 1560 0 1 588
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730767052
transform 1 0 1560 0 -1 556
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730767052
transform 1 0 1560 0 1 588
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730767052
transform 1 0 104 0 -1 696
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730767052
transform 1 0 104 0 -1 696
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_567_6_acx0
timestamp 1730767052
transform 1 0 248 0 -1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_567_6_acx0
timestamp 1730767052
transform 1 0 248 0 -1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_568_6_acx0
timestamp 1730767052
transform 1 0 520 0 -1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_568_6_acx0
timestamp 1730767052
transform 1 0 520 0 -1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_569_6_acx0
timestamp 1730767052
transform 1 0 808 0 -1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_569_6_acx0
timestamp 1730767052
transform 1 0 808 0 -1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_570_6_acx0
timestamp 1730767052
transform 1 0 1104 0 -1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_570_6_acx0
timestamp 1730767052
transform 1 0 1104 0 -1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_513_6_acx0
timestamp 1730767052
transform 1 0 1400 0 -1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_513_6_acx0
timestamp 1730767052
transform 1 0 1400 0 -1 708
box 8 4 79 60
use welltap_svt  __well_tap__15
timestamp 1730767052
transform 1 0 1560 0 -1 696
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1730767052
transform 1 0 1560 0 -1 696
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730767052
transform 1 0 104 0 1 728
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730767052
transform 1 0 104 0 1 728
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_564_6_acx0
timestamp 1730767052
transform 1 0 192 0 1 716
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_564_6_acx0
timestamp 1730767052
transform 1 0 192 0 1 716
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_566_6_acx0
timestamp 1730767052
transform 1 0 480 0 1 716
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_566_6_acx0
timestamp 1730767052
transform 1 0 480 0 1 716
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_565_6_acx0
timestamp 1730767052
transform 1 0 776 0 1 716
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_565_6_acx0
timestamp 1730767052
transform 1 0 776 0 1 716
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_523_6_acx0
timestamp 1730767052
transform 1 0 1080 0 1 716
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_523_6_acx0
timestamp 1730767052
transform 1 0 1080 0 1 716
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_512_6_acx0
timestamp 1730767052
transform 1 0 1392 0 1 716
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_512_6_acx0
timestamp 1730767052
transform 1 0 1392 0 1 716
box 8 4 79 60
use welltap_svt  __well_tap__17
timestamp 1730767052
transform 1 0 1560 0 1 728
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730767052
transform 1 0 1560 0 1 728
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730767052
transform 1 0 104 0 -1 844
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730767052
transform 1 0 104 0 -1 844
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_563_6_acx0
timestamp 1730767052
transform 1 0 248 0 -1 856
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_563_6_acx0
timestamp 1730767052
transform 1 0 248 0 -1 856
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_562_6_acx0
timestamp 1730767052
transform 1 0 528 0 -1 856
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_562_6_acx0
timestamp 1730767052
transform 1 0 528 0 -1 856
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_561_6_acx0
timestamp 1730767052
transform 1 0 816 0 -1 856
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_561_6_acx0
timestamp 1730767052
transform 1 0 816 0 -1 856
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_524_6_acx0
timestamp 1730767052
transform 1 0 1104 0 -1 856
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_524_6_acx0
timestamp 1730767052
transform 1 0 1104 0 -1 856
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_511_6_acx0
timestamp 1730767052
transform 1 0 1400 0 -1 856
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_511_6_acx0
timestamp 1730767052
transform 1 0 1400 0 -1 856
box 8 4 79 60
use welltap_svt  __well_tap__19
timestamp 1730767052
transform 1 0 1560 0 -1 844
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730767052
transform 1 0 1560 0 -1 844
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730767052
transform 1 0 104 0 1 880
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730767052
transform 1 0 104 0 1 880
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_558_6_acx0
timestamp 1730767052
transform 1 0 392 0 1 868
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_558_6_acx0
timestamp 1730767052
transform 1 0 392 0 1 868
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_559_6_acx0
timestamp 1730767052
transform 1 0 656 0 1 868
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_559_6_acx0
timestamp 1730767052
transform 1 0 656 0 1 868
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_560_6_acx0
timestamp 1730767052
transform 1 0 920 0 1 868
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_560_6_acx0
timestamp 1730767052
transform 1 0 920 0 1 868
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_510_6_acx0
timestamp 1730767052
transform 1 0 1192 0 1 868
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_510_6_acx0
timestamp 1730767052
transform 1 0 1192 0 1 868
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_59_6_acx0
timestamp 1730767052
transform 1 0 1464 0 1 868
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_59_6_acx0
timestamp 1730767052
transform 1 0 1464 0 1 868
box 8 4 79 60
use welltap_svt  __well_tap__21
timestamp 1730767052
transform 1 0 1560 0 1 880
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730767052
transform 1 0 1560 0 1 880
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730767052
transform 1 0 104 0 -1 996
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730767052
transform 1 0 104 0 -1 996
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_557_6_acx0
timestamp 1730767052
transform 1 0 544 0 -1 1008
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_557_6_acx0
timestamp 1730767052
transform 1 0 544 0 -1 1008
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_552_6_acx0
timestamp 1730767052
transform 1 0 656 0 1 1024
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_552_6_acx0
timestamp 1730767052
transform 1 0 656 0 1 1024
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_556_6_acx0
timestamp 1730767052
transform 1 0 752 0 -1 1008
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_556_6_acx0
timestamp 1730767052
transform 1 0 752 0 -1 1008
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_553_6_acx0
timestamp 1730767052
transform 1 0 840 0 1 1024
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_553_6_acx0
timestamp 1730767052
transform 1 0 840 0 1 1024
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_554_6_acx0
timestamp 1730767052
transform 1 0 1024 0 1 1024
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_555_6_acx0
timestamp 1730767052
transform 1 0 968 0 -1 1008
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_554_6_acx0
timestamp 1730767052
transform 1 0 1024 0 1 1024
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_555_6_acx0
timestamp 1730767052
transform 1 0 968 0 -1 1008
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_525_6_acx0
timestamp 1730767052
transform 1 0 1192 0 -1 1008
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_525_6_acx0
timestamp 1730767052
transform 1 0 1192 0 -1 1008
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_526_6_acx0
timestamp 1730767052
transform 1 0 1216 0 1 1024
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_526_6_acx0
timestamp 1730767052
transform 1 0 1216 0 1 1024
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_57_6_acx0
timestamp 1730767052
transform 1 0 1416 0 1 1024
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_58_6_acx0
timestamp 1730767052
transform 1 0 1424 0 -1 1008
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_57_6_acx0
timestamp 1730767052
transform 1 0 1416 0 1 1024
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_58_6_acx0
timestamp 1730767052
transform 1 0 1424 0 -1 1008
box 8 4 79 60
use welltap_svt  __well_tap__23
timestamp 1730767052
transform 1 0 1560 0 -1 996
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1730767052
transform 1 0 1560 0 -1 996
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730767052
transform 1 0 104 0 1 1036
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730767052
transform 1 0 104 0 1 1036
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_551_6_acx0
timestamp 1730767052
transform 1 0 648 0 -1 1164
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_551_6_acx0
timestamp 1730767052
transform 1 0 648 0 -1 1164
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_550_6_acx0
timestamp 1730767052
transform 1 0 824 0 -1 1164
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_550_6_acx0
timestamp 1730767052
transform 1 0 824 0 -1 1164
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_549_6_acx0
timestamp 1730767052
transform 1 0 1008 0 -1 1164
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_549_6_acx0
timestamp 1730767052
transform 1 0 1008 0 -1 1164
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_527_6_acx0
timestamp 1730767052
transform 1 0 1200 0 -1 1164
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_527_6_acx0
timestamp 1730767052
transform 1 0 1200 0 -1 1164
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_56_6_acx0
timestamp 1730767052
transform 1 0 1392 0 -1 1164
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_56_6_acx0
timestamp 1730767052
transform 1 0 1392 0 -1 1164
box 8 4 79 60
use welltap_svt  __well_tap__25
timestamp 1730767052
transform 1 0 1560 0 1 1036
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1730767052
transform 1 0 1560 0 1 1036
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730767052
transform 1 0 104 0 -1 1152
box 8 4 12 24
use welltap_svt  __well_tap__28
timestamp 1730767052
transform 1 0 104 0 1 1192
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730767052
transform 1 0 104 0 -1 1152
box 8 4 12 24
use welltap_svt  __well_tap__28
timestamp 1730767052
transform 1 0 104 0 1 1192
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_546_6_acx0
timestamp 1730767052
transform 1 0 528 0 1 1180
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_546_6_acx0
timestamp 1730767052
transform 1 0 528 0 1 1180
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_547_6_acx0
timestamp 1730767052
transform 1 0 736 0 1 1180
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_547_6_acx0
timestamp 1730767052
transform 1 0 736 0 1 1180
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_548_6_acx0
timestamp 1730767052
transform 1 0 952 0 1 1180
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_548_6_acx0
timestamp 1730767052
transform 1 0 952 0 1 1180
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_528_6_acx0
timestamp 1730767052
transform 1 0 1168 0 1 1180
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_528_6_acx0
timestamp 1730767052
transform 1 0 1168 0 1 1180
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_55_6_acx0
timestamp 1730767052
transform 1 0 1392 0 1 1180
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_55_6_acx0
timestamp 1730767052
transform 1 0 1392 0 1 1180
box 8 4 79 60
use welltap_svt  __well_tap__27
timestamp 1730767052
transform 1 0 1560 0 -1 1152
box 8 4 12 24
use welltap_svt  __well_tap__29
timestamp 1730767052
transform 1 0 1560 0 1 1192
box 8 4 12 24
use welltap_svt  __well_tap__27
timestamp 1730767052
transform 1 0 1560 0 -1 1152
box 8 4 12 24
use welltap_svt  __well_tap__29
timestamp 1730767052
transform 1 0 1560 0 1 1192
box 8 4 12 24
use welltap_svt  __well_tap__30
timestamp 1730767052
transform 1 0 104 0 -1 1308
box 8 4 12 24
use welltap_svt  __well_tap__30
timestamp 1730767052
transform 1 0 104 0 -1 1308
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_545_6_acx0
timestamp 1730767052
transform 1 0 480 0 -1 1320
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_545_6_acx0
timestamp 1730767052
transform 1 0 480 0 -1 1320
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_544_6_acx0
timestamp 1730767052
transform 1 0 720 0 -1 1320
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_544_6_acx0
timestamp 1730767052
transform 1 0 720 0 -1 1320
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_529_6_acx0
timestamp 1730767052
transform 1 0 960 0 -1 1320
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_529_6_acx0
timestamp 1730767052
transform 1 0 960 0 -1 1320
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_54_6_acx0
timestamp 1730767052
transform 1 0 1208 0 -1 1320
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_54_6_acx0
timestamp 1730767052
transform 1 0 1208 0 -1 1320
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_53_6_acx0
timestamp 1730767052
transform 1 0 1456 0 -1 1320
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_53_6_acx0
timestamp 1730767052
transform 1 0 1456 0 -1 1320
box 8 4 79 60
use welltap_svt  __well_tap__31
timestamp 1730767052
transform 1 0 1560 0 -1 1308
box 8 4 12 24
use welltap_svt  __well_tap__31
timestamp 1730767052
transform 1 0 1560 0 -1 1308
box 8 4 12 24
use welltap_svt  __well_tap__32
timestamp 1730767052
transform 1 0 104 0 1 1344
box 8 4 12 24
use welltap_svt  __well_tap__32
timestamp 1730767052
transform 1 0 104 0 1 1344
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_541_6_acx0
timestamp 1730767052
transform 1 0 416 0 1 1332
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_541_6_acx0
timestamp 1730767052
transform 1 0 416 0 1 1332
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_542_6_acx0
timestamp 1730767052
transform 1 0 656 0 1 1332
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_542_6_acx0
timestamp 1730767052
transform 1 0 656 0 1 1332
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_543_6_acx0
timestamp 1730767052
transform 1 0 904 0 1 1332
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_543_6_acx0
timestamp 1730767052
transform 1 0 904 0 1 1332
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_530_6_acx0
timestamp 1730767052
transform 1 0 1160 0 1 1332
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_530_6_acx0
timestamp 1730767052
transform 1 0 1160 0 1 1332
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_52_6_acx0
timestamp 1730767052
transform 1 0 1424 0 1 1332
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_52_6_acx0
timestamp 1730767052
transform 1 0 1424 0 1 1332
box 8 4 79 60
use welltap_svt  __well_tap__33
timestamp 1730767052
transform 1 0 1560 0 1 1344
box 8 4 12 24
use welltap_svt  __well_tap__33
timestamp 1730767052
transform 1 0 1560 0 1 1344
box 8 4 12 24
use welltap_svt  __well_tap__34
timestamp 1730767052
transform 1 0 104 0 -1 1452
box 8 4 12 24
use welltap_svt  __well_tap__34
timestamp 1730767052
transform 1 0 104 0 -1 1452
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_540_6_acx0
timestamp 1730767052
transform 1 0 464 0 -1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_540_6_acx0
timestamp 1730767052
transform 1 0 464 0 -1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_539_6_acx0
timestamp 1730767052
transform 1 0 608 0 -1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_539_6_acx0
timestamp 1730767052
transform 1 0 608 0 -1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_538_6_acx0
timestamp 1730767052
transform 1 0 768 0 -1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_538_6_acx0
timestamp 1730767052
transform 1 0 768 0 -1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_532_6_acx0
timestamp 1730767052
transform 1 0 936 0 -1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_532_6_acx0
timestamp 1730767052
transform 1 0 936 0 -1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_531_6_acx0
timestamp 1730767052
transform 1 0 1112 0 -1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_531_6_acx0
timestamp 1730767052
transform 1 0 1112 0 -1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_50_6_acx0
timestamp 1730767052
transform 1 0 1296 0 -1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_50_6_acx0
timestamp 1730767052
transform 1 0 1296 0 -1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_51_6_acx0
timestamp 1730767052
transform 1 0 1464 0 -1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_51_6_acx0
timestamp 1730767052
transform 1 0 1464 0 -1 1464
box 8 4 79 60
use welltap_svt  __well_tap__35
timestamp 1730767052
transform 1 0 1560 0 -1 1452
box 8 4 12 24
use welltap_svt  __well_tap__35
timestamp 1730767052
transform 1 0 1560 0 -1 1452
box 8 4 12 24
use welltap_svt  __well_tap__36
timestamp 1730767052
transform 1 0 104 0 1 1476
box 8 4 12 24
use welltap_svt  __well_tap__36
timestamp 1730767052
transform 1 0 104 0 1 1476
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_537_6_acx0
timestamp 1730767052
transform 1 0 536 0 1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_537_6_acx0
timestamp 1730767052
transform 1 0 536 0 1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_536_6_acx0
timestamp 1730767052
transform 1 0 624 0 1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_536_6_acx0
timestamp 1730767052
transform 1 0 624 0 1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_535_6_acx0
timestamp 1730767052
transform 1 0 712 0 1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_535_6_acx0
timestamp 1730767052
transform 1 0 712 0 1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_534_6_acx0
timestamp 1730767052
transform 1 0 800 0 1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_534_6_acx0
timestamp 1730767052
transform 1 0 800 0 1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_533_6_acx0
timestamp 1730767052
transform 1 0 888 0 1 1464
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_533_6_acx0
timestamp 1730767052
transform 1 0 888 0 1 1464
box 8 4 79 60
use welltap_svt  __well_tap__37
timestamp 1730767052
transform 1 0 1560 0 1 1476
box 8 4 12 24
use welltap_svt  __well_tap__37
timestamp 1730767052
transform 1 0 1560 0 1 1476
box 8 4 12 24
<< end >>
