magic
tech TSMC180
timestamp 1734143631
<< m1 >>
rect 6 57 9 60
rect 24 57 27 60
rect 42 57 45 60
rect 60 57 63 60
rect 6 18 59 51
rect 6 10 9 13
<< labels >>
rlabel m1 s 6 57 9 60 6 in_50_6
port 1 nsew signal input
rlabel m1 s 24 57 27 60 6 in_51_6
port 2 nsew signal input
rlabel m1 s 6 10 9 13 6 out
port 3 nsew signal output
rlabel m1 s 42 57 45 60 6 Vdd
port 4 nsew power input
rlabel m1 s 60 57 63 60 6 GND
port 5 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 66 70
string LEFclass CORE
string LEFsite CoreSite
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
