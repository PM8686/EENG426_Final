magic
tech sky130l
timestamp 1731220307
<< checkpaint >>
rect -19 61 52 69
rect -24 44 52 61
rect -24 -24 60 44
rect -24 -26 52 -24
rect -19 -28 47 -26
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 11 20 12
rect 15 8 16 11
rect 19 8 20 11
rect 15 6 20 8
<< ndc >>
rect 9 7 12 10
rect 16 8 19 11
<< ntransistor >>
rect 13 6 15 12
<< pdiffusion >>
rect 8 28 13 29
rect 8 25 9 28
rect 12 25 13 28
rect 8 19 13 25
rect 15 28 20 29
rect 15 25 16 28
rect 19 25 20 28
rect 15 19 20 25
<< pdc >>
rect 9 25 12 28
rect 16 25 19 28
<< ptransistor >>
rect 13 19 15 29
<< polysilicon >>
rect 13 36 20 37
rect 13 33 16 36
rect 19 33 20 36
rect 13 32 20 33
rect 13 29 15 32
rect 13 12 15 19
rect 13 4 15 6
<< pc >>
rect 16 33 19 36
<< m1 >>
rect 16 36 19 37
rect 9 28 12 29
rect 9 24 12 25
rect 16 28 19 33
rect 16 24 19 25
rect 24 11 28 12
rect 9 10 12 11
rect 15 8 16 11
rect 19 8 28 11
rect 9 6 12 7
<< m2c >>
rect 9 25 12 28
rect 9 7 12 10
<< m2 >>
rect 8 28 13 29
rect 8 25 9 28
rect 12 25 13 28
rect 8 24 13 25
rect 8 10 13 11
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
<< labels >>
rlabel space 0 0 32 40 6 prboundary
rlabel pdiffusion 20 26 20 26 3 x
rlabel polysilicon 20 34 20 34 3 x
rlabel ndiffusion 16 7 16 7 3 Y
rlabel ndiffusion 16 12 16 12 3 Y
rlabel pdiffusion 16 20 16 20 3 x
rlabel pdiffusion 16 26 16 26 3 x
rlabel pdiffusion 16 29 16 29 3 x
rlabel polysilicon 14 5 14 5 3 x
rlabel ntransistor 14 7 14 7 3 x
rlabel polysilicon 14 13 14 13 3 x
rlabel ptransistor 14 20 14 20 3 x
rlabel polysilicon 14 30 14 30 3 x
rlabel polysilicon 14 33 14 33 3 x
rlabel polysilicon 14 34 14 34 3 x
rlabel polysilicon 14 37 14 37 3 x
rlabel pdiffusion 9 20 9 20 3 Vdd
rlabel m1 25 12 25 12 3 Y
port 1 e
rlabel m1 20 9 20 9 3 Y
port 1 e
rlabel ndc 17 9 17 9 3 Y
port 1 e
rlabel m1 17 25 17 25 3 x
rlabel pdc 17 26 17 26 3 x
rlabel m1 17 29 17 29 3 x
rlabel pc 17 34 17 34 3 x
rlabel m1 17 37 17 37 3 x
rlabel m1 16 9 16 9 3 Y
port 1 e
rlabel m1 10 7 10 7 3 GND
rlabel m1 10 11 10 11 3 GND
rlabel m1 10 25 10 25 3 Vdd
rlabel m1 10 29 10 29 3 Vdd
rlabel m2 13 8 13 8 3 GND
rlabel m2 13 26 13 26 3 Vdd
rlabel m2c 10 8 10 8 3 GND
rlabel m2c 10 26 10 26 3 Vdd
rlabel m2 9 7 9 7 3 GND
rlabel m2 9 8 9 8 3 GND
rlabel m2 9 11 9 11 3 GND
rlabel m2 9 25 9 25 3 Vdd
rlabel m2 9 26 9 26 3 Vdd
rlabel m2 9 29 9 29 3 Vdd
<< end >>
