magic
tech sky130l
timestamp 1731220305
<< checkpaint >>
rect -16 81 52 84
rect -16 76 62 81
rect -16 43 84 76
rect -23 40 84 43
rect -24 8 84 40
rect -24 -9 81 8
rect -24 -14 74 -9
rect -24 -16 69 -14
rect -24 -20 68 -16
rect -24 -25 55 -20
rect -24 -28 44 -25
<< ndiffusion >>
rect 16 23 21 24
rect 16 20 17 23
rect 20 20 21 23
rect 16 14 21 20
rect 23 14 28 24
rect 30 22 35 24
rect 30 19 31 22
rect 34 19 35 22
rect 30 18 35 19
rect 37 23 42 24
rect 37 20 38 23
rect 41 20 42 23
rect 37 18 42 20
rect 30 14 34 18
<< ndc >>
rect 17 20 20 23
rect 31 19 34 22
rect 38 20 41 23
<< ntransistor >>
rect 21 14 23 24
rect 28 14 30 24
rect 35 18 37 24
<< pdiffusion >>
rect 16 38 21 39
rect 16 35 17 38
rect 20 35 21 38
rect 16 31 21 35
rect 23 35 28 39
rect 23 32 24 35
rect 27 32 28 35
rect 23 31 28 32
rect 30 38 35 39
rect 30 35 31 38
rect 34 35 35 38
rect 30 31 35 35
rect 37 38 42 39
rect 37 35 38 38
rect 41 35 42 38
rect 37 31 42 35
<< pdc >>
rect 17 35 20 38
rect 24 32 27 35
rect 31 35 34 38
rect 38 35 41 38
<< ptransistor >>
rect 21 31 23 39
rect 28 31 30 39
rect 35 31 37 39
<< polysilicon >>
rect 24 48 30 49
rect 24 45 25 48
rect 28 45 30 48
rect 24 44 30 45
rect 21 39 23 41
rect 28 39 30 44
rect 35 39 37 41
rect 21 24 23 31
rect 28 24 30 31
rect 35 28 37 31
rect 35 27 49 28
rect 35 26 45 27
rect 35 24 37 26
rect 44 24 45 26
rect 48 24 49 27
rect 44 23 49 24
rect 35 16 37 18
rect 21 12 23 14
rect 28 12 30 14
rect 16 11 23 12
rect 16 8 17 11
rect 20 8 23 11
rect 16 7 23 8
<< pc >>
rect 25 45 28 48
rect 45 24 48 27
rect 17 8 20 11
<< m1 >>
rect 16 48 20 52
rect 17 45 25 48
rect 28 45 29 48
rect 48 43 52 44
rect 38 40 52 43
rect 17 38 20 39
rect 31 38 34 39
rect 17 34 20 35
rect 24 35 27 36
rect 31 34 34 35
rect 38 38 41 40
rect 17 27 20 28
rect 17 23 20 24
rect 24 27 27 32
rect 24 23 27 24
rect 38 23 41 35
rect 45 27 48 28
rect 45 23 48 24
rect 17 19 20 20
rect 31 22 34 23
rect 38 19 41 20
rect 31 16 34 19
rect 31 13 32 16
rect 35 13 36 16
rect 31 12 36 13
rect 9 8 17 11
rect 20 8 21 11
rect 8 4 12 8
<< m2c >>
rect 17 35 20 38
rect 31 35 34 38
rect 17 24 20 27
rect 24 24 27 27
rect 45 24 48 27
rect 32 13 35 16
<< m2 >>
rect 16 38 35 39
rect 16 35 17 38
rect 20 35 31 38
rect 34 35 35 38
rect 16 34 35 35
rect 16 27 49 28
rect 16 24 17 27
rect 20 24 24 27
rect 27 24 45 27
rect 48 24 49 27
rect 16 23 49 24
rect 31 16 36 17
rect 31 13 32 16
rect 35 13 36 16
rect 31 12 36 13
<< labels >>
rlabel space 0 0 56 56 6 prboundary
rlabel ndiffusion 42 21 42 21 3 Y
rlabel polysilicon 45 24 45 24 3 _Y
rlabel polysilicon 45 25 45 25 3 _Y
rlabel pdiffusion 42 36 42 36 3 Y
rlabel polysilicon 36 17 36 17 3 _Y
rlabel ndiffusion 38 19 38 19 3 Y
rlabel ndiffusion 38 21 38 21 3 Y
rlabel ndiffusion 38 24 38 24 3 Y
rlabel ndiffusion 35 20 35 20 3 GND
rlabel pdiffusion 38 32 38 32 3 Y
rlabel pdiffusion 38 36 38 36 3 Y
rlabel pdiffusion 38 39 38 39 3 Y
rlabel polysilicon 36 40 36 40 3 _Y
rlabel ntransistor 36 19 36 19 3 _Y
rlabel polysilicon 36 25 36 25 3 _Y
rlabel polysilicon 36 27 36 27 3 _Y
rlabel polysilicon 36 28 36 28 3 _Y
rlabel polysilicon 36 29 36 29 3 _Y
rlabel ptransistor 36 32 36 32 3 _Y
rlabel ndiffusion 31 15 31 15 3 GND
rlabel ndiffusion 31 19 31 19 3 GND
rlabel ndiffusion 31 20 31 20 3 GND
rlabel ndiffusion 31 23 31 23 3 GND
rlabel pdiffusion 31 32 31 32 3 Vdd
rlabel pdiffusion 31 36 31 36 3 Vdd
rlabel pdiffusion 31 39 31 39 3 Vdd
rlabel pdiffusion 28 33 28 33 3 _Y
rlabel polysilicon 29 40 29 40 3 A
rlabel polysilicon 29 13 29 13 3 A
rlabel ntransistor 29 15 29 15 3 A
rlabel polysilicon 29 25 29 25 3 A
rlabel ptransistor 29 32 29 32 3 A
rlabel polysilicon 25 45 25 45 3 A
rlabel polysilicon 25 46 25 46 3 A
rlabel polysilicon 25 49 25 49 3 A
rlabel ndiffusion 21 21 21 21 3 _Y
rlabel pdiffusion 24 32 24 32 3 _Y
rlabel pdiffusion 24 33 24 33 3 _Y
rlabel pdiffusion 24 36 24 36 3 _Y
rlabel polysilicon 22 13 22 13 3 B
rlabel ntransistor 22 15 22 15 3 B
rlabel polysilicon 22 25 22 25 3 B
rlabel ptransistor 22 32 22 32 3 B
rlabel polysilicon 22 40 22 40 3 B
rlabel polysilicon 17 8 17 8 3 B
rlabel polysilicon 17 9 17 9 3 B
rlabel polysilicon 17 12 17 12 3 B
rlabel ndiffusion 17 15 17 15 3 _Y
rlabel ndiffusion 17 21 17 21 3 _Y
rlabel pdiffusion 17 32 17 32 3 Vdd
rlabel m1 49 44 49 44 3 Y
port 1 e
rlabel m1 46 24 46 24 3 _Y
rlabel m1 46 28 46 28 3 _Y
rlabel m1 39 20 39 20 3 Y
port 1 e
rlabel ndc 39 21 39 21 3 Y
port 1 e
rlabel m1 39 24 39 24 3 Y
port 1 e
rlabel pdc 39 36 39 36 3 Y
port 1 e
rlabel m1 39 39 39 39 3 Y
port 1 e
rlabel m1 39 41 39 41 3 Y
port 1 e
rlabel m1 32 35 32 35 3 Vdd
rlabel m1 32 39 32 39 3 Vdd
rlabel m1 32 23 32 23 3 GND
rlabel ndc 32 20 32 20 3 GND
rlabel m1 25 24 25 24 3 _Y
rlabel m1 25 28 25 28 3 _Y
rlabel pdc 25 33 25 33 3 _Y
rlabel m1 25 36 25 36 3 _Y
rlabel m1 29 46 29 46 3 A
port 2 e
rlabel pc 26 46 26 46 3 A
port 2 e
rlabel m1 21 9 21 9 3 B
port 3 e
rlabel m1 18 20 18 20 3 _Y
rlabel ndc 18 21 18 21 3 _Y
rlabel m1 18 24 18 24 3 _Y
rlabel m1 18 28 18 28 3 _Y
rlabel m1 18 35 18 35 3 Vdd
rlabel m1 18 39 18 39 3 Vdd
rlabel m1 18 46 18 46 3 A
port 2 e
rlabel pc 18 9 18 9 3 B
port 3 e
rlabel m1 17 49 17 49 3 A
port 2 e
rlabel m1 10 9 10 9 3 B
port 3 e
rlabel m1 9 5 9 5 3 B
port 3 e
rlabel m2 49 25 49 25 3 _Y
rlabel m2c 46 25 46 25 3 _Y
rlabel m2 36 14 36 14 3 GND
rlabel m2 28 25 28 25 3 _Y
rlabel m2 35 36 35 36 3 Vdd
rlabel m2c 33 14 33 14 3 GND
rlabel m2c 25 25 25 25 3 _Y
rlabel m2c 32 36 32 36 3 Vdd
rlabel m2 32 13 32 13 3 GND
rlabel m2 32 14 32 14 3 GND
rlabel m2 32 17 32 17 3 GND
rlabel m2 21 25 21 25 3 _Y
rlabel m2 21 36 21 36 3 Vdd
rlabel m2c 18 25 18 25 3 _Y
rlabel m2c 18 36 18 36 3 Vdd
rlabel m2 17 24 17 24 3 _Y
rlabel m2 17 25 17 25 3 _Y
rlabel m2 17 28 17 28 3 _Y
rlabel m2 17 35 17 35 3 Vdd
rlabel m2 17 36 17 36 3 Vdd
rlabel m2 17 39 17 39 3 Vdd
<< end >>
