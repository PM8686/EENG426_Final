magic
tech TSMC180
timestamp 1734130717
<< ndiffusion >>
rect 6 15 12 22
rect 6 13 7 15
rect 9 13 12 15
rect 6 12 12 13
rect 14 12 20 22
rect 22 15 28 22
rect 32 21 38 22
rect 32 19 33 21
rect 35 19 38 21
rect 32 17 38 19
rect 40 20 48 22
rect 40 18 43 20
rect 45 18 48 20
rect 40 17 48 18
rect 22 13 25 15
rect 27 13 28 15
rect 22 12 28 13
rect 44 12 48 17
rect 50 21 56 22
rect 50 19 53 21
rect 55 19 56 21
rect 50 12 56 19
rect 60 15 66 22
rect 60 13 63 15
rect 65 13 66 15
rect 60 12 66 13
rect 68 21 74 22
rect 68 19 70 21
rect 72 19 74 21
rect 68 12 74 19
<< ndcontact >>
rect 7 13 9 15
rect 33 19 35 21
rect 43 18 45 20
rect 25 13 27 15
rect 53 19 55 21
rect 63 13 65 15
rect 70 19 72 21
<< ntransistor >>
rect 12 12 14 22
rect 20 12 22 22
rect 38 17 40 22
rect 48 12 50 22
rect 66 12 68 22
<< pdiffusion >>
rect 6 41 12 53
rect 6 39 7 41
rect 9 39 12 41
rect 6 38 12 39
rect 14 52 18 53
rect 14 50 15 52
rect 17 50 18 52
rect 14 46 18 50
rect 14 38 20 46
rect 22 41 28 46
rect 22 39 25 41
rect 27 39 28 41
rect 22 38 28 39
rect 32 43 38 53
rect 32 41 34 43
rect 36 41 38 43
rect 32 38 38 41
rect 40 38 48 53
rect 50 49 56 53
rect 50 47 52 49
rect 54 47 56 49
rect 50 38 56 47
rect 60 38 66 53
rect 68 43 74 53
rect 68 41 70 43
rect 72 41 74 43
rect 68 38 74 41
<< pdcontact >>
rect 7 39 9 41
rect 15 50 17 52
rect 25 39 27 41
rect 34 41 36 43
rect 52 47 54 49
rect 70 41 72 43
<< ptransistor >>
rect 12 38 14 53
rect 20 38 22 46
rect 38 38 40 53
rect 48 38 50 53
rect 66 38 68 53
<< polysilicon >>
rect 6 59 14 60
rect 6 57 7 59
rect 9 57 14 59
rect 6 56 14 57
rect 12 53 14 56
rect 38 59 44 60
rect 38 57 41 59
rect 43 57 44 59
rect 38 56 44 57
rect 48 59 60 60
rect 48 57 57 59
rect 59 57 60 59
rect 48 56 60 57
rect 38 53 40 56
rect 48 53 50 56
rect 66 53 68 56
rect 20 46 22 49
rect 12 22 14 38
rect 20 22 22 38
rect 38 22 40 38
rect 48 22 50 38
rect 66 36 68 38
rect 66 35 70 36
rect 66 33 67 35
rect 69 33 70 35
rect 66 32 70 33
rect 66 22 68 32
rect 12 9 14 12
rect 20 9 22 12
rect 38 9 40 17
rect 48 9 50 12
rect 66 9 68 12
rect 20 7 40 9
rect 20 -4 22 7
rect 20 -5 24 -4
rect 20 -7 21 -5
rect 23 -7 24 -5
rect 20 -8 24 -7
<< polycontact >>
rect 7 57 9 59
rect 41 57 43 59
rect 57 57 59 59
rect 67 33 69 35
rect 21 -7 23 -5
<< m1 >>
rect -3 67 2 68
rect -3 64 -2 67
rect 1 64 2 67
rect -3 63 2 64
rect 6 59 10 76
rect 24 60 27 76
rect 42 60 45 76
rect 6 57 7 59
rect 9 57 10 59
rect 6 56 10 57
rect 15 57 27 60
rect 40 59 45 60
rect 40 57 41 59
rect 43 57 45 59
rect 55 60 58 76
rect 61 67 66 68
rect 61 64 62 67
rect 65 64 66 67
rect 61 63 66 64
rect 55 59 63 60
rect 55 57 57 59
rect 59 57 63 59
rect 15 53 18 57
rect 40 56 44 57
rect 55 56 63 57
rect 14 52 19 53
rect 14 49 15 52
rect 18 49 19 52
rect 61 52 66 53
rect 14 48 19 49
rect 51 50 56 51
rect 51 47 52 50
rect 55 47 56 50
rect 61 49 62 52
rect 65 49 66 52
rect 61 48 66 49
rect 51 46 56 47
rect 33 43 37 44
rect 69 43 73 44
rect -3 42 2 43
rect -3 39 -2 42
rect 1 39 2 42
rect -3 38 2 39
rect 6 42 11 43
rect 6 39 7 42
rect 10 39 11 42
rect 6 38 11 39
rect 24 41 29 43
rect 24 39 25 41
rect 27 39 29 41
rect 33 41 34 43
rect 36 41 70 43
rect 72 41 80 43
rect 33 40 80 41
rect 24 36 29 39
rect 24 33 25 36
rect 28 33 29 36
rect 24 32 29 33
rect 32 36 37 37
rect 32 33 33 36
rect 36 33 37 36
rect 32 21 37 33
rect 65 36 70 37
rect 65 33 66 36
rect 69 33 70 36
rect 65 32 70 33
rect 52 26 57 27
rect 52 23 53 26
rect 56 23 57 26
rect 52 22 57 23
rect 69 26 74 27
rect 69 23 70 26
rect 73 23 74 26
rect 69 22 74 23
rect 52 21 56 22
rect 32 19 33 21
rect 35 19 37 21
rect 32 17 37 19
rect 42 20 46 21
rect 42 18 43 20
rect 45 18 46 20
rect 52 19 53 21
rect 55 19 56 21
rect 52 18 56 19
rect 69 21 73 22
rect 69 19 70 21
rect 72 19 73 21
rect 69 18 73 19
rect 42 17 46 18
rect 6 15 10 16
rect 6 13 7 15
rect 9 13 10 15
rect 6 12 10 13
rect 24 15 29 16
rect 24 12 25 15
rect 28 12 29 15
rect 6 5 9 12
rect 24 11 29 12
rect 43 5 46 17
rect 77 16 80 40
rect 61 15 66 16
rect 61 12 62 15
rect 65 12 66 15
rect 61 11 66 12
rect 76 15 81 16
rect 76 12 77 15
rect 80 12 81 15
rect 76 11 81 12
rect 6 4 11 5
rect 6 1 7 4
rect 10 1 11 4
rect 6 0 11 1
rect 42 4 47 5
rect 42 1 43 4
rect 46 1 47 4
rect 42 0 47 1
rect 20 -5 24 -4
rect 20 -7 21 -5
rect 23 -7 24 -5
rect 20 -8 24 -7
<< m2c >>
rect -2 64 1 67
rect 62 64 65 67
rect 15 50 17 52
rect 17 50 18 52
rect 15 49 18 50
rect 52 49 55 50
rect 52 47 54 49
rect 54 47 55 49
rect 62 49 65 52
rect -2 39 1 42
rect 7 41 10 42
rect 7 39 9 41
rect 9 39 10 41
rect 25 33 28 36
rect 33 33 36 36
rect 66 35 69 36
rect 66 33 67 35
rect 67 33 69 35
rect 53 23 56 26
rect 70 23 73 26
rect 25 13 27 15
rect 27 13 28 15
rect 25 12 28 13
rect 62 13 63 15
rect 63 13 65 15
rect 62 12 65 13
rect 77 12 80 15
rect 7 1 10 4
rect 43 1 46 4
<< m2 >>
rect -3 67 66 68
rect -3 64 -2 67
rect 1 64 62 67
rect 65 64 66 67
rect -3 63 66 64
rect -3 43 2 63
rect 14 52 56 53
rect 14 49 15 52
rect 18 50 56 52
rect 18 49 52 50
rect 14 48 52 49
rect 51 47 52 48
rect 55 47 56 50
rect 61 52 66 63
rect 61 49 62 52
rect 65 49 66 52
rect 61 48 66 49
rect 51 46 56 47
rect -3 42 11 43
rect -3 39 -2 42
rect 1 39 7 42
rect 10 39 11 42
rect -3 38 11 39
rect 24 36 70 37
rect 24 33 25 36
rect 28 33 33 36
rect 36 33 66 36
rect 69 33 70 36
rect 24 32 70 33
rect 52 26 74 27
rect 52 23 53 26
rect 56 23 70 26
rect 73 23 74 26
rect 52 22 74 23
rect 24 15 81 16
rect 24 12 25 15
rect 28 12 62 15
rect 65 12 77 15
rect 80 12 81 15
rect 24 11 81 12
rect 6 4 47 5
rect 6 1 7 4
rect 10 1 43 4
rect 46 1 47 4
rect 6 0 47 1
<< labels >>
rlabel pdiffusion 23 39 23 39 3 _S
rlabel ndiffusion 23 13 23 13 3 Y
rlabel polysilicon 21 23 21 23 3 S
rlabel polysilicon 21 36 21 36 3 S
rlabel pdiffusion 15 39 15 39 3 Vdd
rlabel polysilicon 13 23 13 23 3 A
rlabel polysilicon 13 36 13 36 3 A
rlabel ndiffusion 7 13 7 13 3 GND
rlabel pdiffusion 7 39 7 39 3 #5
rlabel ndiffusion 51 13 51 13 3 #10
rlabel polysilicon 49 23 49 23 3 B
rlabel polysilicon 49 36 49 36 3 B
rlabel pdiffusion 51 39 51 39 3 Vdd
rlabel ndiffusion 41 18 41 18 3 GND
rlabel polysilicon 39 23 39 23 3 S
rlabel polysilicon 39 36 39 36 3 S
rlabel ndiffusion 33 18 33 18 3 _S
rlabel ndiffusion 69 13 69 13 3 #10
rlabel pdiffusion 69 39 69 39 3 Y
rlabel polysilicon 67 23 67 23 3 _S
rlabel polysilicon 67 36 67 36 3 _S
rlabel ndiffusion 61 13 61 13 3 Y
rlabel pdiffusion 61 39 61 39 3 #5
rlabel m1 43 58 43 58 3 S
port 3 e
rlabel m1 7 58 7 58 3 A
port 6 e
rlabel m1 7 11 7 11 2 GND
rlabel pdiffusion 35 48 35 48 1 Y
rlabel m1 61 58 61 58 5 B
rlabel m1 25 58 25 58 5 Vdd
rlabel m1 22 -7 22 -7 1 S
rlabel pdcontact 35 42 35 42 1 Y
rlabel m1 8 74 8 74 5 A
rlabel m1 25 74 25 74 5 Vdd
rlabel m1 44 74 44 74 5 S
rlabel m1 57 74 57 74 5 B
rlabel m1 79 41 79 41 7 Y
<< end >>
