magic
tech sky130l
timestamp 1731220673
<< m1 >>
rect 904 2047 908 2063
rect 1064 2047 1068 2063
rect 344 1823 348 1839
rect 1856 1803 1860 1819
rect 1960 1803 1964 1819
rect 1392 1595 1396 1615
rect 328 1367 332 1383
rect 184 1239 188 1255
rect 1136 1007 1140 1023
rect 1120 895 1124 911
rect 1808 811 1812 827
rect 344 679 348 695
rect 1696 587 1700 603
<< m2c >>
rect 172 2551 176 2555
rect 228 2551 232 2555
rect 284 2551 288 2555
rect 340 2551 344 2555
rect 396 2551 400 2555
rect 188 2531 192 2535
rect 244 2531 248 2535
rect 300 2531 304 2535
rect 356 2531 360 2535
rect 1532 2531 1536 2535
rect 1588 2531 1592 2535
rect 1644 2531 1648 2535
rect 1700 2531 1704 2535
rect 1756 2531 1760 2535
rect 1812 2531 1816 2535
rect 1868 2531 1872 2535
rect 1924 2531 1928 2535
rect 1980 2531 1984 2535
rect 2036 2531 2040 2535
rect 2092 2531 2096 2535
rect 2148 2531 2152 2535
rect 2204 2531 2208 2535
rect 204 2519 208 2523
rect 260 2519 264 2523
rect 324 2519 328 2523
rect 396 2519 400 2523
rect 468 2519 472 2523
rect 532 2519 536 2523
rect 596 2519 600 2523
rect 660 2519 664 2523
rect 724 2519 728 2523
rect 788 2519 792 2523
rect 852 2519 856 2523
rect 916 2519 920 2523
rect 980 2519 984 2523
rect 1044 2519 1048 2523
rect 1492 2511 1496 2515
rect 1548 2511 1552 2515
rect 1604 2511 1608 2515
rect 1660 2511 1664 2515
rect 1716 2511 1720 2515
rect 1772 2511 1776 2515
rect 1828 2511 1832 2515
rect 1884 2511 1888 2515
rect 1940 2511 1944 2515
rect 1996 2511 2000 2515
rect 2052 2511 2056 2515
rect 2108 2511 2112 2515
rect 2164 2511 2168 2515
rect 244 2499 248 2503
rect 300 2499 304 2503
rect 364 2499 368 2503
rect 436 2499 440 2503
rect 508 2499 512 2503
rect 572 2499 576 2503
rect 636 2499 640 2503
rect 700 2499 704 2503
rect 764 2499 768 2503
rect 828 2499 832 2503
rect 892 2499 896 2503
rect 956 2499 960 2503
rect 1020 2499 1024 2503
rect 1084 2499 1088 2503
rect 1524 2499 1528 2503
rect 1588 2499 1592 2503
rect 1660 2499 1664 2503
rect 1732 2499 1736 2503
rect 1804 2499 1808 2503
rect 1876 2499 1880 2503
rect 1948 2499 1952 2503
rect 2020 2499 2024 2503
rect 2092 2499 2096 2503
rect 2164 2499 2168 2503
rect 1564 2479 1568 2483
rect 1628 2479 1632 2483
rect 1700 2479 1704 2483
rect 1772 2479 1776 2483
rect 1844 2479 1848 2483
rect 1916 2479 1920 2483
rect 1988 2479 1992 2483
rect 2060 2479 2064 2483
rect 2132 2479 2136 2483
rect 2204 2479 2208 2483
rect 204 2439 208 2443
rect 260 2439 264 2443
rect 316 2439 320 2443
rect 372 2439 376 2443
rect 428 2439 432 2443
rect 484 2439 488 2443
rect 540 2439 544 2443
rect 596 2439 600 2443
rect 652 2439 656 2443
rect 708 2439 712 2443
rect 764 2439 768 2443
rect 820 2439 824 2443
rect 876 2439 880 2443
rect 932 2439 936 2443
rect 988 2439 992 2443
rect 1044 2439 1048 2443
rect 1100 2439 1104 2443
rect 164 2419 168 2423
rect 220 2419 224 2423
rect 276 2419 280 2423
rect 332 2419 336 2423
rect 388 2419 392 2423
rect 444 2419 448 2423
rect 500 2419 504 2423
rect 556 2419 560 2423
rect 612 2419 616 2423
rect 668 2419 672 2423
rect 724 2419 728 2423
rect 780 2419 784 2423
rect 836 2419 840 2423
rect 892 2419 896 2423
rect 948 2421 952 2425
rect 1004 2421 1008 2425
rect 1580 2423 1584 2427
rect 1644 2423 1648 2427
rect 1708 2423 1712 2427
rect 1780 2423 1784 2427
rect 1852 2423 1856 2427
rect 1916 2423 1920 2427
rect 1988 2423 1992 2427
rect 2060 2423 2064 2427
rect 2132 2423 2136 2427
rect 2204 2423 2208 2427
rect 1060 2419 1064 2423
rect 1540 2405 1544 2409
rect 1604 2405 1608 2409
rect 1668 2405 1672 2409
rect 1740 2405 1744 2409
rect 1812 2403 1816 2407
rect 1876 2403 1880 2407
rect 1948 2403 1952 2407
rect 2020 2405 2024 2409
rect 2092 2405 2096 2409
rect 2164 2403 2168 2407
rect 500 2395 504 2399
rect 556 2395 560 2399
rect 612 2395 616 2399
rect 668 2395 672 2399
rect 1548 2387 1552 2391
rect 1604 2387 1608 2391
rect 1660 2387 1664 2391
rect 1716 2387 1720 2391
rect 1772 2387 1776 2391
rect 1836 2387 1840 2391
rect 1900 2387 1904 2391
rect 1964 2387 1968 2391
rect 2028 2387 2032 2391
rect 2092 2387 2096 2391
rect 540 2375 544 2379
rect 596 2377 600 2381
rect 652 2377 656 2381
rect 708 2377 712 2381
rect 1588 2367 1592 2371
rect 1644 2367 1648 2371
rect 1700 2367 1704 2371
rect 1756 2367 1760 2371
rect 1812 2367 1816 2371
rect 1876 2367 1880 2371
rect 1940 2369 1944 2373
rect 2004 2367 2008 2371
rect 2068 2367 2072 2371
rect 2132 2369 2136 2373
rect 356 2315 360 2319
rect 428 2315 432 2319
rect 500 2315 504 2319
rect 572 2315 576 2319
rect 644 2315 648 2319
rect 716 2315 720 2319
rect 780 2315 784 2319
rect 844 2315 848 2319
rect 900 2315 904 2319
rect 964 2315 968 2319
rect 1028 2315 1032 2319
rect 1092 2315 1096 2319
rect 1148 2315 1152 2319
rect 1204 2315 1208 2319
rect 1260 2315 1264 2319
rect 1508 2307 1512 2311
rect 1572 2307 1576 2311
rect 1644 2307 1648 2311
rect 1724 2307 1728 2311
rect 1796 2307 1800 2311
rect 1868 2307 1872 2311
rect 1940 2307 1944 2311
rect 2020 2307 2024 2311
rect 2100 2307 2104 2311
rect 2180 2307 2184 2311
rect 316 2297 320 2301
rect 388 2295 392 2299
rect 460 2297 464 2301
rect 532 2295 536 2299
rect 604 2295 608 2299
rect 676 2295 680 2299
rect 740 2297 744 2301
rect 804 2297 808 2301
rect 860 2297 864 2301
rect 924 2297 928 2301
rect 988 2295 992 2299
rect 1052 2297 1056 2301
rect 1108 2297 1112 2301
rect 1164 2297 1168 2301
rect 1220 2295 1224 2299
rect 1468 2287 1472 2291
rect 1532 2287 1536 2291
rect 1604 2287 1608 2291
rect 1684 2287 1688 2291
rect 1756 2287 1760 2291
rect 1828 2287 1832 2291
rect 1900 2287 1904 2291
rect 1980 2287 1984 2291
rect 2060 2287 2064 2291
rect 2140 2287 2144 2291
rect 156 2275 160 2279
rect 252 2275 256 2279
rect 356 2275 360 2279
rect 460 2275 464 2279
rect 572 2275 576 2279
rect 684 2275 688 2279
rect 788 2275 792 2279
rect 892 2275 896 2279
rect 996 2275 1000 2279
rect 1108 2275 1112 2279
rect 1220 2275 1224 2279
rect 1364 2275 1368 2279
rect 1460 2275 1464 2279
rect 1564 2275 1568 2279
rect 1668 2275 1672 2279
rect 1772 2275 1776 2279
rect 1884 2275 1888 2279
rect 1996 2275 2000 2279
rect 2108 2275 2112 2279
rect 2220 2275 2224 2279
rect 196 2255 200 2259
rect 292 2257 296 2261
rect 396 2257 400 2261
rect 500 2255 504 2259
rect 612 2257 616 2261
rect 724 2255 728 2259
rect 828 2255 832 2259
rect 932 2255 936 2259
rect 1036 2255 1040 2259
rect 1148 2255 1152 2259
rect 1260 2255 1264 2259
rect 1404 2255 1408 2259
rect 1500 2255 1504 2259
rect 1604 2255 1608 2259
rect 1708 2255 1712 2259
rect 1812 2257 1816 2261
rect 1924 2255 1928 2259
rect 2036 2255 2040 2259
rect 2148 2255 2152 2259
rect 2260 2255 2264 2259
rect 180 2203 184 2207
rect 268 2203 272 2207
rect 356 2203 360 2207
rect 452 2203 456 2207
rect 556 2203 560 2207
rect 660 2203 664 2207
rect 764 2203 768 2207
rect 868 2203 872 2207
rect 972 2203 976 2207
rect 1076 2203 1080 2207
rect 1180 2203 1184 2207
rect 1260 2203 1264 2207
rect 1404 2203 1408 2207
rect 1524 2203 1528 2207
rect 1644 2203 1648 2207
rect 1756 2203 1760 2207
rect 1852 2203 1856 2207
rect 1940 2203 1944 2207
rect 2020 2203 2024 2207
rect 2092 2203 2096 2207
rect 2164 2203 2168 2207
rect 2228 2203 2232 2207
rect 2292 2203 2296 2207
rect 2356 2203 2360 2207
rect 2420 2203 2424 2207
rect 2476 2203 2480 2207
rect 140 2183 144 2187
rect 228 2183 232 2187
rect 316 2183 320 2187
rect 412 2183 416 2187
rect 516 2183 520 2187
rect 620 2183 624 2187
rect 724 2185 728 2189
rect 828 2185 832 2189
rect 932 2183 936 2187
rect 1036 2185 1040 2189
rect 1140 2183 1144 2187
rect 1220 2183 1224 2187
rect 1364 2185 1368 2189
rect 1484 2183 1488 2187
rect 1604 2183 1608 2187
rect 1716 2183 1720 2187
rect 1812 2183 1816 2187
rect 1900 2183 1904 2187
rect 1980 2183 1984 2187
rect 2052 2183 2056 2187
rect 2124 2183 2128 2187
rect 2188 2183 2192 2187
rect 2252 2183 2256 2187
rect 2316 2183 2320 2187
rect 2380 2183 2384 2187
rect 2436 2183 2440 2187
rect 236 2171 240 2175
rect 332 2171 336 2175
rect 436 2171 440 2175
rect 540 2171 544 2175
rect 644 2171 648 2175
rect 748 2171 752 2175
rect 844 2171 848 2175
rect 940 2171 944 2175
rect 1036 2171 1040 2175
rect 1140 2171 1144 2175
rect 1220 2171 1224 2175
rect 276 2151 280 2155
rect 372 2151 376 2155
rect 476 2151 480 2155
rect 580 2151 584 2155
rect 684 2151 688 2155
rect 788 2151 792 2155
rect 884 2151 888 2155
rect 980 2151 984 2155
rect 1076 2151 1080 2155
rect 1180 2153 1184 2157
rect 1260 2153 1264 2157
rect 1388 2151 1392 2155
rect 1604 2151 1608 2155
rect 1796 2151 1800 2155
rect 1972 2151 1976 2155
rect 2140 2151 2144 2155
rect 2300 2151 2304 2155
rect 2436 2151 2440 2155
rect 1428 2131 1432 2135
rect 1644 2133 1648 2137
rect 1836 2131 1840 2135
rect 2012 2131 2016 2135
rect 2180 2133 2184 2137
rect 2340 2133 2344 2137
rect 2476 2133 2480 2137
rect 340 2099 344 2103
rect 396 2099 400 2103
rect 460 2099 464 2103
rect 524 2099 528 2103
rect 596 2099 600 2103
rect 668 2099 672 2103
rect 748 2099 752 2103
rect 836 2099 840 2103
rect 924 2099 928 2103
rect 1012 2099 1016 2103
rect 1100 2099 1104 2103
rect 1188 2099 1192 2103
rect 1260 2099 1264 2103
rect 300 2081 304 2085
rect 356 2079 360 2083
rect 420 2079 424 2083
rect 484 2079 488 2083
rect 556 2079 560 2083
rect 628 2079 632 2083
rect 708 2081 712 2085
rect 796 2079 800 2083
rect 884 2081 888 2085
rect 972 2079 976 2083
rect 1060 2079 1064 2083
rect 1148 2079 1152 2083
rect 1220 2079 1224 2083
rect 1420 2079 1424 2083
rect 1588 2079 1592 2083
rect 1748 2079 1752 2083
rect 1892 2079 1896 2083
rect 2028 2079 2032 2083
rect 2156 2079 2160 2083
rect 2276 2079 2280 2083
rect 2404 2079 2408 2083
rect 380 2065 384 2069
rect 436 2063 440 2067
rect 492 2063 496 2067
rect 556 2063 560 2067
rect 620 2063 624 2067
rect 692 2063 696 2067
rect 772 2063 776 2067
rect 844 2063 848 2067
rect 904 2063 908 2067
rect 924 2063 928 2067
rect 1004 2063 1008 2067
rect 1064 2063 1068 2067
rect 1084 2063 1088 2067
rect 1164 2063 1168 2067
rect 1220 2063 1224 2067
rect 420 2043 424 2047
rect 476 2043 480 2047
rect 532 2045 536 2049
rect 596 2045 600 2049
rect 660 2045 664 2049
rect 732 2043 736 2047
rect 812 2045 816 2049
rect 884 2043 888 2047
rect 904 2043 908 2047
rect 964 2045 968 2049
rect 1380 2059 1384 2063
rect 1548 2059 1552 2063
rect 1708 2059 1712 2063
rect 1852 2061 1856 2065
rect 1988 2061 1992 2065
rect 2116 2059 2120 2063
rect 2236 2059 2240 2063
rect 2364 2059 2368 2063
rect 1044 2043 1048 2047
rect 1064 2043 1068 2047
rect 1124 2043 1128 2047
rect 1204 2043 1208 2047
rect 1260 2045 1264 2049
rect 1428 2043 1432 2047
rect 1532 2043 1536 2047
rect 1636 2043 1640 2047
rect 1732 2043 1736 2047
rect 1820 2043 1824 2047
rect 1908 2043 1912 2047
rect 2004 2043 2008 2047
rect 2100 2043 2104 2047
rect 1468 2023 1472 2027
rect 1572 2023 1576 2027
rect 1676 2025 1680 2029
rect 1772 2023 1776 2027
rect 1860 2025 1864 2029
rect 1948 2023 1952 2027
rect 2044 2023 2048 2027
rect 2140 2025 2144 2029
rect 268 1987 272 1991
rect 324 1987 328 1991
rect 396 1987 400 1991
rect 476 1987 480 1991
rect 572 1987 576 1991
rect 668 1987 672 1991
rect 772 1987 776 1991
rect 884 1987 888 1991
rect 996 1987 1000 1991
rect 1116 1987 1120 1991
rect 1236 1987 1240 1991
rect 228 1967 232 1971
rect 284 1967 288 1971
rect 356 1967 360 1971
rect 436 1967 440 1971
rect 532 1967 536 1971
rect 628 1967 632 1971
rect 732 1967 736 1971
rect 844 1967 848 1971
rect 956 1969 960 1973
rect 1076 1967 1080 1971
rect 1196 1967 1200 1971
rect 1492 1967 1496 1971
rect 1548 1967 1552 1971
rect 1612 1967 1616 1971
rect 1676 1967 1680 1971
rect 1740 1967 1744 1971
rect 1804 1967 1808 1971
rect 1868 1967 1872 1971
rect 1932 1967 1936 1971
rect 1996 1967 2000 1971
rect 2068 1967 2072 1971
rect 132 1951 136 1955
rect 196 1951 200 1955
rect 300 1951 304 1955
rect 420 1951 424 1955
rect 564 1951 568 1955
rect 724 1951 728 1955
rect 900 1951 904 1955
rect 1076 1951 1080 1955
rect 1452 1947 1456 1951
rect 1508 1947 1512 1951
rect 1572 1949 1576 1953
rect 1636 1949 1640 1953
rect 1700 1947 1704 1951
rect 1764 1947 1768 1951
rect 1828 1947 1832 1951
rect 1892 1947 1896 1951
rect 1956 1947 1960 1951
rect 2028 1947 2032 1951
rect 172 1931 176 1935
rect 236 1931 240 1935
rect 340 1931 344 1935
rect 460 1931 464 1935
rect 604 1931 608 1935
rect 764 1931 768 1935
rect 940 1933 944 1937
rect 1116 1931 1120 1935
rect 1548 1931 1552 1935
rect 1612 1931 1616 1935
rect 1684 1931 1688 1935
rect 1756 1931 1760 1935
rect 1828 1931 1832 1935
rect 1900 1933 1904 1937
rect 1980 1931 1984 1935
rect 2068 1931 2072 1935
rect 2164 1931 2168 1935
rect 2260 1931 2264 1935
rect 2356 1931 2360 1935
rect 2436 1931 2440 1935
rect 1588 1911 1592 1915
rect 1652 1911 1656 1915
rect 1724 1911 1728 1915
rect 1796 1911 1800 1915
rect 1868 1913 1872 1917
rect 1940 1911 1944 1915
rect 2020 1911 2024 1915
rect 2108 1911 2112 1915
rect 2204 1911 2208 1915
rect 2300 1911 2304 1915
rect 2396 1911 2400 1915
rect 2476 1911 2480 1915
rect 172 1871 176 1875
rect 228 1871 232 1875
rect 308 1871 312 1875
rect 396 1871 400 1875
rect 492 1871 496 1875
rect 580 1871 584 1875
rect 668 1871 672 1875
rect 756 1871 760 1875
rect 836 1871 840 1875
rect 908 1871 912 1875
rect 980 1871 984 1875
rect 1052 1871 1056 1875
rect 1124 1871 1128 1875
rect 1196 1871 1200 1875
rect 132 1853 136 1857
rect 188 1853 192 1857
rect 268 1853 272 1857
rect 356 1851 360 1855
rect 452 1851 456 1855
rect 540 1853 544 1857
rect 628 1853 632 1857
rect 1644 1855 1648 1859
rect 1700 1855 1704 1859
rect 1764 1855 1768 1859
rect 1836 1855 1840 1859
rect 1908 1855 1912 1859
rect 1980 1855 1984 1859
rect 2044 1855 2048 1859
rect 2108 1855 2112 1859
rect 2172 1855 2176 1859
rect 2236 1855 2240 1859
rect 2300 1855 2304 1859
rect 2364 1855 2368 1859
rect 2420 1855 2424 1859
rect 2476 1855 2480 1859
rect 716 1851 720 1855
rect 796 1851 800 1855
rect 868 1851 872 1855
rect 940 1851 944 1855
rect 1012 1851 1016 1855
rect 1084 1851 1088 1855
rect 1156 1851 1160 1855
rect 132 1839 136 1843
rect 188 1839 192 1843
rect 276 1839 280 1843
rect 344 1839 348 1843
rect 372 1839 376 1843
rect 476 1839 480 1843
rect 572 1839 576 1843
rect 668 1841 672 1845
rect 756 1839 760 1843
rect 836 1839 840 1843
rect 908 1839 912 1843
rect 980 1839 984 1843
rect 1060 1839 1064 1843
rect 1140 1839 1144 1843
rect 1604 1837 1608 1841
rect 1660 1835 1664 1839
rect 1724 1835 1728 1839
rect 1796 1835 1800 1839
rect 1868 1837 1872 1841
rect 1940 1835 1944 1839
rect 2004 1837 2008 1841
rect 2068 1835 2072 1839
rect 2132 1835 2136 1839
rect 2196 1835 2200 1839
rect 2260 1835 2264 1839
rect 2324 1835 2328 1839
rect 2380 1835 2384 1839
rect 2436 1835 2440 1839
rect 172 1819 176 1823
rect 228 1819 232 1823
rect 316 1819 320 1823
rect 344 1819 348 1823
rect 412 1819 416 1823
rect 516 1819 520 1823
rect 612 1819 616 1823
rect 708 1819 712 1823
rect 796 1819 800 1823
rect 876 1821 880 1825
rect 948 1819 952 1823
rect 1020 1819 1024 1823
rect 1100 1819 1104 1823
rect 1180 1819 1184 1823
rect 1612 1819 1616 1823
rect 1700 1819 1704 1823
rect 1796 1819 1800 1823
rect 1856 1819 1860 1823
rect 1908 1819 1912 1823
rect 1960 1819 1964 1823
rect 2036 1819 2040 1823
rect 2172 1819 2176 1823
rect 2316 1819 2320 1823
rect 2436 1819 2440 1823
rect 1652 1799 1656 1803
rect 1740 1799 1744 1803
rect 1836 1799 1840 1803
rect 1856 1799 1860 1803
rect 1948 1799 1952 1803
rect 1960 1799 1964 1803
rect 2076 1801 2080 1805
rect 2212 1799 2216 1803
rect 2356 1801 2360 1805
rect 2476 1799 2480 1803
rect 172 1755 176 1759
rect 236 1755 240 1759
rect 332 1755 336 1759
rect 436 1755 440 1759
rect 540 1755 544 1759
rect 644 1755 648 1759
rect 740 1755 744 1759
rect 836 1755 840 1759
rect 924 1755 928 1759
rect 1012 1755 1016 1759
rect 1100 1755 1104 1759
rect 1188 1755 1192 1759
rect 1564 1747 1568 1751
rect 1644 1747 1648 1751
rect 1732 1747 1736 1751
rect 1828 1747 1832 1751
rect 1916 1747 1920 1751
rect 2004 1747 2008 1751
rect 2092 1747 2096 1751
rect 2172 1747 2176 1751
rect 2252 1747 2256 1751
rect 2332 1747 2336 1751
rect 2412 1747 2416 1751
rect 2476 1747 2480 1751
rect 132 1735 136 1739
rect 196 1735 200 1739
rect 292 1735 296 1739
rect 396 1735 400 1739
rect 500 1737 504 1741
rect 604 1735 608 1739
rect 700 1735 704 1739
rect 796 1735 800 1739
rect 884 1735 888 1739
rect 972 1737 976 1741
rect 1060 1737 1064 1741
rect 1148 1735 1152 1739
rect 1524 1727 1528 1731
rect 1604 1727 1608 1731
rect 1692 1727 1696 1731
rect 1788 1727 1792 1731
rect 1876 1727 1880 1731
rect 1964 1729 1968 1733
rect 2052 1727 2056 1731
rect 2132 1729 2136 1733
rect 2212 1727 2216 1731
rect 2292 1729 2296 1733
rect 2372 1727 2376 1731
rect 2436 1727 2440 1731
rect 148 1721 152 1725
rect 220 1719 224 1723
rect 300 1719 304 1723
rect 388 1719 392 1723
rect 484 1719 488 1723
rect 588 1719 592 1723
rect 692 1719 696 1723
rect 804 1719 808 1723
rect 916 1719 920 1723
rect 1028 1719 1032 1723
rect 1140 1719 1144 1723
rect 1380 1711 1384 1715
rect 1444 1711 1448 1715
rect 1524 1711 1528 1715
rect 1612 1711 1616 1715
rect 1708 1711 1712 1715
rect 1804 1711 1808 1715
rect 1900 1711 1904 1715
rect 1996 1711 2000 1715
rect 2092 1711 2096 1715
rect 2180 1711 2184 1715
rect 2268 1711 2272 1715
rect 2364 1711 2368 1715
rect 2436 1711 2440 1715
rect 188 1699 192 1703
rect 260 1699 264 1703
rect 340 1699 344 1703
rect 428 1699 432 1703
rect 524 1699 528 1703
rect 628 1699 632 1703
rect 732 1699 736 1703
rect 844 1701 848 1705
rect 956 1699 960 1703
rect 1068 1699 1072 1703
rect 1180 1699 1184 1703
rect 1420 1691 1424 1695
rect 1484 1691 1488 1695
rect 1564 1691 1568 1695
rect 1652 1691 1656 1695
rect 1748 1691 1752 1695
rect 1844 1691 1848 1695
rect 1940 1691 1944 1695
rect 2036 1691 2040 1695
rect 2132 1691 2136 1695
rect 2220 1693 2224 1697
rect 2308 1691 2312 1695
rect 2404 1691 2408 1695
rect 2476 1691 2480 1695
rect 292 1643 296 1647
rect 356 1643 360 1647
rect 436 1643 440 1647
rect 524 1643 528 1647
rect 612 1643 616 1647
rect 708 1643 712 1647
rect 804 1643 808 1647
rect 900 1643 904 1647
rect 996 1643 1000 1647
rect 1100 1643 1104 1647
rect 1204 1643 1208 1647
rect 1388 1635 1392 1639
rect 1444 1635 1448 1639
rect 1532 1635 1536 1639
rect 1620 1635 1624 1639
rect 1716 1635 1720 1639
rect 1820 1635 1824 1639
rect 1932 1635 1936 1639
rect 2060 1635 2064 1639
rect 2196 1635 2200 1639
rect 2340 1635 2344 1639
rect 2476 1635 2480 1639
rect 252 1625 256 1629
rect 316 1623 320 1627
rect 396 1623 400 1627
rect 484 1623 488 1627
rect 572 1623 576 1627
rect 668 1623 672 1627
rect 764 1623 768 1627
rect 860 1623 864 1627
rect 956 1625 960 1629
rect 1060 1623 1064 1627
rect 1164 1623 1168 1627
rect 1348 1615 1352 1619
rect 1392 1615 1396 1619
rect 1404 1615 1408 1619
rect 1492 1615 1496 1619
rect 1580 1615 1584 1619
rect 1676 1615 1680 1619
rect 1780 1617 1784 1621
rect 1892 1615 1896 1619
rect 2020 1617 2024 1621
rect 2156 1615 2160 1619
rect 2300 1615 2304 1619
rect 2436 1615 2440 1619
rect 284 1609 288 1613
rect 340 1607 344 1611
rect 412 1607 416 1611
rect 492 1607 496 1611
rect 580 1607 584 1611
rect 676 1607 680 1611
rect 772 1607 776 1611
rect 876 1607 880 1611
rect 988 1607 992 1611
rect 1100 1607 1104 1611
rect 1348 1603 1352 1607
rect 1404 1603 1408 1607
rect 1460 1603 1464 1607
rect 1540 1603 1544 1607
rect 1620 1603 1624 1607
rect 1700 1603 1704 1607
rect 1772 1603 1776 1607
rect 1852 1603 1856 1607
rect 1932 1603 1936 1607
rect 2012 1603 2016 1607
rect 324 1587 328 1591
rect 380 1587 384 1591
rect 452 1587 456 1591
rect 532 1587 536 1591
rect 620 1589 624 1593
rect 716 1587 720 1591
rect 812 1589 816 1593
rect 916 1587 920 1591
rect 1028 1587 1032 1591
rect 1140 1589 1144 1593
rect 1392 1591 1396 1595
rect 1388 1583 1392 1587
rect 1444 1583 1448 1587
rect 1500 1583 1504 1587
rect 1580 1583 1584 1587
rect 1660 1585 1664 1589
rect 1740 1583 1744 1587
rect 1812 1585 1816 1589
rect 1892 1585 1896 1589
rect 1972 1583 1976 1587
rect 2052 1585 2056 1589
rect 284 1535 288 1539
rect 356 1535 360 1539
rect 436 1535 440 1539
rect 524 1535 528 1539
rect 620 1535 624 1539
rect 708 1535 712 1539
rect 796 1535 800 1539
rect 884 1535 888 1539
rect 964 1535 968 1539
rect 1044 1535 1048 1539
rect 1124 1535 1128 1539
rect 1204 1535 1208 1539
rect 1260 1535 1264 1539
rect 1388 1531 1392 1535
rect 1508 1531 1512 1535
rect 1644 1531 1648 1535
rect 1772 1531 1776 1535
rect 1908 1531 1912 1535
rect 2044 1531 2048 1535
rect 244 1515 248 1519
rect 316 1517 320 1521
rect 396 1517 400 1521
rect 484 1515 488 1519
rect 580 1515 584 1519
rect 668 1515 672 1519
rect 756 1515 760 1519
rect 844 1517 848 1521
rect 924 1517 928 1521
rect 1004 1515 1008 1519
rect 1084 1517 1088 1521
rect 1164 1515 1168 1519
rect 1220 1515 1224 1519
rect 1348 1511 1352 1515
rect 1468 1513 1472 1517
rect 1604 1511 1608 1515
rect 1732 1511 1736 1515
rect 1868 1511 1872 1515
rect 2004 1511 2008 1515
rect 1348 1499 1352 1503
rect 1404 1499 1408 1503
rect 1460 1499 1464 1503
rect 1532 1499 1536 1503
rect 1612 1499 1616 1503
rect 1692 1499 1696 1503
rect 1772 1499 1776 1503
rect 1852 1499 1856 1503
rect 1932 1499 1936 1503
rect 2012 1499 2016 1503
rect 2100 1499 2104 1503
rect 260 1495 264 1499
rect 324 1495 328 1499
rect 396 1495 400 1499
rect 476 1495 480 1499
rect 556 1495 560 1499
rect 636 1495 640 1499
rect 716 1495 720 1499
rect 796 1495 800 1499
rect 876 1495 880 1499
rect 956 1495 960 1499
rect 1036 1495 1040 1499
rect 1124 1495 1128 1499
rect 300 1475 304 1479
rect 364 1475 368 1479
rect 436 1475 440 1479
rect 516 1475 520 1479
rect 596 1475 600 1479
rect 676 1475 680 1479
rect 756 1475 760 1479
rect 836 1477 840 1481
rect 1388 1479 1392 1483
rect 1444 1481 1448 1485
rect 1500 1481 1504 1485
rect 1572 1479 1576 1483
rect 1652 1479 1656 1483
rect 1732 1481 1736 1485
rect 1812 1479 1816 1483
rect 1892 1479 1896 1483
rect 1972 1479 1976 1483
rect 2052 1479 2056 1483
rect 2140 1481 2144 1485
rect 916 1475 920 1479
rect 996 1475 1000 1479
rect 1076 1475 1080 1479
rect 1164 1475 1168 1479
rect 228 1419 232 1423
rect 292 1419 296 1423
rect 364 1419 368 1423
rect 444 1419 448 1423
rect 540 1419 544 1423
rect 644 1419 648 1423
rect 748 1419 752 1423
rect 852 1419 856 1423
rect 956 1419 960 1423
rect 1060 1419 1064 1423
rect 1164 1419 1168 1423
rect 1260 1419 1264 1423
rect 1396 1419 1400 1423
rect 1484 1419 1488 1423
rect 1572 1419 1576 1423
rect 1668 1419 1672 1423
rect 1764 1419 1768 1423
rect 1852 1419 1856 1423
rect 1940 1419 1944 1423
rect 2028 1419 2032 1423
rect 2108 1419 2112 1423
rect 2196 1419 2200 1423
rect 2284 1419 2288 1423
rect 188 1401 192 1405
rect 252 1399 256 1403
rect 324 1401 328 1405
rect 404 1401 408 1405
rect 500 1399 504 1403
rect 604 1401 608 1405
rect 708 1399 712 1403
rect 812 1399 816 1403
rect 916 1401 920 1405
rect 1020 1399 1024 1403
rect 1124 1399 1128 1403
rect 1220 1399 1224 1403
rect 1356 1401 1360 1405
rect 1444 1399 1448 1403
rect 1532 1399 1536 1403
rect 1628 1401 1632 1405
rect 1724 1399 1728 1403
rect 1812 1399 1816 1403
rect 1900 1399 1904 1403
rect 1988 1399 1992 1403
rect 2068 1399 2072 1403
rect 2156 1399 2160 1403
rect 2244 1399 2248 1403
rect 132 1385 136 1389
rect 204 1383 208 1387
rect 276 1385 280 1389
rect 1548 1387 1552 1391
rect 1628 1387 1632 1391
rect 1716 1387 1720 1391
rect 1812 1387 1816 1391
rect 1900 1387 1904 1391
rect 1988 1387 1992 1391
rect 2076 1387 2080 1391
rect 2156 1387 2160 1391
rect 2228 1387 2232 1391
rect 2300 1387 2304 1391
rect 2380 1387 2384 1391
rect 2436 1387 2440 1391
rect 328 1383 332 1387
rect 340 1383 344 1387
rect 412 1383 416 1387
rect 484 1383 488 1387
rect 564 1383 568 1387
rect 644 1383 648 1387
rect 732 1383 736 1387
rect 820 1383 824 1387
rect 908 1383 912 1387
rect 996 1383 1000 1387
rect 1084 1383 1088 1387
rect 1180 1383 1184 1387
rect 172 1363 176 1367
rect 244 1363 248 1367
rect 316 1363 320 1367
rect 328 1363 332 1367
rect 380 1363 384 1367
rect 452 1363 456 1367
rect 524 1363 528 1367
rect 604 1363 608 1367
rect 684 1363 688 1367
rect 772 1363 776 1367
rect 860 1363 864 1367
rect 948 1363 952 1367
rect 1036 1365 1040 1369
rect 1124 1365 1128 1369
rect 1220 1365 1224 1369
rect 1588 1367 1592 1371
rect 1668 1367 1672 1371
rect 1756 1367 1760 1371
rect 1852 1369 1856 1373
rect 1940 1369 1944 1373
rect 2028 1367 2032 1371
rect 2116 1367 2120 1371
rect 2196 1367 2200 1371
rect 2268 1367 2272 1371
rect 2340 1367 2344 1371
rect 2420 1367 2424 1371
rect 2476 1367 2480 1371
rect 1620 1315 1624 1319
rect 1684 1315 1688 1319
rect 1764 1315 1768 1319
rect 1844 1315 1848 1319
rect 1932 1315 1936 1319
rect 2020 1315 2024 1319
rect 2100 1315 2104 1319
rect 2180 1315 2184 1319
rect 2260 1315 2264 1319
rect 2340 1315 2344 1319
rect 2420 1315 2424 1319
rect 2476 1315 2480 1319
rect 172 1295 176 1299
rect 276 1295 280 1299
rect 404 1295 408 1299
rect 516 1295 520 1299
rect 620 1295 624 1299
rect 724 1295 728 1299
rect 820 1295 824 1299
rect 916 1295 920 1299
rect 1012 1295 1016 1299
rect 1580 1295 1584 1299
rect 1644 1295 1648 1299
rect 1724 1295 1728 1299
rect 1804 1297 1808 1301
rect 1892 1295 1896 1299
rect 1980 1295 1984 1299
rect 2060 1297 2064 1301
rect 2140 1295 2144 1299
rect 2220 1295 2224 1299
rect 2300 1295 2304 1299
rect 2380 1295 2384 1299
rect 2436 1295 2440 1299
rect 1548 1283 1552 1287
rect 1612 1283 1616 1287
rect 1692 1283 1696 1287
rect 1780 1283 1784 1287
rect 1876 1283 1880 1287
rect 1972 1283 1976 1287
rect 2076 1283 2080 1287
rect 2188 1283 2192 1287
rect 2300 1283 2304 1287
rect 132 1277 136 1281
rect 236 1275 240 1279
rect 364 1275 368 1279
rect 476 1275 480 1279
rect 580 1275 584 1279
rect 684 1275 688 1279
rect 780 1277 784 1281
rect 876 1277 880 1281
rect 972 1275 976 1279
rect 1588 1263 1592 1267
rect 1652 1265 1656 1269
rect 1732 1263 1736 1267
rect 1820 1263 1824 1267
rect 1916 1265 1920 1269
rect 2012 1263 2016 1267
rect 2116 1263 2120 1267
rect 2228 1265 2232 1269
rect 2340 1265 2344 1269
rect 132 1255 136 1259
rect 184 1255 188 1259
rect 196 1255 200 1259
rect 284 1255 288 1259
rect 372 1255 376 1259
rect 452 1255 456 1259
rect 532 1255 536 1259
rect 604 1255 608 1259
rect 676 1255 680 1259
rect 748 1255 752 1259
rect 820 1255 824 1259
rect 900 1255 904 1259
rect 172 1235 176 1239
rect 184 1235 188 1239
rect 236 1235 240 1239
rect 324 1235 328 1239
rect 412 1235 416 1239
rect 492 1235 496 1239
rect 572 1235 576 1239
rect 644 1235 648 1239
rect 716 1237 720 1241
rect 788 1235 792 1239
rect 860 1235 864 1239
rect 940 1237 944 1241
rect 1556 1207 1560 1211
rect 1612 1207 1616 1211
rect 1668 1207 1672 1211
rect 1724 1207 1728 1211
rect 1780 1207 1784 1211
rect 1836 1207 1840 1211
rect 1892 1207 1896 1211
rect 1948 1207 1952 1211
rect 2004 1207 2008 1211
rect 2068 1207 2072 1211
rect 2140 1207 2144 1211
rect 2220 1207 2224 1211
rect 2308 1207 2312 1211
rect 2404 1207 2408 1211
rect 2476 1207 2480 1211
rect 1516 1187 1520 1191
rect 1572 1187 1576 1191
rect 1628 1189 1632 1193
rect 1684 1187 1688 1191
rect 1740 1187 1744 1191
rect 1796 1187 1800 1191
rect 1852 1187 1856 1191
rect 1908 1187 1912 1191
rect 1964 1187 1968 1191
rect 2028 1187 2032 1191
rect 2100 1187 2104 1191
rect 2180 1187 2184 1191
rect 2268 1187 2272 1191
rect 2364 1187 2368 1191
rect 2436 1187 2440 1191
rect 172 1179 176 1183
rect 228 1179 232 1183
rect 308 1179 312 1183
rect 388 1179 392 1183
rect 468 1179 472 1183
rect 548 1179 552 1183
rect 620 1179 624 1183
rect 684 1179 688 1183
rect 756 1179 760 1183
rect 828 1179 832 1183
rect 900 1179 904 1183
rect 1548 1171 1552 1175
rect 1612 1171 1616 1175
rect 1684 1171 1688 1175
rect 1772 1171 1776 1175
rect 1884 1171 1888 1175
rect 2012 1171 2016 1175
rect 2156 1171 2160 1175
rect 2308 1171 2312 1175
rect 2436 1171 2440 1175
rect 132 1161 136 1165
rect 188 1159 192 1163
rect 268 1159 272 1163
rect 348 1159 352 1163
rect 428 1161 432 1165
rect 508 1159 512 1163
rect 580 1159 584 1163
rect 644 1159 648 1163
rect 716 1159 720 1163
rect 788 1159 792 1163
rect 860 1159 864 1163
rect 1588 1151 1592 1155
rect 1652 1151 1656 1155
rect 1724 1151 1728 1155
rect 1812 1151 1816 1155
rect 1924 1151 1928 1155
rect 2052 1153 2056 1157
rect 2196 1153 2200 1157
rect 2348 1153 2352 1157
rect 2476 1151 2480 1155
rect 164 1143 168 1147
rect 260 1143 264 1147
rect 356 1143 360 1147
rect 452 1143 456 1147
rect 548 1143 552 1147
rect 636 1145 640 1149
rect 716 1143 720 1147
rect 788 1143 792 1147
rect 860 1143 864 1147
rect 940 1143 944 1147
rect 1020 1143 1024 1147
rect 204 1123 208 1127
rect 300 1125 304 1129
rect 396 1125 400 1129
rect 492 1123 496 1127
rect 588 1125 592 1129
rect 676 1125 680 1129
rect 756 1123 760 1127
rect 828 1123 832 1127
rect 900 1123 904 1127
rect 980 1123 984 1127
rect 1060 1123 1064 1127
rect 1420 1099 1424 1103
rect 1484 1099 1488 1103
rect 1556 1099 1560 1103
rect 1628 1099 1632 1103
rect 1708 1099 1712 1103
rect 1788 1099 1792 1103
rect 1868 1099 1872 1103
rect 1948 1099 1952 1103
rect 2020 1099 2024 1103
rect 2092 1099 2096 1103
rect 2172 1099 2176 1103
rect 2252 1099 2256 1103
rect 1380 1079 1384 1083
rect 1444 1079 1448 1083
rect 1516 1079 1520 1083
rect 1588 1079 1592 1083
rect 1668 1079 1672 1083
rect 1748 1079 1752 1083
rect 1828 1081 1832 1085
rect 1908 1079 1912 1083
rect 1980 1079 1984 1083
rect 2052 1079 2056 1083
rect 2132 1079 2136 1083
rect 2212 1079 2216 1083
rect 244 1063 248 1067
rect 316 1063 320 1067
rect 396 1063 400 1067
rect 484 1063 488 1067
rect 580 1063 584 1067
rect 676 1063 680 1067
rect 764 1063 768 1067
rect 852 1063 856 1067
rect 932 1063 936 1067
rect 1012 1063 1016 1067
rect 1092 1063 1096 1067
rect 1180 1063 1184 1067
rect 1348 1059 1352 1063
rect 1436 1059 1440 1063
rect 1556 1059 1560 1063
rect 1676 1059 1680 1063
rect 1796 1059 1800 1063
rect 1908 1061 1912 1065
rect 2020 1059 2024 1063
rect 2132 1059 2136 1063
rect 2236 1059 2240 1063
rect 2348 1059 2352 1063
rect 2436 1059 2440 1063
rect 204 1043 208 1047
rect 276 1043 280 1047
rect 356 1043 360 1047
rect 444 1043 448 1047
rect 540 1045 544 1049
rect 636 1043 640 1047
rect 724 1045 728 1049
rect 812 1043 816 1047
rect 892 1043 896 1047
rect 972 1043 976 1047
rect 1052 1043 1056 1047
rect 1140 1043 1144 1047
rect 1388 1039 1392 1043
rect 1476 1039 1480 1043
rect 1596 1039 1600 1043
rect 1716 1039 1720 1043
rect 1836 1039 1840 1043
rect 1948 1039 1952 1043
rect 2060 1039 2064 1043
rect 2172 1039 2176 1043
rect 2276 1039 2280 1043
rect 2388 1039 2392 1043
rect 2476 1039 2480 1043
rect 276 1023 280 1027
rect 364 1023 368 1027
rect 460 1023 464 1027
rect 556 1023 560 1027
rect 652 1023 656 1027
rect 748 1025 752 1029
rect 836 1023 840 1027
rect 924 1023 928 1027
rect 1004 1023 1008 1027
rect 1084 1023 1088 1027
rect 1136 1023 1140 1027
rect 1164 1023 1168 1027
rect 1220 1023 1224 1027
rect 316 1003 320 1007
rect 404 1005 408 1009
rect 500 1005 504 1009
rect 596 1003 600 1007
rect 692 1005 696 1009
rect 788 1003 792 1007
rect 876 1003 880 1007
rect 964 1003 968 1007
rect 1044 1005 1048 1009
rect 1124 1003 1128 1007
rect 1136 1003 1140 1007
rect 1204 1003 1208 1007
rect 1260 1003 1264 1007
rect 1388 983 1392 987
rect 1548 983 1552 987
rect 1716 983 1720 987
rect 1860 983 1864 987
rect 1988 983 1992 987
rect 2108 983 2112 987
rect 2212 983 2216 987
rect 2308 983 2312 987
rect 2404 983 2408 987
rect 2476 983 2480 987
rect 1348 963 1352 967
rect 1508 965 1512 969
rect 1676 963 1680 967
rect 1820 963 1824 967
rect 1948 963 1952 967
rect 2068 963 2072 967
rect 2172 963 2176 967
rect 2268 963 2272 967
rect 2364 963 2368 967
rect 2436 963 2440 967
rect 308 951 312 955
rect 396 951 400 955
rect 492 951 496 955
rect 588 951 592 955
rect 692 951 696 955
rect 788 951 792 955
rect 876 951 880 955
rect 964 951 968 955
rect 1044 951 1048 955
rect 1124 951 1128 955
rect 1204 951 1208 955
rect 1260 953 1264 957
rect 1348 939 1352 943
rect 1404 939 1408 943
rect 1484 939 1488 943
rect 1588 939 1592 943
rect 1700 939 1704 943
rect 1812 939 1816 943
rect 1916 939 1920 943
rect 2012 939 2016 943
rect 2108 939 2112 943
rect 2196 939 2200 943
rect 2276 939 2280 943
rect 2356 939 2360 943
rect 2436 939 2440 943
rect 268 931 272 935
rect 356 931 360 935
rect 452 931 456 935
rect 548 931 552 935
rect 652 931 656 935
rect 748 933 752 937
rect 836 931 840 935
rect 924 931 928 935
rect 1004 931 1008 935
rect 1084 933 1088 937
rect 1164 931 1168 935
rect 1220 931 1224 935
rect 1388 919 1392 923
rect 1444 919 1448 923
rect 1524 919 1528 923
rect 1628 919 1632 923
rect 1740 919 1744 923
rect 1852 921 1856 925
rect 1956 919 1960 923
rect 2052 919 2056 923
rect 2148 919 2152 923
rect 2236 921 2240 925
rect 2316 921 2320 925
rect 2396 921 2400 925
rect 2476 919 2480 923
rect 252 911 256 915
rect 324 911 328 915
rect 404 913 408 917
rect 500 911 504 915
rect 596 911 600 915
rect 692 911 696 915
rect 788 911 792 915
rect 884 911 888 915
rect 972 911 976 915
rect 1068 911 1072 915
rect 1120 911 1124 915
rect 1164 911 1168 915
rect 292 891 296 895
rect 364 893 368 897
rect 444 891 448 895
rect 540 891 544 895
rect 636 891 640 895
rect 732 891 736 895
rect 828 891 832 895
rect 924 891 928 895
rect 1012 891 1016 895
rect 1108 891 1112 895
rect 1120 891 1124 895
rect 1204 891 1208 895
rect 1468 863 1472 867
rect 1524 863 1528 867
rect 1588 863 1592 867
rect 1660 863 1664 867
rect 1740 863 1744 867
rect 1828 863 1832 867
rect 1932 863 1936 867
rect 2052 863 2056 867
rect 2180 863 2184 867
rect 2316 863 2320 867
rect 2460 863 2464 867
rect 1428 843 1432 847
rect 1484 843 1488 847
rect 1548 843 1552 847
rect 1620 843 1624 847
rect 1700 843 1704 847
rect 1788 845 1792 849
rect 1892 843 1896 847
rect 2012 845 2016 849
rect 2140 843 2144 847
rect 2276 843 2280 847
rect 2420 843 2424 847
rect 284 835 288 839
rect 348 835 352 839
rect 412 835 416 839
rect 476 835 480 839
rect 540 835 544 839
rect 604 835 608 839
rect 668 835 672 839
rect 732 835 736 839
rect 796 835 800 839
rect 868 835 872 839
rect 940 835 944 839
rect 1572 829 1576 833
rect 1628 827 1632 831
rect 1684 827 1688 831
rect 1748 827 1752 831
rect 1808 827 1812 831
rect 1828 827 1832 831
rect 1908 827 1912 831
rect 1996 827 2000 831
rect 2084 827 2088 831
rect 2172 827 2176 831
rect 2268 827 2272 831
rect 2364 827 2368 831
rect 2436 827 2440 831
rect 244 817 248 821
rect 308 815 312 819
rect 372 817 376 821
rect 436 815 440 819
rect 500 815 504 819
rect 564 815 568 819
rect 628 815 632 819
rect 692 815 696 819
rect 756 815 760 819
rect 828 815 832 819
rect 900 815 904 819
rect 1612 807 1616 811
rect 1668 807 1672 811
rect 1724 807 1728 811
rect 1788 807 1792 811
rect 1808 807 1812 811
rect 1868 807 1872 811
rect 1948 807 1952 811
rect 2036 807 2040 811
rect 2124 807 2128 811
rect 2212 807 2216 811
rect 2308 807 2312 811
rect 2404 807 2408 811
rect 2476 807 2480 811
rect 196 799 200 803
rect 284 799 288 803
rect 372 801 376 805
rect 460 799 464 803
rect 540 799 544 803
rect 612 799 616 803
rect 684 799 688 803
rect 748 799 752 803
rect 812 799 816 803
rect 876 799 880 803
rect 948 799 952 803
rect 1020 799 1024 803
rect 236 779 240 783
rect 324 779 328 783
rect 412 779 416 783
rect 500 779 504 783
rect 580 779 584 783
rect 652 779 656 783
rect 724 781 728 785
rect 788 779 792 783
rect 852 781 856 785
rect 916 781 920 785
rect 988 781 992 785
rect 1060 781 1064 785
rect 1604 751 1608 755
rect 1660 751 1664 755
rect 1724 751 1728 755
rect 1796 751 1800 755
rect 1868 751 1872 755
rect 1956 751 1960 755
rect 2052 751 2056 755
rect 2156 751 2160 755
rect 2268 751 2272 755
rect 2380 751 2384 755
rect 2476 751 2480 755
rect 1564 731 1568 735
rect 1620 731 1624 735
rect 1684 731 1688 735
rect 1756 733 1760 737
rect 1828 731 1832 735
rect 1916 733 1920 737
rect 2012 731 2016 735
rect 2116 731 2120 735
rect 2228 731 2232 735
rect 2340 731 2344 735
rect 2436 731 2440 735
rect 172 727 176 731
rect 292 727 296 731
rect 428 727 432 731
rect 556 727 560 731
rect 684 727 688 731
rect 812 727 816 731
rect 940 727 944 731
rect 1076 727 1080 731
rect 1348 719 1352 723
rect 1412 719 1416 723
rect 1508 719 1512 723
rect 1612 719 1616 723
rect 1716 719 1720 723
rect 1820 719 1824 723
rect 1924 719 1928 723
rect 2028 719 2032 723
rect 2132 719 2136 723
rect 2236 719 2240 723
rect 2348 719 2352 723
rect 2436 719 2440 723
rect 132 709 136 713
rect 252 709 256 713
rect 388 707 392 711
rect 516 709 520 713
rect 644 707 648 711
rect 772 707 776 711
rect 900 707 904 711
rect 1036 707 1040 711
rect 1388 701 1392 705
rect 1452 701 1456 705
rect 1548 701 1552 705
rect 132 695 136 699
rect 188 695 192 699
rect 276 695 280 699
rect 344 695 348 699
rect 372 695 376 699
rect 484 695 488 699
rect 604 695 608 699
rect 724 695 728 699
rect 852 695 856 699
rect 980 695 984 699
rect 1108 697 1112 701
rect 1652 699 1656 703
rect 1756 701 1760 705
rect 1860 699 1864 703
rect 1964 699 1968 703
rect 2068 699 2072 703
rect 2172 699 2176 703
rect 2276 699 2280 703
rect 2388 699 2392 703
rect 2476 699 2480 703
rect 1220 695 1224 699
rect 172 675 176 679
rect 228 675 232 679
rect 316 675 320 679
rect 344 675 348 679
rect 412 675 416 679
rect 524 677 528 681
rect 644 675 648 679
rect 764 677 768 681
rect 892 675 896 679
rect 1020 677 1024 681
rect 1148 675 1152 679
rect 1260 675 1264 679
rect 1388 635 1392 639
rect 1452 635 1456 639
rect 1548 635 1552 639
rect 1644 635 1648 639
rect 1748 635 1752 639
rect 1860 635 1864 639
rect 1972 635 1976 639
rect 2092 635 2096 639
rect 2220 635 2224 639
rect 2356 635 2360 639
rect 2476 635 2480 639
rect 188 619 192 623
rect 300 619 304 623
rect 404 619 408 623
rect 500 619 504 623
rect 596 619 600 623
rect 692 619 696 623
rect 788 619 792 623
rect 884 619 888 623
rect 980 619 984 623
rect 1076 619 1080 623
rect 1180 619 1184 623
rect 1260 619 1264 623
rect 1348 615 1352 619
rect 1412 615 1416 619
rect 1508 615 1512 619
rect 1604 617 1608 621
rect 1708 615 1712 619
rect 1820 617 1824 621
rect 1932 615 1936 619
rect 2052 615 2056 619
rect 2180 615 2184 619
rect 2316 615 2320 619
rect 2436 615 2440 619
rect 148 599 152 603
rect 260 599 264 603
rect 364 599 368 603
rect 460 601 464 605
rect 556 601 560 605
rect 652 599 656 603
rect 748 599 752 603
rect 844 599 848 603
rect 940 599 944 603
rect 1036 601 1040 605
rect 1364 603 1368 607
rect 1444 605 1448 609
rect 1532 603 1536 607
rect 1628 603 1632 607
rect 1696 603 1700 607
rect 1724 603 1728 607
rect 1828 603 1832 607
rect 1940 603 1944 607
rect 2060 603 2064 607
rect 2188 603 2192 607
rect 2324 603 2328 607
rect 2436 603 2440 607
rect 1140 599 1144 603
rect 1220 599 1224 603
rect 132 587 136 591
rect 220 587 224 591
rect 316 587 320 591
rect 412 587 416 591
rect 516 587 520 591
rect 612 587 616 591
rect 708 587 712 591
rect 804 587 808 591
rect 892 589 896 593
rect 980 587 984 591
rect 1068 587 1072 591
rect 1164 587 1168 591
rect 1404 583 1408 587
rect 1484 585 1488 589
rect 1572 583 1576 587
rect 1668 583 1672 587
rect 1696 583 1700 587
rect 1764 583 1768 587
rect 1868 583 1872 587
rect 1980 583 1984 587
rect 2100 585 2104 589
rect 2228 583 2232 587
rect 2364 585 2368 589
rect 2476 583 2480 587
rect 172 567 176 571
rect 260 569 264 573
rect 356 569 360 573
rect 452 567 456 571
rect 556 567 560 571
rect 652 567 656 571
rect 748 567 752 571
rect 844 567 848 571
rect 932 567 936 571
rect 1020 567 1024 571
rect 1108 569 1112 573
rect 1204 569 1208 573
rect 1412 531 1416 535
rect 1492 531 1496 535
rect 1588 531 1592 535
rect 1684 531 1688 535
rect 1788 531 1792 535
rect 1892 531 1896 535
rect 1996 531 2000 535
rect 2092 531 2096 535
rect 2188 531 2192 535
rect 2292 531 2296 535
rect 2396 531 2400 535
rect 2476 531 2480 535
rect 1372 511 1376 515
rect 1452 511 1456 515
rect 1548 513 1552 517
rect 1644 513 1648 517
rect 1748 511 1752 515
rect 1852 513 1856 517
rect 1956 511 1960 515
rect 2052 513 2056 517
rect 2148 511 2152 515
rect 2252 511 2256 515
rect 2356 511 2360 515
rect 2436 511 2440 515
rect 180 507 184 511
rect 276 507 280 511
rect 372 507 376 511
rect 468 507 472 511
rect 564 507 568 511
rect 660 507 664 511
rect 748 507 752 511
rect 828 507 832 511
rect 908 507 912 511
rect 988 507 992 511
rect 1068 507 1072 511
rect 1348 495 1352 499
rect 1436 495 1440 499
rect 1556 495 1560 499
rect 1676 495 1680 499
rect 1788 495 1792 499
rect 1900 495 1904 499
rect 2004 495 2008 499
rect 2100 495 2104 499
rect 2188 497 2192 501
rect 2276 495 2280 499
rect 2364 495 2368 499
rect 2436 495 2440 499
rect 140 487 144 491
rect 236 487 240 491
rect 332 489 336 493
rect 428 487 432 491
rect 524 489 528 493
rect 620 487 624 491
rect 708 487 712 491
rect 788 489 792 493
rect 868 489 872 493
rect 948 487 952 491
rect 1028 487 1032 491
rect 1388 477 1392 481
rect 1476 477 1480 481
rect 132 471 136 475
rect 188 471 192 475
rect 268 473 272 477
rect 356 471 360 475
rect 444 471 448 475
rect 540 471 544 475
rect 636 471 640 475
rect 732 471 736 475
rect 828 471 832 475
rect 932 471 936 475
rect 1036 471 1040 475
rect 1140 471 1144 475
rect 1220 473 1224 477
rect 1596 475 1600 479
rect 1716 475 1720 479
rect 1828 475 1832 479
rect 1940 475 1944 479
rect 2044 475 2048 479
rect 2140 475 2144 479
rect 2228 477 2232 481
rect 2316 475 2320 479
rect 2404 475 2408 479
rect 2476 477 2480 481
rect 172 451 176 455
rect 228 453 232 457
rect 308 451 312 455
rect 396 451 400 455
rect 484 451 488 455
rect 580 451 584 455
rect 676 451 680 455
rect 772 453 776 457
rect 868 451 872 455
rect 972 451 976 455
rect 1076 453 1080 457
rect 1180 451 1184 455
rect 1260 453 1264 457
rect 1620 411 1624 415
rect 1676 411 1680 415
rect 1732 411 1736 415
rect 1796 411 1800 415
rect 1868 411 1872 415
rect 1948 411 1952 415
rect 2028 411 2032 415
rect 2116 411 2120 415
rect 2212 411 2216 415
rect 2308 411 2312 415
rect 2404 411 2408 415
rect 2476 411 2480 415
rect 172 399 176 403
rect 228 399 232 403
rect 316 399 320 403
rect 420 399 424 403
rect 532 399 536 403
rect 644 399 648 403
rect 756 399 760 403
rect 868 399 872 403
rect 972 399 976 403
rect 1076 399 1080 403
rect 1180 399 1184 403
rect 1260 399 1264 403
rect 1580 393 1584 397
rect 1636 393 1640 397
rect 1692 393 1696 397
rect 1756 393 1760 397
rect 1828 391 1832 395
rect 1908 391 1912 395
rect 1988 391 1992 395
rect 2076 391 2080 395
rect 2172 391 2176 395
rect 2268 391 2272 395
rect 2364 391 2368 395
rect 2436 391 2440 395
rect 132 379 136 383
rect 188 379 192 383
rect 276 379 280 383
rect 380 379 384 383
rect 492 379 496 383
rect 604 379 608 383
rect 716 379 720 383
rect 828 379 832 383
rect 932 379 936 383
rect 1036 381 1040 385
rect 1140 379 1144 383
rect 1220 379 1224 383
rect 1660 375 1664 379
rect 1716 375 1720 379
rect 1780 375 1784 379
rect 1852 375 1856 379
rect 1924 375 1928 379
rect 2004 375 2008 379
rect 2092 375 2096 379
rect 2180 375 2184 379
rect 2268 375 2272 379
rect 2356 375 2360 379
rect 2436 375 2440 379
rect 132 363 136 367
rect 212 363 216 367
rect 316 365 320 369
rect 420 363 424 367
rect 524 363 528 367
rect 628 363 632 367
rect 732 363 736 367
rect 828 363 832 367
rect 916 363 920 367
rect 996 363 1000 367
rect 1076 363 1080 367
rect 1156 363 1160 367
rect 1220 363 1224 367
rect 1700 355 1704 359
rect 1756 355 1760 359
rect 1820 355 1824 359
rect 1892 355 1896 359
rect 1964 355 1968 359
rect 2044 357 2048 361
rect 2132 357 2136 361
rect 2220 355 2224 359
rect 2308 357 2312 361
rect 2396 355 2400 359
rect 2476 357 2480 361
rect 172 343 176 347
rect 252 345 256 349
rect 356 343 360 347
rect 460 343 464 347
rect 564 343 568 347
rect 668 343 672 347
rect 772 343 776 347
rect 868 343 872 347
rect 956 343 960 347
rect 1036 345 1040 349
rect 1116 343 1120 347
rect 1196 343 1200 347
rect 1260 343 1264 347
rect 1388 295 1392 299
rect 1492 295 1496 299
rect 1620 295 1624 299
rect 1748 295 1752 299
rect 1876 295 1880 299
rect 1988 295 1992 299
rect 2100 295 2104 299
rect 2204 295 2208 299
rect 2300 295 2304 299
rect 2396 295 2400 299
rect 2476 295 2480 299
rect 172 287 176 291
rect 252 287 256 291
rect 356 287 360 291
rect 460 287 464 291
rect 572 287 576 291
rect 676 287 680 291
rect 780 287 784 291
rect 884 287 888 291
rect 980 287 984 291
rect 1076 287 1080 291
rect 1180 287 1184 291
rect 1260 287 1264 291
rect 1348 277 1352 281
rect 1452 277 1456 281
rect 1580 275 1584 279
rect 1708 275 1712 279
rect 1836 277 1840 281
rect 1948 275 1952 279
rect 2060 277 2064 281
rect 2164 275 2168 279
rect 2260 277 2264 281
rect 2356 275 2360 279
rect 2436 275 2440 279
rect 132 267 136 271
rect 212 267 216 271
rect 316 269 320 273
rect 420 269 424 273
rect 532 267 536 271
rect 636 269 640 273
rect 740 269 744 273
rect 844 267 848 271
rect 940 267 944 271
rect 1036 267 1040 271
rect 1140 267 1144 271
rect 1220 267 1224 271
rect 132 255 136 259
rect 204 255 208 259
rect 300 255 304 259
rect 404 255 408 259
rect 516 255 520 259
rect 628 255 632 259
rect 740 255 744 259
rect 852 255 856 259
rect 964 255 968 259
rect 1084 255 1088 259
rect 1204 255 1208 259
rect 1348 255 1352 259
rect 1428 255 1432 259
rect 1532 255 1536 259
rect 1636 255 1640 259
rect 1740 255 1744 259
rect 1844 255 1848 259
rect 1948 255 1952 259
rect 2052 255 2056 259
rect 2156 255 2160 259
rect 2252 255 2256 259
rect 2356 255 2360 259
rect 2436 255 2440 259
rect 172 235 176 239
rect 244 237 248 241
rect 340 237 344 241
rect 444 235 448 239
rect 556 235 560 239
rect 668 235 672 239
rect 780 235 784 239
rect 892 235 896 239
rect 1004 235 1008 239
rect 1124 237 1128 241
rect 1244 237 1248 241
rect 1388 235 1392 239
rect 1468 235 1472 239
rect 1572 235 1576 239
rect 1676 235 1680 239
rect 1780 235 1784 239
rect 1884 235 1888 239
rect 1988 235 1992 239
rect 2092 235 2096 239
rect 2196 235 2200 239
rect 2292 235 2296 239
rect 2396 235 2400 239
rect 2476 235 2480 239
rect 220 179 224 183
rect 316 179 320 183
rect 420 179 424 183
rect 524 179 528 183
rect 628 179 632 183
rect 732 179 736 183
rect 836 179 840 183
rect 932 179 936 183
rect 1036 179 1040 183
rect 1140 179 1144 183
rect 1388 179 1392 183
rect 1444 179 1448 183
rect 1508 179 1512 183
rect 1588 179 1592 183
rect 1676 179 1680 183
rect 1756 179 1760 183
rect 1844 179 1848 183
rect 1932 179 1936 183
rect 2028 179 2032 183
rect 2140 179 2144 183
rect 2252 179 2256 183
rect 2372 179 2376 183
rect 2476 179 2480 183
rect 180 159 184 163
rect 276 159 280 163
rect 380 161 384 165
rect 484 161 488 165
rect 588 159 592 163
rect 692 161 696 165
rect 796 159 800 163
rect 892 159 896 163
rect 996 159 1000 163
rect 1100 159 1104 163
rect 1348 161 1352 165
rect 1404 161 1408 165
rect 1468 159 1472 163
rect 1548 161 1552 165
rect 1636 161 1640 165
rect 1716 159 1720 163
rect 1804 161 1808 165
rect 1892 161 1896 165
rect 1988 159 1992 163
rect 2100 161 2104 165
rect 2212 161 2216 165
rect 2332 159 2336 163
rect 2436 159 2440 163
rect 132 139 136 143
rect 188 139 192 143
rect 244 139 248 143
rect 300 139 304 143
rect 356 139 360 143
rect 412 139 416 143
rect 468 139 472 143
rect 524 139 528 143
rect 580 139 584 143
rect 636 139 640 143
rect 692 139 696 143
rect 748 139 752 143
rect 812 139 816 143
rect 876 139 880 143
rect 940 139 944 143
rect 1004 139 1008 143
rect 1068 139 1072 143
rect 1132 139 1136 143
rect 1348 127 1352 131
rect 1404 127 1408 131
rect 1460 127 1464 131
rect 1516 127 1520 131
rect 1572 127 1576 131
rect 1628 127 1632 131
rect 1684 127 1688 131
rect 1740 127 1744 131
rect 1804 127 1808 131
rect 1860 127 1864 131
rect 1924 127 1928 131
rect 1988 127 1992 131
rect 2052 127 2056 131
rect 2124 127 2128 131
rect 2204 127 2208 131
rect 2284 127 2288 131
rect 2372 127 2376 131
rect 2436 127 2440 131
rect 172 119 176 123
rect 228 119 232 123
rect 284 121 288 125
rect 340 121 344 125
rect 396 121 400 125
rect 452 121 456 125
rect 508 119 512 123
rect 564 119 568 123
rect 620 121 624 125
rect 676 119 680 123
rect 732 119 736 123
rect 788 119 792 123
rect 852 121 856 125
rect 916 121 920 125
rect 980 121 984 125
rect 1044 121 1048 125
rect 1108 121 1112 125
rect 1172 121 1176 125
rect 1388 107 1392 111
rect 1444 107 1448 111
rect 1500 107 1504 111
rect 1556 107 1560 111
rect 1612 107 1616 111
rect 1668 107 1672 111
rect 1724 107 1728 111
rect 1780 107 1784 111
rect 1844 107 1848 111
rect 1900 107 1904 111
rect 1964 107 1968 111
rect 2028 109 2032 113
rect 2092 109 2096 113
rect 2164 107 2168 111
rect 2244 107 2248 111
rect 2324 109 2328 113
rect 2476 109 2480 113
<< m2 >>
rect 134 2576 140 2577
rect 110 2573 116 2574
rect 110 2569 111 2573
rect 115 2569 116 2573
rect 134 2572 135 2576
rect 139 2572 140 2576
rect 134 2571 140 2572
rect 190 2576 196 2577
rect 190 2572 191 2576
rect 195 2572 196 2576
rect 190 2571 196 2572
rect 246 2576 252 2577
rect 246 2572 247 2576
rect 251 2572 252 2576
rect 246 2571 252 2572
rect 302 2576 308 2577
rect 302 2572 303 2576
rect 307 2572 308 2576
rect 302 2571 308 2572
rect 358 2576 364 2577
rect 358 2572 359 2576
rect 363 2572 364 2576
rect 358 2571 364 2572
rect 1286 2573 1292 2574
rect 110 2568 116 2569
rect 1286 2569 1287 2573
rect 1291 2569 1292 2573
rect 1286 2568 1292 2569
rect 110 2556 116 2557
rect 1286 2556 1292 2557
rect 110 2552 111 2556
rect 115 2552 116 2556
rect 110 2551 116 2552
rect 150 2555 156 2556
rect 150 2551 151 2555
rect 155 2551 156 2555
rect 150 2550 156 2551
rect 171 2555 177 2556
rect 171 2551 172 2555
rect 176 2554 177 2555
rect 186 2555 192 2556
rect 186 2554 187 2555
rect 176 2552 187 2554
rect 176 2551 177 2552
rect 171 2550 177 2551
rect 186 2551 187 2552
rect 191 2551 192 2555
rect 186 2550 192 2551
rect 206 2555 212 2556
rect 206 2551 207 2555
rect 211 2551 212 2555
rect 206 2550 212 2551
rect 227 2555 233 2556
rect 227 2551 228 2555
rect 232 2554 233 2555
rect 242 2555 248 2556
rect 242 2554 243 2555
rect 232 2552 243 2554
rect 232 2551 233 2552
rect 227 2550 233 2551
rect 242 2551 243 2552
rect 247 2551 248 2555
rect 242 2550 248 2551
rect 262 2555 268 2556
rect 262 2551 263 2555
rect 267 2551 268 2555
rect 262 2550 268 2551
rect 283 2555 289 2556
rect 283 2551 284 2555
rect 288 2554 289 2555
rect 298 2555 304 2556
rect 298 2554 299 2555
rect 288 2552 299 2554
rect 288 2551 289 2552
rect 283 2550 289 2551
rect 298 2551 299 2552
rect 303 2551 304 2555
rect 298 2550 304 2551
rect 318 2555 324 2556
rect 318 2551 319 2555
rect 323 2551 324 2555
rect 318 2550 324 2551
rect 339 2555 345 2556
rect 339 2551 340 2555
rect 344 2554 345 2555
rect 354 2555 360 2556
rect 354 2554 355 2555
rect 344 2552 355 2554
rect 344 2551 345 2552
rect 339 2550 345 2551
rect 354 2551 355 2552
rect 359 2551 360 2555
rect 354 2550 360 2551
rect 374 2555 380 2556
rect 374 2551 375 2555
rect 379 2551 380 2555
rect 374 2550 380 2551
rect 395 2555 401 2556
rect 395 2551 396 2555
rect 400 2551 401 2555
rect 1286 2552 1287 2556
rect 1291 2552 1292 2556
rect 1494 2556 1500 2557
rect 1286 2551 1292 2552
rect 1326 2553 1332 2554
rect 395 2550 401 2551
rect 214 2547 220 2548
rect 214 2543 215 2547
rect 219 2546 220 2547
rect 397 2546 399 2550
rect 1326 2549 1327 2553
rect 1331 2549 1332 2553
rect 1494 2552 1495 2556
rect 1499 2552 1500 2556
rect 1494 2551 1500 2552
rect 1550 2556 1556 2557
rect 1550 2552 1551 2556
rect 1555 2552 1556 2556
rect 1550 2551 1556 2552
rect 1606 2556 1612 2557
rect 1606 2552 1607 2556
rect 1611 2552 1612 2556
rect 1606 2551 1612 2552
rect 1662 2556 1668 2557
rect 1662 2552 1663 2556
rect 1667 2552 1668 2556
rect 1662 2551 1668 2552
rect 1718 2556 1724 2557
rect 1718 2552 1719 2556
rect 1723 2552 1724 2556
rect 1718 2551 1724 2552
rect 1774 2556 1780 2557
rect 1774 2552 1775 2556
rect 1779 2552 1780 2556
rect 1774 2551 1780 2552
rect 1830 2556 1836 2557
rect 1830 2552 1831 2556
rect 1835 2552 1836 2556
rect 1830 2551 1836 2552
rect 1886 2556 1892 2557
rect 1886 2552 1887 2556
rect 1891 2552 1892 2556
rect 1886 2551 1892 2552
rect 1942 2556 1948 2557
rect 1942 2552 1943 2556
rect 1947 2552 1948 2556
rect 1942 2551 1948 2552
rect 1998 2556 2004 2557
rect 1998 2552 1999 2556
rect 2003 2552 2004 2556
rect 1998 2551 2004 2552
rect 2054 2556 2060 2557
rect 2054 2552 2055 2556
rect 2059 2552 2060 2556
rect 2054 2551 2060 2552
rect 2110 2556 2116 2557
rect 2110 2552 2111 2556
rect 2115 2552 2116 2556
rect 2110 2551 2116 2552
rect 2166 2556 2172 2557
rect 2166 2552 2167 2556
rect 2171 2552 2172 2556
rect 2166 2551 2172 2552
rect 2502 2553 2508 2554
rect 1326 2548 1332 2549
rect 2502 2549 2503 2553
rect 2507 2549 2508 2553
rect 2502 2548 2508 2549
rect 219 2544 399 2546
rect 219 2543 220 2544
rect 214 2542 220 2543
rect 1326 2536 1332 2537
rect 2502 2536 2508 2537
rect 186 2535 193 2536
rect 186 2531 187 2535
rect 192 2531 193 2535
rect 186 2530 193 2531
rect 242 2535 249 2536
rect 242 2531 243 2535
rect 248 2531 249 2535
rect 242 2530 249 2531
rect 298 2535 305 2536
rect 298 2531 299 2535
rect 304 2531 305 2535
rect 298 2530 305 2531
rect 354 2535 361 2536
rect 354 2531 355 2535
rect 360 2531 361 2535
rect 1326 2532 1327 2536
rect 1331 2532 1332 2536
rect 1326 2531 1332 2532
rect 1510 2535 1516 2536
rect 1510 2531 1511 2535
rect 1515 2531 1516 2535
rect 354 2530 361 2531
rect 1510 2530 1516 2531
rect 1531 2535 1540 2536
rect 1531 2531 1532 2535
rect 1539 2531 1540 2535
rect 1531 2530 1540 2531
rect 1566 2535 1572 2536
rect 1566 2531 1567 2535
rect 1571 2531 1572 2535
rect 1566 2530 1572 2531
rect 1587 2535 1593 2536
rect 1587 2531 1588 2535
rect 1592 2534 1593 2535
rect 1598 2535 1604 2536
rect 1598 2534 1599 2535
rect 1592 2532 1599 2534
rect 1592 2531 1593 2532
rect 1587 2530 1593 2531
rect 1598 2531 1599 2532
rect 1603 2531 1604 2535
rect 1598 2530 1604 2531
rect 1622 2535 1628 2536
rect 1622 2531 1623 2535
rect 1627 2531 1628 2535
rect 1622 2530 1628 2531
rect 1643 2535 1649 2536
rect 1643 2531 1644 2535
rect 1648 2534 1649 2535
rect 1658 2535 1664 2536
rect 1658 2534 1659 2535
rect 1648 2532 1659 2534
rect 1648 2531 1649 2532
rect 1643 2530 1649 2531
rect 1658 2531 1659 2532
rect 1663 2531 1664 2535
rect 1658 2530 1664 2531
rect 1678 2535 1684 2536
rect 1678 2531 1679 2535
rect 1683 2531 1684 2535
rect 1678 2530 1684 2531
rect 1699 2535 1705 2536
rect 1699 2531 1700 2535
rect 1704 2534 1705 2535
rect 1714 2535 1720 2536
rect 1714 2534 1715 2535
rect 1704 2532 1715 2534
rect 1704 2531 1705 2532
rect 1699 2530 1705 2531
rect 1714 2531 1715 2532
rect 1719 2531 1720 2535
rect 1714 2530 1720 2531
rect 1734 2535 1740 2536
rect 1734 2531 1735 2535
rect 1739 2531 1740 2535
rect 1734 2530 1740 2531
rect 1755 2535 1761 2536
rect 1755 2531 1756 2535
rect 1760 2534 1761 2535
rect 1770 2535 1776 2536
rect 1770 2534 1771 2535
rect 1760 2532 1771 2534
rect 1760 2531 1761 2532
rect 1755 2530 1761 2531
rect 1770 2531 1771 2532
rect 1775 2531 1776 2535
rect 1770 2530 1776 2531
rect 1790 2535 1796 2536
rect 1790 2531 1791 2535
rect 1795 2531 1796 2535
rect 1790 2530 1796 2531
rect 1811 2535 1820 2536
rect 1811 2531 1812 2535
rect 1819 2531 1820 2535
rect 1811 2530 1820 2531
rect 1846 2535 1852 2536
rect 1846 2531 1847 2535
rect 1851 2531 1852 2535
rect 1846 2530 1852 2531
rect 1867 2535 1873 2536
rect 1867 2531 1868 2535
rect 1872 2534 1873 2535
rect 1882 2535 1888 2536
rect 1882 2534 1883 2535
rect 1872 2532 1883 2534
rect 1872 2531 1873 2532
rect 1867 2530 1873 2531
rect 1882 2531 1883 2532
rect 1887 2531 1888 2535
rect 1882 2530 1888 2531
rect 1902 2535 1908 2536
rect 1902 2531 1903 2535
rect 1907 2531 1908 2535
rect 1902 2530 1908 2531
rect 1923 2535 1929 2536
rect 1923 2531 1924 2535
rect 1928 2534 1929 2535
rect 1938 2535 1944 2536
rect 1938 2534 1939 2535
rect 1928 2532 1939 2534
rect 1928 2531 1929 2532
rect 1923 2530 1929 2531
rect 1938 2531 1939 2532
rect 1943 2531 1944 2535
rect 1938 2530 1944 2531
rect 1958 2535 1964 2536
rect 1958 2531 1959 2535
rect 1963 2531 1964 2535
rect 1958 2530 1964 2531
rect 1979 2535 1985 2536
rect 1979 2531 1980 2535
rect 1984 2534 1985 2535
rect 1994 2535 2000 2536
rect 1994 2534 1995 2535
rect 1984 2532 1995 2534
rect 1984 2531 1985 2532
rect 1979 2530 1985 2531
rect 1994 2531 1995 2532
rect 1999 2531 2000 2535
rect 1994 2530 2000 2531
rect 2014 2535 2020 2536
rect 2014 2531 2015 2535
rect 2019 2531 2020 2535
rect 2014 2530 2020 2531
rect 2035 2535 2041 2536
rect 2035 2531 2036 2535
rect 2040 2534 2041 2535
rect 2050 2535 2056 2536
rect 2050 2534 2051 2535
rect 2040 2532 2051 2534
rect 2040 2531 2041 2532
rect 2035 2530 2041 2531
rect 2050 2531 2051 2532
rect 2055 2531 2056 2535
rect 2050 2530 2056 2531
rect 2070 2535 2076 2536
rect 2070 2531 2071 2535
rect 2075 2531 2076 2535
rect 2070 2530 2076 2531
rect 2091 2535 2097 2536
rect 2091 2531 2092 2535
rect 2096 2534 2097 2535
rect 2102 2535 2108 2536
rect 2102 2534 2103 2535
rect 2096 2532 2103 2534
rect 2096 2531 2097 2532
rect 2091 2530 2097 2531
rect 2102 2531 2103 2532
rect 2107 2531 2108 2535
rect 2102 2530 2108 2531
rect 2126 2535 2132 2536
rect 2126 2531 2127 2535
rect 2131 2531 2132 2535
rect 2126 2530 2132 2531
rect 2147 2535 2153 2536
rect 2147 2531 2148 2535
rect 2152 2534 2153 2535
rect 2162 2535 2168 2536
rect 2162 2534 2163 2535
rect 2152 2532 2163 2534
rect 2152 2531 2153 2532
rect 2147 2530 2153 2531
rect 2162 2531 2163 2532
rect 2167 2531 2168 2535
rect 2162 2530 2168 2531
rect 2182 2535 2188 2536
rect 2182 2531 2183 2535
rect 2187 2531 2188 2535
rect 2182 2530 2188 2531
rect 2190 2535 2196 2536
rect 2190 2531 2191 2535
rect 2195 2534 2196 2535
rect 2203 2535 2209 2536
rect 2203 2534 2204 2535
rect 2195 2532 2204 2534
rect 2195 2531 2196 2532
rect 2190 2530 2196 2531
rect 2203 2531 2204 2532
rect 2208 2531 2209 2535
rect 2502 2532 2503 2536
rect 2507 2532 2508 2536
rect 2502 2531 2508 2532
rect 2203 2530 2209 2531
rect 203 2523 209 2524
rect 203 2519 204 2523
rect 208 2522 209 2523
rect 214 2523 220 2524
rect 214 2522 215 2523
rect 208 2520 215 2522
rect 208 2519 209 2520
rect 203 2518 209 2519
rect 214 2519 215 2520
rect 219 2519 220 2523
rect 214 2518 220 2519
rect 246 2523 252 2524
rect 246 2519 247 2523
rect 251 2522 252 2523
rect 259 2523 265 2524
rect 259 2522 260 2523
rect 251 2520 260 2522
rect 251 2519 252 2520
rect 246 2518 252 2519
rect 259 2519 260 2520
rect 264 2519 265 2523
rect 259 2518 265 2519
rect 302 2523 308 2524
rect 302 2519 303 2523
rect 307 2522 308 2523
rect 323 2523 329 2524
rect 323 2522 324 2523
rect 307 2520 324 2522
rect 307 2519 308 2520
rect 302 2518 308 2519
rect 323 2519 324 2520
rect 328 2519 329 2523
rect 323 2518 329 2519
rect 366 2523 372 2524
rect 366 2519 367 2523
rect 371 2522 372 2523
rect 395 2523 401 2524
rect 395 2522 396 2523
rect 371 2520 396 2522
rect 371 2519 372 2520
rect 366 2518 372 2519
rect 395 2519 396 2520
rect 400 2519 401 2523
rect 395 2518 401 2519
rect 438 2523 444 2524
rect 438 2519 439 2523
rect 443 2522 444 2523
rect 467 2523 473 2524
rect 467 2522 468 2523
rect 443 2520 468 2522
rect 443 2519 444 2520
rect 438 2518 444 2519
rect 467 2519 468 2520
rect 472 2519 473 2523
rect 467 2518 473 2519
rect 531 2523 537 2524
rect 531 2519 532 2523
rect 536 2522 537 2523
rect 566 2523 572 2524
rect 566 2522 567 2523
rect 536 2520 567 2522
rect 536 2519 537 2520
rect 531 2518 537 2519
rect 566 2519 567 2520
rect 571 2519 572 2523
rect 566 2518 572 2519
rect 574 2523 580 2524
rect 574 2519 575 2523
rect 579 2522 580 2523
rect 595 2523 601 2524
rect 595 2522 596 2523
rect 579 2520 596 2522
rect 579 2519 580 2520
rect 574 2518 580 2519
rect 595 2519 596 2520
rect 600 2519 601 2523
rect 595 2518 601 2519
rect 638 2523 644 2524
rect 638 2519 639 2523
rect 643 2522 644 2523
rect 659 2523 665 2524
rect 659 2522 660 2523
rect 643 2520 660 2522
rect 643 2519 644 2520
rect 638 2518 644 2519
rect 659 2519 660 2520
rect 664 2519 665 2523
rect 659 2518 665 2519
rect 702 2523 708 2524
rect 702 2519 703 2523
rect 707 2522 708 2523
rect 723 2523 729 2524
rect 723 2522 724 2523
rect 707 2520 724 2522
rect 707 2519 708 2520
rect 702 2518 708 2519
rect 723 2519 724 2520
rect 728 2519 729 2523
rect 723 2518 729 2519
rect 762 2523 768 2524
rect 762 2519 763 2523
rect 767 2522 768 2523
rect 787 2523 793 2524
rect 787 2522 788 2523
rect 767 2520 788 2522
rect 767 2519 768 2520
rect 762 2518 768 2519
rect 787 2519 788 2520
rect 792 2519 793 2523
rect 787 2518 793 2519
rect 826 2523 832 2524
rect 826 2519 827 2523
rect 831 2522 832 2523
rect 851 2523 857 2524
rect 851 2522 852 2523
rect 831 2520 852 2522
rect 831 2519 832 2520
rect 826 2518 832 2519
rect 851 2519 852 2520
rect 856 2519 857 2523
rect 851 2518 857 2519
rect 890 2523 896 2524
rect 890 2519 891 2523
rect 895 2522 896 2523
rect 915 2523 921 2524
rect 915 2522 916 2523
rect 895 2520 916 2522
rect 895 2519 896 2520
rect 890 2518 896 2519
rect 915 2519 916 2520
rect 920 2519 921 2523
rect 915 2518 921 2519
rect 958 2523 964 2524
rect 958 2519 959 2523
rect 963 2522 964 2523
rect 979 2523 985 2524
rect 979 2522 980 2523
rect 963 2520 980 2522
rect 963 2519 964 2520
rect 958 2518 964 2519
rect 979 2519 980 2520
rect 984 2519 985 2523
rect 979 2518 985 2519
rect 1018 2523 1024 2524
rect 1018 2519 1019 2523
rect 1023 2522 1024 2523
rect 1043 2523 1049 2524
rect 1043 2522 1044 2523
rect 1023 2520 1044 2522
rect 1023 2519 1024 2520
rect 1018 2518 1024 2519
rect 1043 2519 1044 2520
rect 1048 2519 1049 2523
rect 1043 2518 1049 2519
rect 1491 2515 1497 2516
rect 1491 2511 1492 2515
rect 1496 2514 1497 2515
rect 1526 2515 1532 2516
rect 1526 2514 1527 2515
rect 1496 2512 1527 2514
rect 1496 2511 1497 2512
rect 1491 2510 1497 2511
rect 1526 2511 1527 2512
rect 1531 2511 1532 2515
rect 1526 2510 1532 2511
rect 1534 2515 1540 2516
rect 1534 2511 1535 2515
rect 1539 2514 1540 2515
rect 1547 2515 1553 2516
rect 1547 2514 1548 2515
rect 1539 2512 1548 2514
rect 1539 2511 1540 2512
rect 1534 2510 1540 2511
rect 1547 2511 1548 2512
rect 1552 2511 1553 2515
rect 1547 2510 1553 2511
rect 1598 2515 1609 2516
rect 1598 2511 1599 2515
rect 1603 2511 1604 2515
rect 1608 2511 1609 2515
rect 1598 2510 1609 2511
rect 1658 2515 1665 2516
rect 1658 2511 1659 2515
rect 1664 2511 1665 2515
rect 1658 2510 1665 2511
rect 1714 2515 1721 2516
rect 1714 2511 1715 2515
rect 1720 2511 1721 2515
rect 1714 2510 1721 2511
rect 1770 2515 1777 2516
rect 1770 2511 1771 2515
rect 1776 2511 1777 2515
rect 1770 2510 1777 2511
rect 1814 2515 1820 2516
rect 1814 2511 1815 2515
rect 1819 2514 1820 2515
rect 1827 2515 1833 2516
rect 1827 2514 1828 2515
rect 1819 2512 1828 2514
rect 1819 2511 1820 2512
rect 1814 2510 1820 2511
rect 1827 2511 1828 2512
rect 1832 2511 1833 2515
rect 1827 2510 1833 2511
rect 1882 2515 1889 2516
rect 1882 2511 1883 2515
rect 1888 2511 1889 2515
rect 1882 2510 1889 2511
rect 1938 2515 1945 2516
rect 1938 2511 1939 2515
rect 1944 2511 1945 2515
rect 1938 2510 1945 2511
rect 1994 2515 2001 2516
rect 1994 2511 1995 2515
rect 2000 2511 2001 2515
rect 1994 2510 2001 2511
rect 2050 2515 2057 2516
rect 2050 2511 2051 2515
rect 2056 2511 2057 2515
rect 2050 2510 2057 2511
rect 2102 2515 2113 2516
rect 2102 2511 2103 2515
rect 2107 2511 2108 2515
rect 2112 2511 2113 2515
rect 2102 2510 2113 2511
rect 2162 2515 2169 2516
rect 2162 2511 2163 2515
rect 2168 2511 2169 2515
rect 2162 2510 2169 2511
rect 222 2505 228 2506
rect 110 2504 116 2505
rect 110 2500 111 2504
rect 115 2500 116 2504
rect 222 2501 223 2505
rect 227 2501 228 2505
rect 278 2505 284 2506
rect 222 2500 228 2501
rect 243 2503 252 2504
rect 110 2499 116 2500
rect 243 2499 244 2503
rect 251 2499 252 2503
rect 278 2501 279 2505
rect 283 2501 284 2505
rect 342 2505 348 2506
rect 278 2500 284 2501
rect 299 2503 308 2504
rect 243 2498 252 2499
rect 299 2499 300 2503
rect 307 2499 308 2503
rect 342 2501 343 2505
rect 347 2501 348 2505
rect 414 2505 420 2506
rect 342 2500 348 2501
rect 363 2503 372 2504
rect 299 2498 308 2499
rect 363 2499 364 2503
rect 371 2499 372 2503
rect 414 2501 415 2505
rect 419 2501 420 2505
rect 486 2505 492 2506
rect 414 2500 420 2501
rect 435 2503 444 2504
rect 363 2498 372 2499
rect 435 2499 436 2503
rect 443 2499 444 2503
rect 486 2501 487 2505
rect 491 2501 492 2505
rect 550 2505 556 2506
rect 486 2500 492 2501
rect 494 2503 500 2504
rect 435 2498 444 2499
rect 494 2499 495 2503
rect 499 2502 500 2503
rect 507 2503 513 2504
rect 507 2502 508 2503
rect 499 2500 508 2502
rect 499 2499 500 2500
rect 494 2498 500 2499
rect 507 2499 508 2500
rect 512 2499 513 2503
rect 550 2501 551 2505
rect 555 2501 556 2505
rect 614 2505 620 2506
rect 550 2500 556 2501
rect 571 2503 580 2504
rect 507 2498 513 2499
rect 571 2499 572 2503
rect 579 2499 580 2503
rect 614 2501 615 2505
rect 619 2501 620 2505
rect 678 2505 684 2506
rect 614 2500 620 2501
rect 635 2503 644 2504
rect 571 2498 580 2499
rect 635 2499 636 2503
rect 643 2499 644 2503
rect 678 2501 679 2505
rect 683 2501 684 2505
rect 742 2505 748 2506
rect 678 2500 684 2501
rect 699 2503 708 2504
rect 635 2498 644 2499
rect 699 2499 700 2503
rect 707 2499 708 2503
rect 742 2501 743 2505
rect 747 2501 748 2505
rect 806 2505 812 2506
rect 742 2500 748 2501
rect 762 2503 769 2504
rect 699 2498 708 2499
rect 762 2499 763 2503
rect 768 2499 769 2503
rect 806 2501 807 2505
rect 811 2501 812 2505
rect 870 2505 876 2506
rect 806 2500 812 2501
rect 826 2503 833 2504
rect 762 2498 769 2499
rect 826 2499 827 2503
rect 832 2499 833 2503
rect 870 2501 871 2505
rect 875 2501 876 2505
rect 934 2505 940 2506
rect 870 2500 876 2501
rect 890 2503 897 2504
rect 826 2498 833 2499
rect 890 2499 891 2503
rect 896 2499 897 2503
rect 934 2501 935 2505
rect 939 2501 940 2505
rect 998 2505 1004 2506
rect 934 2500 940 2501
rect 955 2503 964 2504
rect 890 2498 897 2499
rect 955 2499 956 2503
rect 963 2499 964 2503
rect 998 2501 999 2505
rect 1003 2501 1004 2505
rect 1062 2505 1068 2506
rect 998 2500 1004 2501
rect 1018 2503 1025 2504
rect 955 2498 964 2499
rect 1018 2499 1019 2503
rect 1024 2499 1025 2503
rect 1062 2501 1063 2505
rect 1067 2501 1068 2505
rect 1286 2504 1292 2505
rect 1062 2500 1068 2501
rect 1070 2503 1076 2504
rect 1018 2498 1025 2499
rect 1070 2499 1071 2503
rect 1075 2502 1076 2503
rect 1083 2503 1089 2504
rect 1083 2502 1084 2503
rect 1075 2500 1084 2502
rect 1075 2499 1076 2500
rect 1070 2498 1076 2499
rect 1083 2499 1084 2500
rect 1088 2499 1089 2503
rect 1286 2500 1287 2504
rect 1291 2500 1292 2504
rect 1286 2499 1292 2500
rect 1523 2503 1529 2504
rect 1523 2499 1524 2503
rect 1528 2502 1529 2503
rect 1574 2503 1580 2504
rect 1528 2500 1570 2502
rect 1528 2499 1529 2500
rect 1083 2498 1089 2499
rect 1523 2498 1529 2499
rect 1566 2499 1572 2500
rect 1566 2495 1567 2499
rect 1571 2495 1572 2499
rect 1574 2499 1575 2503
rect 1579 2502 1580 2503
rect 1587 2503 1593 2504
rect 1587 2502 1588 2503
rect 1579 2500 1588 2502
rect 1579 2499 1580 2500
rect 1574 2498 1580 2499
rect 1587 2499 1588 2500
rect 1592 2499 1593 2503
rect 1587 2498 1593 2499
rect 1630 2503 1636 2504
rect 1630 2499 1631 2503
rect 1635 2502 1636 2503
rect 1659 2503 1665 2504
rect 1659 2502 1660 2503
rect 1635 2500 1660 2502
rect 1635 2499 1636 2500
rect 1630 2498 1636 2499
rect 1659 2499 1660 2500
rect 1664 2499 1665 2503
rect 1659 2498 1665 2499
rect 1702 2503 1708 2504
rect 1702 2499 1703 2503
rect 1707 2502 1708 2503
rect 1731 2503 1737 2504
rect 1731 2502 1732 2503
rect 1707 2500 1732 2502
rect 1707 2499 1708 2500
rect 1702 2498 1708 2499
rect 1731 2499 1732 2500
rect 1736 2499 1737 2503
rect 1731 2498 1737 2499
rect 1774 2503 1780 2504
rect 1774 2499 1775 2503
rect 1779 2502 1780 2503
rect 1803 2503 1809 2504
rect 1803 2502 1804 2503
rect 1779 2500 1804 2502
rect 1779 2499 1780 2500
rect 1774 2498 1780 2499
rect 1803 2499 1804 2500
rect 1808 2499 1809 2503
rect 1803 2498 1809 2499
rect 1875 2503 1881 2504
rect 1875 2499 1876 2503
rect 1880 2502 1881 2503
rect 1910 2503 1916 2504
rect 1910 2502 1911 2503
rect 1880 2500 1911 2502
rect 1880 2499 1881 2500
rect 1875 2498 1881 2499
rect 1910 2499 1911 2500
rect 1915 2499 1916 2503
rect 1910 2498 1916 2499
rect 1918 2503 1924 2504
rect 1918 2499 1919 2503
rect 1923 2502 1924 2503
rect 1947 2503 1953 2504
rect 1947 2502 1948 2503
rect 1923 2500 1948 2502
rect 1923 2499 1924 2500
rect 1918 2498 1924 2499
rect 1947 2499 1948 2500
rect 1952 2499 1953 2503
rect 1947 2498 1953 2499
rect 1990 2503 1996 2504
rect 1990 2499 1991 2503
rect 1995 2502 1996 2503
rect 2019 2503 2025 2504
rect 2019 2502 2020 2503
rect 1995 2500 2020 2502
rect 1995 2499 1996 2500
rect 1990 2498 1996 2499
rect 2019 2499 2020 2500
rect 2024 2499 2025 2503
rect 2019 2498 2025 2499
rect 2062 2503 2068 2504
rect 2062 2499 2063 2503
rect 2067 2502 2068 2503
rect 2091 2503 2097 2504
rect 2091 2502 2092 2503
rect 2067 2500 2092 2502
rect 2067 2499 2068 2500
rect 2062 2498 2068 2499
rect 2091 2499 2092 2500
rect 2096 2499 2097 2503
rect 2091 2498 2097 2499
rect 2134 2503 2140 2504
rect 2134 2499 2135 2503
rect 2139 2502 2140 2503
rect 2163 2503 2169 2504
rect 2163 2502 2164 2503
rect 2139 2500 2164 2502
rect 2139 2499 2140 2500
rect 2134 2498 2140 2499
rect 2163 2499 2164 2500
rect 2168 2499 2169 2503
rect 2163 2498 2169 2499
rect 1566 2494 1572 2495
rect 110 2487 116 2488
rect 110 2483 111 2487
rect 115 2483 116 2487
rect 1286 2487 1292 2488
rect 110 2482 116 2483
rect 206 2484 212 2485
rect 206 2480 207 2484
rect 211 2480 212 2484
rect 206 2479 212 2480
rect 262 2484 268 2485
rect 262 2480 263 2484
rect 267 2480 268 2484
rect 262 2479 268 2480
rect 326 2484 332 2485
rect 326 2480 327 2484
rect 331 2480 332 2484
rect 326 2479 332 2480
rect 398 2484 404 2485
rect 398 2480 399 2484
rect 403 2480 404 2484
rect 398 2479 404 2480
rect 470 2484 476 2485
rect 470 2480 471 2484
rect 475 2480 476 2484
rect 470 2479 476 2480
rect 534 2484 540 2485
rect 534 2480 535 2484
rect 539 2480 540 2484
rect 534 2479 540 2480
rect 598 2484 604 2485
rect 598 2480 599 2484
rect 603 2480 604 2484
rect 598 2479 604 2480
rect 662 2484 668 2485
rect 662 2480 663 2484
rect 667 2480 668 2484
rect 662 2479 668 2480
rect 726 2484 732 2485
rect 726 2480 727 2484
rect 731 2480 732 2484
rect 726 2479 732 2480
rect 790 2484 796 2485
rect 790 2480 791 2484
rect 795 2480 796 2484
rect 790 2479 796 2480
rect 854 2484 860 2485
rect 854 2480 855 2484
rect 859 2480 860 2484
rect 854 2479 860 2480
rect 918 2484 924 2485
rect 918 2480 919 2484
rect 923 2480 924 2484
rect 918 2479 924 2480
rect 982 2484 988 2485
rect 982 2480 983 2484
rect 987 2480 988 2484
rect 982 2479 988 2480
rect 1046 2484 1052 2485
rect 1046 2480 1047 2484
rect 1051 2480 1052 2484
rect 1286 2483 1287 2487
rect 1291 2483 1292 2487
rect 1542 2485 1548 2486
rect 1286 2482 1292 2483
rect 1326 2484 1332 2485
rect 1046 2479 1052 2480
rect 1326 2480 1327 2484
rect 1331 2480 1332 2484
rect 1542 2481 1543 2485
rect 1547 2481 1548 2485
rect 1606 2485 1612 2486
rect 1542 2480 1548 2481
rect 1563 2483 1569 2484
rect 1326 2479 1332 2480
rect 1563 2479 1564 2483
rect 1568 2482 1569 2483
rect 1574 2483 1580 2484
rect 1574 2482 1575 2483
rect 1568 2480 1575 2482
rect 1568 2479 1569 2480
rect 1563 2478 1569 2479
rect 1574 2479 1575 2480
rect 1579 2479 1580 2483
rect 1606 2481 1607 2485
rect 1611 2481 1612 2485
rect 1678 2485 1684 2486
rect 1606 2480 1612 2481
rect 1627 2483 1636 2484
rect 1574 2478 1580 2479
rect 1627 2479 1628 2483
rect 1635 2479 1636 2483
rect 1678 2481 1679 2485
rect 1683 2481 1684 2485
rect 1750 2485 1756 2486
rect 1678 2480 1684 2481
rect 1699 2483 1708 2484
rect 1627 2478 1636 2479
rect 1699 2479 1700 2483
rect 1707 2479 1708 2483
rect 1750 2481 1751 2485
rect 1755 2481 1756 2485
rect 1822 2485 1828 2486
rect 1750 2480 1756 2481
rect 1771 2483 1780 2484
rect 1699 2478 1708 2479
rect 1771 2479 1772 2483
rect 1779 2479 1780 2483
rect 1822 2481 1823 2485
rect 1827 2481 1828 2485
rect 1894 2485 1900 2486
rect 1822 2480 1828 2481
rect 1842 2483 1849 2484
rect 1771 2478 1780 2479
rect 1842 2479 1843 2483
rect 1848 2479 1849 2483
rect 1894 2481 1895 2485
rect 1899 2481 1900 2485
rect 1966 2485 1972 2486
rect 1894 2480 1900 2481
rect 1915 2483 1924 2484
rect 1842 2478 1849 2479
rect 1915 2479 1916 2483
rect 1923 2479 1924 2483
rect 1966 2481 1967 2485
rect 1971 2481 1972 2485
rect 2038 2485 2044 2486
rect 1966 2480 1972 2481
rect 1987 2483 1996 2484
rect 1915 2478 1924 2479
rect 1987 2479 1988 2483
rect 1995 2479 1996 2483
rect 2038 2481 2039 2485
rect 2043 2481 2044 2485
rect 2110 2485 2116 2486
rect 2038 2480 2044 2481
rect 2059 2483 2068 2484
rect 1987 2478 1996 2479
rect 2059 2479 2060 2483
rect 2067 2479 2068 2483
rect 2110 2481 2111 2485
rect 2115 2481 2116 2485
rect 2182 2485 2188 2486
rect 2110 2480 2116 2481
rect 2131 2483 2140 2484
rect 2059 2478 2068 2479
rect 2131 2479 2132 2483
rect 2139 2479 2140 2483
rect 2182 2481 2183 2485
rect 2187 2481 2188 2485
rect 2502 2484 2508 2485
rect 2182 2480 2188 2481
rect 2190 2483 2196 2484
rect 2131 2478 2140 2479
rect 2190 2479 2191 2483
rect 2195 2482 2196 2483
rect 2203 2483 2209 2484
rect 2203 2482 2204 2483
rect 2195 2480 2204 2482
rect 2195 2479 2196 2480
rect 2190 2478 2196 2479
rect 2203 2479 2204 2480
rect 2208 2479 2209 2483
rect 2502 2480 2503 2484
rect 2507 2480 2508 2484
rect 2502 2479 2508 2480
rect 2203 2478 2209 2479
rect 1326 2467 1332 2468
rect 166 2464 172 2465
rect 110 2461 116 2462
rect 110 2457 111 2461
rect 115 2457 116 2461
rect 166 2460 167 2464
rect 171 2460 172 2464
rect 166 2459 172 2460
rect 222 2464 228 2465
rect 222 2460 223 2464
rect 227 2460 228 2464
rect 222 2459 228 2460
rect 278 2464 284 2465
rect 278 2460 279 2464
rect 283 2460 284 2464
rect 278 2459 284 2460
rect 334 2464 340 2465
rect 334 2460 335 2464
rect 339 2460 340 2464
rect 334 2459 340 2460
rect 390 2464 396 2465
rect 390 2460 391 2464
rect 395 2460 396 2464
rect 390 2459 396 2460
rect 446 2464 452 2465
rect 446 2460 447 2464
rect 451 2460 452 2464
rect 446 2459 452 2460
rect 502 2464 508 2465
rect 502 2460 503 2464
rect 507 2460 508 2464
rect 502 2459 508 2460
rect 558 2464 564 2465
rect 558 2460 559 2464
rect 563 2460 564 2464
rect 558 2459 564 2460
rect 614 2464 620 2465
rect 614 2460 615 2464
rect 619 2460 620 2464
rect 614 2459 620 2460
rect 670 2464 676 2465
rect 670 2460 671 2464
rect 675 2460 676 2464
rect 670 2459 676 2460
rect 726 2464 732 2465
rect 726 2460 727 2464
rect 731 2460 732 2464
rect 726 2459 732 2460
rect 782 2464 788 2465
rect 782 2460 783 2464
rect 787 2460 788 2464
rect 782 2459 788 2460
rect 838 2464 844 2465
rect 838 2460 839 2464
rect 843 2460 844 2464
rect 838 2459 844 2460
rect 894 2464 900 2465
rect 894 2460 895 2464
rect 899 2460 900 2464
rect 894 2459 900 2460
rect 950 2464 956 2465
rect 950 2460 951 2464
rect 955 2460 956 2464
rect 950 2459 956 2460
rect 1006 2464 1012 2465
rect 1006 2460 1007 2464
rect 1011 2460 1012 2464
rect 1006 2459 1012 2460
rect 1062 2464 1068 2465
rect 1062 2460 1063 2464
rect 1067 2460 1068 2464
rect 1326 2463 1327 2467
rect 1331 2463 1332 2467
rect 2502 2467 2508 2468
rect 1326 2462 1332 2463
rect 1526 2464 1532 2465
rect 1062 2459 1068 2460
rect 1286 2461 1292 2462
rect 110 2456 116 2457
rect 1286 2457 1287 2461
rect 1291 2457 1292 2461
rect 1526 2460 1527 2464
rect 1531 2460 1532 2464
rect 1526 2459 1532 2460
rect 1590 2464 1596 2465
rect 1590 2460 1591 2464
rect 1595 2460 1596 2464
rect 1590 2459 1596 2460
rect 1662 2464 1668 2465
rect 1662 2460 1663 2464
rect 1667 2460 1668 2464
rect 1662 2459 1668 2460
rect 1734 2464 1740 2465
rect 1734 2460 1735 2464
rect 1739 2460 1740 2464
rect 1734 2459 1740 2460
rect 1806 2464 1812 2465
rect 1806 2460 1807 2464
rect 1811 2460 1812 2464
rect 1806 2459 1812 2460
rect 1878 2464 1884 2465
rect 1878 2460 1879 2464
rect 1883 2460 1884 2464
rect 1878 2459 1884 2460
rect 1950 2464 1956 2465
rect 1950 2460 1951 2464
rect 1955 2460 1956 2464
rect 1950 2459 1956 2460
rect 2022 2464 2028 2465
rect 2022 2460 2023 2464
rect 2027 2460 2028 2464
rect 2022 2459 2028 2460
rect 2094 2464 2100 2465
rect 2094 2460 2095 2464
rect 2099 2460 2100 2464
rect 2094 2459 2100 2460
rect 2166 2464 2172 2465
rect 2166 2460 2167 2464
rect 2171 2460 2172 2464
rect 2502 2463 2503 2467
rect 2507 2463 2508 2467
rect 2502 2462 2508 2463
rect 2166 2459 2172 2460
rect 1286 2456 1292 2457
rect 1542 2448 1548 2449
rect 1326 2445 1332 2446
rect 110 2444 116 2445
rect 1286 2444 1292 2445
rect 110 2440 111 2444
rect 115 2440 116 2444
rect 110 2439 116 2440
rect 182 2443 188 2444
rect 182 2439 183 2443
rect 187 2439 188 2443
rect 182 2438 188 2439
rect 203 2443 209 2444
rect 203 2439 204 2443
rect 208 2442 209 2443
rect 218 2443 224 2444
rect 218 2442 219 2443
rect 208 2440 219 2442
rect 208 2439 209 2440
rect 203 2438 209 2439
rect 218 2439 219 2440
rect 223 2439 224 2443
rect 218 2438 224 2439
rect 238 2443 244 2444
rect 238 2439 239 2443
rect 243 2439 244 2443
rect 238 2438 244 2439
rect 259 2443 265 2444
rect 259 2439 260 2443
rect 264 2442 265 2443
rect 274 2443 280 2444
rect 274 2442 275 2443
rect 264 2440 275 2442
rect 264 2439 265 2440
rect 259 2438 265 2439
rect 274 2439 275 2440
rect 279 2439 280 2443
rect 274 2438 280 2439
rect 294 2443 300 2444
rect 294 2439 295 2443
rect 299 2439 300 2443
rect 294 2438 300 2439
rect 315 2443 321 2444
rect 315 2439 316 2443
rect 320 2442 321 2443
rect 330 2443 336 2444
rect 330 2442 331 2443
rect 320 2440 331 2442
rect 320 2439 321 2440
rect 315 2438 321 2439
rect 330 2439 331 2440
rect 335 2439 336 2443
rect 330 2438 336 2439
rect 350 2443 356 2444
rect 350 2439 351 2443
rect 355 2439 356 2443
rect 350 2438 356 2439
rect 371 2443 377 2444
rect 371 2439 372 2443
rect 376 2442 377 2443
rect 386 2443 392 2444
rect 386 2442 387 2443
rect 376 2440 387 2442
rect 376 2439 377 2440
rect 371 2438 377 2439
rect 386 2439 387 2440
rect 391 2439 392 2443
rect 386 2438 392 2439
rect 406 2443 412 2444
rect 406 2439 407 2443
rect 411 2439 412 2443
rect 406 2438 412 2439
rect 427 2443 433 2444
rect 427 2439 428 2443
rect 432 2442 433 2443
rect 442 2443 448 2444
rect 442 2442 443 2443
rect 432 2440 443 2442
rect 432 2439 433 2440
rect 427 2438 433 2439
rect 442 2439 443 2440
rect 447 2439 448 2443
rect 442 2438 448 2439
rect 462 2443 468 2444
rect 462 2439 463 2443
rect 467 2439 468 2443
rect 462 2438 468 2439
rect 483 2443 489 2444
rect 483 2439 484 2443
rect 488 2442 489 2443
rect 498 2443 504 2444
rect 498 2442 499 2443
rect 488 2440 499 2442
rect 488 2439 489 2440
rect 483 2438 489 2439
rect 498 2439 499 2440
rect 503 2439 504 2443
rect 498 2438 504 2439
rect 518 2443 524 2444
rect 518 2439 519 2443
rect 523 2439 524 2443
rect 518 2438 524 2439
rect 539 2443 545 2444
rect 539 2439 540 2443
rect 544 2442 545 2443
rect 554 2443 560 2444
rect 554 2442 555 2443
rect 544 2440 555 2442
rect 544 2439 545 2440
rect 539 2438 545 2439
rect 554 2439 555 2440
rect 559 2439 560 2443
rect 554 2438 560 2439
rect 574 2443 580 2444
rect 574 2439 575 2443
rect 579 2439 580 2443
rect 574 2438 580 2439
rect 595 2443 601 2444
rect 595 2439 596 2443
rect 600 2442 601 2443
rect 610 2443 616 2444
rect 610 2442 611 2443
rect 600 2440 611 2442
rect 600 2439 601 2440
rect 595 2438 601 2439
rect 610 2439 611 2440
rect 615 2439 616 2443
rect 610 2438 616 2439
rect 630 2443 636 2444
rect 630 2439 631 2443
rect 635 2439 636 2443
rect 630 2438 636 2439
rect 651 2443 657 2444
rect 651 2439 652 2443
rect 656 2442 657 2443
rect 666 2443 672 2444
rect 666 2442 667 2443
rect 656 2440 667 2442
rect 656 2439 657 2440
rect 651 2438 657 2439
rect 666 2439 667 2440
rect 671 2439 672 2443
rect 666 2438 672 2439
rect 686 2443 692 2444
rect 686 2439 687 2443
rect 691 2439 692 2443
rect 686 2438 692 2439
rect 707 2443 713 2444
rect 707 2439 708 2443
rect 712 2442 713 2443
rect 722 2443 728 2444
rect 722 2442 723 2443
rect 712 2440 723 2442
rect 712 2439 713 2440
rect 707 2438 713 2439
rect 722 2439 723 2440
rect 727 2439 728 2443
rect 722 2438 728 2439
rect 742 2443 748 2444
rect 742 2439 743 2443
rect 747 2439 748 2443
rect 742 2438 748 2439
rect 763 2443 769 2444
rect 763 2439 764 2443
rect 768 2442 769 2443
rect 778 2443 784 2444
rect 778 2442 779 2443
rect 768 2440 779 2442
rect 768 2439 769 2440
rect 763 2438 769 2439
rect 778 2439 779 2440
rect 783 2439 784 2443
rect 778 2438 784 2439
rect 798 2443 804 2444
rect 798 2439 799 2443
rect 803 2439 804 2443
rect 798 2438 804 2439
rect 819 2443 825 2444
rect 819 2439 820 2443
rect 824 2442 825 2443
rect 834 2443 840 2444
rect 834 2442 835 2443
rect 824 2440 835 2442
rect 824 2439 825 2440
rect 819 2438 825 2439
rect 834 2439 835 2440
rect 839 2439 840 2443
rect 834 2438 840 2439
rect 854 2443 860 2444
rect 854 2439 855 2443
rect 859 2439 860 2443
rect 854 2438 860 2439
rect 874 2443 881 2444
rect 874 2439 875 2443
rect 880 2439 881 2443
rect 874 2438 881 2439
rect 910 2443 916 2444
rect 910 2439 911 2443
rect 915 2439 916 2443
rect 910 2438 916 2439
rect 918 2443 924 2444
rect 918 2439 919 2443
rect 923 2442 924 2443
rect 931 2443 937 2444
rect 931 2442 932 2443
rect 923 2440 932 2442
rect 923 2439 924 2440
rect 918 2438 924 2439
rect 931 2439 932 2440
rect 936 2439 937 2443
rect 931 2438 937 2439
rect 966 2443 972 2444
rect 966 2439 967 2443
rect 971 2439 972 2443
rect 966 2438 972 2439
rect 974 2443 980 2444
rect 974 2439 975 2443
rect 979 2442 980 2443
rect 987 2443 993 2444
rect 987 2442 988 2443
rect 979 2440 988 2442
rect 979 2439 980 2440
rect 974 2438 980 2439
rect 987 2439 988 2440
rect 992 2439 993 2443
rect 987 2438 993 2439
rect 1022 2443 1028 2444
rect 1022 2439 1023 2443
rect 1027 2439 1028 2443
rect 1043 2443 1049 2444
rect 1043 2442 1044 2443
rect 1022 2438 1028 2439
rect 1032 2440 1044 2442
rect 1032 2434 1034 2440
rect 1043 2439 1044 2440
rect 1048 2439 1049 2443
rect 1043 2438 1049 2439
rect 1078 2443 1084 2444
rect 1078 2439 1079 2443
rect 1083 2439 1084 2443
rect 1099 2443 1105 2444
rect 1099 2442 1100 2443
rect 1078 2438 1084 2439
rect 1088 2440 1100 2442
rect 948 2432 1034 2434
rect 948 2426 950 2432
rect 1088 2430 1090 2440
rect 1099 2439 1100 2440
rect 1104 2439 1105 2443
rect 1286 2440 1287 2444
rect 1291 2440 1292 2444
rect 1326 2441 1327 2445
rect 1331 2441 1332 2445
rect 1542 2444 1543 2448
rect 1547 2444 1548 2448
rect 1542 2443 1548 2444
rect 1606 2448 1612 2449
rect 1606 2444 1607 2448
rect 1611 2444 1612 2448
rect 1606 2443 1612 2444
rect 1670 2448 1676 2449
rect 1670 2444 1671 2448
rect 1675 2444 1676 2448
rect 1670 2443 1676 2444
rect 1742 2448 1748 2449
rect 1742 2444 1743 2448
rect 1747 2444 1748 2448
rect 1742 2443 1748 2444
rect 1814 2448 1820 2449
rect 1814 2444 1815 2448
rect 1819 2444 1820 2448
rect 1814 2443 1820 2444
rect 1878 2448 1884 2449
rect 1878 2444 1879 2448
rect 1883 2444 1884 2448
rect 1878 2443 1884 2444
rect 1950 2448 1956 2449
rect 1950 2444 1951 2448
rect 1955 2444 1956 2448
rect 1950 2443 1956 2444
rect 2022 2448 2028 2449
rect 2022 2444 2023 2448
rect 2027 2444 2028 2448
rect 2022 2443 2028 2444
rect 2094 2448 2100 2449
rect 2094 2444 2095 2448
rect 2099 2444 2100 2448
rect 2094 2443 2100 2444
rect 2166 2448 2172 2449
rect 2166 2444 2167 2448
rect 2171 2444 2172 2448
rect 2166 2443 2172 2444
rect 2502 2445 2508 2446
rect 1326 2440 1332 2441
rect 2502 2441 2503 2445
rect 2507 2441 2508 2445
rect 2502 2440 2508 2441
rect 1286 2439 1292 2440
rect 1099 2438 1105 2439
rect 1004 2428 1090 2430
rect 1326 2428 1332 2429
rect 2502 2428 2508 2429
rect 1004 2426 1006 2428
rect 947 2425 953 2426
rect 163 2423 172 2424
rect 163 2419 164 2423
rect 171 2419 172 2423
rect 163 2418 172 2419
rect 218 2423 225 2424
rect 218 2419 219 2423
rect 224 2419 225 2423
rect 218 2418 225 2419
rect 274 2423 281 2424
rect 274 2419 275 2423
rect 280 2419 281 2423
rect 274 2418 281 2419
rect 330 2423 337 2424
rect 330 2419 331 2423
rect 336 2419 337 2423
rect 330 2418 337 2419
rect 386 2423 393 2424
rect 386 2419 387 2423
rect 392 2419 393 2423
rect 386 2418 393 2419
rect 442 2423 449 2424
rect 442 2419 443 2423
rect 448 2419 449 2423
rect 442 2418 449 2419
rect 498 2423 505 2424
rect 498 2419 499 2423
rect 504 2419 505 2423
rect 498 2418 505 2419
rect 554 2423 561 2424
rect 554 2419 555 2423
rect 560 2419 561 2423
rect 554 2418 561 2419
rect 610 2423 617 2424
rect 610 2419 611 2423
rect 616 2419 617 2423
rect 610 2418 617 2419
rect 666 2423 673 2424
rect 666 2419 667 2423
rect 672 2419 673 2423
rect 666 2418 673 2419
rect 722 2423 729 2424
rect 722 2419 723 2423
rect 728 2419 729 2423
rect 722 2418 729 2419
rect 778 2423 785 2424
rect 778 2419 779 2423
rect 784 2419 785 2423
rect 778 2418 785 2419
rect 834 2423 841 2424
rect 834 2419 835 2423
rect 840 2419 841 2423
rect 834 2418 841 2419
rect 891 2423 897 2424
rect 891 2419 892 2423
rect 896 2422 897 2423
rect 896 2420 942 2422
rect 947 2421 948 2425
rect 952 2421 953 2425
rect 947 2420 953 2421
rect 1003 2425 1009 2426
rect 1003 2421 1004 2425
rect 1008 2421 1009 2425
rect 1326 2424 1327 2428
rect 1331 2424 1332 2428
rect 1003 2420 1009 2421
rect 1059 2423 1065 2424
rect 896 2419 897 2420
rect 891 2418 897 2419
rect 940 2418 942 2420
rect 974 2419 980 2420
rect 974 2418 975 2419
rect 940 2416 975 2418
rect 974 2415 975 2416
rect 979 2415 980 2419
rect 1059 2419 1060 2423
rect 1064 2422 1065 2423
rect 1070 2423 1076 2424
rect 1326 2423 1332 2424
rect 1558 2427 1564 2428
rect 1558 2423 1559 2427
rect 1563 2423 1564 2427
rect 1070 2422 1071 2423
rect 1064 2420 1071 2422
rect 1064 2419 1065 2420
rect 1059 2418 1065 2419
rect 1070 2419 1071 2420
rect 1075 2419 1076 2423
rect 1558 2422 1564 2423
rect 1566 2427 1572 2428
rect 1566 2423 1567 2427
rect 1571 2426 1572 2427
rect 1579 2427 1585 2428
rect 1579 2426 1580 2427
rect 1571 2424 1580 2426
rect 1571 2423 1572 2424
rect 1566 2422 1572 2423
rect 1579 2423 1580 2424
rect 1584 2423 1585 2427
rect 1579 2422 1585 2423
rect 1622 2427 1628 2428
rect 1622 2423 1623 2427
rect 1627 2423 1628 2427
rect 1643 2427 1649 2428
rect 1643 2426 1644 2427
rect 1622 2422 1628 2423
rect 1632 2424 1644 2426
rect 1070 2418 1076 2419
rect 1632 2418 1634 2424
rect 1643 2423 1644 2424
rect 1648 2423 1649 2427
rect 1643 2422 1649 2423
rect 1686 2427 1692 2428
rect 1686 2423 1687 2427
rect 1691 2423 1692 2427
rect 1707 2427 1713 2428
rect 1707 2426 1708 2427
rect 1686 2422 1692 2423
rect 1696 2424 1708 2426
rect 974 2414 980 2415
rect 1540 2416 1634 2418
rect 1540 2410 1542 2416
rect 1696 2414 1698 2424
rect 1707 2423 1708 2424
rect 1712 2423 1713 2427
rect 1707 2422 1713 2423
rect 1758 2427 1764 2428
rect 1758 2423 1759 2427
rect 1763 2423 1764 2427
rect 1779 2427 1785 2428
rect 1779 2426 1780 2427
rect 1758 2422 1764 2423
rect 1768 2424 1780 2426
rect 1768 2418 1770 2424
rect 1779 2423 1780 2424
rect 1784 2423 1785 2427
rect 1779 2422 1785 2423
rect 1830 2427 1836 2428
rect 1830 2423 1831 2427
rect 1835 2423 1836 2427
rect 1851 2427 1857 2428
rect 1851 2426 1852 2427
rect 1830 2422 1836 2423
rect 1840 2424 1852 2426
rect 1604 2412 1698 2414
rect 1700 2416 1770 2418
rect 1604 2410 1606 2412
rect 1700 2410 1702 2416
rect 1840 2414 1842 2424
rect 1851 2423 1852 2424
rect 1856 2423 1857 2427
rect 1851 2422 1857 2423
rect 1894 2427 1900 2428
rect 1894 2423 1895 2427
rect 1899 2423 1900 2427
rect 1894 2422 1900 2423
rect 1915 2427 1921 2428
rect 1915 2423 1916 2427
rect 1920 2426 1921 2427
rect 1946 2427 1952 2428
rect 1946 2426 1947 2427
rect 1920 2424 1947 2426
rect 1920 2423 1921 2424
rect 1915 2422 1921 2423
rect 1946 2423 1947 2424
rect 1951 2423 1952 2427
rect 1946 2422 1952 2423
rect 1966 2427 1972 2428
rect 1966 2423 1967 2427
rect 1971 2423 1972 2427
rect 1966 2422 1972 2423
rect 1974 2427 1980 2428
rect 1974 2423 1975 2427
rect 1979 2426 1980 2427
rect 1987 2427 1993 2428
rect 1987 2426 1988 2427
rect 1979 2424 1988 2426
rect 1979 2423 1980 2424
rect 1974 2422 1980 2423
rect 1987 2423 1988 2424
rect 1992 2423 1993 2427
rect 1987 2422 1993 2423
rect 2038 2427 2044 2428
rect 2038 2423 2039 2427
rect 2043 2423 2044 2427
rect 2038 2422 2044 2423
rect 2054 2427 2065 2428
rect 2054 2423 2055 2427
rect 2059 2423 2060 2427
rect 2064 2423 2065 2427
rect 2054 2422 2065 2423
rect 2110 2427 2116 2428
rect 2110 2423 2111 2427
rect 2115 2423 2116 2427
rect 2131 2427 2137 2428
rect 2131 2426 2132 2427
rect 2110 2422 2116 2423
rect 2120 2424 2132 2426
rect 2120 2418 2122 2424
rect 2131 2423 2132 2424
rect 2136 2423 2137 2427
rect 2131 2422 2137 2423
rect 2182 2427 2188 2428
rect 2182 2423 2183 2427
rect 2187 2423 2188 2427
rect 2203 2427 2209 2428
rect 2203 2426 2204 2427
rect 2182 2422 2188 2423
rect 2192 2424 2204 2426
rect 1741 2412 1842 2414
rect 2020 2416 2122 2418
rect 1741 2410 1743 2412
rect 2020 2410 2022 2416
rect 2192 2414 2194 2424
rect 2203 2423 2204 2424
rect 2208 2423 2209 2427
rect 2502 2424 2503 2428
rect 2507 2424 2508 2428
rect 2502 2423 2508 2424
rect 2203 2422 2209 2423
rect 2092 2412 2194 2414
rect 2092 2410 2094 2412
rect 1539 2409 1545 2410
rect 1539 2405 1540 2409
rect 1544 2405 1545 2409
rect 1539 2404 1545 2405
rect 1603 2409 1609 2410
rect 1603 2405 1604 2409
rect 1608 2405 1609 2409
rect 1603 2404 1609 2405
rect 1667 2409 1702 2410
rect 1667 2405 1668 2409
rect 1672 2408 1702 2409
rect 1739 2409 1745 2410
rect 1672 2405 1673 2408
rect 1667 2404 1673 2405
rect 1739 2405 1740 2409
rect 1744 2405 1745 2409
rect 2019 2409 2025 2410
rect 1739 2404 1745 2405
rect 1810 2407 1817 2408
rect 1810 2403 1811 2407
rect 1816 2403 1817 2407
rect 1810 2402 1817 2403
rect 1875 2407 1881 2408
rect 1875 2403 1876 2407
rect 1880 2406 1881 2407
rect 1946 2407 1953 2408
rect 1880 2404 1938 2406
rect 1880 2403 1881 2404
rect 1875 2402 1881 2403
rect 499 2399 505 2400
rect 499 2395 500 2399
rect 504 2398 505 2399
rect 555 2399 561 2400
rect 504 2396 550 2398
rect 504 2395 505 2396
rect 499 2394 505 2395
rect 548 2386 550 2396
rect 555 2395 556 2399
rect 560 2398 561 2399
rect 611 2399 617 2400
rect 560 2396 606 2398
rect 560 2395 561 2396
rect 555 2394 561 2395
rect 604 2386 606 2396
rect 611 2395 612 2399
rect 616 2398 617 2399
rect 667 2399 673 2400
rect 616 2396 662 2398
rect 616 2395 617 2396
rect 611 2394 617 2395
rect 660 2386 662 2396
rect 667 2395 668 2399
rect 672 2398 673 2399
rect 918 2399 924 2400
rect 918 2398 919 2399
rect 672 2396 919 2398
rect 672 2395 673 2396
rect 667 2394 673 2395
rect 918 2395 919 2396
rect 923 2395 924 2399
rect 1936 2398 1938 2404
rect 1946 2403 1947 2407
rect 1952 2403 1953 2407
rect 2019 2405 2020 2409
rect 2024 2405 2025 2409
rect 2019 2404 2025 2405
rect 2091 2409 2097 2410
rect 2091 2405 2092 2409
rect 2096 2405 2097 2409
rect 2091 2404 2097 2405
rect 2163 2407 2169 2408
rect 1946 2402 1953 2403
rect 2163 2403 2164 2407
rect 2168 2406 2169 2407
rect 2190 2407 2196 2408
rect 2190 2406 2191 2407
rect 2168 2404 2191 2406
rect 2168 2403 2169 2404
rect 2163 2402 2169 2403
rect 2190 2403 2191 2404
rect 2195 2403 2196 2407
rect 2190 2402 2196 2403
rect 2054 2399 2060 2400
rect 2054 2398 2055 2399
rect 1936 2396 2055 2398
rect 918 2394 924 2395
rect 2054 2395 2055 2396
rect 2059 2395 2060 2399
rect 2054 2394 2060 2395
rect 1547 2391 1553 2392
rect 1547 2387 1548 2391
rect 1552 2387 1553 2391
rect 1547 2386 1553 2387
rect 1590 2391 1596 2392
rect 1590 2387 1591 2391
rect 1595 2390 1596 2391
rect 1603 2391 1609 2392
rect 1603 2390 1604 2391
rect 1595 2388 1604 2390
rect 1595 2387 1596 2388
rect 1590 2386 1596 2387
rect 1603 2387 1604 2388
rect 1608 2387 1609 2391
rect 1603 2386 1609 2387
rect 1646 2391 1652 2392
rect 1646 2387 1647 2391
rect 1651 2390 1652 2391
rect 1659 2391 1665 2392
rect 1659 2390 1660 2391
rect 1651 2388 1660 2390
rect 1651 2387 1652 2388
rect 1646 2386 1652 2387
rect 1659 2387 1660 2388
rect 1664 2387 1665 2391
rect 1659 2386 1665 2387
rect 1702 2391 1708 2392
rect 1702 2387 1703 2391
rect 1707 2390 1708 2391
rect 1715 2391 1721 2392
rect 1715 2390 1716 2391
rect 1707 2388 1716 2390
rect 1707 2387 1708 2388
rect 1702 2386 1708 2387
rect 1715 2387 1716 2388
rect 1720 2387 1721 2391
rect 1715 2386 1721 2387
rect 1766 2391 1777 2392
rect 1766 2387 1767 2391
rect 1771 2387 1772 2391
rect 1776 2387 1777 2391
rect 1766 2386 1777 2387
rect 1835 2391 1841 2392
rect 1835 2387 1836 2391
rect 1840 2390 1841 2391
rect 1899 2391 1905 2392
rect 1840 2388 1894 2390
rect 1840 2387 1841 2388
rect 1835 2386 1841 2387
rect 548 2384 598 2386
rect 604 2384 654 2386
rect 660 2384 710 2386
rect 596 2382 598 2384
rect 652 2382 654 2384
rect 708 2382 710 2384
rect 1549 2382 1551 2386
rect 1782 2383 1788 2384
rect 1782 2382 1783 2383
rect 518 2381 524 2382
rect 110 2380 116 2381
rect 110 2376 111 2380
rect 115 2376 116 2380
rect 518 2377 519 2381
rect 523 2377 524 2381
rect 574 2381 580 2382
rect 518 2376 524 2377
rect 539 2379 548 2380
rect 110 2375 116 2376
rect 539 2375 540 2379
rect 547 2375 548 2379
rect 574 2377 575 2381
rect 579 2377 580 2381
rect 574 2376 580 2377
rect 595 2381 601 2382
rect 595 2377 596 2381
rect 600 2377 601 2381
rect 595 2376 601 2377
rect 630 2381 636 2382
rect 630 2377 631 2381
rect 635 2377 636 2381
rect 630 2376 636 2377
rect 651 2381 657 2382
rect 651 2377 652 2381
rect 656 2377 657 2381
rect 651 2376 657 2377
rect 686 2381 692 2382
rect 686 2377 687 2381
rect 691 2377 692 2381
rect 686 2376 692 2377
rect 707 2381 713 2382
rect 707 2377 708 2381
rect 712 2377 713 2381
rect 707 2376 713 2377
rect 1286 2380 1292 2381
rect 1549 2380 1783 2382
rect 1286 2376 1287 2380
rect 1291 2376 1292 2380
rect 1782 2379 1783 2380
rect 1787 2379 1788 2383
rect 1782 2378 1788 2379
rect 1892 2378 1894 2388
rect 1899 2387 1900 2391
rect 1904 2390 1905 2391
rect 1963 2391 1969 2392
rect 1904 2388 1954 2390
rect 1904 2387 1905 2388
rect 1899 2386 1905 2387
rect 1952 2378 1954 2388
rect 1963 2387 1964 2391
rect 1968 2390 1969 2391
rect 1974 2391 1980 2392
rect 1974 2390 1975 2391
rect 1968 2388 1975 2390
rect 1968 2387 1969 2388
rect 1963 2386 1969 2387
rect 1974 2387 1975 2388
rect 1979 2387 1980 2391
rect 1974 2386 1980 2387
rect 2006 2391 2012 2392
rect 2006 2387 2007 2391
rect 2011 2390 2012 2391
rect 2027 2391 2033 2392
rect 2027 2390 2028 2391
rect 2011 2388 2028 2390
rect 2011 2387 2012 2388
rect 2006 2386 2012 2387
rect 2027 2387 2028 2388
rect 2032 2387 2033 2391
rect 2027 2386 2033 2387
rect 2070 2391 2076 2392
rect 2070 2387 2071 2391
rect 2075 2390 2076 2391
rect 2091 2391 2097 2392
rect 2091 2390 2092 2391
rect 2075 2388 2092 2390
rect 2075 2387 2076 2388
rect 2070 2386 2076 2387
rect 2091 2387 2092 2388
rect 2096 2387 2097 2391
rect 2091 2386 2097 2387
rect 1892 2376 1942 2378
rect 1952 2376 2134 2378
rect 1286 2375 1292 2376
rect 539 2374 548 2375
rect 1940 2374 1942 2376
rect 2132 2374 2134 2376
rect 1566 2373 1572 2374
rect 1326 2372 1332 2373
rect 1326 2368 1327 2372
rect 1331 2368 1332 2372
rect 1566 2369 1567 2373
rect 1571 2369 1572 2373
rect 1622 2373 1628 2374
rect 1566 2368 1572 2369
rect 1587 2371 1596 2372
rect 1326 2367 1332 2368
rect 1587 2367 1588 2371
rect 1595 2367 1596 2371
rect 1622 2369 1623 2373
rect 1627 2369 1628 2373
rect 1678 2373 1684 2374
rect 1622 2368 1628 2369
rect 1643 2371 1652 2372
rect 1587 2366 1596 2367
rect 1643 2367 1644 2371
rect 1651 2367 1652 2371
rect 1678 2369 1679 2373
rect 1683 2369 1684 2373
rect 1734 2373 1740 2374
rect 1678 2368 1684 2369
rect 1699 2371 1708 2372
rect 1643 2366 1652 2367
rect 1699 2367 1700 2371
rect 1707 2367 1708 2371
rect 1734 2369 1735 2373
rect 1739 2369 1740 2373
rect 1790 2373 1796 2374
rect 1734 2368 1740 2369
rect 1755 2371 1761 2372
rect 1699 2366 1708 2367
rect 1755 2367 1756 2371
rect 1760 2370 1761 2371
rect 1766 2371 1772 2372
rect 1766 2370 1767 2371
rect 1760 2368 1767 2370
rect 1760 2367 1761 2368
rect 1755 2366 1761 2367
rect 1766 2367 1767 2368
rect 1771 2367 1772 2371
rect 1790 2369 1791 2373
rect 1795 2369 1796 2373
rect 1854 2373 1860 2374
rect 1790 2368 1796 2369
rect 1810 2371 1817 2372
rect 1766 2366 1772 2367
rect 1810 2367 1811 2371
rect 1816 2367 1817 2371
rect 1854 2369 1855 2373
rect 1859 2369 1860 2373
rect 1918 2373 1924 2374
rect 1854 2368 1860 2369
rect 1862 2371 1868 2372
rect 1810 2366 1817 2367
rect 1862 2367 1863 2371
rect 1867 2370 1868 2371
rect 1875 2371 1881 2372
rect 1875 2370 1876 2371
rect 1867 2368 1876 2370
rect 1867 2367 1868 2368
rect 1862 2366 1868 2367
rect 1875 2367 1876 2368
rect 1880 2367 1881 2371
rect 1918 2369 1919 2373
rect 1923 2369 1924 2373
rect 1918 2368 1924 2369
rect 1939 2373 1945 2374
rect 1939 2369 1940 2373
rect 1944 2369 1945 2373
rect 1939 2368 1945 2369
rect 1982 2373 1988 2374
rect 1982 2369 1983 2373
rect 1987 2369 1988 2373
rect 2046 2373 2052 2374
rect 1982 2368 1988 2369
rect 2003 2371 2012 2372
rect 1875 2366 1881 2367
rect 2003 2367 2004 2371
rect 2011 2367 2012 2371
rect 2046 2369 2047 2373
rect 2051 2369 2052 2373
rect 2110 2373 2116 2374
rect 2046 2368 2052 2369
rect 2067 2371 2076 2372
rect 2003 2366 2012 2367
rect 2067 2367 2068 2371
rect 2075 2367 2076 2371
rect 2110 2369 2111 2373
rect 2115 2369 2116 2373
rect 2110 2368 2116 2369
rect 2131 2373 2137 2374
rect 2131 2369 2132 2373
rect 2136 2369 2137 2373
rect 2131 2368 2137 2369
rect 2502 2372 2508 2373
rect 2502 2368 2503 2372
rect 2507 2368 2508 2372
rect 2502 2367 2508 2368
rect 2067 2366 2076 2367
rect 110 2363 116 2364
rect 110 2359 111 2363
rect 115 2359 116 2363
rect 1286 2363 1292 2364
rect 110 2358 116 2359
rect 502 2360 508 2361
rect 502 2356 503 2360
rect 507 2356 508 2360
rect 502 2355 508 2356
rect 558 2360 564 2361
rect 558 2356 559 2360
rect 563 2356 564 2360
rect 558 2355 564 2356
rect 614 2360 620 2361
rect 614 2356 615 2360
rect 619 2356 620 2360
rect 614 2355 620 2356
rect 670 2360 676 2361
rect 670 2356 671 2360
rect 675 2356 676 2360
rect 1286 2359 1287 2363
rect 1291 2359 1292 2363
rect 1286 2358 1292 2359
rect 670 2355 676 2356
rect 1326 2355 1332 2356
rect 1326 2351 1327 2355
rect 1331 2351 1332 2355
rect 2502 2355 2508 2356
rect 1326 2350 1332 2351
rect 1550 2352 1556 2353
rect 1550 2348 1551 2352
rect 1555 2348 1556 2352
rect 1550 2347 1556 2348
rect 1606 2352 1612 2353
rect 1606 2348 1607 2352
rect 1611 2348 1612 2352
rect 1606 2347 1612 2348
rect 1662 2352 1668 2353
rect 1662 2348 1663 2352
rect 1667 2348 1668 2352
rect 1662 2347 1668 2348
rect 1718 2352 1724 2353
rect 1718 2348 1719 2352
rect 1723 2348 1724 2352
rect 1718 2347 1724 2348
rect 1774 2352 1780 2353
rect 1774 2348 1775 2352
rect 1779 2348 1780 2352
rect 1774 2347 1780 2348
rect 1838 2352 1844 2353
rect 1838 2348 1839 2352
rect 1843 2348 1844 2352
rect 1838 2347 1844 2348
rect 1902 2352 1908 2353
rect 1902 2348 1903 2352
rect 1907 2348 1908 2352
rect 1902 2347 1908 2348
rect 1966 2352 1972 2353
rect 1966 2348 1967 2352
rect 1971 2348 1972 2352
rect 1966 2347 1972 2348
rect 2030 2352 2036 2353
rect 2030 2348 2031 2352
rect 2035 2348 2036 2352
rect 2030 2347 2036 2348
rect 2094 2352 2100 2353
rect 2094 2348 2095 2352
rect 2099 2348 2100 2352
rect 2502 2351 2503 2355
rect 2507 2351 2508 2355
rect 2502 2350 2508 2351
rect 2094 2347 2100 2348
rect 318 2340 324 2341
rect 110 2337 116 2338
rect 110 2333 111 2337
rect 115 2333 116 2337
rect 318 2336 319 2340
rect 323 2336 324 2340
rect 318 2335 324 2336
rect 390 2340 396 2341
rect 390 2336 391 2340
rect 395 2336 396 2340
rect 390 2335 396 2336
rect 462 2340 468 2341
rect 462 2336 463 2340
rect 467 2336 468 2340
rect 462 2335 468 2336
rect 534 2340 540 2341
rect 534 2336 535 2340
rect 539 2336 540 2340
rect 534 2335 540 2336
rect 606 2340 612 2341
rect 606 2336 607 2340
rect 611 2336 612 2340
rect 606 2335 612 2336
rect 678 2340 684 2341
rect 678 2336 679 2340
rect 683 2336 684 2340
rect 678 2335 684 2336
rect 742 2340 748 2341
rect 742 2336 743 2340
rect 747 2336 748 2340
rect 742 2335 748 2336
rect 806 2340 812 2341
rect 806 2336 807 2340
rect 811 2336 812 2340
rect 806 2335 812 2336
rect 862 2340 868 2341
rect 862 2336 863 2340
rect 867 2336 868 2340
rect 862 2335 868 2336
rect 926 2340 932 2341
rect 926 2336 927 2340
rect 931 2336 932 2340
rect 926 2335 932 2336
rect 990 2340 996 2341
rect 990 2336 991 2340
rect 995 2336 996 2340
rect 990 2335 996 2336
rect 1054 2340 1060 2341
rect 1054 2336 1055 2340
rect 1059 2336 1060 2340
rect 1054 2335 1060 2336
rect 1110 2340 1116 2341
rect 1110 2336 1111 2340
rect 1115 2336 1116 2340
rect 1110 2335 1116 2336
rect 1166 2340 1172 2341
rect 1166 2336 1167 2340
rect 1171 2336 1172 2340
rect 1166 2335 1172 2336
rect 1222 2340 1228 2341
rect 1222 2336 1223 2340
rect 1227 2336 1228 2340
rect 1222 2335 1228 2336
rect 1286 2337 1292 2338
rect 110 2332 116 2333
rect 1286 2333 1287 2337
rect 1291 2333 1292 2337
rect 1286 2332 1292 2333
rect 1470 2332 1476 2333
rect 1326 2329 1332 2330
rect 1326 2325 1327 2329
rect 1331 2325 1332 2329
rect 1470 2328 1471 2332
rect 1475 2328 1476 2332
rect 1470 2327 1476 2328
rect 1534 2332 1540 2333
rect 1534 2328 1535 2332
rect 1539 2328 1540 2332
rect 1534 2327 1540 2328
rect 1606 2332 1612 2333
rect 1606 2328 1607 2332
rect 1611 2328 1612 2332
rect 1606 2327 1612 2328
rect 1686 2332 1692 2333
rect 1686 2328 1687 2332
rect 1691 2328 1692 2332
rect 1686 2327 1692 2328
rect 1758 2332 1764 2333
rect 1758 2328 1759 2332
rect 1763 2328 1764 2332
rect 1758 2327 1764 2328
rect 1830 2332 1836 2333
rect 1830 2328 1831 2332
rect 1835 2328 1836 2332
rect 1830 2327 1836 2328
rect 1902 2332 1908 2333
rect 1902 2328 1903 2332
rect 1907 2328 1908 2332
rect 1902 2327 1908 2328
rect 1982 2332 1988 2333
rect 1982 2328 1983 2332
rect 1987 2328 1988 2332
rect 1982 2327 1988 2328
rect 2062 2332 2068 2333
rect 2062 2328 2063 2332
rect 2067 2328 2068 2332
rect 2062 2327 2068 2328
rect 2142 2332 2148 2333
rect 2142 2328 2143 2332
rect 2147 2328 2148 2332
rect 2142 2327 2148 2328
rect 2502 2329 2508 2330
rect 1326 2324 1332 2325
rect 2502 2325 2503 2329
rect 2507 2325 2508 2329
rect 2502 2324 2508 2325
rect 110 2320 116 2321
rect 1286 2320 1292 2321
rect 110 2316 111 2320
rect 115 2316 116 2320
rect 110 2315 116 2316
rect 334 2319 340 2320
rect 334 2315 335 2319
rect 339 2315 340 2319
rect 334 2314 340 2315
rect 355 2319 361 2320
rect 355 2315 356 2319
rect 360 2318 361 2319
rect 386 2319 392 2320
rect 386 2318 387 2319
rect 360 2316 387 2318
rect 360 2315 361 2316
rect 355 2314 361 2315
rect 386 2315 387 2316
rect 391 2315 392 2319
rect 386 2314 392 2315
rect 406 2319 412 2320
rect 406 2315 407 2319
rect 411 2315 412 2319
rect 406 2314 412 2315
rect 427 2319 433 2320
rect 427 2315 428 2319
rect 432 2318 433 2319
rect 458 2319 464 2320
rect 458 2318 459 2319
rect 432 2316 459 2318
rect 432 2315 433 2316
rect 427 2314 433 2315
rect 458 2315 459 2316
rect 463 2315 464 2319
rect 458 2314 464 2315
rect 478 2319 484 2320
rect 478 2315 479 2319
rect 483 2315 484 2319
rect 499 2319 505 2320
rect 499 2318 500 2319
rect 478 2314 484 2315
rect 488 2316 500 2318
rect 488 2310 490 2316
rect 499 2315 500 2316
rect 504 2315 505 2319
rect 499 2314 505 2315
rect 550 2319 556 2320
rect 550 2315 551 2319
rect 555 2315 556 2319
rect 550 2314 556 2315
rect 571 2319 577 2320
rect 571 2315 572 2319
rect 576 2315 577 2319
rect 571 2314 577 2315
rect 622 2319 628 2320
rect 622 2315 623 2319
rect 627 2315 628 2319
rect 622 2314 628 2315
rect 643 2319 649 2320
rect 643 2315 644 2319
rect 648 2318 649 2319
rect 674 2319 680 2320
rect 674 2318 675 2319
rect 648 2316 675 2318
rect 648 2315 649 2316
rect 643 2314 649 2315
rect 674 2315 675 2316
rect 679 2315 680 2319
rect 674 2314 680 2315
rect 694 2319 700 2320
rect 694 2315 695 2319
rect 699 2315 700 2319
rect 694 2314 700 2315
rect 710 2319 721 2320
rect 710 2315 711 2319
rect 715 2315 716 2319
rect 720 2315 721 2319
rect 710 2314 721 2315
rect 758 2319 764 2320
rect 758 2315 759 2319
rect 763 2315 764 2319
rect 758 2314 764 2315
rect 766 2319 772 2320
rect 766 2315 767 2319
rect 771 2318 772 2319
rect 779 2319 785 2320
rect 779 2318 780 2319
rect 771 2316 780 2318
rect 771 2315 772 2316
rect 766 2314 772 2315
rect 779 2315 780 2316
rect 784 2315 785 2319
rect 779 2314 785 2315
rect 822 2319 828 2320
rect 822 2315 823 2319
rect 827 2315 828 2319
rect 822 2314 828 2315
rect 843 2319 849 2320
rect 843 2315 844 2319
rect 848 2315 849 2319
rect 843 2314 849 2315
rect 878 2319 884 2320
rect 878 2315 879 2319
rect 883 2315 884 2319
rect 899 2319 905 2320
rect 899 2318 900 2319
rect 878 2314 884 2315
rect 888 2316 900 2318
rect 319 2308 490 2310
rect 319 2302 321 2308
rect 573 2306 575 2314
rect 845 2310 847 2314
rect 460 2304 575 2306
rect 740 2308 847 2310
rect 460 2302 462 2304
rect 740 2302 742 2308
rect 888 2306 890 2316
rect 899 2315 900 2316
rect 904 2315 905 2319
rect 899 2314 905 2315
rect 942 2319 948 2320
rect 942 2315 943 2319
rect 947 2315 948 2319
rect 963 2319 969 2320
rect 963 2318 964 2319
rect 942 2314 948 2315
rect 952 2316 964 2318
rect 952 2310 954 2316
rect 963 2315 964 2316
rect 968 2315 969 2319
rect 963 2314 969 2315
rect 1006 2319 1012 2320
rect 1006 2315 1007 2319
rect 1011 2315 1012 2319
rect 1027 2319 1033 2320
rect 1027 2318 1028 2319
rect 1006 2314 1012 2315
rect 1016 2316 1028 2318
rect 804 2304 890 2306
rect 892 2308 954 2310
rect 804 2302 806 2304
rect 892 2302 894 2308
rect 1016 2306 1018 2316
rect 1027 2315 1028 2316
rect 1032 2315 1033 2319
rect 1027 2314 1033 2315
rect 1070 2319 1076 2320
rect 1070 2315 1071 2319
rect 1075 2315 1076 2319
rect 1070 2314 1076 2315
rect 1078 2319 1084 2320
rect 1078 2315 1079 2319
rect 1083 2318 1084 2319
rect 1091 2319 1097 2320
rect 1091 2318 1092 2319
rect 1083 2316 1092 2318
rect 1083 2315 1084 2316
rect 1078 2314 1084 2315
rect 1091 2315 1092 2316
rect 1096 2315 1097 2319
rect 1091 2314 1097 2315
rect 1126 2319 1132 2320
rect 1126 2315 1127 2319
rect 1131 2315 1132 2319
rect 1147 2319 1153 2320
rect 1147 2318 1148 2319
rect 1126 2314 1132 2315
rect 1136 2316 1148 2318
rect 1136 2310 1138 2316
rect 1147 2315 1148 2316
rect 1152 2315 1153 2319
rect 1147 2314 1153 2315
rect 1182 2319 1188 2320
rect 1182 2315 1183 2319
rect 1187 2315 1188 2319
rect 1203 2319 1209 2320
rect 1203 2318 1204 2319
rect 1182 2314 1188 2315
rect 1192 2316 1204 2318
rect 1192 2310 1194 2316
rect 1203 2315 1204 2316
rect 1208 2315 1209 2319
rect 1203 2314 1209 2315
rect 1238 2319 1244 2320
rect 1238 2315 1239 2319
rect 1243 2315 1244 2319
rect 1259 2319 1265 2320
rect 1259 2318 1260 2319
rect 1238 2314 1244 2315
rect 1248 2316 1260 2318
rect 924 2304 1018 2306
rect 1052 2308 1138 2310
rect 1159 2308 1194 2310
rect 924 2302 926 2304
rect 1052 2302 1054 2308
rect 1159 2306 1161 2308
rect 1248 2306 1250 2316
rect 1259 2315 1260 2316
rect 1264 2315 1265 2319
rect 1286 2316 1287 2320
rect 1291 2316 1292 2320
rect 1286 2315 1292 2316
rect 1259 2314 1265 2315
rect 1326 2312 1332 2313
rect 2502 2312 2508 2313
rect 1326 2308 1327 2312
rect 1331 2308 1332 2312
rect 1326 2307 1332 2308
rect 1486 2311 1492 2312
rect 1486 2307 1487 2311
rect 1491 2307 1492 2311
rect 1486 2306 1492 2307
rect 1507 2311 1513 2312
rect 1507 2307 1508 2311
rect 1512 2310 1513 2311
rect 1530 2311 1536 2312
rect 1530 2310 1531 2311
rect 1512 2308 1531 2310
rect 1512 2307 1513 2308
rect 1507 2306 1513 2307
rect 1530 2307 1531 2308
rect 1535 2307 1536 2311
rect 1530 2306 1536 2307
rect 1550 2311 1556 2312
rect 1550 2307 1551 2311
rect 1555 2307 1556 2311
rect 1550 2306 1556 2307
rect 1571 2311 1577 2312
rect 1571 2307 1572 2311
rect 1576 2310 1577 2311
rect 1602 2311 1608 2312
rect 1602 2310 1603 2311
rect 1576 2308 1603 2310
rect 1576 2307 1577 2308
rect 1571 2306 1577 2307
rect 1602 2307 1603 2308
rect 1607 2307 1608 2311
rect 1602 2306 1608 2307
rect 1622 2311 1628 2312
rect 1622 2307 1623 2311
rect 1627 2307 1628 2311
rect 1622 2306 1628 2307
rect 1643 2311 1649 2312
rect 1643 2307 1644 2311
rect 1648 2310 1649 2311
rect 1678 2311 1684 2312
rect 1678 2310 1679 2311
rect 1648 2308 1679 2310
rect 1648 2307 1649 2308
rect 1643 2306 1649 2307
rect 1678 2307 1679 2308
rect 1683 2307 1684 2311
rect 1678 2306 1684 2307
rect 1702 2311 1708 2312
rect 1702 2307 1703 2311
rect 1707 2307 1708 2311
rect 1702 2306 1708 2307
rect 1723 2311 1729 2312
rect 1723 2307 1724 2311
rect 1728 2310 1729 2311
rect 1754 2311 1760 2312
rect 1754 2310 1755 2311
rect 1728 2308 1755 2310
rect 1728 2307 1729 2308
rect 1723 2306 1729 2307
rect 1754 2307 1755 2308
rect 1759 2307 1760 2311
rect 1754 2306 1760 2307
rect 1774 2311 1780 2312
rect 1774 2307 1775 2311
rect 1779 2307 1780 2311
rect 1774 2306 1780 2307
rect 1782 2311 1788 2312
rect 1782 2307 1783 2311
rect 1787 2310 1788 2311
rect 1795 2311 1801 2312
rect 1795 2310 1796 2311
rect 1787 2308 1796 2310
rect 1787 2307 1788 2308
rect 1782 2306 1788 2307
rect 1795 2307 1796 2308
rect 1800 2307 1801 2311
rect 1795 2306 1801 2307
rect 1846 2311 1852 2312
rect 1846 2307 1847 2311
rect 1851 2307 1852 2311
rect 1846 2306 1852 2307
rect 1867 2311 1873 2312
rect 1867 2307 1868 2311
rect 1872 2310 1873 2311
rect 1894 2311 1900 2312
rect 1894 2310 1895 2311
rect 1872 2308 1895 2310
rect 1872 2307 1873 2308
rect 1867 2306 1873 2307
rect 1894 2307 1895 2308
rect 1899 2307 1900 2311
rect 1894 2306 1900 2307
rect 1918 2311 1924 2312
rect 1918 2307 1919 2311
rect 1923 2307 1924 2311
rect 1918 2306 1924 2307
rect 1939 2311 1945 2312
rect 1939 2307 1940 2311
rect 1944 2310 1945 2311
rect 1978 2311 1984 2312
rect 1978 2310 1979 2311
rect 1944 2308 1979 2310
rect 1944 2307 1945 2308
rect 1939 2306 1945 2307
rect 1978 2307 1979 2308
rect 1983 2307 1984 2311
rect 1978 2306 1984 2307
rect 1998 2311 2004 2312
rect 1998 2307 1999 2311
rect 2003 2307 2004 2311
rect 1998 2306 2004 2307
rect 2019 2311 2025 2312
rect 2019 2307 2020 2311
rect 2024 2310 2025 2311
rect 2058 2311 2064 2312
rect 2058 2310 2059 2311
rect 2024 2308 2059 2310
rect 2024 2307 2025 2308
rect 2019 2306 2025 2307
rect 2058 2307 2059 2308
rect 2063 2307 2064 2311
rect 2058 2306 2064 2307
rect 2078 2311 2084 2312
rect 2078 2307 2079 2311
rect 2083 2307 2084 2311
rect 2078 2306 2084 2307
rect 2099 2311 2105 2312
rect 2099 2307 2100 2311
rect 2104 2310 2105 2311
rect 2138 2311 2144 2312
rect 2138 2310 2139 2311
rect 2104 2308 2139 2310
rect 2104 2307 2105 2308
rect 2099 2306 2105 2307
rect 2138 2307 2139 2308
rect 2143 2307 2144 2311
rect 2138 2306 2144 2307
rect 2158 2311 2164 2312
rect 2158 2307 2159 2311
rect 2163 2307 2164 2311
rect 2179 2311 2185 2312
rect 2179 2310 2180 2311
rect 2158 2306 2164 2307
rect 2168 2308 2180 2310
rect 1108 2304 1161 2306
rect 1164 2304 1250 2306
rect 1108 2302 1110 2304
rect 1164 2302 1166 2304
rect 1886 2303 1892 2304
rect 315 2301 321 2302
rect 315 2297 316 2301
rect 320 2297 321 2301
rect 459 2301 465 2302
rect 315 2296 321 2297
rect 386 2299 393 2300
rect 386 2295 387 2299
rect 392 2295 393 2299
rect 459 2297 460 2301
rect 464 2297 465 2301
rect 739 2301 745 2302
rect 459 2296 465 2297
rect 531 2299 537 2300
rect 386 2294 393 2295
rect 531 2295 532 2299
rect 536 2298 537 2299
rect 542 2299 548 2300
rect 542 2298 543 2299
rect 536 2296 543 2298
rect 536 2295 537 2296
rect 531 2294 537 2295
rect 542 2295 543 2296
rect 547 2295 548 2299
rect 542 2294 548 2295
rect 603 2299 609 2300
rect 603 2295 604 2299
rect 608 2298 609 2299
rect 674 2299 681 2300
rect 608 2296 671 2298
rect 608 2295 609 2296
rect 603 2294 609 2295
rect 669 2290 671 2296
rect 674 2295 675 2299
rect 680 2295 681 2299
rect 739 2297 740 2301
rect 744 2297 745 2301
rect 739 2296 745 2297
rect 803 2301 809 2302
rect 803 2297 804 2301
rect 808 2297 809 2301
rect 803 2296 809 2297
rect 859 2301 894 2302
rect 859 2297 860 2301
rect 864 2300 894 2301
rect 923 2301 929 2302
rect 864 2297 865 2300
rect 859 2296 865 2297
rect 923 2297 924 2301
rect 928 2297 929 2301
rect 1051 2301 1057 2302
rect 923 2296 929 2297
rect 987 2299 993 2300
rect 674 2294 681 2295
rect 987 2295 988 2299
rect 992 2298 993 2299
rect 992 2296 1042 2298
rect 1051 2297 1052 2301
rect 1056 2297 1057 2301
rect 1051 2296 1057 2297
rect 1107 2301 1113 2302
rect 1107 2297 1108 2301
rect 1112 2297 1113 2301
rect 1107 2296 1113 2297
rect 1163 2301 1169 2302
rect 1163 2297 1164 2301
rect 1168 2297 1169 2301
rect 1163 2296 1169 2297
rect 1219 2299 1225 2300
rect 992 2295 993 2296
rect 987 2294 993 2295
rect 1040 2294 1042 2296
rect 1078 2295 1084 2296
rect 1078 2294 1079 2295
rect 1040 2292 1079 2294
rect 766 2291 772 2292
rect 766 2290 767 2291
rect 669 2288 767 2290
rect 766 2287 767 2288
rect 771 2287 772 2291
rect 1078 2291 1079 2292
rect 1083 2291 1084 2295
rect 1219 2295 1220 2299
rect 1224 2298 1225 2299
rect 1258 2299 1264 2300
rect 1258 2298 1259 2299
rect 1224 2296 1259 2298
rect 1224 2295 1225 2296
rect 1219 2294 1225 2295
rect 1258 2295 1259 2296
rect 1263 2295 1264 2299
rect 1886 2299 1887 2303
rect 1891 2302 1892 2303
rect 2168 2302 2170 2308
rect 2179 2307 2180 2308
rect 2184 2307 2185 2311
rect 2502 2308 2503 2312
rect 2507 2308 2508 2312
rect 2502 2307 2508 2308
rect 2179 2306 2185 2307
rect 1891 2300 2170 2302
rect 1891 2299 1892 2300
rect 1886 2298 1892 2299
rect 1258 2294 1264 2295
rect 1078 2290 1084 2291
rect 1467 2291 1473 2292
rect 766 2286 772 2287
rect 1467 2287 1468 2291
rect 1472 2290 1473 2291
rect 1522 2291 1528 2292
rect 1522 2290 1523 2291
rect 1472 2288 1523 2290
rect 1472 2287 1473 2288
rect 1467 2286 1473 2287
rect 1522 2287 1523 2288
rect 1527 2287 1528 2291
rect 1522 2286 1528 2287
rect 1530 2291 1537 2292
rect 1530 2287 1531 2291
rect 1536 2287 1537 2291
rect 1530 2286 1537 2287
rect 1602 2291 1609 2292
rect 1602 2287 1603 2291
rect 1608 2287 1609 2291
rect 1602 2286 1609 2287
rect 1678 2291 1689 2292
rect 1678 2287 1679 2291
rect 1683 2287 1684 2291
rect 1688 2287 1689 2291
rect 1678 2286 1689 2287
rect 1754 2291 1761 2292
rect 1754 2287 1755 2291
rect 1760 2287 1761 2291
rect 1754 2286 1761 2287
rect 1827 2291 1833 2292
rect 1827 2287 1828 2291
rect 1832 2290 1833 2291
rect 1862 2291 1868 2292
rect 1862 2290 1863 2291
rect 1832 2288 1863 2290
rect 1832 2287 1833 2288
rect 1827 2286 1833 2287
rect 1862 2287 1863 2288
rect 1867 2287 1868 2291
rect 1862 2286 1868 2287
rect 1894 2291 1905 2292
rect 1894 2287 1895 2291
rect 1899 2287 1900 2291
rect 1904 2287 1905 2291
rect 1894 2286 1905 2287
rect 1978 2291 1985 2292
rect 1978 2287 1979 2291
rect 1984 2287 1985 2291
rect 1978 2286 1985 2287
rect 2058 2291 2065 2292
rect 2058 2287 2059 2291
rect 2064 2287 2065 2291
rect 2058 2286 2065 2287
rect 2138 2291 2145 2292
rect 2138 2287 2139 2291
rect 2144 2287 2145 2291
rect 2138 2286 2145 2287
rect 155 2279 161 2280
rect 155 2275 156 2279
rect 160 2278 161 2279
rect 251 2279 257 2280
rect 160 2276 238 2278
rect 160 2275 161 2276
rect 155 2274 161 2275
rect 236 2266 238 2276
rect 251 2275 252 2279
rect 256 2278 257 2279
rect 355 2279 361 2280
rect 256 2276 321 2278
rect 256 2275 257 2276
rect 251 2274 257 2275
rect 319 2266 321 2276
rect 355 2275 356 2279
rect 360 2275 361 2279
rect 355 2274 361 2275
rect 458 2279 465 2280
rect 458 2275 459 2279
rect 464 2275 465 2279
rect 458 2274 465 2275
rect 502 2279 508 2280
rect 502 2275 503 2279
rect 507 2278 508 2279
rect 571 2279 577 2280
rect 571 2278 572 2279
rect 507 2276 572 2278
rect 507 2275 508 2276
rect 502 2274 508 2275
rect 571 2275 572 2276
rect 576 2275 577 2279
rect 571 2274 577 2275
rect 683 2279 689 2280
rect 683 2275 684 2279
rect 688 2278 689 2279
rect 710 2279 716 2280
rect 710 2278 711 2279
rect 688 2276 711 2278
rect 688 2275 689 2276
rect 683 2274 689 2275
rect 710 2275 711 2276
rect 715 2275 716 2279
rect 710 2274 716 2275
rect 726 2279 732 2280
rect 726 2275 727 2279
rect 731 2278 732 2279
rect 787 2279 793 2280
rect 787 2278 788 2279
rect 731 2276 788 2278
rect 731 2275 732 2276
rect 726 2274 732 2275
rect 787 2275 788 2276
rect 792 2275 793 2279
rect 787 2274 793 2275
rect 830 2279 836 2280
rect 830 2275 831 2279
rect 835 2278 836 2279
rect 891 2279 897 2280
rect 891 2278 892 2279
rect 835 2276 892 2278
rect 835 2275 836 2276
rect 830 2274 836 2275
rect 891 2275 892 2276
rect 896 2275 897 2279
rect 891 2274 897 2275
rect 995 2279 1001 2280
rect 995 2275 996 2279
rect 1000 2275 1001 2279
rect 995 2274 1001 2275
rect 1038 2279 1044 2280
rect 1038 2275 1039 2279
rect 1043 2278 1044 2279
rect 1107 2279 1113 2280
rect 1107 2278 1108 2279
rect 1043 2276 1108 2278
rect 1043 2275 1044 2276
rect 1038 2274 1044 2275
rect 1107 2275 1108 2276
rect 1112 2275 1113 2279
rect 1107 2274 1113 2275
rect 1150 2279 1156 2280
rect 1150 2275 1151 2279
rect 1155 2278 1156 2279
rect 1219 2279 1225 2280
rect 1219 2278 1220 2279
rect 1155 2276 1220 2278
rect 1155 2275 1156 2276
rect 1150 2274 1156 2275
rect 1219 2275 1220 2276
rect 1224 2275 1225 2279
rect 1219 2274 1225 2275
rect 1363 2279 1369 2280
rect 1363 2275 1364 2279
rect 1368 2278 1369 2279
rect 1398 2279 1404 2280
rect 1398 2278 1399 2279
rect 1368 2276 1399 2278
rect 1368 2275 1369 2276
rect 1363 2274 1369 2275
rect 1398 2275 1399 2276
rect 1403 2275 1404 2279
rect 1398 2274 1404 2275
rect 1406 2279 1412 2280
rect 1406 2275 1407 2279
rect 1411 2278 1412 2279
rect 1459 2279 1465 2280
rect 1459 2278 1460 2279
rect 1411 2276 1460 2278
rect 1411 2275 1412 2276
rect 1406 2274 1412 2275
rect 1459 2275 1460 2276
rect 1464 2275 1465 2279
rect 1459 2274 1465 2275
rect 1502 2279 1508 2280
rect 1502 2275 1503 2279
rect 1507 2278 1508 2279
rect 1563 2279 1569 2280
rect 1563 2278 1564 2279
rect 1507 2276 1564 2278
rect 1507 2275 1508 2276
rect 1502 2274 1508 2275
rect 1563 2275 1564 2276
rect 1568 2275 1569 2279
rect 1563 2274 1569 2275
rect 1606 2279 1612 2280
rect 1606 2275 1607 2279
rect 1611 2278 1612 2279
rect 1667 2279 1673 2280
rect 1667 2278 1668 2279
rect 1611 2276 1668 2278
rect 1611 2275 1612 2276
rect 1606 2274 1612 2275
rect 1667 2275 1668 2276
rect 1672 2275 1673 2279
rect 1667 2274 1673 2275
rect 1710 2279 1716 2280
rect 1710 2275 1711 2279
rect 1715 2278 1716 2279
rect 1771 2279 1777 2280
rect 1771 2278 1772 2279
rect 1715 2276 1772 2278
rect 1715 2275 1716 2276
rect 1710 2274 1716 2275
rect 1771 2275 1772 2276
rect 1776 2275 1777 2279
rect 1771 2274 1777 2275
rect 1883 2279 1892 2280
rect 1883 2275 1884 2279
rect 1891 2275 1892 2279
rect 1883 2274 1892 2275
rect 1926 2279 1932 2280
rect 1926 2275 1927 2279
rect 1931 2278 1932 2279
rect 1995 2279 2001 2280
rect 1995 2278 1996 2279
rect 1931 2276 1996 2278
rect 1931 2275 1932 2276
rect 1926 2274 1932 2275
rect 1995 2275 1996 2276
rect 2000 2275 2001 2279
rect 1995 2274 2001 2275
rect 2038 2279 2044 2280
rect 2038 2275 2039 2279
rect 2043 2278 2044 2279
rect 2107 2279 2113 2280
rect 2107 2278 2108 2279
rect 2043 2276 2108 2278
rect 2043 2275 2044 2276
rect 2038 2274 2044 2275
rect 2107 2275 2108 2276
rect 2112 2275 2113 2279
rect 2107 2274 2113 2275
rect 2150 2279 2156 2280
rect 2150 2275 2151 2279
rect 2155 2278 2156 2279
rect 2219 2279 2225 2280
rect 2219 2278 2220 2279
rect 2155 2276 2220 2278
rect 2155 2275 2156 2276
rect 2150 2274 2156 2275
rect 2219 2275 2220 2276
rect 2224 2275 2225 2279
rect 2219 2274 2225 2275
rect 357 2270 359 2274
rect 997 2270 999 2274
rect 1074 2271 1080 2272
rect 1074 2270 1075 2271
rect 357 2268 614 2270
rect 997 2268 1075 2270
rect 236 2264 294 2266
rect 319 2264 399 2266
rect 292 2262 294 2264
rect 397 2262 399 2264
rect 612 2262 614 2268
rect 1074 2267 1075 2268
rect 1079 2267 1080 2271
rect 1074 2266 1080 2267
rect 1522 2267 1528 2268
rect 1522 2263 1523 2267
rect 1527 2266 1528 2267
rect 1527 2264 1814 2266
rect 1527 2263 1528 2264
rect 1522 2262 1528 2263
rect 1812 2262 1814 2264
rect 174 2261 180 2262
rect 110 2260 116 2261
rect 110 2256 111 2260
rect 115 2256 116 2260
rect 174 2257 175 2261
rect 179 2257 180 2261
rect 270 2261 276 2262
rect 174 2256 180 2257
rect 182 2259 188 2260
rect 110 2255 116 2256
rect 182 2255 183 2259
rect 187 2258 188 2259
rect 195 2259 201 2260
rect 195 2258 196 2259
rect 187 2256 196 2258
rect 187 2255 188 2256
rect 182 2254 188 2255
rect 195 2255 196 2256
rect 200 2255 201 2259
rect 270 2257 271 2261
rect 275 2257 276 2261
rect 270 2256 276 2257
rect 291 2261 297 2262
rect 291 2257 292 2261
rect 296 2257 297 2261
rect 291 2256 297 2257
rect 374 2261 380 2262
rect 374 2257 375 2261
rect 379 2257 380 2261
rect 374 2256 380 2257
rect 395 2261 401 2262
rect 395 2257 396 2261
rect 400 2257 401 2261
rect 395 2256 401 2257
rect 478 2261 484 2262
rect 478 2257 479 2261
rect 483 2257 484 2261
rect 590 2261 596 2262
rect 478 2256 484 2257
rect 499 2259 508 2260
rect 195 2254 201 2255
rect 499 2255 500 2259
rect 507 2255 508 2259
rect 590 2257 591 2261
rect 595 2257 596 2261
rect 590 2256 596 2257
rect 611 2261 617 2262
rect 611 2257 612 2261
rect 616 2257 617 2261
rect 611 2256 617 2257
rect 702 2261 708 2262
rect 702 2257 703 2261
rect 707 2257 708 2261
rect 806 2261 812 2262
rect 702 2256 708 2257
rect 723 2259 732 2260
rect 499 2254 508 2255
rect 723 2255 724 2259
rect 731 2255 732 2259
rect 806 2257 807 2261
rect 811 2257 812 2261
rect 910 2261 916 2262
rect 806 2256 812 2257
rect 827 2259 836 2260
rect 723 2254 732 2255
rect 827 2255 828 2259
rect 835 2255 836 2259
rect 910 2257 911 2261
rect 915 2257 916 2261
rect 1014 2261 1020 2262
rect 910 2256 916 2257
rect 926 2259 937 2260
rect 827 2254 836 2255
rect 926 2255 927 2259
rect 931 2255 932 2259
rect 936 2255 937 2259
rect 1014 2257 1015 2261
rect 1019 2257 1020 2261
rect 1126 2261 1132 2262
rect 1014 2256 1020 2257
rect 1035 2259 1044 2260
rect 926 2254 937 2255
rect 1035 2255 1036 2259
rect 1043 2255 1044 2259
rect 1126 2257 1127 2261
rect 1131 2257 1132 2261
rect 1238 2261 1244 2262
rect 1382 2261 1388 2262
rect 1126 2256 1132 2257
rect 1147 2259 1156 2260
rect 1035 2254 1044 2255
rect 1147 2255 1148 2259
rect 1155 2255 1156 2259
rect 1238 2257 1239 2261
rect 1243 2257 1244 2261
rect 1286 2260 1292 2261
rect 1238 2256 1244 2257
rect 1258 2259 1265 2260
rect 1147 2254 1156 2255
rect 1258 2255 1259 2259
rect 1264 2255 1265 2259
rect 1286 2256 1287 2260
rect 1291 2256 1292 2260
rect 1286 2255 1292 2256
rect 1326 2260 1332 2261
rect 1326 2256 1327 2260
rect 1331 2256 1332 2260
rect 1382 2257 1383 2261
rect 1387 2257 1388 2261
rect 1478 2261 1484 2262
rect 1382 2256 1388 2257
rect 1403 2259 1412 2260
rect 1326 2255 1332 2256
rect 1403 2255 1404 2259
rect 1411 2255 1412 2259
rect 1478 2257 1479 2261
rect 1483 2257 1484 2261
rect 1582 2261 1588 2262
rect 1478 2256 1484 2257
rect 1499 2259 1508 2260
rect 1258 2254 1265 2255
rect 1403 2254 1412 2255
rect 1499 2255 1500 2259
rect 1507 2255 1508 2259
rect 1582 2257 1583 2261
rect 1587 2257 1588 2261
rect 1686 2261 1692 2262
rect 1582 2256 1588 2257
rect 1603 2259 1612 2260
rect 1499 2254 1508 2255
rect 1603 2255 1604 2259
rect 1611 2255 1612 2259
rect 1686 2257 1687 2261
rect 1691 2257 1692 2261
rect 1790 2261 1796 2262
rect 1686 2256 1692 2257
rect 1707 2259 1716 2260
rect 1603 2254 1612 2255
rect 1707 2255 1708 2259
rect 1715 2255 1716 2259
rect 1790 2257 1791 2261
rect 1795 2257 1796 2261
rect 1790 2256 1796 2257
rect 1811 2261 1817 2262
rect 1811 2257 1812 2261
rect 1816 2257 1817 2261
rect 1811 2256 1817 2257
rect 1902 2261 1908 2262
rect 1902 2257 1903 2261
rect 1907 2257 1908 2261
rect 2014 2261 2020 2262
rect 1902 2256 1908 2257
rect 1923 2259 1932 2260
rect 1707 2254 1716 2255
rect 1923 2255 1924 2259
rect 1931 2255 1932 2259
rect 2014 2257 2015 2261
rect 2019 2257 2020 2261
rect 2126 2261 2132 2262
rect 2014 2256 2020 2257
rect 2035 2259 2044 2260
rect 1923 2254 1932 2255
rect 2035 2255 2036 2259
rect 2043 2255 2044 2259
rect 2126 2257 2127 2261
rect 2131 2257 2132 2261
rect 2238 2261 2244 2262
rect 2126 2256 2132 2257
rect 2147 2259 2156 2260
rect 2035 2254 2044 2255
rect 2147 2255 2148 2259
rect 2155 2255 2156 2259
rect 2238 2257 2239 2261
rect 2243 2257 2244 2261
rect 2502 2260 2508 2261
rect 2238 2256 2244 2257
rect 2246 2259 2252 2260
rect 2147 2254 2156 2255
rect 2246 2255 2247 2259
rect 2251 2258 2252 2259
rect 2259 2259 2265 2260
rect 2259 2258 2260 2259
rect 2251 2256 2260 2258
rect 2251 2255 2252 2256
rect 2246 2254 2252 2255
rect 2259 2255 2260 2256
rect 2264 2255 2265 2259
rect 2502 2256 2503 2260
rect 2507 2256 2508 2260
rect 2502 2255 2508 2256
rect 2259 2254 2265 2255
rect 110 2243 116 2244
rect 110 2239 111 2243
rect 115 2239 116 2243
rect 1286 2243 1292 2244
rect 110 2238 116 2239
rect 158 2240 164 2241
rect 158 2236 159 2240
rect 163 2236 164 2240
rect 158 2235 164 2236
rect 254 2240 260 2241
rect 254 2236 255 2240
rect 259 2236 260 2240
rect 254 2235 260 2236
rect 358 2240 364 2241
rect 358 2236 359 2240
rect 363 2236 364 2240
rect 358 2235 364 2236
rect 462 2240 468 2241
rect 462 2236 463 2240
rect 467 2236 468 2240
rect 462 2235 468 2236
rect 574 2240 580 2241
rect 574 2236 575 2240
rect 579 2236 580 2240
rect 574 2235 580 2236
rect 686 2240 692 2241
rect 686 2236 687 2240
rect 691 2236 692 2240
rect 686 2235 692 2236
rect 790 2240 796 2241
rect 790 2236 791 2240
rect 795 2236 796 2240
rect 790 2235 796 2236
rect 894 2240 900 2241
rect 894 2236 895 2240
rect 899 2236 900 2240
rect 894 2235 900 2236
rect 998 2240 1004 2241
rect 998 2236 999 2240
rect 1003 2236 1004 2240
rect 998 2235 1004 2236
rect 1110 2240 1116 2241
rect 1110 2236 1111 2240
rect 1115 2236 1116 2240
rect 1110 2235 1116 2236
rect 1222 2240 1228 2241
rect 1222 2236 1223 2240
rect 1227 2236 1228 2240
rect 1286 2239 1287 2243
rect 1291 2239 1292 2243
rect 1286 2238 1292 2239
rect 1326 2243 1332 2244
rect 1326 2239 1327 2243
rect 1331 2239 1332 2243
rect 2502 2243 2508 2244
rect 1326 2238 1332 2239
rect 1366 2240 1372 2241
rect 1222 2235 1228 2236
rect 1366 2236 1367 2240
rect 1371 2236 1372 2240
rect 1366 2235 1372 2236
rect 1462 2240 1468 2241
rect 1462 2236 1463 2240
rect 1467 2236 1468 2240
rect 1462 2235 1468 2236
rect 1566 2240 1572 2241
rect 1566 2236 1567 2240
rect 1571 2236 1572 2240
rect 1566 2235 1572 2236
rect 1670 2240 1676 2241
rect 1670 2236 1671 2240
rect 1675 2236 1676 2240
rect 1670 2235 1676 2236
rect 1774 2240 1780 2241
rect 1774 2236 1775 2240
rect 1779 2236 1780 2240
rect 1774 2235 1780 2236
rect 1886 2240 1892 2241
rect 1886 2236 1887 2240
rect 1891 2236 1892 2240
rect 1886 2235 1892 2236
rect 1998 2240 2004 2241
rect 1998 2236 1999 2240
rect 2003 2236 2004 2240
rect 1998 2235 2004 2236
rect 2110 2240 2116 2241
rect 2110 2236 2111 2240
rect 2115 2236 2116 2240
rect 2110 2235 2116 2236
rect 2222 2240 2228 2241
rect 2222 2236 2223 2240
rect 2227 2236 2228 2240
rect 2502 2239 2503 2243
rect 2507 2239 2508 2243
rect 2502 2238 2508 2239
rect 2222 2235 2228 2236
rect 142 2228 148 2229
rect 110 2225 116 2226
rect 110 2221 111 2225
rect 115 2221 116 2225
rect 142 2224 143 2228
rect 147 2224 148 2228
rect 142 2223 148 2224
rect 230 2228 236 2229
rect 230 2224 231 2228
rect 235 2224 236 2228
rect 230 2223 236 2224
rect 318 2228 324 2229
rect 318 2224 319 2228
rect 323 2224 324 2228
rect 318 2223 324 2224
rect 414 2228 420 2229
rect 414 2224 415 2228
rect 419 2224 420 2228
rect 414 2223 420 2224
rect 518 2228 524 2229
rect 518 2224 519 2228
rect 523 2224 524 2228
rect 518 2223 524 2224
rect 622 2228 628 2229
rect 622 2224 623 2228
rect 627 2224 628 2228
rect 622 2223 628 2224
rect 726 2228 732 2229
rect 726 2224 727 2228
rect 731 2224 732 2228
rect 726 2223 732 2224
rect 830 2228 836 2229
rect 830 2224 831 2228
rect 835 2224 836 2228
rect 830 2223 836 2224
rect 934 2228 940 2229
rect 934 2224 935 2228
rect 939 2224 940 2228
rect 934 2223 940 2224
rect 1038 2228 1044 2229
rect 1038 2224 1039 2228
rect 1043 2224 1044 2228
rect 1038 2223 1044 2224
rect 1142 2228 1148 2229
rect 1142 2224 1143 2228
rect 1147 2224 1148 2228
rect 1142 2223 1148 2224
rect 1222 2228 1228 2229
rect 1222 2224 1223 2228
rect 1227 2224 1228 2228
rect 1366 2228 1372 2229
rect 1222 2223 1228 2224
rect 1286 2225 1292 2226
rect 110 2220 116 2221
rect 1286 2221 1287 2225
rect 1291 2221 1292 2225
rect 1286 2220 1292 2221
rect 1326 2225 1332 2226
rect 1326 2221 1327 2225
rect 1331 2221 1332 2225
rect 1366 2224 1367 2228
rect 1371 2224 1372 2228
rect 1366 2223 1372 2224
rect 1486 2228 1492 2229
rect 1486 2224 1487 2228
rect 1491 2224 1492 2228
rect 1486 2223 1492 2224
rect 1606 2228 1612 2229
rect 1606 2224 1607 2228
rect 1611 2224 1612 2228
rect 1606 2223 1612 2224
rect 1718 2228 1724 2229
rect 1718 2224 1719 2228
rect 1723 2224 1724 2228
rect 1718 2223 1724 2224
rect 1814 2228 1820 2229
rect 1814 2224 1815 2228
rect 1819 2224 1820 2228
rect 1814 2223 1820 2224
rect 1902 2228 1908 2229
rect 1902 2224 1903 2228
rect 1907 2224 1908 2228
rect 1902 2223 1908 2224
rect 1982 2228 1988 2229
rect 1982 2224 1983 2228
rect 1987 2224 1988 2228
rect 1982 2223 1988 2224
rect 2054 2228 2060 2229
rect 2054 2224 2055 2228
rect 2059 2224 2060 2228
rect 2054 2223 2060 2224
rect 2126 2228 2132 2229
rect 2126 2224 2127 2228
rect 2131 2224 2132 2228
rect 2126 2223 2132 2224
rect 2190 2228 2196 2229
rect 2190 2224 2191 2228
rect 2195 2224 2196 2228
rect 2190 2223 2196 2224
rect 2254 2228 2260 2229
rect 2254 2224 2255 2228
rect 2259 2224 2260 2228
rect 2254 2223 2260 2224
rect 2318 2228 2324 2229
rect 2318 2224 2319 2228
rect 2323 2224 2324 2228
rect 2318 2223 2324 2224
rect 2382 2228 2388 2229
rect 2382 2224 2383 2228
rect 2387 2224 2388 2228
rect 2382 2223 2388 2224
rect 2438 2228 2444 2229
rect 2438 2224 2439 2228
rect 2443 2224 2444 2228
rect 2438 2223 2444 2224
rect 2502 2225 2508 2226
rect 1326 2220 1332 2221
rect 2502 2221 2503 2225
rect 2507 2221 2508 2225
rect 2502 2220 2508 2221
rect 110 2208 116 2209
rect 1286 2208 1292 2209
rect 110 2204 111 2208
rect 115 2204 116 2208
rect 110 2203 116 2204
rect 158 2207 164 2208
rect 158 2203 159 2207
rect 163 2203 164 2207
rect 158 2202 164 2203
rect 179 2207 185 2208
rect 179 2203 180 2207
rect 184 2206 185 2207
rect 226 2207 232 2208
rect 226 2206 227 2207
rect 184 2204 227 2206
rect 184 2203 185 2204
rect 179 2202 185 2203
rect 226 2203 227 2204
rect 231 2203 232 2207
rect 226 2202 232 2203
rect 246 2207 252 2208
rect 246 2203 247 2207
rect 251 2203 252 2207
rect 246 2202 252 2203
rect 267 2207 273 2208
rect 267 2203 268 2207
rect 272 2206 273 2207
rect 314 2207 320 2208
rect 314 2206 315 2207
rect 272 2204 315 2206
rect 272 2203 273 2204
rect 267 2202 273 2203
rect 314 2203 315 2204
rect 319 2203 320 2207
rect 314 2202 320 2203
rect 334 2207 340 2208
rect 334 2203 335 2207
rect 339 2203 340 2207
rect 334 2202 340 2203
rect 355 2207 361 2208
rect 355 2203 356 2207
rect 360 2206 361 2207
rect 410 2207 416 2208
rect 410 2206 411 2207
rect 360 2204 411 2206
rect 360 2203 361 2204
rect 355 2202 361 2203
rect 410 2203 411 2204
rect 415 2203 416 2207
rect 410 2202 416 2203
rect 430 2207 436 2208
rect 430 2203 431 2207
rect 435 2203 436 2207
rect 430 2202 436 2203
rect 451 2207 457 2208
rect 451 2203 452 2207
rect 456 2206 457 2207
rect 514 2207 520 2208
rect 514 2206 515 2207
rect 456 2204 515 2206
rect 456 2203 457 2204
rect 451 2202 457 2203
rect 514 2203 515 2204
rect 519 2203 520 2207
rect 514 2202 520 2203
rect 534 2207 540 2208
rect 534 2203 535 2207
rect 539 2203 540 2207
rect 555 2207 561 2208
rect 555 2206 556 2207
rect 534 2202 540 2203
rect 544 2204 556 2206
rect 238 2199 244 2200
rect 238 2195 239 2199
rect 243 2198 244 2199
rect 544 2198 546 2204
rect 555 2203 556 2204
rect 560 2203 561 2207
rect 555 2202 561 2203
rect 638 2207 644 2208
rect 638 2203 639 2207
rect 643 2203 644 2207
rect 638 2202 644 2203
rect 646 2207 652 2208
rect 646 2203 647 2207
rect 651 2206 652 2207
rect 659 2207 665 2208
rect 659 2206 660 2207
rect 651 2204 660 2206
rect 651 2203 652 2204
rect 646 2202 652 2203
rect 659 2203 660 2204
rect 664 2203 665 2207
rect 659 2202 665 2203
rect 742 2207 748 2208
rect 742 2203 743 2207
rect 747 2203 748 2207
rect 742 2202 748 2203
rect 750 2207 756 2208
rect 750 2203 751 2207
rect 755 2206 756 2207
rect 763 2207 769 2208
rect 763 2206 764 2207
rect 755 2204 764 2206
rect 755 2203 756 2204
rect 750 2202 756 2203
rect 763 2203 764 2204
rect 768 2203 769 2207
rect 763 2202 769 2203
rect 846 2207 852 2208
rect 846 2203 847 2207
rect 851 2203 852 2207
rect 867 2207 873 2208
rect 867 2206 868 2207
rect 846 2202 852 2203
rect 856 2204 868 2206
rect 856 2198 858 2204
rect 867 2203 868 2204
rect 872 2203 873 2207
rect 867 2202 873 2203
rect 950 2207 956 2208
rect 950 2203 951 2207
rect 955 2203 956 2207
rect 971 2207 977 2208
rect 971 2206 972 2207
rect 950 2202 956 2203
rect 960 2204 972 2206
rect 243 2196 546 2198
rect 724 2196 858 2198
rect 243 2195 244 2196
rect 238 2194 244 2195
rect 724 2190 726 2196
rect 960 2194 962 2204
rect 971 2203 972 2204
rect 976 2203 977 2207
rect 971 2202 977 2203
rect 1054 2207 1060 2208
rect 1054 2203 1055 2207
rect 1059 2203 1060 2207
rect 1054 2202 1060 2203
rect 1074 2207 1081 2208
rect 1074 2203 1075 2207
rect 1080 2203 1081 2207
rect 1074 2202 1081 2203
rect 1158 2207 1164 2208
rect 1158 2203 1159 2207
rect 1163 2203 1164 2207
rect 1158 2202 1164 2203
rect 1179 2207 1185 2208
rect 1179 2203 1180 2207
rect 1184 2206 1185 2207
rect 1218 2207 1224 2208
rect 1218 2206 1219 2207
rect 1184 2204 1219 2206
rect 1184 2203 1185 2204
rect 1179 2202 1185 2203
rect 1218 2203 1219 2204
rect 1223 2203 1224 2207
rect 1218 2202 1224 2203
rect 1238 2207 1244 2208
rect 1238 2203 1239 2207
rect 1243 2203 1244 2207
rect 1259 2207 1265 2208
rect 1259 2206 1260 2207
rect 1238 2202 1244 2203
rect 1248 2204 1260 2206
rect 1248 2194 1250 2204
rect 1259 2203 1260 2204
rect 1264 2203 1265 2207
rect 1286 2204 1287 2208
rect 1291 2204 1292 2208
rect 1286 2203 1292 2204
rect 1326 2208 1332 2209
rect 2502 2208 2508 2209
rect 1326 2204 1327 2208
rect 1331 2204 1332 2208
rect 1326 2203 1332 2204
rect 1382 2207 1388 2208
rect 1382 2203 1383 2207
rect 1387 2203 1388 2207
rect 1259 2202 1265 2203
rect 1382 2202 1388 2203
rect 1398 2207 1409 2208
rect 1398 2203 1399 2207
rect 1403 2203 1404 2207
rect 1408 2203 1409 2207
rect 1398 2202 1409 2203
rect 1502 2207 1508 2208
rect 1502 2203 1503 2207
rect 1507 2203 1508 2207
rect 1502 2202 1508 2203
rect 1523 2207 1529 2208
rect 1523 2203 1524 2207
rect 1528 2206 1529 2207
rect 1602 2207 1608 2208
rect 1602 2206 1603 2207
rect 1528 2204 1603 2206
rect 1528 2203 1529 2204
rect 1523 2202 1529 2203
rect 1602 2203 1603 2204
rect 1607 2203 1608 2207
rect 1602 2202 1608 2203
rect 1622 2207 1628 2208
rect 1622 2203 1623 2207
rect 1627 2203 1628 2207
rect 1643 2207 1649 2208
rect 1643 2206 1644 2207
rect 1622 2202 1628 2203
rect 1632 2204 1644 2206
rect 1632 2194 1634 2204
rect 1643 2203 1644 2204
rect 1648 2203 1649 2207
rect 1643 2202 1649 2203
rect 1734 2207 1740 2208
rect 1734 2203 1735 2207
rect 1739 2203 1740 2207
rect 1734 2202 1740 2203
rect 1755 2207 1761 2208
rect 1755 2203 1756 2207
rect 1760 2206 1761 2207
rect 1810 2207 1816 2208
rect 1810 2206 1811 2207
rect 1760 2204 1811 2206
rect 1760 2203 1761 2204
rect 1755 2202 1761 2203
rect 1810 2203 1811 2204
rect 1815 2203 1816 2207
rect 1810 2202 1816 2203
rect 1830 2207 1836 2208
rect 1830 2203 1831 2207
rect 1835 2203 1836 2207
rect 1830 2202 1836 2203
rect 1851 2207 1857 2208
rect 1851 2203 1852 2207
rect 1856 2206 1857 2207
rect 1898 2207 1904 2208
rect 1898 2206 1899 2207
rect 1856 2204 1899 2206
rect 1856 2203 1857 2204
rect 1851 2202 1857 2203
rect 1898 2203 1899 2204
rect 1903 2203 1904 2207
rect 1898 2202 1904 2203
rect 1918 2207 1924 2208
rect 1918 2203 1919 2207
rect 1923 2203 1924 2207
rect 1918 2202 1924 2203
rect 1939 2207 1945 2208
rect 1939 2203 1940 2207
rect 1944 2206 1945 2207
rect 1978 2207 1984 2208
rect 1978 2206 1979 2207
rect 1944 2204 1979 2206
rect 1944 2203 1945 2204
rect 1939 2202 1945 2203
rect 1978 2203 1979 2204
rect 1983 2203 1984 2207
rect 1978 2202 1984 2203
rect 1998 2207 2004 2208
rect 1998 2203 1999 2207
rect 2003 2203 2004 2207
rect 1998 2202 2004 2203
rect 2019 2207 2025 2208
rect 2019 2203 2020 2207
rect 2024 2206 2025 2207
rect 2050 2207 2056 2208
rect 2050 2206 2051 2207
rect 2024 2204 2051 2206
rect 2024 2203 2025 2204
rect 2019 2202 2025 2203
rect 2050 2203 2051 2204
rect 2055 2203 2056 2207
rect 2050 2202 2056 2203
rect 2070 2207 2076 2208
rect 2070 2203 2071 2207
rect 2075 2203 2076 2207
rect 2070 2202 2076 2203
rect 2091 2207 2097 2208
rect 2091 2203 2092 2207
rect 2096 2206 2097 2207
rect 2122 2207 2128 2208
rect 2122 2206 2123 2207
rect 2096 2204 2123 2206
rect 2096 2203 2097 2204
rect 2091 2202 2097 2203
rect 2122 2203 2123 2204
rect 2127 2203 2128 2207
rect 2122 2202 2128 2203
rect 2142 2207 2148 2208
rect 2142 2203 2143 2207
rect 2147 2203 2148 2207
rect 2142 2202 2148 2203
rect 2163 2207 2169 2208
rect 2163 2203 2164 2207
rect 2168 2206 2169 2207
rect 2186 2207 2192 2208
rect 2186 2206 2187 2207
rect 2168 2204 2187 2206
rect 2168 2203 2169 2204
rect 2163 2202 2169 2203
rect 2186 2203 2187 2204
rect 2191 2203 2192 2207
rect 2186 2202 2192 2203
rect 2206 2207 2212 2208
rect 2206 2203 2207 2207
rect 2211 2203 2212 2207
rect 2206 2202 2212 2203
rect 2227 2207 2233 2208
rect 2227 2203 2228 2207
rect 2232 2206 2233 2207
rect 2250 2207 2256 2208
rect 2250 2206 2251 2207
rect 2232 2204 2251 2206
rect 2232 2203 2233 2204
rect 2227 2202 2233 2203
rect 2250 2203 2251 2204
rect 2255 2203 2256 2207
rect 2250 2202 2256 2203
rect 2270 2207 2276 2208
rect 2270 2203 2271 2207
rect 2275 2203 2276 2207
rect 2270 2202 2276 2203
rect 2291 2207 2297 2208
rect 2291 2203 2292 2207
rect 2296 2206 2297 2207
rect 2314 2207 2320 2208
rect 2314 2206 2315 2207
rect 2296 2204 2315 2206
rect 2296 2203 2297 2204
rect 2291 2202 2297 2203
rect 2314 2203 2315 2204
rect 2319 2203 2320 2207
rect 2314 2202 2320 2203
rect 2334 2207 2340 2208
rect 2334 2203 2335 2207
rect 2339 2203 2340 2207
rect 2334 2202 2340 2203
rect 2355 2207 2361 2208
rect 2355 2203 2356 2207
rect 2360 2206 2361 2207
rect 2378 2207 2384 2208
rect 2378 2206 2379 2207
rect 2360 2204 2379 2206
rect 2360 2203 2361 2204
rect 2355 2202 2361 2203
rect 2378 2203 2379 2204
rect 2383 2203 2384 2207
rect 2378 2202 2384 2203
rect 2398 2207 2404 2208
rect 2398 2203 2399 2207
rect 2403 2203 2404 2207
rect 2398 2202 2404 2203
rect 2419 2207 2425 2208
rect 2419 2203 2420 2207
rect 2424 2206 2425 2207
rect 2434 2207 2440 2208
rect 2434 2206 2435 2207
rect 2424 2204 2435 2206
rect 2424 2203 2425 2204
rect 2419 2202 2425 2203
rect 2434 2203 2435 2204
rect 2439 2203 2440 2207
rect 2434 2202 2440 2203
rect 2454 2207 2460 2208
rect 2454 2203 2455 2207
rect 2459 2203 2460 2207
rect 2454 2202 2460 2203
rect 2462 2207 2468 2208
rect 2462 2203 2463 2207
rect 2467 2206 2468 2207
rect 2475 2207 2481 2208
rect 2475 2206 2476 2207
rect 2467 2204 2476 2206
rect 2467 2203 2468 2204
rect 2462 2202 2468 2203
rect 2475 2203 2476 2204
rect 2480 2203 2481 2207
rect 2502 2204 2503 2208
rect 2507 2204 2508 2208
rect 2502 2203 2508 2204
rect 2475 2202 2481 2203
rect 828 2192 962 2194
rect 1036 2192 1250 2194
rect 1364 2192 1634 2194
rect 828 2190 830 2192
rect 1036 2190 1038 2192
rect 1364 2190 1366 2192
rect 723 2189 729 2190
rect 139 2187 145 2188
rect 139 2183 140 2187
rect 144 2186 145 2187
rect 182 2187 188 2188
rect 182 2186 183 2187
rect 144 2184 183 2186
rect 144 2183 145 2184
rect 139 2182 145 2183
rect 182 2183 183 2184
rect 187 2183 188 2187
rect 182 2182 188 2183
rect 226 2187 233 2188
rect 226 2183 227 2187
rect 232 2183 233 2187
rect 226 2182 233 2183
rect 314 2187 321 2188
rect 314 2183 315 2187
rect 320 2183 321 2187
rect 314 2182 321 2183
rect 410 2187 417 2188
rect 410 2183 411 2187
rect 416 2183 417 2187
rect 410 2182 417 2183
rect 514 2187 521 2188
rect 514 2183 515 2187
rect 520 2183 521 2187
rect 514 2182 521 2183
rect 619 2187 625 2188
rect 619 2183 620 2187
rect 624 2186 625 2187
rect 624 2184 694 2186
rect 723 2185 724 2189
rect 728 2185 729 2189
rect 723 2184 729 2185
rect 827 2189 833 2190
rect 827 2185 828 2189
rect 832 2185 833 2189
rect 1035 2189 1041 2190
rect 827 2184 833 2185
rect 926 2187 937 2188
rect 624 2183 625 2184
rect 619 2182 625 2183
rect 692 2182 694 2184
rect 750 2183 756 2184
rect 750 2182 751 2183
rect 692 2180 751 2182
rect 750 2179 751 2180
rect 755 2179 756 2183
rect 926 2183 927 2187
rect 931 2183 932 2187
rect 936 2183 937 2187
rect 1035 2185 1036 2189
rect 1040 2185 1041 2189
rect 1363 2189 1369 2190
rect 1035 2184 1041 2185
rect 1078 2187 1084 2188
rect 926 2182 937 2183
rect 1078 2183 1079 2187
rect 1083 2186 1084 2187
rect 1139 2187 1145 2188
rect 1139 2186 1140 2187
rect 1083 2184 1140 2186
rect 1083 2183 1084 2184
rect 1078 2182 1084 2183
rect 1139 2183 1140 2184
rect 1144 2183 1145 2187
rect 1139 2182 1145 2183
rect 1218 2187 1225 2188
rect 1218 2183 1219 2187
rect 1224 2183 1225 2187
rect 1363 2185 1364 2189
rect 1368 2185 1369 2189
rect 1363 2184 1369 2185
rect 1430 2187 1436 2188
rect 1218 2182 1225 2183
rect 1430 2183 1431 2187
rect 1435 2186 1436 2187
rect 1483 2187 1489 2188
rect 1483 2186 1484 2187
rect 1435 2184 1484 2186
rect 1435 2183 1436 2184
rect 1430 2182 1436 2183
rect 1483 2183 1484 2184
rect 1488 2183 1489 2187
rect 1483 2182 1489 2183
rect 1602 2187 1609 2188
rect 1602 2183 1603 2187
rect 1608 2183 1609 2187
rect 1602 2182 1609 2183
rect 1715 2187 1724 2188
rect 1715 2183 1716 2187
rect 1723 2183 1724 2187
rect 1715 2182 1724 2183
rect 1810 2187 1817 2188
rect 1810 2183 1811 2187
rect 1816 2183 1817 2187
rect 1810 2182 1817 2183
rect 1898 2187 1905 2188
rect 1898 2183 1899 2187
rect 1904 2183 1905 2187
rect 1898 2182 1905 2183
rect 1978 2187 1985 2188
rect 1978 2183 1979 2187
rect 1984 2183 1985 2187
rect 1978 2182 1985 2183
rect 2050 2187 2057 2188
rect 2050 2183 2051 2187
rect 2056 2183 2057 2187
rect 2050 2182 2057 2183
rect 2122 2187 2129 2188
rect 2122 2183 2123 2187
rect 2128 2183 2129 2187
rect 2122 2182 2129 2183
rect 2186 2187 2193 2188
rect 2186 2183 2187 2187
rect 2192 2183 2193 2187
rect 2186 2182 2193 2183
rect 2250 2187 2257 2188
rect 2250 2183 2251 2187
rect 2256 2183 2257 2187
rect 2250 2182 2257 2183
rect 2314 2187 2321 2188
rect 2314 2183 2315 2187
rect 2320 2183 2321 2187
rect 2314 2182 2321 2183
rect 2378 2187 2385 2188
rect 2378 2183 2379 2187
rect 2384 2183 2385 2187
rect 2378 2182 2385 2183
rect 2434 2187 2441 2188
rect 2434 2183 2435 2187
rect 2440 2183 2441 2187
rect 2434 2182 2441 2183
rect 750 2178 756 2179
rect 235 2175 244 2176
rect 235 2171 236 2175
rect 243 2171 244 2175
rect 235 2170 244 2171
rect 278 2175 284 2176
rect 278 2171 279 2175
rect 283 2174 284 2175
rect 331 2175 337 2176
rect 331 2174 332 2175
rect 283 2172 332 2174
rect 283 2171 284 2172
rect 278 2170 284 2171
rect 331 2171 332 2172
rect 336 2171 337 2175
rect 331 2170 337 2171
rect 374 2175 380 2176
rect 374 2171 375 2175
rect 379 2174 380 2175
rect 435 2175 441 2176
rect 435 2174 436 2175
rect 379 2172 436 2174
rect 379 2171 380 2172
rect 374 2170 380 2171
rect 435 2171 436 2172
rect 440 2171 441 2175
rect 435 2170 441 2171
rect 478 2175 484 2176
rect 478 2171 479 2175
rect 483 2174 484 2175
rect 539 2175 545 2176
rect 539 2174 540 2175
rect 483 2172 540 2174
rect 483 2171 484 2172
rect 478 2170 484 2171
rect 539 2171 540 2172
rect 544 2171 545 2175
rect 539 2170 545 2171
rect 643 2175 652 2176
rect 643 2171 644 2175
rect 651 2171 652 2175
rect 643 2170 652 2171
rect 686 2175 692 2176
rect 686 2171 687 2175
rect 691 2174 692 2175
rect 747 2175 753 2176
rect 747 2174 748 2175
rect 691 2172 748 2174
rect 691 2171 692 2172
rect 686 2170 692 2171
rect 747 2171 748 2172
rect 752 2171 753 2175
rect 747 2170 753 2171
rect 790 2175 796 2176
rect 790 2171 791 2175
rect 795 2174 796 2175
rect 843 2175 849 2176
rect 843 2174 844 2175
rect 795 2172 844 2174
rect 795 2171 796 2172
rect 790 2170 796 2171
rect 843 2171 844 2172
rect 848 2171 849 2175
rect 843 2170 849 2171
rect 886 2175 892 2176
rect 886 2171 887 2175
rect 891 2174 892 2175
rect 939 2175 945 2176
rect 939 2174 940 2175
rect 891 2172 940 2174
rect 891 2171 892 2172
rect 886 2170 892 2171
rect 939 2171 940 2172
rect 944 2171 945 2175
rect 939 2170 945 2171
rect 1035 2175 1041 2176
rect 1035 2171 1036 2175
rect 1040 2174 1041 2175
rect 1139 2175 1145 2176
rect 1040 2172 1102 2174
rect 1040 2171 1041 2172
rect 1035 2170 1041 2171
rect 1100 2162 1102 2172
rect 1139 2171 1140 2175
rect 1144 2174 1145 2175
rect 1219 2175 1225 2176
rect 1144 2172 1161 2174
rect 1144 2171 1145 2172
rect 1139 2170 1145 2171
rect 1159 2166 1161 2172
rect 1219 2171 1220 2175
rect 1224 2174 1225 2175
rect 1258 2175 1264 2176
rect 1258 2174 1259 2175
rect 1224 2172 1259 2174
rect 1224 2171 1225 2172
rect 1219 2170 1225 2171
rect 1258 2171 1259 2172
rect 1263 2171 1264 2175
rect 1258 2170 1264 2171
rect 1159 2164 1262 2166
rect 1100 2160 1182 2162
rect 1180 2158 1182 2160
rect 1260 2158 1262 2164
rect 254 2157 260 2158
rect 110 2156 116 2157
rect 110 2152 111 2156
rect 115 2152 116 2156
rect 254 2153 255 2157
rect 259 2153 260 2157
rect 350 2157 356 2158
rect 254 2152 260 2153
rect 275 2155 284 2156
rect 110 2151 116 2152
rect 275 2151 276 2155
rect 283 2151 284 2155
rect 350 2153 351 2157
rect 355 2153 356 2157
rect 454 2157 460 2158
rect 350 2152 356 2153
rect 371 2155 380 2156
rect 275 2150 284 2151
rect 371 2151 372 2155
rect 379 2151 380 2155
rect 454 2153 455 2157
rect 459 2153 460 2157
rect 558 2157 564 2158
rect 454 2152 460 2153
rect 475 2155 484 2156
rect 371 2150 380 2151
rect 475 2151 476 2155
rect 483 2151 484 2155
rect 558 2153 559 2157
rect 563 2153 564 2157
rect 662 2157 668 2158
rect 558 2152 564 2153
rect 566 2155 572 2156
rect 475 2150 484 2151
rect 566 2151 567 2155
rect 571 2154 572 2155
rect 579 2155 585 2156
rect 579 2154 580 2155
rect 571 2152 580 2154
rect 571 2151 572 2152
rect 566 2150 572 2151
rect 579 2151 580 2152
rect 584 2151 585 2155
rect 662 2153 663 2157
rect 667 2153 668 2157
rect 766 2157 772 2158
rect 662 2152 668 2153
rect 683 2155 692 2156
rect 579 2150 585 2151
rect 683 2151 684 2155
rect 691 2151 692 2155
rect 766 2153 767 2157
rect 771 2153 772 2157
rect 862 2157 868 2158
rect 766 2152 772 2153
rect 787 2155 796 2156
rect 683 2150 692 2151
rect 787 2151 788 2155
rect 795 2151 796 2155
rect 862 2153 863 2157
rect 867 2153 868 2157
rect 958 2157 964 2158
rect 862 2152 868 2153
rect 883 2155 892 2156
rect 787 2150 796 2151
rect 883 2151 884 2155
rect 891 2151 892 2155
rect 958 2153 959 2157
rect 963 2153 964 2157
rect 1054 2157 1060 2158
rect 958 2152 964 2153
rect 979 2155 988 2156
rect 883 2150 892 2151
rect 979 2151 980 2155
rect 987 2151 988 2155
rect 1054 2153 1055 2157
rect 1059 2153 1060 2157
rect 1158 2157 1164 2158
rect 1054 2152 1060 2153
rect 1075 2155 1084 2156
rect 979 2150 988 2151
rect 1075 2151 1076 2155
rect 1083 2151 1084 2155
rect 1158 2153 1159 2157
rect 1163 2153 1164 2157
rect 1158 2152 1164 2153
rect 1179 2157 1185 2158
rect 1179 2153 1180 2157
rect 1184 2153 1185 2157
rect 1179 2152 1185 2153
rect 1238 2157 1244 2158
rect 1238 2153 1239 2157
rect 1243 2153 1244 2157
rect 1238 2152 1244 2153
rect 1259 2157 1265 2158
rect 1259 2153 1260 2157
rect 1264 2153 1265 2157
rect 1259 2152 1265 2153
rect 1286 2156 1292 2157
rect 1286 2152 1287 2156
rect 1291 2152 1292 2156
rect 1286 2151 1292 2152
rect 1387 2155 1393 2156
rect 1387 2151 1388 2155
rect 1392 2154 1393 2155
rect 1603 2155 1609 2156
rect 1392 2152 1598 2154
rect 1392 2151 1393 2152
rect 1075 2150 1084 2151
rect 1387 2150 1393 2151
rect 1596 2142 1598 2152
rect 1603 2151 1604 2155
rect 1608 2154 1609 2155
rect 1746 2155 1752 2156
rect 1746 2154 1747 2155
rect 1608 2152 1747 2154
rect 1608 2151 1609 2152
rect 1603 2150 1609 2151
rect 1746 2151 1747 2152
rect 1751 2151 1752 2155
rect 1746 2150 1752 2151
rect 1795 2155 1801 2156
rect 1795 2151 1796 2155
rect 1800 2154 1801 2155
rect 1838 2155 1844 2156
rect 1800 2152 1834 2154
rect 1800 2151 1801 2152
rect 1795 2150 1801 2151
rect 1832 2142 1834 2152
rect 1838 2151 1839 2155
rect 1843 2154 1844 2155
rect 1971 2155 1977 2156
rect 1971 2154 1972 2155
rect 1843 2152 1972 2154
rect 1843 2151 1844 2152
rect 1838 2150 1844 2151
rect 1971 2151 1972 2152
rect 1976 2151 1977 2155
rect 1971 2150 1977 2151
rect 2139 2155 2145 2156
rect 2139 2151 2140 2155
rect 2144 2154 2145 2155
rect 2299 2155 2305 2156
rect 2144 2152 2294 2154
rect 2144 2151 2145 2152
rect 2139 2150 2145 2151
rect 2292 2142 2294 2152
rect 2299 2151 2300 2155
rect 2304 2154 2305 2155
rect 2435 2155 2441 2156
rect 2304 2152 2422 2154
rect 2304 2151 2305 2152
rect 2299 2150 2305 2151
rect 2420 2142 2422 2152
rect 2435 2151 2436 2155
rect 2440 2154 2441 2155
rect 2462 2155 2468 2156
rect 2462 2154 2463 2155
rect 2440 2152 2463 2154
rect 2440 2151 2441 2152
rect 2435 2150 2441 2151
rect 2462 2151 2463 2152
rect 2467 2151 2468 2155
rect 2462 2150 2468 2151
rect 1596 2140 1646 2142
rect 1832 2140 2182 2142
rect 2292 2140 2342 2142
rect 2420 2140 2478 2142
rect 110 2139 116 2140
rect 110 2135 111 2139
rect 115 2135 116 2139
rect 1286 2139 1292 2140
rect 110 2134 116 2135
rect 238 2136 244 2137
rect 238 2132 239 2136
rect 243 2132 244 2136
rect 238 2131 244 2132
rect 334 2136 340 2137
rect 334 2132 335 2136
rect 339 2132 340 2136
rect 334 2131 340 2132
rect 438 2136 444 2137
rect 438 2132 439 2136
rect 443 2132 444 2136
rect 438 2131 444 2132
rect 542 2136 548 2137
rect 542 2132 543 2136
rect 547 2132 548 2136
rect 542 2131 548 2132
rect 646 2136 652 2137
rect 646 2132 647 2136
rect 651 2132 652 2136
rect 646 2131 652 2132
rect 750 2136 756 2137
rect 750 2132 751 2136
rect 755 2132 756 2136
rect 750 2131 756 2132
rect 846 2136 852 2137
rect 846 2132 847 2136
rect 851 2132 852 2136
rect 846 2131 852 2132
rect 942 2136 948 2137
rect 942 2132 943 2136
rect 947 2132 948 2136
rect 942 2131 948 2132
rect 1038 2136 1044 2137
rect 1038 2132 1039 2136
rect 1043 2132 1044 2136
rect 1038 2131 1044 2132
rect 1142 2136 1148 2137
rect 1142 2132 1143 2136
rect 1147 2132 1148 2136
rect 1142 2131 1148 2132
rect 1222 2136 1228 2137
rect 1222 2132 1223 2136
rect 1227 2132 1228 2136
rect 1286 2135 1287 2139
rect 1291 2135 1292 2139
rect 1644 2138 1646 2140
rect 2180 2138 2182 2140
rect 2340 2138 2342 2140
rect 2476 2138 2478 2140
rect 1406 2137 1412 2138
rect 1286 2134 1292 2135
rect 1326 2136 1332 2137
rect 1222 2131 1228 2132
rect 1326 2132 1327 2136
rect 1331 2132 1332 2136
rect 1406 2133 1407 2137
rect 1411 2133 1412 2137
rect 1622 2137 1628 2138
rect 1406 2132 1412 2133
rect 1427 2135 1436 2136
rect 1326 2131 1332 2132
rect 1427 2131 1428 2135
rect 1435 2131 1436 2135
rect 1622 2133 1623 2137
rect 1627 2133 1628 2137
rect 1622 2132 1628 2133
rect 1643 2137 1649 2138
rect 1643 2133 1644 2137
rect 1648 2133 1649 2137
rect 1643 2132 1649 2133
rect 1814 2137 1820 2138
rect 1814 2133 1815 2137
rect 1819 2133 1820 2137
rect 1990 2137 1996 2138
rect 1814 2132 1820 2133
rect 1835 2135 1844 2136
rect 1427 2130 1436 2131
rect 1835 2131 1836 2135
rect 1843 2131 1844 2135
rect 1990 2133 1991 2137
rect 1995 2133 1996 2137
rect 2158 2137 2164 2138
rect 1990 2132 1996 2133
rect 2011 2135 2017 2136
rect 1835 2130 1844 2131
rect 2011 2131 2012 2135
rect 2016 2134 2017 2135
rect 2110 2135 2116 2136
rect 2110 2134 2111 2135
rect 2016 2132 2111 2134
rect 2016 2131 2017 2132
rect 2011 2130 2017 2131
rect 2110 2131 2111 2132
rect 2115 2131 2116 2135
rect 2158 2133 2159 2137
rect 2163 2133 2164 2137
rect 2158 2132 2164 2133
rect 2179 2137 2185 2138
rect 2179 2133 2180 2137
rect 2184 2133 2185 2137
rect 2179 2132 2185 2133
rect 2318 2137 2324 2138
rect 2318 2133 2319 2137
rect 2323 2133 2324 2137
rect 2318 2132 2324 2133
rect 2339 2137 2345 2138
rect 2339 2133 2340 2137
rect 2344 2133 2345 2137
rect 2339 2132 2345 2133
rect 2454 2137 2460 2138
rect 2454 2133 2455 2137
rect 2459 2133 2460 2137
rect 2454 2132 2460 2133
rect 2475 2137 2481 2138
rect 2475 2133 2476 2137
rect 2480 2133 2481 2137
rect 2475 2132 2481 2133
rect 2502 2136 2508 2137
rect 2502 2132 2503 2136
rect 2507 2132 2508 2136
rect 2502 2131 2508 2132
rect 2110 2130 2116 2131
rect 302 2124 308 2125
rect 110 2121 116 2122
rect 110 2117 111 2121
rect 115 2117 116 2121
rect 302 2120 303 2124
rect 307 2120 308 2124
rect 302 2119 308 2120
rect 358 2124 364 2125
rect 358 2120 359 2124
rect 363 2120 364 2124
rect 358 2119 364 2120
rect 422 2124 428 2125
rect 422 2120 423 2124
rect 427 2120 428 2124
rect 422 2119 428 2120
rect 486 2124 492 2125
rect 486 2120 487 2124
rect 491 2120 492 2124
rect 486 2119 492 2120
rect 558 2124 564 2125
rect 558 2120 559 2124
rect 563 2120 564 2124
rect 558 2119 564 2120
rect 630 2124 636 2125
rect 630 2120 631 2124
rect 635 2120 636 2124
rect 630 2119 636 2120
rect 710 2124 716 2125
rect 710 2120 711 2124
rect 715 2120 716 2124
rect 710 2119 716 2120
rect 798 2124 804 2125
rect 798 2120 799 2124
rect 803 2120 804 2124
rect 798 2119 804 2120
rect 886 2124 892 2125
rect 886 2120 887 2124
rect 891 2120 892 2124
rect 886 2119 892 2120
rect 974 2124 980 2125
rect 974 2120 975 2124
rect 979 2120 980 2124
rect 974 2119 980 2120
rect 1062 2124 1068 2125
rect 1062 2120 1063 2124
rect 1067 2120 1068 2124
rect 1062 2119 1068 2120
rect 1150 2124 1156 2125
rect 1150 2120 1151 2124
rect 1155 2120 1156 2124
rect 1150 2119 1156 2120
rect 1222 2124 1228 2125
rect 1222 2120 1223 2124
rect 1227 2120 1228 2124
rect 1222 2119 1228 2120
rect 1286 2121 1292 2122
rect 110 2116 116 2117
rect 1286 2117 1287 2121
rect 1291 2117 1292 2121
rect 1286 2116 1292 2117
rect 1326 2119 1332 2120
rect 1326 2115 1327 2119
rect 1331 2115 1332 2119
rect 2502 2119 2508 2120
rect 1326 2114 1332 2115
rect 1390 2116 1396 2117
rect 1390 2112 1391 2116
rect 1395 2112 1396 2116
rect 1390 2111 1396 2112
rect 1606 2116 1612 2117
rect 1606 2112 1607 2116
rect 1611 2112 1612 2116
rect 1606 2111 1612 2112
rect 1798 2116 1804 2117
rect 1798 2112 1799 2116
rect 1803 2112 1804 2116
rect 1798 2111 1804 2112
rect 1974 2116 1980 2117
rect 1974 2112 1975 2116
rect 1979 2112 1980 2116
rect 1974 2111 1980 2112
rect 2142 2116 2148 2117
rect 2142 2112 2143 2116
rect 2147 2112 2148 2116
rect 2142 2111 2148 2112
rect 2302 2116 2308 2117
rect 2302 2112 2303 2116
rect 2307 2112 2308 2116
rect 2302 2111 2308 2112
rect 2438 2116 2444 2117
rect 2438 2112 2439 2116
rect 2443 2112 2444 2116
rect 2502 2115 2503 2119
rect 2507 2115 2508 2119
rect 2502 2114 2508 2115
rect 2438 2111 2444 2112
rect 110 2104 116 2105
rect 1286 2104 1292 2105
rect 110 2100 111 2104
rect 115 2100 116 2104
rect 110 2099 116 2100
rect 318 2103 324 2104
rect 318 2099 319 2103
rect 323 2099 324 2103
rect 318 2098 324 2099
rect 339 2103 345 2104
rect 339 2099 340 2103
rect 344 2102 345 2103
rect 354 2103 360 2104
rect 354 2102 355 2103
rect 344 2100 355 2102
rect 344 2099 345 2100
rect 339 2098 345 2099
rect 354 2099 355 2100
rect 359 2099 360 2103
rect 354 2098 360 2099
rect 374 2103 380 2104
rect 374 2099 375 2103
rect 379 2099 380 2103
rect 374 2098 380 2099
rect 395 2103 401 2104
rect 395 2099 396 2103
rect 400 2102 401 2103
rect 418 2103 424 2104
rect 418 2102 419 2103
rect 400 2100 419 2102
rect 400 2099 401 2100
rect 395 2098 401 2099
rect 418 2099 419 2100
rect 423 2099 424 2103
rect 418 2098 424 2099
rect 438 2103 444 2104
rect 438 2099 439 2103
rect 443 2099 444 2103
rect 438 2098 444 2099
rect 459 2103 465 2104
rect 459 2099 460 2103
rect 464 2102 465 2103
rect 482 2103 488 2104
rect 482 2102 483 2103
rect 464 2100 483 2102
rect 464 2099 465 2100
rect 459 2098 465 2099
rect 482 2099 483 2100
rect 487 2099 488 2103
rect 482 2098 488 2099
rect 502 2103 508 2104
rect 502 2099 503 2103
rect 507 2099 508 2103
rect 502 2098 508 2099
rect 523 2103 529 2104
rect 523 2099 524 2103
rect 528 2102 529 2103
rect 554 2103 560 2104
rect 554 2102 555 2103
rect 528 2100 555 2102
rect 528 2099 529 2100
rect 523 2098 529 2099
rect 554 2099 555 2100
rect 559 2099 560 2103
rect 554 2098 560 2099
rect 574 2103 580 2104
rect 574 2099 575 2103
rect 579 2099 580 2103
rect 574 2098 580 2099
rect 595 2103 601 2104
rect 595 2099 596 2103
rect 600 2102 601 2103
rect 626 2103 632 2104
rect 626 2102 627 2103
rect 600 2100 627 2102
rect 600 2099 601 2100
rect 595 2098 601 2099
rect 626 2099 627 2100
rect 631 2099 632 2103
rect 626 2098 632 2099
rect 646 2103 652 2104
rect 646 2099 647 2103
rect 651 2099 652 2103
rect 646 2098 652 2099
rect 654 2103 660 2104
rect 654 2099 655 2103
rect 659 2102 660 2103
rect 667 2103 673 2104
rect 667 2102 668 2103
rect 659 2100 668 2102
rect 659 2099 660 2100
rect 654 2098 660 2099
rect 667 2099 668 2100
rect 672 2099 673 2103
rect 667 2098 673 2099
rect 726 2103 732 2104
rect 726 2099 727 2103
rect 731 2099 732 2103
rect 726 2098 732 2099
rect 747 2103 753 2104
rect 747 2099 748 2103
rect 752 2102 753 2103
rect 794 2103 800 2104
rect 794 2102 795 2103
rect 752 2100 795 2102
rect 752 2099 753 2100
rect 747 2098 753 2099
rect 794 2099 795 2100
rect 799 2099 800 2103
rect 794 2098 800 2099
rect 814 2103 820 2104
rect 814 2099 815 2103
rect 819 2099 820 2103
rect 814 2098 820 2099
rect 835 2103 844 2104
rect 835 2099 836 2103
rect 843 2099 844 2103
rect 835 2098 844 2099
rect 902 2103 908 2104
rect 902 2099 903 2103
rect 907 2099 908 2103
rect 923 2103 929 2104
rect 923 2102 924 2103
rect 902 2098 908 2099
rect 912 2100 924 2102
rect 912 2094 914 2100
rect 923 2099 924 2100
rect 928 2099 929 2103
rect 923 2098 929 2099
rect 990 2103 996 2104
rect 990 2099 991 2103
rect 995 2099 996 2103
rect 1011 2103 1017 2104
rect 1011 2102 1012 2103
rect 990 2098 996 2099
rect 1000 2100 1012 2102
rect 708 2092 914 2094
rect 566 2091 572 2092
rect 566 2090 567 2091
rect 300 2088 567 2090
rect 300 2086 302 2088
rect 566 2087 567 2088
rect 571 2087 572 2091
rect 566 2086 572 2087
rect 708 2086 710 2092
rect 1000 2090 1002 2100
rect 1011 2099 1012 2100
rect 1016 2099 1017 2103
rect 1011 2098 1017 2099
rect 1078 2103 1084 2104
rect 1078 2099 1079 2103
rect 1083 2099 1084 2103
rect 1078 2098 1084 2099
rect 1099 2103 1105 2104
rect 1099 2099 1100 2103
rect 1104 2102 1105 2103
rect 1146 2103 1152 2104
rect 1146 2102 1147 2103
rect 1104 2100 1147 2102
rect 1104 2099 1105 2100
rect 1099 2098 1105 2099
rect 1146 2099 1147 2100
rect 1151 2099 1152 2103
rect 1146 2098 1152 2099
rect 1166 2103 1172 2104
rect 1166 2099 1167 2103
rect 1171 2099 1172 2103
rect 1166 2098 1172 2099
rect 1187 2103 1193 2104
rect 1187 2099 1188 2103
rect 1192 2102 1193 2103
rect 1218 2103 1224 2104
rect 1218 2102 1219 2103
rect 1192 2100 1219 2102
rect 1192 2099 1193 2100
rect 1187 2098 1193 2099
rect 1218 2099 1219 2100
rect 1223 2099 1224 2103
rect 1218 2098 1224 2099
rect 1238 2103 1244 2104
rect 1238 2099 1239 2103
rect 1243 2099 1244 2103
rect 1238 2098 1244 2099
rect 1258 2103 1265 2104
rect 1258 2099 1259 2103
rect 1264 2099 1265 2103
rect 1286 2100 1287 2104
rect 1291 2100 1292 2104
rect 1382 2104 1388 2105
rect 1286 2099 1292 2100
rect 1326 2101 1332 2102
rect 1258 2098 1265 2099
rect 1326 2097 1327 2101
rect 1331 2097 1332 2101
rect 1382 2100 1383 2104
rect 1387 2100 1388 2104
rect 1382 2099 1388 2100
rect 1550 2104 1556 2105
rect 1550 2100 1551 2104
rect 1555 2100 1556 2104
rect 1550 2099 1556 2100
rect 1710 2104 1716 2105
rect 1710 2100 1711 2104
rect 1715 2100 1716 2104
rect 1710 2099 1716 2100
rect 1854 2104 1860 2105
rect 1854 2100 1855 2104
rect 1859 2100 1860 2104
rect 1854 2099 1860 2100
rect 1990 2104 1996 2105
rect 1990 2100 1991 2104
rect 1995 2100 1996 2104
rect 1990 2099 1996 2100
rect 2118 2104 2124 2105
rect 2118 2100 2119 2104
rect 2123 2100 2124 2104
rect 2118 2099 2124 2100
rect 2238 2104 2244 2105
rect 2238 2100 2239 2104
rect 2243 2100 2244 2104
rect 2238 2099 2244 2100
rect 2366 2104 2372 2105
rect 2366 2100 2367 2104
rect 2371 2100 2372 2104
rect 2366 2099 2372 2100
rect 2502 2101 2508 2102
rect 1326 2096 1332 2097
rect 2502 2097 2503 2101
rect 2507 2097 2508 2101
rect 2502 2096 2508 2097
rect 885 2088 1002 2090
rect 885 2086 887 2088
rect 299 2085 305 2086
rect 299 2081 300 2085
rect 304 2081 305 2085
rect 707 2085 713 2086
rect 299 2080 305 2081
rect 354 2083 361 2084
rect 354 2079 355 2083
rect 360 2079 361 2083
rect 354 2078 361 2079
rect 418 2083 425 2084
rect 418 2079 419 2083
rect 424 2079 425 2083
rect 418 2078 425 2079
rect 482 2083 489 2084
rect 482 2079 483 2083
rect 488 2079 489 2083
rect 482 2078 489 2079
rect 554 2083 561 2084
rect 554 2079 555 2083
rect 560 2079 561 2083
rect 554 2078 561 2079
rect 626 2083 633 2084
rect 626 2079 627 2083
rect 632 2079 633 2083
rect 707 2081 708 2085
rect 712 2081 713 2085
rect 883 2085 889 2086
rect 707 2080 713 2081
rect 794 2083 801 2084
rect 626 2078 633 2079
rect 794 2079 795 2083
rect 800 2079 801 2083
rect 883 2081 884 2085
rect 888 2081 889 2085
rect 1326 2084 1332 2085
rect 2502 2084 2508 2085
rect 883 2080 889 2081
rect 971 2083 977 2084
rect 794 2078 801 2079
rect 971 2079 972 2083
rect 976 2082 977 2083
rect 982 2083 988 2084
rect 982 2082 983 2083
rect 976 2080 983 2082
rect 976 2079 977 2080
rect 971 2078 977 2079
rect 982 2079 983 2080
rect 987 2079 988 2083
rect 982 2078 988 2079
rect 1059 2083 1065 2084
rect 1059 2079 1060 2083
rect 1064 2082 1065 2083
rect 1110 2083 1116 2084
rect 1110 2082 1111 2083
rect 1064 2080 1111 2082
rect 1064 2079 1065 2080
rect 1059 2078 1065 2079
rect 1110 2079 1111 2080
rect 1115 2079 1116 2083
rect 1110 2078 1116 2079
rect 1146 2083 1153 2084
rect 1146 2079 1147 2083
rect 1152 2079 1153 2083
rect 1146 2078 1153 2079
rect 1218 2083 1225 2084
rect 1218 2079 1219 2083
rect 1224 2079 1225 2083
rect 1326 2080 1327 2084
rect 1331 2080 1332 2084
rect 1326 2079 1332 2080
rect 1398 2083 1404 2084
rect 1398 2079 1399 2083
rect 1403 2079 1404 2083
rect 1218 2078 1225 2079
rect 1398 2078 1404 2079
rect 1419 2083 1425 2084
rect 1419 2079 1420 2083
rect 1424 2082 1425 2083
rect 1546 2083 1552 2084
rect 1546 2082 1547 2083
rect 1424 2080 1547 2082
rect 1424 2079 1425 2080
rect 1419 2078 1425 2079
rect 1546 2079 1547 2080
rect 1551 2079 1552 2083
rect 1546 2078 1552 2079
rect 1566 2083 1572 2084
rect 1566 2079 1567 2083
rect 1571 2079 1572 2083
rect 1566 2078 1572 2079
rect 1587 2083 1593 2084
rect 1587 2079 1588 2083
rect 1592 2082 1593 2083
rect 1706 2083 1712 2084
rect 1706 2082 1707 2083
rect 1592 2080 1707 2082
rect 1592 2079 1593 2080
rect 1587 2078 1593 2079
rect 1706 2079 1707 2080
rect 1711 2079 1712 2083
rect 1706 2078 1712 2079
rect 1726 2083 1732 2084
rect 1726 2079 1727 2083
rect 1731 2079 1732 2083
rect 1726 2078 1732 2079
rect 1746 2083 1753 2084
rect 1746 2079 1747 2083
rect 1752 2079 1753 2083
rect 1746 2078 1753 2079
rect 1870 2083 1876 2084
rect 1870 2079 1871 2083
rect 1875 2079 1876 2083
rect 1870 2078 1876 2079
rect 1891 2083 1897 2084
rect 1891 2079 1892 2083
rect 1896 2082 1897 2083
rect 1906 2083 1912 2084
rect 1906 2082 1907 2083
rect 1896 2080 1907 2082
rect 1896 2079 1897 2080
rect 1891 2078 1897 2079
rect 1906 2079 1907 2080
rect 1911 2079 1912 2083
rect 1906 2078 1912 2079
rect 2006 2083 2012 2084
rect 2006 2079 2007 2083
rect 2011 2079 2012 2083
rect 2027 2083 2033 2084
rect 2027 2082 2028 2083
rect 2006 2078 2012 2079
rect 2016 2080 2028 2082
rect 474 2075 480 2076
rect 474 2074 475 2075
rect 380 2072 475 2074
rect 380 2070 382 2072
rect 474 2071 475 2072
rect 479 2071 480 2075
rect 2016 2074 2018 2080
rect 2027 2079 2028 2080
rect 2032 2079 2033 2083
rect 2027 2078 2033 2079
rect 2134 2083 2140 2084
rect 2134 2079 2135 2083
rect 2139 2079 2140 2083
rect 2134 2078 2140 2079
rect 2155 2083 2161 2084
rect 2155 2079 2156 2083
rect 2160 2082 2161 2083
rect 2234 2083 2240 2084
rect 2234 2082 2235 2083
rect 2160 2080 2235 2082
rect 2160 2079 2161 2080
rect 2155 2078 2161 2079
rect 2234 2079 2235 2080
rect 2239 2079 2240 2083
rect 2234 2078 2240 2079
rect 2254 2083 2260 2084
rect 2254 2079 2255 2083
rect 2259 2079 2260 2083
rect 2254 2078 2260 2079
rect 2275 2083 2281 2084
rect 2275 2079 2276 2083
rect 2280 2082 2281 2083
rect 2362 2083 2368 2084
rect 2362 2082 2363 2083
rect 2280 2080 2363 2082
rect 2280 2079 2281 2080
rect 2275 2078 2281 2079
rect 2362 2079 2363 2080
rect 2367 2079 2368 2083
rect 2362 2078 2368 2079
rect 2382 2083 2388 2084
rect 2382 2079 2383 2083
rect 2387 2079 2388 2083
rect 2403 2083 2409 2084
rect 2403 2082 2404 2083
rect 2382 2078 2388 2079
rect 2392 2080 2404 2082
rect 474 2070 480 2071
rect 1852 2072 2018 2074
rect 379 2069 385 2070
rect 379 2065 380 2069
rect 384 2065 385 2069
rect 379 2064 385 2065
rect 435 2067 441 2068
rect 435 2063 436 2067
rect 440 2063 441 2067
rect 435 2062 441 2063
rect 491 2067 497 2068
rect 491 2063 492 2067
rect 496 2066 497 2067
rect 555 2067 561 2068
rect 496 2064 546 2066
rect 496 2063 497 2064
rect 491 2062 497 2063
rect 437 2054 439 2062
rect 544 2054 546 2064
rect 555 2063 556 2067
rect 560 2066 561 2067
rect 619 2067 625 2068
rect 560 2064 614 2066
rect 560 2063 561 2064
rect 555 2062 561 2063
rect 612 2054 614 2064
rect 619 2063 620 2067
rect 624 2066 625 2067
rect 654 2067 660 2068
rect 654 2066 655 2067
rect 624 2064 655 2066
rect 624 2063 625 2064
rect 619 2062 625 2063
rect 654 2063 655 2064
rect 659 2063 660 2067
rect 654 2062 660 2063
rect 691 2067 697 2068
rect 691 2063 692 2067
rect 696 2066 697 2067
rect 771 2067 777 2068
rect 696 2064 766 2066
rect 696 2063 697 2064
rect 691 2062 697 2063
rect 764 2054 766 2064
rect 771 2063 772 2067
rect 776 2063 777 2067
rect 771 2062 777 2063
rect 838 2067 849 2068
rect 838 2063 839 2067
rect 843 2063 844 2067
rect 848 2063 849 2067
rect 838 2062 849 2063
rect 903 2067 909 2068
rect 903 2063 904 2067
rect 908 2066 909 2067
rect 923 2067 929 2068
rect 923 2066 924 2067
rect 908 2064 924 2066
rect 908 2063 909 2064
rect 903 2062 909 2063
rect 923 2063 924 2064
rect 928 2063 929 2067
rect 923 2062 929 2063
rect 998 2067 1009 2068
rect 998 2063 999 2067
rect 1003 2063 1004 2067
rect 1008 2063 1009 2067
rect 998 2062 1009 2063
rect 1063 2067 1069 2068
rect 1063 2063 1064 2067
rect 1068 2066 1069 2067
rect 1083 2067 1089 2068
rect 1083 2066 1084 2067
rect 1068 2064 1084 2066
rect 1068 2063 1069 2064
rect 1063 2062 1069 2063
rect 1083 2063 1084 2064
rect 1088 2063 1089 2067
rect 1083 2062 1089 2063
rect 1126 2067 1132 2068
rect 1126 2063 1127 2067
rect 1131 2066 1132 2067
rect 1163 2067 1169 2068
rect 1163 2066 1164 2067
rect 1131 2064 1164 2066
rect 1131 2063 1132 2064
rect 1126 2062 1132 2063
rect 1163 2063 1164 2064
rect 1168 2063 1169 2067
rect 1163 2062 1169 2063
rect 1206 2067 1212 2068
rect 1206 2063 1207 2067
rect 1211 2066 1212 2067
rect 1219 2067 1225 2068
rect 1219 2066 1220 2067
rect 1211 2064 1220 2066
rect 1211 2063 1212 2064
rect 1206 2062 1212 2063
rect 1219 2063 1220 2064
rect 1224 2063 1225 2067
rect 1852 2066 1854 2072
rect 2392 2070 2394 2080
rect 2403 2079 2404 2080
rect 2408 2079 2409 2083
rect 2502 2080 2503 2084
rect 2507 2080 2508 2084
rect 2502 2079 2508 2080
rect 2403 2078 2409 2079
rect 1988 2068 2394 2070
rect 1988 2066 1990 2068
rect 1851 2065 1857 2066
rect 1219 2062 1225 2063
rect 1379 2063 1385 2064
rect 773 2058 775 2062
rect 1379 2059 1380 2063
rect 1384 2062 1385 2063
rect 1466 2063 1472 2064
rect 1466 2062 1467 2063
rect 1384 2060 1467 2062
rect 1384 2059 1385 2060
rect 1379 2058 1385 2059
rect 1466 2059 1467 2060
rect 1471 2059 1472 2063
rect 1466 2058 1472 2059
rect 1546 2063 1553 2064
rect 1546 2059 1547 2063
rect 1552 2059 1553 2063
rect 1546 2058 1553 2059
rect 1706 2063 1713 2064
rect 1706 2059 1707 2063
rect 1712 2059 1713 2063
rect 1851 2061 1852 2065
rect 1856 2061 1857 2065
rect 1851 2060 1857 2061
rect 1987 2065 1993 2066
rect 1987 2061 1988 2065
rect 1992 2061 1993 2065
rect 1987 2060 1993 2061
rect 2110 2063 2121 2064
rect 1706 2058 1713 2059
rect 2110 2059 2111 2063
rect 2115 2059 2116 2063
rect 2120 2059 2121 2063
rect 2110 2058 2121 2059
rect 2234 2063 2241 2064
rect 2234 2059 2235 2063
rect 2240 2059 2241 2063
rect 2234 2058 2241 2059
rect 2362 2063 2369 2064
rect 2362 2059 2363 2063
rect 2368 2059 2369 2063
rect 2362 2058 2369 2059
rect 773 2056 954 2058
rect 437 2052 535 2054
rect 544 2052 598 2054
rect 612 2052 662 2054
rect 764 2052 814 2054
rect 533 2050 535 2052
rect 596 2050 598 2052
rect 660 2050 662 2052
rect 812 2050 814 2052
rect 952 2050 954 2056
rect 1110 2055 1116 2056
rect 1110 2051 1111 2055
rect 1115 2054 1116 2055
rect 1115 2052 1262 2054
rect 1115 2051 1116 2052
rect 1110 2050 1116 2051
rect 1260 2050 1262 2052
rect 398 2049 404 2050
rect 110 2048 116 2049
rect 110 2044 111 2048
rect 115 2044 116 2048
rect 398 2045 399 2049
rect 403 2045 404 2049
rect 454 2049 460 2050
rect 398 2044 404 2045
rect 419 2047 425 2048
rect 110 2043 116 2044
rect 419 2043 420 2047
rect 424 2046 425 2047
rect 430 2047 436 2048
rect 430 2046 431 2047
rect 424 2044 431 2046
rect 424 2043 425 2044
rect 419 2042 425 2043
rect 430 2043 431 2044
rect 435 2043 436 2047
rect 454 2045 455 2049
rect 459 2045 460 2049
rect 510 2049 516 2050
rect 454 2044 460 2045
rect 474 2047 481 2048
rect 430 2042 436 2043
rect 474 2043 475 2047
rect 480 2043 481 2047
rect 510 2045 511 2049
rect 515 2045 516 2049
rect 510 2044 516 2045
rect 531 2049 537 2050
rect 531 2045 532 2049
rect 536 2045 537 2049
rect 531 2044 537 2045
rect 574 2049 580 2050
rect 574 2045 575 2049
rect 579 2045 580 2049
rect 574 2044 580 2045
rect 595 2049 601 2050
rect 595 2045 596 2049
rect 600 2045 601 2049
rect 595 2044 601 2045
rect 638 2049 644 2050
rect 638 2045 639 2049
rect 643 2045 644 2049
rect 638 2044 644 2045
rect 659 2049 665 2050
rect 659 2045 660 2049
rect 664 2045 665 2049
rect 659 2044 665 2045
rect 710 2049 716 2050
rect 710 2045 711 2049
rect 715 2045 716 2049
rect 790 2049 796 2050
rect 710 2044 716 2045
rect 726 2047 737 2048
rect 474 2042 481 2043
rect 726 2043 727 2047
rect 731 2043 732 2047
rect 736 2043 737 2047
rect 790 2045 791 2049
rect 795 2045 796 2049
rect 790 2044 796 2045
rect 811 2049 817 2050
rect 811 2045 812 2049
rect 816 2045 817 2049
rect 811 2044 817 2045
rect 862 2049 868 2050
rect 862 2045 863 2049
rect 867 2045 868 2049
rect 942 2049 948 2050
rect 862 2044 868 2045
rect 883 2047 889 2048
rect 726 2042 737 2043
rect 883 2043 884 2047
rect 888 2046 889 2047
rect 903 2047 909 2048
rect 903 2046 904 2047
rect 888 2044 904 2046
rect 888 2043 889 2044
rect 883 2042 889 2043
rect 903 2043 904 2044
rect 908 2043 909 2047
rect 942 2045 943 2049
rect 947 2045 948 2049
rect 952 2049 969 2050
rect 952 2048 964 2049
rect 942 2044 948 2045
rect 963 2045 964 2048
rect 968 2045 969 2049
rect 963 2044 969 2045
rect 1022 2049 1028 2050
rect 1022 2045 1023 2049
rect 1027 2045 1028 2049
rect 1102 2049 1108 2050
rect 1022 2044 1028 2045
rect 1043 2047 1049 2048
rect 903 2042 909 2043
rect 1043 2043 1044 2047
rect 1048 2046 1049 2047
rect 1063 2047 1069 2048
rect 1063 2046 1064 2047
rect 1048 2044 1064 2046
rect 1048 2043 1049 2044
rect 1043 2042 1049 2043
rect 1063 2043 1064 2044
rect 1068 2043 1069 2047
rect 1102 2045 1103 2049
rect 1107 2045 1108 2049
rect 1182 2049 1188 2050
rect 1102 2044 1108 2045
rect 1123 2047 1132 2048
rect 1063 2042 1069 2043
rect 1123 2043 1124 2047
rect 1131 2043 1132 2047
rect 1182 2045 1183 2049
rect 1187 2045 1188 2049
rect 1238 2049 1244 2050
rect 1182 2044 1188 2045
rect 1203 2047 1212 2048
rect 1123 2042 1132 2043
rect 1203 2043 1204 2047
rect 1211 2043 1212 2047
rect 1238 2045 1239 2049
rect 1243 2045 1244 2049
rect 1238 2044 1244 2045
rect 1259 2049 1265 2050
rect 1259 2045 1260 2049
rect 1264 2045 1265 2049
rect 1259 2044 1265 2045
rect 1286 2048 1292 2049
rect 1286 2044 1287 2048
rect 1291 2044 1292 2048
rect 1286 2043 1292 2044
rect 1427 2047 1433 2048
rect 1427 2043 1428 2047
rect 1432 2046 1433 2047
rect 1531 2047 1537 2048
rect 1432 2044 1526 2046
rect 1432 2043 1433 2044
rect 1203 2042 1212 2043
rect 1427 2042 1433 2043
rect 1524 2034 1526 2044
rect 1531 2043 1532 2047
rect 1536 2046 1537 2047
rect 1542 2047 1548 2048
rect 1542 2046 1543 2047
rect 1536 2044 1543 2046
rect 1536 2043 1537 2044
rect 1531 2042 1537 2043
rect 1542 2043 1543 2044
rect 1547 2043 1548 2047
rect 1542 2042 1548 2043
rect 1574 2047 1580 2048
rect 1574 2043 1575 2047
rect 1579 2046 1580 2047
rect 1635 2047 1641 2048
rect 1635 2046 1636 2047
rect 1579 2044 1636 2046
rect 1579 2043 1580 2044
rect 1574 2042 1580 2043
rect 1635 2043 1636 2044
rect 1640 2043 1641 2047
rect 1635 2042 1641 2043
rect 1731 2047 1737 2048
rect 1731 2043 1732 2047
rect 1736 2046 1737 2047
rect 1819 2047 1825 2048
rect 1736 2044 1814 2046
rect 1736 2043 1737 2044
rect 1731 2042 1737 2043
rect 1812 2034 1814 2044
rect 1819 2043 1820 2047
rect 1824 2046 1825 2047
rect 1906 2047 1913 2048
rect 1824 2044 1902 2046
rect 1824 2043 1825 2044
rect 1819 2042 1825 2043
rect 1900 2034 1902 2044
rect 1906 2043 1907 2047
rect 1912 2043 1913 2047
rect 1906 2042 1913 2043
rect 1950 2047 1956 2048
rect 1950 2043 1951 2047
rect 1955 2046 1956 2047
rect 2003 2047 2009 2048
rect 2003 2046 2004 2047
rect 1955 2044 2004 2046
rect 1955 2043 1956 2044
rect 1950 2042 1956 2043
rect 2003 2043 2004 2044
rect 2008 2043 2009 2047
rect 2003 2042 2009 2043
rect 2046 2047 2052 2048
rect 2046 2043 2047 2047
rect 2051 2046 2052 2047
rect 2099 2047 2105 2048
rect 2099 2046 2100 2047
rect 2051 2044 2100 2046
rect 2051 2043 2052 2044
rect 2046 2042 2052 2043
rect 2099 2043 2100 2044
rect 2104 2043 2105 2047
rect 2099 2042 2105 2043
rect 1524 2032 1679 2034
rect 1812 2032 1862 2034
rect 1900 2032 2142 2034
rect 110 2031 116 2032
rect 110 2027 111 2031
rect 115 2027 116 2031
rect 1286 2031 1292 2032
rect 110 2026 116 2027
rect 382 2028 388 2029
rect 382 2024 383 2028
rect 387 2024 388 2028
rect 382 2023 388 2024
rect 438 2028 444 2029
rect 438 2024 439 2028
rect 443 2024 444 2028
rect 438 2023 444 2024
rect 494 2028 500 2029
rect 494 2024 495 2028
rect 499 2024 500 2028
rect 494 2023 500 2024
rect 558 2028 564 2029
rect 558 2024 559 2028
rect 563 2024 564 2028
rect 558 2023 564 2024
rect 622 2028 628 2029
rect 622 2024 623 2028
rect 627 2024 628 2028
rect 622 2023 628 2024
rect 694 2028 700 2029
rect 694 2024 695 2028
rect 699 2024 700 2028
rect 694 2023 700 2024
rect 774 2028 780 2029
rect 774 2024 775 2028
rect 779 2024 780 2028
rect 774 2023 780 2024
rect 846 2028 852 2029
rect 846 2024 847 2028
rect 851 2024 852 2028
rect 846 2023 852 2024
rect 926 2028 932 2029
rect 926 2024 927 2028
rect 931 2024 932 2028
rect 926 2023 932 2024
rect 1006 2028 1012 2029
rect 1006 2024 1007 2028
rect 1011 2024 1012 2028
rect 1006 2023 1012 2024
rect 1086 2028 1092 2029
rect 1086 2024 1087 2028
rect 1091 2024 1092 2028
rect 1086 2023 1092 2024
rect 1166 2028 1172 2029
rect 1166 2024 1167 2028
rect 1171 2024 1172 2028
rect 1166 2023 1172 2024
rect 1222 2028 1228 2029
rect 1222 2024 1223 2028
rect 1227 2024 1228 2028
rect 1286 2027 1287 2031
rect 1291 2027 1292 2031
rect 1677 2030 1679 2032
rect 1860 2030 1862 2032
rect 2140 2030 2142 2032
rect 1446 2029 1452 2030
rect 1286 2026 1292 2027
rect 1326 2028 1332 2029
rect 1222 2023 1228 2024
rect 1326 2024 1327 2028
rect 1331 2024 1332 2028
rect 1446 2025 1447 2029
rect 1451 2025 1452 2029
rect 1550 2029 1556 2030
rect 1446 2024 1452 2025
rect 1466 2027 1473 2028
rect 1326 2023 1332 2024
rect 1466 2023 1467 2027
rect 1472 2023 1473 2027
rect 1550 2025 1551 2029
rect 1555 2025 1556 2029
rect 1654 2029 1660 2030
rect 1550 2024 1556 2025
rect 1571 2027 1580 2028
rect 1466 2022 1473 2023
rect 1571 2023 1572 2027
rect 1579 2023 1580 2027
rect 1654 2025 1655 2029
rect 1659 2025 1660 2029
rect 1654 2024 1660 2025
rect 1675 2029 1681 2030
rect 1675 2025 1676 2029
rect 1680 2025 1681 2029
rect 1675 2024 1681 2025
rect 1750 2029 1756 2030
rect 1750 2025 1751 2029
rect 1755 2025 1756 2029
rect 1838 2029 1844 2030
rect 1750 2024 1756 2025
rect 1771 2027 1780 2028
rect 1571 2022 1580 2023
rect 1771 2023 1772 2027
rect 1779 2023 1780 2027
rect 1838 2025 1839 2029
rect 1843 2025 1844 2029
rect 1838 2024 1844 2025
rect 1859 2029 1865 2030
rect 1859 2025 1860 2029
rect 1864 2025 1865 2029
rect 1859 2024 1865 2025
rect 1926 2029 1932 2030
rect 1926 2025 1927 2029
rect 1931 2025 1932 2029
rect 2022 2029 2028 2030
rect 1926 2024 1932 2025
rect 1947 2027 1956 2028
rect 1771 2022 1780 2023
rect 1947 2023 1948 2027
rect 1955 2023 1956 2027
rect 2022 2025 2023 2029
rect 2027 2025 2028 2029
rect 2118 2029 2124 2030
rect 2022 2024 2028 2025
rect 2043 2027 2052 2028
rect 1947 2022 1956 2023
rect 2043 2023 2044 2027
rect 2051 2023 2052 2027
rect 2118 2025 2119 2029
rect 2123 2025 2124 2029
rect 2118 2024 2124 2025
rect 2139 2029 2145 2030
rect 2139 2025 2140 2029
rect 2144 2025 2145 2029
rect 2139 2024 2145 2025
rect 2502 2028 2508 2029
rect 2502 2024 2503 2028
rect 2507 2024 2508 2028
rect 2502 2023 2508 2024
rect 2043 2022 2052 2023
rect 230 2012 236 2013
rect 110 2009 116 2010
rect 110 2005 111 2009
rect 115 2005 116 2009
rect 230 2008 231 2012
rect 235 2008 236 2012
rect 230 2007 236 2008
rect 286 2012 292 2013
rect 286 2008 287 2012
rect 291 2008 292 2012
rect 286 2007 292 2008
rect 358 2012 364 2013
rect 358 2008 359 2012
rect 363 2008 364 2012
rect 358 2007 364 2008
rect 438 2012 444 2013
rect 438 2008 439 2012
rect 443 2008 444 2012
rect 438 2007 444 2008
rect 534 2012 540 2013
rect 534 2008 535 2012
rect 539 2008 540 2012
rect 534 2007 540 2008
rect 630 2012 636 2013
rect 630 2008 631 2012
rect 635 2008 636 2012
rect 630 2007 636 2008
rect 734 2012 740 2013
rect 734 2008 735 2012
rect 739 2008 740 2012
rect 734 2007 740 2008
rect 846 2012 852 2013
rect 846 2008 847 2012
rect 851 2008 852 2012
rect 846 2007 852 2008
rect 958 2012 964 2013
rect 958 2008 959 2012
rect 963 2008 964 2012
rect 958 2007 964 2008
rect 1078 2012 1084 2013
rect 1078 2008 1079 2012
rect 1083 2008 1084 2012
rect 1078 2007 1084 2008
rect 1198 2012 1204 2013
rect 1198 2008 1199 2012
rect 1203 2008 1204 2012
rect 1326 2011 1332 2012
rect 1198 2007 1204 2008
rect 1286 2009 1292 2010
rect 110 2004 116 2005
rect 1286 2005 1287 2009
rect 1291 2005 1292 2009
rect 1326 2007 1327 2011
rect 1331 2007 1332 2011
rect 2502 2011 2508 2012
rect 1326 2006 1332 2007
rect 1430 2008 1436 2009
rect 1286 2004 1292 2005
rect 1430 2004 1431 2008
rect 1435 2004 1436 2008
rect 1430 2003 1436 2004
rect 1534 2008 1540 2009
rect 1534 2004 1535 2008
rect 1539 2004 1540 2008
rect 1534 2003 1540 2004
rect 1638 2008 1644 2009
rect 1638 2004 1639 2008
rect 1643 2004 1644 2008
rect 1638 2003 1644 2004
rect 1734 2008 1740 2009
rect 1734 2004 1735 2008
rect 1739 2004 1740 2008
rect 1734 2003 1740 2004
rect 1822 2008 1828 2009
rect 1822 2004 1823 2008
rect 1827 2004 1828 2008
rect 1822 2003 1828 2004
rect 1910 2008 1916 2009
rect 1910 2004 1911 2008
rect 1915 2004 1916 2008
rect 1910 2003 1916 2004
rect 2006 2008 2012 2009
rect 2006 2004 2007 2008
rect 2011 2004 2012 2008
rect 2006 2003 2012 2004
rect 2102 2008 2108 2009
rect 2102 2004 2103 2008
rect 2107 2004 2108 2008
rect 2502 2007 2503 2011
rect 2507 2007 2508 2011
rect 2502 2006 2508 2007
rect 2102 2003 2108 2004
rect 110 1992 116 1993
rect 1286 1992 1292 1993
rect 110 1988 111 1992
rect 115 1988 116 1992
rect 110 1987 116 1988
rect 246 1991 252 1992
rect 246 1987 247 1991
rect 251 1987 252 1991
rect 246 1986 252 1987
rect 267 1991 273 1992
rect 267 1987 268 1991
rect 272 1990 273 1991
rect 282 1991 288 1992
rect 282 1990 283 1991
rect 272 1988 283 1990
rect 272 1987 273 1988
rect 267 1986 273 1987
rect 282 1987 283 1988
rect 287 1987 288 1991
rect 282 1986 288 1987
rect 302 1991 308 1992
rect 302 1987 303 1991
rect 307 1987 308 1991
rect 302 1986 308 1987
rect 323 1991 329 1992
rect 323 1987 324 1991
rect 328 1990 329 1991
rect 354 1991 360 1992
rect 354 1990 355 1991
rect 328 1988 355 1990
rect 328 1987 329 1988
rect 323 1986 329 1987
rect 354 1987 355 1988
rect 359 1987 360 1991
rect 354 1986 360 1987
rect 374 1991 380 1992
rect 374 1987 375 1991
rect 379 1987 380 1991
rect 374 1986 380 1987
rect 395 1991 401 1992
rect 395 1987 396 1991
rect 400 1990 401 1991
rect 418 1991 424 1992
rect 418 1990 419 1991
rect 400 1988 419 1990
rect 400 1987 401 1988
rect 395 1986 401 1987
rect 418 1987 419 1988
rect 423 1987 424 1991
rect 418 1986 424 1987
rect 454 1991 460 1992
rect 454 1987 455 1991
rect 459 1987 460 1991
rect 454 1986 460 1987
rect 475 1991 481 1992
rect 475 1987 476 1991
rect 480 1990 481 1991
rect 530 1991 536 1992
rect 530 1990 531 1991
rect 480 1988 531 1990
rect 480 1987 481 1988
rect 475 1986 481 1987
rect 530 1987 531 1988
rect 535 1987 536 1991
rect 530 1986 536 1987
rect 550 1991 556 1992
rect 550 1987 551 1991
rect 555 1987 556 1991
rect 550 1986 556 1987
rect 571 1991 577 1992
rect 571 1987 572 1991
rect 576 1990 577 1991
rect 626 1991 632 1992
rect 626 1990 627 1991
rect 576 1988 627 1990
rect 576 1987 577 1988
rect 571 1986 577 1987
rect 626 1987 627 1988
rect 631 1987 632 1991
rect 626 1986 632 1987
rect 646 1991 652 1992
rect 646 1987 647 1991
rect 651 1987 652 1991
rect 646 1986 652 1987
rect 654 1991 660 1992
rect 654 1987 655 1991
rect 659 1990 660 1991
rect 667 1991 673 1992
rect 667 1990 668 1991
rect 659 1988 668 1990
rect 659 1987 660 1988
rect 654 1986 660 1987
rect 667 1987 668 1988
rect 672 1987 673 1991
rect 667 1986 673 1987
rect 750 1991 756 1992
rect 750 1987 751 1991
rect 755 1987 756 1991
rect 750 1986 756 1987
rect 771 1991 777 1992
rect 771 1987 772 1991
rect 776 1990 777 1991
rect 842 1991 848 1992
rect 842 1990 843 1991
rect 776 1988 843 1990
rect 776 1987 777 1988
rect 771 1986 777 1987
rect 842 1987 843 1988
rect 847 1987 848 1991
rect 842 1986 848 1987
rect 862 1991 868 1992
rect 862 1987 863 1991
rect 867 1987 868 1991
rect 862 1986 868 1987
rect 883 1991 889 1992
rect 883 1987 884 1991
rect 888 1990 889 1991
rect 898 1991 904 1992
rect 898 1990 899 1991
rect 888 1988 899 1990
rect 888 1987 889 1988
rect 883 1986 889 1987
rect 898 1987 899 1988
rect 903 1987 904 1991
rect 898 1986 904 1987
rect 974 1991 980 1992
rect 974 1987 975 1991
rect 979 1987 980 1991
rect 974 1986 980 1987
rect 995 1991 1004 1992
rect 995 1987 996 1991
rect 1003 1987 1004 1991
rect 995 1986 1004 1987
rect 1094 1991 1100 1992
rect 1094 1987 1095 1991
rect 1099 1987 1100 1991
rect 1094 1986 1100 1987
rect 1115 1991 1121 1992
rect 1115 1987 1116 1991
rect 1120 1990 1121 1991
rect 1194 1991 1200 1992
rect 1194 1990 1195 1991
rect 1120 1988 1195 1990
rect 1120 1987 1121 1988
rect 1115 1986 1121 1987
rect 1194 1987 1195 1988
rect 1199 1987 1200 1991
rect 1194 1986 1200 1987
rect 1214 1991 1220 1992
rect 1214 1987 1215 1991
rect 1219 1987 1220 1991
rect 1235 1991 1241 1992
rect 1235 1990 1236 1991
rect 1214 1986 1220 1987
rect 1224 1988 1236 1990
rect 1224 1978 1226 1988
rect 1235 1987 1236 1988
rect 1240 1987 1241 1991
rect 1286 1988 1287 1992
rect 1291 1988 1292 1992
rect 1454 1992 1460 1993
rect 1286 1987 1292 1988
rect 1326 1989 1332 1990
rect 1235 1986 1241 1987
rect 1326 1985 1327 1989
rect 1331 1985 1332 1989
rect 1454 1988 1455 1992
rect 1459 1988 1460 1992
rect 1454 1987 1460 1988
rect 1510 1992 1516 1993
rect 1510 1988 1511 1992
rect 1515 1988 1516 1992
rect 1510 1987 1516 1988
rect 1574 1992 1580 1993
rect 1574 1988 1575 1992
rect 1579 1988 1580 1992
rect 1574 1987 1580 1988
rect 1638 1992 1644 1993
rect 1638 1988 1639 1992
rect 1643 1988 1644 1992
rect 1638 1987 1644 1988
rect 1702 1992 1708 1993
rect 1702 1988 1703 1992
rect 1707 1988 1708 1992
rect 1702 1987 1708 1988
rect 1766 1992 1772 1993
rect 1766 1988 1767 1992
rect 1771 1988 1772 1992
rect 1766 1987 1772 1988
rect 1830 1992 1836 1993
rect 1830 1988 1831 1992
rect 1835 1988 1836 1992
rect 1830 1987 1836 1988
rect 1894 1992 1900 1993
rect 1894 1988 1895 1992
rect 1899 1988 1900 1992
rect 1894 1987 1900 1988
rect 1958 1992 1964 1993
rect 1958 1988 1959 1992
rect 1963 1988 1964 1992
rect 1958 1987 1964 1988
rect 2030 1992 2036 1993
rect 2030 1988 2031 1992
rect 2035 1988 2036 1992
rect 2030 1987 2036 1988
rect 2502 1989 2508 1990
rect 1326 1984 1332 1985
rect 2502 1985 2503 1989
rect 2507 1985 2508 1989
rect 2502 1984 2508 1985
rect 956 1976 1226 1978
rect 956 1974 958 1976
rect 955 1973 961 1974
rect 227 1971 236 1972
rect 227 1967 228 1971
rect 235 1967 236 1971
rect 227 1966 236 1967
rect 282 1971 289 1972
rect 282 1967 283 1971
rect 288 1967 289 1971
rect 282 1966 289 1967
rect 354 1971 361 1972
rect 354 1967 355 1971
rect 360 1967 361 1971
rect 354 1966 361 1967
rect 430 1971 441 1972
rect 430 1967 431 1971
rect 435 1967 436 1971
rect 440 1967 441 1971
rect 430 1966 441 1967
rect 530 1971 537 1972
rect 530 1967 531 1971
rect 536 1967 537 1971
rect 530 1966 537 1967
rect 626 1971 633 1972
rect 626 1967 627 1971
rect 632 1967 633 1971
rect 626 1966 633 1967
rect 726 1971 737 1972
rect 726 1967 727 1971
rect 731 1967 732 1971
rect 736 1967 737 1971
rect 726 1966 737 1967
rect 842 1971 849 1972
rect 842 1967 843 1971
rect 848 1967 849 1971
rect 955 1969 956 1973
rect 960 1969 961 1973
rect 1326 1972 1332 1973
rect 2502 1972 2508 1973
rect 955 1968 961 1969
rect 1075 1971 1081 1972
rect 842 1966 849 1967
rect 1075 1967 1076 1971
rect 1080 1970 1081 1971
rect 1114 1971 1120 1972
rect 1114 1970 1115 1971
rect 1080 1968 1115 1970
rect 1080 1967 1081 1968
rect 1075 1966 1081 1967
rect 1114 1967 1115 1968
rect 1119 1967 1120 1971
rect 1114 1966 1120 1967
rect 1194 1971 1201 1972
rect 1194 1967 1195 1971
rect 1200 1967 1201 1971
rect 1326 1968 1327 1972
rect 1331 1968 1332 1972
rect 1326 1967 1332 1968
rect 1470 1971 1476 1972
rect 1470 1967 1471 1971
rect 1475 1967 1476 1971
rect 1194 1966 1201 1967
rect 1470 1966 1476 1967
rect 1491 1971 1497 1972
rect 1491 1967 1492 1971
rect 1496 1970 1497 1971
rect 1506 1971 1512 1972
rect 1506 1970 1507 1971
rect 1496 1968 1507 1970
rect 1496 1967 1497 1968
rect 1491 1966 1497 1967
rect 1506 1967 1507 1968
rect 1511 1967 1512 1971
rect 1506 1966 1512 1967
rect 1526 1971 1532 1972
rect 1526 1967 1527 1971
rect 1531 1967 1532 1971
rect 1526 1966 1532 1967
rect 1542 1971 1553 1972
rect 1542 1967 1543 1971
rect 1547 1967 1548 1971
rect 1552 1967 1553 1971
rect 1542 1966 1553 1967
rect 1590 1971 1596 1972
rect 1590 1967 1591 1971
rect 1595 1967 1596 1971
rect 1590 1966 1596 1967
rect 1598 1971 1604 1972
rect 1598 1967 1599 1971
rect 1603 1970 1604 1971
rect 1611 1971 1617 1972
rect 1611 1970 1612 1971
rect 1603 1968 1612 1970
rect 1603 1967 1604 1968
rect 1598 1966 1604 1967
rect 1611 1967 1612 1968
rect 1616 1967 1617 1971
rect 1611 1966 1617 1967
rect 1654 1971 1660 1972
rect 1654 1967 1655 1971
rect 1659 1967 1660 1971
rect 1675 1971 1681 1972
rect 1675 1970 1676 1971
rect 1654 1966 1660 1967
rect 1664 1968 1676 1970
rect 1664 1962 1666 1968
rect 1675 1967 1676 1968
rect 1680 1967 1681 1971
rect 1675 1966 1681 1967
rect 1718 1971 1724 1972
rect 1718 1967 1719 1971
rect 1723 1967 1724 1971
rect 1739 1971 1745 1972
rect 1739 1970 1740 1971
rect 1718 1966 1724 1967
rect 1728 1968 1740 1970
rect 1572 1960 1666 1962
rect 131 1955 137 1956
rect 131 1951 132 1955
rect 136 1954 137 1955
rect 166 1955 172 1956
rect 166 1954 167 1955
rect 136 1952 167 1954
rect 136 1951 137 1952
rect 131 1950 137 1951
rect 166 1951 167 1952
rect 171 1951 172 1955
rect 166 1950 172 1951
rect 174 1955 180 1956
rect 174 1951 175 1955
rect 179 1954 180 1955
rect 195 1955 201 1956
rect 195 1954 196 1955
rect 179 1952 196 1954
rect 179 1951 180 1952
rect 174 1950 180 1951
rect 195 1951 196 1952
rect 200 1951 201 1955
rect 195 1950 201 1951
rect 238 1955 244 1956
rect 238 1951 239 1955
rect 243 1954 244 1955
rect 299 1955 305 1956
rect 299 1954 300 1955
rect 243 1952 300 1954
rect 243 1951 244 1952
rect 238 1950 244 1951
rect 299 1951 300 1952
rect 304 1951 305 1955
rect 299 1950 305 1951
rect 418 1955 425 1956
rect 418 1951 419 1955
rect 424 1951 425 1955
rect 418 1950 425 1951
rect 462 1955 468 1956
rect 462 1951 463 1955
rect 467 1954 468 1955
rect 563 1955 569 1956
rect 563 1954 564 1955
rect 467 1952 564 1954
rect 467 1951 468 1952
rect 462 1950 468 1951
rect 563 1951 564 1952
rect 568 1951 569 1955
rect 563 1950 569 1951
rect 723 1955 729 1956
rect 723 1951 724 1955
rect 728 1954 729 1955
rect 898 1955 905 1956
rect 728 1952 890 1954
rect 728 1951 729 1952
rect 723 1950 729 1951
rect 888 1942 890 1952
rect 898 1951 899 1955
rect 904 1951 905 1955
rect 898 1950 905 1951
rect 1054 1955 1060 1956
rect 1054 1951 1055 1955
rect 1059 1954 1060 1955
rect 1075 1955 1081 1956
rect 1075 1954 1076 1955
rect 1059 1952 1076 1954
rect 1059 1951 1060 1952
rect 1054 1950 1060 1951
rect 1075 1951 1076 1952
rect 1080 1951 1081 1955
rect 1572 1954 1574 1960
rect 1728 1958 1730 1968
rect 1739 1967 1740 1968
rect 1744 1967 1745 1971
rect 1739 1966 1745 1967
rect 1782 1971 1788 1972
rect 1782 1967 1783 1971
rect 1787 1967 1788 1971
rect 1782 1966 1788 1967
rect 1803 1971 1809 1972
rect 1803 1967 1804 1971
rect 1808 1970 1809 1971
rect 1826 1971 1832 1972
rect 1826 1970 1827 1971
rect 1808 1968 1827 1970
rect 1808 1967 1809 1968
rect 1803 1966 1809 1967
rect 1826 1967 1827 1968
rect 1831 1967 1832 1971
rect 1826 1966 1832 1967
rect 1846 1971 1852 1972
rect 1846 1967 1847 1971
rect 1851 1967 1852 1971
rect 1846 1966 1852 1967
rect 1867 1971 1873 1972
rect 1867 1967 1868 1971
rect 1872 1970 1873 1971
rect 1890 1971 1896 1972
rect 1890 1970 1891 1971
rect 1872 1968 1891 1970
rect 1872 1967 1873 1968
rect 1867 1966 1873 1967
rect 1890 1967 1891 1968
rect 1895 1967 1896 1971
rect 1890 1966 1896 1967
rect 1910 1971 1916 1972
rect 1910 1967 1911 1971
rect 1915 1967 1916 1971
rect 1910 1966 1916 1967
rect 1931 1971 1937 1972
rect 1931 1967 1932 1971
rect 1936 1970 1937 1971
rect 1954 1971 1960 1972
rect 1954 1970 1955 1971
rect 1936 1968 1955 1970
rect 1936 1967 1937 1968
rect 1931 1966 1937 1967
rect 1954 1967 1955 1968
rect 1959 1967 1960 1971
rect 1954 1966 1960 1967
rect 1974 1971 1980 1972
rect 1974 1967 1975 1971
rect 1979 1967 1980 1971
rect 1974 1966 1980 1967
rect 1995 1971 2001 1972
rect 1995 1967 1996 1971
rect 2000 1970 2001 1971
rect 2026 1971 2032 1972
rect 2026 1970 2027 1971
rect 2000 1968 2027 1970
rect 2000 1967 2001 1968
rect 1995 1966 2001 1967
rect 2026 1967 2027 1968
rect 2031 1967 2032 1971
rect 2026 1966 2032 1967
rect 2046 1971 2052 1972
rect 2046 1967 2047 1971
rect 2051 1967 2052 1971
rect 2046 1966 2052 1967
rect 2054 1971 2060 1972
rect 2054 1967 2055 1971
rect 2059 1970 2060 1971
rect 2067 1971 2073 1972
rect 2067 1970 2068 1971
rect 2059 1968 2068 1970
rect 2059 1967 2060 1968
rect 2054 1966 2060 1967
rect 2067 1967 2068 1968
rect 2072 1967 2073 1971
rect 2502 1968 2503 1972
rect 2507 1968 2508 1972
rect 2502 1967 2508 1968
rect 2067 1966 2073 1967
rect 1636 1956 1730 1958
rect 1636 1954 1638 1956
rect 1571 1953 1577 1954
rect 1075 1950 1081 1951
rect 1451 1951 1457 1952
rect 1451 1947 1452 1951
rect 1456 1950 1457 1951
rect 1506 1951 1513 1952
rect 1456 1948 1502 1950
rect 1456 1947 1457 1948
rect 1451 1946 1457 1947
rect 1500 1942 1502 1948
rect 1506 1947 1507 1951
rect 1512 1947 1513 1951
rect 1571 1949 1572 1953
rect 1576 1949 1577 1953
rect 1571 1948 1577 1949
rect 1635 1953 1641 1954
rect 1635 1949 1636 1953
rect 1640 1949 1641 1953
rect 1635 1948 1641 1949
rect 1699 1951 1705 1952
rect 1506 1946 1513 1947
rect 1699 1947 1700 1951
rect 1704 1950 1705 1951
rect 1710 1951 1716 1952
rect 1710 1950 1711 1951
rect 1704 1948 1711 1950
rect 1704 1947 1705 1948
rect 1699 1946 1705 1947
rect 1710 1947 1711 1948
rect 1715 1947 1716 1951
rect 1710 1946 1716 1947
rect 1763 1951 1769 1952
rect 1763 1947 1764 1951
rect 1768 1950 1769 1951
rect 1774 1951 1780 1952
rect 1774 1950 1775 1951
rect 1768 1948 1775 1950
rect 1768 1947 1769 1948
rect 1763 1946 1769 1947
rect 1774 1947 1775 1948
rect 1779 1947 1780 1951
rect 1774 1946 1780 1947
rect 1826 1951 1833 1952
rect 1826 1947 1827 1951
rect 1832 1947 1833 1951
rect 1826 1946 1833 1947
rect 1890 1951 1897 1952
rect 1890 1947 1891 1951
rect 1896 1947 1897 1951
rect 1890 1946 1897 1947
rect 1954 1951 1961 1952
rect 1954 1947 1955 1951
rect 1960 1947 1961 1951
rect 1954 1946 1961 1947
rect 2026 1951 2033 1952
rect 2026 1947 2027 1951
rect 2032 1947 2033 1951
rect 2026 1946 2033 1947
rect 1598 1943 1604 1944
rect 1598 1942 1599 1943
rect 888 1940 943 1942
rect 1500 1940 1599 1942
rect 941 1938 943 1940
rect 1598 1939 1599 1940
rect 1603 1939 1604 1943
rect 2054 1943 2060 1944
rect 2054 1942 2055 1943
rect 1598 1938 1604 1939
rect 1900 1940 2055 1942
rect 1900 1938 1902 1940
rect 2054 1939 2055 1940
rect 2059 1939 2060 1943
rect 2054 1938 2060 1939
rect 150 1937 156 1938
rect 110 1936 116 1937
rect 110 1932 111 1936
rect 115 1932 116 1936
rect 150 1933 151 1937
rect 155 1933 156 1937
rect 214 1937 220 1938
rect 150 1932 156 1933
rect 171 1935 180 1936
rect 110 1931 116 1932
rect 171 1931 172 1935
rect 179 1931 180 1935
rect 214 1933 215 1937
rect 219 1933 220 1937
rect 318 1937 324 1938
rect 214 1932 220 1933
rect 235 1935 244 1936
rect 171 1930 180 1931
rect 235 1931 236 1935
rect 243 1931 244 1935
rect 318 1933 319 1937
rect 323 1933 324 1937
rect 438 1937 444 1938
rect 318 1932 324 1933
rect 339 1935 345 1936
rect 235 1930 244 1931
rect 339 1931 340 1935
rect 344 1934 345 1935
rect 350 1935 356 1936
rect 350 1934 351 1935
rect 344 1932 351 1934
rect 344 1931 345 1932
rect 339 1930 345 1931
rect 350 1931 351 1932
rect 355 1931 356 1935
rect 438 1933 439 1937
rect 443 1933 444 1937
rect 582 1937 588 1938
rect 438 1932 444 1933
rect 459 1935 468 1936
rect 350 1930 356 1931
rect 459 1931 460 1935
rect 467 1931 468 1935
rect 582 1933 583 1937
rect 587 1933 588 1937
rect 742 1937 748 1938
rect 582 1932 588 1933
rect 602 1935 609 1936
rect 459 1930 468 1931
rect 602 1931 603 1935
rect 608 1931 609 1935
rect 742 1933 743 1937
rect 747 1933 748 1937
rect 918 1937 924 1938
rect 742 1932 748 1933
rect 750 1935 756 1936
rect 602 1930 609 1931
rect 750 1931 751 1935
rect 755 1934 756 1935
rect 763 1935 769 1936
rect 763 1934 764 1935
rect 755 1932 764 1934
rect 755 1931 756 1932
rect 750 1930 756 1931
rect 763 1931 764 1932
rect 768 1931 769 1935
rect 918 1933 919 1937
rect 923 1933 924 1937
rect 918 1932 924 1933
rect 939 1937 945 1938
rect 939 1933 940 1937
rect 944 1933 945 1937
rect 939 1932 945 1933
rect 1094 1937 1100 1938
rect 1899 1937 1905 1938
rect 1094 1933 1095 1937
rect 1099 1933 1100 1937
rect 1286 1936 1292 1937
rect 1094 1932 1100 1933
rect 1114 1935 1121 1936
rect 763 1930 769 1931
rect 1114 1931 1115 1935
rect 1120 1931 1121 1935
rect 1286 1932 1287 1936
rect 1291 1932 1292 1936
rect 1286 1931 1292 1932
rect 1547 1935 1553 1936
rect 1547 1931 1548 1935
rect 1552 1934 1553 1935
rect 1598 1935 1604 1936
rect 1552 1932 1594 1934
rect 1552 1931 1553 1932
rect 1114 1930 1121 1931
rect 1547 1930 1553 1931
rect 1592 1922 1594 1932
rect 1598 1931 1599 1935
rect 1603 1934 1604 1935
rect 1611 1935 1617 1936
rect 1611 1934 1612 1935
rect 1603 1932 1612 1934
rect 1603 1931 1604 1932
rect 1598 1930 1604 1931
rect 1611 1931 1612 1932
rect 1616 1931 1617 1935
rect 1611 1930 1617 1931
rect 1662 1935 1668 1936
rect 1662 1931 1663 1935
rect 1667 1934 1668 1935
rect 1683 1935 1689 1936
rect 1683 1934 1684 1935
rect 1667 1932 1684 1934
rect 1667 1931 1668 1932
rect 1662 1930 1668 1931
rect 1683 1931 1684 1932
rect 1688 1931 1689 1935
rect 1683 1930 1689 1931
rect 1755 1935 1761 1936
rect 1755 1931 1756 1935
rect 1760 1934 1761 1935
rect 1766 1935 1772 1936
rect 1766 1934 1767 1935
rect 1760 1932 1767 1934
rect 1760 1931 1761 1932
rect 1755 1930 1761 1931
rect 1766 1931 1767 1932
rect 1771 1931 1772 1935
rect 1766 1930 1772 1931
rect 1814 1935 1820 1936
rect 1814 1931 1815 1935
rect 1819 1934 1820 1935
rect 1827 1935 1833 1936
rect 1827 1934 1828 1935
rect 1819 1932 1828 1934
rect 1819 1931 1820 1932
rect 1814 1930 1820 1931
rect 1827 1931 1828 1932
rect 1832 1931 1833 1935
rect 1899 1933 1900 1937
rect 1904 1933 1905 1937
rect 1899 1932 1905 1933
rect 1942 1935 1948 1936
rect 1827 1930 1833 1931
rect 1942 1931 1943 1935
rect 1947 1934 1948 1935
rect 1979 1935 1985 1936
rect 1979 1934 1980 1935
rect 1947 1932 1980 1934
rect 1947 1931 1948 1932
rect 1942 1930 1948 1931
rect 1979 1931 1980 1932
rect 1984 1931 1985 1935
rect 1979 1930 1985 1931
rect 2022 1935 2028 1936
rect 2022 1931 2023 1935
rect 2027 1934 2028 1935
rect 2067 1935 2073 1936
rect 2067 1934 2068 1935
rect 2027 1932 2068 1934
rect 2027 1931 2028 1932
rect 2022 1930 2028 1931
rect 2067 1931 2068 1932
rect 2072 1931 2073 1935
rect 2067 1930 2073 1931
rect 2110 1935 2116 1936
rect 2110 1931 2111 1935
rect 2115 1934 2116 1935
rect 2163 1935 2169 1936
rect 2163 1934 2164 1935
rect 2115 1932 2164 1934
rect 2115 1931 2116 1932
rect 2110 1930 2116 1931
rect 2163 1931 2164 1932
rect 2168 1931 2169 1935
rect 2163 1930 2169 1931
rect 2206 1935 2212 1936
rect 2206 1931 2207 1935
rect 2211 1934 2212 1935
rect 2259 1935 2265 1936
rect 2259 1934 2260 1935
rect 2211 1932 2260 1934
rect 2211 1931 2212 1932
rect 2206 1930 2212 1931
rect 2259 1931 2260 1932
rect 2264 1931 2265 1935
rect 2259 1930 2265 1931
rect 2355 1935 2361 1936
rect 2355 1931 2356 1935
rect 2360 1934 2361 1935
rect 2398 1935 2404 1936
rect 2360 1932 2394 1934
rect 2360 1931 2361 1932
rect 2355 1930 2361 1931
rect 2392 1926 2394 1932
rect 2398 1931 2399 1935
rect 2403 1934 2404 1935
rect 2435 1935 2441 1936
rect 2435 1934 2436 1935
rect 2403 1932 2436 1934
rect 2403 1931 2404 1932
rect 2398 1930 2404 1931
rect 2435 1931 2436 1932
rect 2440 1931 2441 1935
rect 2435 1930 2441 1931
rect 2418 1927 2424 1928
rect 2418 1926 2419 1927
rect 2392 1924 2419 1926
rect 2418 1923 2419 1924
rect 2423 1923 2424 1927
rect 2418 1922 2424 1923
rect 1592 1920 1870 1922
rect 110 1919 116 1920
rect 110 1915 111 1919
rect 115 1915 116 1919
rect 1286 1919 1292 1920
rect 110 1914 116 1915
rect 134 1916 140 1917
rect 134 1912 135 1916
rect 139 1912 140 1916
rect 134 1911 140 1912
rect 198 1916 204 1917
rect 198 1912 199 1916
rect 203 1912 204 1916
rect 198 1911 204 1912
rect 302 1916 308 1917
rect 302 1912 303 1916
rect 307 1912 308 1916
rect 302 1911 308 1912
rect 422 1916 428 1917
rect 422 1912 423 1916
rect 427 1912 428 1916
rect 422 1911 428 1912
rect 566 1916 572 1917
rect 566 1912 567 1916
rect 571 1912 572 1916
rect 566 1911 572 1912
rect 726 1916 732 1917
rect 726 1912 727 1916
rect 731 1912 732 1916
rect 726 1911 732 1912
rect 902 1916 908 1917
rect 902 1912 903 1916
rect 907 1912 908 1916
rect 902 1911 908 1912
rect 1078 1916 1084 1917
rect 1078 1912 1079 1916
rect 1083 1912 1084 1916
rect 1286 1915 1287 1919
rect 1291 1915 1292 1919
rect 1868 1918 1870 1920
rect 1566 1917 1572 1918
rect 1286 1914 1292 1915
rect 1326 1916 1332 1917
rect 1078 1911 1084 1912
rect 1326 1912 1327 1916
rect 1331 1912 1332 1916
rect 1566 1913 1567 1917
rect 1571 1913 1572 1917
rect 1630 1917 1636 1918
rect 1566 1912 1572 1913
rect 1587 1915 1593 1916
rect 1326 1911 1332 1912
rect 1587 1911 1588 1915
rect 1592 1914 1593 1915
rect 1598 1915 1604 1916
rect 1598 1914 1599 1915
rect 1592 1912 1599 1914
rect 1592 1911 1593 1912
rect 1587 1910 1593 1911
rect 1598 1911 1599 1912
rect 1603 1911 1604 1915
rect 1630 1913 1631 1917
rect 1635 1913 1636 1917
rect 1702 1917 1708 1918
rect 1630 1912 1636 1913
rect 1651 1915 1657 1916
rect 1598 1910 1604 1911
rect 1651 1911 1652 1915
rect 1656 1914 1657 1915
rect 1662 1915 1668 1916
rect 1662 1914 1663 1915
rect 1656 1912 1663 1914
rect 1656 1911 1657 1912
rect 1651 1910 1657 1911
rect 1662 1911 1663 1912
rect 1667 1911 1668 1915
rect 1702 1913 1703 1917
rect 1707 1913 1708 1917
rect 1774 1917 1780 1918
rect 1702 1912 1708 1913
rect 1710 1915 1716 1916
rect 1662 1910 1668 1911
rect 1710 1911 1711 1915
rect 1715 1914 1716 1915
rect 1723 1915 1729 1916
rect 1723 1914 1724 1915
rect 1715 1912 1724 1914
rect 1715 1911 1716 1912
rect 1710 1910 1716 1911
rect 1723 1911 1724 1912
rect 1728 1911 1729 1915
rect 1774 1913 1775 1917
rect 1779 1913 1780 1917
rect 1846 1917 1852 1918
rect 1774 1912 1780 1913
rect 1795 1915 1801 1916
rect 1723 1910 1729 1911
rect 1795 1911 1796 1915
rect 1800 1914 1801 1915
rect 1814 1915 1820 1916
rect 1814 1914 1815 1915
rect 1800 1912 1815 1914
rect 1800 1911 1801 1912
rect 1795 1910 1801 1911
rect 1814 1911 1815 1912
rect 1819 1911 1820 1915
rect 1846 1913 1847 1917
rect 1851 1913 1852 1917
rect 1846 1912 1852 1913
rect 1867 1917 1873 1918
rect 1867 1913 1868 1917
rect 1872 1913 1873 1917
rect 1867 1912 1873 1913
rect 1918 1917 1924 1918
rect 1918 1913 1919 1917
rect 1923 1913 1924 1917
rect 1998 1917 2004 1918
rect 1918 1912 1924 1913
rect 1939 1915 1948 1916
rect 1814 1910 1820 1911
rect 1939 1911 1940 1915
rect 1947 1911 1948 1915
rect 1998 1913 1999 1917
rect 2003 1913 2004 1917
rect 2086 1917 2092 1918
rect 1998 1912 2004 1913
rect 2019 1915 2028 1916
rect 1939 1910 1948 1911
rect 2019 1911 2020 1915
rect 2027 1911 2028 1915
rect 2086 1913 2087 1917
rect 2091 1913 2092 1917
rect 2182 1917 2188 1918
rect 2086 1912 2092 1913
rect 2107 1915 2116 1916
rect 2019 1910 2028 1911
rect 2107 1911 2108 1915
rect 2115 1911 2116 1915
rect 2182 1913 2183 1917
rect 2187 1913 2188 1917
rect 2278 1917 2284 1918
rect 2182 1912 2188 1913
rect 2203 1915 2212 1916
rect 2107 1910 2116 1911
rect 2203 1911 2204 1915
rect 2211 1911 2212 1915
rect 2278 1913 2279 1917
rect 2283 1913 2284 1917
rect 2374 1917 2380 1918
rect 2278 1912 2284 1913
rect 2286 1915 2292 1916
rect 2203 1910 2212 1911
rect 2286 1911 2287 1915
rect 2291 1914 2292 1915
rect 2299 1915 2305 1916
rect 2299 1914 2300 1915
rect 2291 1912 2300 1914
rect 2291 1911 2292 1912
rect 2286 1910 2292 1911
rect 2299 1911 2300 1912
rect 2304 1911 2305 1915
rect 2374 1913 2375 1917
rect 2379 1913 2380 1917
rect 2454 1917 2460 1918
rect 2374 1912 2380 1913
rect 2395 1915 2404 1916
rect 2299 1910 2305 1911
rect 2395 1911 2396 1915
rect 2403 1911 2404 1915
rect 2454 1913 2455 1917
rect 2459 1913 2460 1917
rect 2502 1916 2508 1917
rect 2454 1912 2460 1913
rect 2470 1915 2481 1916
rect 2395 1910 2404 1911
rect 2470 1911 2471 1915
rect 2475 1911 2476 1915
rect 2480 1911 2481 1915
rect 2502 1912 2503 1916
rect 2507 1912 2508 1916
rect 2502 1911 2508 1912
rect 2470 1910 2481 1911
rect 1326 1899 1332 1900
rect 134 1896 140 1897
rect 110 1893 116 1894
rect 110 1889 111 1893
rect 115 1889 116 1893
rect 134 1892 135 1896
rect 139 1892 140 1896
rect 134 1891 140 1892
rect 190 1896 196 1897
rect 190 1892 191 1896
rect 195 1892 196 1896
rect 190 1891 196 1892
rect 270 1896 276 1897
rect 270 1892 271 1896
rect 275 1892 276 1896
rect 270 1891 276 1892
rect 358 1896 364 1897
rect 358 1892 359 1896
rect 363 1892 364 1896
rect 358 1891 364 1892
rect 454 1896 460 1897
rect 454 1892 455 1896
rect 459 1892 460 1896
rect 454 1891 460 1892
rect 542 1896 548 1897
rect 542 1892 543 1896
rect 547 1892 548 1896
rect 542 1891 548 1892
rect 630 1896 636 1897
rect 630 1892 631 1896
rect 635 1892 636 1896
rect 630 1891 636 1892
rect 718 1896 724 1897
rect 718 1892 719 1896
rect 723 1892 724 1896
rect 718 1891 724 1892
rect 798 1896 804 1897
rect 798 1892 799 1896
rect 803 1892 804 1896
rect 798 1891 804 1892
rect 870 1896 876 1897
rect 870 1892 871 1896
rect 875 1892 876 1896
rect 870 1891 876 1892
rect 942 1896 948 1897
rect 942 1892 943 1896
rect 947 1892 948 1896
rect 942 1891 948 1892
rect 1014 1896 1020 1897
rect 1014 1892 1015 1896
rect 1019 1892 1020 1896
rect 1014 1891 1020 1892
rect 1086 1896 1092 1897
rect 1086 1892 1087 1896
rect 1091 1892 1092 1896
rect 1086 1891 1092 1892
rect 1158 1896 1164 1897
rect 1158 1892 1159 1896
rect 1163 1892 1164 1896
rect 1326 1895 1327 1899
rect 1331 1895 1332 1899
rect 2502 1899 2508 1900
rect 1326 1894 1332 1895
rect 1550 1896 1556 1897
rect 1158 1891 1164 1892
rect 1286 1893 1292 1894
rect 110 1888 116 1889
rect 1286 1889 1287 1893
rect 1291 1889 1292 1893
rect 1550 1892 1551 1896
rect 1555 1892 1556 1896
rect 1550 1891 1556 1892
rect 1614 1896 1620 1897
rect 1614 1892 1615 1896
rect 1619 1892 1620 1896
rect 1614 1891 1620 1892
rect 1686 1896 1692 1897
rect 1686 1892 1687 1896
rect 1691 1892 1692 1896
rect 1686 1891 1692 1892
rect 1758 1896 1764 1897
rect 1758 1892 1759 1896
rect 1763 1892 1764 1896
rect 1758 1891 1764 1892
rect 1830 1896 1836 1897
rect 1830 1892 1831 1896
rect 1835 1892 1836 1896
rect 1830 1891 1836 1892
rect 1902 1896 1908 1897
rect 1902 1892 1903 1896
rect 1907 1892 1908 1896
rect 1902 1891 1908 1892
rect 1982 1896 1988 1897
rect 1982 1892 1983 1896
rect 1987 1892 1988 1896
rect 1982 1891 1988 1892
rect 2070 1896 2076 1897
rect 2070 1892 2071 1896
rect 2075 1892 2076 1896
rect 2070 1891 2076 1892
rect 2166 1896 2172 1897
rect 2166 1892 2167 1896
rect 2171 1892 2172 1896
rect 2166 1891 2172 1892
rect 2262 1896 2268 1897
rect 2262 1892 2263 1896
rect 2267 1892 2268 1896
rect 2262 1891 2268 1892
rect 2358 1896 2364 1897
rect 2358 1892 2359 1896
rect 2363 1892 2364 1896
rect 2358 1891 2364 1892
rect 2438 1896 2444 1897
rect 2438 1892 2439 1896
rect 2443 1892 2444 1896
rect 2502 1895 2503 1899
rect 2507 1895 2508 1899
rect 2502 1894 2508 1895
rect 2438 1891 2444 1892
rect 1286 1888 1292 1889
rect 1606 1880 1612 1881
rect 1326 1877 1332 1878
rect 110 1876 116 1877
rect 1286 1876 1292 1877
rect 110 1872 111 1876
rect 115 1872 116 1876
rect 110 1871 116 1872
rect 150 1875 156 1876
rect 150 1871 151 1875
rect 155 1871 156 1875
rect 150 1870 156 1871
rect 158 1875 164 1876
rect 158 1871 159 1875
rect 163 1874 164 1875
rect 171 1875 177 1876
rect 171 1874 172 1875
rect 163 1872 172 1874
rect 163 1871 164 1872
rect 158 1870 164 1871
rect 171 1871 172 1872
rect 176 1871 177 1875
rect 171 1870 177 1871
rect 206 1875 212 1876
rect 206 1871 207 1875
rect 211 1871 212 1875
rect 227 1875 233 1876
rect 227 1874 228 1875
rect 206 1870 212 1871
rect 216 1872 228 1874
rect 216 1862 218 1872
rect 227 1871 228 1872
rect 232 1871 233 1875
rect 227 1870 233 1871
rect 286 1875 292 1876
rect 286 1871 287 1875
rect 291 1871 292 1875
rect 307 1875 313 1876
rect 307 1874 308 1875
rect 286 1870 292 1871
rect 296 1872 308 1874
rect 296 1866 298 1872
rect 307 1871 308 1872
rect 312 1871 313 1875
rect 307 1870 313 1871
rect 374 1875 380 1876
rect 374 1871 375 1875
rect 379 1871 380 1875
rect 374 1870 380 1871
rect 395 1875 401 1876
rect 395 1871 396 1875
rect 400 1874 401 1875
rect 450 1875 456 1876
rect 450 1874 451 1875
rect 400 1872 451 1874
rect 400 1871 401 1872
rect 395 1870 401 1871
rect 450 1871 451 1872
rect 455 1871 456 1875
rect 450 1870 456 1871
rect 470 1875 476 1876
rect 470 1871 471 1875
rect 475 1871 476 1875
rect 470 1870 476 1871
rect 491 1875 497 1876
rect 491 1871 492 1875
rect 496 1871 497 1875
rect 491 1870 497 1871
rect 558 1875 564 1876
rect 558 1871 559 1875
rect 563 1871 564 1875
rect 558 1870 564 1871
rect 574 1875 585 1876
rect 574 1871 575 1875
rect 579 1871 580 1875
rect 584 1871 585 1875
rect 574 1870 585 1871
rect 646 1875 652 1876
rect 646 1871 647 1875
rect 651 1871 652 1875
rect 667 1875 673 1876
rect 667 1874 668 1875
rect 646 1870 652 1871
rect 656 1872 668 1874
rect 132 1860 218 1862
rect 220 1864 298 1866
rect 132 1858 134 1860
rect 220 1858 222 1864
rect 493 1862 495 1870
rect 656 1862 658 1872
rect 667 1871 668 1872
rect 672 1871 673 1875
rect 667 1870 673 1871
rect 734 1875 740 1876
rect 734 1871 735 1875
rect 739 1871 740 1875
rect 734 1870 740 1871
rect 755 1875 761 1876
rect 755 1871 756 1875
rect 760 1874 761 1875
rect 794 1875 800 1876
rect 794 1874 795 1875
rect 760 1872 795 1874
rect 760 1871 761 1872
rect 755 1870 761 1871
rect 794 1871 795 1872
rect 799 1871 800 1875
rect 794 1870 800 1871
rect 814 1875 820 1876
rect 814 1871 815 1875
rect 819 1871 820 1875
rect 814 1870 820 1871
rect 835 1875 841 1876
rect 835 1871 836 1875
rect 840 1874 841 1875
rect 866 1875 872 1876
rect 866 1874 867 1875
rect 840 1872 867 1874
rect 840 1871 841 1872
rect 835 1870 841 1871
rect 866 1871 867 1872
rect 871 1871 872 1875
rect 866 1870 872 1871
rect 886 1875 892 1876
rect 886 1871 887 1875
rect 891 1871 892 1875
rect 886 1870 892 1871
rect 907 1875 913 1876
rect 907 1871 908 1875
rect 912 1874 913 1875
rect 938 1875 944 1876
rect 938 1874 939 1875
rect 912 1872 939 1874
rect 912 1871 913 1872
rect 907 1870 913 1871
rect 938 1871 939 1872
rect 943 1871 944 1875
rect 938 1870 944 1871
rect 958 1875 964 1876
rect 958 1871 959 1875
rect 963 1871 964 1875
rect 958 1870 964 1871
rect 979 1875 985 1876
rect 979 1871 980 1875
rect 984 1874 985 1875
rect 1022 1875 1028 1876
rect 1022 1874 1023 1875
rect 984 1872 1023 1874
rect 984 1871 985 1872
rect 979 1870 985 1871
rect 1022 1871 1023 1872
rect 1027 1871 1028 1875
rect 1022 1870 1028 1871
rect 1030 1875 1036 1876
rect 1030 1871 1031 1875
rect 1035 1871 1036 1875
rect 1030 1870 1036 1871
rect 1051 1875 1060 1876
rect 1051 1871 1052 1875
rect 1059 1871 1060 1875
rect 1051 1870 1060 1871
rect 1102 1875 1108 1876
rect 1102 1871 1103 1875
rect 1107 1871 1108 1875
rect 1102 1870 1108 1871
rect 1123 1875 1129 1876
rect 1123 1871 1124 1875
rect 1128 1874 1129 1875
rect 1150 1875 1156 1876
rect 1150 1874 1151 1875
rect 1128 1872 1151 1874
rect 1128 1871 1129 1872
rect 1123 1870 1129 1871
rect 1150 1871 1151 1872
rect 1155 1871 1156 1875
rect 1150 1870 1156 1871
rect 1174 1875 1180 1876
rect 1174 1871 1175 1875
rect 1179 1871 1180 1875
rect 1195 1875 1201 1876
rect 1195 1874 1196 1875
rect 1174 1870 1180 1871
rect 1184 1872 1196 1874
rect 982 1867 988 1868
rect 750 1863 756 1864
rect 750 1862 751 1863
rect 268 1860 495 1862
rect 540 1860 658 1862
rect 660 1860 751 1862
rect 268 1858 270 1860
rect 540 1858 542 1860
rect 660 1858 662 1860
rect 750 1859 751 1860
rect 755 1859 756 1863
rect 982 1863 983 1867
rect 987 1866 988 1867
rect 1184 1866 1186 1872
rect 1195 1871 1196 1872
rect 1200 1871 1201 1875
rect 1286 1872 1287 1876
rect 1291 1872 1292 1876
rect 1326 1873 1327 1877
rect 1331 1873 1332 1877
rect 1606 1876 1607 1880
rect 1611 1876 1612 1880
rect 1606 1875 1612 1876
rect 1662 1880 1668 1881
rect 1662 1876 1663 1880
rect 1667 1876 1668 1880
rect 1662 1875 1668 1876
rect 1726 1880 1732 1881
rect 1726 1876 1727 1880
rect 1731 1876 1732 1880
rect 1726 1875 1732 1876
rect 1798 1880 1804 1881
rect 1798 1876 1799 1880
rect 1803 1876 1804 1880
rect 1798 1875 1804 1876
rect 1870 1880 1876 1881
rect 1870 1876 1871 1880
rect 1875 1876 1876 1880
rect 1870 1875 1876 1876
rect 1942 1880 1948 1881
rect 1942 1876 1943 1880
rect 1947 1876 1948 1880
rect 1942 1875 1948 1876
rect 2006 1880 2012 1881
rect 2006 1876 2007 1880
rect 2011 1876 2012 1880
rect 2006 1875 2012 1876
rect 2070 1880 2076 1881
rect 2070 1876 2071 1880
rect 2075 1876 2076 1880
rect 2070 1875 2076 1876
rect 2134 1880 2140 1881
rect 2134 1876 2135 1880
rect 2139 1876 2140 1880
rect 2134 1875 2140 1876
rect 2198 1880 2204 1881
rect 2198 1876 2199 1880
rect 2203 1876 2204 1880
rect 2198 1875 2204 1876
rect 2262 1880 2268 1881
rect 2262 1876 2263 1880
rect 2267 1876 2268 1880
rect 2262 1875 2268 1876
rect 2326 1880 2332 1881
rect 2326 1876 2327 1880
rect 2331 1876 2332 1880
rect 2326 1875 2332 1876
rect 2382 1880 2388 1881
rect 2382 1876 2383 1880
rect 2387 1876 2388 1880
rect 2382 1875 2388 1876
rect 2438 1880 2444 1881
rect 2438 1876 2439 1880
rect 2443 1876 2444 1880
rect 2438 1875 2444 1876
rect 2502 1877 2508 1878
rect 1326 1872 1332 1873
rect 2502 1873 2503 1877
rect 2507 1873 2508 1877
rect 2502 1872 2508 1873
rect 1286 1871 1292 1872
rect 1195 1870 1201 1871
rect 987 1864 1186 1866
rect 987 1863 988 1864
rect 982 1862 988 1863
rect 750 1858 756 1859
rect 1326 1860 1332 1861
rect 2502 1860 2508 1861
rect 131 1857 137 1858
rect 131 1853 132 1857
rect 136 1853 137 1857
rect 131 1852 137 1853
rect 187 1857 222 1858
rect 187 1853 188 1857
rect 192 1856 222 1857
rect 267 1857 273 1858
rect 192 1853 193 1856
rect 187 1852 193 1853
rect 267 1853 268 1857
rect 272 1853 273 1857
rect 539 1857 545 1858
rect 267 1852 273 1853
rect 350 1855 361 1856
rect 350 1851 351 1855
rect 355 1851 356 1855
rect 360 1851 361 1855
rect 350 1850 361 1851
rect 450 1855 457 1856
rect 450 1851 451 1855
rect 456 1851 457 1855
rect 539 1853 540 1857
rect 544 1853 545 1857
rect 539 1852 545 1853
rect 627 1857 662 1858
rect 627 1853 628 1857
rect 632 1856 662 1857
rect 1326 1856 1327 1860
rect 1331 1856 1332 1860
rect 632 1853 633 1856
rect 627 1852 633 1853
rect 710 1855 721 1856
rect 450 1850 457 1851
rect 710 1851 711 1855
rect 715 1851 716 1855
rect 720 1851 721 1855
rect 794 1855 801 1856
rect 710 1850 721 1851
rect 786 1851 792 1852
rect 786 1850 787 1851
rect 748 1848 787 1850
rect 748 1846 750 1848
rect 786 1847 787 1848
rect 791 1847 792 1851
rect 794 1851 795 1855
rect 800 1851 801 1855
rect 794 1850 801 1851
rect 866 1855 873 1856
rect 866 1851 867 1855
rect 872 1851 873 1855
rect 866 1850 873 1851
rect 938 1855 945 1856
rect 938 1851 939 1855
rect 944 1851 945 1855
rect 938 1850 945 1851
rect 950 1855 956 1856
rect 950 1851 951 1855
rect 955 1854 956 1855
rect 1011 1855 1017 1856
rect 1011 1854 1012 1855
rect 955 1852 1012 1854
rect 955 1851 956 1852
rect 950 1850 956 1851
rect 1011 1851 1012 1852
rect 1016 1851 1017 1855
rect 1011 1850 1017 1851
rect 1022 1855 1028 1856
rect 1022 1851 1023 1855
rect 1027 1854 1028 1855
rect 1083 1855 1089 1856
rect 1083 1854 1084 1855
rect 1027 1852 1084 1854
rect 1027 1851 1028 1852
rect 1022 1850 1028 1851
rect 1083 1851 1084 1852
rect 1088 1851 1089 1855
rect 1083 1850 1089 1851
rect 1150 1855 1161 1856
rect 1326 1855 1332 1856
rect 1622 1859 1628 1860
rect 1622 1855 1623 1859
rect 1627 1855 1628 1859
rect 1150 1851 1151 1855
rect 1155 1851 1156 1855
rect 1160 1851 1161 1855
rect 1622 1854 1628 1855
rect 1643 1859 1649 1860
rect 1643 1855 1644 1859
rect 1648 1858 1649 1859
rect 1658 1859 1664 1860
rect 1658 1858 1659 1859
rect 1648 1856 1659 1858
rect 1648 1855 1649 1856
rect 1643 1854 1649 1855
rect 1658 1855 1659 1856
rect 1663 1855 1664 1859
rect 1658 1854 1664 1855
rect 1678 1859 1684 1860
rect 1678 1855 1679 1859
rect 1683 1855 1684 1859
rect 1678 1854 1684 1855
rect 1699 1859 1705 1860
rect 1699 1855 1700 1859
rect 1704 1858 1705 1859
rect 1722 1859 1728 1860
rect 1722 1858 1723 1859
rect 1704 1856 1723 1858
rect 1704 1855 1705 1856
rect 1699 1854 1705 1855
rect 1722 1855 1723 1856
rect 1727 1855 1728 1859
rect 1722 1854 1728 1855
rect 1742 1859 1748 1860
rect 1742 1855 1743 1859
rect 1747 1855 1748 1859
rect 1742 1854 1748 1855
rect 1763 1859 1772 1860
rect 1763 1855 1764 1859
rect 1771 1855 1772 1859
rect 1763 1854 1772 1855
rect 1814 1859 1820 1860
rect 1814 1855 1815 1859
rect 1819 1855 1820 1859
rect 1835 1859 1841 1860
rect 1835 1858 1836 1859
rect 1814 1854 1820 1855
rect 1824 1856 1836 1858
rect 1150 1850 1161 1851
rect 1824 1850 1826 1856
rect 1835 1855 1836 1856
rect 1840 1855 1841 1859
rect 1835 1854 1841 1855
rect 1886 1859 1892 1860
rect 1886 1855 1887 1859
rect 1891 1855 1892 1859
rect 1886 1854 1892 1855
rect 1894 1859 1900 1860
rect 1894 1855 1895 1859
rect 1899 1858 1900 1859
rect 1907 1859 1913 1860
rect 1907 1858 1908 1859
rect 1899 1856 1908 1858
rect 1899 1855 1900 1856
rect 1894 1854 1900 1855
rect 1907 1855 1908 1856
rect 1912 1855 1913 1859
rect 1907 1854 1913 1855
rect 1958 1859 1964 1860
rect 1958 1855 1959 1859
rect 1963 1855 1964 1859
rect 1979 1859 1985 1860
rect 1979 1858 1980 1859
rect 1958 1854 1964 1855
rect 1968 1856 1980 1858
rect 1968 1850 1970 1856
rect 1979 1855 1980 1856
rect 1984 1855 1985 1859
rect 1979 1854 1985 1855
rect 2022 1859 2028 1860
rect 2022 1855 2023 1859
rect 2027 1855 2028 1859
rect 2022 1854 2028 1855
rect 2043 1859 2049 1860
rect 2043 1855 2044 1859
rect 2048 1858 2049 1859
rect 2066 1859 2072 1860
rect 2066 1858 2067 1859
rect 2048 1856 2067 1858
rect 2048 1855 2049 1856
rect 2043 1854 2049 1855
rect 2066 1855 2067 1856
rect 2071 1855 2072 1859
rect 2066 1854 2072 1855
rect 2086 1859 2092 1860
rect 2086 1855 2087 1859
rect 2091 1855 2092 1859
rect 2086 1854 2092 1855
rect 2107 1859 2113 1860
rect 2107 1855 2108 1859
rect 2112 1858 2113 1859
rect 2130 1859 2136 1860
rect 2130 1858 2131 1859
rect 2112 1856 2131 1858
rect 2112 1855 2113 1856
rect 2107 1854 2113 1855
rect 2130 1855 2131 1856
rect 2135 1855 2136 1859
rect 2130 1854 2136 1855
rect 2150 1859 2156 1860
rect 2150 1855 2151 1859
rect 2155 1855 2156 1859
rect 2150 1854 2156 1855
rect 2171 1859 2177 1860
rect 2171 1855 2172 1859
rect 2176 1858 2177 1859
rect 2194 1859 2200 1860
rect 2194 1858 2195 1859
rect 2176 1856 2195 1858
rect 2176 1855 2177 1856
rect 2171 1854 2177 1855
rect 2194 1855 2195 1856
rect 2199 1855 2200 1859
rect 2194 1854 2200 1855
rect 2214 1859 2220 1860
rect 2214 1855 2215 1859
rect 2219 1855 2220 1859
rect 2214 1854 2220 1855
rect 2235 1859 2241 1860
rect 2235 1855 2236 1859
rect 2240 1858 2241 1859
rect 2258 1859 2264 1860
rect 2258 1858 2259 1859
rect 2240 1856 2259 1858
rect 2240 1855 2241 1856
rect 2235 1854 2241 1855
rect 2258 1855 2259 1856
rect 2263 1855 2264 1859
rect 2258 1854 2264 1855
rect 2278 1859 2284 1860
rect 2278 1855 2279 1859
rect 2283 1855 2284 1859
rect 2278 1854 2284 1855
rect 2299 1859 2305 1860
rect 2299 1855 2300 1859
rect 2304 1858 2305 1859
rect 2322 1859 2328 1860
rect 2322 1858 2323 1859
rect 2304 1856 2323 1858
rect 2304 1855 2305 1856
rect 2299 1854 2305 1855
rect 2322 1855 2323 1856
rect 2327 1855 2328 1859
rect 2322 1854 2328 1855
rect 2342 1859 2348 1860
rect 2342 1855 2343 1859
rect 2347 1855 2348 1859
rect 2342 1854 2348 1855
rect 2363 1859 2369 1860
rect 2363 1855 2364 1859
rect 2368 1858 2369 1859
rect 2378 1859 2384 1860
rect 2378 1858 2379 1859
rect 2368 1856 2379 1858
rect 2368 1855 2369 1856
rect 2363 1854 2369 1855
rect 2378 1855 2379 1856
rect 2383 1855 2384 1859
rect 2378 1854 2384 1855
rect 2398 1859 2404 1860
rect 2398 1855 2399 1859
rect 2403 1855 2404 1859
rect 2398 1854 2404 1855
rect 2418 1859 2425 1860
rect 2418 1855 2419 1859
rect 2424 1855 2425 1859
rect 2418 1854 2425 1855
rect 2454 1859 2460 1860
rect 2454 1855 2455 1859
rect 2459 1855 2460 1859
rect 2454 1854 2460 1855
rect 2462 1859 2468 1860
rect 2462 1855 2463 1859
rect 2467 1858 2468 1859
rect 2475 1859 2481 1860
rect 2475 1858 2476 1859
rect 2467 1856 2476 1858
rect 2467 1855 2468 1856
rect 2462 1854 2468 1855
rect 2475 1855 2476 1856
rect 2480 1855 2481 1859
rect 2502 1856 2503 1860
rect 2507 1856 2508 1860
rect 2502 1855 2508 1856
rect 2475 1854 2481 1855
rect 786 1846 792 1847
rect 1604 1848 1826 1850
rect 1868 1848 1970 1850
rect 667 1845 750 1846
rect 131 1843 137 1844
rect 131 1839 132 1843
rect 136 1842 137 1843
rect 158 1843 164 1844
rect 158 1842 159 1843
rect 136 1840 159 1842
rect 136 1839 137 1840
rect 131 1838 137 1839
rect 158 1839 159 1840
rect 163 1839 164 1843
rect 158 1838 164 1839
rect 174 1843 180 1844
rect 174 1839 175 1843
rect 179 1842 180 1843
rect 187 1843 193 1844
rect 187 1842 188 1843
rect 179 1840 188 1842
rect 179 1839 180 1840
rect 174 1838 180 1839
rect 187 1839 188 1840
rect 192 1839 193 1843
rect 187 1838 193 1839
rect 230 1843 236 1844
rect 230 1839 231 1843
rect 235 1842 236 1843
rect 275 1843 281 1844
rect 275 1842 276 1843
rect 235 1840 276 1842
rect 235 1839 236 1840
rect 230 1838 236 1839
rect 275 1839 276 1840
rect 280 1839 281 1843
rect 275 1838 281 1839
rect 343 1843 349 1844
rect 343 1839 344 1843
rect 348 1842 349 1843
rect 371 1843 377 1844
rect 371 1842 372 1843
rect 348 1840 372 1842
rect 348 1839 349 1840
rect 343 1838 349 1839
rect 371 1839 372 1840
rect 376 1839 377 1843
rect 371 1838 377 1839
rect 410 1843 416 1844
rect 410 1839 411 1843
rect 415 1842 416 1843
rect 475 1843 481 1844
rect 475 1842 476 1843
rect 415 1840 476 1842
rect 415 1839 416 1840
rect 410 1838 416 1839
rect 475 1839 476 1840
rect 480 1839 481 1843
rect 475 1838 481 1839
rect 571 1843 580 1844
rect 571 1839 572 1843
rect 579 1839 580 1843
rect 667 1841 668 1845
rect 672 1844 750 1845
rect 672 1841 673 1844
rect 667 1840 673 1841
rect 755 1843 761 1844
rect 571 1838 580 1839
rect 755 1839 756 1843
rect 760 1839 761 1843
rect 755 1838 761 1839
rect 830 1843 841 1844
rect 830 1839 831 1843
rect 835 1839 836 1843
rect 840 1839 841 1843
rect 830 1838 841 1839
rect 907 1843 913 1844
rect 907 1839 908 1843
rect 912 1842 913 1843
rect 918 1843 924 1844
rect 918 1842 919 1843
rect 912 1840 919 1842
rect 912 1839 913 1840
rect 907 1838 913 1839
rect 918 1839 919 1840
rect 923 1839 924 1843
rect 918 1838 924 1839
rect 979 1843 988 1844
rect 979 1839 980 1843
rect 987 1839 988 1843
rect 979 1838 988 1839
rect 1022 1843 1028 1844
rect 1022 1839 1023 1843
rect 1027 1842 1028 1843
rect 1059 1843 1065 1844
rect 1059 1842 1060 1843
rect 1027 1840 1060 1842
rect 1027 1839 1028 1840
rect 1022 1838 1028 1839
rect 1059 1839 1060 1840
rect 1064 1839 1065 1843
rect 1059 1838 1065 1839
rect 1110 1843 1116 1844
rect 1110 1839 1111 1843
rect 1115 1842 1116 1843
rect 1139 1843 1145 1844
rect 1139 1842 1140 1843
rect 1115 1840 1140 1842
rect 1115 1839 1116 1840
rect 1110 1838 1116 1839
rect 1139 1839 1140 1840
rect 1144 1839 1145 1843
rect 1604 1842 1606 1848
rect 1868 1842 1870 1848
rect 2286 1847 2292 1848
rect 2286 1846 2287 1847
rect 2004 1844 2287 1846
rect 2004 1842 2006 1844
rect 2286 1843 2287 1844
rect 2291 1843 2292 1847
rect 2286 1842 2292 1843
rect 1139 1838 1145 1839
rect 1603 1841 1609 1842
rect 757 1830 759 1838
rect 1603 1837 1604 1841
rect 1608 1837 1609 1841
rect 1867 1841 1873 1842
rect 1603 1836 1609 1837
rect 1658 1839 1665 1840
rect 1658 1835 1659 1839
rect 1664 1835 1665 1839
rect 1658 1834 1665 1835
rect 1722 1839 1729 1840
rect 1722 1835 1723 1839
rect 1728 1835 1729 1839
rect 1722 1834 1729 1835
rect 1795 1839 1801 1840
rect 1795 1835 1796 1839
rect 1800 1838 1801 1839
rect 1800 1836 1854 1838
rect 1867 1837 1868 1841
rect 1872 1837 1873 1841
rect 2003 1841 2009 1842
rect 1867 1836 1873 1837
rect 1939 1839 1945 1840
rect 1800 1835 1801 1836
rect 1795 1834 1801 1835
rect 1852 1834 1854 1836
rect 1894 1835 1900 1836
rect 1894 1834 1895 1835
rect 1852 1832 1895 1834
rect 1894 1831 1895 1832
rect 1899 1831 1900 1835
rect 1939 1835 1940 1839
rect 1944 1838 1945 1839
rect 1970 1839 1976 1840
rect 1970 1838 1971 1839
rect 1944 1836 1971 1838
rect 1944 1835 1945 1836
rect 1939 1834 1945 1835
rect 1970 1835 1971 1836
rect 1975 1835 1976 1839
rect 2003 1837 2004 1841
rect 2008 1837 2009 1841
rect 2003 1836 2009 1837
rect 2066 1839 2073 1840
rect 1970 1834 1976 1835
rect 2066 1835 2067 1839
rect 2072 1835 2073 1839
rect 2066 1834 2073 1835
rect 2130 1839 2137 1840
rect 2130 1835 2131 1839
rect 2136 1835 2137 1839
rect 2130 1834 2137 1835
rect 2194 1839 2201 1840
rect 2194 1835 2195 1839
rect 2200 1835 2201 1839
rect 2194 1834 2201 1835
rect 2258 1839 2265 1840
rect 2258 1835 2259 1839
rect 2264 1835 2265 1839
rect 2258 1834 2265 1835
rect 2322 1839 2329 1840
rect 2322 1835 2323 1839
rect 2328 1835 2329 1839
rect 2322 1834 2329 1835
rect 2378 1839 2385 1840
rect 2378 1835 2379 1839
rect 2384 1835 2385 1839
rect 2378 1834 2385 1835
rect 2435 1839 2441 1840
rect 2435 1835 2436 1839
rect 2440 1838 2441 1839
rect 2470 1839 2476 1840
rect 2470 1838 2471 1839
rect 2440 1836 2471 1838
rect 2440 1835 2441 1836
rect 2435 1834 2441 1835
rect 2470 1835 2471 1836
rect 2475 1835 2476 1839
rect 2470 1834 2476 1835
rect 1894 1830 1900 1831
rect 757 1828 878 1830
rect 876 1826 878 1828
rect 150 1825 156 1826
rect 110 1824 116 1825
rect 110 1820 111 1824
rect 115 1820 116 1824
rect 150 1821 151 1825
rect 155 1821 156 1825
rect 206 1825 212 1826
rect 150 1820 156 1821
rect 171 1823 180 1824
rect 110 1819 116 1820
rect 171 1819 172 1823
rect 179 1819 180 1823
rect 206 1821 207 1825
rect 211 1821 212 1825
rect 294 1825 300 1826
rect 206 1820 212 1821
rect 227 1823 236 1824
rect 171 1818 180 1819
rect 227 1819 228 1823
rect 235 1819 236 1823
rect 294 1821 295 1825
rect 299 1821 300 1825
rect 390 1825 396 1826
rect 294 1820 300 1821
rect 315 1823 321 1824
rect 227 1818 236 1819
rect 315 1819 316 1823
rect 320 1822 321 1823
rect 343 1823 349 1824
rect 343 1822 344 1823
rect 320 1820 344 1822
rect 320 1819 321 1820
rect 315 1818 321 1819
rect 343 1819 344 1820
rect 348 1819 349 1823
rect 390 1821 391 1825
rect 395 1821 396 1825
rect 494 1825 500 1826
rect 390 1820 396 1821
rect 410 1823 417 1824
rect 343 1818 349 1819
rect 410 1819 411 1823
rect 416 1819 417 1823
rect 494 1821 495 1825
rect 499 1821 500 1825
rect 590 1825 596 1826
rect 494 1820 500 1821
rect 510 1823 521 1824
rect 410 1818 417 1819
rect 510 1819 511 1823
rect 515 1819 516 1823
rect 520 1819 521 1823
rect 590 1821 591 1825
rect 595 1821 596 1825
rect 686 1825 692 1826
rect 590 1820 596 1821
rect 611 1823 620 1824
rect 510 1818 521 1819
rect 611 1819 612 1823
rect 619 1819 620 1823
rect 686 1821 687 1825
rect 691 1821 692 1825
rect 774 1825 780 1826
rect 686 1820 692 1821
rect 707 1823 716 1824
rect 611 1818 620 1819
rect 707 1819 708 1823
rect 715 1819 716 1823
rect 774 1821 775 1825
rect 779 1821 780 1825
rect 854 1825 860 1826
rect 774 1820 780 1821
rect 786 1823 792 1824
rect 707 1818 716 1819
rect 786 1819 787 1823
rect 791 1822 792 1823
rect 795 1823 801 1824
rect 795 1822 796 1823
rect 791 1820 796 1822
rect 791 1819 792 1820
rect 786 1818 792 1819
rect 795 1819 796 1820
rect 800 1819 801 1823
rect 854 1821 855 1825
rect 859 1821 860 1825
rect 854 1820 860 1821
rect 875 1825 881 1826
rect 875 1821 876 1825
rect 880 1821 881 1825
rect 875 1820 881 1821
rect 926 1825 932 1826
rect 926 1821 927 1825
rect 931 1821 932 1825
rect 998 1825 1004 1826
rect 926 1820 932 1821
rect 947 1823 956 1824
rect 795 1818 801 1819
rect 947 1819 948 1823
rect 955 1819 956 1823
rect 998 1821 999 1825
rect 1003 1821 1004 1825
rect 1078 1825 1084 1826
rect 998 1820 1004 1821
rect 1019 1823 1028 1824
rect 947 1818 956 1819
rect 1019 1819 1020 1823
rect 1027 1819 1028 1823
rect 1078 1821 1079 1825
rect 1083 1821 1084 1825
rect 1158 1825 1164 1826
rect 1078 1820 1084 1821
rect 1099 1823 1105 1824
rect 1019 1818 1028 1819
rect 1099 1819 1100 1823
rect 1104 1822 1105 1823
rect 1110 1823 1116 1824
rect 1110 1822 1111 1823
rect 1104 1820 1111 1822
rect 1104 1819 1105 1820
rect 1099 1818 1105 1819
rect 1110 1819 1111 1820
rect 1115 1819 1116 1823
rect 1158 1821 1159 1825
rect 1163 1821 1164 1825
rect 1286 1824 1292 1825
rect 1158 1820 1164 1821
rect 1174 1823 1185 1824
rect 1110 1818 1116 1819
rect 1174 1819 1175 1823
rect 1179 1819 1180 1823
rect 1184 1819 1185 1823
rect 1286 1820 1287 1824
rect 1291 1820 1292 1824
rect 1286 1819 1292 1820
rect 1611 1823 1617 1824
rect 1611 1819 1612 1823
rect 1616 1822 1617 1823
rect 1654 1823 1660 1824
rect 1654 1822 1655 1823
rect 1616 1820 1655 1822
rect 1616 1819 1617 1820
rect 1174 1818 1185 1819
rect 1611 1818 1617 1819
rect 1654 1819 1655 1820
rect 1659 1819 1660 1823
rect 1654 1818 1660 1819
rect 1662 1823 1668 1824
rect 1662 1819 1663 1823
rect 1667 1822 1668 1823
rect 1699 1823 1705 1824
rect 1699 1822 1700 1823
rect 1667 1820 1700 1822
rect 1667 1819 1668 1820
rect 1662 1818 1668 1819
rect 1699 1819 1700 1820
rect 1704 1819 1705 1823
rect 1699 1818 1705 1819
rect 1750 1823 1756 1824
rect 1750 1819 1751 1823
rect 1755 1822 1756 1823
rect 1795 1823 1801 1824
rect 1795 1822 1796 1823
rect 1755 1820 1796 1822
rect 1755 1819 1756 1820
rect 1750 1818 1756 1819
rect 1795 1819 1796 1820
rect 1800 1819 1801 1823
rect 1795 1818 1801 1819
rect 1855 1823 1861 1824
rect 1855 1819 1856 1823
rect 1860 1822 1861 1823
rect 1907 1823 1913 1824
rect 1907 1822 1908 1823
rect 1860 1820 1908 1822
rect 1860 1819 1861 1820
rect 1855 1818 1861 1819
rect 1907 1819 1908 1820
rect 1912 1819 1913 1823
rect 1907 1818 1913 1819
rect 1959 1823 1965 1824
rect 1959 1819 1960 1823
rect 1964 1822 1965 1823
rect 2035 1823 2041 1824
rect 2035 1822 2036 1823
rect 1964 1820 2036 1822
rect 1964 1819 1965 1820
rect 1959 1818 1965 1819
rect 2035 1819 2036 1820
rect 2040 1819 2041 1823
rect 2035 1818 2041 1819
rect 2171 1823 2177 1824
rect 2171 1819 2172 1823
rect 2176 1822 2177 1823
rect 2315 1823 2321 1824
rect 2176 1820 2310 1822
rect 2176 1819 2177 1820
rect 2171 1818 2177 1819
rect 1970 1811 1976 1812
rect 110 1807 116 1808
rect 110 1803 111 1807
rect 115 1803 116 1807
rect 1286 1807 1292 1808
rect 110 1802 116 1803
rect 134 1804 140 1805
rect 134 1800 135 1804
rect 139 1800 140 1804
rect 134 1799 140 1800
rect 190 1804 196 1805
rect 190 1800 191 1804
rect 195 1800 196 1804
rect 190 1799 196 1800
rect 278 1804 284 1805
rect 278 1800 279 1804
rect 283 1800 284 1804
rect 278 1799 284 1800
rect 374 1804 380 1805
rect 374 1800 375 1804
rect 379 1800 380 1804
rect 374 1799 380 1800
rect 478 1804 484 1805
rect 478 1800 479 1804
rect 483 1800 484 1804
rect 478 1799 484 1800
rect 574 1804 580 1805
rect 574 1800 575 1804
rect 579 1800 580 1804
rect 574 1799 580 1800
rect 670 1804 676 1805
rect 670 1800 671 1804
rect 675 1800 676 1804
rect 670 1799 676 1800
rect 758 1804 764 1805
rect 758 1800 759 1804
rect 763 1800 764 1804
rect 758 1799 764 1800
rect 838 1804 844 1805
rect 838 1800 839 1804
rect 843 1800 844 1804
rect 838 1799 844 1800
rect 910 1804 916 1805
rect 910 1800 911 1804
rect 915 1800 916 1804
rect 910 1799 916 1800
rect 982 1804 988 1805
rect 982 1800 983 1804
rect 987 1800 988 1804
rect 982 1799 988 1800
rect 1062 1804 1068 1805
rect 1062 1800 1063 1804
rect 1067 1800 1068 1804
rect 1062 1799 1068 1800
rect 1142 1804 1148 1805
rect 1142 1800 1143 1804
rect 1147 1800 1148 1804
rect 1286 1803 1287 1807
rect 1291 1803 1292 1807
rect 1970 1807 1971 1811
rect 1975 1810 1976 1811
rect 2308 1810 2310 1820
rect 2315 1819 2316 1823
rect 2320 1822 2321 1823
rect 2326 1823 2332 1824
rect 2326 1822 2327 1823
rect 2320 1820 2327 1822
rect 2320 1819 2321 1820
rect 2315 1818 2321 1819
rect 2326 1819 2327 1820
rect 2331 1819 2332 1823
rect 2326 1818 2332 1819
rect 2435 1823 2441 1824
rect 2435 1819 2436 1823
rect 2440 1822 2441 1823
rect 2462 1823 2468 1824
rect 2462 1822 2463 1823
rect 2440 1820 2463 1822
rect 2440 1819 2441 1820
rect 2435 1818 2441 1819
rect 2462 1819 2463 1820
rect 2467 1819 2468 1823
rect 2462 1818 2468 1819
rect 1975 1808 2078 1810
rect 2308 1808 2358 1810
rect 1975 1807 1976 1808
rect 1970 1806 1976 1807
rect 2076 1806 2078 1808
rect 2356 1806 2358 1808
rect 1630 1805 1636 1806
rect 1286 1802 1292 1803
rect 1326 1804 1332 1805
rect 1142 1799 1148 1800
rect 1326 1800 1327 1804
rect 1331 1800 1332 1804
rect 1630 1801 1631 1805
rect 1635 1801 1636 1805
rect 1718 1805 1724 1806
rect 1630 1800 1636 1801
rect 1651 1803 1657 1804
rect 1326 1799 1332 1800
rect 1651 1799 1652 1803
rect 1656 1802 1657 1803
rect 1662 1803 1668 1804
rect 1662 1802 1663 1803
rect 1656 1800 1663 1802
rect 1656 1799 1657 1800
rect 1651 1798 1657 1799
rect 1662 1799 1663 1800
rect 1667 1799 1668 1803
rect 1718 1801 1719 1805
rect 1723 1801 1724 1805
rect 1814 1805 1820 1806
rect 1718 1800 1724 1801
rect 1739 1803 1745 1804
rect 1662 1798 1668 1799
rect 1739 1799 1740 1803
rect 1744 1802 1745 1803
rect 1750 1803 1756 1804
rect 1750 1802 1751 1803
rect 1744 1800 1751 1802
rect 1744 1799 1745 1800
rect 1739 1798 1745 1799
rect 1750 1799 1751 1800
rect 1755 1799 1756 1803
rect 1814 1801 1815 1805
rect 1819 1801 1820 1805
rect 1926 1805 1932 1806
rect 1814 1800 1820 1801
rect 1835 1803 1841 1804
rect 1750 1798 1756 1799
rect 1835 1799 1836 1803
rect 1840 1802 1841 1803
rect 1855 1803 1861 1804
rect 1855 1802 1856 1803
rect 1840 1800 1856 1802
rect 1840 1799 1841 1800
rect 1835 1798 1841 1799
rect 1855 1799 1856 1800
rect 1860 1799 1861 1803
rect 1926 1801 1927 1805
rect 1931 1801 1932 1805
rect 2054 1805 2060 1806
rect 1926 1800 1932 1801
rect 1947 1803 1953 1804
rect 1855 1798 1861 1799
rect 1947 1799 1948 1803
rect 1952 1802 1953 1803
rect 1959 1803 1965 1804
rect 1959 1802 1960 1803
rect 1952 1800 1960 1802
rect 1952 1799 1953 1800
rect 1947 1798 1953 1799
rect 1959 1799 1960 1800
rect 1964 1799 1965 1803
rect 2054 1801 2055 1805
rect 2059 1801 2060 1805
rect 2054 1800 2060 1801
rect 2075 1805 2081 1806
rect 2075 1801 2076 1805
rect 2080 1801 2081 1805
rect 2075 1800 2081 1801
rect 2190 1805 2196 1806
rect 2190 1801 2191 1805
rect 2195 1801 2196 1805
rect 2334 1805 2340 1806
rect 2190 1800 2196 1801
rect 2206 1803 2217 1804
rect 1959 1798 1965 1799
rect 2206 1799 2207 1803
rect 2211 1799 2212 1803
rect 2216 1799 2217 1803
rect 2334 1801 2335 1805
rect 2339 1801 2340 1805
rect 2334 1800 2340 1801
rect 2355 1805 2361 1806
rect 2355 1801 2356 1805
rect 2360 1801 2361 1805
rect 2355 1800 2361 1801
rect 2454 1805 2460 1806
rect 2454 1801 2455 1805
rect 2459 1801 2460 1805
rect 2502 1804 2508 1805
rect 2454 1800 2460 1801
rect 2470 1803 2481 1804
rect 2206 1798 2217 1799
rect 2470 1799 2471 1803
rect 2475 1799 2476 1803
rect 2480 1799 2481 1803
rect 2502 1800 2503 1804
rect 2507 1800 2508 1804
rect 2502 1799 2508 1800
rect 2470 1798 2481 1799
rect 1326 1787 1332 1788
rect 1326 1783 1327 1787
rect 1331 1783 1332 1787
rect 2502 1787 2508 1788
rect 1326 1782 1332 1783
rect 1614 1784 1620 1785
rect 134 1780 140 1781
rect 110 1777 116 1778
rect 110 1773 111 1777
rect 115 1773 116 1777
rect 134 1776 135 1780
rect 139 1776 140 1780
rect 134 1775 140 1776
rect 198 1780 204 1781
rect 198 1776 199 1780
rect 203 1776 204 1780
rect 198 1775 204 1776
rect 294 1780 300 1781
rect 294 1776 295 1780
rect 299 1776 300 1780
rect 294 1775 300 1776
rect 398 1780 404 1781
rect 398 1776 399 1780
rect 403 1776 404 1780
rect 398 1775 404 1776
rect 502 1780 508 1781
rect 502 1776 503 1780
rect 507 1776 508 1780
rect 502 1775 508 1776
rect 606 1780 612 1781
rect 606 1776 607 1780
rect 611 1776 612 1780
rect 606 1775 612 1776
rect 702 1780 708 1781
rect 702 1776 703 1780
rect 707 1776 708 1780
rect 702 1775 708 1776
rect 798 1780 804 1781
rect 798 1776 799 1780
rect 803 1776 804 1780
rect 798 1775 804 1776
rect 886 1780 892 1781
rect 886 1776 887 1780
rect 891 1776 892 1780
rect 886 1775 892 1776
rect 974 1780 980 1781
rect 974 1776 975 1780
rect 979 1776 980 1780
rect 974 1775 980 1776
rect 1062 1780 1068 1781
rect 1062 1776 1063 1780
rect 1067 1776 1068 1780
rect 1062 1775 1068 1776
rect 1150 1780 1156 1781
rect 1150 1776 1151 1780
rect 1155 1776 1156 1780
rect 1614 1780 1615 1784
rect 1619 1780 1620 1784
rect 1614 1779 1620 1780
rect 1702 1784 1708 1785
rect 1702 1780 1703 1784
rect 1707 1780 1708 1784
rect 1702 1779 1708 1780
rect 1798 1784 1804 1785
rect 1798 1780 1799 1784
rect 1803 1780 1804 1784
rect 1798 1779 1804 1780
rect 1910 1784 1916 1785
rect 1910 1780 1911 1784
rect 1915 1780 1916 1784
rect 1910 1779 1916 1780
rect 2038 1784 2044 1785
rect 2038 1780 2039 1784
rect 2043 1780 2044 1784
rect 2038 1779 2044 1780
rect 2174 1784 2180 1785
rect 2174 1780 2175 1784
rect 2179 1780 2180 1784
rect 2174 1779 2180 1780
rect 2318 1784 2324 1785
rect 2318 1780 2319 1784
rect 2323 1780 2324 1784
rect 2318 1779 2324 1780
rect 2438 1784 2444 1785
rect 2438 1780 2439 1784
rect 2443 1780 2444 1784
rect 2502 1783 2503 1787
rect 2507 1783 2508 1787
rect 2502 1782 2508 1783
rect 2438 1779 2444 1780
rect 1150 1775 1156 1776
rect 1286 1777 1292 1778
rect 110 1772 116 1773
rect 1286 1773 1287 1777
rect 1291 1773 1292 1777
rect 1286 1772 1292 1773
rect 1526 1772 1532 1773
rect 1326 1769 1332 1770
rect 1326 1765 1327 1769
rect 1331 1765 1332 1769
rect 1526 1768 1527 1772
rect 1531 1768 1532 1772
rect 1526 1767 1532 1768
rect 1606 1772 1612 1773
rect 1606 1768 1607 1772
rect 1611 1768 1612 1772
rect 1606 1767 1612 1768
rect 1694 1772 1700 1773
rect 1694 1768 1695 1772
rect 1699 1768 1700 1772
rect 1694 1767 1700 1768
rect 1790 1772 1796 1773
rect 1790 1768 1791 1772
rect 1795 1768 1796 1772
rect 1790 1767 1796 1768
rect 1878 1772 1884 1773
rect 1878 1768 1879 1772
rect 1883 1768 1884 1772
rect 1878 1767 1884 1768
rect 1966 1772 1972 1773
rect 1966 1768 1967 1772
rect 1971 1768 1972 1772
rect 1966 1767 1972 1768
rect 2054 1772 2060 1773
rect 2054 1768 2055 1772
rect 2059 1768 2060 1772
rect 2054 1767 2060 1768
rect 2134 1772 2140 1773
rect 2134 1768 2135 1772
rect 2139 1768 2140 1772
rect 2134 1767 2140 1768
rect 2214 1772 2220 1773
rect 2214 1768 2215 1772
rect 2219 1768 2220 1772
rect 2214 1767 2220 1768
rect 2294 1772 2300 1773
rect 2294 1768 2295 1772
rect 2299 1768 2300 1772
rect 2294 1767 2300 1768
rect 2374 1772 2380 1773
rect 2374 1768 2375 1772
rect 2379 1768 2380 1772
rect 2374 1767 2380 1768
rect 2438 1772 2444 1773
rect 2438 1768 2439 1772
rect 2443 1768 2444 1772
rect 2438 1767 2444 1768
rect 2502 1769 2508 1770
rect 1326 1764 1332 1765
rect 2502 1765 2503 1769
rect 2507 1765 2508 1769
rect 2502 1764 2508 1765
rect 110 1760 116 1761
rect 1286 1760 1292 1761
rect 110 1756 111 1760
rect 115 1756 116 1760
rect 110 1755 116 1756
rect 150 1759 156 1760
rect 150 1755 151 1759
rect 155 1755 156 1759
rect 150 1754 156 1755
rect 171 1759 177 1760
rect 171 1755 172 1759
rect 176 1758 177 1759
rect 194 1759 200 1760
rect 194 1758 195 1759
rect 176 1756 195 1758
rect 176 1755 177 1756
rect 171 1754 177 1755
rect 194 1755 195 1756
rect 199 1755 200 1759
rect 194 1754 200 1755
rect 214 1759 220 1760
rect 214 1755 215 1759
rect 219 1755 220 1759
rect 214 1754 220 1755
rect 235 1759 241 1760
rect 235 1755 236 1759
rect 240 1758 241 1759
rect 290 1759 296 1760
rect 290 1758 291 1759
rect 240 1756 291 1758
rect 240 1755 241 1756
rect 235 1754 241 1755
rect 290 1755 291 1756
rect 295 1755 296 1759
rect 290 1754 296 1755
rect 310 1759 316 1760
rect 310 1755 311 1759
rect 315 1755 316 1759
rect 310 1754 316 1755
rect 331 1759 337 1760
rect 331 1755 332 1759
rect 336 1758 337 1759
rect 394 1759 400 1760
rect 394 1758 395 1759
rect 336 1756 395 1758
rect 336 1755 337 1756
rect 331 1754 337 1755
rect 394 1755 395 1756
rect 399 1755 400 1759
rect 394 1754 400 1755
rect 414 1759 420 1760
rect 414 1755 415 1759
rect 419 1755 420 1759
rect 414 1754 420 1755
rect 422 1759 428 1760
rect 422 1755 423 1759
rect 427 1758 428 1759
rect 435 1759 441 1760
rect 435 1758 436 1759
rect 427 1756 436 1758
rect 427 1755 428 1756
rect 422 1754 428 1755
rect 435 1755 436 1756
rect 440 1755 441 1759
rect 435 1754 441 1755
rect 518 1759 524 1760
rect 518 1755 519 1759
rect 523 1755 524 1759
rect 518 1754 524 1755
rect 539 1759 545 1760
rect 539 1755 540 1759
rect 544 1758 545 1759
rect 586 1759 592 1760
rect 586 1758 587 1759
rect 544 1756 587 1758
rect 544 1755 545 1756
rect 539 1754 545 1755
rect 586 1755 587 1756
rect 591 1755 592 1759
rect 586 1754 592 1755
rect 622 1759 628 1760
rect 622 1755 623 1759
rect 627 1755 628 1759
rect 643 1759 649 1760
rect 643 1758 644 1759
rect 622 1754 628 1755
rect 632 1756 644 1758
rect 632 1746 634 1756
rect 643 1755 644 1756
rect 648 1755 649 1759
rect 643 1754 649 1755
rect 718 1759 724 1760
rect 718 1755 719 1759
rect 723 1755 724 1759
rect 718 1754 724 1755
rect 739 1759 745 1760
rect 739 1755 740 1759
rect 744 1758 745 1759
rect 794 1759 800 1760
rect 794 1758 795 1759
rect 744 1756 795 1758
rect 744 1755 745 1756
rect 739 1754 745 1755
rect 794 1755 795 1756
rect 799 1755 800 1759
rect 794 1754 800 1755
rect 814 1759 820 1760
rect 814 1755 815 1759
rect 819 1755 820 1759
rect 814 1754 820 1755
rect 830 1759 841 1760
rect 830 1755 831 1759
rect 835 1755 836 1759
rect 840 1755 841 1759
rect 830 1754 841 1755
rect 902 1759 908 1760
rect 902 1755 903 1759
rect 907 1755 908 1759
rect 902 1754 908 1755
rect 918 1759 929 1760
rect 918 1755 919 1759
rect 923 1755 924 1759
rect 928 1755 929 1759
rect 918 1754 929 1755
rect 990 1759 996 1760
rect 990 1755 991 1759
rect 995 1755 996 1759
rect 990 1754 996 1755
rect 1011 1759 1017 1760
rect 1011 1755 1012 1759
rect 1016 1758 1017 1759
rect 1026 1759 1032 1760
rect 1026 1758 1027 1759
rect 1016 1756 1027 1758
rect 1016 1755 1017 1756
rect 1011 1754 1017 1755
rect 1026 1755 1027 1756
rect 1031 1755 1032 1759
rect 1026 1754 1032 1755
rect 1078 1759 1084 1760
rect 1078 1755 1079 1759
rect 1083 1755 1084 1759
rect 1099 1759 1105 1760
rect 1099 1758 1100 1759
rect 1078 1754 1084 1755
rect 1088 1756 1100 1758
rect 1088 1750 1090 1756
rect 1099 1755 1100 1756
rect 1104 1755 1105 1759
rect 1099 1754 1105 1755
rect 1166 1759 1172 1760
rect 1166 1755 1167 1759
rect 1171 1755 1172 1759
rect 1187 1759 1193 1760
rect 1187 1758 1188 1759
rect 1166 1754 1172 1755
rect 1176 1756 1188 1758
rect 500 1744 634 1746
rect 972 1748 1090 1750
rect 500 1742 502 1744
rect 972 1742 974 1748
rect 1176 1746 1178 1756
rect 1187 1755 1188 1756
rect 1192 1755 1193 1759
rect 1286 1756 1287 1760
rect 1291 1756 1292 1760
rect 1286 1755 1292 1756
rect 1187 1754 1193 1755
rect 1326 1752 1332 1753
rect 2502 1752 2508 1753
rect 1326 1748 1327 1752
rect 1331 1748 1332 1752
rect 1326 1747 1332 1748
rect 1542 1751 1548 1752
rect 1542 1747 1543 1751
rect 1547 1747 1548 1751
rect 1542 1746 1548 1747
rect 1563 1751 1569 1752
rect 1563 1747 1564 1751
rect 1568 1750 1569 1751
rect 1602 1751 1608 1752
rect 1602 1750 1603 1751
rect 1568 1748 1603 1750
rect 1568 1747 1569 1748
rect 1563 1746 1569 1747
rect 1602 1747 1603 1748
rect 1607 1747 1608 1751
rect 1602 1746 1608 1747
rect 1622 1751 1628 1752
rect 1622 1747 1623 1751
rect 1627 1747 1628 1751
rect 1622 1746 1628 1747
rect 1643 1751 1649 1752
rect 1643 1747 1644 1751
rect 1648 1750 1649 1751
rect 1690 1751 1696 1752
rect 1690 1750 1691 1751
rect 1648 1748 1691 1750
rect 1648 1747 1649 1748
rect 1643 1746 1649 1747
rect 1690 1747 1691 1748
rect 1695 1747 1696 1751
rect 1690 1746 1696 1747
rect 1710 1751 1716 1752
rect 1710 1747 1711 1751
rect 1715 1747 1716 1751
rect 1710 1746 1716 1747
rect 1731 1751 1737 1752
rect 1731 1747 1732 1751
rect 1736 1750 1737 1751
rect 1786 1751 1792 1752
rect 1786 1750 1787 1751
rect 1736 1748 1787 1750
rect 1736 1747 1737 1748
rect 1731 1746 1737 1747
rect 1786 1747 1787 1748
rect 1791 1747 1792 1751
rect 1786 1746 1792 1747
rect 1806 1751 1812 1752
rect 1806 1747 1807 1751
rect 1811 1747 1812 1751
rect 1806 1746 1812 1747
rect 1827 1751 1833 1752
rect 1827 1747 1828 1751
rect 1832 1750 1833 1751
rect 1874 1751 1880 1752
rect 1874 1750 1875 1751
rect 1832 1748 1875 1750
rect 1832 1747 1833 1748
rect 1827 1746 1833 1747
rect 1874 1747 1875 1748
rect 1879 1747 1880 1751
rect 1874 1746 1880 1747
rect 1894 1751 1900 1752
rect 1894 1747 1895 1751
rect 1899 1747 1900 1751
rect 1894 1746 1900 1747
rect 1914 1751 1921 1752
rect 1914 1747 1915 1751
rect 1920 1747 1921 1751
rect 1914 1746 1921 1747
rect 1982 1751 1988 1752
rect 1982 1747 1983 1751
rect 1987 1747 1988 1751
rect 1982 1746 1988 1747
rect 2003 1751 2009 1752
rect 2003 1747 2004 1751
rect 2008 1750 2009 1751
rect 2050 1751 2056 1752
rect 2050 1750 2051 1751
rect 2008 1748 2051 1750
rect 2008 1747 2009 1748
rect 2003 1746 2009 1747
rect 2050 1747 2051 1748
rect 2055 1747 2056 1751
rect 2050 1746 2056 1747
rect 2070 1751 2076 1752
rect 2070 1747 2071 1751
rect 2075 1747 2076 1751
rect 2070 1746 2076 1747
rect 2090 1751 2097 1752
rect 2090 1747 2091 1751
rect 2096 1747 2097 1751
rect 2090 1746 2097 1747
rect 2150 1751 2156 1752
rect 2150 1747 2151 1751
rect 2155 1747 2156 1751
rect 2171 1751 2177 1752
rect 2171 1750 2172 1751
rect 2150 1746 2156 1747
rect 2160 1748 2172 1750
rect 1061 1744 1178 1746
rect 1061 1742 1063 1744
rect 2160 1742 2162 1748
rect 2171 1747 2172 1748
rect 2176 1747 2177 1751
rect 2171 1746 2177 1747
rect 2230 1751 2236 1752
rect 2230 1747 2231 1751
rect 2235 1747 2236 1751
rect 2251 1751 2257 1752
rect 2251 1750 2252 1751
rect 2230 1746 2236 1747
rect 2240 1748 2252 1750
rect 499 1741 505 1742
rect 131 1739 140 1740
rect 131 1735 132 1739
rect 139 1735 140 1739
rect 131 1734 140 1735
rect 194 1739 201 1740
rect 194 1735 195 1739
rect 200 1735 201 1739
rect 194 1734 201 1735
rect 290 1739 297 1740
rect 290 1735 291 1739
rect 296 1735 297 1739
rect 290 1734 297 1735
rect 394 1739 401 1740
rect 394 1735 395 1739
rect 400 1735 401 1739
rect 499 1737 500 1741
rect 504 1737 505 1741
rect 971 1741 977 1742
rect 499 1736 505 1737
rect 603 1739 609 1740
rect 394 1734 401 1735
rect 603 1735 604 1739
rect 608 1738 609 1739
rect 614 1739 620 1740
rect 614 1738 615 1739
rect 608 1736 615 1738
rect 608 1735 609 1736
rect 603 1734 609 1735
rect 614 1735 615 1736
rect 619 1735 620 1739
rect 614 1734 620 1735
rect 699 1739 705 1740
rect 699 1735 700 1739
rect 704 1738 705 1739
rect 730 1739 736 1740
rect 730 1738 731 1739
rect 704 1736 731 1738
rect 704 1735 705 1736
rect 699 1734 705 1735
rect 730 1735 731 1736
rect 735 1735 736 1739
rect 730 1734 736 1735
rect 794 1739 801 1740
rect 794 1735 795 1739
rect 800 1735 801 1739
rect 794 1734 801 1735
rect 883 1739 889 1740
rect 883 1735 884 1739
rect 888 1738 889 1739
rect 954 1739 960 1740
rect 954 1738 955 1739
rect 888 1736 955 1738
rect 888 1735 889 1736
rect 883 1734 889 1735
rect 954 1735 955 1736
rect 959 1735 960 1739
rect 971 1737 972 1741
rect 976 1737 977 1741
rect 971 1736 977 1737
rect 1059 1741 1065 1742
rect 1059 1737 1060 1741
rect 1064 1737 1065 1741
rect 1999 1740 2162 1742
rect 1059 1736 1065 1737
rect 1147 1739 1153 1740
rect 954 1734 960 1735
rect 1147 1735 1148 1739
rect 1152 1738 1153 1739
rect 1174 1739 1180 1740
rect 1174 1738 1175 1739
rect 1152 1736 1175 1738
rect 1152 1735 1153 1736
rect 1147 1734 1153 1735
rect 1174 1735 1175 1736
rect 1179 1735 1180 1739
rect 1174 1734 1180 1735
rect 1999 1734 2001 1740
rect 2240 1738 2242 1748
rect 2251 1747 2252 1748
rect 2256 1747 2257 1751
rect 2251 1746 2257 1747
rect 2310 1751 2316 1752
rect 2310 1747 2311 1751
rect 2315 1747 2316 1751
rect 2310 1746 2316 1747
rect 2326 1751 2337 1752
rect 2326 1747 2327 1751
rect 2331 1747 2332 1751
rect 2336 1747 2337 1751
rect 2326 1746 2337 1747
rect 2390 1751 2396 1752
rect 2390 1747 2391 1751
rect 2395 1747 2396 1751
rect 2411 1751 2417 1752
rect 2411 1750 2412 1751
rect 2390 1746 2396 1747
rect 2400 1748 2412 1750
rect 2400 1738 2402 1748
rect 2411 1747 2412 1748
rect 2416 1747 2417 1751
rect 2411 1746 2417 1747
rect 2454 1751 2460 1752
rect 2454 1747 2455 1751
rect 2459 1747 2460 1751
rect 2454 1746 2460 1747
rect 2462 1751 2468 1752
rect 2462 1747 2463 1751
rect 2467 1750 2468 1751
rect 2475 1751 2481 1752
rect 2475 1750 2476 1751
rect 2467 1748 2476 1750
rect 2467 1747 2468 1748
rect 2462 1746 2468 1747
rect 2475 1747 2476 1748
rect 2480 1747 2481 1751
rect 2502 1748 2503 1752
rect 2507 1748 2508 1752
rect 2502 1747 2508 1748
rect 2475 1746 2481 1747
rect 2132 1736 2242 1738
rect 2292 1736 2402 1738
rect 2132 1734 2134 1736
rect 2292 1734 2294 1736
rect 1963 1733 2001 1734
rect 422 1731 428 1732
rect 422 1730 423 1731
rect 148 1728 423 1730
rect 148 1726 150 1728
rect 422 1727 423 1728
rect 427 1727 428 1731
rect 422 1726 428 1727
rect 1523 1731 1529 1732
rect 1523 1727 1524 1731
rect 1528 1730 1529 1731
rect 1594 1731 1600 1732
rect 1594 1730 1595 1731
rect 1528 1728 1595 1730
rect 1528 1727 1529 1728
rect 1523 1726 1529 1727
rect 1594 1727 1595 1728
rect 1599 1727 1600 1731
rect 1594 1726 1600 1727
rect 1602 1731 1609 1732
rect 1602 1727 1603 1731
rect 1608 1727 1609 1731
rect 1602 1726 1609 1727
rect 1690 1731 1697 1732
rect 1690 1727 1691 1731
rect 1696 1727 1697 1731
rect 1690 1726 1697 1727
rect 1786 1731 1793 1732
rect 1786 1727 1787 1731
rect 1792 1727 1793 1731
rect 1786 1726 1793 1727
rect 1874 1731 1881 1732
rect 1874 1727 1875 1731
rect 1880 1727 1881 1731
rect 1963 1729 1964 1733
rect 1968 1732 2001 1733
rect 2131 1733 2137 1734
rect 1968 1729 1969 1732
rect 1963 1728 1969 1729
rect 2050 1731 2057 1732
rect 1874 1726 1881 1727
rect 2050 1727 2051 1731
rect 2056 1727 2057 1731
rect 2131 1729 2132 1733
rect 2136 1729 2137 1733
rect 2291 1733 2297 1734
rect 2131 1728 2137 1729
rect 2206 1731 2217 1732
rect 2050 1726 2057 1727
rect 2206 1727 2207 1731
rect 2211 1727 2212 1731
rect 2216 1727 2217 1731
rect 2291 1729 2292 1733
rect 2296 1729 2297 1733
rect 2291 1728 2297 1729
rect 2371 1731 2377 1732
rect 2206 1726 2217 1727
rect 2371 1727 2372 1731
rect 2376 1730 2377 1731
rect 2402 1731 2408 1732
rect 2402 1730 2403 1731
rect 2376 1728 2403 1730
rect 2376 1727 2377 1728
rect 2371 1726 2377 1727
rect 2402 1727 2403 1728
rect 2407 1727 2408 1731
rect 2402 1726 2408 1727
rect 2435 1731 2441 1732
rect 2435 1727 2436 1731
rect 2440 1730 2441 1731
rect 2470 1731 2476 1732
rect 2470 1730 2471 1731
rect 2440 1728 2471 1730
rect 2440 1727 2441 1728
rect 2435 1726 2441 1727
rect 2470 1727 2471 1728
rect 2475 1727 2476 1731
rect 2470 1726 2476 1727
rect 147 1725 153 1726
rect 147 1721 148 1725
rect 152 1721 153 1725
rect 147 1720 153 1721
rect 190 1723 196 1724
rect 190 1719 191 1723
rect 195 1722 196 1723
rect 219 1723 225 1724
rect 219 1722 220 1723
rect 195 1720 220 1722
rect 195 1719 196 1720
rect 190 1718 196 1719
rect 219 1719 220 1720
rect 224 1719 225 1723
rect 219 1718 225 1719
rect 262 1723 268 1724
rect 262 1719 263 1723
rect 267 1722 268 1723
rect 299 1723 305 1724
rect 299 1722 300 1723
rect 267 1720 300 1722
rect 267 1719 268 1720
rect 262 1718 268 1719
rect 299 1719 300 1720
rect 304 1719 305 1723
rect 299 1718 305 1719
rect 342 1723 348 1724
rect 342 1719 343 1723
rect 347 1722 348 1723
rect 387 1723 393 1724
rect 387 1722 388 1723
rect 347 1720 388 1722
rect 347 1719 348 1720
rect 342 1718 348 1719
rect 387 1719 388 1720
rect 392 1719 393 1723
rect 387 1718 393 1719
rect 430 1723 436 1724
rect 430 1719 431 1723
rect 435 1722 436 1723
rect 483 1723 489 1724
rect 483 1722 484 1723
rect 435 1720 484 1722
rect 435 1719 436 1720
rect 430 1718 436 1719
rect 483 1719 484 1720
rect 488 1719 489 1723
rect 483 1718 489 1719
rect 586 1723 593 1724
rect 586 1719 587 1723
rect 592 1719 593 1723
rect 586 1718 593 1719
rect 691 1723 697 1724
rect 691 1719 692 1723
rect 696 1722 697 1723
rect 798 1723 809 1724
rect 696 1720 790 1722
rect 696 1719 697 1720
rect 691 1718 697 1719
rect 788 1710 790 1720
rect 798 1719 799 1723
rect 803 1719 804 1723
rect 808 1719 809 1723
rect 798 1718 809 1719
rect 910 1723 921 1724
rect 910 1719 911 1723
rect 915 1719 916 1723
rect 920 1719 921 1723
rect 910 1718 921 1719
rect 1026 1723 1033 1724
rect 1026 1719 1027 1723
rect 1032 1719 1033 1723
rect 1026 1718 1033 1719
rect 1070 1723 1076 1724
rect 1070 1719 1071 1723
rect 1075 1722 1076 1723
rect 1139 1723 1145 1724
rect 1139 1722 1140 1723
rect 1075 1720 1140 1722
rect 1075 1719 1076 1720
rect 1070 1718 1076 1719
rect 1139 1719 1140 1720
rect 1144 1719 1145 1723
rect 1139 1718 1145 1719
rect 1379 1715 1385 1716
rect 1379 1711 1380 1715
rect 1384 1714 1385 1715
rect 1414 1715 1420 1716
rect 1414 1714 1415 1715
rect 1384 1712 1415 1714
rect 1384 1711 1385 1712
rect 1379 1710 1385 1711
rect 1414 1711 1415 1712
rect 1419 1711 1420 1715
rect 1414 1710 1420 1711
rect 1422 1715 1428 1716
rect 1422 1711 1423 1715
rect 1427 1714 1428 1715
rect 1443 1715 1449 1716
rect 1443 1714 1444 1715
rect 1427 1712 1444 1714
rect 1427 1711 1428 1712
rect 1422 1710 1428 1711
rect 1443 1711 1444 1712
rect 1448 1711 1449 1715
rect 1443 1710 1449 1711
rect 1486 1715 1492 1716
rect 1486 1711 1487 1715
rect 1491 1714 1492 1715
rect 1523 1715 1529 1716
rect 1523 1714 1524 1715
rect 1491 1712 1524 1714
rect 1491 1711 1492 1712
rect 1486 1710 1492 1711
rect 1523 1711 1524 1712
rect 1528 1711 1529 1715
rect 1523 1710 1529 1711
rect 1566 1715 1572 1716
rect 1566 1711 1567 1715
rect 1571 1714 1572 1715
rect 1611 1715 1617 1716
rect 1611 1714 1612 1715
rect 1571 1712 1612 1714
rect 1571 1711 1572 1712
rect 1566 1710 1572 1711
rect 1611 1711 1612 1712
rect 1616 1711 1617 1715
rect 1611 1710 1617 1711
rect 1654 1715 1660 1716
rect 1654 1711 1655 1715
rect 1659 1714 1660 1715
rect 1707 1715 1713 1716
rect 1707 1714 1708 1715
rect 1659 1712 1708 1714
rect 1659 1711 1660 1712
rect 1654 1710 1660 1711
rect 1707 1711 1708 1712
rect 1712 1711 1713 1715
rect 1707 1710 1713 1711
rect 1750 1715 1756 1716
rect 1750 1711 1751 1715
rect 1755 1714 1756 1715
rect 1803 1715 1809 1716
rect 1803 1714 1804 1715
rect 1755 1712 1804 1714
rect 1755 1711 1756 1712
rect 1750 1710 1756 1711
rect 1803 1711 1804 1712
rect 1808 1711 1809 1715
rect 1803 1710 1809 1711
rect 1899 1715 1905 1716
rect 1899 1711 1900 1715
rect 1904 1714 1905 1715
rect 1942 1715 1948 1716
rect 1904 1712 1938 1714
rect 1904 1711 1905 1712
rect 1899 1710 1905 1711
rect 788 1708 846 1710
rect 844 1706 846 1708
rect 166 1705 172 1706
rect 110 1704 116 1705
rect 110 1700 111 1704
rect 115 1700 116 1704
rect 166 1701 167 1705
rect 171 1701 172 1705
rect 238 1705 244 1706
rect 166 1700 172 1701
rect 187 1703 196 1704
rect 110 1699 116 1700
rect 187 1699 188 1703
rect 195 1699 196 1703
rect 238 1701 239 1705
rect 243 1701 244 1705
rect 318 1705 324 1706
rect 238 1700 244 1701
rect 259 1703 268 1704
rect 187 1698 196 1699
rect 259 1699 260 1703
rect 267 1699 268 1703
rect 318 1701 319 1705
rect 323 1701 324 1705
rect 406 1705 412 1706
rect 318 1700 324 1701
rect 339 1703 348 1704
rect 259 1698 268 1699
rect 339 1699 340 1703
rect 347 1699 348 1703
rect 406 1701 407 1705
rect 411 1701 412 1705
rect 502 1705 508 1706
rect 406 1700 412 1701
rect 427 1703 436 1704
rect 339 1698 348 1699
rect 427 1699 428 1703
rect 435 1699 436 1703
rect 502 1701 503 1705
rect 507 1701 508 1705
rect 606 1705 612 1706
rect 502 1700 508 1701
rect 510 1703 516 1704
rect 427 1698 436 1699
rect 510 1699 511 1703
rect 515 1702 516 1703
rect 523 1703 529 1704
rect 523 1702 524 1703
rect 515 1700 524 1702
rect 515 1699 516 1700
rect 510 1698 516 1699
rect 523 1699 524 1700
rect 528 1699 529 1703
rect 606 1701 607 1705
rect 611 1701 612 1705
rect 710 1705 716 1706
rect 606 1700 612 1701
rect 614 1703 620 1704
rect 523 1698 529 1699
rect 614 1699 615 1703
rect 619 1702 620 1703
rect 627 1703 633 1704
rect 627 1702 628 1703
rect 619 1700 628 1702
rect 619 1699 620 1700
rect 614 1698 620 1699
rect 627 1699 628 1700
rect 632 1699 633 1703
rect 710 1701 711 1705
rect 715 1701 716 1705
rect 822 1705 828 1706
rect 710 1700 716 1701
rect 730 1703 737 1704
rect 627 1698 633 1699
rect 730 1699 731 1703
rect 736 1699 737 1703
rect 822 1701 823 1705
rect 827 1701 828 1705
rect 822 1700 828 1701
rect 843 1705 849 1706
rect 843 1701 844 1705
rect 848 1701 849 1705
rect 843 1700 849 1701
rect 934 1705 940 1706
rect 934 1701 935 1705
rect 939 1701 940 1705
rect 1046 1705 1052 1706
rect 934 1700 940 1701
rect 954 1703 961 1704
rect 730 1698 737 1699
rect 954 1699 955 1703
rect 960 1699 961 1703
rect 1046 1701 1047 1705
rect 1051 1701 1052 1705
rect 1158 1705 1164 1706
rect 1046 1700 1052 1701
rect 1067 1703 1076 1704
rect 954 1698 961 1699
rect 1067 1699 1068 1703
rect 1075 1699 1076 1703
rect 1158 1701 1159 1705
rect 1163 1701 1164 1705
rect 1286 1704 1292 1705
rect 1158 1700 1164 1701
rect 1174 1703 1185 1704
rect 1067 1698 1076 1699
rect 1174 1699 1175 1703
rect 1179 1699 1180 1703
rect 1184 1699 1185 1703
rect 1286 1700 1287 1704
rect 1291 1700 1292 1704
rect 1936 1702 1938 1712
rect 1942 1711 1943 1715
rect 1947 1714 1948 1715
rect 1995 1715 2001 1716
rect 1995 1714 1996 1715
rect 1947 1712 1996 1714
rect 1947 1711 1948 1712
rect 1942 1710 1948 1711
rect 1995 1711 1996 1712
rect 2000 1711 2001 1715
rect 1995 1710 2001 1711
rect 2090 1715 2097 1716
rect 2090 1711 2091 1715
rect 2096 1711 2097 1715
rect 2090 1710 2097 1711
rect 2134 1715 2140 1716
rect 2134 1711 2135 1715
rect 2139 1714 2140 1715
rect 2179 1715 2185 1716
rect 2179 1714 2180 1715
rect 2139 1712 2180 1714
rect 2139 1711 2140 1712
rect 2134 1710 2140 1711
rect 2179 1711 2180 1712
rect 2184 1711 2185 1715
rect 2179 1710 2185 1711
rect 2267 1715 2273 1716
rect 2267 1711 2268 1715
rect 2272 1714 2273 1715
rect 2318 1715 2324 1716
rect 2272 1712 2314 1714
rect 2272 1711 2273 1712
rect 2267 1710 2273 1711
rect 2312 1706 2314 1712
rect 2318 1711 2319 1715
rect 2323 1714 2324 1715
rect 2363 1715 2369 1716
rect 2363 1714 2364 1715
rect 2323 1712 2364 1714
rect 2323 1711 2324 1712
rect 2318 1710 2324 1711
rect 2363 1711 2364 1712
rect 2368 1711 2369 1715
rect 2363 1710 2369 1711
rect 2435 1715 2441 1716
rect 2435 1711 2436 1715
rect 2440 1714 2441 1715
rect 2462 1715 2468 1716
rect 2462 1714 2463 1715
rect 2440 1712 2463 1714
rect 2440 1711 2441 1712
rect 2435 1710 2441 1711
rect 2462 1711 2463 1712
rect 2467 1711 2468 1715
rect 2462 1710 2468 1711
rect 2474 1707 2480 1708
rect 2474 1706 2475 1707
rect 2312 1704 2475 1706
rect 2474 1703 2475 1704
rect 2479 1703 2480 1707
rect 2474 1702 2480 1703
rect 1936 1700 2222 1702
rect 1286 1699 1292 1700
rect 1174 1698 1185 1699
rect 2220 1698 2222 1700
rect 1398 1697 1404 1698
rect 1326 1696 1332 1697
rect 1326 1692 1327 1696
rect 1331 1692 1332 1696
rect 1398 1693 1399 1697
rect 1403 1693 1404 1697
rect 1462 1697 1468 1698
rect 1398 1692 1404 1693
rect 1419 1695 1428 1696
rect 1326 1691 1332 1692
rect 1419 1691 1420 1695
rect 1427 1691 1428 1695
rect 1462 1693 1463 1697
rect 1467 1693 1468 1697
rect 1542 1697 1548 1698
rect 1462 1692 1468 1693
rect 1483 1695 1492 1696
rect 1419 1690 1428 1691
rect 1483 1691 1484 1695
rect 1491 1691 1492 1695
rect 1542 1693 1543 1697
rect 1547 1693 1548 1697
rect 1630 1697 1636 1698
rect 1542 1692 1548 1693
rect 1563 1695 1572 1696
rect 1483 1690 1492 1691
rect 1563 1691 1564 1695
rect 1571 1691 1572 1695
rect 1630 1693 1631 1697
rect 1635 1693 1636 1697
rect 1726 1697 1732 1698
rect 1630 1692 1636 1693
rect 1651 1695 1660 1696
rect 1563 1690 1572 1691
rect 1651 1691 1652 1695
rect 1659 1691 1660 1695
rect 1726 1693 1727 1697
rect 1731 1693 1732 1697
rect 1822 1697 1828 1698
rect 1726 1692 1732 1693
rect 1747 1695 1756 1696
rect 1651 1690 1660 1691
rect 1747 1691 1748 1695
rect 1755 1691 1756 1695
rect 1822 1693 1823 1697
rect 1827 1693 1828 1697
rect 1918 1697 1924 1698
rect 1822 1692 1828 1693
rect 1842 1695 1849 1696
rect 1747 1690 1756 1691
rect 1842 1691 1843 1695
rect 1848 1691 1849 1695
rect 1918 1693 1919 1697
rect 1923 1693 1924 1697
rect 2014 1697 2020 1698
rect 1918 1692 1924 1693
rect 1939 1695 1948 1696
rect 1842 1690 1849 1691
rect 1939 1691 1940 1695
rect 1947 1691 1948 1695
rect 2014 1693 2015 1697
rect 2019 1693 2020 1697
rect 2110 1697 2116 1698
rect 2014 1692 2020 1693
rect 2030 1695 2041 1696
rect 1939 1690 1948 1691
rect 2030 1691 2031 1695
rect 2035 1691 2036 1695
rect 2040 1691 2041 1695
rect 2110 1693 2111 1697
rect 2115 1693 2116 1697
rect 2198 1697 2204 1698
rect 2110 1692 2116 1693
rect 2131 1695 2140 1696
rect 2030 1690 2041 1691
rect 2131 1691 2132 1695
rect 2139 1691 2140 1695
rect 2198 1693 2199 1697
rect 2203 1693 2204 1697
rect 2198 1692 2204 1693
rect 2219 1697 2225 1698
rect 2219 1693 2220 1697
rect 2224 1693 2225 1697
rect 2219 1692 2225 1693
rect 2286 1697 2292 1698
rect 2286 1693 2287 1697
rect 2291 1693 2292 1697
rect 2382 1697 2388 1698
rect 2286 1692 2292 1693
rect 2307 1695 2313 1696
rect 2131 1690 2140 1691
rect 2307 1691 2308 1695
rect 2312 1694 2313 1695
rect 2318 1695 2324 1696
rect 2318 1694 2319 1695
rect 2312 1692 2319 1694
rect 2312 1691 2313 1692
rect 2307 1690 2313 1691
rect 2318 1691 2319 1692
rect 2323 1691 2324 1695
rect 2382 1693 2383 1697
rect 2387 1693 2388 1697
rect 2454 1697 2460 1698
rect 2382 1692 2388 1693
rect 2402 1695 2409 1696
rect 2318 1690 2324 1691
rect 2402 1691 2403 1695
rect 2408 1691 2409 1695
rect 2454 1693 2455 1697
rect 2459 1693 2460 1697
rect 2502 1696 2508 1697
rect 2454 1692 2460 1693
rect 2462 1695 2468 1696
rect 2402 1690 2409 1691
rect 2462 1691 2463 1695
rect 2467 1694 2468 1695
rect 2475 1695 2481 1696
rect 2475 1694 2476 1695
rect 2467 1692 2476 1694
rect 2467 1691 2468 1692
rect 2462 1690 2468 1691
rect 2475 1691 2476 1692
rect 2480 1691 2481 1695
rect 2502 1692 2503 1696
rect 2507 1692 2508 1696
rect 2502 1691 2508 1692
rect 2475 1690 2481 1691
rect 110 1687 116 1688
rect 110 1683 111 1687
rect 115 1683 116 1687
rect 1286 1687 1292 1688
rect 110 1682 116 1683
rect 150 1684 156 1685
rect 150 1680 151 1684
rect 155 1680 156 1684
rect 150 1679 156 1680
rect 222 1684 228 1685
rect 222 1680 223 1684
rect 227 1680 228 1684
rect 222 1679 228 1680
rect 302 1684 308 1685
rect 302 1680 303 1684
rect 307 1680 308 1684
rect 302 1679 308 1680
rect 390 1684 396 1685
rect 390 1680 391 1684
rect 395 1680 396 1684
rect 390 1679 396 1680
rect 486 1684 492 1685
rect 486 1680 487 1684
rect 491 1680 492 1684
rect 486 1679 492 1680
rect 590 1684 596 1685
rect 590 1680 591 1684
rect 595 1680 596 1684
rect 590 1679 596 1680
rect 694 1684 700 1685
rect 694 1680 695 1684
rect 699 1680 700 1684
rect 694 1679 700 1680
rect 806 1684 812 1685
rect 806 1680 807 1684
rect 811 1680 812 1684
rect 806 1679 812 1680
rect 918 1684 924 1685
rect 918 1680 919 1684
rect 923 1680 924 1684
rect 918 1679 924 1680
rect 1030 1684 1036 1685
rect 1030 1680 1031 1684
rect 1035 1680 1036 1684
rect 1030 1679 1036 1680
rect 1142 1684 1148 1685
rect 1142 1680 1143 1684
rect 1147 1680 1148 1684
rect 1286 1683 1287 1687
rect 1291 1683 1292 1687
rect 1286 1682 1292 1683
rect 1142 1679 1148 1680
rect 1326 1679 1332 1680
rect 1326 1675 1327 1679
rect 1331 1675 1332 1679
rect 2502 1679 2508 1680
rect 1326 1674 1332 1675
rect 1382 1676 1388 1677
rect 1382 1672 1383 1676
rect 1387 1672 1388 1676
rect 1382 1671 1388 1672
rect 1446 1676 1452 1677
rect 1446 1672 1447 1676
rect 1451 1672 1452 1676
rect 1446 1671 1452 1672
rect 1526 1676 1532 1677
rect 1526 1672 1527 1676
rect 1531 1672 1532 1676
rect 1526 1671 1532 1672
rect 1614 1676 1620 1677
rect 1614 1672 1615 1676
rect 1619 1672 1620 1676
rect 1614 1671 1620 1672
rect 1710 1676 1716 1677
rect 1710 1672 1711 1676
rect 1715 1672 1716 1676
rect 1710 1671 1716 1672
rect 1806 1676 1812 1677
rect 1806 1672 1807 1676
rect 1811 1672 1812 1676
rect 1806 1671 1812 1672
rect 1902 1676 1908 1677
rect 1902 1672 1903 1676
rect 1907 1672 1908 1676
rect 1902 1671 1908 1672
rect 1998 1676 2004 1677
rect 1998 1672 1999 1676
rect 2003 1672 2004 1676
rect 1998 1671 2004 1672
rect 2094 1676 2100 1677
rect 2094 1672 2095 1676
rect 2099 1672 2100 1676
rect 2094 1671 2100 1672
rect 2182 1676 2188 1677
rect 2182 1672 2183 1676
rect 2187 1672 2188 1676
rect 2182 1671 2188 1672
rect 2270 1676 2276 1677
rect 2270 1672 2271 1676
rect 2275 1672 2276 1676
rect 2270 1671 2276 1672
rect 2366 1676 2372 1677
rect 2366 1672 2367 1676
rect 2371 1672 2372 1676
rect 2366 1671 2372 1672
rect 2438 1676 2444 1677
rect 2438 1672 2439 1676
rect 2443 1672 2444 1676
rect 2502 1675 2503 1679
rect 2507 1675 2508 1679
rect 2502 1674 2508 1675
rect 2438 1671 2444 1672
rect 254 1668 260 1669
rect 110 1665 116 1666
rect 110 1661 111 1665
rect 115 1661 116 1665
rect 254 1664 255 1668
rect 259 1664 260 1668
rect 254 1663 260 1664
rect 318 1668 324 1669
rect 318 1664 319 1668
rect 323 1664 324 1668
rect 318 1663 324 1664
rect 398 1668 404 1669
rect 398 1664 399 1668
rect 403 1664 404 1668
rect 398 1663 404 1664
rect 486 1668 492 1669
rect 486 1664 487 1668
rect 491 1664 492 1668
rect 486 1663 492 1664
rect 574 1668 580 1669
rect 574 1664 575 1668
rect 579 1664 580 1668
rect 574 1663 580 1664
rect 670 1668 676 1669
rect 670 1664 671 1668
rect 675 1664 676 1668
rect 670 1663 676 1664
rect 766 1668 772 1669
rect 766 1664 767 1668
rect 771 1664 772 1668
rect 766 1663 772 1664
rect 862 1668 868 1669
rect 862 1664 863 1668
rect 867 1664 868 1668
rect 862 1663 868 1664
rect 958 1668 964 1669
rect 958 1664 959 1668
rect 963 1664 964 1668
rect 958 1663 964 1664
rect 1062 1668 1068 1669
rect 1062 1664 1063 1668
rect 1067 1664 1068 1668
rect 1062 1663 1068 1664
rect 1166 1668 1172 1669
rect 1166 1664 1167 1668
rect 1171 1664 1172 1668
rect 1166 1663 1172 1664
rect 1286 1665 1292 1666
rect 110 1660 116 1661
rect 1286 1661 1287 1665
rect 1291 1661 1292 1665
rect 1286 1660 1292 1661
rect 1350 1660 1356 1661
rect 1326 1657 1332 1658
rect 1326 1653 1327 1657
rect 1331 1653 1332 1657
rect 1350 1656 1351 1660
rect 1355 1656 1356 1660
rect 1350 1655 1356 1656
rect 1406 1660 1412 1661
rect 1406 1656 1407 1660
rect 1411 1656 1412 1660
rect 1406 1655 1412 1656
rect 1494 1660 1500 1661
rect 1494 1656 1495 1660
rect 1499 1656 1500 1660
rect 1494 1655 1500 1656
rect 1582 1660 1588 1661
rect 1582 1656 1583 1660
rect 1587 1656 1588 1660
rect 1582 1655 1588 1656
rect 1678 1660 1684 1661
rect 1678 1656 1679 1660
rect 1683 1656 1684 1660
rect 1678 1655 1684 1656
rect 1782 1660 1788 1661
rect 1782 1656 1783 1660
rect 1787 1656 1788 1660
rect 1782 1655 1788 1656
rect 1894 1660 1900 1661
rect 1894 1656 1895 1660
rect 1899 1656 1900 1660
rect 1894 1655 1900 1656
rect 2022 1660 2028 1661
rect 2022 1656 2023 1660
rect 2027 1656 2028 1660
rect 2022 1655 2028 1656
rect 2158 1660 2164 1661
rect 2158 1656 2159 1660
rect 2163 1656 2164 1660
rect 2158 1655 2164 1656
rect 2302 1660 2308 1661
rect 2302 1656 2303 1660
rect 2307 1656 2308 1660
rect 2302 1655 2308 1656
rect 2438 1660 2444 1661
rect 2438 1656 2439 1660
rect 2443 1656 2444 1660
rect 2438 1655 2444 1656
rect 2502 1657 2508 1658
rect 1326 1652 1332 1653
rect 2502 1653 2503 1657
rect 2507 1653 2508 1657
rect 2502 1652 2508 1653
rect 110 1648 116 1649
rect 1286 1648 1292 1649
rect 110 1644 111 1648
rect 115 1644 116 1648
rect 110 1643 116 1644
rect 270 1647 276 1648
rect 270 1643 271 1647
rect 275 1643 276 1647
rect 270 1642 276 1643
rect 291 1647 297 1648
rect 291 1643 292 1647
rect 296 1646 297 1647
rect 314 1647 320 1648
rect 314 1646 315 1647
rect 296 1644 315 1646
rect 296 1643 297 1644
rect 291 1642 297 1643
rect 314 1643 315 1644
rect 319 1643 320 1647
rect 314 1642 320 1643
rect 334 1647 340 1648
rect 334 1643 335 1647
rect 339 1643 340 1647
rect 334 1642 340 1643
rect 355 1647 361 1648
rect 355 1643 356 1647
rect 360 1646 361 1647
rect 394 1647 400 1648
rect 394 1646 395 1647
rect 360 1644 395 1646
rect 360 1643 361 1644
rect 355 1642 361 1643
rect 394 1643 395 1644
rect 399 1643 400 1647
rect 394 1642 400 1643
rect 414 1647 420 1648
rect 414 1643 415 1647
rect 419 1643 420 1647
rect 414 1642 420 1643
rect 435 1647 441 1648
rect 435 1643 436 1647
rect 440 1646 441 1647
rect 482 1647 488 1648
rect 482 1646 483 1647
rect 440 1644 483 1646
rect 440 1643 441 1644
rect 435 1642 441 1643
rect 482 1643 483 1644
rect 487 1643 488 1647
rect 482 1642 488 1643
rect 502 1647 508 1648
rect 502 1643 503 1647
rect 507 1643 508 1647
rect 502 1642 508 1643
rect 518 1647 529 1648
rect 518 1643 519 1647
rect 523 1643 524 1647
rect 528 1643 529 1647
rect 518 1642 529 1643
rect 590 1647 596 1648
rect 590 1643 591 1647
rect 595 1643 596 1647
rect 590 1642 596 1643
rect 606 1647 617 1648
rect 606 1643 607 1647
rect 611 1643 612 1647
rect 616 1643 617 1647
rect 606 1642 617 1643
rect 686 1647 692 1648
rect 686 1643 687 1647
rect 691 1643 692 1647
rect 686 1642 692 1643
rect 707 1647 713 1648
rect 707 1643 708 1647
rect 712 1646 713 1647
rect 762 1647 768 1648
rect 762 1646 763 1647
rect 712 1644 763 1646
rect 712 1643 713 1644
rect 707 1642 713 1643
rect 762 1643 763 1644
rect 767 1643 768 1647
rect 762 1642 768 1643
rect 782 1647 788 1648
rect 782 1643 783 1647
rect 787 1643 788 1647
rect 782 1642 788 1643
rect 798 1647 809 1648
rect 798 1643 799 1647
rect 803 1643 804 1647
rect 808 1643 809 1647
rect 798 1642 809 1643
rect 878 1647 884 1648
rect 878 1643 879 1647
rect 883 1643 884 1647
rect 878 1642 884 1643
rect 899 1647 905 1648
rect 899 1643 900 1647
rect 904 1646 905 1647
rect 910 1647 916 1648
rect 910 1646 911 1647
rect 904 1644 911 1646
rect 904 1643 905 1644
rect 899 1642 905 1643
rect 910 1643 911 1644
rect 915 1643 916 1647
rect 910 1642 916 1643
rect 974 1647 980 1648
rect 974 1643 975 1647
rect 979 1643 980 1647
rect 974 1642 980 1643
rect 995 1647 1001 1648
rect 995 1643 996 1647
rect 1000 1646 1001 1647
rect 1058 1647 1064 1648
rect 1058 1646 1059 1647
rect 1000 1644 1059 1646
rect 1000 1643 1001 1644
rect 995 1642 1001 1643
rect 1058 1643 1059 1644
rect 1063 1643 1064 1647
rect 1058 1642 1064 1643
rect 1078 1647 1084 1648
rect 1078 1643 1079 1647
rect 1083 1643 1084 1647
rect 1078 1642 1084 1643
rect 1098 1647 1105 1648
rect 1098 1643 1099 1647
rect 1104 1643 1105 1647
rect 1098 1642 1105 1643
rect 1182 1647 1188 1648
rect 1182 1643 1183 1647
rect 1187 1643 1188 1647
rect 1203 1647 1209 1648
rect 1203 1646 1204 1647
rect 1182 1642 1188 1643
rect 1192 1644 1204 1646
rect 510 1635 516 1636
rect 510 1634 511 1635
rect 252 1632 511 1634
rect 252 1630 254 1632
rect 510 1631 511 1632
rect 515 1631 516 1635
rect 1192 1634 1194 1644
rect 1203 1643 1204 1644
rect 1208 1643 1209 1647
rect 1286 1644 1287 1648
rect 1291 1644 1292 1648
rect 1286 1643 1292 1644
rect 1203 1642 1209 1643
rect 1326 1640 1332 1641
rect 2502 1640 2508 1641
rect 1326 1636 1327 1640
rect 1331 1636 1332 1640
rect 1326 1635 1332 1636
rect 1366 1639 1372 1640
rect 1366 1635 1367 1639
rect 1371 1635 1372 1639
rect 1366 1634 1372 1635
rect 1387 1639 1393 1640
rect 1387 1635 1388 1639
rect 1392 1638 1393 1639
rect 1402 1639 1408 1640
rect 1402 1638 1403 1639
rect 1392 1636 1403 1638
rect 1392 1635 1393 1636
rect 1387 1634 1393 1635
rect 1402 1635 1403 1636
rect 1407 1635 1408 1639
rect 1402 1634 1408 1635
rect 1422 1639 1428 1640
rect 1422 1635 1423 1639
rect 1427 1635 1428 1639
rect 1422 1634 1428 1635
rect 1443 1639 1449 1640
rect 1443 1635 1444 1639
rect 1448 1638 1449 1639
rect 1490 1639 1496 1640
rect 1490 1638 1491 1639
rect 1448 1636 1491 1638
rect 1448 1635 1449 1636
rect 1443 1634 1449 1635
rect 1490 1635 1491 1636
rect 1495 1635 1496 1639
rect 1490 1634 1496 1635
rect 1510 1639 1516 1640
rect 1510 1635 1511 1639
rect 1515 1635 1516 1639
rect 1510 1634 1516 1635
rect 1531 1639 1537 1640
rect 1531 1635 1532 1639
rect 1536 1638 1537 1639
rect 1578 1639 1584 1640
rect 1578 1638 1579 1639
rect 1536 1636 1579 1638
rect 1536 1635 1537 1636
rect 1531 1634 1537 1635
rect 1578 1635 1579 1636
rect 1583 1635 1584 1639
rect 1578 1634 1584 1635
rect 1598 1639 1604 1640
rect 1598 1635 1599 1639
rect 1603 1635 1604 1639
rect 1598 1634 1604 1635
rect 1619 1639 1625 1640
rect 1619 1635 1620 1639
rect 1624 1638 1625 1639
rect 1674 1639 1680 1640
rect 1674 1638 1675 1639
rect 1624 1636 1675 1638
rect 1624 1635 1625 1636
rect 1619 1634 1625 1635
rect 1674 1635 1675 1636
rect 1679 1635 1680 1639
rect 1674 1634 1680 1635
rect 1694 1639 1700 1640
rect 1694 1635 1695 1639
rect 1699 1635 1700 1639
rect 1694 1634 1700 1635
rect 1702 1639 1708 1640
rect 1702 1635 1703 1639
rect 1707 1638 1708 1639
rect 1715 1639 1721 1640
rect 1715 1638 1716 1639
rect 1707 1636 1716 1638
rect 1707 1635 1708 1636
rect 1702 1634 1708 1635
rect 1715 1635 1716 1636
rect 1720 1635 1721 1639
rect 1715 1634 1721 1635
rect 1798 1639 1804 1640
rect 1798 1635 1799 1639
rect 1803 1635 1804 1639
rect 1798 1634 1804 1635
rect 1819 1639 1825 1640
rect 1819 1635 1820 1639
rect 1824 1638 1825 1639
rect 1890 1639 1896 1640
rect 1890 1638 1891 1639
rect 1824 1636 1891 1638
rect 1824 1635 1825 1636
rect 1819 1634 1825 1635
rect 1890 1635 1891 1636
rect 1895 1635 1896 1639
rect 1890 1634 1896 1635
rect 1910 1639 1916 1640
rect 1910 1635 1911 1639
rect 1915 1635 1916 1639
rect 1910 1634 1916 1635
rect 1930 1639 1937 1640
rect 1930 1635 1931 1639
rect 1936 1635 1937 1639
rect 1930 1634 1937 1635
rect 2038 1639 2044 1640
rect 2038 1635 2039 1639
rect 2043 1635 2044 1639
rect 2038 1634 2044 1635
rect 2059 1639 2065 1640
rect 2059 1635 2060 1639
rect 2064 1638 2065 1639
rect 2154 1639 2160 1640
rect 2154 1638 2155 1639
rect 2064 1636 2155 1638
rect 2064 1635 2065 1636
rect 2059 1634 2065 1635
rect 2154 1635 2155 1636
rect 2159 1635 2160 1639
rect 2154 1634 2160 1635
rect 2174 1639 2180 1640
rect 2174 1635 2175 1639
rect 2179 1635 2180 1639
rect 2174 1634 2180 1635
rect 2195 1639 2201 1640
rect 2195 1635 2196 1639
rect 2200 1638 2201 1639
rect 2298 1639 2304 1640
rect 2298 1638 2299 1639
rect 2200 1636 2299 1638
rect 2200 1635 2201 1636
rect 2195 1634 2201 1635
rect 2298 1635 2299 1636
rect 2303 1635 2304 1639
rect 2298 1634 2304 1635
rect 2318 1639 2324 1640
rect 2318 1635 2319 1639
rect 2323 1635 2324 1639
rect 2339 1639 2345 1640
rect 2339 1638 2340 1639
rect 2318 1634 2324 1635
rect 2328 1636 2340 1638
rect 510 1630 516 1631
rect 956 1632 1194 1634
rect 956 1630 958 1632
rect 2328 1630 2330 1636
rect 2339 1635 2340 1636
rect 2344 1635 2345 1639
rect 2339 1634 2345 1635
rect 2454 1639 2460 1640
rect 2454 1635 2455 1639
rect 2459 1635 2460 1639
rect 2454 1634 2460 1635
rect 2474 1639 2481 1640
rect 2474 1635 2475 1639
rect 2480 1635 2481 1639
rect 2502 1636 2503 1640
rect 2507 1636 2508 1640
rect 2502 1635 2508 1636
rect 2474 1634 2481 1635
rect 251 1629 257 1630
rect 251 1625 252 1629
rect 256 1625 257 1629
rect 955 1629 961 1630
rect 251 1624 257 1625
rect 314 1627 321 1628
rect 314 1623 315 1627
rect 320 1623 321 1627
rect 314 1622 321 1623
rect 394 1627 401 1628
rect 394 1623 395 1627
rect 400 1623 401 1627
rect 394 1622 401 1623
rect 482 1627 489 1628
rect 482 1623 483 1627
rect 488 1623 489 1627
rect 482 1622 489 1623
rect 571 1627 577 1628
rect 571 1623 572 1627
rect 576 1626 577 1627
rect 614 1627 620 1628
rect 614 1626 615 1627
rect 576 1624 615 1626
rect 576 1623 577 1624
rect 571 1622 577 1623
rect 614 1623 615 1624
rect 619 1623 620 1627
rect 614 1622 620 1623
rect 667 1627 673 1628
rect 667 1623 668 1627
rect 672 1626 673 1627
rect 754 1627 760 1628
rect 754 1626 755 1627
rect 672 1624 755 1626
rect 672 1623 673 1624
rect 667 1622 673 1623
rect 754 1623 755 1624
rect 759 1623 760 1627
rect 754 1622 760 1623
rect 762 1627 769 1628
rect 762 1623 763 1627
rect 768 1623 769 1627
rect 762 1622 769 1623
rect 859 1627 865 1628
rect 859 1623 860 1627
rect 864 1626 865 1627
rect 914 1627 920 1628
rect 914 1626 915 1627
rect 864 1624 915 1626
rect 864 1623 865 1624
rect 859 1622 865 1623
rect 914 1623 915 1624
rect 919 1623 920 1627
rect 955 1625 956 1629
rect 960 1625 961 1629
rect 1780 1628 2330 1630
rect 955 1624 961 1625
rect 1058 1627 1065 1628
rect 914 1622 920 1623
rect 1058 1623 1059 1627
rect 1064 1623 1065 1627
rect 1058 1622 1065 1623
rect 1163 1627 1169 1628
rect 1163 1623 1164 1627
rect 1168 1626 1169 1627
rect 1174 1627 1180 1628
rect 1174 1626 1175 1627
rect 1168 1624 1175 1626
rect 1168 1623 1169 1624
rect 1163 1622 1169 1623
rect 1174 1623 1175 1624
rect 1179 1623 1180 1627
rect 1174 1622 1180 1623
rect 1780 1622 1782 1628
rect 2030 1623 2036 1624
rect 2030 1622 2031 1623
rect 1779 1621 1785 1622
rect 518 1619 524 1620
rect 518 1618 519 1619
rect 284 1616 519 1618
rect 284 1614 286 1616
rect 518 1615 519 1616
rect 523 1615 524 1619
rect 518 1614 524 1615
rect 1347 1619 1353 1620
rect 1347 1615 1348 1619
rect 1352 1618 1353 1619
rect 1391 1619 1397 1620
rect 1391 1618 1392 1619
rect 1352 1616 1392 1618
rect 1352 1615 1353 1616
rect 1347 1614 1353 1615
rect 1391 1615 1392 1616
rect 1396 1615 1397 1619
rect 1391 1614 1397 1615
rect 1402 1619 1409 1620
rect 1402 1615 1403 1619
rect 1408 1615 1409 1619
rect 1402 1614 1409 1615
rect 1490 1619 1497 1620
rect 1490 1615 1491 1619
rect 1496 1615 1497 1619
rect 1490 1614 1497 1615
rect 1578 1619 1585 1620
rect 1578 1615 1579 1619
rect 1584 1615 1585 1619
rect 1578 1614 1585 1615
rect 1674 1619 1681 1620
rect 1674 1615 1675 1619
rect 1680 1615 1681 1619
rect 1779 1617 1780 1621
rect 1784 1617 1785 1621
rect 2019 1621 2031 1622
rect 1779 1616 1785 1617
rect 1890 1619 1897 1620
rect 1674 1614 1681 1615
rect 1890 1615 1891 1619
rect 1896 1615 1897 1619
rect 2019 1617 2020 1621
rect 2024 1620 2031 1621
rect 2024 1617 2025 1620
rect 2030 1619 2031 1620
rect 2035 1619 2036 1623
rect 2030 1618 2036 1619
rect 2154 1619 2161 1620
rect 2019 1616 2025 1617
rect 1890 1614 1897 1615
rect 2154 1615 2155 1619
rect 2160 1615 2161 1619
rect 2154 1614 2161 1615
rect 2298 1619 2305 1620
rect 2298 1615 2299 1619
rect 2304 1615 2305 1619
rect 2298 1614 2305 1615
rect 2435 1619 2441 1620
rect 2435 1615 2436 1619
rect 2440 1618 2441 1619
rect 2462 1619 2468 1620
rect 2462 1618 2463 1619
rect 2440 1616 2463 1618
rect 2440 1615 2441 1616
rect 2435 1614 2441 1615
rect 2462 1615 2463 1616
rect 2467 1615 2468 1619
rect 2462 1614 2468 1615
rect 283 1613 289 1614
rect 283 1609 284 1613
rect 288 1609 289 1613
rect 283 1608 289 1609
rect 326 1611 332 1612
rect 326 1607 327 1611
rect 331 1610 332 1611
rect 339 1611 345 1612
rect 339 1610 340 1611
rect 331 1608 340 1610
rect 331 1607 332 1608
rect 326 1606 332 1607
rect 339 1607 340 1608
rect 344 1607 345 1611
rect 339 1606 345 1607
rect 382 1611 388 1612
rect 382 1607 383 1611
rect 387 1610 388 1611
rect 411 1611 417 1612
rect 411 1610 412 1611
rect 387 1608 412 1610
rect 387 1607 388 1608
rect 382 1606 388 1607
rect 411 1607 412 1608
rect 416 1607 417 1611
rect 411 1606 417 1607
rect 491 1611 497 1612
rect 491 1607 492 1611
rect 496 1607 497 1611
rect 491 1606 497 1607
rect 579 1611 585 1612
rect 579 1607 580 1611
rect 584 1610 585 1611
rect 606 1611 612 1612
rect 606 1610 607 1611
rect 584 1608 607 1610
rect 584 1607 585 1608
rect 579 1606 585 1607
rect 606 1607 607 1608
rect 611 1607 612 1611
rect 606 1606 612 1607
rect 675 1611 681 1612
rect 675 1607 676 1611
rect 680 1610 681 1611
rect 706 1611 712 1612
rect 706 1610 707 1611
rect 680 1608 707 1610
rect 680 1607 681 1608
rect 675 1606 681 1607
rect 706 1607 707 1608
rect 711 1607 712 1611
rect 706 1606 712 1607
rect 718 1611 724 1612
rect 718 1607 719 1611
rect 723 1610 724 1611
rect 771 1611 777 1612
rect 771 1610 772 1611
rect 723 1608 772 1610
rect 723 1607 724 1608
rect 718 1606 724 1607
rect 771 1607 772 1608
rect 776 1607 777 1611
rect 771 1606 777 1607
rect 798 1611 804 1612
rect 798 1607 799 1611
rect 803 1610 804 1611
rect 875 1611 881 1612
rect 875 1610 876 1611
rect 803 1608 876 1610
rect 803 1607 804 1608
rect 798 1606 804 1607
rect 875 1607 876 1608
rect 880 1607 881 1611
rect 875 1606 881 1607
rect 987 1611 993 1612
rect 987 1607 988 1611
rect 992 1610 993 1611
rect 1098 1611 1105 1612
rect 992 1608 1086 1610
rect 992 1607 993 1608
rect 987 1606 993 1607
rect 254 1599 260 1600
rect 254 1595 255 1599
rect 259 1598 260 1599
rect 493 1598 495 1606
rect 754 1599 760 1600
rect 259 1596 490 1598
rect 493 1596 622 1598
rect 259 1595 260 1596
rect 254 1594 260 1595
rect 302 1593 308 1594
rect 110 1592 116 1593
rect 110 1588 111 1592
rect 115 1588 116 1592
rect 302 1589 303 1593
rect 307 1589 308 1593
rect 358 1593 364 1594
rect 302 1588 308 1589
rect 323 1591 332 1592
rect 110 1587 116 1588
rect 323 1587 324 1591
rect 331 1587 332 1591
rect 358 1589 359 1593
rect 363 1589 364 1593
rect 430 1593 436 1594
rect 358 1588 364 1589
rect 379 1591 388 1592
rect 323 1586 332 1587
rect 379 1587 380 1591
rect 387 1587 388 1591
rect 430 1589 431 1593
rect 435 1589 436 1593
rect 430 1588 436 1589
rect 451 1591 457 1592
rect 379 1586 388 1587
rect 451 1587 452 1591
rect 456 1590 457 1591
rect 478 1591 484 1592
rect 478 1590 479 1591
rect 456 1588 479 1590
rect 456 1587 457 1588
rect 451 1586 457 1587
rect 478 1587 479 1588
rect 483 1587 484 1591
rect 488 1590 490 1596
rect 620 1594 622 1596
rect 754 1595 755 1599
rect 759 1598 760 1599
rect 1084 1598 1086 1608
rect 1098 1607 1099 1611
rect 1104 1607 1105 1611
rect 1098 1606 1105 1607
rect 1262 1607 1268 1608
rect 1262 1603 1263 1607
rect 1267 1606 1268 1607
rect 1347 1607 1353 1608
rect 1347 1606 1348 1607
rect 1267 1604 1348 1606
rect 1267 1603 1268 1604
rect 1262 1602 1268 1603
rect 1347 1603 1348 1604
rect 1352 1603 1353 1607
rect 1347 1602 1353 1603
rect 1390 1607 1396 1608
rect 1390 1603 1391 1607
rect 1395 1606 1396 1607
rect 1403 1607 1409 1608
rect 1403 1606 1404 1607
rect 1395 1604 1404 1606
rect 1395 1603 1396 1604
rect 1390 1602 1396 1603
rect 1403 1603 1404 1604
rect 1408 1603 1409 1607
rect 1403 1602 1409 1603
rect 1446 1607 1452 1608
rect 1446 1603 1447 1607
rect 1451 1606 1452 1607
rect 1459 1607 1465 1608
rect 1459 1606 1460 1607
rect 1451 1604 1460 1606
rect 1451 1603 1452 1604
rect 1446 1602 1452 1603
rect 1459 1603 1460 1604
rect 1464 1603 1465 1607
rect 1459 1602 1465 1603
rect 1502 1607 1508 1608
rect 1502 1603 1503 1607
rect 1507 1606 1508 1607
rect 1539 1607 1545 1608
rect 1539 1606 1540 1607
rect 1507 1604 1540 1606
rect 1507 1603 1508 1604
rect 1502 1602 1508 1603
rect 1539 1603 1540 1604
rect 1544 1603 1545 1607
rect 1539 1602 1545 1603
rect 1582 1607 1588 1608
rect 1582 1603 1583 1607
rect 1587 1606 1588 1607
rect 1619 1607 1625 1608
rect 1619 1606 1620 1607
rect 1587 1604 1620 1606
rect 1587 1603 1588 1604
rect 1582 1602 1588 1603
rect 1619 1603 1620 1604
rect 1624 1603 1625 1607
rect 1619 1602 1625 1603
rect 1699 1607 1705 1608
rect 1699 1603 1700 1607
rect 1704 1606 1705 1607
rect 1771 1607 1777 1608
rect 1704 1604 1766 1606
rect 1704 1603 1705 1604
rect 1699 1602 1705 1603
rect 759 1596 814 1598
rect 1084 1596 1142 1598
rect 759 1595 760 1596
rect 754 1594 760 1595
rect 812 1594 814 1596
rect 1140 1594 1142 1596
rect 1391 1595 1397 1596
rect 510 1593 516 1594
rect 502 1591 508 1592
rect 502 1590 503 1591
rect 488 1588 503 1590
rect 478 1586 484 1587
rect 502 1587 503 1588
rect 507 1587 508 1591
rect 510 1589 511 1593
rect 515 1589 516 1593
rect 598 1593 604 1594
rect 510 1588 516 1589
rect 518 1591 524 1592
rect 502 1586 508 1587
rect 518 1587 519 1591
rect 523 1590 524 1591
rect 531 1591 537 1592
rect 531 1590 532 1591
rect 523 1588 532 1590
rect 523 1587 524 1588
rect 518 1586 524 1587
rect 531 1587 532 1588
rect 536 1587 537 1591
rect 598 1589 599 1593
rect 603 1589 604 1593
rect 598 1588 604 1589
rect 619 1593 625 1594
rect 619 1589 620 1593
rect 624 1589 625 1593
rect 619 1588 625 1589
rect 694 1593 700 1594
rect 694 1589 695 1593
rect 699 1589 700 1593
rect 790 1593 796 1594
rect 694 1588 700 1589
rect 715 1591 724 1592
rect 531 1586 537 1587
rect 715 1587 716 1591
rect 723 1587 724 1591
rect 790 1589 791 1593
rect 795 1589 796 1593
rect 790 1588 796 1589
rect 811 1593 817 1594
rect 811 1589 812 1593
rect 816 1589 817 1593
rect 811 1588 817 1589
rect 894 1593 900 1594
rect 894 1589 895 1593
rect 899 1589 900 1593
rect 1006 1593 1012 1594
rect 894 1588 900 1589
rect 914 1591 921 1592
rect 715 1586 724 1587
rect 914 1587 915 1591
rect 920 1587 921 1591
rect 1006 1589 1007 1593
rect 1011 1589 1012 1593
rect 1118 1593 1124 1594
rect 1006 1588 1012 1589
rect 1014 1591 1020 1592
rect 914 1586 921 1587
rect 1014 1587 1015 1591
rect 1019 1590 1020 1591
rect 1027 1591 1033 1592
rect 1027 1590 1028 1591
rect 1019 1588 1028 1590
rect 1019 1587 1020 1588
rect 1014 1586 1020 1587
rect 1027 1587 1028 1588
rect 1032 1587 1033 1591
rect 1118 1589 1119 1593
rect 1123 1589 1124 1593
rect 1118 1588 1124 1589
rect 1139 1593 1145 1594
rect 1139 1589 1140 1593
rect 1144 1589 1145 1593
rect 1139 1588 1145 1589
rect 1286 1592 1292 1593
rect 1286 1588 1287 1592
rect 1291 1588 1292 1592
rect 1391 1591 1392 1595
rect 1396 1594 1397 1595
rect 1764 1594 1766 1604
rect 1771 1603 1772 1607
rect 1776 1606 1777 1607
rect 1851 1607 1857 1608
rect 1776 1604 1846 1606
rect 1776 1603 1777 1604
rect 1771 1602 1777 1603
rect 1844 1594 1846 1604
rect 1851 1603 1852 1607
rect 1856 1606 1857 1607
rect 1930 1607 1937 1608
rect 1856 1604 1926 1606
rect 1856 1603 1857 1604
rect 1851 1602 1857 1603
rect 1924 1594 1926 1604
rect 1930 1603 1931 1607
rect 1936 1603 1937 1607
rect 1930 1602 1937 1603
rect 1974 1607 1980 1608
rect 1974 1603 1975 1607
rect 1979 1606 1980 1607
rect 2011 1607 2017 1608
rect 2011 1606 2012 1607
rect 1979 1604 2012 1606
rect 1979 1603 1980 1604
rect 1974 1602 1980 1603
rect 2011 1603 2012 1604
rect 2016 1603 2017 1607
rect 2011 1602 2017 1603
rect 1396 1592 1662 1594
rect 1764 1592 1814 1594
rect 1844 1592 1894 1594
rect 1924 1592 2054 1594
rect 1396 1591 1397 1592
rect 1391 1590 1397 1591
rect 1660 1590 1662 1592
rect 1812 1590 1814 1592
rect 1892 1590 1894 1592
rect 2052 1590 2054 1592
rect 1366 1589 1372 1590
rect 1286 1587 1292 1588
rect 1326 1588 1332 1589
rect 1027 1586 1033 1587
rect 1326 1584 1327 1588
rect 1331 1584 1332 1588
rect 1366 1585 1367 1589
rect 1371 1585 1372 1589
rect 1422 1589 1428 1590
rect 1366 1584 1372 1585
rect 1387 1587 1396 1588
rect 1326 1583 1332 1584
rect 1387 1583 1388 1587
rect 1395 1583 1396 1587
rect 1422 1585 1423 1589
rect 1427 1585 1428 1589
rect 1478 1589 1484 1590
rect 1422 1584 1428 1585
rect 1443 1587 1452 1588
rect 1387 1582 1396 1583
rect 1443 1583 1444 1587
rect 1451 1583 1452 1587
rect 1478 1585 1479 1589
rect 1483 1585 1484 1589
rect 1558 1589 1564 1590
rect 1478 1584 1484 1585
rect 1499 1587 1508 1588
rect 1443 1582 1452 1583
rect 1499 1583 1500 1587
rect 1507 1583 1508 1587
rect 1558 1585 1559 1589
rect 1563 1585 1564 1589
rect 1638 1589 1644 1590
rect 1558 1584 1564 1585
rect 1579 1587 1588 1588
rect 1499 1582 1508 1583
rect 1579 1583 1580 1587
rect 1587 1583 1588 1587
rect 1638 1585 1639 1589
rect 1643 1585 1644 1589
rect 1638 1584 1644 1585
rect 1659 1589 1665 1590
rect 1659 1585 1660 1589
rect 1664 1585 1665 1589
rect 1659 1584 1665 1585
rect 1718 1589 1724 1590
rect 1718 1585 1719 1589
rect 1723 1585 1724 1589
rect 1790 1589 1796 1590
rect 1718 1584 1724 1585
rect 1739 1587 1748 1588
rect 1579 1582 1588 1583
rect 1739 1583 1740 1587
rect 1747 1583 1748 1587
rect 1790 1585 1791 1589
rect 1795 1585 1796 1589
rect 1790 1584 1796 1585
rect 1811 1589 1817 1590
rect 1811 1585 1812 1589
rect 1816 1585 1817 1589
rect 1811 1584 1817 1585
rect 1870 1589 1876 1590
rect 1870 1585 1871 1589
rect 1875 1585 1876 1589
rect 1870 1584 1876 1585
rect 1891 1589 1897 1590
rect 1891 1585 1892 1589
rect 1896 1585 1897 1589
rect 1891 1584 1897 1585
rect 1950 1589 1956 1590
rect 1950 1585 1951 1589
rect 1955 1585 1956 1589
rect 2030 1589 2036 1590
rect 1950 1584 1956 1585
rect 1971 1587 1980 1588
rect 1739 1582 1748 1583
rect 1971 1583 1972 1587
rect 1979 1583 1980 1587
rect 2030 1585 2031 1589
rect 2035 1585 2036 1589
rect 2030 1584 2036 1585
rect 2051 1589 2057 1590
rect 2051 1585 2052 1589
rect 2056 1585 2057 1589
rect 2051 1584 2057 1585
rect 2502 1588 2508 1589
rect 2502 1584 2503 1588
rect 2507 1584 2508 1588
rect 2502 1583 2508 1584
rect 1971 1582 1980 1583
rect 110 1575 116 1576
rect 110 1571 111 1575
rect 115 1571 116 1575
rect 1286 1575 1292 1576
rect 110 1570 116 1571
rect 286 1572 292 1573
rect 286 1568 287 1572
rect 291 1568 292 1572
rect 286 1567 292 1568
rect 342 1572 348 1573
rect 342 1568 343 1572
rect 347 1568 348 1572
rect 342 1567 348 1568
rect 414 1572 420 1573
rect 414 1568 415 1572
rect 419 1568 420 1572
rect 414 1567 420 1568
rect 494 1572 500 1573
rect 494 1568 495 1572
rect 499 1568 500 1572
rect 494 1567 500 1568
rect 582 1572 588 1573
rect 582 1568 583 1572
rect 587 1568 588 1572
rect 582 1567 588 1568
rect 678 1572 684 1573
rect 678 1568 679 1572
rect 683 1568 684 1572
rect 678 1567 684 1568
rect 774 1572 780 1573
rect 774 1568 775 1572
rect 779 1568 780 1572
rect 774 1567 780 1568
rect 878 1572 884 1573
rect 878 1568 879 1572
rect 883 1568 884 1572
rect 878 1567 884 1568
rect 990 1572 996 1573
rect 990 1568 991 1572
rect 995 1568 996 1572
rect 990 1567 996 1568
rect 1102 1572 1108 1573
rect 1102 1568 1103 1572
rect 1107 1568 1108 1572
rect 1286 1571 1287 1575
rect 1291 1571 1292 1575
rect 1286 1570 1292 1571
rect 1326 1571 1332 1572
rect 1102 1567 1108 1568
rect 1326 1567 1327 1571
rect 1331 1567 1332 1571
rect 2502 1571 2508 1572
rect 1326 1566 1332 1567
rect 1350 1568 1356 1569
rect 1350 1564 1351 1568
rect 1355 1564 1356 1568
rect 1350 1563 1356 1564
rect 1406 1568 1412 1569
rect 1406 1564 1407 1568
rect 1411 1564 1412 1568
rect 1406 1563 1412 1564
rect 1462 1568 1468 1569
rect 1462 1564 1463 1568
rect 1467 1564 1468 1568
rect 1462 1563 1468 1564
rect 1542 1568 1548 1569
rect 1542 1564 1543 1568
rect 1547 1564 1548 1568
rect 1542 1563 1548 1564
rect 1622 1568 1628 1569
rect 1622 1564 1623 1568
rect 1627 1564 1628 1568
rect 1622 1563 1628 1564
rect 1702 1568 1708 1569
rect 1702 1564 1703 1568
rect 1707 1564 1708 1568
rect 1702 1563 1708 1564
rect 1774 1568 1780 1569
rect 1774 1564 1775 1568
rect 1779 1564 1780 1568
rect 1774 1563 1780 1564
rect 1854 1568 1860 1569
rect 1854 1564 1855 1568
rect 1859 1564 1860 1568
rect 1854 1563 1860 1564
rect 1934 1568 1940 1569
rect 1934 1564 1935 1568
rect 1939 1564 1940 1568
rect 1934 1563 1940 1564
rect 2014 1568 2020 1569
rect 2014 1564 2015 1568
rect 2019 1564 2020 1568
rect 2502 1567 2503 1571
rect 2507 1567 2508 1571
rect 2502 1566 2508 1567
rect 2014 1563 2020 1564
rect 246 1560 252 1561
rect 110 1557 116 1558
rect 110 1553 111 1557
rect 115 1553 116 1557
rect 246 1556 247 1560
rect 251 1556 252 1560
rect 246 1555 252 1556
rect 318 1560 324 1561
rect 318 1556 319 1560
rect 323 1556 324 1560
rect 318 1555 324 1556
rect 398 1560 404 1561
rect 398 1556 399 1560
rect 403 1556 404 1560
rect 398 1555 404 1556
rect 486 1560 492 1561
rect 486 1556 487 1560
rect 491 1556 492 1560
rect 486 1555 492 1556
rect 582 1560 588 1561
rect 582 1556 583 1560
rect 587 1556 588 1560
rect 582 1555 588 1556
rect 670 1560 676 1561
rect 670 1556 671 1560
rect 675 1556 676 1560
rect 670 1555 676 1556
rect 758 1560 764 1561
rect 758 1556 759 1560
rect 763 1556 764 1560
rect 758 1555 764 1556
rect 846 1560 852 1561
rect 846 1556 847 1560
rect 851 1556 852 1560
rect 846 1555 852 1556
rect 926 1560 932 1561
rect 926 1556 927 1560
rect 931 1556 932 1560
rect 926 1555 932 1556
rect 1006 1560 1012 1561
rect 1006 1556 1007 1560
rect 1011 1556 1012 1560
rect 1006 1555 1012 1556
rect 1086 1560 1092 1561
rect 1086 1556 1087 1560
rect 1091 1556 1092 1560
rect 1086 1555 1092 1556
rect 1166 1560 1172 1561
rect 1166 1556 1167 1560
rect 1171 1556 1172 1560
rect 1166 1555 1172 1556
rect 1222 1560 1228 1561
rect 1222 1556 1223 1560
rect 1227 1556 1228 1560
rect 1222 1555 1228 1556
rect 1286 1557 1292 1558
rect 110 1552 116 1553
rect 1286 1553 1287 1557
rect 1291 1553 1292 1557
rect 1350 1556 1356 1557
rect 1286 1552 1292 1553
rect 1326 1553 1332 1554
rect 1326 1549 1327 1553
rect 1331 1549 1332 1553
rect 1350 1552 1351 1556
rect 1355 1552 1356 1556
rect 1350 1551 1356 1552
rect 1470 1556 1476 1557
rect 1470 1552 1471 1556
rect 1475 1552 1476 1556
rect 1470 1551 1476 1552
rect 1606 1556 1612 1557
rect 1606 1552 1607 1556
rect 1611 1552 1612 1556
rect 1606 1551 1612 1552
rect 1734 1556 1740 1557
rect 1734 1552 1735 1556
rect 1739 1552 1740 1556
rect 1734 1551 1740 1552
rect 1870 1556 1876 1557
rect 1870 1552 1871 1556
rect 1875 1552 1876 1556
rect 1870 1551 1876 1552
rect 2006 1556 2012 1557
rect 2006 1552 2007 1556
rect 2011 1552 2012 1556
rect 2006 1551 2012 1552
rect 2502 1553 2508 1554
rect 1326 1548 1332 1549
rect 2502 1549 2503 1553
rect 2507 1549 2508 1553
rect 2502 1548 2508 1549
rect 110 1540 116 1541
rect 1286 1540 1292 1541
rect 110 1536 111 1540
rect 115 1536 116 1540
rect 110 1535 116 1536
rect 262 1539 268 1540
rect 262 1535 263 1539
rect 267 1535 268 1539
rect 262 1534 268 1535
rect 270 1539 276 1540
rect 270 1535 271 1539
rect 275 1538 276 1539
rect 283 1539 289 1540
rect 283 1538 284 1539
rect 275 1536 284 1538
rect 275 1535 276 1536
rect 270 1534 276 1535
rect 283 1535 284 1536
rect 288 1535 289 1539
rect 283 1534 289 1535
rect 334 1539 340 1540
rect 334 1535 335 1539
rect 339 1535 340 1539
rect 334 1534 340 1535
rect 350 1539 361 1540
rect 350 1535 351 1539
rect 355 1535 356 1539
rect 360 1535 361 1539
rect 350 1534 361 1535
rect 414 1539 420 1540
rect 414 1535 415 1539
rect 419 1535 420 1539
rect 435 1539 441 1540
rect 435 1538 436 1539
rect 414 1534 420 1535
rect 424 1536 436 1538
rect 424 1530 426 1536
rect 435 1535 436 1536
rect 440 1535 441 1539
rect 435 1534 441 1535
rect 502 1539 508 1540
rect 502 1535 503 1539
rect 507 1535 508 1539
rect 502 1534 508 1535
rect 523 1539 529 1540
rect 523 1535 524 1539
rect 528 1538 529 1539
rect 578 1539 584 1540
rect 578 1538 579 1539
rect 528 1536 579 1538
rect 528 1535 529 1536
rect 523 1534 529 1535
rect 578 1535 579 1536
rect 583 1535 584 1539
rect 578 1534 584 1535
rect 598 1539 604 1540
rect 598 1535 599 1539
rect 603 1535 604 1539
rect 619 1539 625 1540
rect 619 1538 620 1539
rect 598 1534 604 1535
rect 608 1536 620 1538
rect 319 1528 426 1530
rect 319 1522 321 1528
rect 608 1526 610 1536
rect 619 1535 620 1536
rect 624 1535 625 1539
rect 619 1534 625 1535
rect 686 1539 692 1540
rect 686 1535 687 1539
rect 691 1535 692 1539
rect 686 1534 692 1535
rect 706 1539 713 1540
rect 706 1535 707 1539
rect 712 1535 713 1539
rect 706 1534 713 1535
rect 774 1539 780 1540
rect 774 1535 775 1539
rect 779 1535 780 1539
rect 774 1534 780 1535
rect 795 1539 804 1540
rect 795 1535 796 1539
rect 803 1535 804 1539
rect 795 1534 804 1535
rect 862 1539 868 1540
rect 862 1535 863 1539
rect 867 1535 868 1539
rect 862 1534 868 1535
rect 878 1539 889 1540
rect 878 1535 879 1539
rect 883 1535 884 1539
rect 888 1535 889 1539
rect 878 1534 889 1535
rect 942 1539 948 1540
rect 942 1535 943 1539
rect 947 1535 948 1539
rect 963 1539 969 1540
rect 963 1538 964 1539
rect 942 1534 948 1535
rect 952 1536 964 1538
rect 952 1530 954 1536
rect 963 1535 964 1536
rect 968 1535 969 1539
rect 963 1534 969 1535
rect 1022 1539 1028 1540
rect 1022 1535 1023 1539
rect 1027 1535 1028 1539
rect 1043 1539 1049 1540
rect 1043 1538 1044 1539
rect 1022 1534 1028 1535
rect 1032 1536 1044 1538
rect 397 1524 610 1526
rect 844 1528 954 1530
rect 397 1522 399 1524
rect 844 1522 846 1528
rect 1032 1526 1034 1536
rect 1043 1535 1044 1536
rect 1048 1535 1049 1539
rect 1043 1534 1049 1535
rect 1102 1539 1108 1540
rect 1102 1535 1103 1539
rect 1107 1535 1108 1539
rect 1102 1534 1108 1535
rect 1123 1539 1129 1540
rect 1123 1535 1124 1539
rect 1128 1538 1129 1539
rect 1162 1539 1168 1540
rect 1162 1538 1163 1539
rect 1128 1536 1163 1538
rect 1128 1535 1129 1536
rect 1123 1534 1129 1535
rect 1162 1535 1163 1536
rect 1167 1535 1168 1539
rect 1162 1534 1168 1535
rect 1182 1539 1188 1540
rect 1182 1535 1183 1539
rect 1187 1535 1188 1539
rect 1182 1534 1188 1535
rect 1203 1539 1209 1540
rect 1203 1535 1204 1539
rect 1208 1538 1209 1539
rect 1218 1539 1224 1540
rect 1218 1538 1219 1539
rect 1208 1536 1219 1538
rect 1208 1535 1209 1536
rect 1203 1534 1209 1535
rect 1218 1535 1219 1536
rect 1223 1535 1224 1539
rect 1218 1534 1224 1535
rect 1238 1539 1244 1540
rect 1238 1535 1239 1539
rect 1243 1535 1244 1539
rect 1238 1534 1244 1535
rect 1259 1539 1268 1540
rect 1259 1535 1260 1539
rect 1267 1535 1268 1539
rect 1286 1536 1287 1540
rect 1291 1536 1292 1540
rect 1286 1535 1292 1536
rect 1326 1536 1332 1537
rect 2502 1536 2508 1537
rect 1259 1534 1268 1535
rect 1326 1532 1327 1536
rect 1331 1532 1332 1536
rect 1326 1531 1332 1532
rect 1366 1535 1372 1536
rect 1366 1531 1367 1535
rect 1371 1531 1372 1535
rect 1387 1535 1393 1536
rect 1387 1534 1388 1535
rect 1366 1530 1372 1531
rect 1376 1532 1388 1534
rect 1376 1526 1378 1532
rect 1387 1531 1388 1532
rect 1392 1531 1393 1535
rect 1387 1530 1393 1531
rect 1486 1535 1492 1536
rect 1486 1531 1487 1535
rect 1491 1531 1492 1535
rect 1486 1530 1492 1531
rect 1507 1535 1513 1536
rect 1507 1531 1508 1535
rect 1512 1534 1513 1535
rect 1602 1535 1608 1536
rect 1602 1534 1603 1535
rect 1512 1532 1603 1534
rect 1512 1531 1513 1532
rect 1507 1530 1513 1531
rect 1602 1531 1603 1532
rect 1607 1531 1608 1535
rect 1602 1530 1608 1531
rect 1622 1535 1628 1536
rect 1622 1531 1623 1535
rect 1627 1531 1628 1535
rect 1622 1530 1628 1531
rect 1643 1535 1649 1536
rect 1643 1531 1644 1535
rect 1648 1534 1649 1535
rect 1730 1535 1736 1536
rect 1730 1534 1731 1535
rect 1648 1532 1731 1534
rect 1648 1531 1649 1532
rect 1643 1530 1649 1531
rect 1730 1531 1731 1532
rect 1735 1531 1736 1535
rect 1730 1530 1736 1531
rect 1750 1535 1756 1536
rect 1750 1531 1751 1535
rect 1755 1531 1756 1535
rect 1750 1530 1756 1531
rect 1771 1535 1777 1536
rect 1771 1531 1772 1535
rect 1776 1534 1777 1535
rect 1862 1535 1868 1536
rect 1862 1534 1863 1535
rect 1776 1532 1863 1534
rect 1776 1531 1777 1532
rect 1771 1530 1777 1531
rect 1862 1531 1863 1532
rect 1867 1531 1868 1535
rect 1862 1530 1868 1531
rect 1886 1535 1892 1536
rect 1886 1531 1887 1535
rect 1891 1531 1892 1535
rect 1886 1530 1892 1531
rect 1907 1535 1913 1536
rect 1907 1531 1908 1535
rect 1912 1534 1913 1535
rect 2002 1535 2008 1536
rect 2002 1534 2003 1535
rect 1912 1532 2003 1534
rect 1912 1531 1913 1532
rect 1907 1530 1913 1531
rect 2002 1531 2003 1532
rect 2007 1531 2008 1535
rect 2002 1530 2008 1531
rect 2022 1535 2028 1536
rect 2022 1531 2023 1535
rect 2027 1531 2028 1535
rect 2043 1535 2049 1536
rect 2043 1534 2044 1535
rect 2022 1530 2028 1531
rect 2032 1532 2044 1534
rect 924 1524 1034 1526
rect 1084 1524 1378 1526
rect 1774 1527 1780 1528
rect 924 1522 926 1524
rect 1084 1522 1086 1524
rect 1742 1523 1748 1524
rect 1742 1522 1743 1523
rect 315 1521 321 1522
rect 243 1519 249 1520
rect 243 1515 244 1519
rect 248 1518 249 1519
rect 254 1519 260 1520
rect 254 1518 255 1519
rect 248 1516 255 1518
rect 248 1515 249 1516
rect 243 1514 249 1515
rect 254 1515 255 1516
rect 259 1515 260 1519
rect 315 1517 316 1521
rect 320 1517 321 1521
rect 315 1516 321 1517
rect 395 1521 401 1522
rect 395 1517 396 1521
rect 400 1517 401 1521
rect 843 1521 849 1522
rect 395 1516 401 1517
rect 478 1519 489 1520
rect 254 1514 260 1515
rect 478 1515 479 1519
rect 483 1515 484 1519
rect 488 1515 489 1519
rect 478 1514 489 1515
rect 578 1519 585 1520
rect 578 1515 579 1519
rect 584 1515 585 1519
rect 578 1514 585 1515
rect 667 1519 676 1520
rect 667 1515 668 1519
rect 675 1515 676 1519
rect 667 1514 676 1515
rect 754 1519 761 1520
rect 754 1515 755 1519
rect 760 1515 761 1519
rect 843 1517 844 1521
rect 848 1517 849 1521
rect 843 1516 849 1517
rect 923 1521 929 1522
rect 923 1517 924 1521
rect 928 1517 929 1521
rect 1083 1521 1089 1522
rect 923 1516 929 1517
rect 1003 1519 1009 1520
rect 754 1514 761 1515
rect 1003 1515 1004 1519
rect 1008 1518 1009 1519
rect 1014 1519 1020 1520
rect 1014 1518 1015 1519
rect 1008 1516 1015 1518
rect 1008 1515 1009 1516
rect 1003 1514 1009 1515
rect 1014 1515 1015 1516
rect 1019 1515 1020 1519
rect 1083 1517 1084 1521
rect 1088 1517 1089 1521
rect 1468 1520 1743 1522
rect 1083 1516 1089 1517
rect 1162 1519 1169 1520
rect 1014 1514 1020 1515
rect 1162 1515 1163 1519
rect 1168 1515 1169 1519
rect 1162 1514 1169 1515
rect 1218 1519 1225 1520
rect 1218 1515 1219 1519
rect 1224 1515 1225 1519
rect 1468 1518 1470 1520
rect 1742 1519 1743 1520
rect 1747 1519 1748 1523
rect 1774 1523 1775 1527
rect 1779 1526 1780 1527
rect 2032 1526 2034 1532
rect 2043 1531 2044 1532
rect 2048 1531 2049 1535
rect 2502 1532 2503 1536
rect 2507 1532 2508 1536
rect 2502 1531 2508 1532
rect 2043 1530 2049 1531
rect 1779 1524 2034 1526
rect 1779 1523 1780 1524
rect 1774 1522 1780 1523
rect 1742 1518 1748 1519
rect 1467 1517 1473 1518
rect 1218 1514 1225 1515
rect 1347 1515 1353 1516
rect 1347 1511 1348 1515
rect 1352 1514 1353 1515
rect 1386 1515 1392 1516
rect 1386 1514 1387 1515
rect 1352 1512 1387 1514
rect 1352 1511 1353 1512
rect 1347 1510 1353 1511
rect 1386 1511 1387 1512
rect 1391 1511 1392 1515
rect 1467 1513 1468 1517
rect 1472 1513 1473 1517
rect 1467 1512 1473 1513
rect 1602 1515 1609 1516
rect 1386 1510 1392 1511
rect 1602 1511 1603 1515
rect 1608 1511 1609 1515
rect 1602 1510 1609 1511
rect 1730 1515 1737 1516
rect 1730 1511 1731 1515
rect 1736 1511 1737 1515
rect 1730 1510 1737 1511
rect 1862 1515 1873 1516
rect 1862 1511 1863 1515
rect 1867 1511 1868 1515
rect 1872 1511 1873 1515
rect 1862 1510 1873 1511
rect 2002 1515 2009 1516
rect 2002 1511 2003 1515
rect 2008 1511 2009 1515
rect 2002 1510 2009 1511
rect 1347 1503 1353 1504
rect 259 1499 265 1500
rect 259 1495 260 1499
rect 264 1498 265 1499
rect 270 1499 276 1500
rect 270 1498 271 1499
rect 264 1496 271 1498
rect 264 1495 265 1496
rect 259 1494 265 1495
rect 270 1495 271 1496
rect 275 1495 276 1499
rect 270 1494 276 1495
rect 323 1499 329 1500
rect 323 1495 324 1499
rect 328 1498 329 1499
rect 350 1499 356 1500
rect 350 1498 351 1499
rect 328 1496 351 1498
rect 328 1495 329 1496
rect 323 1494 329 1495
rect 350 1495 351 1496
rect 355 1495 356 1499
rect 350 1494 356 1495
rect 366 1499 372 1500
rect 366 1495 367 1499
rect 371 1498 372 1499
rect 395 1499 401 1500
rect 395 1498 396 1499
rect 371 1496 396 1498
rect 371 1495 372 1496
rect 366 1494 372 1495
rect 395 1495 396 1496
rect 400 1495 401 1499
rect 395 1494 401 1495
rect 438 1499 444 1500
rect 438 1495 439 1499
rect 443 1498 444 1499
rect 475 1499 481 1500
rect 475 1498 476 1499
rect 443 1496 476 1498
rect 443 1495 444 1496
rect 438 1494 444 1495
rect 475 1495 476 1496
rect 480 1495 481 1499
rect 475 1494 481 1495
rect 555 1499 561 1500
rect 555 1495 556 1499
rect 560 1498 561 1499
rect 606 1499 612 1500
rect 560 1496 602 1498
rect 560 1495 561 1496
rect 555 1494 561 1495
rect 600 1490 602 1496
rect 606 1495 607 1499
rect 611 1498 612 1499
rect 635 1499 641 1500
rect 635 1498 636 1499
rect 611 1496 636 1498
rect 611 1495 612 1496
rect 606 1494 612 1495
rect 635 1495 636 1496
rect 640 1495 641 1499
rect 635 1494 641 1495
rect 715 1499 721 1500
rect 715 1495 716 1499
rect 720 1495 721 1499
rect 715 1494 721 1495
rect 795 1499 801 1500
rect 795 1495 796 1499
rect 800 1498 801 1499
rect 850 1499 856 1500
rect 850 1498 851 1499
rect 800 1496 851 1498
rect 800 1495 801 1496
rect 795 1494 801 1495
rect 850 1495 851 1496
rect 855 1495 856 1499
rect 850 1494 856 1495
rect 875 1499 884 1500
rect 875 1495 876 1499
rect 883 1495 884 1499
rect 875 1494 884 1495
rect 934 1499 940 1500
rect 934 1495 935 1499
rect 939 1498 940 1499
rect 955 1499 961 1500
rect 955 1498 956 1499
rect 939 1496 956 1498
rect 939 1495 940 1496
rect 934 1494 940 1495
rect 955 1495 956 1496
rect 960 1495 961 1499
rect 955 1494 961 1495
rect 998 1499 1004 1500
rect 998 1495 999 1499
rect 1003 1498 1004 1499
rect 1035 1499 1041 1500
rect 1035 1498 1036 1499
rect 1003 1496 1036 1498
rect 1003 1495 1004 1496
rect 998 1494 1004 1495
rect 1035 1495 1036 1496
rect 1040 1495 1041 1499
rect 1035 1494 1041 1495
rect 1078 1499 1084 1500
rect 1078 1495 1079 1499
rect 1083 1498 1084 1499
rect 1123 1499 1129 1500
rect 1123 1498 1124 1499
rect 1083 1496 1124 1498
rect 1083 1495 1084 1496
rect 1078 1494 1084 1495
rect 1123 1495 1124 1496
rect 1128 1495 1129 1499
rect 1347 1499 1348 1503
rect 1352 1502 1353 1503
rect 1403 1503 1409 1504
rect 1352 1500 1398 1502
rect 1352 1499 1353 1500
rect 1347 1498 1353 1499
rect 1123 1494 1129 1495
rect 630 1491 636 1492
rect 630 1490 631 1491
rect 600 1488 631 1490
rect 630 1487 631 1488
rect 635 1487 636 1491
rect 630 1486 636 1487
rect 717 1486 719 1494
rect 1396 1490 1398 1500
rect 1403 1499 1404 1503
rect 1408 1502 1409 1503
rect 1459 1503 1465 1504
rect 1408 1500 1454 1502
rect 1408 1499 1409 1500
rect 1403 1498 1409 1499
rect 1452 1490 1454 1500
rect 1459 1499 1460 1503
rect 1464 1502 1465 1503
rect 1531 1503 1537 1504
rect 1464 1500 1526 1502
rect 1464 1499 1465 1500
rect 1459 1498 1465 1499
rect 1524 1490 1526 1500
rect 1531 1499 1532 1503
rect 1536 1502 1537 1503
rect 1566 1503 1572 1504
rect 1566 1502 1567 1503
rect 1536 1500 1567 1502
rect 1536 1499 1537 1500
rect 1531 1498 1537 1499
rect 1566 1499 1567 1500
rect 1571 1499 1572 1503
rect 1566 1498 1572 1499
rect 1574 1503 1580 1504
rect 1574 1499 1575 1503
rect 1579 1502 1580 1503
rect 1611 1503 1617 1504
rect 1611 1502 1612 1503
rect 1579 1500 1612 1502
rect 1579 1499 1580 1500
rect 1574 1498 1580 1499
rect 1611 1499 1612 1500
rect 1616 1499 1617 1503
rect 1611 1498 1617 1499
rect 1654 1503 1660 1504
rect 1654 1499 1655 1503
rect 1659 1502 1660 1503
rect 1691 1503 1697 1504
rect 1691 1502 1692 1503
rect 1659 1500 1692 1502
rect 1659 1499 1660 1500
rect 1654 1498 1660 1499
rect 1691 1499 1692 1500
rect 1696 1499 1697 1503
rect 1691 1498 1697 1499
rect 1771 1503 1780 1504
rect 1771 1499 1772 1503
rect 1779 1499 1780 1503
rect 1771 1498 1780 1499
rect 1814 1503 1820 1504
rect 1814 1499 1815 1503
rect 1819 1502 1820 1503
rect 1851 1503 1857 1504
rect 1851 1502 1852 1503
rect 1819 1500 1852 1502
rect 1819 1499 1820 1500
rect 1814 1498 1820 1499
rect 1851 1499 1852 1500
rect 1856 1499 1857 1503
rect 1851 1498 1857 1499
rect 1894 1503 1900 1504
rect 1894 1499 1895 1503
rect 1899 1502 1900 1503
rect 1931 1503 1937 1504
rect 1931 1502 1932 1503
rect 1899 1500 1932 1502
rect 1899 1499 1900 1500
rect 1894 1498 1900 1499
rect 1931 1499 1932 1500
rect 1936 1499 1937 1503
rect 1931 1498 1937 1499
rect 1974 1503 1980 1504
rect 1974 1499 1975 1503
rect 1979 1502 1980 1503
rect 2011 1503 2017 1504
rect 2011 1502 2012 1503
rect 1979 1500 2012 1502
rect 1979 1499 1980 1500
rect 1974 1498 1980 1499
rect 2011 1499 2012 1500
rect 2016 1499 2017 1503
rect 2011 1498 2017 1499
rect 2054 1503 2060 1504
rect 2054 1499 2055 1503
rect 2059 1502 2060 1503
rect 2099 1503 2105 1504
rect 2099 1502 2100 1503
rect 2059 1500 2100 1502
rect 2059 1499 2060 1500
rect 2054 1498 2060 1499
rect 2099 1499 2100 1500
rect 2104 1499 2105 1503
rect 2099 1498 2105 1499
rect 1822 1491 1828 1492
rect 1396 1488 1446 1490
rect 1452 1488 1502 1490
rect 1524 1488 1734 1490
rect 1444 1486 1446 1488
rect 1500 1486 1502 1488
rect 1732 1486 1734 1488
rect 1822 1487 1823 1491
rect 1827 1490 1828 1491
rect 1827 1488 2142 1490
rect 1827 1487 1828 1488
rect 1822 1486 1828 1487
rect 2140 1486 2142 1488
rect 717 1484 831 1486
rect 1366 1485 1372 1486
rect 829 1482 831 1484
rect 1326 1484 1332 1485
rect 278 1481 284 1482
rect 110 1480 116 1481
rect 110 1476 111 1480
rect 115 1476 116 1480
rect 278 1477 279 1481
rect 283 1477 284 1481
rect 342 1481 348 1482
rect 278 1476 284 1477
rect 286 1479 292 1480
rect 110 1475 116 1476
rect 286 1475 287 1479
rect 291 1478 292 1479
rect 299 1479 305 1480
rect 299 1478 300 1479
rect 291 1476 300 1478
rect 291 1475 292 1476
rect 286 1474 292 1475
rect 299 1475 300 1476
rect 304 1475 305 1479
rect 342 1477 343 1481
rect 347 1477 348 1481
rect 414 1481 420 1482
rect 342 1476 348 1477
rect 363 1479 372 1480
rect 299 1474 305 1475
rect 363 1475 364 1479
rect 371 1475 372 1479
rect 414 1477 415 1481
rect 419 1477 420 1481
rect 494 1481 500 1482
rect 414 1476 420 1477
rect 435 1479 444 1480
rect 363 1474 372 1475
rect 435 1475 436 1479
rect 443 1475 444 1479
rect 494 1477 495 1481
rect 499 1477 500 1481
rect 574 1481 580 1482
rect 494 1476 500 1477
rect 510 1479 521 1480
rect 435 1474 444 1475
rect 510 1475 511 1479
rect 515 1475 516 1479
rect 520 1475 521 1479
rect 574 1477 575 1481
rect 579 1477 580 1481
rect 654 1481 660 1482
rect 574 1476 580 1477
rect 595 1479 601 1480
rect 510 1474 521 1475
rect 595 1475 596 1479
rect 600 1478 601 1479
rect 606 1479 612 1480
rect 606 1478 607 1479
rect 600 1476 607 1478
rect 600 1475 601 1476
rect 595 1474 601 1475
rect 606 1475 607 1476
rect 611 1475 612 1479
rect 654 1477 655 1481
rect 659 1477 660 1481
rect 734 1481 740 1482
rect 654 1476 660 1477
rect 670 1479 681 1480
rect 606 1474 612 1475
rect 670 1475 671 1479
rect 675 1475 676 1479
rect 680 1475 681 1479
rect 734 1477 735 1481
rect 739 1477 740 1481
rect 814 1481 820 1482
rect 734 1476 740 1477
rect 754 1479 761 1480
rect 670 1474 681 1475
rect 754 1475 755 1479
rect 760 1475 761 1479
rect 814 1477 815 1481
rect 819 1477 820 1481
rect 829 1481 841 1482
rect 829 1480 836 1481
rect 814 1476 820 1477
rect 835 1477 836 1480
rect 840 1477 841 1481
rect 835 1476 841 1477
rect 894 1481 900 1482
rect 894 1477 895 1481
rect 899 1477 900 1481
rect 974 1481 980 1482
rect 894 1476 900 1477
rect 915 1479 921 1480
rect 754 1474 761 1475
rect 915 1475 916 1479
rect 920 1478 921 1479
rect 934 1479 940 1480
rect 934 1478 935 1479
rect 920 1476 935 1478
rect 920 1475 921 1476
rect 915 1474 921 1475
rect 934 1475 935 1476
rect 939 1475 940 1479
rect 974 1477 975 1481
rect 979 1477 980 1481
rect 1054 1481 1060 1482
rect 974 1476 980 1477
rect 995 1479 1004 1480
rect 934 1474 940 1475
rect 995 1475 996 1479
rect 1003 1475 1004 1479
rect 1054 1477 1055 1481
rect 1059 1477 1060 1481
rect 1142 1481 1148 1482
rect 1054 1476 1060 1477
rect 1075 1479 1084 1480
rect 995 1474 1004 1475
rect 1075 1475 1076 1479
rect 1083 1475 1084 1479
rect 1142 1477 1143 1481
rect 1147 1477 1148 1481
rect 1286 1480 1292 1481
rect 1142 1476 1148 1477
rect 1150 1479 1156 1480
rect 1075 1474 1084 1475
rect 1150 1475 1151 1479
rect 1155 1478 1156 1479
rect 1163 1479 1169 1480
rect 1163 1478 1164 1479
rect 1155 1476 1164 1478
rect 1155 1475 1156 1476
rect 1150 1474 1156 1475
rect 1163 1475 1164 1476
rect 1168 1475 1169 1479
rect 1286 1476 1287 1480
rect 1291 1476 1292 1480
rect 1326 1480 1327 1484
rect 1331 1480 1332 1484
rect 1366 1481 1367 1485
rect 1371 1481 1372 1485
rect 1422 1485 1428 1486
rect 1366 1480 1372 1481
rect 1386 1483 1393 1484
rect 1326 1479 1332 1480
rect 1386 1479 1387 1483
rect 1392 1479 1393 1483
rect 1422 1481 1423 1485
rect 1427 1481 1428 1485
rect 1422 1480 1428 1481
rect 1443 1485 1449 1486
rect 1443 1481 1444 1485
rect 1448 1481 1449 1485
rect 1443 1480 1449 1481
rect 1478 1485 1484 1486
rect 1478 1481 1479 1485
rect 1483 1481 1484 1485
rect 1478 1480 1484 1481
rect 1499 1485 1505 1486
rect 1499 1481 1500 1485
rect 1504 1481 1505 1485
rect 1499 1480 1505 1481
rect 1550 1485 1556 1486
rect 1550 1481 1551 1485
rect 1555 1481 1556 1485
rect 1630 1485 1636 1486
rect 1550 1480 1556 1481
rect 1571 1483 1580 1484
rect 1386 1478 1393 1479
rect 1571 1479 1572 1483
rect 1579 1479 1580 1483
rect 1630 1481 1631 1485
rect 1635 1481 1636 1485
rect 1710 1485 1716 1486
rect 1630 1480 1636 1481
rect 1651 1483 1660 1484
rect 1571 1478 1580 1479
rect 1651 1479 1652 1483
rect 1659 1479 1660 1483
rect 1710 1481 1711 1485
rect 1715 1481 1716 1485
rect 1710 1480 1716 1481
rect 1731 1485 1737 1486
rect 1731 1481 1732 1485
rect 1736 1481 1737 1485
rect 1731 1480 1737 1481
rect 1790 1485 1796 1486
rect 1790 1481 1791 1485
rect 1795 1481 1796 1485
rect 1870 1485 1876 1486
rect 1790 1480 1796 1481
rect 1811 1483 1820 1484
rect 1651 1478 1660 1479
rect 1811 1479 1812 1483
rect 1819 1479 1820 1483
rect 1870 1481 1871 1485
rect 1875 1481 1876 1485
rect 1950 1485 1956 1486
rect 1870 1480 1876 1481
rect 1891 1483 1900 1484
rect 1811 1478 1820 1479
rect 1891 1479 1892 1483
rect 1899 1479 1900 1483
rect 1950 1481 1951 1485
rect 1955 1481 1956 1485
rect 2030 1485 2036 1486
rect 1950 1480 1956 1481
rect 1971 1483 1980 1484
rect 1891 1478 1900 1479
rect 1971 1479 1972 1483
rect 1979 1479 1980 1483
rect 2030 1481 2031 1485
rect 2035 1481 2036 1485
rect 2118 1485 2124 1486
rect 2030 1480 2036 1481
rect 2051 1483 2060 1484
rect 1971 1478 1980 1479
rect 2051 1479 2052 1483
rect 2059 1479 2060 1483
rect 2118 1481 2119 1485
rect 2123 1481 2124 1485
rect 2118 1480 2124 1481
rect 2139 1485 2145 1486
rect 2139 1481 2140 1485
rect 2144 1481 2145 1485
rect 2139 1480 2145 1481
rect 2502 1484 2508 1485
rect 2502 1480 2503 1484
rect 2507 1480 2508 1484
rect 2502 1479 2508 1480
rect 2051 1478 2060 1479
rect 1286 1475 1292 1476
rect 1163 1474 1169 1475
rect 1326 1467 1332 1468
rect 110 1463 116 1464
rect 110 1459 111 1463
rect 115 1459 116 1463
rect 1286 1463 1292 1464
rect 110 1458 116 1459
rect 262 1460 268 1461
rect 262 1456 263 1460
rect 267 1456 268 1460
rect 262 1455 268 1456
rect 326 1460 332 1461
rect 326 1456 327 1460
rect 331 1456 332 1460
rect 326 1455 332 1456
rect 398 1460 404 1461
rect 398 1456 399 1460
rect 403 1456 404 1460
rect 398 1455 404 1456
rect 478 1460 484 1461
rect 478 1456 479 1460
rect 483 1456 484 1460
rect 478 1455 484 1456
rect 558 1460 564 1461
rect 558 1456 559 1460
rect 563 1456 564 1460
rect 558 1455 564 1456
rect 638 1460 644 1461
rect 638 1456 639 1460
rect 643 1456 644 1460
rect 638 1455 644 1456
rect 718 1460 724 1461
rect 718 1456 719 1460
rect 723 1456 724 1460
rect 718 1455 724 1456
rect 798 1460 804 1461
rect 798 1456 799 1460
rect 803 1456 804 1460
rect 798 1455 804 1456
rect 878 1460 884 1461
rect 878 1456 879 1460
rect 883 1456 884 1460
rect 878 1455 884 1456
rect 958 1460 964 1461
rect 958 1456 959 1460
rect 963 1456 964 1460
rect 958 1455 964 1456
rect 1038 1460 1044 1461
rect 1038 1456 1039 1460
rect 1043 1456 1044 1460
rect 1038 1455 1044 1456
rect 1126 1460 1132 1461
rect 1126 1456 1127 1460
rect 1131 1456 1132 1460
rect 1286 1459 1287 1463
rect 1291 1459 1292 1463
rect 1326 1463 1327 1467
rect 1331 1463 1332 1467
rect 2502 1467 2508 1468
rect 1326 1462 1332 1463
rect 1350 1464 1356 1465
rect 1350 1460 1351 1464
rect 1355 1460 1356 1464
rect 1350 1459 1356 1460
rect 1406 1464 1412 1465
rect 1406 1460 1407 1464
rect 1411 1460 1412 1464
rect 1406 1459 1412 1460
rect 1462 1464 1468 1465
rect 1462 1460 1463 1464
rect 1467 1460 1468 1464
rect 1462 1459 1468 1460
rect 1534 1464 1540 1465
rect 1534 1460 1535 1464
rect 1539 1460 1540 1464
rect 1534 1459 1540 1460
rect 1614 1464 1620 1465
rect 1614 1460 1615 1464
rect 1619 1460 1620 1464
rect 1614 1459 1620 1460
rect 1694 1464 1700 1465
rect 1694 1460 1695 1464
rect 1699 1460 1700 1464
rect 1694 1459 1700 1460
rect 1774 1464 1780 1465
rect 1774 1460 1775 1464
rect 1779 1460 1780 1464
rect 1774 1459 1780 1460
rect 1854 1464 1860 1465
rect 1854 1460 1855 1464
rect 1859 1460 1860 1464
rect 1854 1459 1860 1460
rect 1934 1464 1940 1465
rect 1934 1460 1935 1464
rect 1939 1460 1940 1464
rect 1934 1459 1940 1460
rect 2014 1464 2020 1465
rect 2014 1460 2015 1464
rect 2019 1460 2020 1464
rect 2014 1459 2020 1460
rect 2102 1464 2108 1465
rect 2102 1460 2103 1464
rect 2107 1460 2108 1464
rect 2502 1463 2503 1467
rect 2507 1463 2508 1467
rect 2502 1462 2508 1463
rect 2102 1459 2108 1460
rect 1286 1458 1292 1459
rect 1126 1455 1132 1456
rect 190 1444 196 1445
rect 110 1441 116 1442
rect 110 1437 111 1441
rect 115 1437 116 1441
rect 190 1440 191 1444
rect 195 1440 196 1444
rect 190 1439 196 1440
rect 254 1444 260 1445
rect 254 1440 255 1444
rect 259 1440 260 1444
rect 254 1439 260 1440
rect 326 1444 332 1445
rect 326 1440 327 1444
rect 331 1440 332 1444
rect 326 1439 332 1440
rect 406 1444 412 1445
rect 406 1440 407 1444
rect 411 1440 412 1444
rect 406 1439 412 1440
rect 502 1444 508 1445
rect 502 1440 503 1444
rect 507 1440 508 1444
rect 502 1439 508 1440
rect 606 1444 612 1445
rect 606 1440 607 1444
rect 611 1440 612 1444
rect 606 1439 612 1440
rect 710 1444 716 1445
rect 710 1440 711 1444
rect 715 1440 716 1444
rect 710 1439 716 1440
rect 814 1444 820 1445
rect 814 1440 815 1444
rect 819 1440 820 1444
rect 814 1439 820 1440
rect 918 1444 924 1445
rect 918 1440 919 1444
rect 923 1440 924 1444
rect 918 1439 924 1440
rect 1022 1444 1028 1445
rect 1022 1440 1023 1444
rect 1027 1440 1028 1444
rect 1022 1439 1028 1440
rect 1126 1444 1132 1445
rect 1126 1440 1127 1444
rect 1131 1440 1132 1444
rect 1126 1439 1132 1440
rect 1222 1444 1228 1445
rect 1222 1440 1223 1444
rect 1227 1440 1228 1444
rect 1358 1444 1364 1445
rect 1222 1439 1228 1440
rect 1286 1441 1292 1442
rect 110 1436 116 1437
rect 1286 1437 1287 1441
rect 1291 1437 1292 1441
rect 1286 1436 1292 1437
rect 1326 1441 1332 1442
rect 1326 1437 1327 1441
rect 1331 1437 1332 1441
rect 1358 1440 1359 1444
rect 1363 1440 1364 1444
rect 1358 1439 1364 1440
rect 1446 1444 1452 1445
rect 1446 1440 1447 1444
rect 1451 1440 1452 1444
rect 1446 1439 1452 1440
rect 1534 1444 1540 1445
rect 1534 1440 1535 1444
rect 1539 1440 1540 1444
rect 1534 1439 1540 1440
rect 1630 1444 1636 1445
rect 1630 1440 1631 1444
rect 1635 1440 1636 1444
rect 1630 1439 1636 1440
rect 1726 1444 1732 1445
rect 1726 1440 1727 1444
rect 1731 1440 1732 1444
rect 1726 1439 1732 1440
rect 1814 1444 1820 1445
rect 1814 1440 1815 1444
rect 1819 1440 1820 1444
rect 1814 1439 1820 1440
rect 1902 1444 1908 1445
rect 1902 1440 1903 1444
rect 1907 1440 1908 1444
rect 1902 1439 1908 1440
rect 1990 1444 1996 1445
rect 1990 1440 1991 1444
rect 1995 1440 1996 1444
rect 1990 1439 1996 1440
rect 2070 1444 2076 1445
rect 2070 1440 2071 1444
rect 2075 1440 2076 1444
rect 2070 1439 2076 1440
rect 2158 1444 2164 1445
rect 2158 1440 2159 1444
rect 2163 1440 2164 1444
rect 2158 1439 2164 1440
rect 2246 1444 2252 1445
rect 2246 1440 2247 1444
rect 2251 1440 2252 1444
rect 2246 1439 2252 1440
rect 2502 1441 2508 1442
rect 1326 1436 1332 1437
rect 2502 1437 2503 1441
rect 2507 1437 2508 1441
rect 2502 1436 2508 1437
rect 110 1424 116 1425
rect 1286 1424 1292 1425
rect 110 1420 111 1424
rect 115 1420 116 1424
rect 110 1419 116 1420
rect 206 1423 212 1424
rect 206 1419 207 1423
rect 211 1419 212 1423
rect 206 1418 212 1419
rect 214 1423 220 1424
rect 214 1419 215 1423
rect 219 1422 220 1423
rect 227 1423 233 1424
rect 227 1422 228 1423
rect 219 1420 228 1422
rect 219 1419 220 1420
rect 214 1418 220 1419
rect 227 1419 228 1420
rect 232 1419 233 1423
rect 227 1418 233 1419
rect 270 1423 276 1424
rect 270 1419 271 1423
rect 275 1419 276 1423
rect 291 1423 297 1424
rect 291 1422 292 1423
rect 270 1418 276 1419
rect 280 1420 292 1422
rect 280 1410 282 1420
rect 291 1419 292 1420
rect 296 1419 297 1423
rect 291 1418 297 1419
rect 342 1423 348 1424
rect 342 1419 343 1423
rect 347 1419 348 1423
rect 342 1418 348 1419
rect 350 1423 356 1424
rect 350 1419 351 1423
rect 355 1422 356 1423
rect 363 1423 369 1424
rect 363 1422 364 1423
rect 355 1420 364 1422
rect 355 1419 356 1420
rect 350 1418 356 1419
rect 363 1419 364 1420
rect 368 1419 369 1423
rect 363 1418 369 1419
rect 422 1423 428 1424
rect 422 1419 423 1423
rect 427 1419 428 1423
rect 443 1423 449 1424
rect 443 1422 444 1423
rect 422 1418 428 1419
rect 432 1420 444 1422
rect 432 1410 434 1420
rect 443 1419 444 1420
rect 448 1419 449 1423
rect 443 1418 449 1419
rect 518 1423 524 1424
rect 518 1419 519 1423
rect 523 1419 524 1423
rect 539 1423 545 1424
rect 539 1422 540 1423
rect 518 1418 524 1419
rect 528 1420 540 1422
rect 528 1410 530 1420
rect 539 1419 540 1420
rect 544 1419 545 1423
rect 539 1418 545 1419
rect 622 1423 628 1424
rect 622 1419 623 1423
rect 627 1419 628 1423
rect 622 1418 628 1419
rect 630 1423 636 1424
rect 630 1419 631 1423
rect 635 1422 636 1423
rect 643 1423 649 1424
rect 643 1422 644 1423
rect 635 1420 644 1422
rect 635 1419 636 1420
rect 630 1418 636 1419
rect 643 1419 644 1420
rect 648 1419 649 1423
rect 643 1418 649 1419
rect 726 1423 732 1424
rect 726 1419 727 1423
rect 731 1419 732 1423
rect 747 1423 753 1424
rect 747 1422 748 1423
rect 726 1418 732 1419
rect 736 1420 748 1422
rect 736 1410 738 1420
rect 747 1419 748 1420
rect 752 1419 753 1423
rect 747 1418 753 1419
rect 830 1423 836 1424
rect 830 1419 831 1423
rect 835 1419 836 1423
rect 830 1418 836 1419
rect 850 1423 857 1424
rect 850 1419 851 1423
rect 856 1419 857 1423
rect 850 1418 857 1419
rect 934 1423 940 1424
rect 934 1419 935 1423
rect 939 1419 940 1423
rect 934 1418 940 1419
rect 955 1423 961 1424
rect 955 1419 956 1423
rect 960 1422 961 1423
rect 1018 1423 1024 1424
rect 1018 1422 1019 1423
rect 960 1420 1019 1422
rect 960 1419 961 1420
rect 955 1418 961 1419
rect 1018 1419 1019 1420
rect 1023 1419 1024 1423
rect 1018 1418 1024 1419
rect 1038 1423 1044 1424
rect 1038 1419 1039 1423
rect 1043 1419 1044 1423
rect 1038 1418 1044 1419
rect 1059 1423 1065 1424
rect 1059 1419 1060 1423
rect 1064 1422 1065 1423
rect 1122 1423 1128 1424
rect 1122 1422 1123 1423
rect 1064 1420 1123 1422
rect 1064 1419 1065 1420
rect 1059 1418 1065 1419
rect 1122 1419 1123 1420
rect 1127 1419 1128 1423
rect 1122 1418 1128 1419
rect 1142 1423 1148 1424
rect 1142 1419 1143 1423
rect 1147 1419 1148 1423
rect 1142 1418 1148 1419
rect 1163 1423 1169 1424
rect 1163 1419 1164 1423
rect 1168 1422 1169 1423
rect 1218 1423 1224 1424
rect 1218 1422 1219 1423
rect 1168 1420 1219 1422
rect 1168 1419 1169 1420
rect 1163 1418 1169 1419
rect 1218 1419 1219 1420
rect 1223 1419 1224 1423
rect 1218 1418 1224 1419
rect 1238 1423 1244 1424
rect 1238 1419 1239 1423
rect 1243 1419 1244 1423
rect 1238 1418 1244 1419
rect 1246 1423 1252 1424
rect 1246 1419 1247 1423
rect 1251 1422 1252 1423
rect 1259 1423 1265 1424
rect 1259 1422 1260 1423
rect 1251 1420 1260 1422
rect 1251 1419 1252 1420
rect 1246 1418 1252 1419
rect 1259 1419 1260 1420
rect 1264 1419 1265 1423
rect 1286 1420 1287 1424
rect 1291 1420 1292 1424
rect 1286 1419 1292 1420
rect 1326 1424 1332 1425
rect 2502 1424 2508 1425
rect 1326 1420 1327 1424
rect 1331 1420 1332 1424
rect 1326 1419 1332 1420
rect 1374 1423 1380 1424
rect 1374 1419 1375 1423
rect 1379 1419 1380 1423
rect 1259 1418 1265 1419
rect 1374 1418 1380 1419
rect 1395 1423 1401 1424
rect 1395 1419 1396 1423
rect 1400 1422 1401 1423
rect 1442 1423 1448 1424
rect 1442 1422 1443 1423
rect 1400 1420 1443 1422
rect 1400 1419 1401 1420
rect 1395 1418 1401 1419
rect 1442 1419 1443 1420
rect 1447 1419 1448 1423
rect 1442 1418 1448 1419
rect 1462 1423 1468 1424
rect 1462 1419 1463 1423
rect 1467 1419 1468 1423
rect 1462 1418 1468 1419
rect 1483 1423 1489 1424
rect 1483 1419 1484 1423
rect 1488 1422 1489 1423
rect 1530 1423 1536 1424
rect 1530 1422 1531 1423
rect 1488 1420 1531 1422
rect 1488 1419 1489 1420
rect 1483 1418 1489 1419
rect 1530 1419 1531 1420
rect 1535 1419 1536 1423
rect 1530 1418 1536 1419
rect 1550 1423 1556 1424
rect 1550 1419 1551 1423
rect 1555 1419 1556 1423
rect 1550 1418 1556 1419
rect 1566 1423 1577 1424
rect 1566 1419 1567 1423
rect 1571 1419 1572 1423
rect 1576 1419 1577 1423
rect 1566 1418 1577 1419
rect 1646 1423 1652 1424
rect 1646 1419 1647 1423
rect 1651 1419 1652 1423
rect 1667 1423 1673 1424
rect 1667 1422 1668 1423
rect 1646 1418 1652 1419
rect 1656 1420 1668 1422
rect 1656 1414 1658 1420
rect 1667 1419 1668 1420
rect 1672 1419 1673 1423
rect 1667 1418 1673 1419
rect 1742 1423 1748 1424
rect 1742 1419 1743 1423
rect 1747 1419 1748 1423
rect 1763 1423 1769 1424
rect 1763 1422 1764 1423
rect 1742 1418 1748 1419
rect 1752 1420 1764 1422
rect 1356 1412 1658 1414
rect 1150 1411 1156 1412
rect 1150 1410 1151 1411
rect 188 1408 282 1410
rect 324 1408 434 1410
rect 436 1408 530 1410
rect 604 1408 738 1410
rect 916 1408 1151 1410
rect 188 1406 190 1408
rect 324 1406 326 1408
rect 436 1406 438 1408
rect 604 1406 606 1408
rect 916 1406 918 1408
rect 1150 1407 1151 1408
rect 1155 1407 1156 1411
rect 1150 1406 1156 1407
rect 1356 1406 1358 1412
rect 1752 1410 1754 1420
rect 1763 1419 1764 1420
rect 1768 1419 1769 1423
rect 1763 1418 1769 1419
rect 1830 1423 1836 1424
rect 1830 1419 1831 1423
rect 1835 1419 1836 1423
rect 1830 1418 1836 1419
rect 1851 1423 1857 1424
rect 1851 1419 1852 1423
rect 1856 1422 1857 1423
rect 1898 1423 1904 1424
rect 1898 1422 1899 1423
rect 1856 1420 1899 1422
rect 1856 1419 1857 1420
rect 1851 1418 1857 1419
rect 1898 1419 1899 1420
rect 1903 1419 1904 1423
rect 1898 1418 1904 1419
rect 1918 1423 1924 1424
rect 1918 1419 1919 1423
rect 1923 1419 1924 1423
rect 1918 1418 1924 1419
rect 1939 1423 1945 1424
rect 1939 1419 1940 1423
rect 1944 1422 1945 1423
rect 1986 1423 1992 1424
rect 1986 1422 1987 1423
rect 1944 1420 1987 1422
rect 1944 1419 1945 1420
rect 1939 1418 1945 1419
rect 1986 1419 1987 1420
rect 1991 1419 1992 1423
rect 1986 1418 1992 1419
rect 2006 1423 2012 1424
rect 2006 1419 2007 1423
rect 2011 1419 2012 1423
rect 2006 1418 2012 1419
rect 2027 1423 2033 1424
rect 2027 1419 2028 1423
rect 2032 1422 2033 1423
rect 2066 1423 2072 1424
rect 2066 1422 2067 1423
rect 2032 1420 2067 1422
rect 2032 1419 2033 1420
rect 2027 1418 2033 1419
rect 2066 1419 2067 1420
rect 2071 1419 2072 1423
rect 2066 1418 2072 1419
rect 2086 1423 2092 1424
rect 2086 1419 2087 1423
rect 2091 1419 2092 1423
rect 2086 1418 2092 1419
rect 2107 1423 2113 1424
rect 2107 1419 2108 1423
rect 2112 1422 2113 1423
rect 2154 1423 2160 1424
rect 2154 1422 2155 1423
rect 2112 1420 2155 1422
rect 2112 1419 2113 1420
rect 2107 1418 2113 1419
rect 2154 1419 2155 1420
rect 2159 1419 2160 1423
rect 2154 1418 2160 1419
rect 2174 1423 2180 1424
rect 2174 1419 2175 1423
rect 2179 1419 2180 1423
rect 2174 1418 2180 1419
rect 2195 1423 2201 1424
rect 2195 1419 2196 1423
rect 2200 1422 2201 1423
rect 2238 1423 2244 1424
rect 2238 1422 2239 1423
rect 2200 1420 2239 1422
rect 2200 1419 2201 1420
rect 2195 1418 2201 1419
rect 2238 1419 2239 1420
rect 2243 1419 2244 1423
rect 2238 1418 2244 1419
rect 2262 1423 2268 1424
rect 2262 1419 2263 1423
rect 2267 1419 2268 1423
rect 2262 1418 2268 1419
rect 2283 1423 2289 1424
rect 2283 1419 2284 1423
rect 2288 1419 2289 1423
rect 2502 1420 2503 1424
rect 2507 1420 2508 1424
rect 2502 1419 2508 1420
rect 2283 1418 2289 1419
rect 1994 1415 2000 1416
rect 1994 1411 1995 1415
rect 1999 1414 2000 1415
rect 2285 1414 2287 1418
rect 1999 1412 2287 1414
rect 1999 1411 2000 1412
rect 1994 1410 2000 1411
rect 1628 1408 1754 1410
rect 1628 1406 1630 1408
rect 187 1405 193 1406
rect 187 1401 188 1405
rect 192 1401 193 1405
rect 323 1405 329 1406
rect 187 1400 193 1401
rect 251 1403 257 1404
rect 251 1399 252 1403
rect 256 1402 257 1403
rect 286 1403 292 1404
rect 286 1402 287 1403
rect 256 1400 287 1402
rect 256 1399 257 1400
rect 251 1398 257 1399
rect 286 1399 287 1400
rect 291 1399 292 1403
rect 323 1401 324 1405
rect 328 1401 329 1405
rect 323 1400 329 1401
rect 403 1405 438 1406
rect 403 1401 404 1405
rect 408 1404 438 1405
rect 603 1405 609 1406
rect 408 1401 409 1404
rect 403 1400 409 1401
rect 499 1403 505 1404
rect 286 1398 292 1399
rect 499 1399 500 1403
rect 504 1402 505 1403
rect 510 1403 516 1404
rect 510 1402 511 1403
rect 504 1400 511 1402
rect 504 1399 505 1400
rect 499 1398 505 1399
rect 510 1399 511 1400
rect 515 1399 516 1403
rect 603 1401 604 1405
rect 608 1401 609 1405
rect 915 1405 921 1406
rect 603 1400 609 1401
rect 686 1403 692 1404
rect 510 1398 516 1399
rect 686 1399 687 1403
rect 691 1402 692 1403
rect 707 1403 713 1404
rect 707 1402 708 1403
rect 691 1400 708 1402
rect 691 1399 692 1400
rect 686 1398 692 1399
rect 707 1399 708 1400
rect 712 1399 713 1403
rect 707 1398 713 1399
rect 811 1403 817 1404
rect 811 1399 812 1403
rect 816 1402 817 1403
rect 858 1403 864 1404
rect 858 1402 859 1403
rect 816 1400 859 1402
rect 816 1399 817 1400
rect 811 1398 817 1399
rect 858 1399 859 1400
rect 863 1399 864 1403
rect 915 1401 916 1405
rect 920 1401 921 1405
rect 1355 1405 1361 1406
rect 915 1400 921 1401
rect 1018 1403 1025 1404
rect 858 1398 864 1399
rect 1018 1399 1019 1403
rect 1024 1399 1025 1403
rect 1018 1398 1025 1399
rect 1122 1403 1129 1404
rect 1122 1399 1123 1403
rect 1128 1399 1129 1403
rect 1122 1398 1129 1399
rect 1218 1403 1225 1404
rect 1218 1399 1219 1403
rect 1224 1399 1225 1403
rect 1355 1401 1356 1405
rect 1360 1401 1361 1405
rect 1627 1405 1633 1406
rect 1355 1400 1361 1401
rect 1442 1403 1449 1404
rect 1218 1398 1225 1399
rect 1442 1399 1443 1403
rect 1448 1399 1449 1403
rect 1442 1398 1449 1399
rect 1530 1403 1537 1404
rect 1530 1399 1531 1403
rect 1536 1399 1537 1403
rect 1627 1401 1628 1405
rect 1632 1401 1633 1405
rect 1627 1400 1633 1401
rect 1723 1403 1729 1404
rect 1530 1398 1537 1399
rect 1723 1399 1724 1403
rect 1728 1402 1729 1403
rect 1754 1403 1760 1404
rect 1754 1402 1755 1403
rect 1728 1400 1755 1402
rect 1728 1399 1729 1400
rect 1723 1398 1729 1399
rect 1754 1399 1755 1400
rect 1759 1399 1760 1403
rect 1754 1398 1760 1399
rect 1811 1403 1817 1404
rect 1811 1399 1812 1403
rect 1816 1402 1817 1403
rect 1822 1403 1828 1404
rect 1822 1402 1823 1403
rect 1816 1400 1823 1402
rect 1816 1399 1817 1400
rect 1811 1398 1817 1399
rect 1822 1399 1823 1400
rect 1827 1399 1828 1403
rect 1822 1398 1828 1399
rect 1898 1403 1905 1404
rect 1898 1399 1899 1403
rect 1904 1399 1905 1403
rect 1898 1398 1905 1399
rect 1986 1403 1993 1404
rect 1986 1399 1987 1403
rect 1992 1399 1993 1403
rect 1986 1398 1993 1399
rect 2066 1403 2073 1404
rect 2066 1399 2067 1403
rect 2072 1399 2073 1403
rect 2066 1398 2073 1399
rect 2154 1403 2161 1404
rect 2154 1399 2155 1403
rect 2160 1399 2161 1403
rect 2154 1398 2161 1399
rect 2238 1403 2249 1404
rect 2238 1399 2239 1403
rect 2243 1399 2244 1403
rect 2248 1399 2249 1403
rect 2238 1398 2249 1399
rect 214 1395 220 1396
rect 214 1394 215 1395
rect 132 1392 215 1394
rect 132 1390 134 1392
rect 214 1391 215 1392
rect 219 1391 220 1395
rect 350 1395 356 1396
rect 350 1394 351 1395
rect 214 1390 220 1391
rect 276 1392 351 1394
rect 276 1390 278 1392
rect 350 1391 351 1392
rect 355 1391 356 1395
rect 350 1390 356 1391
rect 1547 1391 1553 1392
rect 131 1389 137 1390
rect 131 1385 132 1389
rect 136 1385 137 1389
rect 275 1389 281 1390
rect 131 1384 137 1385
rect 174 1387 180 1388
rect 174 1383 175 1387
rect 179 1386 180 1387
rect 203 1387 209 1388
rect 203 1386 204 1387
rect 179 1384 204 1386
rect 179 1383 180 1384
rect 174 1382 180 1383
rect 203 1383 204 1384
rect 208 1383 209 1387
rect 275 1385 276 1389
rect 280 1385 281 1389
rect 275 1384 281 1385
rect 327 1387 333 1388
rect 203 1382 209 1383
rect 327 1383 328 1387
rect 332 1386 333 1387
rect 339 1387 345 1388
rect 339 1386 340 1387
rect 332 1384 340 1386
rect 332 1383 333 1384
rect 327 1382 333 1383
rect 339 1383 340 1384
rect 344 1383 345 1387
rect 339 1382 345 1383
rect 382 1387 388 1388
rect 382 1383 383 1387
rect 387 1386 388 1387
rect 411 1387 417 1388
rect 411 1386 412 1387
rect 387 1384 412 1386
rect 387 1383 388 1384
rect 382 1382 388 1383
rect 411 1383 412 1384
rect 416 1383 417 1387
rect 411 1382 417 1383
rect 462 1387 468 1388
rect 462 1383 463 1387
rect 467 1386 468 1387
rect 483 1387 489 1388
rect 483 1386 484 1387
rect 467 1384 484 1386
rect 467 1383 468 1384
rect 462 1382 468 1383
rect 483 1383 484 1384
rect 488 1383 489 1387
rect 483 1382 489 1383
rect 526 1387 532 1388
rect 526 1383 527 1387
rect 531 1386 532 1387
rect 563 1387 569 1388
rect 563 1386 564 1387
rect 531 1384 564 1386
rect 531 1383 532 1384
rect 526 1382 532 1383
rect 563 1383 564 1384
rect 568 1383 569 1387
rect 563 1382 569 1383
rect 606 1387 612 1388
rect 606 1383 607 1387
rect 611 1386 612 1387
rect 643 1387 649 1388
rect 643 1386 644 1387
rect 611 1384 644 1386
rect 611 1383 612 1384
rect 606 1382 612 1383
rect 643 1383 644 1384
rect 648 1383 649 1387
rect 643 1382 649 1383
rect 654 1387 660 1388
rect 654 1383 655 1387
rect 659 1386 660 1387
rect 731 1387 737 1388
rect 731 1386 732 1387
rect 659 1384 732 1386
rect 659 1383 660 1384
rect 654 1382 660 1383
rect 731 1383 732 1384
rect 736 1383 737 1387
rect 731 1382 737 1383
rect 774 1387 780 1388
rect 774 1383 775 1387
rect 779 1386 780 1387
rect 819 1387 825 1388
rect 819 1386 820 1387
rect 779 1384 820 1386
rect 779 1383 780 1384
rect 774 1382 780 1383
rect 819 1383 820 1384
rect 824 1383 825 1387
rect 819 1382 825 1383
rect 907 1387 913 1388
rect 907 1383 908 1387
rect 912 1386 913 1387
rect 995 1387 1001 1388
rect 912 1384 990 1386
rect 912 1383 913 1384
rect 907 1382 913 1383
rect 988 1374 990 1384
rect 995 1383 996 1387
rect 1000 1386 1001 1387
rect 1083 1387 1089 1388
rect 1000 1384 1078 1386
rect 1000 1383 1001 1384
rect 995 1382 1001 1383
rect 1076 1374 1078 1384
rect 1083 1383 1084 1387
rect 1088 1386 1089 1387
rect 1179 1387 1185 1388
rect 1088 1384 1161 1386
rect 1088 1383 1089 1384
rect 1083 1382 1089 1383
rect 1159 1374 1161 1384
rect 1179 1383 1180 1387
rect 1184 1386 1185 1387
rect 1246 1387 1252 1388
rect 1246 1386 1247 1387
rect 1184 1384 1247 1386
rect 1184 1383 1185 1384
rect 1179 1382 1185 1383
rect 1246 1383 1247 1384
rect 1251 1383 1252 1387
rect 1547 1387 1548 1391
rect 1552 1390 1553 1391
rect 1590 1391 1596 1392
rect 1552 1388 1586 1390
rect 1552 1387 1553 1388
rect 1547 1386 1553 1387
rect 1246 1382 1252 1383
rect 1584 1378 1586 1388
rect 1590 1387 1591 1391
rect 1595 1390 1596 1391
rect 1627 1391 1633 1392
rect 1627 1390 1628 1391
rect 1595 1388 1628 1390
rect 1595 1387 1596 1388
rect 1590 1386 1596 1387
rect 1627 1387 1628 1388
rect 1632 1387 1633 1391
rect 1627 1386 1633 1387
rect 1670 1391 1676 1392
rect 1670 1387 1671 1391
rect 1675 1390 1676 1391
rect 1715 1391 1721 1392
rect 1715 1390 1716 1391
rect 1675 1388 1716 1390
rect 1675 1387 1676 1388
rect 1670 1386 1676 1387
rect 1715 1387 1716 1388
rect 1720 1387 1721 1391
rect 1715 1386 1721 1387
rect 1811 1391 1817 1392
rect 1811 1387 1812 1391
rect 1816 1390 1817 1391
rect 1899 1391 1905 1392
rect 1816 1388 1890 1390
rect 1816 1387 1817 1388
rect 1811 1386 1817 1387
rect 1888 1378 1890 1388
rect 1899 1387 1900 1391
rect 1904 1390 1905 1391
rect 1930 1391 1936 1392
rect 1930 1390 1931 1391
rect 1904 1388 1931 1390
rect 1904 1387 1905 1388
rect 1899 1386 1905 1387
rect 1930 1387 1931 1388
rect 1935 1387 1936 1391
rect 1930 1386 1936 1387
rect 1987 1391 1996 1392
rect 1987 1387 1988 1391
rect 1995 1387 1996 1391
rect 1987 1386 1996 1387
rect 2030 1391 2036 1392
rect 2030 1387 2031 1391
rect 2035 1390 2036 1391
rect 2075 1391 2081 1392
rect 2075 1390 2076 1391
rect 2035 1388 2076 1390
rect 2035 1387 2036 1388
rect 2030 1386 2036 1387
rect 2075 1387 2076 1388
rect 2080 1387 2081 1391
rect 2075 1386 2081 1387
rect 2118 1391 2124 1392
rect 2118 1387 2119 1391
rect 2123 1390 2124 1391
rect 2155 1391 2161 1392
rect 2155 1390 2156 1391
rect 2123 1388 2156 1390
rect 2123 1387 2124 1388
rect 2118 1386 2124 1387
rect 2155 1387 2156 1388
rect 2160 1387 2161 1391
rect 2155 1386 2161 1387
rect 2214 1391 2220 1392
rect 2214 1387 2215 1391
rect 2219 1390 2220 1391
rect 2227 1391 2233 1392
rect 2227 1390 2228 1391
rect 2219 1388 2228 1390
rect 2219 1387 2220 1388
rect 2214 1386 2220 1387
rect 2227 1387 2228 1388
rect 2232 1387 2233 1391
rect 2227 1386 2233 1387
rect 2270 1391 2276 1392
rect 2270 1387 2271 1391
rect 2275 1390 2276 1391
rect 2299 1391 2305 1392
rect 2299 1390 2300 1391
rect 2275 1388 2300 1390
rect 2275 1387 2276 1388
rect 2270 1386 2276 1387
rect 2299 1387 2300 1388
rect 2304 1387 2305 1391
rect 2299 1386 2305 1387
rect 2379 1391 2385 1392
rect 2379 1387 2380 1391
rect 2384 1390 2385 1391
rect 2414 1391 2420 1392
rect 2414 1390 2415 1391
rect 2384 1388 2415 1390
rect 2384 1387 2385 1388
rect 2379 1386 2385 1387
rect 2414 1387 2415 1388
rect 2419 1387 2420 1391
rect 2414 1386 2420 1387
rect 2422 1391 2428 1392
rect 2422 1387 2423 1391
rect 2427 1390 2428 1391
rect 2435 1391 2441 1392
rect 2435 1390 2436 1391
rect 2427 1388 2436 1390
rect 2427 1387 2428 1388
rect 2422 1386 2428 1387
rect 2435 1387 2436 1388
rect 2440 1387 2441 1391
rect 2435 1386 2441 1387
rect 1584 1376 1854 1378
rect 1888 1376 1942 1378
rect 1852 1374 1854 1376
rect 1940 1374 1942 1376
rect 988 1372 1038 1374
rect 1076 1372 1126 1374
rect 1159 1372 1222 1374
rect 1566 1373 1572 1374
rect 1036 1370 1038 1372
rect 1124 1370 1126 1372
rect 1220 1370 1222 1372
rect 1326 1372 1332 1373
rect 150 1369 156 1370
rect 110 1368 116 1369
rect 110 1364 111 1368
rect 115 1364 116 1368
rect 150 1365 151 1369
rect 155 1365 156 1369
rect 222 1369 228 1370
rect 150 1364 156 1365
rect 171 1367 180 1368
rect 110 1363 116 1364
rect 171 1363 172 1367
rect 179 1363 180 1367
rect 222 1365 223 1369
rect 227 1365 228 1369
rect 294 1369 300 1370
rect 222 1364 228 1365
rect 243 1367 252 1368
rect 171 1362 180 1363
rect 243 1363 244 1367
rect 251 1363 252 1367
rect 294 1365 295 1369
rect 299 1365 300 1369
rect 358 1369 364 1370
rect 294 1364 300 1365
rect 315 1367 321 1368
rect 243 1362 252 1363
rect 315 1363 316 1367
rect 320 1366 321 1367
rect 327 1367 333 1368
rect 327 1366 328 1367
rect 320 1364 328 1366
rect 320 1363 321 1364
rect 315 1362 321 1363
rect 327 1363 328 1364
rect 332 1363 333 1367
rect 358 1365 359 1369
rect 363 1365 364 1369
rect 430 1369 436 1370
rect 358 1364 364 1365
rect 379 1367 388 1368
rect 327 1362 333 1363
rect 379 1363 380 1367
rect 387 1363 388 1367
rect 430 1365 431 1369
rect 435 1365 436 1369
rect 502 1369 508 1370
rect 430 1364 436 1365
rect 451 1367 457 1368
rect 379 1362 388 1363
rect 451 1363 452 1367
rect 456 1366 457 1367
rect 462 1367 468 1368
rect 462 1366 463 1367
rect 456 1364 463 1366
rect 456 1363 457 1364
rect 451 1362 457 1363
rect 462 1363 463 1364
rect 467 1363 468 1367
rect 502 1365 503 1369
rect 507 1365 508 1369
rect 582 1369 588 1370
rect 502 1364 508 1365
rect 523 1367 532 1368
rect 462 1362 468 1363
rect 523 1363 524 1367
rect 531 1363 532 1367
rect 582 1365 583 1369
rect 587 1365 588 1369
rect 662 1369 668 1370
rect 582 1364 588 1365
rect 603 1367 612 1368
rect 523 1362 532 1363
rect 603 1363 604 1367
rect 611 1363 612 1367
rect 662 1365 663 1369
rect 667 1365 668 1369
rect 750 1369 756 1370
rect 662 1364 668 1365
rect 683 1367 692 1368
rect 603 1362 612 1363
rect 683 1363 684 1367
rect 691 1363 692 1367
rect 750 1365 751 1369
rect 755 1365 756 1369
rect 838 1369 844 1370
rect 750 1364 756 1365
rect 771 1367 780 1368
rect 683 1362 692 1363
rect 771 1363 772 1367
rect 779 1363 780 1367
rect 838 1365 839 1369
rect 843 1365 844 1369
rect 926 1369 932 1370
rect 838 1364 844 1365
rect 858 1367 865 1368
rect 771 1362 780 1363
rect 858 1363 859 1367
rect 864 1363 865 1367
rect 926 1365 927 1369
rect 931 1365 932 1369
rect 1014 1369 1020 1370
rect 926 1364 932 1365
rect 947 1367 953 1368
rect 858 1362 865 1363
rect 947 1363 948 1367
rect 952 1366 953 1367
rect 966 1367 972 1368
rect 966 1366 967 1367
rect 952 1364 967 1366
rect 952 1363 953 1364
rect 947 1362 953 1363
rect 966 1363 967 1364
rect 971 1363 972 1367
rect 1014 1365 1015 1369
rect 1019 1365 1020 1369
rect 1014 1364 1020 1365
rect 1035 1369 1041 1370
rect 1035 1365 1036 1369
rect 1040 1365 1041 1369
rect 1035 1364 1041 1365
rect 1102 1369 1108 1370
rect 1102 1365 1103 1369
rect 1107 1365 1108 1369
rect 1102 1364 1108 1365
rect 1123 1369 1129 1370
rect 1123 1365 1124 1369
rect 1128 1365 1129 1369
rect 1123 1364 1129 1365
rect 1198 1369 1204 1370
rect 1198 1365 1199 1369
rect 1203 1365 1204 1369
rect 1198 1364 1204 1365
rect 1219 1369 1225 1370
rect 1219 1365 1220 1369
rect 1224 1365 1225 1369
rect 1219 1364 1225 1365
rect 1286 1368 1292 1369
rect 1286 1364 1287 1368
rect 1291 1364 1292 1368
rect 1326 1368 1327 1372
rect 1331 1368 1332 1372
rect 1566 1369 1567 1373
rect 1571 1369 1572 1373
rect 1646 1373 1652 1374
rect 1566 1368 1572 1369
rect 1587 1371 1596 1372
rect 1326 1367 1332 1368
rect 1587 1367 1588 1371
rect 1595 1367 1596 1371
rect 1646 1369 1647 1373
rect 1651 1369 1652 1373
rect 1734 1373 1740 1374
rect 1646 1368 1652 1369
rect 1667 1371 1676 1372
rect 1587 1366 1596 1367
rect 1667 1367 1668 1371
rect 1675 1367 1676 1371
rect 1734 1369 1735 1373
rect 1739 1369 1740 1373
rect 1830 1373 1836 1374
rect 1734 1368 1740 1369
rect 1754 1371 1761 1372
rect 1667 1366 1676 1367
rect 1754 1367 1755 1371
rect 1760 1367 1761 1371
rect 1830 1369 1831 1373
rect 1835 1369 1836 1373
rect 1830 1368 1836 1369
rect 1851 1373 1857 1374
rect 1851 1369 1852 1373
rect 1856 1369 1857 1373
rect 1851 1368 1857 1369
rect 1918 1373 1924 1374
rect 1918 1369 1919 1373
rect 1923 1369 1924 1373
rect 1918 1368 1924 1369
rect 1939 1373 1945 1374
rect 1939 1369 1940 1373
rect 1944 1369 1945 1373
rect 1939 1368 1945 1369
rect 2006 1373 2012 1374
rect 2006 1369 2007 1373
rect 2011 1369 2012 1373
rect 2094 1373 2100 1374
rect 2006 1368 2012 1369
rect 2027 1371 2036 1372
rect 1754 1366 1761 1367
rect 2027 1367 2028 1371
rect 2035 1367 2036 1371
rect 2094 1369 2095 1373
rect 2099 1369 2100 1373
rect 2174 1373 2180 1374
rect 2094 1368 2100 1369
rect 2115 1371 2124 1372
rect 2027 1366 2036 1367
rect 2115 1367 2116 1371
rect 2123 1367 2124 1371
rect 2174 1369 2175 1373
rect 2179 1369 2180 1373
rect 2246 1373 2252 1374
rect 2174 1368 2180 1369
rect 2195 1371 2201 1372
rect 2115 1366 2124 1367
rect 2195 1367 2196 1371
rect 2200 1370 2201 1371
rect 2214 1371 2220 1372
rect 2214 1370 2215 1371
rect 2200 1368 2215 1370
rect 2200 1367 2201 1368
rect 2195 1366 2201 1367
rect 2214 1367 2215 1368
rect 2219 1367 2220 1371
rect 2246 1369 2247 1373
rect 2251 1369 2252 1373
rect 2318 1373 2324 1374
rect 2246 1368 2252 1369
rect 2267 1371 2276 1372
rect 2214 1366 2220 1367
rect 2267 1367 2268 1371
rect 2275 1367 2276 1371
rect 2318 1369 2319 1373
rect 2323 1369 2324 1373
rect 2398 1373 2404 1374
rect 2318 1368 2324 1369
rect 2326 1371 2332 1372
rect 2267 1366 2276 1367
rect 2326 1367 2327 1371
rect 2331 1370 2332 1371
rect 2339 1371 2345 1372
rect 2339 1370 2340 1371
rect 2331 1368 2340 1370
rect 2331 1367 2332 1368
rect 2326 1366 2332 1367
rect 2339 1367 2340 1368
rect 2344 1367 2345 1371
rect 2398 1369 2399 1373
rect 2403 1369 2404 1373
rect 2454 1373 2460 1374
rect 2398 1368 2404 1369
rect 2419 1371 2428 1372
rect 2339 1366 2345 1367
rect 2419 1367 2420 1371
rect 2427 1367 2428 1371
rect 2454 1369 2455 1373
rect 2459 1369 2460 1373
rect 2502 1372 2508 1373
rect 2454 1368 2460 1369
rect 2462 1371 2468 1372
rect 2419 1366 2428 1367
rect 2462 1367 2463 1371
rect 2467 1370 2468 1371
rect 2475 1371 2481 1372
rect 2475 1370 2476 1371
rect 2467 1368 2476 1370
rect 2467 1367 2468 1368
rect 2462 1366 2468 1367
rect 2475 1367 2476 1368
rect 2480 1367 2481 1371
rect 2502 1368 2503 1372
rect 2507 1368 2508 1372
rect 2502 1367 2508 1368
rect 2475 1366 2481 1367
rect 1286 1363 1292 1364
rect 966 1362 972 1363
rect 1326 1355 1332 1356
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 1286 1351 1292 1352
rect 110 1346 116 1347
rect 134 1348 140 1349
rect 134 1344 135 1348
rect 139 1344 140 1348
rect 134 1343 140 1344
rect 206 1348 212 1349
rect 206 1344 207 1348
rect 211 1344 212 1348
rect 206 1343 212 1344
rect 278 1348 284 1349
rect 278 1344 279 1348
rect 283 1344 284 1348
rect 278 1343 284 1344
rect 342 1348 348 1349
rect 342 1344 343 1348
rect 347 1344 348 1348
rect 342 1343 348 1344
rect 414 1348 420 1349
rect 414 1344 415 1348
rect 419 1344 420 1348
rect 414 1343 420 1344
rect 486 1348 492 1349
rect 486 1344 487 1348
rect 491 1344 492 1348
rect 486 1343 492 1344
rect 566 1348 572 1349
rect 566 1344 567 1348
rect 571 1344 572 1348
rect 566 1343 572 1344
rect 646 1348 652 1349
rect 646 1344 647 1348
rect 651 1344 652 1348
rect 646 1343 652 1344
rect 734 1348 740 1349
rect 734 1344 735 1348
rect 739 1344 740 1348
rect 734 1343 740 1344
rect 822 1348 828 1349
rect 822 1344 823 1348
rect 827 1344 828 1348
rect 822 1343 828 1344
rect 910 1348 916 1349
rect 910 1344 911 1348
rect 915 1344 916 1348
rect 910 1343 916 1344
rect 998 1348 1004 1349
rect 998 1344 999 1348
rect 1003 1344 1004 1348
rect 998 1343 1004 1344
rect 1086 1348 1092 1349
rect 1086 1344 1087 1348
rect 1091 1344 1092 1348
rect 1086 1343 1092 1344
rect 1182 1348 1188 1349
rect 1182 1344 1183 1348
rect 1187 1344 1188 1348
rect 1286 1347 1287 1351
rect 1291 1347 1292 1351
rect 1326 1351 1327 1355
rect 1331 1351 1332 1355
rect 2502 1355 2508 1356
rect 1326 1350 1332 1351
rect 1550 1352 1556 1353
rect 1550 1348 1551 1352
rect 1555 1348 1556 1352
rect 1550 1347 1556 1348
rect 1630 1352 1636 1353
rect 1630 1348 1631 1352
rect 1635 1348 1636 1352
rect 1630 1347 1636 1348
rect 1718 1352 1724 1353
rect 1718 1348 1719 1352
rect 1723 1348 1724 1352
rect 1718 1347 1724 1348
rect 1814 1352 1820 1353
rect 1814 1348 1815 1352
rect 1819 1348 1820 1352
rect 1814 1347 1820 1348
rect 1902 1352 1908 1353
rect 1902 1348 1903 1352
rect 1907 1348 1908 1352
rect 1902 1347 1908 1348
rect 1990 1352 1996 1353
rect 1990 1348 1991 1352
rect 1995 1348 1996 1352
rect 1990 1347 1996 1348
rect 2078 1352 2084 1353
rect 2078 1348 2079 1352
rect 2083 1348 2084 1352
rect 2078 1347 2084 1348
rect 2158 1352 2164 1353
rect 2158 1348 2159 1352
rect 2163 1348 2164 1352
rect 2158 1347 2164 1348
rect 2230 1352 2236 1353
rect 2230 1348 2231 1352
rect 2235 1348 2236 1352
rect 2230 1347 2236 1348
rect 2302 1352 2308 1353
rect 2302 1348 2303 1352
rect 2307 1348 2308 1352
rect 2302 1347 2308 1348
rect 2382 1352 2388 1353
rect 2382 1348 2383 1352
rect 2387 1348 2388 1352
rect 2382 1347 2388 1348
rect 2438 1352 2444 1353
rect 2438 1348 2439 1352
rect 2443 1348 2444 1352
rect 2502 1351 2503 1355
rect 2507 1351 2508 1355
rect 2502 1350 2508 1351
rect 2438 1347 2444 1348
rect 1286 1346 1292 1347
rect 1182 1343 1188 1344
rect 1582 1340 1588 1341
rect 1326 1337 1332 1338
rect 1326 1333 1327 1337
rect 1331 1333 1332 1337
rect 1582 1336 1583 1340
rect 1587 1336 1588 1340
rect 1582 1335 1588 1336
rect 1646 1340 1652 1341
rect 1646 1336 1647 1340
rect 1651 1336 1652 1340
rect 1646 1335 1652 1336
rect 1726 1340 1732 1341
rect 1726 1336 1727 1340
rect 1731 1336 1732 1340
rect 1726 1335 1732 1336
rect 1806 1340 1812 1341
rect 1806 1336 1807 1340
rect 1811 1336 1812 1340
rect 1806 1335 1812 1336
rect 1894 1340 1900 1341
rect 1894 1336 1895 1340
rect 1899 1336 1900 1340
rect 1894 1335 1900 1336
rect 1982 1340 1988 1341
rect 1982 1336 1983 1340
rect 1987 1336 1988 1340
rect 1982 1335 1988 1336
rect 2062 1340 2068 1341
rect 2062 1336 2063 1340
rect 2067 1336 2068 1340
rect 2062 1335 2068 1336
rect 2142 1340 2148 1341
rect 2142 1336 2143 1340
rect 2147 1336 2148 1340
rect 2142 1335 2148 1336
rect 2222 1340 2228 1341
rect 2222 1336 2223 1340
rect 2227 1336 2228 1340
rect 2222 1335 2228 1336
rect 2302 1340 2308 1341
rect 2302 1336 2303 1340
rect 2307 1336 2308 1340
rect 2302 1335 2308 1336
rect 2382 1340 2388 1341
rect 2382 1336 2383 1340
rect 2387 1336 2388 1340
rect 2382 1335 2388 1336
rect 2438 1340 2444 1341
rect 2438 1336 2439 1340
rect 2443 1336 2444 1340
rect 2438 1335 2444 1336
rect 2502 1337 2508 1338
rect 1326 1332 1332 1333
rect 2502 1333 2503 1337
rect 2507 1333 2508 1337
rect 2502 1332 2508 1333
rect 134 1320 140 1321
rect 110 1317 116 1318
rect 110 1313 111 1317
rect 115 1313 116 1317
rect 134 1316 135 1320
rect 139 1316 140 1320
rect 134 1315 140 1316
rect 238 1320 244 1321
rect 238 1316 239 1320
rect 243 1316 244 1320
rect 238 1315 244 1316
rect 366 1320 372 1321
rect 366 1316 367 1320
rect 371 1316 372 1320
rect 366 1315 372 1316
rect 478 1320 484 1321
rect 478 1316 479 1320
rect 483 1316 484 1320
rect 478 1315 484 1316
rect 582 1320 588 1321
rect 582 1316 583 1320
rect 587 1316 588 1320
rect 582 1315 588 1316
rect 686 1320 692 1321
rect 686 1316 687 1320
rect 691 1316 692 1320
rect 686 1315 692 1316
rect 782 1320 788 1321
rect 782 1316 783 1320
rect 787 1316 788 1320
rect 782 1315 788 1316
rect 878 1320 884 1321
rect 878 1316 879 1320
rect 883 1316 884 1320
rect 878 1315 884 1316
rect 974 1320 980 1321
rect 974 1316 975 1320
rect 979 1316 980 1320
rect 1326 1320 1332 1321
rect 2502 1320 2508 1321
rect 974 1315 980 1316
rect 1286 1317 1292 1318
rect 110 1312 116 1313
rect 1286 1313 1287 1317
rect 1291 1313 1292 1317
rect 1326 1316 1327 1320
rect 1331 1316 1332 1320
rect 1326 1315 1332 1316
rect 1598 1319 1604 1320
rect 1598 1315 1599 1319
rect 1603 1315 1604 1319
rect 1598 1314 1604 1315
rect 1619 1319 1625 1320
rect 1619 1315 1620 1319
rect 1624 1318 1625 1319
rect 1642 1319 1648 1320
rect 1642 1318 1643 1319
rect 1624 1316 1643 1318
rect 1624 1315 1625 1316
rect 1619 1314 1625 1315
rect 1642 1315 1643 1316
rect 1647 1315 1648 1319
rect 1642 1314 1648 1315
rect 1662 1319 1668 1320
rect 1662 1315 1663 1319
rect 1667 1315 1668 1319
rect 1662 1314 1668 1315
rect 1683 1319 1689 1320
rect 1683 1315 1684 1319
rect 1688 1318 1689 1319
rect 1722 1319 1728 1320
rect 1722 1318 1723 1319
rect 1688 1316 1723 1318
rect 1688 1315 1689 1316
rect 1683 1314 1689 1315
rect 1722 1315 1723 1316
rect 1727 1315 1728 1319
rect 1722 1314 1728 1315
rect 1742 1319 1748 1320
rect 1742 1315 1743 1319
rect 1747 1315 1748 1319
rect 1742 1314 1748 1315
rect 1763 1319 1769 1320
rect 1763 1315 1764 1319
rect 1768 1318 1769 1319
rect 1778 1319 1784 1320
rect 1778 1318 1779 1319
rect 1768 1316 1779 1318
rect 1768 1315 1769 1316
rect 1763 1314 1769 1315
rect 1778 1315 1779 1316
rect 1783 1315 1784 1319
rect 1778 1314 1784 1315
rect 1822 1319 1828 1320
rect 1822 1315 1823 1319
rect 1827 1315 1828 1319
rect 1822 1314 1828 1315
rect 1843 1319 1849 1320
rect 1843 1315 1844 1319
rect 1848 1318 1849 1319
rect 1886 1319 1892 1320
rect 1886 1318 1887 1319
rect 1848 1316 1887 1318
rect 1848 1315 1849 1316
rect 1843 1314 1849 1315
rect 1886 1315 1887 1316
rect 1891 1315 1892 1319
rect 1886 1314 1892 1315
rect 1910 1319 1916 1320
rect 1910 1315 1911 1319
rect 1915 1315 1916 1319
rect 1910 1314 1916 1315
rect 1930 1319 1937 1320
rect 1930 1315 1931 1319
rect 1936 1315 1937 1319
rect 1930 1314 1937 1315
rect 1998 1319 2004 1320
rect 1998 1315 1999 1319
rect 2003 1315 2004 1319
rect 2019 1319 2025 1320
rect 2019 1318 2020 1319
rect 1998 1314 2004 1315
rect 2008 1316 2020 1318
rect 1286 1312 1292 1313
rect 2008 1306 2010 1316
rect 2019 1315 2020 1316
rect 2024 1315 2025 1319
rect 2019 1314 2025 1315
rect 2078 1319 2084 1320
rect 2078 1315 2079 1319
rect 2083 1315 2084 1319
rect 2078 1314 2084 1315
rect 2099 1319 2105 1320
rect 2099 1315 2100 1319
rect 2104 1318 2105 1319
rect 2138 1319 2144 1320
rect 2138 1318 2139 1319
rect 2104 1316 2139 1318
rect 2104 1315 2105 1316
rect 2099 1314 2105 1315
rect 2138 1315 2139 1316
rect 2143 1315 2144 1319
rect 2138 1314 2144 1315
rect 2158 1319 2164 1320
rect 2158 1315 2159 1319
rect 2163 1315 2164 1319
rect 2158 1314 2164 1315
rect 2179 1319 2185 1320
rect 2179 1315 2180 1319
rect 2184 1318 2185 1319
rect 2218 1319 2224 1320
rect 2218 1318 2219 1319
rect 2184 1316 2219 1318
rect 2184 1315 2185 1316
rect 2179 1314 2185 1315
rect 2218 1315 2219 1316
rect 2223 1315 2224 1319
rect 2218 1314 2224 1315
rect 2238 1319 2244 1320
rect 2238 1315 2239 1319
rect 2243 1315 2244 1319
rect 2238 1314 2244 1315
rect 2259 1319 2265 1320
rect 2259 1315 2260 1319
rect 2264 1318 2265 1319
rect 2298 1319 2304 1320
rect 2298 1318 2299 1319
rect 2264 1316 2299 1318
rect 2264 1315 2265 1316
rect 2259 1314 2265 1315
rect 2298 1315 2299 1316
rect 2303 1315 2304 1319
rect 2298 1314 2304 1315
rect 2318 1319 2324 1320
rect 2318 1315 2319 1319
rect 2323 1315 2324 1319
rect 2339 1319 2345 1320
rect 2339 1318 2340 1319
rect 2318 1314 2324 1315
rect 2328 1316 2340 1318
rect 2328 1306 2330 1316
rect 2339 1315 2340 1316
rect 2344 1315 2345 1319
rect 2339 1314 2345 1315
rect 2398 1319 2404 1320
rect 2398 1315 2399 1319
rect 2403 1315 2404 1319
rect 2398 1314 2404 1315
rect 2414 1319 2425 1320
rect 2414 1315 2415 1319
rect 2419 1315 2420 1319
rect 2424 1315 2425 1319
rect 2414 1314 2425 1315
rect 2454 1319 2460 1320
rect 2454 1315 2455 1319
rect 2459 1315 2460 1319
rect 2454 1314 2460 1315
rect 2470 1319 2481 1320
rect 2470 1315 2471 1319
rect 2475 1315 2476 1319
rect 2480 1315 2481 1319
rect 2502 1316 2503 1320
rect 2507 1316 2508 1320
rect 2502 1315 2508 1316
rect 2470 1314 2481 1315
rect 1804 1304 2010 1306
rect 2060 1304 2330 1306
rect 1804 1302 1806 1304
rect 2060 1302 2062 1304
rect 1803 1301 1809 1302
rect 110 1300 116 1301
rect 1286 1300 1292 1301
rect 110 1296 111 1300
rect 115 1296 116 1300
rect 110 1295 116 1296
rect 150 1299 156 1300
rect 150 1295 151 1299
rect 155 1295 156 1299
rect 150 1294 156 1295
rect 158 1299 164 1300
rect 158 1295 159 1299
rect 163 1298 164 1299
rect 171 1299 177 1300
rect 171 1298 172 1299
rect 163 1296 172 1298
rect 163 1295 164 1296
rect 158 1294 164 1295
rect 171 1295 172 1296
rect 176 1295 177 1299
rect 171 1294 177 1295
rect 254 1299 260 1300
rect 254 1295 255 1299
rect 259 1295 260 1299
rect 254 1294 260 1295
rect 275 1299 281 1300
rect 275 1295 276 1299
rect 280 1298 281 1299
rect 362 1299 368 1300
rect 362 1298 363 1299
rect 280 1296 363 1298
rect 280 1295 281 1296
rect 275 1294 281 1295
rect 362 1295 363 1296
rect 367 1295 368 1299
rect 362 1294 368 1295
rect 382 1299 388 1300
rect 382 1295 383 1299
rect 387 1295 388 1299
rect 403 1299 409 1300
rect 403 1298 404 1299
rect 382 1294 388 1295
rect 392 1296 404 1298
rect 392 1286 394 1296
rect 403 1295 404 1296
rect 408 1295 409 1299
rect 403 1294 409 1295
rect 494 1299 500 1300
rect 494 1295 495 1299
rect 499 1295 500 1299
rect 494 1294 500 1295
rect 515 1299 521 1300
rect 515 1295 516 1299
rect 520 1298 521 1299
rect 578 1299 584 1300
rect 578 1298 579 1299
rect 520 1296 579 1298
rect 520 1295 521 1296
rect 515 1294 521 1295
rect 578 1295 579 1296
rect 583 1295 584 1299
rect 578 1294 584 1295
rect 598 1299 604 1300
rect 598 1295 599 1299
rect 603 1295 604 1299
rect 598 1294 604 1295
rect 619 1299 625 1300
rect 619 1295 620 1299
rect 624 1298 625 1299
rect 654 1299 660 1300
rect 654 1298 655 1299
rect 624 1296 655 1298
rect 624 1295 625 1296
rect 619 1294 625 1295
rect 654 1295 655 1296
rect 659 1295 660 1299
rect 654 1294 660 1295
rect 702 1299 708 1300
rect 702 1295 703 1299
rect 707 1295 708 1299
rect 702 1294 708 1295
rect 723 1299 729 1300
rect 723 1295 724 1299
rect 728 1298 729 1299
rect 746 1299 752 1300
rect 746 1298 747 1299
rect 728 1296 747 1298
rect 728 1295 729 1296
rect 723 1294 729 1295
rect 746 1295 747 1296
rect 751 1295 752 1299
rect 746 1294 752 1295
rect 798 1299 804 1300
rect 798 1295 799 1299
rect 803 1295 804 1299
rect 798 1294 804 1295
rect 806 1299 812 1300
rect 806 1295 807 1299
rect 811 1298 812 1299
rect 819 1299 825 1300
rect 819 1298 820 1299
rect 811 1296 820 1298
rect 811 1295 812 1296
rect 806 1294 812 1295
rect 819 1295 820 1296
rect 824 1295 825 1299
rect 819 1294 825 1295
rect 894 1299 900 1300
rect 894 1295 895 1299
rect 899 1295 900 1299
rect 915 1299 921 1300
rect 915 1298 916 1299
rect 894 1294 900 1295
rect 904 1296 916 1298
rect 904 1290 906 1296
rect 915 1295 916 1296
rect 920 1295 921 1299
rect 915 1294 921 1295
rect 990 1299 996 1300
rect 990 1295 991 1299
rect 995 1295 996 1299
rect 1011 1299 1017 1300
rect 1011 1298 1012 1299
rect 990 1294 996 1295
rect 1000 1296 1012 1298
rect 132 1284 394 1286
rect 780 1288 906 1290
rect 132 1282 134 1284
rect 780 1282 782 1288
rect 1000 1286 1002 1296
rect 1011 1295 1012 1296
rect 1016 1295 1017 1299
rect 1286 1296 1287 1300
rect 1291 1296 1292 1300
rect 1286 1295 1292 1296
rect 1579 1299 1588 1300
rect 1579 1295 1580 1299
rect 1587 1295 1588 1299
rect 1011 1294 1017 1295
rect 1579 1294 1588 1295
rect 1642 1299 1649 1300
rect 1642 1295 1643 1299
rect 1648 1295 1649 1299
rect 1642 1294 1649 1295
rect 1722 1299 1729 1300
rect 1722 1295 1723 1299
rect 1728 1295 1729 1299
rect 1803 1297 1804 1301
rect 1808 1297 1809 1301
rect 2059 1301 2065 1302
rect 1803 1296 1809 1297
rect 1886 1299 1897 1300
rect 1722 1294 1729 1295
rect 1886 1295 1887 1299
rect 1891 1295 1892 1299
rect 1896 1295 1897 1299
rect 1886 1294 1897 1295
rect 1979 1299 1985 1300
rect 1979 1295 1980 1299
rect 1984 1298 1985 1299
rect 2010 1299 2016 1300
rect 2010 1298 2011 1299
rect 1984 1296 2011 1298
rect 1984 1295 1985 1296
rect 1979 1294 1985 1295
rect 2010 1295 2011 1296
rect 2015 1295 2016 1299
rect 2059 1297 2060 1301
rect 2064 1297 2065 1301
rect 2059 1296 2065 1297
rect 2138 1299 2145 1300
rect 2010 1294 2016 1295
rect 2138 1295 2139 1299
rect 2144 1295 2145 1299
rect 2138 1294 2145 1295
rect 2218 1299 2225 1300
rect 2218 1295 2219 1299
rect 2224 1295 2225 1299
rect 2218 1294 2225 1295
rect 2299 1299 2305 1300
rect 2299 1295 2300 1299
rect 2304 1298 2305 1299
rect 2326 1299 2332 1300
rect 2326 1298 2327 1299
rect 2304 1296 2327 1298
rect 2304 1295 2305 1296
rect 2299 1294 2305 1295
rect 2326 1295 2327 1296
rect 2331 1295 2332 1299
rect 2326 1294 2332 1295
rect 2379 1299 2385 1300
rect 2379 1295 2380 1299
rect 2384 1298 2385 1299
rect 2390 1299 2396 1300
rect 2390 1298 2391 1299
rect 2384 1296 2391 1298
rect 2384 1295 2385 1296
rect 2379 1294 2385 1295
rect 2390 1295 2391 1296
rect 2395 1295 2396 1299
rect 2390 1294 2396 1295
rect 2435 1299 2441 1300
rect 2435 1295 2436 1299
rect 2440 1298 2441 1299
rect 2462 1299 2468 1300
rect 2462 1298 2463 1299
rect 2440 1296 2463 1298
rect 2440 1295 2441 1296
rect 2435 1294 2441 1295
rect 2462 1295 2463 1296
rect 2467 1295 2468 1299
rect 2462 1294 2468 1295
rect 876 1284 1002 1286
rect 1547 1287 1553 1288
rect 876 1282 878 1284
rect 1547 1283 1548 1287
rect 1552 1286 1553 1287
rect 1606 1287 1617 1288
rect 1552 1284 1602 1286
rect 1552 1283 1553 1284
rect 1547 1282 1553 1283
rect 131 1281 137 1282
rect 131 1277 132 1281
rect 136 1277 137 1281
rect 779 1281 785 1282
rect 131 1276 137 1277
rect 235 1279 241 1280
rect 235 1275 236 1279
rect 240 1278 241 1279
rect 246 1279 252 1280
rect 246 1278 247 1279
rect 240 1276 247 1278
rect 240 1275 241 1276
rect 235 1274 241 1275
rect 246 1275 247 1276
rect 251 1275 252 1279
rect 246 1274 252 1275
rect 362 1279 369 1280
rect 362 1275 363 1279
rect 368 1275 369 1279
rect 362 1274 369 1275
rect 475 1279 481 1280
rect 475 1275 476 1279
rect 480 1278 481 1279
rect 570 1279 576 1280
rect 570 1278 571 1279
rect 480 1276 571 1278
rect 480 1275 481 1276
rect 475 1274 481 1275
rect 570 1275 571 1276
rect 575 1275 576 1279
rect 570 1274 576 1275
rect 578 1279 585 1280
rect 578 1275 579 1279
rect 584 1275 585 1279
rect 578 1274 585 1275
rect 683 1279 689 1280
rect 683 1275 684 1279
rect 688 1278 689 1279
rect 688 1276 754 1278
rect 779 1277 780 1281
rect 784 1277 785 1281
rect 779 1276 785 1277
rect 875 1281 881 1282
rect 875 1277 876 1281
rect 880 1277 881 1281
rect 875 1276 881 1277
rect 966 1279 977 1280
rect 688 1275 689 1276
rect 683 1274 689 1275
rect 752 1274 754 1276
rect 806 1275 812 1276
rect 806 1274 807 1275
rect 752 1272 807 1274
rect 806 1271 807 1272
rect 811 1271 812 1275
rect 966 1275 967 1279
rect 971 1275 972 1279
rect 976 1275 977 1279
rect 966 1274 977 1275
rect 1600 1274 1602 1284
rect 1606 1283 1607 1287
rect 1611 1283 1612 1287
rect 1616 1283 1617 1287
rect 1606 1282 1617 1283
rect 1691 1287 1697 1288
rect 1691 1283 1692 1287
rect 1696 1286 1697 1287
rect 1778 1287 1785 1288
rect 1696 1284 1774 1286
rect 1696 1283 1697 1284
rect 1691 1282 1697 1283
rect 1772 1274 1774 1284
rect 1778 1283 1779 1287
rect 1784 1283 1785 1287
rect 1778 1282 1785 1283
rect 1830 1287 1836 1288
rect 1830 1283 1831 1287
rect 1835 1286 1836 1287
rect 1875 1287 1881 1288
rect 1875 1286 1876 1287
rect 1835 1284 1876 1286
rect 1835 1283 1836 1284
rect 1830 1282 1836 1283
rect 1875 1283 1876 1284
rect 1880 1283 1881 1287
rect 1875 1282 1881 1283
rect 1971 1287 1977 1288
rect 1971 1283 1972 1287
rect 1976 1286 1977 1287
rect 2066 1287 2072 1288
rect 2066 1286 2067 1287
rect 1976 1284 2067 1286
rect 1976 1283 1977 1284
rect 1971 1282 1977 1283
rect 2066 1283 2067 1284
rect 2071 1283 2072 1287
rect 2066 1282 2072 1283
rect 2075 1287 2081 1288
rect 2075 1283 2076 1287
rect 2080 1286 2081 1287
rect 2187 1287 2193 1288
rect 2080 1284 2182 1286
rect 2080 1283 2081 1284
rect 2075 1282 2081 1283
rect 2180 1274 2182 1284
rect 2187 1283 2188 1287
rect 2192 1286 2193 1287
rect 2298 1287 2305 1288
rect 2192 1284 2294 1286
rect 2192 1283 2193 1284
rect 2187 1282 2193 1283
rect 2292 1274 2294 1284
rect 2298 1283 2299 1287
rect 2304 1283 2305 1287
rect 2298 1282 2305 1283
rect 1600 1272 1654 1274
rect 1772 1272 1918 1274
rect 2180 1272 2230 1274
rect 2292 1272 2342 1274
rect 806 1270 812 1271
rect 1652 1270 1654 1272
rect 1916 1270 1918 1272
rect 2228 1270 2230 1272
rect 2340 1270 2342 1272
rect 1566 1269 1572 1270
rect 1326 1268 1332 1269
rect 1326 1264 1327 1268
rect 1331 1264 1332 1268
rect 1566 1265 1567 1269
rect 1571 1265 1572 1269
rect 1630 1269 1636 1270
rect 1566 1264 1572 1265
rect 1582 1267 1593 1268
rect 1326 1263 1332 1264
rect 1582 1263 1583 1267
rect 1587 1263 1588 1267
rect 1592 1263 1593 1267
rect 1630 1265 1631 1269
rect 1635 1265 1636 1269
rect 1630 1264 1636 1265
rect 1651 1269 1657 1270
rect 1651 1265 1652 1269
rect 1656 1265 1657 1269
rect 1651 1264 1657 1265
rect 1710 1269 1716 1270
rect 1710 1265 1711 1269
rect 1715 1265 1716 1269
rect 1798 1269 1804 1270
rect 1710 1264 1716 1265
rect 1718 1267 1724 1268
rect 1582 1262 1593 1263
rect 1718 1263 1719 1267
rect 1723 1266 1724 1267
rect 1731 1267 1737 1268
rect 1731 1266 1732 1267
rect 1723 1264 1732 1266
rect 1723 1263 1724 1264
rect 1718 1262 1724 1263
rect 1731 1263 1732 1264
rect 1736 1263 1737 1267
rect 1798 1265 1799 1269
rect 1803 1265 1804 1269
rect 1894 1269 1900 1270
rect 1798 1264 1804 1265
rect 1819 1267 1825 1268
rect 1731 1262 1737 1263
rect 1819 1263 1820 1267
rect 1824 1266 1825 1267
rect 1830 1267 1836 1268
rect 1830 1266 1831 1267
rect 1824 1264 1831 1266
rect 1824 1263 1825 1264
rect 1819 1262 1825 1263
rect 1830 1263 1831 1264
rect 1835 1263 1836 1267
rect 1894 1265 1895 1269
rect 1899 1265 1900 1269
rect 1894 1264 1900 1265
rect 1915 1269 1921 1270
rect 1915 1265 1916 1269
rect 1920 1265 1921 1269
rect 1915 1264 1921 1265
rect 1990 1269 1996 1270
rect 1990 1265 1991 1269
rect 1995 1265 1996 1269
rect 2094 1269 2100 1270
rect 1990 1264 1996 1265
rect 2010 1267 2017 1268
rect 1830 1262 1836 1263
rect 2010 1263 2011 1267
rect 2016 1263 2017 1267
rect 2094 1265 2095 1269
rect 2099 1265 2100 1269
rect 2206 1269 2212 1270
rect 2094 1264 2100 1265
rect 2110 1267 2121 1268
rect 2010 1262 2017 1263
rect 2110 1263 2111 1267
rect 2115 1263 2116 1267
rect 2120 1263 2121 1267
rect 2206 1265 2207 1269
rect 2211 1265 2212 1269
rect 2206 1264 2212 1265
rect 2227 1269 2233 1270
rect 2227 1265 2228 1269
rect 2232 1265 2233 1269
rect 2227 1264 2233 1265
rect 2318 1269 2324 1270
rect 2318 1265 2319 1269
rect 2323 1265 2324 1269
rect 2318 1264 2324 1265
rect 2339 1269 2345 1270
rect 2339 1265 2340 1269
rect 2344 1265 2345 1269
rect 2339 1264 2345 1265
rect 2502 1268 2508 1269
rect 2502 1264 2503 1268
rect 2507 1264 2508 1268
rect 2502 1263 2508 1264
rect 2110 1262 2121 1263
rect 131 1259 137 1260
rect 131 1255 132 1259
rect 136 1258 137 1259
rect 158 1259 164 1260
rect 158 1258 159 1259
rect 136 1256 159 1258
rect 136 1255 137 1256
rect 131 1254 137 1255
rect 158 1255 159 1256
rect 163 1255 164 1259
rect 158 1254 164 1255
rect 183 1259 189 1260
rect 183 1255 184 1259
rect 188 1258 189 1259
rect 195 1259 201 1260
rect 195 1258 196 1259
rect 188 1256 196 1258
rect 188 1255 189 1256
rect 183 1254 189 1255
rect 195 1255 196 1256
rect 200 1255 201 1259
rect 195 1254 201 1255
rect 238 1259 244 1260
rect 238 1255 239 1259
rect 243 1258 244 1259
rect 283 1259 289 1260
rect 283 1258 284 1259
rect 243 1256 284 1258
rect 243 1255 244 1256
rect 238 1254 244 1255
rect 283 1255 284 1256
rect 288 1255 289 1259
rect 283 1254 289 1255
rect 326 1259 332 1260
rect 326 1255 327 1259
rect 331 1258 332 1259
rect 371 1259 377 1260
rect 371 1258 372 1259
rect 331 1256 372 1258
rect 331 1255 332 1256
rect 326 1254 332 1255
rect 371 1255 372 1256
rect 376 1255 377 1259
rect 371 1254 377 1255
rect 451 1259 457 1260
rect 451 1255 452 1259
rect 456 1258 457 1259
rect 462 1259 468 1260
rect 462 1258 463 1259
rect 456 1256 463 1258
rect 456 1255 457 1256
rect 451 1254 457 1255
rect 462 1255 463 1256
rect 467 1255 468 1259
rect 462 1254 468 1255
rect 502 1259 508 1260
rect 502 1255 503 1259
rect 507 1258 508 1259
rect 531 1259 537 1260
rect 531 1258 532 1259
rect 507 1256 532 1258
rect 507 1255 508 1256
rect 502 1254 508 1255
rect 531 1255 532 1256
rect 536 1255 537 1259
rect 531 1254 537 1255
rect 603 1259 609 1260
rect 603 1255 604 1259
rect 608 1258 609 1259
rect 675 1259 681 1260
rect 608 1256 670 1258
rect 608 1255 609 1256
rect 603 1254 609 1255
rect 668 1246 670 1256
rect 675 1255 676 1259
rect 680 1255 681 1259
rect 675 1254 681 1255
rect 746 1259 753 1260
rect 746 1255 747 1259
rect 752 1255 753 1259
rect 746 1254 753 1255
rect 790 1259 796 1260
rect 790 1255 791 1259
rect 795 1258 796 1259
rect 819 1259 825 1260
rect 819 1258 820 1259
rect 795 1256 820 1258
rect 795 1255 796 1256
rect 790 1254 796 1255
rect 819 1255 820 1256
rect 824 1255 825 1259
rect 819 1254 825 1255
rect 862 1259 868 1260
rect 862 1255 863 1259
rect 867 1258 868 1259
rect 899 1259 905 1260
rect 899 1258 900 1259
rect 867 1256 900 1258
rect 867 1255 868 1256
rect 862 1254 868 1255
rect 899 1255 900 1256
rect 904 1255 905 1259
rect 899 1254 905 1255
rect 677 1250 679 1254
rect 1326 1251 1332 1252
rect 677 1248 943 1250
rect 668 1244 719 1246
rect 717 1242 719 1244
rect 941 1242 943 1248
rect 1326 1247 1327 1251
rect 1331 1247 1332 1251
rect 2502 1251 2508 1252
rect 1326 1246 1332 1247
rect 1550 1248 1556 1249
rect 1550 1244 1551 1248
rect 1555 1244 1556 1248
rect 1550 1243 1556 1244
rect 1614 1248 1620 1249
rect 1614 1244 1615 1248
rect 1619 1244 1620 1248
rect 1614 1243 1620 1244
rect 1694 1248 1700 1249
rect 1694 1244 1695 1248
rect 1699 1244 1700 1248
rect 1694 1243 1700 1244
rect 1782 1248 1788 1249
rect 1782 1244 1783 1248
rect 1787 1244 1788 1248
rect 1782 1243 1788 1244
rect 1878 1248 1884 1249
rect 1878 1244 1879 1248
rect 1883 1244 1884 1248
rect 1878 1243 1884 1244
rect 1974 1248 1980 1249
rect 1974 1244 1975 1248
rect 1979 1244 1980 1248
rect 1974 1243 1980 1244
rect 2078 1248 2084 1249
rect 2078 1244 2079 1248
rect 2083 1244 2084 1248
rect 2078 1243 2084 1244
rect 2190 1248 2196 1249
rect 2190 1244 2191 1248
rect 2195 1244 2196 1248
rect 2190 1243 2196 1244
rect 2302 1248 2308 1249
rect 2302 1244 2303 1248
rect 2307 1244 2308 1248
rect 2502 1247 2503 1251
rect 2507 1247 2508 1251
rect 2502 1246 2508 1247
rect 2302 1243 2308 1244
rect 150 1241 156 1242
rect 110 1240 116 1241
rect 110 1236 111 1240
rect 115 1236 116 1240
rect 150 1237 151 1241
rect 155 1237 156 1241
rect 214 1241 220 1242
rect 150 1236 156 1237
rect 171 1239 177 1240
rect 110 1235 116 1236
rect 171 1235 172 1239
rect 176 1238 177 1239
rect 183 1239 189 1240
rect 183 1238 184 1239
rect 176 1236 184 1238
rect 176 1235 177 1236
rect 171 1234 177 1235
rect 183 1235 184 1236
rect 188 1235 189 1239
rect 214 1237 215 1241
rect 219 1237 220 1241
rect 302 1241 308 1242
rect 214 1236 220 1237
rect 235 1239 244 1240
rect 183 1234 189 1235
rect 235 1235 236 1239
rect 243 1235 244 1239
rect 302 1237 303 1241
rect 307 1237 308 1241
rect 390 1241 396 1242
rect 302 1236 308 1237
rect 323 1239 332 1240
rect 235 1234 244 1235
rect 323 1235 324 1239
rect 331 1235 332 1239
rect 390 1237 391 1241
rect 395 1237 396 1241
rect 470 1241 476 1242
rect 390 1236 396 1237
rect 398 1239 404 1240
rect 323 1234 332 1235
rect 398 1235 399 1239
rect 403 1238 404 1239
rect 411 1239 417 1240
rect 411 1238 412 1239
rect 403 1236 412 1238
rect 403 1235 404 1236
rect 398 1234 404 1235
rect 411 1235 412 1236
rect 416 1235 417 1239
rect 470 1237 471 1241
rect 475 1237 476 1241
rect 550 1241 556 1242
rect 470 1236 476 1237
rect 491 1239 497 1240
rect 411 1234 417 1235
rect 491 1235 492 1239
rect 496 1238 497 1239
rect 502 1239 508 1240
rect 502 1238 503 1239
rect 496 1236 503 1238
rect 496 1235 497 1236
rect 491 1234 497 1235
rect 502 1235 503 1236
rect 507 1235 508 1239
rect 550 1237 551 1241
rect 555 1237 556 1241
rect 622 1241 628 1242
rect 550 1236 556 1237
rect 570 1239 577 1240
rect 502 1234 508 1235
rect 570 1235 571 1239
rect 576 1235 577 1239
rect 622 1237 623 1241
rect 627 1237 628 1241
rect 694 1241 700 1242
rect 622 1236 628 1237
rect 630 1239 636 1240
rect 570 1234 577 1235
rect 630 1235 631 1239
rect 635 1238 636 1239
rect 643 1239 649 1240
rect 643 1238 644 1239
rect 635 1236 644 1238
rect 635 1235 636 1236
rect 630 1234 636 1235
rect 643 1235 644 1236
rect 648 1235 649 1239
rect 694 1237 695 1241
rect 699 1237 700 1241
rect 694 1236 700 1237
rect 715 1241 721 1242
rect 715 1237 716 1241
rect 720 1237 721 1241
rect 715 1236 721 1237
rect 766 1241 772 1242
rect 766 1237 767 1241
rect 771 1237 772 1241
rect 838 1241 844 1242
rect 766 1236 772 1237
rect 787 1239 796 1240
rect 643 1234 649 1235
rect 787 1235 788 1239
rect 795 1235 796 1239
rect 838 1237 839 1241
rect 843 1237 844 1241
rect 918 1241 924 1242
rect 838 1236 844 1237
rect 859 1239 868 1240
rect 787 1234 796 1235
rect 859 1235 860 1239
rect 867 1235 868 1239
rect 918 1237 919 1241
rect 923 1237 924 1241
rect 918 1236 924 1237
rect 939 1241 945 1242
rect 939 1237 940 1241
rect 944 1237 945 1241
rect 939 1236 945 1237
rect 1286 1240 1292 1241
rect 1286 1236 1287 1240
rect 1291 1236 1292 1240
rect 1286 1235 1292 1236
rect 859 1234 868 1235
rect 1518 1232 1524 1233
rect 1326 1229 1332 1230
rect 1326 1225 1327 1229
rect 1331 1225 1332 1229
rect 1518 1228 1519 1232
rect 1523 1228 1524 1232
rect 1518 1227 1524 1228
rect 1574 1232 1580 1233
rect 1574 1228 1575 1232
rect 1579 1228 1580 1232
rect 1574 1227 1580 1228
rect 1630 1232 1636 1233
rect 1630 1228 1631 1232
rect 1635 1228 1636 1232
rect 1630 1227 1636 1228
rect 1686 1232 1692 1233
rect 1686 1228 1687 1232
rect 1691 1228 1692 1232
rect 1686 1227 1692 1228
rect 1742 1232 1748 1233
rect 1742 1228 1743 1232
rect 1747 1228 1748 1232
rect 1742 1227 1748 1228
rect 1798 1232 1804 1233
rect 1798 1228 1799 1232
rect 1803 1228 1804 1232
rect 1798 1227 1804 1228
rect 1854 1232 1860 1233
rect 1854 1228 1855 1232
rect 1859 1228 1860 1232
rect 1854 1227 1860 1228
rect 1910 1232 1916 1233
rect 1910 1228 1911 1232
rect 1915 1228 1916 1232
rect 1910 1227 1916 1228
rect 1966 1232 1972 1233
rect 1966 1228 1967 1232
rect 1971 1228 1972 1232
rect 1966 1227 1972 1228
rect 2030 1232 2036 1233
rect 2030 1228 2031 1232
rect 2035 1228 2036 1232
rect 2030 1227 2036 1228
rect 2102 1232 2108 1233
rect 2102 1228 2103 1232
rect 2107 1228 2108 1232
rect 2102 1227 2108 1228
rect 2182 1232 2188 1233
rect 2182 1228 2183 1232
rect 2187 1228 2188 1232
rect 2182 1227 2188 1228
rect 2270 1232 2276 1233
rect 2270 1228 2271 1232
rect 2275 1228 2276 1232
rect 2270 1227 2276 1228
rect 2366 1232 2372 1233
rect 2366 1228 2367 1232
rect 2371 1228 2372 1232
rect 2366 1227 2372 1228
rect 2438 1232 2444 1233
rect 2438 1228 2439 1232
rect 2443 1228 2444 1232
rect 2438 1227 2444 1228
rect 2502 1229 2508 1230
rect 1326 1224 1332 1225
rect 2502 1225 2503 1229
rect 2507 1225 2508 1229
rect 2502 1224 2508 1225
rect 110 1223 116 1224
rect 110 1219 111 1223
rect 115 1219 116 1223
rect 1286 1223 1292 1224
rect 110 1218 116 1219
rect 134 1220 140 1221
rect 134 1216 135 1220
rect 139 1216 140 1220
rect 134 1215 140 1216
rect 198 1220 204 1221
rect 198 1216 199 1220
rect 203 1216 204 1220
rect 198 1215 204 1216
rect 286 1220 292 1221
rect 286 1216 287 1220
rect 291 1216 292 1220
rect 286 1215 292 1216
rect 374 1220 380 1221
rect 374 1216 375 1220
rect 379 1216 380 1220
rect 374 1215 380 1216
rect 454 1220 460 1221
rect 454 1216 455 1220
rect 459 1216 460 1220
rect 454 1215 460 1216
rect 534 1220 540 1221
rect 534 1216 535 1220
rect 539 1216 540 1220
rect 534 1215 540 1216
rect 606 1220 612 1221
rect 606 1216 607 1220
rect 611 1216 612 1220
rect 606 1215 612 1216
rect 678 1220 684 1221
rect 678 1216 679 1220
rect 683 1216 684 1220
rect 678 1215 684 1216
rect 750 1220 756 1221
rect 750 1216 751 1220
rect 755 1216 756 1220
rect 750 1215 756 1216
rect 822 1220 828 1221
rect 822 1216 823 1220
rect 827 1216 828 1220
rect 822 1215 828 1216
rect 902 1220 908 1221
rect 902 1216 903 1220
rect 907 1216 908 1220
rect 1286 1219 1287 1223
rect 1291 1219 1292 1223
rect 1286 1218 1292 1219
rect 902 1215 908 1216
rect 1326 1212 1332 1213
rect 2502 1212 2508 1213
rect 1326 1208 1327 1212
rect 1331 1208 1332 1212
rect 1326 1207 1332 1208
rect 1534 1211 1540 1212
rect 1534 1207 1535 1211
rect 1539 1207 1540 1211
rect 1534 1206 1540 1207
rect 1555 1211 1561 1212
rect 1555 1207 1556 1211
rect 1560 1210 1561 1211
rect 1570 1211 1576 1212
rect 1570 1210 1571 1211
rect 1560 1208 1571 1210
rect 1560 1207 1561 1208
rect 1555 1206 1561 1207
rect 1570 1207 1571 1208
rect 1575 1207 1576 1211
rect 1570 1206 1576 1207
rect 1590 1211 1596 1212
rect 1590 1207 1591 1211
rect 1595 1207 1596 1211
rect 1590 1206 1596 1207
rect 1606 1211 1617 1212
rect 1606 1207 1607 1211
rect 1611 1207 1612 1211
rect 1616 1207 1617 1211
rect 1606 1206 1617 1207
rect 1646 1211 1652 1212
rect 1646 1207 1647 1211
rect 1651 1207 1652 1211
rect 1646 1206 1652 1207
rect 1667 1211 1673 1212
rect 1667 1207 1668 1211
rect 1672 1210 1673 1211
rect 1682 1211 1688 1212
rect 1682 1210 1683 1211
rect 1672 1208 1683 1210
rect 1672 1207 1673 1208
rect 1667 1206 1673 1207
rect 1682 1207 1683 1208
rect 1687 1207 1688 1211
rect 1682 1206 1688 1207
rect 1702 1211 1708 1212
rect 1702 1207 1703 1211
rect 1707 1207 1708 1211
rect 1702 1206 1708 1207
rect 1723 1211 1729 1212
rect 1723 1207 1724 1211
rect 1728 1210 1729 1211
rect 1738 1211 1744 1212
rect 1738 1210 1739 1211
rect 1728 1208 1739 1210
rect 1728 1207 1729 1208
rect 1723 1206 1729 1207
rect 1738 1207 1739 1208
rect 1743 1207 1744 1211
rect 1738 1206 1744 1207
rect 1758 1211 1764 1212
rect 1758 1207 1759 1211
rect 1763 1207 1764 1211
rect 1758 1206 1764 1207
rect 1779 1211 1785 1212
rect 1779 1207 1780 1211
rect 1784 1210 1785 1211
rect 1794 1211 1800 1212
rect 1794 1210 1795 1211
rect 1784 1208 1795 1210
rect 1784 1207 1785 1208
rect 1779 1206 1785 1207
rect 1794 1207 1795 1208
rect 1799 1207 1800 1211
rect 1794 1206 1800 1207
rect 1814 1211 1820 1212
rect 1814 1207 1815 1211
rect 1819 1207 1820 1211
rect 1814 1206 1820 1207
rect 1835 1211 1841 1212
rect 1835 1207 1836 1211
rect 1840 1210 1841 1211
rect 1850 1211 1856 1212
rect 1850 1210 1851 1211
rect 1840 1208 1851 1210
rect 1840 1207 1841 1208
rect 1835 1206 1841 1207
rect 1850 1207 1851 1208
rect 1855 1207 1856 1211
rect 1850 1206 1856 1207
rect 1870 1211 1876 1212
rect 1870 1207 1871 1211
rect 1875 1207 1876 1211
rect 1870 1206 1876 1207
rect 1891 1211 1897 1212
rect 1891 1207 1892 1211
rect 1896 1210 1897 1211
rect 1906 1211 1912 1212
rect 1906 1210 1907 1211
rect 1896 1208 1907 1210
rect 1896 1207 1897 1208
rect 1891 1206 1897 1207
rect 1906 1207 1907 1208
rect 1911 1207 1912 1211
rect 1906 1206 1912 1207
rect 1926 1211 1932 1212
rect 1926 1207 1927 1211
rect 1931 1207 1932 1211
rect 1926 1206 1932 1207
rect 1947 1211 1953 1212
rect 1947 1207 1948 1211
rect 1952 1210 1953 1211
rect 1962 1211 1968 1212
rect 1962 1210 1963 1211
rect 1952 1208 1963 1210
rect 1952 1207 1953 1208
rect 1947 1206 1953 1207
rect 1962 1207 1963 1208
rect 1967 1207 1968 1211
rect 1962 1206 1968 1207
rect 1982 1211 1988 1212
rect 1982 1207 1983 1211
rect 1987 1207 1988 1211
rect 1982 1206 1988 1207
rect 2003 1211 2009 1212
rect 2003 1207 2004 1211
rect 2008 1210 2009 1211
rect 2026 1211 2032 1212
rect 2026 1210 2027 1211
rect 2008 1208 2027 1210
rect 2008 1207 2009 1208
rect 2003 1206 2009 1207
rect 2026 1207 2027 1208
rect 2031 1207 2032 1211
rect 2026 1206 2032 1207
rect 2046 1211 2052 1212
rect 2046 1207 2047 1211
rect 2051 1207 2052 1211
rect 2046 1206 2052 1207
rect 2066 1211 2073 1212
rect 2066 1207 2067 1211
rect 2072 1207 2073 1211
rect 2066 1206 2073 1207
rect 2118 1211 2124 1212
rect 2118 1207 2119 1211
rect 2123 1207 2124 1211
rect 2118 1206 2124 1207
rect 2139 1211 2145 1212
rect 2139 1207 2140 1211
rect 2144 1210 2145 1211
rect 2178 1211 2184 1212
rect 2178 1210 2179 1211
rect 2144 1208 2179 1210
rect 2144 1207 2145 1208
rect 2139 1206 2145 1207
rect 2178 1207 2179 1208
rect 2183 1207 2184 1211
rect 2178 1206 2184 1207
rect 2198 1211 2204 1212
rect 2198 1207 2199 1211
rect 2203 1207 2204 1211
rect 2198 1206 2204 1207
rect 2219 1211 2225 1212
rect 2219 1207 2220 1211
rect 2224 1210 2225 1211
rect 2266 1211 2272 1212
rect 2266 1210 2267 1211
rect 2224 1208 2267 1210
rect 2224 1207 2225 1208
rect 2219 1206 2225 1207
rect 2266 1207 2267 1208
rect 2271 1207 2272 1211
rect 2266 1206 2272 1207
rect 2286 1211 2292 1212
rect 2286 1207 2287 1211
rect 2291 1207 2292 1211
rect 2286 1206 2292 1207
rect 2306 1211 2313 1212
rect 2306 1207 2307 1211
rect 2312 1207 2313 1211
rect 2306 1206 2313 1207
rect 2382 1211 2388 1212
rect 2382 1207 2383 1211
rect 2387 1207 2388 1211
rect 2382 1206 2388 1207
rect 2390 1211 2396 1212
rect 2390 1207 2391 1211
rect 2395 1210 2396 1211
rect 2403 1211 2409 1212
rect 2403 1210 2404 1211
rect 2395 1208 2404 1210
rect 2395 1207 2396 1208
rect 2390 1206 2396 1207
rect 2403 1207 2404 1208
rect 2408 1207 2409 1211
rect 2403 1206 2409 1207
rect 2454 1211 2460 1212
rect 2454 1207 2455 1211
rect 2459 1207 2460 1211
rect 2454 1206 2460 1207
rect 2462 1211 2468 1212
rect 2462 1207 2463 1211
rect 2467 1210 2468 1211
rect 2475 1211 2481 1212
rect 2475 1210 2476 1211
rect 2467 1208 2476 1210
rect 2467 1207 2468 1208
rect 2462 1206 2468 1207
rect 2475 1207 2476 1208
rect 2480 1207 2481 1211
rect 2502 1208 2503 1212
rect 2507 1208 2508 1212
rect 2502 1207 2508 1208
rect 2475 1206 2481 1207
rect 134 1204 140 1205
rect 110 1201 116 1202
rect 110 1197 111 1201
rect 115 1197 116 1201
rect 134 1200 135 1204
rect 139 1200 140 1204
rect 134 1199 140 1200
rect 190 1204 196 1205
rect 190 1200 191 1204
rect 195 1200 196 1204
rect 190 1199 196 1200
rect 270 1204 276 1205
rect 270 1200 271 1204
rect 275 1200 276 1204
rect 270 1199 276 1200
rect 350 1204 356 1205
rect 350 1200 351 1204
rect 355 1200 356 1204
rect 350 1199 356 1200
rect 430 1204 436 1205
rect 430 1200 431 1204
rect 435 1200 436 1204
rect 430 1199 436 1200
rect 510 1204 516 1205
rect 510 1200 511 1204
rect 515 1200 516 1204
rect 510 1199 516 1200
rect 582 1204 588 1205
rect 582 1200 583 1204
rect 587 1200 588 1204
rect 582 1199 588 1200
rect 646 1204 652 1205
rect 646 1200 647 1204
rect 651 1200 652 1204
rect 646 1199 652 1200
rect 718 1204 724 1205
rect 718 1200 719 1204
rect 723 1200 724 1204
rect 718 1199 724 1200
rect 790 1204 796 1205
rect 790 1200 791 1204
rect 795 1200 796 1204
rect 790 1199 796 1200
rect 862 1204 868 1205
rect 862 1200 863 1204
rect 867 1200 868 1204
rect 862 1199 868 1200
rect 1286 1201 1292 1202
rect 110 1196 116 1197
rect 1286 1197 1287 1201
rect 1291 1197 1292 1201
rect 1718 1199 1724 1200
rect 1718 1198 1719 1199
rect 1286 1196 1292 1197
rect 1628 1196 1719 1198
rect 1628 1194 1630 1196
rect 1718 1195 1719 1196
rect 1723 1195 1724 1199
rect 1718 1194 1724 1195
rect 1627 1193 1633 1194
rect 1515 1191 1521 1192
rect 1515 1187 1516 1191
rect 1520 1190 1521 1191
rect 1570 1191 1577 1192
rect 1520 1188 1566 1190
rect 1520 1187 1521 1188
rect 1515 1186 1521 1187
rect 110 1184 116 1185
rect 1286 1184 1292 1185
rect 110 1180 111 1184
rect 115 1180 116 1184
rect 110 1179 116 1180
rect 150 1183 156 1184
rect 150 1179 151 1183
rect 155 1179 156 1183
rect 150 1178 156 1179
rect 171 1183 177 1184
rect 171 1179 172 1183
rect 176 1182 177 1183
rect 186 1183 192 1184
rect 186 1182 187 1183
rect 176 1180 187 1182
rect 176 1179 177 1180
rect 171 1178 177 1179
rect 186 1179 187 1180
rect 191 1179 192 1183
rect 186 1178 192 1179
rect 206 1183 212 1184
rect 206 1179 207 1183
rect 211 1179 212 1183
rect 206 1178 212 1179
rect 227 1183 233 1184
rect 227 1179 228 1183
rect 232 1182 233 1183
rect 266 1183 272 1184
rect 266 1182 267 1183
rect 232 1180 267 1182
rect 232 1179 233 1180
rect 227 1178 233 1179
rect 266 1179 267 1180
rect 271 1179 272 1183
rect 266 1178 272 1179
rect 286 1183 292 1184
rect 286 1179 287 1183
rect 291 1179 292 1183
rect 286 1178 292 1179
rect 307 1183 313 1184
rect 307 1179 308 1183
rect 312 1182 313 1183
rect 346 1183 352 1184
rect 346 1182 347 1183
rect 312 1180 347 1182
rect 312 1179 313 1180
rect 307 1178 313 1179
rect 346 1179 347 1180
rect 351 1179 352 1183
rect 346 1178 352 1179
rect 366 1183 372 1184
rect 366 1179 367 1183
rect 371 1179 372 1183
rect 366 1178 372 1179
rect 382 1183 393 1184
rect 382 1179 383 1183
rect 387 1179 388 1183
rect 392 1179 393 1183
rect 382 1178 393 1179
rect 446 1183 452 1184
rect 446 1179 447 1183
rect 451 1179 452 1183
rect 446 1178 452 1179
rect 462 1183 473 1184
rect 462 1179 463 1183
rect 467 1179 468 1183
rect 472 1179 473 1183
rect 462 1178 473 1179
rect 526 1183 532 1184
rect 526 1179 527 1183
rect 531 1179 532 1183
rect 526 1178 532 1179
rect 547 1183 553 1184
rect 547 1179 548 1183
rect 552 1179 553 1183
rect 547 1178 553 1179
rect 598 1183 604 1184
rect 598 1179 599 1183
rect 603 1179 604 1183
rect 598 1178 604 1179
rect 619 1183 625 1184
rect 619 1179 620 1183
rect 624 1182 625 1183
rect 642 1183 648 1184
rect 642 1182 643 1183
rect 624 1180 643 1182
rect 624 1179 625 1180
rect 619 1178 625 1179
rect 642 1179 643 1180
rect 647 1179 648 1183
rect 642 1178 648 1179
rect 662 1183 668 1184
rect 662 1179 663 1183
rect 667 1179 668 1183
rect 662 1178 668 1179
rect 683 1183 689 1184
rect 683 1179 684 1183
rect 688 1182 689 1183
rect 714 1183 720 1184
rect 714 1182 715 1183
rect 688 1180 715 1182
rect 688 1179 689 1180
rect 683 1178 689 1179
rect 714 1179 715 1180
rect 719 1179 720 1183
rect 714 1178 720 1179
rect 734 1183 740 1184
rect 734 1179 735 1183
rect 739 1179 740 1183
rect 734 1178 740 1179
rect 755 1183 761 1184
rect 755 1179 756 1183
rect 760 1182 761 1183
rect 786 1183 792 1184
rect 786 1182 787 1183
rect 760 1180 787 1182
rect 760 1179 761 1180
rect 755 1178 761 1179
rect 786 1179 787 1180
rect 791 1179 792 1183
rect 786 1178 792 1179
rect 806 1183 812 1184
rect 806 1179 807 1183
rect 811 1179 812 1183
rect 806 1178 812 1179
rect 827 1183 833 1184
rect 827 1179 828 1183
rect 832 1182 833 1183
rect 858 1183 864 1184
rect 858 1182 859 1183
rect 832 1180 859 1182
rect 832 1179 833 1180
rect 827 1178 833 1179
rect 858 1179 859 1180
rect 863 1179 864 1183
rect 858 1178 864 1179
rect 878 1183 884 1184
rect 878 1179 879 1183
rect 883 1179 884 1183
rect 878 1178 884 1179
rect 886 1183 892 1184
rect 886 1179 887 1183
rect 891 1182 892 1183
rect 899 1183 905 1184
rect 899 1182 900 1183
rect 891 1180 900 1182
rect 891 1179 892 1180
rect 886 1178 892 1179
rect 899 1179 900 1180
rect 904 1179 905 1183
rect 1286 1180 1287 1184
rect 1291 1180 1292 1184
rect 1564 1182 1566 1188
rect 1570 1187 1571 1191
rect 1576 1187 1577 1191
rect 1627 1189 1628 1193
rect 1632 1189 1633 1193
rect 1627 1188 1633 1189
rect 1682 1191 1689 1192
rect 1570 1186 1577 1187
rect 1682 1187 1683 1191
rect 1688 1187 1689 1191
rect 1682 1186 1689 1187
rect 1738 1191 1745 1192
rect 1738 1187 1739 1191
rect 1744 1187 1745 1191
rect 1738 1186 1745 1187
rect 1794 1191 1801 1192
rect 1794 1187 1795 1191
rect 1800 1187 1801 1191
rect 1794 1186 1801 1187
rect 1850 1191 1857 1192
rect 1850 1187 1851 1191
rect 1856 1187 1857 1191
rect 1850 1186 1857 1187
rect 1906 1191 1913 1192
rect 1906 1187 1907 1191
rect 1912 1187 1913 1191
rect 1906 1186 1913 1187
rect 1962 1191 1969 1192
rect 1962 1187 1963 1191
rect 1968 1187 1969 1191
rect 1962 1186 1969 1187
rect 2026 1191 2033 1192
rect 2026 1187 2027 1191
rect 2032 1187 2033 1191
rect 2026 1186 2033 1187
rect 2099 1191 2105 1192
rect 2099 1187 2100 1191
rect 2104 1190 2105 1191
rect 2110 1191 2116 1192
rect 2110 1190 2111 1191
rect 2104 1188 2111 1190
rect 2104 1187 2105 1188
rect 2099 1186 2105 1187
rect 2110 1187 2111 1188
rect 2115 1187 2116 1191
rect 2110 1186 2116 1187
rect 2178 1191 2185 1192
rect 2178 1187 2179 1191
rect 2184 1187 2185 1191
rect 2178 1186 2185 1187
rect 2266 1191 2273 1192
rect 2266 1187 2267 1191
rect 2272 1187 2273 1191
rect 2266 1186 2273 1187
rect 2363 1191 2369 1192
rect 2363 1187 2364 1191
rect 2368 1190 2369 1191
rect 2435 1191 2441 1192
rect 2368 1188 2430 1190
rect 2368 1187 2369 1188
rect 2363 1186 2369 1187
rect 1806 1183 1812 1184
rect 1806 1182 1807 1183
rect 1564 1180 1807 1182
rect 1286 1179 1292 1180
rect 1806 1179 1807 1180
rect 1811 1179 1812 1183
rect 2428 1182 2430 1188
rect 2435 1187 2436 1191
rect 2440 1190 2441 1191
rect 2470 1191 2476 1192
rect 2470 1190 2471 1191
rect 2440 1188 2471 1190
rect 2440 1187 2441 1188
rect 2435 1186 2441 1187
rect 2470 1187 2471 1188
rect 2475 1187 2476 1191
rect 2470 1186 2476 1187
rect 2474 1183 2480 1184
rect 2474 1182 2475 1183
rect 2428 1180 2475 1182
rect 899 1178 905 1179
rect 1806 1178 1812 1179
rect 2474 1179 2475 1180
rect 2479 1179 2480 1183
rect 2474 1178 2480 1179
rect 398 1171 404 1172
rect 398 1170 399 1171
rect 132 1168 399 1170
rect 132 1166 134 1168
rect 398 1167 399 1168
rect 403 1167 404 1171
rect 549 1170 551 1178
rect 1547 1175 1553 1176
rect 1547 1171 1548 1175
rect 1552 1174 1553 1175
rect 1598 1175 1604 1176
rect 1552 1172 1594 1174
rect 1552 1171 1553 1172
rect 1547 1170 1553 1171
rect 398 1166 404 1167
rect 428 1168 551 1170
rect 428 1166 430 1168
rect 1592 1166 1594 1172
rect 1598 1171 1599 1175
rect 1603 1174 1604 1175
rect 1611 1175 1617 1176
rect 1611 1174 1612 1175
rect 1603 1172 1612 1174
rect 1603 1171 1604 1172
rect 1598 1170 1604 1171
rect 1611 1171 1612 1172
rect 1616 1171 1617 1175
rect 1611 1170 1617 1171
rect 1654 1175 1660 1176
rect 1654 1171 1655 1175
rect 1659 1174 1660 1175
rect 1683 1175 1689 1176
rect 1683 1174 1684 1175
rect 1659 1172 1684 1174
rect 1659 1171 1660 1172
rect 1654 1170 1660 1171
rect 1683 1171 1684 1172
rect 1688 1171 1689 1175
rect 1683 1170 1689 1171
rect 1726 1175 1732 1176
rect 1726 1171 1727 1175
rect 1731 1174 1732 1175
rect 1771 1175 1777 1176
rect 1771 1174 1772 1175
rect 1731 1172 1772 1174
rect 1731 1171 1732 1172
rect 1726 1170 1732 1171
rect 1771 1171 1772 1172
rect 1776 1171 1777 1175
rect 1771 1170 1777 1171
rect 1883 1175 1889 1176
rect 1883 1171 1884 1175
rect 1888 1174 1889 1175
rect 2011 1175 2017 1176
rect 1888 1172 2001 1174
rect 1888 1171 1889 1172
rect 1883 1170 1889 1171
rect 1782 1167 1788 1168
rect 1782 1166 1783 1167
rect 131 1165 137 1166
rect 131 1161 132 1165
rect 136 1161 137 1165
rect 427 1165 433 1166
rect 131 1160 137 1161
rect 186 1163 193 1164
rect 186 1159 187 1163
rect 192 1159 193 1163
rect 186 1158 193 1159
rect 266 1163 273 1164
rect 266 1159 267 1163
rect 272 1159 273 1163
rect 266 1158 273 1159
rect 346 1163 353 1164
rect 346 1159 347 1163
rect 352 1159 353 1163
rect 427 1161 428 1165
rect 432 1161 433 1165
rect 1592 1164 1783 1166
rect 427 1160 433 1161
rect 494 1163 500 1164
rect 346 1158 353 1159
rect 494 1159 495 1163
rect 499 1162 500 1163
rect 507 1163 513 1164
rect 507 1162 508 1163
rect 499 1160 508 1162
rect 499 1159 500 1160
rect 494 1158 500 1159
rect 507 1159 508 1160
rect 512 1159 513 1163
rect 507 1158 513 1159
rect 579 1163 585 1164
rect 579 1159 580 1163
rect 584 1162 585 1163
rect 630 1163 636 1164
rect 630 1162 631 1163
rect 584 1160 631 1162
rect 584 1159 585 1160
rect 579 1158 585 1159
rect 630 1159 631 1160
rect 635 1159 636 1163
rect 630 1158 636 1159
rect 642 1163 649 1164
rect 642 1159 643 1163
rect 648 1159 649 1163
rect 642 1158 649 1159
rect 714 1163 721 1164
rect 714 1159 715 1163
rect 720 1159 721 1163
rect 714 1158 721 1159
rect 786 1163 793 1164
rect 786 1159 787 1163
rect 792 1159 793 1163
rect 786 1158 793 1159
rect 858 1163 865 1164
rect 858 1159 859 1163
rect 864 1159 865 1163
rect 1782 1163 1783 1164
rect 1787 1163 1788 1167
rect 1782 1162 1788 1163
rect 1999 1162 2001 1172
rect 2011 1171 2012 1175
rect 2016 1174 2017 1175
rect 2155 1175 2161 1176
rect 2016 1172 2146 1174
rect 2016 1171 2017 1172
rect 2011 1170 2017 1171
rect 2144 1162 2146 1172
rect 2155 1171 2156 1175
rect 2160 1174 2161 1175
rect 2306 1175 2313 1176
rect 2160 1172 2302 1174
rect 2160 1171 2161 1172
rect 2155 1170 2161 1171
rect 2300 1162 2302 1172
rect 2306 1171 2307 1175
rect 2312 1171 2313 1175
rect 2306 1170 2313 1171
rect 2435 1175 2441 1176
rect 2435 1171 2436 1175
rect 2440 1174 2441 1175
rect 2462 1175 2468 1176
rect 2462 1174 2463 1175
rect 2440 1172 2463 1174
rect 2440 1171 2441 1172
rect 2435 1170 2441 1171
rect 2462 1171 2463 1172
rect 2467 1171 2468 1175
rect 2462 1170 2468 1171
rect 1999 1160 2042 1162
rect 2144 1160 2198 1162
rect 2300 1160 2350 1162
rect 858 1158 865 1159
rect 2040 1158 2042 1160
rect 2196 1158 2198 1160
rect 2348 1158 2350 1160
rect 1566 1157 1572 1158
rect 1326 1156 1332 1157
rect 886 1155 892 1156
rect 886 1154 887 1155
rect 636 1152 887 1154
rect 636 1150 638 1152
rect 886 1151 887 1152
rect 891 1151 892 1155
rect 1326 1152 1327 1156
rect 1331 1152 1332 1156
rect 1566 1153 1567 1157
rect 1571 1153 1572 1157
rect 1630 1157 1636 1158
rect 1566 1152 1572 1153
rect 1587 1155 1593 1156
rect 1326 1151 1332 1152
rect 1587 1151 1588 1155
rect 1592 1154 1593 1155
rect 1598 1155 1604 1156
rect 1598 1154 1599 1155
rect 1592 1152 1599 1154
rect 1592 1151 1593 1152
rect 886 1150 892 1151
rect 1587 1150 1593 1151
rect 1598 1151 1599 1152
rect 1603 1151 1604 1155
rect 1630 1153 1631 1157
rect 1635 1153 1636 1157
rect 1702 1157 1708 1158
rect 1630 1152 1636 1153
rect 1651 1155 1660 1156
rect 1598 1150 1604 1151
rect 1651 1151 1652 1155
rect 1659 1151 1660 1155
rect 1702 1153 1703 1157
rect 1707 1153 1708 1157
rect 1790 1157 1796 1158
rect 1702 1152 1708 1153
rect 1723 1155 1732 1156
rect 1651 1150 1660 1151
rect 1723 1151 1724 1155
rect 1731 1151 1732 1155
rect 1790 1153 1791 1157
rect 1795 1153 1796 1157
rect 1902 1157 1908 1158
rect 1790 1152 1796 1153
rect 1806 1155 1817 1156
rect 1723 1150 1732 1151
rect 1806 1151 1807 1155
rect 1811 1151 1812 1155
rect 1816 1151 1817 1155
rect 1902 1153 1903 1157
rect 1907 1153 1908 1157
rect 2030 1157 2036 1158
rect 1902 1152 1908 1153
rect 1918 1155 1929 1156
rect 1806 1150 1817 1151
rect 1918 1151 1919 1155
rect 1923 1151 1924 1155
rect 1928 1151 1929 1155
rect 2030 1153 2031 1157
rect 2035 1153 2036 1157
rect 2040 1157 2057 1158
rect 2040 1156 2052 1157
rect 2030 1152 2036 1153
rect 2051 1153 2052 1156
rect 2056 1153 2057 1157
rect 2051 1152 2057 1153
rect 2174 1157 2180 1158
rect 2174 1153 2175 1157
rect 2179 1153 2180 1157
rect 2174 1152 2180 1153
rect 2195 1157 2201 1158
rect 2195 1153 2196 1157
rect 2200 1153 2201 1157
rect 2195 1152 2201 1153
rect 2326 1157 2332 1158
rect 2326 1153 2327 1157
rect 2331 1153 2332 1157
rect 2326 1152 2332 1153
rect 2347 1157 2353 1158
rect 2347 1153 2348 1157
rect 2352 1153 2353 1157
rect 2347 1152 2353 1153
rect 2454 1157 2460 1158
rect 2454 1153 2455 1157
rect 2459 1153 2460 1157
rect 2502 1156 2508 1157
rect 2454 1152 2460 1153
rect 2462 1155 2468 1156
rect 1918 1150 1929 1151
rect 2462 1151 2463 1155
rect 2467 1154 2468 1155
rect 2475 1155 2481 1156
rect 2475 1154 2476 1155
rect 2467 1152 2476 1154
rect 2467 1151 2468 1152
rect 2462 1150 2468 1151
rect 2475 1151 2476 1152
rect 2480 1151 2481 1155
rect 2502 1152 2503 1156
rect 2507 1152 2508 1156
rect 2502 1151 2508 1152
rect 2475 1150 2481 1151
rect 635 1149 641 1150
rect 163 1147 169 1148
rect 163 1143 164 1147
rect 168 1146 169 1147
rect 259 1147 265 1148
rect 168 1144 254 1146
rect 168 1143 169 1144
rect 163 1142 169 1143
rect 252 1134 254 1144
rect 259 1143 260 1147
rect 264 1146 265 1147
rect 355 1147 361 1148
rect 264 1144 321 1146
rect 264 1143 265 1144
rect 259 1142 265 1143
rect 319 1134 321 1144
rect 355 1143 356 1147
rect 360 1146 361 1147
rect 382 1147 388 1148
rect 382 1146 383 1147
rect 360 1144 383 1146
rect 360 1143 361 1144
rect 355 1142 361 1143
rect 382 1143 383 1144
rect 387 1143 388 1147
rect 382 1142 388 1143
rect 451 1147 457 1148
rect 451 1143 452 1147
rect 456 1146 457 1147
rect 547 1147 553 1148
rect 456 1144 538 1146
rect 456 1143 457 1144
rect 451 1142 457 1143
rect 536 1134 538 1144
rect 547 1143 548 1147
rect 552 1146 553 1147
rect 578 1147 584 1148
rect 578 1146 579 1147
rect 552 1144 579 1146
rect 552 1143 553 1144
rect 547 1142 553 1143
rect 578 1143 579 1144
rect 583 1143 584 1147
rect 635 1145 636 1149
rect 640 1145 641 1149
rect 635 1144 641 1145
rect 715 1147 721 1148
rect 578 1142 584 1143
rect 715 1143 716 1147
rect 720 1143 721 1147
rect 715 1142 721 1143
rect 758 1147 764 1148
rect 758 1143 759 1147
rect 763 1146 764 1147
rect 787 1147 793 1148
rect 787 1146 788 1147
rect 763 1144 788 1146
rect 763 1143 764 1144
rect 758 1142 764 1143
rect 787 1143 788 1144
rect 792 1143 793 1147
rect 787 1142 793 1143
rect 826 1147 832 1148
rect 826 1143 827 1147
rect 831 1146 832 1147
rect 859 1147 865 1148
rect 859 1146 860 1147
rect 831 1144 860 1146
rect 831 1143 832 1144
rect 826 1142 832 1143
rect 859 1143 860 1144
rect 864 1143 865 1147
rect 859 1142 865 1143
rect 902 1147 908 1148
rect 902 1143 903 1147
rect 907 1146 908 1147
rect 939 1147 945 1148
rect 939 1146 940 1147
rect 907 1144 940 1146
rect 907 1143 908 1144
rect 902 1142 908 1143
rect 939 1143 940 1144
rect 944 1143 945 1147
rect 939 1142 945 1143
rect 982 1147 988 1148
rect 982 1143 983 1147
rect 987 1146 988 1147
rect 1019 1147 1025 1148
rect 1019 1146 1020 1147
rect 987 1144 1020 1146
rect 987 1143 988 1144
rect 982 1142 988 1143
rect 1019 1143 1020 1144
rect 1024 1143 1025 1147
rect 1019 1142 1025 1143
rect 252 1132 302 1134
rect 319 1132 398 1134
rect 536 1132 590 1134
rect 300 1130 302 1132
rect 396 1130 398 1132
rect 588 1130 590 1132
rect 717 1130 719 1142
rect 1326 1139 1332 1140
rect 1326 1135 1327 1139
rect 1331 1135 1332 1139
rect 2502 1139 2508 1140
rect 1326 1134 1332 1135
rect 1550 1136 1556 1137
rect 1550 1132 1551 1136
rect 1555 1132 1556 1136
rect 1550 1131 1556 1132
rect 1614 1136 1620 1137
rect 1614 1132 1615 1136
rect 1619 1132 1620 1136
rect 1614 1131 1620 1132
rect 1686 1136 1692 1137
rect 1686 1132 1687 1136
rect 1691 1132 1692 1136
rect 1686 1131 1692 1132
rect 1774 1136 1780 1137
rect 1774 1132 1775 1136
rect 1779 1132 1780 1136
rect 1774 1131 1780 1132
rect 1886 1136 1892 1137
rect 1886 1132 1887 1136
rect 1891 1132 1892 1136
rect 1886 1131 1892 1132
rect 2014 1136 2020 1137
rect 2014 1132 2015 1136
rect 2019 1132 2020 1136
rect 2014 1131 2020 1132
rect 2158 1136 2164 1137
rect 2158 1132 2159 1136
rect 2163 1132 2164 1136
rect 2158 1131 2164 1132
rect 2310 1136 2316 1137
rect 2310 1132 2311 1136
rect 2315 1132 2316 1136
rect 2310 1131 2316 1132
rect 2438 1136 2444 1137
rect 2438 1132 2439 1136
rect 2443 1132 2444 1136
rect 2502 1135 2503 1139
rect 2507 1135 2508 1139
rect 2502 1134 2508 1135
rect 2438 1131 2444 1132
rect 182 1129 188 1130
rect 110 1128 116 1129
rect 110 1124 111 1128
rect 115 1124 116 1128
rect 182 1125 183 1129
rect 187 1125 188 1129
rect 278 1129 284 1130
rect 182 1124 188 1125
rect 198 1127 209 1128
rect 110 1123 116 1124
rect 198 1123 199 1127
rect 203 1123 204 1127
rect 208 1123 209 1127
rect 278 1125 279 1129
rect 283 1125 284 1129
rect 278 1124 284 1125
rect 299 1129 305 1130
rect 299 1125 300 1129
rect 304 1125 305 1129
rect 299 1124 305 1125
rect 374 1129 380 1130
rect 374 1125 375 1129
rect 379 1125 380 1129
rect 374 1124 380 1125
rect 395 1129 401 1130
rect 395 1125 396 1129
rect 400 1125 401 1129
rect 395 1124 401 1125
rect 470 1129 476 1130
rect 470 1125 471 1129
rect 475 1125 476 1129
rect 566 1129 572 1130
rect 470 1124 476 1125
rect 491 1127 500 1128
rect 198 1122 209 1123
rect 491 1123 492 1127
rect 499 1123 500 1127
rect 566 1125 567 1129
rect 571 1125 572 1129
rect 566 1124 572 1125
rect 587 1129 593 1130
rect 587 1125 588 1129
rect 592 1125 593 1129
rect 587 1124 593 1125
rect 654 1129 660 1130
rect 654 1125 655 1129
rect 659 1125 660 1129
rect 654 1124 660 1125
rect 675 1129 719 1130
rect 675 1125 676 1129
rect 680 1128 719 1129
rect 734 1129 740 1130
rect 680 1125 681 1128
rect 675 1124 681 1125
rect 734 1125 735 1129
rect 739 1125 740 1129
rect 806 1129 812 1130
rect 734 1124 740 1125
rect 755 1127 764 1128
rect 491 1122 500 1123
rect 755 1123 756 1127
rect 763 1123 764 1127
rect 806 1125 807 1129
rect 811 1125 812 1129
rect 878 1129 884 1130
rect 806 1124 812 1125
rect 826 1127 833 1128
rect 755 1122 764 1123
rect 826 1123 827 1127
rect 832 1123 833 1127
rect 878 1125 879 1129
rect 883 1125 884 1129
rect 958 1129 964 1130
rect 878 1124 884 1125
rect 899 1127 908 1128
rect 826 1122 833 1123
rect 899 1123 900 1127
rect 907 1123 908 1127
rect 958 1125 959 1129
rect 963 1125 964 1129
rect 1038 1129 1044 1130
rect 958 1124 964 1125
rect 979 1127 988 1128
rect 899 1122 908 1123
rect 979 1123 980 1127
rect 987 1123 988 1127
rect 1038 1125 1039 1129
rect 1043 1125 1044 1129
rect 1286 1128 1292 1129
rect 1038 1124 1044 1125
rect 1059 1127 1068 1128
rect 979 1122 988 1123
rect 1059 1123 1060 1127
rect 1067 1123 1068 1127
rect 1286 1124 1287 1128
rect 1291 1124 1292 1128
rect 1286 1123 1292 1124
rect 1382 1124 1388 1125
rect 1059 1122 1068 1123
rect 1326 1121 1332 1122
rect 1326 1117 1327 1121
rect 1331 1117 1332 1121
rect 1382 1120 1383 1124
rect 1387 1120 1388 1124
rect 1382 1119 1388 1120
rect 1446 1124 1452 1125
rect 1446 1120 1447 1124
rect 1451 1120 1452 1124
rect 1446 1119 1452 1120
rect 1518 1124 1524 1125
rect 1518 1120 1519 1124
rect 1523 1120 1524 1124
rect 1518 1119 1524 1120
rect 1590 1124 1596 1125
rect 1590 1120 1591 1124
rect 1595 1120 1596 1124
rect 1590 1119 1596 1120
rect 1670 1124 1676 1125
rect 1670 1120 1671 1124
rect 1675 1120 1676 1124
rect 1670 1119 1676 1120
rect 1750 1124 1756 1125
rect 1750 1120 1751 1124
rect 1755 1120 1756 1124
rect 1750 1119 1756 1120
rect 1830 1124 1836 1125
rect 1830 1120 1831 1124
rect 1835 1120 1836 1124
rect 1830 1119 1836 1120
rect 1910 1124 1916 1125
rect 1910 1120 1911 1124
rect 1915 1120 1916 1124
rect 1910 1119 1916 1120
rect 1982 1124 1988 1125
rect 1982 1120 1983 1124
rect 1987 1120 1988 1124
rect 1982 1119 1988 1120
rect 2054 1124 2060 1125
rect 2054 1120 2055 1124
rect 2059 1120 2060 1124
rect 2054 1119 2060 1120
rect 2134 1124 2140 1125
rect 2134 1120 2135 1124
rect 2139 1120 2140 1124
rect 2134 1119 2140 1120
rect 2214 1124 2220 1125
rect 2214 1120 2215 1124
rect 2219 1120 2220 1124
rect 2214 1119 2220 1120
rect 2502 1121 2508 1122
rect 1326 1116 1332 1117
rect 2502 1117 2503 1121
rect 2507 1117 2508 1121
rect 2502 1116 2508 1117
rect 110 1111 116 1112
rect 110 1107 111 1111
rect 115 1107 116 1111
rect 1286 1111 1292 1112
rect 110 1106 116 1107
rect 166 1108 172 1109
rect 166 1104 167 1108
rect 171 1104 172 1108
rect 166 1103 172 1104
rect 262 1108 268 1109
rect 262 1104 263 1108
rect 267 1104 268 1108
rect 262 1103 268 1104
rect 358 1108 364 1109
rect 358 1104 359 1108
rect 363 1104 364 1108
rect 358 1103 364 1104
rect 454 1108 460 1109
rect 454 1104 455 1108
rect 459 1104 460 1108
rect 454 1103 460 1104
rect 550 1108 556 1109
rect 550 1104 551 1108
rect 555 1104 556 1108
rect 550 1103 556 1104
rect 638 1108 644 1109
rect 638 1104 639 1108
rect 643 1104 644 1108
rect 638 1103 644 1104
rect 718 1108 724 1109
rect 718 1104 719 1108
rect 723 1104 724 1108
rect 718 1103 724 1104
rect 790 1108 796 1109
rect 790 1104 791 1108
rect 795 1104 796 1108
rect 790 1103 796 1104
rect 862 1108 868 1109
rect 862 1104 863 1108
rect 867 1104 868 1108
rect 862 1103 868 1104
rect 942 1108 948 1109
rect 942 1104 943 1108
rect 947 1104 948 1108
rect 942 1103 948 1104
rect 1022 1108 1028 1109
rect 1022 1104 1023 1108
rect 1027 1104 1028 1108
rect 1286 1107 1287 1111
rect 1291 1107 1292 1111
rect 1286 1106 1292 1107
rect 1022 1103 1028 1104
rect 1326 1104 1332 1105
rect 2502 1104 2508 1105
rect 1326 1100 1327 1104
rect 1331 1100 1332 1104
rect 1326 1099 1332 1100
rect 1398 1103 1404 1104
rect 1398 1099 1399 1103
rect 1403 1099 1404 1103
rect 1398 1098 1404 1099
rect 1419 1103 1425 1104
rect 1419 1099 1420 1103
rect 1424 1102 1425 1103
rect 1442 1103 1448 1104
rect 1442 1102 1443 1103
rect 1424 1100 1443 1102
rect 1424 1099 1425 1100
rect 1419 1098 1425 1099
rect 1442 1099 1443 1100
rect 1447 1099 1448 1103
rect 1442 1098 1448 1099
rect 1462 1103 1468 1104
rect 1462 1099 1463 1103
rect 1467 1099 1468 1103
rect 1462 1098 1468 1099
rect 1483 1103 1489 1104
rect 1483 1099 1484 1103
rect 1488 1102 1489 1103
rect 1514 1103 1520 1104
rect 1514 1102 1515 1103
rect 1488 1100 1515 1102
rect 1488 1099 1489 1100
rect 1483 1098 1489 1099
rect 1514 1099 1515 1100
rect 1519 1099 1520 1103
rect 1514 1098 1520 1099
rect 1534 1103 1540 1104
rect 1534 1099 1535 1103
rect 1539 1099 1540 1103
rect 1534 1098 1540 1099
rect 1555 1103 1561 1104
rect 1555 1099 1556 1103
rect 1560 1102 1561 1103
rect 1586 1103 1592 1104
rect 1586 1102 1587 1103
rect 1560 1100 1587 1102
rect 1560 1099 1561 1100
rect 1555 1098 1561 1099
rect 1586 1099 1587 1100
rect 1591 1099 1592 1103
rect 1586 1098 1592 1099
rect 1606 1103 1612 1104
rect 1606 1099 1607 1103
rect 1611 1099 1612 1103
rect 1606 1098 1612 1099
rect 1627 1103 1633 1104
rect 1627 1099 1628 1103
rect 1632 1102 1633 1103
rect 1666 1103 1672 1104
rect 1666 1102 1667 1103
rect 1632 1100 1667 1102
rect 1632 1099 1633 1100
rect 1627 1098 1633 1099
rect 1666 1099 1667 1100
rect 1671 1099 1672 1103
rect 1666 1098 1672 1099
rect 1686 1103 1692 1104
rect 1686 1099 1687 1103
rect 1691 1099 1692 1103
rect 1686 1098 1692 1099
rect 1707 1103 1713 1104
rect 1707 1099 1708 1103
rect 1712 1102 1713 1103
rect 1746 1103 1752 1104
rect 1746 1102 1747 1103
rect 1712 1100 1747 1102
rect 1712 1099 1713 1100
rect 1707 1098 1713 1099
rect 1746 1099 1747 1100
rect 1751 1099 1752 1103
rect 1746 1098 1752 1099
rect 1766 1103 1772 1104
rect 1766 1099 1767 1103
rect 1771 1099 1772 1103
rect 1766 1098 1772 1099
rect 1782 1103 1793 1104
rect 1782 1099 1783 1103
rect 1787 1099 1788 1103
rect 1792 1099 1793 1103
rect 1782 1098 1793 1099
rect 1846 1103 1852 1104
rect 1846 1099 1847 1103
rect 1851 1099 1852 1103
rect 1846 1098 1852 1099
rect 1867 1103 1873 1104
rect 1867 1099 1868 1103
rect 1872 1102 1873 1103
rect 1906 1103 1912 1104
rect 1906 1102 1907 1103
rect 1872 1100 1907 1102
rect 1872 1099 1873 1100
rect 1867 1098 1873 1099
rect 1906 1099 1907 1100
rect 1911 1099 1912 1103
rect 1906 1098 1912 1099
rect 1926 1103 1932 1104
rect 1926 1099 1927 1103
rect 1931 1099 1932 1103
rect 1926 1098 1932 1099
rect 1947 1103 1953 1104
rect 1947 1099 1948 1103
rect 1952 1102 1953 1103
rect 1978 1103 1984 1104
rect 1978 1102 1979 1103
rect 1952 1100 1979 1102
rect 1952 1099 1953 1100
rect 1947 1098 1953 1099
rect 1978 1099 1979 1100
rect 1983 1099 1984 1103
rect 1978 1098 1984 1099
rect 1998 1103 2004 1104
rect 1998 1099 1999 1103
rect 2003 1099 2004 1103
rect 1998 1098 2004 1099
rect 2019 1103 2025 1104
rect 2019 1099 2020 1103
rect 2024 1102 2025 1103
rect 2050 1103 2056 1104
rect 2050 1102 2051 1103
rect 2024 1100 2051 1102
rect 2024 1099 2025 1100
rect 2019 1098 2025 1099
rect 2050 1099 2051 1100
rect 2055 1099 2056 1103
rect 2050 1098 2056 1099
rect 2070 1103 2076 1104
rect 2070 1099 2071 1103
rect 2075 1099 2076 1103
rect 2070 1098 2076 1099
rect 2091 1103 2097 1104
rect 2091 1099 2092 1103
rect 2096 1102 2097 1103
rect 2130 1103 2136 1104
rect 2130 1102 2131 1103
rect 2096 1100 2131 1102
rect 2096 1099 2097 1100
rect 2091 1098 2097 1099
rect 2130 1099 2131 1100
rect 2135 1099 2136 1103
rect 2130 1098 2136 1099
rect 2150 1103 2156 1104
rect 2150 1099 2151 1103
rect 2155 1099 2156 1103
rect 2150 1098 2156 1099
rect 2171 1103 2177 1104
rect 2171 1099 2172 1103
rect 2176 1102 2177 1103
rect 2210 1103 2216 1104
rect 2210 1102 2211 1103
rect 2176 1100 2211 1102
rect 2176 1099 2177 1100
rect 2171 1098 2177 1099
rect 2210 1099 2211 1100
rect 2215 1099 2216 1103
rect 2210 1098 2216 1099
rect 2230 1103 2236 1104
rect 2230 1099 2231 1103
rect 2235 1099 2236 1103
rect 2230 1098 2236 1099
rect 2238 1103 2244 1104
rect 2238 1099 2239 1103
rect 2243 1102 2244 1103
rect 2251 1103 2257 1104
rect 2251 1102 2252 1103
rect 2243 1100 2252 1102
rect 2243 1099 2244 1100
rect 2238 1098 2244 1099
rect 2251 1099 2252 1100
rect 2256 1099 2257 1103
rect 2502 1100 2503 1104
rect 2507 1100 2508 1104
rect 2502 1099 2508 1100
rect 2251 1098 2257 1099
rect 1918 1091 1924 1092
rect 1918 1090 1919 1091
rect 206 1088 212 1089
rect 110 1085 116 1086
rect 110 1081 111 1085
rect 115 1081 116 1085
rect 206 1084 207 1088
rect 211 1084 212 1088
rect 206 1083 212 1084
rect 278 1088 284 1089
rect 278 1084 279 1088
rect 283 1084 284 1088
rect 278 1083 284 1084
rect 358 1088 364 1089
rect 358 1084 359 1088
rect 363 1084 364 1088
rect 358 1083 364 1084
rect 446 1088 452 1089
rect 446 1084 447 1088
rect 451 1084 452 1088
rect 446 1083 452 1084
rect 542 1088 548 1089
rect 542 1084 543 1088
rect 547 1084 548 1088
rect 542 1083 548 1084
rect 638 1088 644 1089
rect 638 1084 639 1088
rect 643 1084 644 1088
rect 638 1083 644 1084
rect 726 1088 732 1089
rect 726 1084 727 1088
rect 731 1084 732 1088
rect 726 1083 732 1084
rect 814 1088 820 1089
rect 814 1084 815 1088
rect 819 1084 820 1088
rect 814 1083 820 1084
rect 894 1088 900 1089
rect 894 1084 895 1088
rect 899 1084 900 1088
rect 894 1083 900 1084
rect 974 1088 980 1089
rect 974 1084 975 1088
rect 979 1084 980 1088
rect 974 1083 980 1084
rect 1054 1088 1060 1089
rect 1054 1084 1055 1088
rect 1059 1084 1060 1088
rect 1054 1083 1060 1084
rect 1142 1088 1148 1089
rect 1142 1084 1143 1088
rect 1147 1084 1148 1088
rect 1828 1088 1919 1090
rect 1828 1086 1830 1088
rect 1918 1087 1919 1088
rect 1923 1087 1924 1091
rect 1918 1086 1924 1087
rect 1142 1083 1148 1084
rect 1286 1085 1292 1086
rect 110 1080 116 1081
rect 1286 1081 1287 1085
rect 1291 1081 1292 1085
rect 1827 1085 1833 1086
rect 1286 1080 1292 1081
rect 1379 1083 1385 1084
rect 1379 1079 1380 1083
rect 1384 1082 1385 1083
rect 1442 1083 1449 1084
rect 1384 1080 1438 1082
rect 1384 1079 1385 1080
rect 1379 1078 1385 1079
rect 1436 1074 1438 1080
rect 1442 1079 1443 1083
rect 1448 1079 1449 1083
rect 1442 1078 1449 1079
rect 1514 1083 1521 1084
rect 1514 1079 1515 1083
rect 1520 1079 1521 1083
rect 1514 1078 1521 1079
rect 1586 1083 1593 1084
rect 1586 1079 1587 1083
rect 1592 1079 1593 1083
rect 1586 1078 1593 1079
rect 1666 1083 1673 1084
rect 1666 1079 1667 1083
rect 1672 1079 1673 1083
rect 1666 1078 1673 1079
rect 1746 1083 1753 1084
rect 1746 1079 1747 1083
rect 1752 1079 1753 1083
rect 1827 1081 1828 1085
rect 1832 1081 1833 1085
rect 1827 1080 1833 1081
rect 1906 1083 1913 1084
rect 1746 1078 1753 1079
rect 1906 1079 1907 1083
rect 1912 1079 1913 1083
rect 1906 1078 1913 1079
rect 1978 1083 1985 1084
rect 1978 1079 1979 1083
rect 1984 1079 1985 1083
rect 1978 1078 1985 1079
rect 2050 1083 2057 1084
rect 2050 1079 2051 1083
rect 2056 1079 2057 1083
rect 2050 1078 2057 1079
rect 2130 1083 2137 1084
rect 2130 1079 2131 1083
rect 2136 1079 2137 1083
rect 2130 1078 2137 1079
rect 2210 1083 2217 1084
rect 2210 1079 2211 1083
rect 2216 1079 2217 1083
rect 2210 1078 2217 1079
rect 1834 1075 1840 1076
rect 1834 1074 1835 1075
rect 1436 1072 1835 1074
rect 1834 1071 1835 1072
rect 1839 1071 1840 1075
rect 1834 1070 1840 1071
rect 2238 1071 2244 1072
rect 2238 1070 2239 1071
rect 110 1068 116 1069
rect 1286 1068 1292 1069
rect 110 1064 111 1068
rect 115 1064 116 1068
rect 110 1063 116 1064
rect 222 1067 228 1068
rect 222 1063 223 1067
rect 227 1063 228 1067
rect 222 1062 228 1063
rect 243 1067 249 1068
rect 243 1063 244 1067
rect 248 1066 249 1067
rect 274 1067 280 1068
rect 274 1066 275 1067
rect 248 1064 275 1066
rect 248 1063 249 1064
rect 243 1062 249 1063
rect 274 1063 275 1064
rect 279 1063 280 1067
rect 274 1062 280 1063
rect 294 1067 300 1068
rect 294 1063 295 1067
rect 299 1063 300 1067
rect 294 1062 300 1063
rect 315 1067 321 1068
rect 315 1063 316 1067
rect 320 1066 321 1067
rect 354 1067 360 1068
rect 354 1066 355 1067
rect 320 1064 355 1066
rect 320 1063 321 1064
rect 315 1062 321 1063
rect 354 1063 355 1064
rect 359 1063 360 1067
rect 354 1062 360 1063
rect 374 1067 380 1068
rect 374 1063 375 1067
rect 379 1063 380 1067
rect 374 1062 380 1063
rect 395 1067 401 1068
rect 395 1063 396 1067
rect 400 1066 401 1067
rect 442 1067 448 1068
rect 442 1066 443 1067
rect 400 1064 443 1066
rect 400 1063 401 1064
rect 395 1062 401 1063
rect 442 1063 443 1064
rect 447 1063 448 1067
rect 442 1062 448 1063
rect 462 1067 468 1068
rect 462 1063 463 1067
rect 467 1063 468 1067
rect 462 1062 468 1063
rect 470 1067 476 1068
rect 470 1063 471 1067
rect 475 1066 476 1067
rect 483 1067 489 1068
rect 483 1066 484 1067
rect 475 1064 484 1066
rect 475 1063 476 1064
rect 470 1062 476 1063
rect 483 1063 484 1064
rect 488 1063 489 1067
rect 483 1062 489 1063
rect 558 1067 564 1068
rect 558 1063 559 1067
rect 563 1063 564 1067
rect 558 1062 564 1063
rect 578 1067 585 1068
rect 578 1063 579 1067
rect 584 1063 585 1067
rect 578 1062 585 1063
rect 654 1067 660 1068
rect 654 1063 655 1067
rect 659 1063 660 1067
rect 654 1062 660 1063
rect 675 1067 681 1068
rect 675 1063 676 1067
rect 680 1063 681 1067
rect 675 1062 681 1063
rect 742 1067 748 1068
rect 742 1063 743 1067
rect 747 1063 748 1067
rect 742 1062 748 1063
rect 763 1067 769 1068
rect 763 1063 764 1067
rect 768 1066 769 1067
rect 810 1067 816 1068
rect 810 1066 811 1067
rect 768 1064 811 1066
rect 768 1063 769 1064
rect 763 1062 769 1063
rect 810 1063 811 1064
rect 815 1063 816 1067
rect 810 1062 816 1063
rect 830 1067 836 1068
rect 830 1063 831 1067
rect 835 1063 836 1067
rect 830 1062 836 1063
rect 851 1067 857 1068
rect 851 1063 852 1067
rect 856 1066 857 1067
rect 890 1067 896 1068
rect 890 1066 891 1067
rect 856 1064 891 1066
rect 856 1063 857 1064
rect 851 1062 857 1063
rect 890 1063 891 1064
rect 895 1063 896 1067
rect 890 1062 896 1063
rect 910 1067 916 1068
rect 910 1063 911 1067
rect 915 1063 916 1067
rect 910 1062 916 1063
rect 931 1067 937 1068
rect 931 1063 932 1067
rect 936 1066 937 1067
rect 970 1067 976 1068
rect 970 1066 971 1067
rect 936 1064 971 1066
rect 936 1063 937 1064
rect 931 1062 937 1063
rect 970 1063 971 1064
rect 975 1063 976 1067
rect 970 1062 976 1063
rect 990 1067 996 1068
rect 990 1063 991 1067
rect 995 1063 996 1067
rect 990 1062 996 1063
rect 1011 1067 1017 1068
rect 1011 1063 1012 1067
rect 1016 1066 1017 1067
rect 1050 1067 1056 1068
rect 1050 1066 1051 1067
rect 1016 1064 1051 1066
rect 1016 1063 1017 1064
rect 1011 1062 1017 1063
rect 1050 1063 1051 1064
rect 1055 1063 1056 1067
rect 1050 1062 1056 1063
rect 1070 1067 1076 1068
rect 1070 1063 1071 1067
rect 1075 1063 1076 1067
rect 1070 1062 1076 1063
rect 1091 1067 1097 1068
rect 1091 1063 1092 1067
rect 1096 1066 1097 1067
rect 1138 1067 1144 1068
rect 1138 1066 1139 1067
rect 1096 1064 1139 1066
rect 1096 1063 1097 1064
rect 1091 1062 1097 1063
rect 1138 1063 1139 1064
rect 1143 1063 1144 1067
rect 1138 1062 1144 1063
rect 1158 1067 1164 1068
rect 1158 1063 1159 1067
rect 1163 1063 1164 1067
rect 1158 1062 1164 1063
rect 1166 1067 1172 1068
rect 1166 1063 1167 1067
rect 1171 1066 1172 1067
rect 1179 1067 1185 1068
rect 1179 1066 1180 1067
rect 1171 1064 1180 1066
rect 1171 1063 1172 1064
rect 1166 1062 1172 1063
rect 1179 1063 1180 1064
rect 1184 1063 1185 1067
rect 1286 1064 1287 1068
rect 1291 1064 1292 1068
rect 1908 1068 2239 1070
rect 1908 1066 1910 1068
rect 2238 1067 2239 1068
rect 2243 1067 2244 1071
rect 2238 1066 2244 1067
rect 1907 1065 1913 1066
rect 1286 1063 1292 1064
rect 1347 1063 1353 1064
rect 1179 1062 1185 1063
rect 677 1058 679 1062
rect 1347 1059 1348 1063
rect 1352 1062 1353 1063
rect 1390 1063 1396 1064
rect 1352 1060 1386 1062
rect 1352 1059 1353 1060
rect 1347 1058 1353 1059
rect 540 1056 679 1058
rect 540 1050 542 1056
rect 1062 1055 1068 1056
rect 1062 1054 1063 1055
rect 724 1052 1063 1054
rect 724 1050 726 1052
rect 1062 1051 1063 1052
rect 1067 1051 1068 1055
rect 1384 1054 1386 1060
rect 1390 1059 1391 1063
rect 1395 1062 1396 1063
rect 1435 1063 1441 1064
rect 1435 1062 1436 1063
rect 1395 1060 1436 1062
rect 1395 1059 1396 1060
rect 1390 1058 1396 1059
rect 1435 1059 1436 1060
rect 1440 1059 1441 1063
rect 1435 1058 1441 1059
rect 1478 1063 1484 1064
rect 1478 1059 1479 1063
rect 1483 1062 1484 1063
rect 1555 1063 1561 1064
rect 1555 1062 1556 1063
rect 1483 1060 1556 1062
rect 1483 1059 1484 1060
rect 1478 1058 1484 1059
rect 1555 1059 1556 1060
rect 1560 1059 1561 1063
rect 1555 1058 1561 1059
rect 1598 1063 1604 1064
rect 1598 1059 1599 1063
rect 1603 1062 1604 1063
rect 1675 1063 1681 1064
rect 1675 1062 1676 1063
rect 1603 1060 1676 1062
rect 1603 1059 1604 1060
rect 1598 1058 1604 1059
rect 1675 1059 1676 1060
rect 1680 1059 1681 1063
rect 1675 1058 1681 1059
rect 1718 1063 1724 1064
rect 1718 1059 1719 1063
rect 1723 1062 1724 1063
rect 1795 1063 1801 1064
rect 1795 1062 1796 1063
rect 1723 1060 1796 1062
rect 1723 1059 1724 1060
rect 1718 1058 1724 1059
rect 1795 1059 1796 1060
rect 1800 1059 1801 1063
rect 1907 1061 1908 1065
rect 1912 1061 1913 1065
rect 1907 1060 1913 1061
rect 1950 1063 1956 1064
rect 1795 1058 1801 1059
rect 1950 1059 1951 1063
rect 1955 1062 1956 1063
rect 2019 1063 2025 1064
rect 2019 1062 2020 1063
rect 1955 1060 2020 1062
rect 1955 1059 1956 1060
rect 1950 1058 1956 1059
rect 2019 1059 2020 1060
rect 2024 1059 2025 1063
rect 2019 1058 2025 1059
rect 2062 1063 2068 1064
rect 2062 1059 2063 1063
rect 2067 1062 2068 1063
rect 2131 1063 2137 1064
rect 2131 1062 2132 1063
rect 2067 1060 2132 1062
rect 2067 1059 2068 1060
rect 2062 1058 2068 1059
rect 2131 1059 2132 1060
rect 2136 1059 2137 1063
rect 2131 1058 2137 1059
rect 2174 1063 2180 1064
rect 2174 1059 2175 1063
rect 2179 1062 2180 1063
rect 2235 1063 2241 1064
rect 2235 1062 2236 1063
rect 2179 1060 2236 1062
rect 2179 1059 2180 1060
rect 2174 1058 2180 1059
rect 2235 1059 2236 1060
rect 2240 1059 2241 1063
rect 2235 1058 2241 1059
rect 2278 1063 2284 1064
rect 2278 1059 2279 1063
rect 2283 1062 2284 1063
rect 2347 1063 2353 1064
rect 2347 1062 2348 1063
rect 2283 1060 2348 1062
rect 2283 1059 2284 1060
rect 2278 1058 2284 1059
rect 2347 1059 2348 1060
rect 2352 1059 2353 1063
rect 2347 1058 2353 1059
rect 2435 1063 2441 1064
rect 2435 1059 2436 1063
rect 2440 1062 2441 1063
rect 2462 1063 2468 1064
rect 2462 1062 2463 1063
rect 2440 1060 2463 1062
rect 2440 1059 2441 1060
rect 2435 1058 2441 1059
rect 2462 1059 2463 1060
rect 2467 1059 2468 1063
rect 2462 1058 2468 1059
rect 1710 1055 1716 1056
rect 1710 1054 1711 1055
rect 1384 1052 1711 1054
rect 1062 1050 1068 1051
rect 1710 1051 1711 1052
rect 1715 1051 1716 1055
rect 1710 1050 1716 1051
rect 539 1049 545 1050
rect 198 1047 209 1048
rect 198 1043 199 1047
rect 203 1043 204 1047
rect 208 1043 209 1047
rect 198 1042 209 1043
rect 274 1047 281 1048
rect 274 1043 275 1047
rect 280 1043 281 1047
rect 274 1042 281 1043
rect 354 1047 361 1048
rect 354 1043 355 1047
rect 360 1043 361 1047
rect 354 1042 361 1043
rect 442 1047 449 1048
rect 442 1043 443 1047
rect 448 1043 449 1047
rect 539 1045 540 1049
rect 544 1045 545 1049
rect 723 1049 729 1050
rect 539 1044 545 1045
rect 598 1047 604 1048
rect 442 1042 449 1043
rect 598 1043 599 1047
rect 603 1046 604 1047
rect 635 1047 641 1048
rect 635 1046 636 1047
rect 603 1044 636 1046
rect 603 1043 604 1044
rect 598 1042 604 1043
rect 635 1043 636 1044
rect 640 1043 641 1047
rect 723 1045 724 1049
rect 728 1045 729 1049
rect 723 1044 729 1045
rect 810 1047 817 1048
rect 635 1042 641 1043
rect 810 1043 811 1047
rect 816 1043 817 1047
rect 810 1042 817 1043
rect 890 1047 897 1048
rect 890 1043 891 1047
rect 896 1043 897 1047
rect 890 1042 897 1043
rect 970 1047 977 1048
rect 970 1043 971 1047
rect 976 1043 977 1047
rect 970 1042 977 1043
rect 1050 1047 1057 1048
rect 1050 1043 1051 1047
rect 1056 1043 1057 1047
rect 1050 1042 1057 1043
rect 1138 1047 1145 1048
rect 1138 1043 1139 1047
rect 1144 1043 1145 1047
rect 1366 1045 1372 1046
rect 1138 1042 1145 1043
rect 1326 1044 1332 1045
rect 1326 1040 1327 1044
rect 1331 1040 1332 1044
rect 1366 1041 1367 1045
rect 1371 1041 1372 1045
rect 1454 1045 1460 1046
rect 1366 1040 1372 1041
rect 1387 1043 1396 1044
rect 1326 1039 1332 1040
rect 1387 1039 1388 1043
rect 1395 1039 1396 1043
rect 1454 1041 1455 1045
rect 1459 1041 1460 1045
rect 1574 1045 1580 1046
rect 1454 1040 1460 1041
rect 1475 1043 1484 1044
rect 1387 1038 1396 1039
rect 1475 1039 1476 1043
rect 1483 1039 1484 1043
rect 1574 1041 1575 1045
rect 1579 1041 1580 1045
rect 1694 1045 1700 1046
rect 1574 1040 1580 1041
rect 1595 1043 1604 1044
rect 1475 1038 1484 1039
rect 1595 1039 1596 1043
rect 1603 1039 1604 1043
rect 1694 1041 1695 1045
rect 1699 1041 1700 1045
rect 1814 1045 1820 1046
rect 1694 1040 1700 1041
rect 1715 1043 1724 1044
rect 1595 1038 1604 1039
rect 1715 1039 1716 1043
rect 1723 1039 1724 1043
rect 1814 1041 1815 1045
rect 1819 1041 1820 1045
rect 1926 1045 1932 1046
rect 1814 1040 1820 1041
rect 1834 1043 1841 1044
rect 1715 1038 1724 1039
rect 1834 1039 1835 1043
rect 1840 1039 1841 1043
rect 1926 1041 1927 1045
rect 1931 1041 1932 1045
rect 2038 1045 2044 1046
rect 1926 1040 1932 1041
rect 1947 1043 1956 1044
rect 1834 1038 1841 1039
rect 1947 1039 1948 1043
rect 1955 1039 1956 1043
rect 2038 1041 2039 1045
rect 2043 1041 2044 1045
rect 2150 1045 2156 1046
rect 2038 1040 2044 1041
rect 2059 1043 2068 1044
rect 1947 1038 1956 1039
rect 2059 1039 2060 1043
rect 2067 1039 2068 1043
rect 2150 1041 2151 1045
rect 2155 1041 2156 1045
rect 2254 1045 2260 1046
rect 2150 1040 2156 1041
rect 2171 1043 2180 1044
rect 2059 1038 2068 1039
rect 2171 1039 2172 1043
rect 2179 1039 2180 1043
rect 2254 1041 2255 1045
rect 2259 1041 2260 1045
rect 2366 1045 2372 1046
rect 2254 1040 2260 1041
rect 2275 1043 2284 1044
rect 2171 1038 2180 1039
rect 2275 1039 2276 1043
rect 2283 1039 2284 1043
rect 2366 1041 2367 1045
rect 2371 1041 2372 1045
rect 2454 1045 2460 1046
rect 2366 1040 2372 1041
rect 2374 1043 2380 1044
rect 2275 1038 2284 1039
rect 2374 1039 2375 1043
rect 2379 1042 2380 1043
rect 2387 1043 2393 1044
rect 2387 1042 2388 1043
rect 2379 1040 2388 1042
rect 2379 1039 2380 1040
rect 2374 1038 2380 1039
rect 2387 1039 2388 1040
rect 2392 1039 2393 1043
rect 2454 1041 2455 1045
rect 2459 1041 2460 1045
rect 2502 1044 2508 1045
rect 2454 1040 2460 1041
rect 2462 1043 2468 1044
rect 2387 1038 2393 1039
rect 2462 1039 2463 1043
rect 2467 1042 2468 1043
rect 2475 1043 2481 1044
rect 2475 1042 2476 1043
rect 2467 1040 2476 1042
rect 2467 1039 2468 1040
rect 2462 1038 2468 1039
rect 2475 1039 2476 1040
rect 2480 1039 2481 1043
rect 2502 1040 2503 1044
rect 2507 1040 2508 1044
rect 2502 1039 2508 1040
rect 2475 1038 2481 1039
rect 1166 1035 1172 1036
rect 1166 1034 1167 1035
rect 748 1032 1167 1034
rect 748 1030 750 1032
rect 1166 1031 1167 1032
rect 1171 1031 1172 1035
rect 1166 1030 1172 1031
rect 747 1029 753 1030
rect 275 1027 281 1028
rect 275 1023 276 1027
rect 280 1026 281 1027
rect 363 1027 369 1028
rect 280 1024 321 1026
rect 280 1023 281 1024
rect 275 1022 281 1023
rect 319 1014 321 1024
rect 363 1023 364 1027
rect 368 1026 369 1027
rect 459 1027 465 1028
rect 368 1024 454 1026
rect 368 1023 369 1024
rect 363 1022 369 1023
rect 452 1014 454 1024
rect 459 1023 460 1027
rect 464 1026 465 1027
rect 470 1027 476 1028
rect 470 1026 471 1027
rect 464 1024 471 1026
rect 464 1023 465 1024
rect 459 1022 465 1023
rect 470 1023 471 1024
rect 475 1023 476 1027
rect 470 1022 476 1023
rect 555 1027 561 1028
rect 555 1023 556 1027
rect 560 1026 561 1027
rect 651 1027 657 1028
rect 560 1024 646 1026
rect 560 1023 561 1024
rect 555 1022 561 1023
rect 644 1014 646 1024
rect 651 1023 652 1027
rect 656 1026 657 1027
rect 690 1027 696 1028
rect 690 1026 691 1027
rect 656 1024 691 1026
rect 656 1023 657 1024
rect 651 1022 657 1023
rect 690 1023 691 1024
rect 695 1023 696 1027
rect 747 1025 748 1029
rect 752 1025 753 1029
rect 747 1024 753 1025
rect 790 1027 796 1028
rect 690 1022 696 1023
rect 790 1023 791 1027
rect 795 1026 796 1027
rect 835 1027 841 1028
rect 835 1026 836 1027
rect 795 1024 836 1026
rect 795 1023 796 1024
rect 790 1022 796 1023
rect 835 1023 836 1024
rect 840 1023 841 1027
rect 835 1022 841 1023
rect 878 1027 884 1028
rect 878 1023 879 1027
rect 883 1026 884 1027
rect 923 1027 929 1028
rect 923 1026 924 1027
rect 883 1024 924 1026
rect 883 1023 884 1024
rect 878 1022 884 1023
rect 923 1023 924 1024
rect 928 1023 929 1027
rect 923 1022 929 1023
rect 966 1027 972 1028
rect 966 1023 967 1027
rect 971 1026 972 1027
rect 1003 1027 1009 1028
rect 1003 1026 1004 1027
rect 971 1024 1004 1026
rect 971 1023 972 1024
rect 966 1022 972 1023
rect 1003 1023 1004 1024
rect 1008 1023 1009 1027
rect 1003 1022 1009 1023
rect 1046 1027 1052 1028
rect 1046 1023 1047 1027
rect 1051 1026 1052 1027
rect 1083 1027 1089 1028
rect 1083 1026 1084 1027
rect 1051 1024 1084 1026
rect 1051 1023 1052 1024
rect 1046 1022 1052 1023
rect 1083 1023 1084 1024
rect 1088 1023 1089 1027
rect 1083 1022 1089 1023
rect 1135 1027 1141 1028
rect 1135 1023 1136 1027
rect 1140 1026 1141 1027
rect 1163 1027 1169 1028
rect 1163 1026 1164 1027
rect 1140 1024 1164 1026
rect 1140 1023 1141 1024
rect 1135 1022 1141 1023
rect 1163 1023 1164 1024
rect 1168 1023 1169 1027
rect 1163 1022 1169 1023
rect 1206 1027 1212 1028
rect 1206 1023 1207 1027
rect 1211 1026 1212 1027
rect 1219 1027 1225 1028
rect 1219 1026 1220 1027
rect 1211 1024 1220 1026
rect 1211 1023 1212 1024
rect 1206 1022 1212 1023
rect 1219 1023 1220 1024
rect 1224 1023 1225 1027
rect 1219 1022 1225 1023
rect 1326 1027 1332 1028
rect 1326 1023 1327 1027
rect 1331 1023 1332 1027
rect 2502 1027 2508 1028
rect 1326 1022 1332 1023
rect 1350 1024 1356 1025
rect 1350 1020 1351 1024
rect 1355 1020 1356 1024
rect 1350 1019 1356 1020
rect 1438 1024 1444 1025
rect 1438 1020 1439 1024
rect 1443 1020 1444 1024
rect 1438 1019 1444 1020
rect 1558 1024 1564 1025
rect 1558 1020 1559 1024
rect 1563 1020 1564 1024
rect 1558 1019 1564 1020
rect 1678 1024 1684 1025
rect 1678 1020 1679 1024
rect 1683 1020 1684 1024
rect 1678 1019 1684 1020
rect 1798 1024 1804 1025
rect 1798 1020 1799 1024
rect 1803 1020 1804 1024
rect 1798 1019 1804 1020
rect 1910 1024 1916 1025
rect 1910 1020 1911 1024
rect 1915 1020 1916 1024
rect 1910 1019 1916 1020
rect 2022 1024 2028 1025
rect 2022 1020 2023 1024
rect 2027 1020 2028 1024
rect 2022 1019 2028 1020
rect 2134 1024 2140 1025
rect 2134 1020 2135 1024
rect 2139 1020 2140 1024
rect 2134 1019 2140 1020
rect 2238 1024 2244 1025
rect 2238 1020 2239 1024
rect 2243 1020 2244 1024
rect 2238 1019 2244 1020
rect 2350 1024 2356 1025
rect 2350 1020 2351 1024
rect 2355 1020 2356 1024
rect 2350 1019 2356 1020
rect 2438 1024 2444 1025
rect 2438 1020 2439 1024
rect 2443 1020 2444 1024
rect 2502 1023 2503 1027
rect 2507 1023 2508 1027
rect 2502 1022 2508 1023
rect 2438 1019 2444 1020
rect 1214 1015 1220 1016
rect 1214 1014 1215 1015
rect 319 1012 406 1014
rect 452 1012 502 1014
rect 644 1012 694 1014
rect 404 1010 406 1012
rect 500 1010 502 1012
rect 692 1010 694 1012
rect 1044 1012 1215 1014
rect 1044 1010 1046 1012
rect 1214 1011 1215 1012
rect 1219 1011 1220 1015
rect 1214 1010 1220 1011
rect 294 1009 300 1010
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 294 1005 295 1009
rect 299 1005 300 1009
rect 382 1009 388 1010
rect 294 1004 300 1005
rect 302 1007 308 1008
rect 110 1003 116 1004
rect 302 1003 303 1007
rect 307 1006 308 1007
rect 315 1007 321 1008
rect 315 1006 316 1007
rect 307 1004 316 1006
rect 307 1003 308 1004
rect 302 1002 308 1003
rect 315 1003 316 1004
rect 320 1003 321 1007
rect 382 1005 383 1009
rect 387 1005 388 1009
rect 382 1004 388 1005
rect 403 1009 409 1010
rect 403 1005 404 1009
rect 408 1005 409 1009
rect 403 1004 409 1005
rect 478 1009 484 1010
rect 478 1005 479 1009
rect 483 1005 484 1009
rect 478 1004 484 1005
rect 499 1009 505 1010
rect 499 1005 500 1009
rect 504 1005 505 1009
rect 499 1004 505 1005
rect 574 1009 580 1010
rect 574 1005 575 1009
rect 579 1005 580 1009
rect 670 1009 676 1010
rect 574 1004 580 1005
rect 595 1007 604 1008
rect 315 1002 321 1003
rect 595 1003 596 1007
rect 603 1003 604 1007
rect 670 1005 671 1009
rect 675 1005 676 1009
rect 670 1004 676 1005
rect 691 1009 697 1010
rect 691 1005 692 1009
rect 696 1005 697 1009
rect 691 1004 697 1005
rect 766 1009 772 1010
rect 766 1005 767 1009
rect 771 1005 772 1009
rect 854 1009 860 1010
rect 766 1004 772 1005
rect 787 1007 796 1008
rect 595 1002 604 1003
rect 787 1003 788 1007
rect 795 1003 796 1007
rect 854 1005 855 1009
rect 859 1005 860 1009
rect 942 1009 948 1010
rect 854 1004 860 1005
rect 875 1007 884 1008
rect 787 1002 796 1003
rect 875 1003 876 1007
rect 883 1003 884 1007
rect 942 1005 943 1009
rect 947 1005 948 1009
rect 1022 1009 1028 1010
rect 942 1004 948 1005
rect 963 1007 972 1008
rect 875 1002 884 1003
rect 963 1003 964 1007
rect 971 1003 972 1007
rect 1022 1005 1023 1009
rect 1027 1005 1028 1009
rect 1022 1004 1028 1005
rect 1043 1009 1049 1010
rect 1043 1005 1044 1009
rect 1048 1005 1049 1009
rect 1043 1004 1049 1005
rect 1102 1009 1108 1010
rect 1102 1005 1103 1009
rect 1107 1005 1108 1009
rect 1182 1009 1188 1010
rect 1102 1004 1108 1005
rect 1123 1007 1129 1008
rect 963 1002 972 1003
rect 1123 1003 1124 1007
rect 1128 1006 1129 1007
rect 1135 1007 1141 1008
rect 1135 1006 1136 1007
rect 1128 1004 1136 1006
rect 1128 1003 1129 1004
rect 1123 1002 1129 1003
rect 1135 1003 1136 1004
rect 1140 1003 1141 1007
rect 1182 1005 1183 1009
rect 1187 1005 1188 1009
rect 1238 1009 1244 1010
rect 1182 1004 1188 1005
rect 1203 1007 1212 1008
rect 1135 1002 1141 1003
rect 1203 1003 1204 1007
rect 1211 1003 1212 1007
rect 1238 1005 1239 1009
rect 1243 1005 1244 1009
rect 1286 1008 1292 1009
rect 1238 1004 1244 1005
rect 1259 1007 1265 1008
rect 1203 1002 1212 1003
rect 1259 1003 1260 1007
rect 1264 1006 1265 1007
rect 1278 1007 1284 1008
rect 1278 1006 1279 1007
rect 1264 1004 1279 1006
rect 1264 1003 1265 1004
rect 1259 1002 1265 1003
rect 1278 1003 1279 1004
rect 1283 1003 1284 1007
rect 1286 1004 1287 1008
rect 1291 1004 1292 1008
rect 1350 1008 1356 1009
rect 1286 1003 1292 1004
rect 1326 1005 1332 1006
rect 1278 1002 1284 1003
rect 1326 1001 1327 1005
rect 1331 1001 1332 1005
rect 1350 1004 1351 1008
rect 1355 1004 1356 1008
rect 1350 1003 1356 1004
rect 1510 1008 1516 1009
rect 1510 1004 1511 1008
rect 1515 1004 1516 1008
rect 1510 1003 1516 1004
rect 1678 1008 1684 1009
rect 1678 1004 1679 1008
rect 1683 1004 1684 1008
rect 1678 1003 1684 1004
rect 1822 1008 1828 1009
rect 1822 1004 1823 1008
rect 1827 1004 1828 1008
rect 1822 1003 1828 1004
rect 1950 1008 1956 1009
rect 1950 1004 1951 1008
rect 1955 1004 1956 1008
rect 1950 1003 1956 1004
rect 2070 1008 2076 1009
rect 2070 1004 2071 1008
rect 2075 1004 2076 1008
rect 2070 1003 2076 1004
rect 2174 1008 2180 1009
rect 2174 1004 2175 1008
rect 2179 1004 2180 1008
rect 2174 1003 2180 1004
rect 2270 1008 2276 1009
rect 2270 1004 2271 1008
rect 2275 1004 2276 1008
rect 2270 1003 2276 1004
rect 2366 1008 2372 1009
rect 2366 1004 2367 1008
rect 2371 1004 2372 1008
rect 2366 1003 2372 1004
rect 2438 1008 2444 1009
rect 2438 1004 2439 1008
rect 2443 1004 2444 1008
rect 2438 1003 2444 1004
rect 2502 1005 2508 1006
rect 1326 1000 1332 1001
rect 2502 1001 2503 1005
rect 2507 1001 2508 1005
rect 2502 1000 2508 1001
rect 110 991 116 992
rect 110 987 111 991
rect 115 987 116 991
rect 1286 991 1292 992
rect 110 986 116 987
rect 278 988 284 989
rect 278 984 279 988
rect 283 984 284 988
rect 278 983 284 984
rect 366 988 372 989
rect 366 984 367 988
rect 371 984 372 988
rect 366 983 372 984
rect 462 988 468 989
rect 462 984 463 988
rect 467 984 468 988
rect 462 983 468 984
rect 558 988 564 989
rect 558 984 559 988
rect 563 984 564 988
rect 558 983 564 984
rect 654 988 660 989
rect 654 984 655 988
rect 659 984 660 988
rect 654 983 660 984
rect 750 988 756 989
rect 750 984 751 988
rect 755 984 756 988
rect 750 983 756 984
rect 838 988 844 989
rect 838 984 839 988
rect 843 984 844 988
rect 838 983 844 984
rect 926 988 932 989
rect 926 984 927 988
rect 931 984 932 988
rect 926 983 932 984
rect 1006 988 1012 989
rect 1006 984 1007 988
rect 1011 984 1012 988
rect 1006 983 1012 984
rect 1086 988 1092 989
rect 1086 984 1087 988
rect 1091 984 1092 988
rect 1086 983 1092 984
rect 1166 988 1172 989
rect 1166 984 1167 988
rect 1171 984 1172 988
rect 1166 983 1172 984
rect 1222 988 1228 989
rect 1222 984 1223 988
rect 1227 984 1228 988
rect 1286 987 1287 991
rect 1291 987 1292 991
rect 1286 986 1292 987
rect 1326 988 1332 989
rect 2502 988 2508 989
rect 1222 983 1228 984
rect 1326 984 1327 988
rect 1331 984 1332 988
rect 1326 983 1332 984
rect 1366 987 1372 988
rect 1366 983 1367 987
rect 1371 983 1372 987
rect 1366 982 1372 983
rect 1374 987 1380 988
rect 1374 983 1375 987
rect 1379 986 1380 987
rect 1387 987 1393 988
rect 1387 986 1388 987
rect 1379 984 1388 986
rect 1379 983 1380 984
rect 1374 982 1380 983
rect 1387 983 1388 984
rect 1392 983 1393 987
rect 1387 982 1393 983
rect 1526 987 1532 988
rect 1526 983 1527 987
rect 1531 983 1532 987
rect 1526 982 1532 983
rect 1547 987 1553 988
rect 1547 983 1548 987
rect 1552 986 1553 987
rect 1674 987 1680 988
rect 1674 986 1675 987
rect 1552 984 1675 986
rect 1552 983 1553 984
rect 1547 982 1553 983
rect 1674 983 1675 984
rect 1679 983 1680 987
rect 1674 982 1680 983
rect 1694 987 1700 988
rect 1694 983 1695 987
rect 1699 983 1700 987
rect 1694 982 1700 983
rect 1710 987 1721 988
rect 1710 983 1711 987
rect 1715 983 1716 987
rect 1720 983 1721 987
rect 1710 982 1721 983
rect 1838 987 1844 988
rect 1838 983 1839 987
rect 1843 983 1844 987
rect 1838 982 1844 983
rect 1859 987 1865 988
rect 1859 983 1860 987
rect 1864 986 1865 987
rect 1946 987 1952 988
rect 1946 986 1947 987
rect 1864 984 1947 986
rect 1864 983 1865 984
rect 1859 982 1865 983
rect 1946 983 1947 984
rect 1951 983 1952 987
rect 1946 982 1952 983
rect 1966 987 1972 988
rect 1966 983 1967 987
rect 1971 983 1972 987
rect 1966 982 1972 983
rect 1987 987 1993 988
rect 1987 983 1988 987
rect 1992 986 1993 987
rect 2066 987 2072 988
rect 2066 986 2067 987
rect 1992 984 2067 986
rect 1992 983 1993 984
rect 1987 982 1993 983
rect 2066 983 2067 984
rect 2071 983 2072 987
rect 2066 982 2072 983
rect 2086 987 2092 988
rect 2086 983 2087 987
rect 2091 983 2092 987
rect 2086 982 2092 983
rect 2107 987 2113 988
rect 2107 983 2108 987
rect 2112 986 2113 987
rect 2170 987 2176 988
rect 2170 986 2171 987
rect 2112 984 2171 986
rect 2112 983 2113 984
rect 2107 982 2113 983
rect 2170 983 2171 984
rect 2175 983 2176 987
rect 2170 982 2176 983
rect 2190 987 2196 988
rect 2190 983 2191 987
rect 2195 983 2196 987
rect 2190 982 2196 983
rect 2211 987 2217 988
rect 2211 983 2212 987
rect 2216 986 2217 987
rect 2266 987 2272 988
rect 2266 986 2267 987
rect 2216 984 2267 986
rect 2216 983 2217 984
rect 2211 982 2217 983
rect 2266 983 2267 984
rect 2271 983 2272 987
rect 2266 982 2272 983
rect 2286 987 2292 988
rect 2286 983 2287 987
rect 2291 983 2292 987
rect 2286 982 2292 983
rect 2307 987 2313 988
rect 2307 983 2308 987
rect 2312 986 2313 987
rect 2362 987 2368 988
rect 2362 986 2363 987
rect 2312 984 2363 986
rect 2312 983 2313 984
rect 2307 982 2313 983
rect 2362 983 2363 984
rect 2367 983 2368 987
rect 2362 982 2368 983
rect 2382 987 2388 988
rect 2382 983 2383 987
rect 2387 983 2388 987
rect 2382 982 2388 983
rect 2390 987 2396 988
rect 2390 983 2391 987
rect 2395 986 2396 987
rect 2403 987 2409 988
rect 2403 986 2404 987
rect 2395 984 2404 986
rect 2395 983 2396 984
rect 2390 982 2396 983
rect 2403 983 2404 984
rect 2408 983 2409 987
rect 2403 982 2409 983
rect 2454 987 2460 988
rect 2454 983 2455 987
rect 2459 983 2460 987
rect 2454 982 2460 983
rect 2474 987 2481 988
rect 2474 983 2475 987
rect 2480 983 2481 987
rect 2502 984 2503 988
rect 2507 984 2508 988
rect 2502 983 2508 984
rect 2474 982 2481 983
rect 1278 979 1284 980
rect 270 976 276 977
rect 110 973 116 974
rect 110 969 111 973
rect 115 969 116 973
rect 270 972 271 976
rect 275 972 276 976
rect 270 971 276 972
rect 358 976 364 977
rect 358 972 359 976
rect 363 972 364 976
rect 358 971 364 972
rect 454 976 460 977
rect 454 972 455 976
rect 459 972 460 976
rect 454 971 460 972
rect 550 976 556 977
rect 550 972 551 976
rect 555 972 556 976
rect 550 971 556 972
rect 654 976 660 977
rect 654 972 655 976
rect 659 972 660 976
rect 654 971 660 972
rect 750 976 756 977
rect 750 972 751 976
rect 755 972 756 976
rect 750 971 756 972
rect 838 976 844 977
rect 838 972 839 976
rect 843 972 844 976
rect 838 971 844 972
rect 926 976 932 977
rect 926 972 927 976
rect 931 972 932 976
rect 926 971 932 972
rect 1006 976 1012 977
rect 1006 972 1007 976
rect 1011 972 1012 976
rect 1006 971 1012 972
rect 1086 976 1092 977
rect 1086 972 1087 976
rect 1091 972 1092 976
rect 1086 971 1092 972
rect 1166 976 1172 977
rect 1166 972 1167 976
rect 1171 972 1172 976
rect 1166 971 1172 972
rect 1222 976 1228 977
rect 1222 972 1223 976
rect 1227 972 1228 976
rect 1278 975 1279 979
rect 1283 978 1284 979
rect 1283 976 1510 978
rect 1283 975 1284 976
rect 1278 974 1284 975
rect 1222 971 1228 972
rect 1286 973 1292 974
rect 110 968 116 969
rect 1286 969 1287 973
rect 1291 969 1292 973
rect 1508 970 1510 976
rect 1286 968 1292 969
rect 1507 969 1513 970
rect 1347 967 1353 968
rect 1347 966 1348 967
rect 1261 964 1348 966
rect 1261 958 1263 964
rect 1347 963 1348 964
rect 1352 963 1353 967
rect 1507 965 1508 969
rect 1512 965 1513 969
rect 1507 964 1513 965
rect 1674 967 1681 968
rect 1347 962 1353 963
rect 1674 963 1675 967
rect 1680 963 1681 967
rect 1674 962 1681 963
rect 1819 967 1828 968
rect 1819 963 1820 967
rect 1827 963 1828 967
rect 1819 962 1828 963
rect 1946 967 1953 968
rect 1946 963 1947 967
rect 1952 963 1953 967
rect 1946 962 1953 963
rect 2066 967 2073 968
rect 2066 963 2067 967
rect 2072 963 2073 967
rect 2066 962 2073 963
rect 2170 967 2177 968
rect 2170 963 2171 967
rect 2176 963 2177 967
rect 2170 962 2177 963
rect 2266 967 2273 968
rect 2266 963 2267 967
rect 2272 963 2273 967
rect 2266 962 2273 963
rect 2362 967 2369 968
rect 2362 963 2363 967
rect 2368 963 2369 967
rect 2362 962 2369 963
rect 2435 967 2441 968
rect 2435 963 2436 967
rect 2440 966 2441 967
rect 2446 967 2452 968
rect 2446 966 2447 967
rect 2440 964 2447 966
rect 2440 963 2441 964
rect 2435 962 2441 963
rect 2446 963 2447 964
rect 2451 963 2452 967
rect 2446 962 2452 963
rect 1259 957 1265 958
rect 110 956 116 957
rect 110 952 111 956
rect 115 952 116 956
rect 110 951 116 952
rect 286 955 292 956
rect 286 951 287 955
rect 291 951 292 955
rect 286 950 292 951
rect 307 955 313 956
rect 307 951 308 955
rect 312 954 313 955
rect 354 955 360 956
rect 354 954 355 955
rect 312 952 355 954
rect 312 951 313 952
rect 307 950 313 951
rect 354 951 355 952
rect 359 951 360 955
rect 354 950 360 951
rect 374 955 380 956
rect 374 951 375 955
rect 379 951 380 955
rect 374 950 380 951
rect 395 955 401 956
rect 395 951 396 955
rect 400 954 401 955
rect 450 955 456 956
rect 450 954 451 955
rect 400 952 451 954
rect 400 951 401 952
rect 395 950 401 951
rect 450 951 451 952
rect 455 951 456 955
rect 450 950 456 951
rect 470 955 476 956
rect 470 951 471 955
rect 475 951 476 955
rect 470 950 476 951
rect 478 955 484 956
rect 478 951 479 955
rect 483 954 484 955
rect 491 955 497 956
rect 491 954 492 955
rect 483 952 492 954
rect 483 951 484 952
rect 478 950 484 951
rect 491 951 492 952
rect 496 951 497 955
rect 491 950 497 951
rect 566 955 572 956
rect 566 951 567 955
rect 571 951 572 955
rect 566 950 572 951
rect 587 955 593 956
rect 587 951 588 955
rect 592 954 593 955
rect 650 955 656 956
rect 650 954 651 955
rect 592 952 651 954
rect 592 951 593 952
rect 587 950 593 951
rect 650 951 651 952
rect 655 951 656 955
rect 650 950 656 951
rect 670 955 676 956
rect 670 951 671 955
rect 675 951 676 955
rect 670 950 676 951
rect 690 955 697 956
rect 690 951 691 955
rect 696 951 697 955
rect 690 950 697 951
rect 766 955 772 956
rect 766 951 767 955
rect 771 951 772 955
rect 766 950 772 951
rect 787 955 793 956
rect 787 951 788 955
rect 792 954 793 955
rect 834 955 840 956
rect 834 954 835 955
rect 792 952 835 954
rect 792 951 793 952
rect 787 950 793 951
rect 834 951 835 952
rect 839 951 840 955
rect 834 950 840 951
rect 854 955 860 956
rect 854 951 855 955
rect 859 951 860 955
rect 854 950 860 951
rect 875 955 881 956
rect 875 951 876 955
rect 880 954 881 955
rect 922 955 928 956
rect 922 954 923 955
rect 880 952 923 954
rect 880 951 881 952
rect 875 950 881 951
rect 922 951 923 952
rect 927 951 928 955
rect 922 950 928 951
rect 942 955 948 956
rect 942 951 943 955
rect 947 951 948 955
rect 942 950 948 951
rect 963 955 969 956
rect 963 951 964 955
rect 968 954 969 955
rect 1002 955 1008 956
rect 1002 954 1003 955
rect 968 952 1003 954
rect 968 951 969 952
rect 963 950 969 951
rect 1002 951 1003 952
rect 1007 951 1008 955
rect 1002 950 1008 951
rect 1022 955 1028 956
rect 1022 951 1023 955
rect 1027 951 1028 955
rect 1022 950 1028 951
rect 1043 955 1052 956
rect 1043 951 1044 955
rect 1051 951 1052 955
rect 1043 950 1052 951
rect 1102 955 1108 956
rect 1102 951 1103 955
rect 1107 951 1108 955
rect 1123 955 1129 956
rect 1123 954 1124 955
rect 1102 950 1108 951
rect 1112 952 1124 954
rect 1112 946 1114 952
rect 1123 951 1124 952
rect 1128 951 1129 955
rect 1123 950 1129 951
rect 1182 955 1188 956
rect 1182 951 1183 955
rect 1187 951 1188 955
rect 1203 955 1209 956
rect 1203 954 1204 955
rect 1182 950 1188 951
rect 1192 952 1204 954
rect 748 944 1114 946
rect 748 938 750 944
rect 1192 942 1194 952
rect 1203 951 1204 952
rect 1208 951 1209 955
rect 1203 950 1209 951
rect 1238 955 1244 956
rect 1238 951 1239 955
rect 1243 951 1244 955
rect 1259 953 1260 957
rect 1264 953 1265 957
rect 1259 952 1265 953
rect 1286 956 1292 957
rect 1286 952 1287 956
rect 1291 952 1292 956
rect 1286 951 1292 952
rect 1238 950 1244 951
rect 1084 940 1194 942
rect 1347 943 1353 944
rect 1084 938 1086 940
rect 1347 939 1348 943
rect 1352 942 1353 943
rect 1374 943 1380 944
rect 1374 942 1375 943
rect 1352 940 1375 942
rect 1352 939 1353 940
rect 1347 938 1353 939
rect 1374 939 1375 940
rect 1379 939 1380 943
rect 1374 938 1380 939
rect 1390 943 1396 944
rect 1390 939 1391 943
rect 1395 942 1396 943
rect 1403 943 1409 944
rect 1403 942 1404 943
rect 1395 940 1404 942
rect 1395 939 1396 940
rect 1390 938 1396 939
rect 1403 939 1404 940
rect 1408 939 1409 943
rect 1403 938 1409 939
rect 1446 943 1452 944
rect 1446 939 1447 943
rect 1451 942 1452 943
rect 1483 943 1489 944
rect 1483 942 1484 943
rect 1451 940 1484 942
rect 1451 939 1452 940
rect 1446 938 1452 939
rect 1483 939 1484 940
rect 1488 939 1489 943
rect 1483 938 1489 939
rect 1534 943 1540 944
rect 1534 939 1535 943
rect 1539 942 1540 943
rect 1587 943 1593 944
rect 1587 942 1588 943
rect 1539 940 1588 942
rect 1539 939 1540 940
rect 1534 938 1540 939
rect 1587 939 1588 940
rect 1592 939 1593 943
rect 1587 938 1593 939
rect 1630 943 1636 944
rect 1630 939 1631 943
rect 1635 942 1636 943
rect 1699 943 1705 944
rect 1699 942 1700 943
rect 1635 940 1700 942
rect 1635 939 1636 940
rect 1630 938 1636 939
rect 1699 939 1700 940
rect 1704 939 1705 943
rect 1699 938 1705 939
rect 1742 943 1748 944
rect 1742 939 1743 943
rect 1747 942 1748 943
rect 1811 943 1817 944
rect 1811 942 1812 943
rect 1747 940 1812 942
rect 1747 939 1748 940
rect 1742 938 1748 939
rect 1811 939 1812 940
rect 1816 939 1817 943
rect 1811 938 1817 939
rect 1915 943 1921 944
rect 1915 939 1916 943
rect 1920 942 1921 943
rect 1958 943 1964 944
rect 1920 940 1954 942
rect 1920 939 1921 940
rect 1915 938 1921 939
rect 747 937 753 938
rect 267 935 273 936
rect 267 931 268 935
rect 272 934 273 935
rect 302 935 308 936
rect 302 934 303 935
rect 272 932 303 934
rect 272 931 273 932
rect 267 930 273 931
rect 302 931 303 932
rect 307 931 308 935
rect 302 930 308 931
rect 354 935 361 936
rect 354 931 355 935
rect 360 931 361 935
rect 354 930 361 931
rect 450 935 457 936
rect 450 931 451 935
rect 456 931 457 935
rect 450 930 457 931
rect 462 935 468 936
rect 462 931 463 935
rect 467 934 468 935
rect 547 935 553 936
rect 547 934 548 935
rect 467 932 548 934
rect 467 931 468 932
rect 462 930 468 931
rect 547 931 548 932
rect 552 931 553 935
rect 547 930 553 931
rect 650 935 657 936
rect 650 931 651 935
rect 656 931 657 935
rect 747 933 748 937
rect 752 933 753 937
rect 1083 937 1089 938
rect 747 932 753 933
rect 834 935 841 936
rect 650 930 657 931
rect 834 931 835 935
rect 840 931 841 935
rect 834 930 841 931
rect 922 935 929 936
rect 922 931 923 935
rect 928 931 929 935
rect 922 930 929 931
rect 1002 935 1009 936
rect 1002 931 1003 935
rect 1008 931 1009 935
rect 1083 933 1084 937
rect 1088 933 1089 937
rect 1083 932 1089 933
rect 1163 935 1169 936
rect 1002 930 1009 931
rect 1163 931 1164 935
rect 1168 934 1169 935
rect 1202 935 1208 936
rect 1202 934 1203 935
rect 1168 932 1203 934
rect 1168 931 1169 932
rect 1163 930 1169 931
rect 1202 931 1203 932
rect 1207 931 1208 935
rect 1202 930 1208 931
rect 1214 935 1225 936
rect 1214 931 1215 935
rect 1219 931 1220 935
rect 1224 931 1225 935
rect 1214 930 1225 931
rect 1438 931 1444 932
rect 1438 927 1439 931
rect 1443 930 1444 931
rect 1952 930 1954 940
rect 1958 939 1959 943
rect 1963 942 1964 943
rect 2011 943 2017 944
rect 2011 942 2012 943
rect 1963 940 2012 942
rect 1963 939 1964 940
rect 1958 938 1964 939
rect 2011 939 2012 940
rect 2016 939 2017 943
rect 2011 938 2017 939
rect 2054 943 2060 944
rect 2054 939 2055 943
rect 2059 942 2060 943
rect 2107 943 2113 944
rect 2107 942 2108 943
rect 2059 940 2108 942
rect 2059 939 2060 940
rect 2054 938 2060 939
rect 2107 939 2108 940
rect 2112 939 2113 943
rect 2107 938 2113 939
rect 2195 943 2201 944
rect 2195 939 2196 943
rect 2200 939 2201 943
rect 2195 938 2201 939
rect 2275 943 2281 944
rect 2275 939 2276 943
rect 2280 942 2281 943
rect 2355 943 2361 944
rect 2280 940 2350 942
rect 2280 939 2281 940
rect 2275 938 2281 939
rect 2197 934 2199 938
rect 2197 932 2318 934
rect 1443 928 1854 930
rect 1952 928 2238 930
rect 1443 927 1444 928
rect 1438 926 1444 927
rect 1852 926 1854 928
rect 2236 926 2238 928
rect 2316 926 2318 932
rect 2348 930 2350 940
rect 2355 939 2356 943
rect 2360 942 2361 943
rect 2390 943 2396 944
rect 2390 942 2391 943
rect 2360 940 2391 942
rect 2360 939 2361 940
rect 2355 938 2361 939
rect 2390 939 2391 940
rect 2395 939 2396 943
rect 2390 938 2396 939
rect 2435 943 2441 944
rect 2435 939 2436 943
rect 2440 942 2441 943
rect 2462 943 2468 944
rect 2462 942 2463 943
rect 2440 940 2463 942
rect 2440 939 2441 940
rect 2435 938 2441 939
rect 2462 939 2463 940
rect 2467 939 2468 943
rect 2462 938 2468 939
rect 2348 928 2399 930
rect 2397 926 2399 928
rect 1366 925 1372 926
rect 1326 924 1332 925
rect 478 923 484 924
rect 478 922 479 923
rect 404 920 479 922
rect 404 918 406 920
rect 478 919 479 920
rect 483 919 484 923
rect 1326 920 1327 924
rect 1331 920 1332 924
rect 1366 921 1367 925
rect 1371 921 1372 925
rect 1422 925 1428 926
rect 1366 920 1372 921
rect 1387 923 1396 924
rect 1326 919 1332 920
rect 1387 919 1388 923
rect 1395 919 1396 923
rect 1422 921 1423 925
rect 1427 921 1428 925
rect 1502 925 1508 926
rect 1422 920 1428 921
rect 1443 923 1452 924
rect 478 918 484 919
rect 1387 918 1396 919
rect 1443 919 1444 923
rect 1451 919 1452 923
rect 1502 921 1503 925
rect 1507 921 1508 925
rect 1606 925 1612 926
rect 1502 920 1508 921
rect 1523 923 1529 924
rect 1443 918 1452 919
rect 1523 919 1524 923
rect 1528 922 1529 923
rect 1534 923 1540 924
rect 1534 922 1535 923
rect 1528 920 1535 922
rect 1528 919 1529 920
rect 1523 918 1529 919
rect 1534 919 1535 920
rect 1539 919 1540 923
rect 1606 921 1607 925
rect 1611 921 1612 925
rect 1718 925 1724 926
rect 1606 920 1612 921
rect 1627 923 1636 924
rect 1534 918 1540 919
rect 1627 919 1628 923
rect 1635 919 1636 923
rect 1718 921 1719 925
rect 1723 921 1724 925
rect 1830 925 1836 926
rect 1718 920 1724 921
rect 1739 923 1748 924
rect 1627 918 1636 919
rect 1739 919 1740 923
rect 1747 919 1748 923
rect 1830 921 1831 925
rect 1835 921 1836 925
rect 1830 920 1836 921
rect 1851 925 1857 926
rect 1851 921 1852 925
rect 1856 921 1857 925
rect 1851 920 1857 921
rect 1934 925 1940 926
rect 1934 921 1935 925
rect 1939 921 1940 925
rect 2030 925 2036 926
rect 1934 920 1940 921
rect 1955 923 1964 924
rect 1739 918 1748 919
rect 1955 919 1956 923
rect 1963 919 1964 923
rect 2030 921 2031 925
rect 2035 921 2036 925
rect 2126 925 2132 926
rect 2030 920 2036 921
rect 2051 923 2060 924
rect 1955 918 1964 919
rect 2051 919 2052 923
rect 2059 919 2060 923
rect 2126 921 2127 925
rect 2131 921 2132 925
rect 2214 925 2220 926
rect 2126 920 2132 921
rect 2147 923 2156 924
rect 2051 918 2060 919
rect 2147 919 2148 923
rect 2155 919 2156 923
rect 2214 921 2215 925
rect 2219 921 2220 925
rect 2214 920 2220 921
rect 2235 925 2241 926
rect 2235 921 2236 925
rect 2240 921 2241 925
rect 2235 920 2241 921
rect 2294 925 2300 926
rect 2294 921 2295 925
rect 2299 921 2300 925
rect 2294 920 2300 921
rect 2315 925 2321 926
rect 2315 921 2316 925
rect 2320 921 2321 925
rect 2315 920 2321 921
rect 2374 925 2380 926
rect 2374 921 2375 925
rect 2379 921 2380 925
rect 2374 920 2380 921
rect 2395 925 2401 926
rect 2395 921 2396 925
rect 2400 921 2401 925
rect 2395 920 2401 921
rect 2454 925 2460 926
rect 2454 921 2455 925
rect 2459 921 2460 925
rect 2502 924 2508 925
rect 2454 920 2460 921
rect 2462 923 2468 924
rect 2147 918 2156 919
rect 2462 919 2463 923
rect 2467 922 2468 923
rect 2475 923 2481 924
rect 2475 922 2476 923
rect 2467 920 2476 922
rect 2467 919 2468 920
rect 2462 918 2468 919
rect 2475 919 2476 920
rect 2480 919 2481 923
rect 2502 920 2503 924
rect 2507 920 2508 924
rect 2502 919 2508 920
rect 2475 918 2481 919
rect 403 917 409 918
rect 251 915 257 916
rect 251 911 252 915
rect 256 914 257 915
rect 278 915 284 916
rect 278 914 279 915
rect 256 912 279 914
rect 256 911 257 912
rect 251 910 257 911
rect 278 911 279 912
rect 283 911 284 915
rect 278 910 284 911
rect 294 915 300 916
rect 294 911 295 915
rect 299 914 300 915
rect 323 915 329 916
rect 323 914 324 915
rect 299 912 324 914
rect 299 911 300 912
rect 294 910 300 911
rect 323 911 324 912
rect 328 911 329 915
rect 403 913 404 917
rect 408 913 409 917
rect 403 912 409 913
rect 446 915 452 916
rect 323 910 329 911
rect 446 911 447 915
rect 451 914 452 915
rect 499 915 505 916
rect 499 914 500 915
rect 451 912 500 914
rect 451 911 452 912
rect 446 910 452 911
rect 499 911 500 912
rect 504 911 505 915
rect 499 910 505 911
rect 542 915 548 916
rect 542 911 543 915
rect 547 914 548 915
rect 595 915 601 916
rect 595 914 596 915
rect 547 912 596 914
rect 547 911 548 912
rect 542 910 548 911
rect 595 911 596 912
rect 600 911 601 915
rect 595 910 601 911
rect 638 915 644 916
rect 638 911 639 915
rect 643 914 644 915
rect 691 915 697 916
rect 691 914 692 915
rect 643 912 692 914
rect 643 911 644 912
rect 638 910 644 911
rect 691 911 692 912
rect 696 911 697 915
rect 691 910 697 911
rect 787 915 793 916
rect 787 911 788 915
rect 792 911 793 915
rect 787 910 793 911
rect 830 915 836 916
rect 830 911 831 915
rect 835 914 836 915
rect 883 915 889 916
rect 883 914 884 915
rect 835 912 884 914
rect 835 911 836 912
rect 830 910 836 911
rect 883 911 884 912
rect 888 911 889 915
rect 883 910 889 911
rect 926 915 932 916
rect 926 911 927 915
rect 931 914 932 915
rect 971 915 977 916
rect 971 914 972 915
rect 931 912 972 914
rect 931 911 932 912
rect 926 910 932 911
rect 971 911 972 912
rect 976 911 977 915
rect 971 910 977 911
rect 1014 915 1020 916
rect 1014 911 1015 915
rect 1019 914 1020 915
rect 1067 915 1073 916
rect 1067 914 1068 915
rect 1019 912 1068 914
rect 1019 911 1020 912
rect 1014 910 1020 911
rect 1067 911 1068 912
rect 1072 911 1073 915
rect 1067 910 1073 911
rect 1119 915 1125 916
rect 1119 911 1120 915
rect 1124 914 1125 915
rect 1163 915 1169 916
rect 1163 914 1164 915
rect 1124 912 1164 914
rect 1124 911 1125 912
rect 1119 910 1125 911
rect 1163 911 1164 912
rect 1168 911 1169 915
rect 1163 910 1169 911
rect 789 906 791 910
rect 938 907 944 908
rect 938 906 939 907
rect 789 904 939 906
rect 462 903 468 904
rect 462 902 463 903
rect 364 900 463 902
rect 364 898 366 900
rect 462 899 463 900
rect 467 899 468 903
rect 938 903 939 904
rect 943 903 944 907
rect 938 902 944 903
rect 1326 907 1332 908
rect 1326 903 1327 907
rect 1331 903 1332 907
rect 2502 907 2508 908
rect 1326 902 1332 903
rect 1350 904 1356 905
rect 1350 900 1351 904
rect 1355 900 1356 904
rect 1350 899 1356 900
rect 1406 904 1412 905
rect 1406 900 1407 904
rect 1411 900 1412 904
rect 1406 899 1412 900
rect 1486 904 1492 905
rect 1486 900 1487 904
rect 1491 900 1492 904
rect 1486 899 1492 900
rect 1590 904 1596 905
rect 1590 900 1591 904
rect 1595 900 1596 904
rect 1590 899 1596 900
rect 1702 904 1708 905
rect 1702 900 1703 904
rect 1707 900 1708 904
rect 1702 899 1708 900
rect 1814 904 1820 905
rect 1814 900 1815 904
rect 1819 900 1820 904
rect 1814 899 1820 900
rect 1918 904 1924 905
rect 1918 900 1919 904
rect 1923 900 1924 904
rect 1918 899 1924 900
rect 2014 904 2020 905
rect 2014 900 2015 904
rect 2019 900 2020 904
rect 2014 899 2020 900
rect 2110 904 2116 905
rect 2110 900 2111 904
rect 2115 900 2116 904
rect 2110 899 2116 900
rect 2198 904 2204 905
rect 2198 900 2199 904
rect 2203 900 2204 904
rect 2198 899 2204 900
rect 2278 904 2284 905
rect 2278 900 2279 904
rect 2283 900 2284 904
rect 2278 899 2284 900
rect 2358 904 2364 905
rect 2358 900 2359 904
rect 2363 900 2364 904
rect 2358 899 2364 900
rect 2438 904 2444 905
rect 2438 900 2439 904
rect 2443 900 2444 904
rect 2502 903 2503 907
rect 2507 903 2508 907
rect 2502 902 2508 903
rect 2438 899 2444 900
rect 462 898 468 899
rect 270 897 276 898
rect 110 896 116 897
rect 110 892 111 896
rect 115 892 116 896
rect 270 893 271 897
rect 275 893 276 897
rect 342 897 348 898
rect 270 892 276 893
rect 291 895 300 896
rect 110 891 116 892
rect 291 891 292 895
rect 299 891 300 895
rect 342 893 343 897
rect 347 893 348 897
rect 342 892 348 893
rect 363 897 369 898
rect 363 893 364 897
rect 368 893 369 897
rect 363 892 369 893
rect 422 897 428 898
rect 422 893 423 897
rect 427 893 428 897
rect 518 897 524 898
rect 422 892 428 893
rect 443 895 452 896
rect 291 890 300 891
rect 443 891 444 895
rect 451 891 452 895
rect 518 893 519 897
rect 523 893 524 897
rect 614 897 620 898
rect 518 892 524 893
rect 539 895 548 896
rect 443 890 452 891
rect 539 891 540 895
rect 547 891 548 895
rect 614 893 615 897
rect 619 893 620 897
rect 710 897 716 898
rect 614 892 620 893
rect 635 895 644 896
rect 539 890 548 891
rect 635 891 636 895
rect 643 891 644 895
rect 710 893 711 897
rect 715 893 716 897
rect 806 897 812 898
rect 710 892 716 893
rect 718 895 724 896
rect 635 890 644 891
rect 718 891 719 895
rect 723 894 724 895
rect 731 895 737 896
rect 731 894 732 895
rect 723 892 732 894
rect 723 891 724 892
rect 718 890 724 891
rect 731 891 732 892
rect 736 891 737 895
rect 806 893 807 897
rect 811 893 812 897
rect 902 897 908 898
rect 806 892 812 893
rect 827 895 836 896
rect 731 890 737 891
rect 827 891 828 895
rect 835 891 836 895
rect 902 893 903 897
rect 907 893 908 897
rect 990 897 996 898
rect 902 892 908 893
rect 923 895 932 896
rect 827 890 836 891
rect 923 891 924 895
rect 931 891 932 895
rect 990 893 991 897
rect 995 893 996 897
rect 1086 897 1092 898
rect 990 892 996 893
rect 1011 895 1020 896
rect 923 890 932 891
rect 1011 891 1012 895
rect 1019 891 1020 895
rect 1086 893 1087 897
rect 1091 893 1092 897
rect 1182 897 1188 898
rect 1086 892 1092 893
rect 1107 895 1113 896
rect 1011 890 1020 891
rect 1107 891 1108 895
rect 1112 894 1113 895
rect 1119 895 1125 896
rect 1119 894 1120 895
rect 1112 892 1120 894
rect 1112 891 1113 892
rect 1107 890 1113 891
rect 1119 891 1120 892
rect 1124 891 1125 895
rect 1182 893 1183 897
rect 1187 893 1188 897
rect 1286 896 1292 897
rect 1182 892 1188 893
rect 1202 895 1209 896
rect 1119 890 1125 891
rect 1202 891 1203 895
rect 1208 891 1209 895
rect 1286 892 1287 896
rect 1291 892 1292 896
rect 1286 891 1292 892
rect 1202 890 1209 891
rect 1430 888 1436 889
rect 1326 885 1332 886
rect 1326 881 1327 885
rect 1331 881 1332 885
rect 1430 884 1431 888
rect 1435 884 1436 888
rect 1430 883 1436 884
rect 1486 888 1492 889
rect 1486 884 1487 888
rect 1491 884 1492 888
rect 1486 883 1492 884
rect 1550 888 1556 889
rect 1550 884 1551 888
rect 1555 884 1556 888
rect 1550 883 1556 884
rect 1622 888 1628 889
rect 1622 884 1623 888
rect 1627 884 1628 888
rect 1622 883 1628 884
rect 1702 888 1708 889
rect 1702 884 1703 888
rect 1707 884 1708 888
rect 1702 883 1708 884
rect 1790 888 1796 889
rect 1790 884 1791 888
rect 1795 884 1796 888
rect 1790 883 1796 884
rect 1894 888 1900 889
rect 1894 884 1895 888
rect 1899 884 1900 888
rect 1894 883 1900 884
rect 2014 888 2020 889
rect 2014 884 2015 888
rect 2019 884 2020 888
rect 2014 883 2020 884
rect 2142 888 2148 889
rect 2142 884 2143 888
rect 2147 884 2148 888
rect 2142 883 2148 884
rect 2278 888 2284 889
rect 2278 884 2279 888
rect 2283 884 2284 888
rect 2278 883 2284 884
rect 2422 888 2428 889
rect 2422 884 2423 888
rect 2427 884 2428 888
rect 2422 883 2428 884
rect 2502 885 2508 886
rect 1326 880 1332 881
rect 2502 881 2503 885
rect 2507 881 2508 885
rect 2502 880 2508 881
rect 110 879 116 880
rect 110 875 111 879
rect 115 875 116 879
rect 1286 879 1292 880
rect 110 874 116 875
rect 254 876 260 877
rect 254 872 255 876
rect 259 872 260 876
rect 254 871 260 872
rect 326 876 332 877
rect 326 872 327 876
rect 331 872 332 876
rect 326 871 332 872
rect 406 876 412 877
rect 406 872 407 876
rect 411 872 412 876
rect 406 871 412 872
rect 502 876 508 877
rect 502 872 503 876
rect 507 872 508 876
rect 502 871 508 872
rect 598 876 604 877
rect 598 872 599 876
rect 603 872 604 876
rect 598 871 604 872
rect 694 876 700 877
rect 694 872 695 876
rect 699 872 700 876
rect 694 871 700 872
rect 790 876 796 877
rect 790 872 791 876
rect 795 872 796 876
rect 790 871 796 872
rect 886 876 892 877
rect 886 872 887 876
rect 891 872 892 876
rect 886 871 892 872
rect 974 876 980 877
rect 974 872 975 876
rect 979 872 980 876
rect 974 871 980 872
rect 1070 876 1076 877
rect 1070 872 1071 876
rect 1075 872 1076 876
rect 1070 871 1076 872
rect 1166 876 1172 877
rect 1166 872 1167 876
rect 1171 872 1172 876
rect 1286 875 1287 879
rect 1291 875 1292 879
rect 1286 874 1292 875
rect 1166 871 1172 872
rect 1326 868 1332 869
rect 2502 868 2508 869
rect 1326 864 1327 868
rect 1331 864 1332 868
rect 1326 863 1332 864
rect 1446 867 1452 868
rect 1446 863 1447 867
rect 1451 863 1452 867
rect 1446 862 1452 863
rect 1467 867 1473 868
rect 1467 863 1468 867
rect 1472 866 1473 867
rect 1482 867 1488 868
rect 1482 866 1483 867
rect 1472 864 1483 866
rect 1472 863 1473 864
rect 1467 862 1473 863
rect 1482 863 1483 864
rect 1487 863 1488 867
rect 1482 862 1488 863
rect 1502 867 1508 868
rect 1502 863 1503 867
rect 1507 863 1508 867
rect 1502 862 1508 863
rect 1523 867 1529 868
rect 1523 863 1524 867
rect 1528 866 1529 867
rect 1546 867 1552 868
rect 1546 866 1547 867
rect 1528 864 1547 866
rect 1528 863 1529 864
rect 1523 862 1529 863
rect 1546 863 1547 864
rect 1551 863 1552 867
rect 1546 862 1552 863
rect 1566 867 1572 868
rect 1566 863 1567 867
rect 1571 863 1572 867
rect 1566 862 1572 863
rect 1587 867 1593 868
rect 1587 863 1588 867
rect 1592 866 1593 867
rect 1618 867 1624 868
rect 1618 866 1619 867
rect 1592 864 1619 866
rect 1592 863 1593 864
rect 1587 862 1593 863
rect 1618 863 1619 864
rect 1623 863 1624 867
rect 1618 862 1624 863
rect 1638 867 1644 868
rect 1638 863 1639 867
rect 1643 863 1644 867
rect 1638 862 1644 863
rect 1659 867 1665 868
rect 1659 863 1660 867
rect 1664 866 1665 867
rect 1698 867 1704 868
rect 1698 866 1699 867
rect 1664 864 1699 866
rect 1664 863 1665 864
rect 1659 862 1665 863
rect 1698 863 1699 864
rect 1703 863 1704 867
rect 1698 862 1704 863
rect 1718 867 1724 868
rect 1718 863 1719 867
rect 1723 863 1724 867
rect 1718 862 1724 863
rect 1726 867 1732 868
rect 1726 863 1727 867
rect 1731 866 1732 867
rect 1739 867 1745 868
rect 1739 866 1740 867
rect 1731 864 1740 866
rect 1731 863 1732 864
rect 1726 862 1732 863
rect 1739 863 1740 864
rect 1744 863 1745 867
rect 1739 862 1745 863
rect 1806 867 1812 868
rect 1806 863 1807 867
rect 1811 863 1812 867
rect 1806 862 1812 863
rect 1827 867 1833 868
rect 1827 863 1828 867
rect 1832 866 1833 867
rect 1890 867 1896 868
rect 1890 866 1891 867
rect 1832 864 1891 866
rect 1832 863 1833 864
rect 1827 862 1833 863
rect 1890 863 1891 864
rect 1895 863 1896 867
rect 1890 862 1896 863
rect 1910 867 1916 868
rect 1910 863 1911 867
rect 1915 863 1916 867
rect 1910 862 1916 863
rect 1918 867 1924 868
rect 1918 863 1919 867
rect 1923 866 1924 867
rect 1931 867 1937 868
rect 1931 866 1932 867
rect 1923 864 1932 866
rect 1923 863 1924 864
rect 1918 862 1924 863
rect 1931 863 1932 864
rect 1936 863 1937 867
rect 1931 862 1937 863
rect 2030 867 2036 868
rect 2030 863 2031 867
rect 2035 863 2036 867
rect 2030 862 2036 863
rect 2051 867 2057 868
rect 2051 863 2052 867
rect 2056 863 2057 867
rect 2051 862 2057 863
rect 2158 867 2164 868
rect 2158 863 2159 867
rect 2163 863 2164 867
rect 2158 862 2164 863
rect 2179 867 2185 868
rect 2179 863 2180 867
rect 2184 866 2185 867
rect 2274 867 2280 868
rect 2274 866 2275 867
rect 2184 864 2275 866
rect 2184 863 2185 864
rect 2179 862 2185 863
rect 2274 863 2275 864
rect 2279 863 2280 867
rect 2274 862 2280 863
rect 2294 867 2300 868
rect 2294 863 2295 867
rect 2299 863 2300 867
rect 2315 867 2321 868
rect 2315 866 2316 867
rect 2294 862 2300 863
rect 2304 864 2316 866
rect 246 860 252 861
rect 110 857 116 858
rect 110 853 111 857
rect 115 853 116 857
rect 246 856 247 860
rect 251 856 252 860
rect 246 855 252 856
rect 310 860 316 861
rect 310 856 311 860
rect 315 856 316 860
rect 310 855 316 856
rect 374 860 380 861
rect 374 856 375 860
rect 379 856 380 860
rect 374 855 380 856
rect 438 860 444 861
rect 438 856 439 860
rect 443 856 444 860
rect 438 855 444 856
rect 502 860 508 861
rect 502 856 503 860
rect 507 856 508 860
rect 502 855 508 856
rect 566 860 572 861
rect 566 856 567 860
rect 571 856 572 860
rect 566 855 572 856
rect 630 860 636 861
rect 630 856 631 860
rect 635 856 636 860
rect 630 855 636 856
rect 694 860 700 861
rect 694 856 695 860
rect 699 856 700 860
rect 694 855 700 856
rect 758 860 764 861
rect 758 856 759 860
rect 763 856 764 860
rect 758 855 764 856
rect 830 860 836 861
rect 830 856 831 860
rect 835 856 836 860
rect 830 855 836 856
rect 902 860 908 861
rect 902 856 903 860
rect 907 856 908 860
rect 902 855 908 856
rect 1286 857 1292 858
rect 110 852 116 853
rect 1286 853 1287 857
rect 1291 853 1292 857
rect 2053 854 2055 862
rect 2304 854 2306 864
rect 2315 863 2316 864
rect 2320 863 2321 867
rect 2315 862 2321 863
rect 2438 867 2444 868
rect 2438 863 2439 867
rect 2443 863 2444 867
rect 2438 862 2444 863
rect 2446 867 2452 868
rect 2446 863 2447 867
rect 2451 866 2452 867
rect 2459 867 2465 868
rect 2459 866 2460 867
rect 2451 864 2460 866
rect 2451 863 2452 864
rect 2446 862 2452 863
rect 2459 863 2460 864
rect 2464 863 2465 867
rect 2502 864 2503 868
rect 2507 864 2508 868
rect 2502 863 2508 864
rect 2459 862 2465 863
rect 1286 852 1292 853
rect 1788 852 2055 854
rect 2064 852 2306 854
rect 1788 850 1790 852
rect 2064 850 2066 852
rect 1787 849 1793 850
rect 1427 847 1433 848
rect 1427 843 1428 847
rect 1432 846 1433 847
rect 1438 847 1444 848
rect 1438 846 1439 847
rect 1432 844 1439 846
rect 1432 843 1433 844
rect 1427 842 1433 843
rect 1438 843 1439 844
rect 1443 843 1444 847
rect 1438 842 1444 843
rect 1482 847 1489 848
rect 1482 843 1483 847
rect 1488 843 1489 847
rect 1482 842 1489 843
rect 1546 847 1553 848
rect 1546 843 1547 847
rect 1552 843 1553 847
rect 1546 842 1553 843
rect 1618 847 1625 848
rect 1618 843 1619 847
rect 1624 843 1625 847
rect 1618 842 1625 843
rect 1698 847 1705 848
rect 1698 843 1699 847
rect 1704 843 1705 847
rect 1787 845 1788 849
rect 1792 845 1793 849
rect 2011 849 2066 850
rect 1787 844 1793 845
rect 1890 847 1897 848
rect 1698 842 1705 843
rect 1890 843 1891 847
rect 1896 843 1897 847
rect 2011 845 2012 849
rect 2016 848 2066 849
rect 2016 845 2017 848
rect 2011 844 2017 845
rect 2139 847 2145 848
rect 1890 842 1897 843
rect 2139 843 2140 847
rect 2144 846 2145 847
rect 2150 847 2156 848
rect 2150 846 2151 847
rect 2144 844 2151 846
rect 2144 843 2145 844
rect 2139 842 2145 843
rect 2150 843 2151 844
rect 2155 843 2156 847
rect 2150 842 2156 843
rect 2274 847 2281 848
rect 2274 843 2275 847
rect 2280 843 2281 847
rect 2274 842 2281 843
rect 2406 847 2412 848
rect 2406 843 2407 847
rect 2411 846 2412 847
rect 2419 847 2425 848
rect 2419 846 2420 847
rect 2411 844 2420 846
rect 2411 843 2412 844
rect 2406 842 2412 843
rect 2419 843 2420 844
rect 2424 843 2425 847
rect 2419 842 2425 843
rect 110 840 116 841
rect 1286 840 1292 841
rect 110 836 111 840
rect 115 836 116 840
rect 110 835 116 836
rect 262 839 268 840
rect 262 835 263 839
rect 267 835 268 839
rect 262 834 268 835
rect 278 839 289 840
rect 278 835 279 839
rect 283 835 284 839
rect 288 835 289 839
rect 278 834 289 835
rect 326 839 332 840
rect 326 835 327 839
rect 331 835 332 839
rect 326 834 332 835
rect 347 839 353 840
rect 347 835 348 839
rect 352 835 353 839
rect 347 834 353 835
rect 390 839 396 840
rect 390 835 391 839
rect 395 835 396 839
rect 390 834 396 835
rect 411 839 417 840
rect 411 835 412 839
rect 416 838 417 839
rect 434 839 440 840
rect 434 838 435 839
rect 416 836 435 838
rect 416 835 417 836
rect 411 834 417 835
rect 434 835 435 836
rect 439 835 440 839
rect 434 834 440 835
rect 454 839 460 840
rect 454 835 455 839
rect 459 835 460 839
rect 454 834 460 835
rect 475 839 481 840
rect 475 835 476 839
rect 480 838 481 839
rect 498 839 504 840
rect 498 838 499 839
rect 480 836 499 838
rect 480 835 481 836
rect 475 834 481 835
rect 498 835 499 836
rect 503 835 504 839
rect 498 834 504 835
rect 518 839 524 840
rect 518 835 519 839
rect 523 835 524 839
rect 518 834 524 835
rect 539 839 545 840
rect 539 835 540 839
rect 544 838 545 839
rect 562 839 568 840
rect 562 838 563 839
rect 544 836 563 838
rect 544 835 545 836
rect 539 834 545 835
rect 562 835 563 836
rect 567 835 568 839
rect 562 834 568 835
rect 582 839 588 840
rect 582 835 583 839
rect 587 835 588 839
rect 582 834 588 835
rect 590 839 596 840
rect 590 835 591 839
rect 595 838 596 839
rect 603 839 609 840
rect 603 838 604 839
rect 595 836 604 838
rect 595 835 596 836
rect 590 834 596 835
rect 603 835 604 836
rect 608 835 609 839
rect 603 834 609 835
rect 646 839 652 840
rect 646 835 647 839
rect 651 835 652 839
rect 646 834 652 835
rect 667 839 673 840
rect 667 835 668 839
rect 672 838 673 839
rect 690 839 696 840
rect 690 838 691 839
rect 672 836 691 838
rect 672 835 673 836
rect 667 834 673 835
rect 690 835 691 836
rect 695 835 696 839
rect 690 834 696 835
rect 710 839 716 840
rect 710 835 711 839
rect 715 835 716 839
rect 710 834 716 835
rect 731 839 737 840
rect 731 835 732 839
rect 736 838 737 839
rect 754 839 760 840
rect 754 838 755 839
rect 736 836 755 838
rect 736 835 737 836
rect 731 834 737 835
rect 754 835 755 836
rect 759 835 760 839
rect 754 834 760 835
rect 774 839 780 840
rect 774 835 775 839
rect 779 835 780 839
rect 774 834 780 835
rect 795 839 801 840
rect 795 835 796 839
rect 800 838 801 839
rect 826 839 832 840
rect 826 838 827 839
rect 800 836 827 838
rect 800 835 801 836
rect 795 834 801 835
rect 826 835 827 836
rect 831 835 832 839
rect 826 834 832 835
rect 846 839 852 840
rect 846 835 847 839
rect 851 835 852 839
rect 846 834 852 835
rect 867 839 873 840
rect 867 835 868 839
rect 872 838 873 839
rect 898 839 904 840
rect 898 838 899 839
rect 872 836 899 838
rect 872 835 873 836
rect 867 834 873 835
rect 898 835 899 836
rect 903 835 904 839
rect 898 834 904 835
rect 918 839 924 840
rect 918 835 919 839
rect 923 835 924 839
rect 918 834 924 835
rect 938 839 945 840
rect 938 835 939 839
rect 944 835 945 839
rect 1286 836 1287 840
rect 1291 836 1292 840
rect 1726 839 1732 840
rect 1726 838 1727 839
rect 1286 835 1292 836
rect 1572 836 1727 838
rect 938 834 945 835
rect 1572 834 1574 836
rect 1726 835 1727 836
rect 1731 835 1732 839
rect 1726 834 1732 835
rect 349 826 351 834
rect 1571 833 1577 834
rect 1571 829 1572 833
rect 1576 829 1577 833
rect 1571 828 1577 829
rect 1614 831 1620 832
rect 718 827 724 828
rect 718 826 719 827
rect 244 824 351 826
rect 372 824 719 826
rect 244 822 246 824
rect 372 822 374 824
rect 718 823 719 824
rect 723 823 724 827
rect 1614 827 1615 831
rect 1619 830 1620 831
rect 1627 831 1633 832
rect 1627 830 1628 831
rect 1619 828 1628 830
rect 1619 827 1620 828
rect 1614 826 1620 827
rect 1627 827 1628 828
rect 1632 827 1633 831
rect 1627 826 1633 827
rect 1670 831 1676 832
rect 1670 827 1671 831
rect 1675 830 1676 831
rect 1683 831 1689 832
rect 1683 830 1684 831
rect 1675 828 1684 830
rect 1675 827 1676 828
rect 1670 826 1676 827
rect 1683 827 1684 828
rect 1688 827 1689 831
rect 1683 826 1689 827
rect 1726 831 1732 832
rect 1726 827 1727 831
rect 1731 830 1732 831
rect 1747 831 1753 832
rect 1747 830 1748 831
rect 1731 828 1748 830
rect 1731 827 1732 828
rect 1726 826 1732 827
rect 1747 827 1748 828
rect 1752 827 1753 831
rect 1747 826 1753 827
rect 1807 831 1813 832
rect 1807 827 1808 831
rect 1812 830 1813 831
rect 1827 831 1833 832
rect 1827 830 1828 831
rect 1812 828 1828 830
rect 1812 827 1813 828
rect 1807 826 1813 827
rect 1827 827 1828 828
rect 1832 827 1833 831
rect 1827 826 1833 827
rect 1907 831 1913 832
rect 1907 827 1908 831
rect 1912 830 1913 831
rect 1918 831 1924 832
rect 1918 830 1919 831
rect 1912 828 1919 830
rect 1912 827 1913 828
rect 1907 826 1913 827
rect 1918 827 1919 828
rect 1923 827 1924 831
rect 1918 826 1924 827
rect 1950 831 1956 832
rect 1950 827 1951 831
rect 1955 830 1956 831
rect 1995 831 2001 832
rect 1995 830 1996 831
rect 1955 828 1996 830
rect 1955 827 1956 828
rect 1950 826 1956 827
rect 1995 827 1996 828
rect 2000 827 2001 831
rect 1995 826 2001 827
rect 2038 831 2044 832
rect 2038 827 2039 831
rect 2043 830 2044 831
rect 2083 831 2089 832
rect 2083 830 2084 831
rect 2043 828 2084 830
rect 2043 827 2044 828
rect 2038 826 2044 827
rect 2083 827 2084 828
rect 2088 827 2089 831
rect 2083 826 2089 827
rect 2171 831 2177 832
rect 2171 827 2172 831
rect 2176 830 2177 831
rect 2214 831 2220 832
rect 2176 828 2210 830
rect 2176 827 2177 828
rect 2171 826 2177 827
rect 718 822 724 823
rect 2208 822 2210 828
rect 2214 827 2215 831
rect 2219 830 2220 831
rect 2267 831 2273 832
rect 2267 830 2268 831
rect 2219 828 2268 830
rect 2219 827 2220 828
rect 2214 826 2220 827
rect 2267 827 2268 828
rect 2272 827 2273 831
rect 2267 826 2273 827
rect 2310 831 2316 832
rect 2310 827 2311 831
rect 2315 830 2316 831
rect 2363 831 2369 832
rect 2363 830 2364 831
rect 2315 828 2364 830
rect 2315 827 2316 828
rect 2310 826 2316 827
rect 2363 827 2364 828
rect 2368 827 2369 831
rect 2363 826 2369 827
rect 2435 831 2441 832
rect 2435 827 2436 831
rect 2440 830 2441 831
rect 2462 831 2468 832
rect 2462 830 2463 831
rect 2440 828 2463 830
rect 2440 827 2441 828
rect 2435 826 2441 827
rect 2462 827 2463 828
rect 2467 827 2468 831
rect 2462 826 2468 827
rect 2374 823 2380 824
rect 2374 822 2375 823
rect 243 821 249 822
rect 243 817 244 821
rect 248 817 249 821
rect 371 821 377 822
rect 243 816 249 817
rect 307 819 313 820
rect 307 815 308 819
rect 312 818 313 819
rect 318 819 324 820
rect 318 818 319 819
rect 312 816 319 818
rect 312 815 313 816
rect 307 814 313 815
rect 318 815 319 816
rect 323 815 324 819
rect 371 817 372 821
rect 376 817 377 821
rect 2208 820 2375 822
rect 371 816 377 817
rect 434 819 441 820
rect 318 814 324 815
rect 434 815 435 819
rect 440 815 441 819
rect 434 814 441 815
rect 498 819 505 820
rect 498 815 499 819
rect 504 815 505 819
rect 498 814 505 815
rect 562 819 569 820
rect 562 815 563 819
rect 568 815 569 819
rect 562 814 569 815
rect 627 819 633 820
rect 627 815 628 819
rect 632 818 633 819
rect 682 819 688 820
rect 682 818 683 819
rect 632 816 683 818
rect 632 815 633 816
rect 627 814 633 815
rect 682 815 683 816
rect 687 815 688 819
rect 682 814 688 815
rect 690 819 697 820
rect 690 815 691 819
rect 696 815 697 819
rect 690 814 697 815
rect 754 819 761 820
rect 754 815 755 819
rect 760 815 761 819
rect 754 814 761 815
rect 826 819 833 820
rect 826 815 827 819
rect 832 815 833 819
rect 826 814 833 815
rect 898 819 905 820
rect 898 815 899 819
rect 904 815 905 819
rect 2374 819 2375 820
rect 2379 819 2380 823
rect 2374 818 2380 819
rect 898 814 905 815
rect 1590 813 1596 814
rect 1326 812 1332 813
rect 590 811 596 812
rect 590 810 591 811
rect 372 808 591 810
rect 372 806 374 808
rect 590 807 591 808
rect 595 807 596 811
rect 1326 808 1327 812
rect 1331 808 1332 812
rect 1590 809 1591 813
rect 1595 809 1596 813
rect 1646 813 1652 814
rect 1590 808 1596 809
rect 1611 811 1620 812
rect 1326 807 1332 808
rect 1611 807 1612 811
rect 1619 807 1620 811
rect 1646 809 1647 813
rect 1651 809 1652 813
rect 1702 813 1708 814
rect 1646 808 1652 809
rect 1667 811 1676 812
rect 590 806 596 807
rect 1611 806 1620 807
rect 1667 807 1668 811
rect 1675 807 1676 811
rect 1702 809 1703 813
rect 1707 809 1708 813
rect 1766 813 1772 814
rect 1702 808 1708 809
rect 1723 811 1732 812
rect 1667 806 1676 807
rect 1723 807 1724 811
rect 1731 807 1732 811
rect 1766 809 1767 813
rect 1771 809 1772 813
rect 1846 813 1852 814
rect 1766 808 1772 809
rect 1787 811 1793 812
rect 1723 806 1732 807
rect 1787 807 1788 811
rect 1792 810 1793 811
rect 1807 811 1813 812
rect 1807 810 1808 811
rect 1792 808 1808 810
rect 1792 807 1793 808
rect 1787 806 1793 807
rect 1807 807 1808 808
rect 1812 807 1813 811
rect 1846 809 1847 813
rect 1851 809 1852 813
rect 1926 813 1932 814
rect 1846 808 1852 809
rect 1854 811 1860 812
rect 1807 806 1813 807
rect 1854 807 1855 811
rect 1859 810 1860 811
rect 1867 811 1873 812
rect 1867 810 1868 811
rect 1859 808 1868 810
rect 1859 807 1860 808
rect 1854 806 1860 807
rect 1867 807 1868 808
rect 1872 807 1873 811
rect 1926 809 1927 813
rect 1931 809 1932 813
rect 2014 813 2020 814
rect 1926 808 1932 809
rect 1947 811 1956 812
rect 1867 806 1873 807
rect 1947 807 1948 811
rect 1955 807 1956 811
rect 2014 809 2015 813
rect 2019 809 2020 813
rect 2102 813 2108 814
rect 2014 808 2020 809
rect 2035 811 2044 812
rect 1947 806 1956 807
rect 2035 807 2036 811
rect 2043 807 2044 811
rect 2102 809 2103 813
rect 2107 809 2108 813
rect 2190 813 2196 814
rect 2102 808 2108 809
rect 2123 811 2132 812
rect 2035 806 2044 807
rect 2123 807 2124 811
rect 2131 807 2132 811
rect 2190 809 2191 813
rect 2195 809 2196 813
rect 2286 813 2292 814
rect 2190 808 2196 809
rect 2211 811 2220 812
rect 2123 806 2132 807
rect 2211 807 2212 811
rect 2219 807 2220 811
rect 2286 809 2287 813
rect 2291 809 2292 813
rect 2382 813 2388 814
rect 2286 808 2292 809
rect 2307 811 2316 812
rect 2211 806 2220 807
rect 2307 807 2308 811
rect 2315 807 2316 811
rect 2382 809 2383 813
rect 2387 809 2388 813
rect 2454 813 2460 814
rect 2382 808 2388 809
rect 2403 811 2412 812
rect 2307 806 2316 807
rect 2403 807 2404 811
rect 2411 807 2412 811
rect 2454 809 2455 813
rect 2459 809 2460 813
rect 2502 812 2508 813
rect 2454 808 2460 809
rect 2470 811 2481 812
rect 2403 806 2412 807
rect 2470 807 2471 811
rect 2475 807 2476 811
rect 2480 807 2481 811
rect 2502 808 2503 812
rect 2507 808 2508 812
rect 2502 807 2508 808
rect 2470 806 2481 807
rect 371 805 377 806
rect 174 803 180 804
rect 174 799 175 803
rect 179 802 180 803
rect 195 803 201 804
rect 195 802 196 803
rect 179 800 196 802
rect 179 799 180 800
rect 174 798 180 799
rect 195 799 196 800
rect 200 799 201 803
rect 195 798 201 799
rect 238 803 244 804
rect 238 799 239 803
rect 243 802 244 803
rect 283 803 289 804
rect 283 802 284 803
rect 243 800 284 802
rect 243 799 244 800
rect 238 798 244 799
rect 283 799 284 800
rect 288 799 289 803
rect 371 801 372 805
rect 376 801 377 805
rect 371 800 377 801
rect 414 803 420 804
rect 283 798 289 799
rect 414 799 415 803
rect 419 802 420 803
rect 459 803 465 804
rect 459 802 460 803
rect 419 800 460 802
rect 419 799 420 800
rect 414 798 420 799
rect 459 799 460 800
rect 464 799 465 803
rect 459 798 465 799
rect 502 803 508 804
rect 502 799 503 803
rect 507 802 508 803
rect 539 803 545 804
rect 539 802 540 803
rect 507 800 540 802
rect 507 799 508 800
rect 502 798 508 799
rect 539 799 540 800
rect 544 799 545 803
rect 539 798 545 799
rect 590 803 596 804
rect 590 799 591 803
rect 595 802 596 803
rect 611 803 617 804
rect 611 802 612 803
rect 595 800 612 802
rect 595 799 596 800
rect 590 798 596 799
rect 611 799 612 800
rect 616 799 617 803
rect 611 798 617 799
rect 654 803 660 804
rect 654 799 655 803
rect 659 802 660 803
rect 683 803 689 804
rect 683 802 684 803
rect 659 800 684 802
rect 659 799 660 800
rect 654 798 660 799
rect 683 799 684 800
rect 688 799 689 803
rect 683 798 689 799
rect 747 803 753 804
rect 747 799 748 803
rect 752 802 753 803
rect 811 803 817 804
rect 752 800 806 802
rect 752 799 753 800
rect 747 798 753 799
rect 682 791 688 792
rect 682 787 683 791
rect 687 790 688 791
rect 804 790 806 800
rect 811 799 812 803
rect 816 802 817 803
rect 875 803 881 804
rect 816 800 870 802
rect 816 799 817 800
rect 811 798 817 799
rect 868 790 870 800
rect 875 799 876 803
rect 880 802 881 803
rect 947 803 953 804
rect 880 800 942 802
rect 880 799 881 800
rect 875 798 881 799
rect 940 790 942 800
rect 947 799 948 803
rect 952 802 953 803
rect 1019 803 1025 804
rect 952 800 1014 802
rect 952 799 953 800
rect 947 798 953 799
rect 1012 790 1014 800
rect 1019 799 1020 803
rect 1024 802 1025 803
rect 1074 803 1080 804
rect 1074 802 1075 803
rect 1024 800 1075 802
rect 1024 799 1025 800
rect 1019 798 1025 799
rect 1074 799 1075 800
rect 1079 799 1080 803
rect 1074 798 1080 799
rect 1326 795 1332 796
rect 1326 791 1327 795
rect 1331 791 1332 795
rect 2502 795 2508 796
rect 1326 790 1332 791
rect 1574 792 1580 793
rect 687 788 726 790
rect 804 788 854 790
rect 868 788 918 790
rect 940 788 990 790
rect 1012 788 1062 790
rect 687 787 688 788
rect 682 786 688 787
rect 724 786 726 788
rect 852 786 854 788
rect 916 786 918 788
rect 988 786 990 788
rect 1060 786 1062 788
rect 1574 788 1575 792
rect 1579 788 1580 792
rect 1574 787 1580 788
rect 1630 792 1636 793
rect 1630 788 1631 792
rect 1635 788 1636 792
rect 1630 787 1636 788
rect 1686 792 1692 793
rect 1686 788 1687 792
rect 1691 788 1692 792
rect 1686 787 1692 788
rect 1750 792 1756 793
rect 1750 788 1751 792
rect 1755 788 1756 792
rect 1750 787 1756 788
rect 1830 792 1836 793
rect 1830 788 1831 792
rect 1835 788 1836 792
rect 1830 787 1836 788
rect 1910 792 1916 793
rect 1910 788 1911 792
rect 1915 788 1916 792
rect 1910 787 1916 788
rect 1998 792 2004 793
rect 1998 788 1999 792
rect 2003 788 2004 792
rect 1998 787 2004 788
rect 2086 792 2092 793
rect 2086 788 2087 792
rect 2091 788 2092 792
rect 2086 787 2092 788
rect 2174 792 2180 793
rect 2174 788 2175 792
rect 2179 788 2180 792
rect 2174 787 2180 788
rect 2270 792 2276 793
rect 2270 788 2271 792
rect 2275 788 2276 792
rect 2270 787 2276 788
rect 2366 792 2372 793
rect 2366 788 2367 792
rect 2371 788 2372 792
rect 2366 787 2372 788
rect 2438 792 2444 793
rect 2438 788 2439 792
rect 2443 788 2444 792
rect 2502 791 2503 795
rect 2507 791 2508 795
rect 2502 790 2508 791
rect 2438 787 2444 788
rect 214 785 220 786
rect 110 784 116 785
rect 110 780 111 784
rect 115 780 116 784
rect 214 781 215 785
rect 219 781 220 785
rect 302 785 308 786
rect 214 780 220 781
rect 235 783 244 784
rect 110 779 116 780
rect 235 779 236 783
rect 243 779 244 783
rect 302 781 303 785
rect 307 781 308 785
rect 390 785 396 786
rect 302 780 308 781
rect 318 783 329 784
rect 235 778 244 779
rect 318 779 319 783
rect 323 779 324 783
rect 328 779 329 783
rect 390 781 391 785
rect 395 781 396 785
rect 478 785 484 786
rect 390 780 396 781
rect 411 783 420 784
rect 318 778 329 779
rect 411 779 412 783
rect 419 779 420 783
rect 478 781 479 785
rect 483 781 484 785
rect 558 785 564 786
rect 478 780 484 781
rect 499 783 508 784
rect 411 778 420 779
rect 499 779 500 783
rect 507 779 508 783
rect 558 781 559 785
rect 563 781 564 785
rect 630 785 636 786
rect 558 780 564 781
rect 579 783 585 784
rect 499 778 508 779
rect 579 779 580 783
rect 584 782 585 783
rect 590 783 596 784
rect 590 782 591 783
rect 584 780 591 782
rect 584 779 585 780
rect 579 778 585 779
rect 590 779 591 780
rect 595 779 596 783
rect 630 781 631 785
rect 635 781 636 785
rect 702 785 708 786
rect 630 780 636 781
rect 651 783 660 784
rect 590 778 596 779
rect 651 779 652 783
rect 659 779 660 783
rect 702 781 703 785
rect 707 781 708 785
rect 702 780 708 781
rect 723 785 729 786
rect 723 781 724 785
rect 728 781 729 785
rect 723 780 729 781
rect 766 785 772 786
rect 766 781 767 785
rect 771 781 772 785
rect 830 785 836 786
rect 766 780 772 781
rect 782 783 793 784
rect 651 778 660 779
rect 782 779 783 783
rect 787 779 788 783
rect 792 779 793 783
rect 830 781 831 785
rect 835 781 836 785
rect 830 780 836 781
rect 851 785 857 786
rect 851 781 852 785
rect 856 781 857 785
rect 851 780 857 781
rect 894 785 900 786
rect 894 781 895 785
rect 899 781 900 785
rect 894 780 900 781
rect 915 785 921 786
rect 915 781 916 785
rect 920 781 921 785
rect 915 780 921 781
rect 966 785 972 786
rect 966 781 967 785
rect 971 781 972 785
rect 966 780 972 781
rect 987 785 993 786
rect 987 781 988 785
rect 992 781 993 785
rect 987 780 993 781
rect 1038 785 1044 786
rect 1038 781 1039 785
rect 1043 781 1044 785
rect 1038 780 1044 781
rect 1059 785 1065 786
rect 1059 781 1060 785
rect 1064 781 1065 785
rect 1059 780 1065 781
rect 1286 784 1292 785
rect 1286 780 1287 784
rect 1291 780 1292 784
rect 1286 779 1292 780
rect 782 778 793 779
rect 1566 776 1572 777
rect 1326 773 1332 774
rect 1326 769 1327 773
rect 1331 769 1332 773
rect 1566 772 1567 776
rect 1571 772 1572 776
rect 1566 771 1572 772
rect 1622 776 1628 777
rect 1622 772 1623 776
rect 1627 772 1628 776
rect 1622 771 1628 772
rect 1686 776 1692 777
rect 1686 772 1687 776
rect 1691 772 1692 776
rect 1686 771 1692 772
rect 1758 776 1764 777
rect 1758 772 1759 776
rect 1763 772 1764 776
rect 1758 771 1764 772
rect 1830 776 1836 777
rect 1830 772 1831 776
rect 1835 772 1836 776
rect 1830 771 1836 772
rect 1918 776 1924 777
rect 1918 772 1919 776
rect 1923 772 1924 776
rect 1918 771 1924 772
rect 2014 776 2020 777
rect 2014 772 2015 776
rect 2019 772 2020 776
rect 2014 771 2020 772
rect 2118 776 2124 777
rect 2118 772 2119 776
rect 2123 772 2124 776
rect 2118 771 2124 772
rect 2230 776 2236 777
rect 2230 772 2231 776
rect 2235 772 2236 776
rect 2230 771 2236 772
rect 2342 776 2348 777
rect 2342 772 2343 776
rect 2347 772 2348 776
rect 2342 771 2348 772
rect 2438 776 2444 777
rect 2438 772 2439 776
rect 2443 772 2444 776
rect 2438 771 2444 772
rect 2502 773 2508 774
rect 1326 768 1332 769
rect 2502 769 2503 773
rect 2507 769 2508 773
rect 2502 768 2508 769
rect 110 767 116 768
rect 110 763 111 767
rect 115 763 116 767
rect 1286 767 1292 768
rect 110 762 116 763
rect 198 764 204 765
rect 198 760 199 764
rect 203 760 204 764
rect 198 759 204 760
rect 286 764 292 765
rect 286 760 287 764
rect 291 760 292 764
rect 286 759 292 760
rect 374 764 380 765
rect 374 760 375 764
rect 379 760 380 764
rect 374 759 380 760
rect 462 764 468 765
rect 462 760 463 764
rect 467 760 468 764
rect 462 759 468 760
rect 542 764 548 765
rect 542 760 543 764
rect 547 760 548 764
rect 542 759 548 760
rect 614 764 620 765
rect 614 760 615 764
rect 619 760 620 764
rect 614 759 620 760
rect 686 764 692 765
rect 686 760 687 764
rect 691 760 692 764
rect 686 759 692 760
rect 750 764 756 765
rect 750 760 751 764
rect 755 760 756 764
rect 750 759 756 760
rect 814 764 820 765
rect 814 760 815 764
rect 819 760 820 764
rect 814 759 820 760
rect 878 764 884 765
rect 878 760 879 764
rect 883 760 884 764
rect 878 759 884 760
rect 950 764 956 765
rect 950 760 951 764
rect 955 760 956 764
rect 950 759 956 760
rect 1022 764 1028 765
rect 1022 760 1023 764
rect 1027 760 1028 764
rect 1286 763 1287 767
rect 1291 763 1292 767
rect 1286 762 1292 763
rect 1022 759 1028 760
rect 1326 756 1332 757
rect 2502 756 2508 757
rect 134 752 140 753
rect 110 749 116 750
rect 110 745 111 749
rect 115 745 116 749
rect 134 748 135 752
rect 139 748 140 752
rect 134 747 140 748
rect 254 752 260 753
rect 254 748 255 752
rect 259 748 260 752
rect 254 747 260 748
rect 390 752 396 753
rect 390 748 391 752
rect 395 748 396 752
rect 390 747 396 748
rect 518 752 524 753
rect 518 748 519 752
rect 523 748 524 752
rect 518 747 524 748
rect 646 752 652 753
rect 646 748 647 752
rect 651 748 652 752
rect 646 747 652 748
rect 774 752 780 753
rect 774 748 775 752
rect 779 748 780 752
rect 774 747 780 748
rect 902 752 908 753
rect 902 748 903 752
rect 907 748 908 752
rect 902 747 908 748
rect 1038 752 1044 753
rect 1038 748 1039 752
rect 1043 748 1044 752
rect 1326 752 1327 756
rect 1331 752 1332 756
rect 1326 751 1332 752
rect 1582 755 1588 756
rect 1582 751 1583 755
rect 1587 751 1588 755
rect 1582 750 1588 751
rect 1603 755 1609 756
rect 1603 751 1604 755
rect 1608 754 1609 755
rect 1618 755 1624 756
rect 1618 754 1619 755
rect 1608 752 1619 754
rect 1608 751 1609 752
rect 1603 750 1609 751
rect 1618 751 1619 752
rect 1623 751 1624 755
rect 1618 750 1624 751
rect 1638 755 1644 756
rect 1638 751 1639 755
rect 1643 751 1644 755
rect 1638 750 1644 751
rect 1659 755 1665 756
rect 1659 751 1660 755
rect 1664 754 1665 755
rect 1682 755 1688 756
rect 1682 754 1683 755
rect 1664 752 1683 754
rect 1664 751 1665 752
rect 1659 750 1665 751
rect 1682 751 1683 752
rect 1687 751 1688 755
rect 1682 750 1688 751
rect 1702 755 1708 756
rect 1702 751 1703 755
rect 1707 751 1708 755
rect 1702 750 1708 751
rect 1718 755 1729 756
rect 1718 751 1719 755
rect 1723 751 1724 755
rect 1728 751 1729 755
rect 1718 750 1729 751
rect 1774 755 1780 756
rect 1774 751 1775 755
rect 1779 751 1780 755
rect 1774 750 1780 751
rect 1782 755 1788 756
rect 1782 751 1783 755
rect 1787 754 1788 755
rect 1795 755 1801 756
rect 1795 754 1796 755
rect 1787 752 1796 754
rect 1787 751 1788 752
rect 1782 750 1788 751
rect 1795 751 1796 752
rect 1800 751 1801 755
rect 1795 750 1801 751
rect 1846 755 1852 756
rect 1846 751 1847 755
rect 1851 751 1852 755
rect 1867 755 1873 756
rect 1867 754 1868 755
rect 1846 750 1852 751
rect 1856 752 1868 754
rect 1038 747 1044 748
rect 1286 749 1292 750
rect 110 744 116 745
rect 1286 745 1287 749
rect 1291 745 1292 749
rect 1286 744 1292 745
rect 1602 743 1608 744
rect 1602 739 1603 743
rect 1607 742 1608 743
rect 1650 743 1656 744
rect 1650 742 1651 743
rect 1607 740 1651 742
rect 1607 739 1608 740
rect 1602 738 1608 739
rect 1650 739 1651 740
rect 1655 739 1656 743
rect 1856 742 1858 752
rect 1867 751 1868 752
rect 1872 751 1873 755
rect 1867 750 1873 751
rect 1934 755 1940 756
rect 1934 751 1935 755
rect 1939 751 1940 755
rect 1934 750 1940 751
rect 1955 755 1961 756
rect 1955 751 1956 755
rect 1960 754 1961 755
rect 2010 755 2016 756
rect 2010 754 2011 755
rect 1960 752 2011 754
rect 1960 751 1961 752
rect 1955 750 1961 751
rect 2010 751 2011 752
rect 2015 751 2016 755
rect 2010 750 2016 751
rect 2030 755 2036 756
rect 2030 751 2031 755
rect 2035 751 2036 755
rect 2030 750 2036 751
rect 2051 755 2057 756
rect 2051 751 2052 755
rect 2056 754 2057 755
rect 2114 755 2120 756
rect 2114 754 2115 755
rect 2056 752 2115 754
rect 2056 751 2057 752
rect 2051 750 2057 751
rect 2114 751 2115 752
rect 2119 751 2120 755
rect 2114 750 2120 751
rect 2134 755 2140 756
rect 2134 751 2135 755
rect 2139 751 2140 755
rect 2134 750 2140 751
rect 2155 755 2161 756
rect 2155 751 2156 755
rect 2160 754 2161 755
rect 2226 755 2232 756
rect 2226 754 2227 755
rect 2160 752 2227 754
rect 2160 751 2161 752
rect 2155 750 2161 751
rect 2226 751 2227 752
rect 2231 751 2232 755
rect 2226 750 2232 751
rect 2246 755 2252 756
rect 2246 751 2247 755
rect 2251 751 2252 755
rect 2267 755 2273 756
rect 2267 754 2268 755
rect 2246 750 2252 751
rect 2256 752 2268 754
rect 2142 747 2148 748
rect 2126 743 2132 744
rect 2126 742 2127 743
rect 1650 738 1656 739
rect 1756 740 1858 742
rect 1916 740 2127 742
rect 1756 738 1758 740
rect 1916 738 1918 740
rect 2126 739 2127 740
rect 2131 739 2132 743
rect 2142 743 2143 747
rect 2147 746 2148 747
rect 2256 746 2258 752
rect 2267 751 2268 752
rect 2272 751 2273 755
rect 2267 750 2273 751
rect 2358 755 2364 756
rect 2358 751 2359 755
rect 2363 751 2364 755
rect 2358 750 2364 751
rect 2374 755 2385 756
rect 2374 751 2375 755
rect 2379 751 2380 755
rect 2384 751 2385 755
rect 2374 750 2385 751
rect 2454 755 2460 756
rect 2454 751 2455 755
rect 2459 751 2460 755
rect 2454 750 2460 751
rect 2462 755 2468 756
rect 2462 751 2463 755
rect 2467 754 2468 755
rect 2475 755 2481 756
rect 2475 754 2476 755
rect 2467 752 2476 754
rect 2467 751 2468 752
rect 2462 750 2468 751
rect 2475 751 2476 752
rect 2480 751 2481 755
rect 2502 752 2503 756
rect 2507 752 2508 756
rect 2502 751 2508 752
rect 2475 750 2481 751
rect 2147 744 2258 746
rect 2147 743 2148 744
rect 2142 742 2148 743
rect 2126 738 2132 739
rect 1755 737 1761 738
rect 1563 735 1569 736
rect 110 732 116 733
rect 1286 732 1292 733
rect 110 728 111 732
rect 115 728 116 732
rect 110 727 116 728
rect 150 731 156 732
rect 150 727 151 731
rect 155 727 156 731
rect 150 726 156 727
rect 171 731 180 732
rect 171 727 172 731
rect 179 727 180 731
rect 171 726 180 727
rect 270 731 276 732
rect 270 727 271 731
rect 275 727 276 731
rect 291 731 297 732
rect 291 730 292 731
rect 270 726 276 727
rect 280 728 292 730
rect 280 718 282 728
rect 291 727 292 728
rect 296 727 297 731
rect 291 726 297 727
rect 406 731 412 732
rect 406 727 407 731
rect 411 727 412 731
rect 406 726 412 727
rect 427 731 433 732
rect 427 727 428 731
rect 432 727 433 731
rect 427 726 433 727
rect 534 731 540 732
rect 534 727 535 731
rect 539 727 540 731
rect 534 726 540 727
rect 555 731 561 732
rect 555 727 556 731
rect 560 730 561 731
rect 642 731 648 732
rect 642 730 643 731
rect 560 728 643 730
rect 560 727 561 728
rect 555 726 561 727
rect 642 727 643 728
rect 647 727 648 731
rect 642 726 648 727
rect 662 731 668 732
rect 662 727 663 731
rect 667 727 668 731
rect 662 726 668 727
rect 683 731 689 732
rect 683 727 684 731
rect 688 730 689 731
rect 722 731 728 732
rect 722 730 723 731
rect 688 728 723 730
rect 688 727 689 728
rect 683 726 689 727
rect 722 727 723 728
rect 727 727 728 731
rect 722 726 728 727
rect 790 731 796 732
rect 790 727 791 731
rect 795 727 796 731
rect 811 731 817 732
rect 811 730 812 731
rect 790 726 796 727
rect 800 728 812 730
rect 429 722 431 726
rect 133 716 282 718
rect 319 720 431 722
rect 133 714 135 716
rect 319 714 321 720
rect 800 718 802 728
rect 811 727 812 728
rect 816 727 817 731
rect 811 726 817 727
rect 918 731 924 732
rect 918 727 919 731
rect 923 727 924 731
rect 918 726 924 727
rect 939 731 945 732
rect 939 727 940 731
rect 944 730 945 731
rect 1034 731 1040 732
rect 1034 730 1035 731
rect 944 728 1035 730
rect 944 727 945 728
rect 939 726 945 727
rect 1034 727 1035 728
rect 1039 727 1040 731
rect 1034 726 1040 727
rect 1054 731 1060 732
rect 1054 727 1055 731
rect 1059 727 1060 731
rect 1054 726 1060 727
rect 1074 731 1081 732
rect 1074 727 1075 731
rect 1080 727 1081 731
rect 1286 728 1287 732
rect 1291 728 1292 732
rect 1563 731 1564 735
rect 1568 734 1569 735
rect 1610 735 1616 736
rect 1610 734 1611 735
rect 1568 732 1611 734
rect 1568 731 1569 732
rect 1563 730 1569 731
rect 1610 731 1611 732
rect 1615 731 1616 735
rect 1610 730 1616 731
rect 1618 735 1625 736
rect 1618 731 1619 735
rect 1624 731 1625 735
rect 1618 730 1625 731
rect 1682 735 1689 736
rect 1682 731 1683 735
rect 1688 731 1689 735
rect 1755 733 1756 737
rect 1760 733 1761 737
rect 1915 737 1921 738
rect 1755 732 1761 733
rect 1827 735 1833 736
rect 1682 730 1689 731
rect 1782 731 1788 732
rect 1782 730 1783 731
rect 1692 728 1783 730
rect 1286 727 1292 728
rect 1622 727 1628 728
rect 1074 726 1081 727
rect 1347 723 1353 724
rect 1347 719 1348 723
rect 1352 722 1353 723
rect 1411 723 1417 724
rect 1352 720 1406 722
rect 1352 719 1353 720
rect 1347 718 1353 719
rect 516 716 802 718
rect 516 714 518 716
rect 131 713 137 714
rect 131 709 132 713
rect 136 709 137 713
rect 131 708 137 709
rect 251 713 321 714
rect 251 709 252 713
rect 256 712 321 713
rect 515 713 521 714
rect 256 709 257 712
rect 251 708 257 709
rect 387 711 393 712
rect 387 707 388 711
rect 392 710 393 711
rect 494 711 500 712
rect 494 710 495 711
rect 392 708 495 710
rect 392 707 393 708
rect 387 706 393 707
rect 494 707 495 708
rect 499 707 500 711
rect 515 709 516 713
rect 520 709 521 713
rect 515 708 521 709
rect 642 711 649 712
rect 494 706 500 707
rect 642 707 643 711
rect 648 707 649 711
rect 642 706 649 707
rect 771 711 777 712
rect 771 707 772 711
rect 776 710 777 711
rect 782 711 788 712
rect 782 710 783 711
rect 776 708 783 710
rect 776 707 777 708
rect 771 706 777 707
rect 782 707 783 708
rect 787 707 788 711
rect 782 706 788 707
rect 894 711 905 712
rect 894 707 895 711
rect 899 707 900 711
rect 904 707 905 711
rect 894 706 905 707
rect 1034 711 1041 712
rect 1034 707 1035 711
rect 1040 707 1041 711
rect 1404 710 1406 720
rect 1411 719 1412 723
rect 1416 722 1417 723
rect 1507 723 1513 724
rect 1416 720 1494 722
rect 1416 719 1417 720
rect 1411 718 1417 719
rect 1492 710 1494 720
rect 1507 719 1508 723
rect 1512 722 1513 723
rect 1602 723 1608 724
rect 1602 722 1603 723
rect 1512 720 1603 722
rect 1512 719 1513 720
rect 1507 718 1513 719
rect 1602 719 1603 720
rect 1607 719 1608 723
rect 1602 718 1608 719
rect 1611 723 1617 724
rect 1611 719 1612 723
rect 1616 719 1617 723
rect 1622 723 1623 727
rect 1627 726 1628 727
rect 1692 726 1694 728
rect 1782 727 1783 728
rect 1787 727 1788 731
rect 1827 731 1828 735
rect 1832 734 1833 735
rect 1854 735 1860 736
rect 1854 734 1855 735
rect 1832 732 1855 734
rect 1832 731 1833 732
rect 1827 730 1833 731
rect 1854 731 1855 732
rect 1859 731 1860 735
rect 1915 733 1916 737
rect 1920 733 1921 737
rect 1915 732 1921 733
rect 2010 735 2017 736
rect 1854 730 1860 731
rect 2010 731 2011 735
rect 2016 731 2017 735
rect 2010 730 2017 731
rect 2114 735 2121 736
rect 2114 731 2115 735
rect 2120 731 2121 735
rect 2114 730 2121 731
rect 2226 735 2233 736
rect 2226 731 2227 735
rect 2232 731 2233 735
rect 2226 730 2233 731
rect 2339 735 2345 736
rect 2339 731 2340 735
rect 2344 734 2345 735
rect 2386 735 2392 736
rect 2386 734 2387 735
rect 2344 732 2387 734
rect 2344 731 2345 732
rect 2339 730 2345 731
rect 2386 731 2387 732
rect 2391 731 2392 735
rect 2386 730 2392 731
rect 2435 735 2441 736
rect 2435 731 2436 735
rect 2440 734 2441 735
rect 2470 735 2476 736
rect 2470 734 2471 735
rect 2440 732 2471 734
rect 2440 731 2441 732
rect 2435 730 2441 731
rect 2470 731 2471 732
rect 2475 731 2476 735
rect 2470 730 2476 731
rect 1782 726 1788 727
rect 1627 724 1694 726
rect 1627 723 1628 724
rect 1622 722 1628 723
rect 1715 723 1724 724
rect 1611 718 1617 719
rect 1715 719 1716 723
rect 1723 719 1724 723
rect 1715 718 1724 719
rect 1819 723 1825 724
rect 1819 719 1820 723
rect 1824 722 1825 723
rect 1854 723 1860 724
rect 1854 722 1855 723
rect 1824 720 1855 722
rect 1824 719 1825 720
rect 1819 718 1825 719
rect 1854 719 1855 720
rect 1859 719 1860 723
rect 1854 718 1860 719
rect 1862 723 1868 724
rect 1862 719 1863 723
rect 1867 722 1868 723
rect 1923 723 1929 724
rect 1923 722 1924 723
rect 1867 720 1924 722
rect 1867 719 1868 720
rect 1862 718 1868 719
rect 1923 719 1924 720
rect 1928 719 1929 723
rect 1923 718 1929 719
rect 1966 723 1972 724
rect 1966 719 1967 723
rect 1971 722 1972 723
rect 2027 723 2033 724
rect 2027 722 2028 723
rect 1971 720 2028 722
rect 1971 719 1972 720
rect 1966 718 1972 719
rect 2027 719 2028 720
rect 2032 719 2033 723
rect 2027 718 2033 719
rect 2131 723 2137 724
rect 2131 719 2132 723
rect 2136 722 2137 723
rect 2142 723 2148 724
rect 2142 722 2143 723
rect 2136 720 2143 722
rect 2136 719 2137 720
rect 2131 718 2137 719
rect 2142 719 2143 720
rect 2147 719 2148 723
rect 2142 718 2148 719
rect 2174 723 2180 724
rect 2174 719 2175 723
rect 2179 722 2180 723
rect 2235 723 2241 724
rect 2235 722 2236 723
rect 2179 720 2236 722
rect 2179 719 2180 720
rect 2174 718 2180 719
rect 2235 719 2236 720
rect 2240 719 2241 723
rect 2235 718 2241 719
rect 2278 723 2284 724
rect 2278 719 2279 723
rect 2283 722 2284 723
rect 2347 723 2353 724
rect 2347 722 2348 723
rect 2283 720 2348 722
rect 2283 719 2284 720
rect 2278 718 2284 719
rect 2347 719 2348 720
rect 2352 719 2353 723
rect 2347 718 2353 719
rect 2435 723 2441 724
rect 2435 719 2436 723
rect 2440 722 2441 723
rect 2462 723 2468 724
rect 2462 722 2463 723
rect 2440 720 2463 722
rect 2440 719 2441 720
rect 2435 718 2441 719
rect 2462 719 2463 720
rect 2467 719 2468 723
rect 2462 718 2468 719
rect 1613 710 1615 718
rect 1034 706 1041 707
rect 1159 708 1391 710
rect 1404 708 1454 710
rect 1492 708 1551 710
rect 1613 708 1758 710
rect 1159 706 1161 708
rect 1389 706 1391 708
rect 1452 706 1454 708
rect 1549 706 1551 708
rect 1756 706 1758 708
rect 1108 704 1161 706
rect 1366 705 1372 706
rect 1326 704 1332 705
rect 1108 702 1110 704
rect 1107 701 1113 702
rect 131 699 137 700
rect 131 695 132 699
rect 136 695 137 699
rect 131 694 137 695
rect 174 699 180 700
rect 174 695 175 699
rect 179 698 180 699
rect 187 699 193 700
rect 187 698 188 699
rect 179 696 188 698
rect 179 695 180 696
rect 174 694 180 695
rect 187 695 188 696
rect 192 695 193 699
rect 187 694 193 695
rect 230 699 236 700
rect 230 695 231 699
rect 235 698 236 699
rect 275 699 281 700
rect 275 698 276 699
rect 235 696 276 698
rect 235 695 236 696
rect 230 694 236 695
rect 275 695 276 696
rect 280 695 281 699
rect 275 694 281 695
rect 343 699 349 700
rect 343 695 344 699
rect 348 698 349 699
rect 371 699 377 700
rect 371 698 372 699
rect 348 696 372 698
rect 348 695 349 696
rect 343 694 349 695
rect 371 695 372 696
rect 376 695 377 699
rect 371 694 377 695
rect 414 699 420 700
rect 414 695 415 699
rect 419 698 420 699
rect 483 699 489 700
rect 483 698 484 699
rect 419 696 484 698
rect 419 695 420 696
rect 414 694 420 695
rect 483 695 484 696
rect 488 695 489 699
rect 483 694 489 695
rect 603 699 609 700
rect 603 695 604 699
rect 608 698 609 699
rect 722 699 729 700
rect 608 696 719 698
rect 608 695 609 696
rect 603 694 609 695
rect 133 690 135 694
rect 286 691 292 692
rect 286 690 287 691
rect 133 688 287 690
rect 286 687 287 688
rect 291 687 292 691
rect 286 686 292 687
rect 494 687 500 688
rect 494 683 495 687
rect 499 686 500 687
rect 717 686 719 696
rect 722 695 723 699
rect 728 695 729 699
rect 722 694 729 695
rect 851 699 857 700
rect 851 695 852 699
rect 856 698 857 699
rect 974 699 985 700
rect 856 696 950 698
rect 856 695 857 696
rect 851 694 857 695
rect 948 686 950 696
rect 974 695 975 699
rect 979 695 980 699
rect 984 695 985 699
rect 1107 697 1108 701
rect 1112 697 1113 701
rect 1326 700 1327 704
rect 1331 700 1332 704
rect 1366 701 1367 705
rect 1371 701 1372 705
rect 1366 700 1372 701
rect 1387 705 1393 706
rect 1387 701 1388 705
rect 1392 701 1393 705
rect 1387 700 1393 701
rect 1430 705 1436 706
rect 1430 701 1431 705
rect 1435 701 1436 705
rect 1430 700 1436 701
rect 1451 705 1457 706
rect 1451 701 1452 705
rect 1456 701 1457 705
rect 1451 700 1457 701
rect 1526 705 1532 706
rect 1526 701 1527 705
rect 1531 701 1532 705
rect 1526 700 1532 701
rect 1547 705 1553 706
rect 1547 701 1548 705
rect 1552 701 1553 705
rect 1547 700 1553 701
rect 1630 705 1636 706
rect 1630 701 1631 705
rect 1635 701 1636 705
rect 1734 705 1740 706
rect 1630 700 1636 701
rect 1650 703 1657 704
rect 1107 696 1113 697
rect 1150 699 1156 700
rect 974 694 985 695
rect 1150 695 1151 699
rect 1155 698 1156 699
rect 1219 699 1225 700
rect 1326 699 1332 700
rect 1650 699 1651 703
rect 1656 699 1657 703
rect 1734 701 1735 705
rect 1739 701 1740 705
rect 1734 700 1740 701
rect 1755 705 1761 706
rect 1755 701 1756 705
rect 1760 701 1761 705
rect 1755 700 1761 701
rect 1838 705 1844 706
rect 1838 701 1839 705
rect 1843 701 1844 705
rect 1942 705 1948 706
rect 1838 700 1844 701
rect 1859 703 1868 704
rect 1219 698 1220 699
rect 1155 696 1220 698
rect 1155 695 1156 696
rect 1150 694 1156 695
rect 1219 695 1220 696
rect 1224 695 1225 699
rect 1650 698 1657 699
rect 1859 699 1860 703
rect 1867 699 1868 703
rect 1942 701 1943 705
rect 1947 701 1948 705
rect 2046 705 2052 706
rect 1942 700 1948 701
rect 1963 703 1972 704
rect 1859 698 1868 699
rect 1963 699 1964 703
rect 1971 699 1972 703
rect 2046 701 2047 705
rect 2051 701 2052 705
rect 2150 705 2156 706
rect 2046 700 2052 701
rect 2062 703 2073 704
rect 1963 698 1972 699
rect 2062 699 2063 703
rect 2067 699 2068 703
rect 2072 699 2073 703
rect 2150 701 2151 705
rect 2155 701 2156 705
rect 2254 705 2260 706
rect 2150 700 2156 701
rect 2171 703 2180 704
rect 2062 698 2073 699
rect 2171 699 2172 703
rect 2179 699 2180 703
rect 2254 701 2255 705
rect 2259 701 2260 705
rect 2366 705 2372 706
rect 2254 700 2260 701
rect 2275 703 2284 704
rect 2171 698 2180 699
rect 2275 699 2276 703
rect 2283 699 2284 703
rect 2366 701 2367 705
rect 2371 701 2372 705
rect 2454 705 2460 706
rect 2366 700 2372 701
rect 2386 703 2393 704
rect 2275 698 2284 699
rect 2386 699 2387 703
rect 2392 699 2393 703
rect 2454 701 2455 705
rect 2459 701 2460 705
rect 2502 704 2508 705
rect 2454 700 2460 701
rect 2470 703 2481 704
rect 2386 698 2393 699
rect 2470 699 2471 703
rect 2475 699 2476 703
rect 2480 699 2481 703
rect 2502 700 2503 704
rect 2507 700 2508 704
rect 2502 699 2508 700
rect 2470 698 2481 699
rect 1219 694 1225 695
rect 1326 687 1332 688
rect 499 684 526 686
rect 717 684 766 686
rect 948 684 1022 686
rect 499 683 500 684
rect 494 682 500 683
rect 524 682 526 684
rect 764 682 766 684
rect 1020 682 1022 684
rect 1326 683 1327 687
rect 1331 683 1332 687
rect 2502 687 2508 688
rect 1326 682 1332 683
rect 1350 684 1356 685
rect 150 681 156 682
rect 110 680 116 681
rect 110 676 111 680
rect 115 676 116 680
rect 150 677 151 681
rect 155 677 156 681
rect 206 681 212 682
rect 150 676 156 677
rect 171 679 180 680
rect 110 675 116 676
rect 171 675 172 679
rect 179 675 180 679
rect 206 677 207 681
rect 211 677 212 681
rect 294 681 300 682
rect 206 676 212 677
rect 227 679 236 680
rect 171 674 180 675
rect 227 675 228 679
rect 235 675 236 679
rect 294 677 295 681
rect 299 677 300 681
rect 390 681 396 682
rect 294 676 300 677
rect 315 679 321 680
rect 227 674 236 675
rect 315 675 316 679
rect 320 678 321 679
rect 343 679 349 680
rect 343 678 344 679
rect 320 676 344 678
rect 320 675 321 676
rect 315 674 321 675
rect 343 675 344 676
rect 348 675 349 679
rect 390 677 391 681
rect 395 677 396 681
rect 502 681 508 682
rect 390 676 396 677
rect 411 679 420 680
rect 343 674 349 675
rect 411 675 412 679
rect 419 675 420 679
rect 502 677 503 681
rect 507 677 508 681
rect 502 676 508 677
rect 523 681 529 682
rect 523 677 524 681
rect 528 677 529 681
rect 523 676 529 677
rect 622 681 628 682
rect 622 677 623 681
rect 627 677 628 681
rect 742 681 748 682
rect 622 676 628 677
rect 643 679 652 680
rect 411 674 420 675
rect 643 675 644 679
rect 651 675 652 679
rect 742 677 743 681
rect 747 677 748 681
rect 742 676 748 677
rect 763 681 769 682
rect 763 677 764 681
rect 768 677 769 681
rect 763 676 769 677
rect 870 681 876 682
rect 870 677 871 681
rect 875 677 876 681
rect 998 681 1004 682
rect 870 676 876 677
rect 891 679 900 680
rect 643 674 652 675
rect 891 675 892 679
rect 899 675 900 679
rect 998 677 999 681
rect 1003 677 1004 681
rect 998 676 1004 677
rect 1019 681 1025 682
rect 1019 677 1020 681
rect 1024 677 1025 681
rect 1019 676 1025 677
rect 1126 681 1132 682
rect 1126 677 1127 681
rect 1131 677 1132 681
rect 1238 681 1244 682
rect 1126 676 1132 677
rect 1147 679 1156 680
rect 891 674 900 675
rect 1147 675 1148 679
rect 1155 675 1156 679
rect 1238 677 1239 681
rect 1243 677 1244 681
rect 1286 680 1292 681
rect 1238 676 1244 677
rect 1259 679 1265 680
rect 1147 674 1156 675
rect 1259 675 1260 679
rect 1264 675 1265 679
rect 1286 676 1287 680
rect 1291 676 1292 680
rect 1350 680 1351 684
rect 1355 680 1356 684
rect 1350 679 1356 680
rect 1414 684 1420 685
rect 1414 680 1415 684
rect 1419 680 1420 684
rect 1414 679 1420 680
rect 1510 684 1516 685
rect 1510 680 1511 684
rect 1515 680 1516 684
rect 1510 679 1516 680
rect 1614 684 1620 685
rect 1614 680 1615 684
rect 1619 680 1620 684
rect 1614 679 1620 680
rect 1718 684 1724 685
rect 1718 680 1719 684
rect 1723 680 1724 684
rect 1718 679 1724 680
rect 1822 684 1828 685
rect 1822 680 1823 684
rect 1827 680 1828 684
rect 1822 679 1828 680
rect 1926 684 1932 685
rect 1926 680 1927 684
rect 1931 680 1932 684
rect 1926 679 1932 680
rect 2030 684 2036 685
rect 2030 680 2031 684
rect 2035 680 2036 684
rect 2030 679 2036 680
rect 2134 684 2140 685
rect 2134 680 2135 684
rect 2139 680 2140 684
rect 2134 679 2140 680
rect 2238 684 2244 685
rect 2238 680 2239 684
rect 2243 680 2244 684
rect 2238 679 2244 680
rect 2350 684 2356 685
rect 2350 680 2351 684
rect 2355 680 2356 684
rect 2350 679 2356 680
rect 2438 684 2444 685
rect 2438 680 2439 684
rect 2443 680 2444 684
rect 2502 683 2503 687
rect 2507 683 2508 687
rect 2502 682 2508 683
rect 2438 679 2444 680
rect 1286 675 1292 676
rect 1259 674 1265 675
rect 1261 670 1263 674
rect 1342 671 1348 672
rect 1342 670 1343 671
rect 1261 668 1343 670
rect 1342 667 1343 668
rect 1347 667 1348 671
rect 1342 666 1348 667
rect 110 663 116 664
rect 110 659 111 663
rect 115 659 116 663
rect 1286 663 1292 664
rect 110 658 116 659
rect 134 660 140 661
rect 134 656 135 660
rect 139 656 140 660
rect 134 655 140 656
rect 190 660 196 661
rect 190 656 191 660
rect 195 656 196 660
rect 190 655 196 656
rect 278 660 284 661
rect 278 656 279 660
rect 283 656 284 660
rect 278 655 284 656
rect 374 660 380 661
rect 374 656 375 660
rect 379 656 380 660
rect 374 655 380 656
rect 486 660 492 661
rect 486 656 487 660
rect 491 656 492 660
rect 486 655 492 656
rect 606 660 612 661
rect 606 656 607 660
rect 611 656 612 660
rect 606 655 612 656
rect 726 660 732 661
rect 726 656 727 660
rect 731 656 732 660
rect 726 655 732 656
rect 854 660 860 661
rect 854 656 855 660
rect 859 656 860 660
rect 854 655 860 656
rect 982 660 988 661
rect 982 656 983 660
rect 987 656 988 660
rect 982 655 988 656
rect 1110 660 1116 661
rect 1110 656 1111 660
rect 1115 656 1116 660
rect 1110 655 1116 656
rect 1222 660 1228 661
rect 1222 656 1223 660
rect 1227 656 1228 660
rect 1286 659 1287 663
rect 1291 659 1292 663
rect 1286 658 1292 659
rect 1350 660 1356 661
rect 1222 655 1228 656
rect 1326 657 1332 658
rect 1326 653 1327 657
rect 1331 653 1332 657
rect 1350 656 1351 660
rect 1355 656 1356 660
rect 1350 655 1356 656
rect 1414 660 1420 661
rect 1414 656 1415 660
rect 1419 656 1420 660
rect 1414 655 1420 656
rect 1510 660 1516 661
rect 1510 656 1511 660
rect 1515 656 1516 660
rect 1510 655 1516 656
rect 1606 660 1612 661
rect 1606 656 1607 660
rect 1611 656 1612 660
rect 1606 655 1612 656
rect 1710 660 1716 661
rect 1710 656 1711 660
rect 1715 656 1716 660
rect 1710 655 1716 656
rect 1822 660 1828 661
rect 1822 656 1823 660
rect 1827 656 1828 660
rect 1822 655 1828 656
rect 1934 660 1940 661
rect 1934 656 1935 660
rect 1939 656 1940 660
rect 1934 655 1940 656
rect 2054 660 2060 661
rect 2054 656 2055 660
rect 2059 656 2060 660
rect 2054 655 2060 656
rect 2182 660 2188 661
rect 2182 656 2183 660
rect 2187 656 2188 660
rect 2182 655 2188 656
rect 2318 660 2324 661
rect 2318 656 2319 660
rect 2323 656 2324 660
rect 2318 655 2324 656
rect 2438 660 2444 661
rect 2438 656 2439 660
rect 2443 656 2444 660
rect 2438 655 2444 656
rect 2502 657 2508 658
rect 1326 652 1332 653
rect 2502 653 2503 657
rect 2507 653 2508 657
rect 2502 652 2508 653
rect 150 644 156 645
rect 110 641 116 642
rect 110 637 111 641
rect 115 637 116 641
rect 150 640 151 644
rect 155 640 156 644
rect 150 639 156 640
rect 262 644 268 645
rect 262 640 263 644
rect 267 640 268 644
rect 262 639 268 640
rect 366 644 372 645
rect 366 640 367 644
rect 371 640 372 644
rect 366 639 372 640
rect 462 644 468 645
rect 462 640 463 644
rect 467 640 468 644
rect 462 639 468 640
rect 558 644 564 645
rect 558 640 559 644
rect 563 640 564 644
rect 558 639 564 640
rect 654 644 660 645
rect 654 640 655 644
rect 659 640 660 644
rect 654 639 660 640
rect 750 644 756 645
rect 750 640 751 644
rect 755 640 756 644
rect 750 639 756 640
rect 846 644 852 645
rect 846 640 847 644
rect 851 640 852 644
rect 846 639 852 640
rect 942 644 948 645
rect 942 640 943 644
rect 947 640 948 644
rect 942 639 948 640
rect 1038 644 1044 645
rect 1038 640 1039 644
rect 1043 640 1044 644
rect 1038 639 1044 640
rect 1142 644 1148 645
rect 1142 640 1143 644
rect 1147 640 1148 644
rect 1142 639 1148 640
rect 1222 644 1228 645
rect 1222 640 1223 644
rect 1227 640 1228 644
rect 1222 639 1228 640
rect 1286 641 1292 642
rect 110 636 116 637
rect 1286 637 1287 641
rect 1291 637 1292 641
rect 1286 636 1292 637
rect 1326 640 1332 641
rect 2502 640 2508 641
rect 1326 636 1327 640
rect 1331 636 1332 640
rect 1326 635 1332 636
rect 1366 639 1372 640
rect 1366 635 1367 639
rect 1371 635 1372 639
rect 1366 634 1372 635
rect 1387 639 1393 640
rect 1387 635 1388 639
rect 1392 638 1393 639
rect 1410 639 1416 640
rect 1410 638 1411 639
rect 1392 636 1411 638
rect 1392 635 1393 636
rect 1387 634 1393 635
rect 1410 635 1411 636
rect 1415 635 1416 639
rect 1410 634 1416 635
rect 1430 639 1436 640
rect 1430 635 1431 639
rect 1435 635 1436 639
rect 1430 634 1436 635
rect 1451 639 1457 640
rect 1451 635 1452 639
rect 1456 638 1457 639
rect 1506 639 1512 640
rect 1506 638 1507 639
rect 1456 636 1507 638
rect 1456 635 1457 636
rect 1451 634 1457 635
rect 1506 635 1507 636
rect 1511 635 1512 639
rect 1506 634 1512 635
rect 1526 639 1532 640
rect 1526 635 1527 639
rect 1531 635 1532 639
rect 1526 634 1532 635
rect 1534 639 1540 640
rect 1534 635 1535 639
rect 1539 638 1540 639
rect 1547 639 1553 640
rect 1547 638 1548 639
rect 1539 636 1548 638
rect 1539 635 1540 636
rect 1534 634 1540 635
rect 1547 635 1548 636
rect 1552 635 1553 639
rect 1547 634 1553 635
rect 1622 639 1628 640
rect 1622 635 1623 639
rect 1627 635 1628 639
rect 1643 639 1649 640
rect 1643 638 1644 639
rect 1622 634 1628 635
rect 1632 636 1644 638
rect 1262 631 1268 632
rect 1262 627 1263 631
rect 1267 630 1268 631
rect 1632 630 1634 636
rect 1643 635 1644 636
rect 1648 635 1649 639
rect 1643 634 1649 635
rect 1726 639 1732 640
rect 1726 635 1727 639
rect 1731 635 1732 639
rect 1726 634 1732 635
rect 1747 639 1753 640
rect 1747 635 1748 639
rect 1752 635 1753 639
rect 1747 634 1753 635
rect 1838 639 1844 640
rect 1838 635 1839 639
rect 1843 635 1844 639
rect 1838 634 1844 635
rect 1854 639 1865 640
rect 1854 635 1855 639
rect 1859 635 1860 639
rect 1864 635 1865 639
rect 1854 634 1865 635
rect 1950 639 1956 640
rect 1950 635 1951 639
rect 1955 635 1956 639
rect 1971 639 1977 640
rect 1971 638 1972 639
rect 1950 634 1956 635
rect 1960 636 1972 638
rect 1267 628 1634 630
rect 1267 627 1268 628
rect 1262 626 1268 627
rect 1749 626 1751 634
rect 1960 626 1962 636
rect 1971 635 1972 636
rect 1976 635 1977 639
rect 1971 634 1977 635
rect 2070 639 2076 640
rect 2070 635 2071 639
rect 2075 635 2076 639
rect 2070 634 2076 635
rect 2091 639 2097 640
rect 2091 635 2092 639
rect 2096 638 2097 639
rect 2178 639 2184 640
rect 2178 638 2179 639
rect 2096 636 2179 638
rect 2096 635 2097 636
rect 2091 634 2097 635
rect 2178 635 2179 636
rect 2183 635 2184 639
rect 2178 634 2184 635
rect 2198 639 2204 640
rect 2198 635 2199 639
rect 2203 635 2204 639
rect 2198 634 2204 635
rect 2219 639 2225 640
rect 2219 635 2220 639
rect 2224 638 2225 639
rect 2314 639 2320 640
rect 2314 638 2315 639
rect 2224 636 2315 638
rect 2224 635 2225 636
rect 2219 634 2225 635
rect 2314 635 2315 636
rect 2319 635 2320 639
rect 2314 634 2320 635
rect 2334 639 2340 640
rect 2334 635 2335 639
rect 2339 635 2340 639
rect 2334 634 2340 635
rect 2350 639 2361 640
rect 2350 635 2351 639
rect 2355 635 2356 639
rect 2360 635 2361 639
rect 2350 634 2361 635
rect 2454 639 2460 640
rect 2454 635 2455 639
rect 2459 635 2460 639
rect 2454 634 2460 635
rect 2462 639 2468 640
rect 2462 635 2463 639
rect 2467 638 2468 639
rect 2475 639 2481 640
rect 2475 638 2476 639
rect 2467 636 2476 638
rect 2467 635 2468 636
rect 2462 634 2468 635
rect 2475 635 2476 636
rect 2480 635 2481 639
rect 2502 636 2503 640
rect 2507 636 2508 640
rect 2502 635 2508 636
rect 2475 634 2481 635
rect 110 624 116 625
rect 1286 624 1292 625
rect 110 620 111 624
rect 115 620 116 624
rect 110 619 116 620
rect 166 623 172 624
rect 166 619 167 623
rect 171 619 172 623
rect 166 618 172 619
rect 187 623 193 624
rect 187 619 188 623
rect 192 622 193 623
rect 258 623 264 624
rect 258 622 259 623
rect 192 620 259 622
rect 192 619 193 620
rect 187 618 193 619
rect 258 619 259 620
rect 263 619 264 623
rect 258 618 264 619
rect 278 623 284 624
rect 278 619 279 623
rect 283 619 284 623
rect 278 618 284 619
rect 286 623 292 624
rect 286 619 287 623
rect 291 622 292 623
rect 299 623 305 624
rect 299 622 300 623
rect 291 620 300 622
rect 291 619 292 620
rect 286 618 292 619
rect 299 619 300 620
rect 304 619 305 623
rect 299 618 305 619
rect 382 623 388 624
rect 382 619 383 623
rect 387 619 388 623
rect 382 618 388 619
rect 403 623 412 624
rect 403 619 404 623
rect 411 619 412 623
rect 403 618 412 619
rect 478 623 484 624
rect 478 619 479 623
rect 483 619 484 623
rect 478 618 484 619
rect 486 623 492 624
rect 486 619 487 623
rect 491 622 492 623
rect 499 623 505 624
rect 499 622 500 623
rect 491 620 500 622
rect 491 619 492 620
rect 486 618 492 619
rect 499 619 500 620
rect 504 619 505 623
rect 499 618 505 619
rect 574 623 580 624
rect 574 619 575 623
rect 579 619 580 623
rect 595 623 601 624
rect 595 622 596 623
rect 574 618 580 619
rect 584 620 596 622
rect 584 614 586 620
rect 595 619 596 620
rect 600 619 601 623
rect 595 618 601 619
rect 670 623 676 624
rect 670 619 671 623
rect 675 619 676 623
rect 691 623 697 624
rect 691 622 692 623
rect 670 618 676 619
rect 680 620 692 622
rect 461 612 586 614
rect 461 606 463 612
rect 680 610 682 620
rect 691 619 692 620
rect 696 619 697 623
rect 691 618 697 619
rect 766 623 772 624
rect 766 619 767 623
rect 771 619 772 623
rect 766 618 772 619
rect 787 623 793 624
rect 787 619 788 623
rect 792 622 793 623
rect 842 623 848 624
rect 842 622 843 623
rect 792 620 843 622
rect 792 619 793 620
rect 787 618 793 619
rect 842 619 843 620
rect 847 619 848 623
rect 842 618 848 619
rect 862 623 868 624
rect 862 619 863 623
rect 867 619 868 623
rect 862 618 868 619
rect 883 623 889 624
rect 883 619 884 623
rect 888 622 889 623
rect 938 623 944 624
rect 938 622 939 623
rect 888 620 939 622
rect 888 619 889 620
rect 883 618 889 619
rect 938 619 939 620
rect 943 619 944 623
rect 938 618 944 619
rect 958 623 964 624
rect 958 619 959 623
rect 963 619 964 623
rect 958 618 964 619
rect 974 623 985 624
rect 974 619 975 623
rect 979 619 980 623
rect 984 619 985 623
rect 974 618 985 619
rect 1054 623 1060 624
rect 1054 619 1055 623
rect 1059 619 1060 623
rect 1054 618 1060 619
rect 1075 623 1081 624
rect 1075 619 1076 623
rect 1080 622 1081 623
rect 1138 623 1144 624
rect 1138 622 1139 623
rect 1080 620 1139 622
rect 1080 619 1081 620
rect 1075 618 1081 619
rect 1138 619 1139 620
rect 1143 619 1144 623
rect 1138 618 1144 619
rect 1158 623 1164 624
rect 1158 619 1159 623
rect 1163 619 1164 623
rect 1158 618 1164 619
rect 1166 623 1172 624
rect 1166 619 1167 623
rect 1171 622 1172 623
rect 1179 623 1185 624
rect 1179 622 1180 623
rect 1171 620 1180 622
rect 1171 619 1172 620
rect 1166 618 1172 619
rect 1179 619 1180 620
rect 1184 619 1185 623
rect 1179 618 1185 619
rect 1238 623 1244 624
rect 1238 619 1239 623
rect 1243 619 1244 623
rect 1238 618 1244 619
rect 1259 623 1265 624
rect 1259 619 1260 623
rect 1264 619 1265 623
rect 1286 620 1287 624
rect 1291 620 1292 624
rect 1604 624 1751 626
rect 1820 624 1962 626
rect 1604 622 1606 624
rect 1820 622 1822 624
rect 1603 621 1609 622
rect 1286 619 1292 620
rect 1342 619 1353 620
rect 1259 618 1265 619
rect 1261 614 1263 618
rect 1342 615 1343 619
rect 1347 615 1348 619
rect 1352 615 1353 619
rect 1342 614 1353 615
rect 1410 619 1417 620
rect 1410 615 1411 619
rect 1416 615 1417 619
rect 1410 614 1417 615
rect 1506 619 1513 620
rect 1506 615 1507 619
rect 1512 615 1513 619
rect 1603 617 1604 621
rect 1608 617 1609 621
rect 1819 621 1825 622
rect 1603 616 1609 617
rect 1707 619 1713 620
rect 1506 614 1513 615
rect 1534 615 1540 616
rect 1534 614 1535 615
rect 1159 612 1263 614
rect 1516 612 1535 614
rect 1159 610 1161 612
rect 1516 610 1518 612
rect 1534 611 1535 612
rect 1539 611 1540 615
rect 1707 615 1708 619
rect 1712 618 1713 619
rect 1762 619 1768 620
rect 1762 618 1763 619
rect 1712 616 1763 618
rect 1712 615 1713 616
rect 1707 614 1713 615
rect 1762 615 1763 616
rect 1767 615 1768 619
rect 1819 617 1820 621
rect 1824 617 1825 621
rect 1819 616 1825 617
rect 1931 619 1937 620
rect 1762 614 1768 615
rect 1931 615 1932 619
rect 1936 618 1937 619
rect 2042 619 2048 620
rect 2042 618 2043 619
rect 1936 616 2043 618
rect 1936 615 1937 616
rect 1931 614 1937 615
rect 2042 615 2043 616
rect 2047 615 2048 619
rect 2042 614 2048 615
rect 2051 619 2057 620
rect 2051 615 2052 619
rect 2056 618 2057 619
rect 2062 619 2068 620
rect 2062 618 2063 619
rect 2056 616 2063 618
rect 2056 615 2057 616
rect 2051 614 2057 615
rect 2062 615 2063 616
rect 2067 615 2068 619
rect 2062 614 2068 615
rect 2178 619 2185 620
rect 2178 615 2179 619
rect 2184 615 2185 619
rect 2178 614 2185 615
rect 2314 619 2321 620
rect 2314 615 2315 619
rect 2320 615 2321 619
rect 2314 614 2321 615
rect 2435 619 2441 620
rect 2435 615 2436 619
rect 2440 618 2441 619
rect 2470 619 2476 620
rect 2470 618 2471 619
rect 2440 616 2471 618
rect 2440 615 2441 616
rect 2435 614 2441 615
rect 2470 615 2471 616
rect 2475 615 2476 619
rect 2470 614 2476 615
rect 1534 610 1540 611
rect 556 608 682 610
rect 1036 608 1161 610
rect 1443 609 1518 610
rect 556 606 558 608
rect 1036 606 1038 608
rect 1363 607 1369 608
rect 459 605 465 606
rect 147 603 153 604
rect 147 599 148 603
rect 152 602 153 603
rect 158 603 164 604
rect 158 602 159 603
rect 152 600 159 602
rect 152 599 153 600
rect 147 598 153 599
rect 158 599 159 600
rect 163 599 164 603
rect 158 598 164 599
rect 258 603 265 604
rect 258 599 259 603
rect 264 599 265 603
rect 258 598 265 599
rect 363 603 369 604
rect 363 599 364 603
rect 368 602 369 603
rect 368 600 434 602
rect 459 601 460 605
rect 464 601 465 605
rect 459 600 465 601
rect 555 605 561 606
rect 555 601 556 605
rect 560 601 561 605
rect 1035 605 1041 606
rect 555 600 561 601
rect 646 603 657 604
rect 368 599 369 600
rect 363 598 369 599
rect 432 598 434 600
rect 486 599 492 600
rect 486 598 487 599
rect 432 596 487 598
rect 486 595 487 596
rect 491 595 492 599
rect 646 599 647 603
rect 651 599 652 603
rect 656 599 657 603
rect 646 598 657 599
rect 747 603 753 604
rect 747 599 748 603
rect 752 602 753 603
rect 834 603 840 604
rect 834 602 835 603
rect 752 600 835 602
rect 752 599 753 600
rect 747 598 753 599
rect 834 599 835 600
rect 839 599 840 603
rect 834 598 840 599
rect 842 603 849 604
rect 842 599 843 603
rect 848 599 849 603
rect 842 598 849 599
rect 938 603 945 604
rect 938 599 939 603
rect 944 599 945 603
rect 1035 601 1036 605
rect 1040 601 1041 605
rect 1035 600 1041 601
rect 1138 603 1145 604
rect 938 598 945 599
rect 1018 599 1024 600
rect 1018 598 1019 599
rect 486 594 492 595
rect 972 596 1019 598
rect 972 594 974 596
rect 1018 595 1019 596
rect 1023 595 1024 599
rect 1138 599 1139 603
rect 1144 599 1145 603
rect 1138 598 1145 599
rect 1219 603 1225 604
rect 1219 599 1220 603
rect 1224 602 1225 603
rect 1262 603 1268 604
rect 1262 602 1263 603
rect 1224 600 1263 602
rect 1224 599 1225 600
rect 1219 598 1225 599
rect 1262 599 1263 600
rect 1267 599 1268 603
rect 1363 603 1364 607
rect 1368 606 1369 607
rect 1368 604 1438 606
rect 1443 605 1444 609
rect 1448 608 1518 609
rect 1448 605 1449 608
rect 1443 604 1449 605
rect 1531 607 1537 608
rect 1368 603 1369 604
rect 1363 602 1369 603
rect 1262 598 1268 599
rect 1018 594 1024 595
rect 1436 594 1438 604
rect 1531 603 1532 607
rect 1536 606 1537 607
rect 1574 607 1580 608
rect 1536 604 1570 606
rect 1536 603 1537 604
rect 1531 602 1537 603
rect 1568 598 1570 604
rect 1574 603 1575 607
rect 1579 606 1580 607
rect 1627 607 1633 608
rect 1627 606 1628 607
rect 1579 604 1628 606
rect 1579 603 1580 604
rect 1574 602 1580 603
rect 1627 603 1628 604
rect 1632 603 1633 607
rect 1627 602 1633 603
rect 1695 607 1701 608
rect 1695 603 1696 607
rect 1700 606 1701 607
rect 1723 607 1729 608
rect 1723 606 1724 607
rect 1700 604 1724 606
rect 1700 603 1701 604
rect 1695 602 1701 603
rect 1723 603 1724 604
rect 1728 603 1729 607
rect 1723 602 1729 603
rect 1827 607 1833 608
rect 1827 603 1828 607
rect 1832 606 1833 607
rect 1870 607 1876 608
rect 1832 604 1866 606
rect 1832 603 1833 604
rect 1827 602 1833 603
rect 1586 599 1592 600
rect 1586 598 1587 599
rect 1568 596 1587 598
rect 1586 595 1587 596
rect 1591 595 1592 599
rect 1864 598 1866 604
rect 1870 603 1871 607
rect 1875 606 1876 607
rect 1939 607 1945 608
rect 1939 606 1940 607
rect 1875 604 1940 606
rect 1875 603 1876 604
rect 1870 602 1876 603
rect 1939 603 1940 604
rect 1944 603 1945 607
rect 1939 602 1945 603
rect 1982 607 1988 608
rect 1982 603 1983 607
rect 1987 606 1988 607
rect 2059 607 2065 608
rect 2059 606 2060 607
rect 1987 604 2060 606
rect 1987 603 1988 604
rect 1982 602 1988 603
rect 2059 603 2060 604
rect 2064 603 2065 607
rect 2059 602 2065 603
rect 2187 607 2193 608
rect 2187 603 2188 607
rect 2192 606 2193 607
rect 2323 607 2329 608
rect 2192 604 2318 606
rect 2192 603 2193 604
rect 2187 602 2193 603
rect 1890 599 1896 600
rect 1890 598 1891 599
rect 1864 596 1891 598
rect 1586 594 1592 595
rect 1890 595 1891 596
rect 1895 595 1896 599
rect 1890 594 1896 595
rect 2042 595 2048 596
rect 891 593 974 594
rect 131 591 137 592
rect 131 587 132 591
rect 136 587 137 591
rect 131 586 137 587
rect 219 591 225 592
rect 219 587 220 591
rect 224 590 225 591
rect 286 591 292 592
rect 224 588 271 590
rect 224 587 225 588
rect 219 586 225 587
rect 133 578 135 586
rect 269 578 271 588
rect 286 587 287 591
rect 291 590 292 591
rect 315 591 321 592
rect 315 590 316 591
rect 291 588 316 590
rect 291 587 292 588
rect 286 586 292 587
rect 315 587 316 588
rect 320 587 321 591
rect 315 586 321 587
rect 406 591 417 592
rect 406 587 407 591
rect 411 587 412 591
rect 416 587 417 591
rect 406 586 417 587
rect 454 591 460 592
rect 454 587 455 591
rect 459 590 460 591
rect 515 591 521 592
rect 515 590 516 591
rect 459 588 516 590
rect 459 587 460 588
rect 454 586 460 587
rect 515 587 516 588
rect 520 587 521 591
rect 515 586 521 587
rect 558 591 564 592
rect 558 587 559 591
rect 563 590 564 591
rect 611 591 617 592
rect 611 590 612 591
rect 563 588 612 590
rect 563 587 564 588
rect 558 586 564 587
rect 611 587 612 588
rect 616 587 617 591
rect 611 586 617 587
rect 707 591 713 592
rect 707 587 708 591
rect 712 590 713 591
rect 742 591 748 592
rect 742 590 743 591
rect 712 588 743 590
rect 712 587 713 588
rect 707 586 713 587
rect 742 587 743 588
rect 747 587 748 591
rect 742 586 748 587
rect 750 591 756 592
rect 750 587 751 591
rect 755 590 756 591
rect 803 591 809 592
rect 803 590 804 591
rect 755 588 804 590
rect 755 587 756 588
rect 750 586 756 587
rect 803 587 804 588
rect 808 587 809 591
rect 891 589 892 593
rect 896 592 974 593
rect 1436 592 1486 594
rect 896 589 897 592
rect 891 588 897 589
rect 979 591 985 592
rect 803 586 809 587
rect 979 587 980 591
rect 984 587 985 591
rect 979 586 985 587
rect 1067 591 1073 592
rect 1067 587 1068 591
rect 1072 590 1073 591
rect 1163 591 1172 592
rect 1072 588 1161 590
rect 1072 587 1073 588
rect 1067 586 1073 587
rect 981 578 983 586
rect 1159 578 1161 588
rect 1163 587 1164 591
rect 1171 587 1172 591
rect 1484 590 1486 592
rect 2042 591 2043 595
rect 2047 594 2048 595
rect 2316 594 2318 604
rect 2323 603 2324 607
rect 2328 606 2329 607
rect 2350 607 2356 608
rect 2350 606 2351 607
rect 2328 604 2351 606
rect 2328 603 2329 604
rect 2323 602 2329 603
rect 2350 603 2351 604
rect 2355 603 2356 607
rect 2350 602 2356 603
rect 2435 607 2441 608
rect 2435 603 2436 607
rect 2440 606 2441 607
rect 2462 607 2468 608
rect 2462 606 2463 607
rect 2440 604 2463 606
rect 2440 603 2441 604
rect 2435 602 2441 603
rect 2462 603 2463 604
rect 2467 603 2468 607
rect 2462 602 2468 603
rect 2047 592 2103 594
rect 2316 592 2366 594
rect 2047 591 2048 592
rect 2042 590 2048 591
rect 2101 590 2103 592
rect 2364 590 2366 592
rect 1382 589 1388 590
rect 1163 586 1172 587
rect 1326 588 1332 589
rect 1326 584 1327 588
rect 1331 584 1332 588
rect 1382 585 1383 589
rect 1387 585 1388 589
rect 1462 589 1468 590
rect 1382 584 1388 585
rect 1398 587 1409 588
rect 1326 583 1332 584
rect 1398 583 1399 587
rect 1403 583 1404 587
rect 1408 583 1409 587
rect 1462 585 1463 589
rect 1467 585 1468 589
rect 1462 584 1468 585
rect 1483 589 1489 590
rect 1483 585 1484 589
rect 1488 585 1489 589
rect 1483 584 1489 585
rect 1550 589 1556 590
rect 1550 585 1551 589
rect 1555 585 1556 589
rect 1646 589 1652 590
rect 1550 584 1556 585
rect 1571 587 1580 588
rect 1398 582 1409 583
rect 1571 583 1572 587
rect 1579 583 1580 587
rect 1646 585 1647 589
rect 1651 585 1652 589
rect 1742 589 1748 590
rect 1646 584 1652 585
rect 1667 587 1673 588
rect 1571 582 1580 583
rect 1667 583 1668 587
rect 1672 586 1673 587
rect 1695 587 1701 588
rect 1695 586 1696 587
rect 1672 584 1696 586
rect 1672 583 1673 584
rect 1667 582 1673 583
rect 1695 583 1696 584
rect 1700 583 1701 587
rect 1742 585 1743 589
rect 1747 585 1748 589
rect 1846 589 1852 590
rect 1742 584 1748 585
rect 1762 587 1769 588
rect 1695 582 1701 583
rect 1762 583 1763 587
rect 1768 583 1769 587
rect 1846 585 1847 589
rect 1851 585 1852 589
rect 1958 589 1964 590
rect 1846 584 1852 585
rect 1867 587 1876 588
rect 1762 582 1769 583
rect 1867 583 1868 587
rect 1875 583 1876 587
rect 1958 585 1959 589
rect 1963 585 1964 589
rect 2078 589 2084 590
rect 1958 584 1964 585
rect 1979 587 1988 588
rect 1867 582 1876 583
rect 1979 583 1980 587
rect 1987 583 1988 587
rect 2078 585 2079 589
rect 2083 585 2084 589
rect 2078 584 2084 585
rect 2099 589 2105 590
rect 2099 585 2100 589
rect 2104 585 2105 589
rect 2099 584 2105 585
rect 2206 589 2212 590
rect 2206 585 2207 589
rect 2211 585 2212 589
rect 2342 589 2348 590
rect 2206 584 2212 585
rect 2214 587 2220 588
rect 1979 582 1988 583
rect 2214 583 2215 587
rect 2219 586 2220 587
rect 2227 587 2233 588
rect 2227 586 2228 587
rect 2219 584 2228 586
rect 2219 583 2220 584
rect 2214 582 2220 583
rect 2227 583 2228 584
rect 2232 583 2233 587
rect 2342 585 2343 589
rect 2347 585 2348 589
rect 2342 584 2348 585
rect 2363 589 2369 590
rect 2363 585 2364 589
rect 2368 585 2369 589
rect 2363 584 2369 585
rect 2454 589 2460 590
rect 2454 585 2455 589
rect 2459 585 2460 589
rect 2502 588 2508 589
rect 2454 584 2460 585
rect 2462 587 2468 588
rect 2227 582 2233 583
rect 2462 583 2463 587
rect 2467 586 2468 587
rect 2475 587 2481 588
rect 2475 586 2476 587
rect 2467 584 2476 586
rect 2467 583 2468 584
rect 2462 582 2468 583
rect 2475 583 2476 584
rect 2480 583 2481 587
rect 2502 584 2503 588
rect 2507 584 2508 588
rect 2502 583 2508 584
rect 2475 582 2481 583
rect 133 576 262 578
rect 269 576 359 578
rect 981 576 1110 578
rect 1159 576 1206 578
rect 260 574 262 576
rect 357 574 359 576
rect 1108 574 1110 576
rect 1204 574 1206 576
rect 150 573 156 574
rect 110 572 116 573
rect 110 568 111 572
rect 115 568 116 572
rect 150 569 151 573
rect 155 569 156 573
rect 238 573 244 574
rect 150 568 156 569
rect 158 571 164 572
rect 110 567 116 568
rect 158 567 159 571
rect 163 570 164 571
rect 171 571 177 572
rect 171 570 172 571
rect 163 568 172 570
rect 163 567 164 568
rect 158 566 164 567
rect 171 567 172 568
rect 176 567 177 571
rect 238 569 239 573
rect 243 569 244 573
rect 238 568 244 569
rect 259 573 265 574
rect 259 569 260 573
rect 264 569 265 573
rect 259 568 265 569
rect 334 573 340 574
rect 334 569 335 573
rect 339 569 340 573
rect 334 568 340 569
rect 355 573 361 574
rect 355 569 356 573
rect 360 569 361 573
rect 355 568 361 569
rect 430 573 436 574
rect 430 569 431 573
rect 435 569 436 573
rect 534 573 540 574
rect 430 568 436 569
rect 451 571 460 572
rect 171 566 177 567
rect 451 567 452 571
rect 459 567 460 571
rect 534 569 535 573
rect 539 569 540 573
rect 630 573 636 574
rect 534 568 540 569
rect 555 571 564 572
rect 451 566 460 567
rect 555 567 556 571
rect 563 567 564 571
rect 630 569 631 573
rect 635 569 636 573
rect 726 573 732 574
rect 630 568 636 569
rect 646 571 657 572
rect 555 566 564 567
rect 646 567 647 571
rect 651 567 652 571
rect 656 567 657 571
rect 726 569 727 573
rect 731 569 732 573
rect 822 573 828 574
rect 726 568 732 569
rect 747 571 756 572
rect 646 566 657 567
rect 747 567 748 571
rect 755 567 756 571
rect 822 569 823 573
rect 827 569 828 573
rect 910 573 916 574
rect 822 568 828 569
rect 834 571 840 572
rect 747 566 756 567
rect 834 567 835 571
rect 839 570 840 571
rect 843 571 849 572
rect 843 570 844 571
rect 839 568 844 570
rect 839 567 840 568
rect 834 566 840 567
rect 843 567 844 568
rect 848 567 849 571
rect 910 569 911 573
rect 915 569 916 573
rect 998 573 1004 574
rect 910 568 916 569
rect 931 571 937 572
rect 843 566 849 567
rect 931 567 932 571
rect 936 570 937 571
rect 942 571 948 572
rect 942 570 943 571
rect 936 568 943 570
rect 936 567 937 568
rect 931 566 937 567
rect 942 567 943 568
rect 947 567 948 571
rect 998 569 999 573
rect 1003 569 1004 573
rect 1086 573 1092 574
rect 998 568 1004 569
rect 1018 571 1025 572
rect 942 566 948 567
rect 1018 567 1019 571
rect 1024 567 1025 571
rect 1086 569 1087 573
rect 1091 569 1092 573
rect 1086 568 1092 569
rect 1107 573 1113 574
rect 1107 569 1108 573
rect 1112 569 1113 573
rect 1107 568 1113 569
rect 1182 573 1188 574
rect 1182 569 1183 573
rect 1187 569 1188 573
rect 1182 568 1188 569
rect 1203 573 1209 574
rect 1203 569 1204 573
rect 1208 569 1209 573
rect 1203 568 1209 569
rect 1286 572 1292 573
rect 1286 568 1287 572
rect 1291 568 1292 572
rect 1286 567 1292 568
rect 1326 571 1332 572
rect 1326 567 1327 571
rect 1331 567 1332 571
rect 2502 571 2508 572
rect 1018 566 1025 567
rect 1326 566 1332 567
rect 1366 568 1372 569
rect 1366 564 1367 568
rect 1371 564 1372 568
rect 1366 563 1372 564
rect 1446 568 1452 569
rect 1446 564 1447 568
rect 1451 564 1452 568
rect 1446 563 1452 564
rect 1534 568 1540 569
rect 1534 564 1535 568
rect 1539 564 1540 568
rect 1534 563 1540 564
rect 1630 568 1636 569
rect 1630 564 1631 568
rect 1635 564 1636 568
rect 1630 563 1636 564
rect 1726 568 1732 569
rect 1726 564 1727 568
rect 1731 564 1732 568
rect 1726 563 1732 564
rect 1830 568 1836 569
rect 1830 564 1831 568
rect 1835 564 1836 568
rect 1830 563 1836 564
rect 1942 568 1948 569
rect 1942 564 1943 568
rect 1947 564 1948 568
rect 1942 563 1948 564
rect 2062 568 2068 569
rect 2062 564 2063 568
rect 2067 564 2068 568
rect 2062 563 2068 564
rect 2190 568 2196 569
rect 2190 564 2191 568
rect 2195 564 2196 568
rect 2190 563 2196 564
rect 2326 568 2332 569
rect 2326 564 2327 568
rect 2331 564 2332 568
rect 2326 563 2332 564
rect 2438 568 2444 569
rect 2438 564 2439 568
rect 2443 564 2444 568
rect 2502 567 2503 571
rect 2507 567 2508 571
rect 2502 566 2508 567
rect 2438 563 2444 564
rect 1374 556 1380 557
rect 110 555 116 556
rect 110 551 111 555
rect 115 551 116 555
rect 1286 555 1292 556
rect 110 550 116 551
rect 134 552 140 553
rect 134 548 135 552
rect 139 548 140 552
rect 134 547 140 548
rect 222 552 228 553
rect 222 548 223 552
rect 227 548 228 552
rect 222 547 228 548
rect 318 552 324 553
rect 318 548 319 552
rect 323 548 324 552
rect 318 547 324 548
rect 414 552 420 553
rect 414 548 415 552
rect 419 548 420 552
rect 414 547 420 548
rect 518 552 524 553
rect 518 548 519 552
rect 523 548 524 552
rect 518 547 524 548
rect 614 552 620 553
rect 614 548 615 552
rect 619 548 620 552
rect 614 547 620 548
rect 710 552 716 553
rect 710 548 711 552
rect 715 548 716 552
rect 710 547 716 548
rect 806 552 812 553
rect 806 548 807 552
rect 811 548 812 552
rect 806 547 812 548
rect 894 552 900 553
rect 894 548 895 552
rect 899 548 900 552
rect 894 547 900 548
rect 982 552 988 553
rect 982 548 983 552
rect 987 548 988 552
rect 982 547 988 548
rect 1070 552 1076 553
rect 1070 548 1071 552
rect 1075 548 1076 552
rect 1070 547 1076 548
rect 1166 552 1172 553
rect 1166 548 1167 552
rect 1171 548 1172 552
rect 1286 551 1287 555
rect 1291 551 1292 555
rect 1286 550 1292 551
rect 1326 553 1332 554
rect 1326 549 1327 553
rect 1331 549 1332 553
rect 1374 552 1375 556
rect 1379 552 1380 556
rect 1374 551 1380 552
rect 1454 556 1460 557
rect 1454 552 1455 556
rect 1459 552 1460 556
rect 1454 551 1460 552
rect 1550 556 1556 557
rect 1550 552 1551 556
rect 1555 552 1556 556
rect 1550 551 1556 552
rect 1646 556 1652 557
rect 1646 552 1647 556
rect 1651 552 1652 556
rect 1646 551 1652 552
rect 1750 556 1756 557
rect 1750 552 1751 556
rect 1755 552 1756 556
rect 1750 551 1756 552
rect 1854 556 1860 557
rect 1854 552 1855 556
rect 1859 552 1860 556
rect 1854 551 1860 552
rect 1958 556 1964 557
rect 1958 552 1959 556
rect 1963 552 1964 556
rect 1958 551 1964 552
rect 2054 556 2060 557
rect 2054 552 2055 556
rect 2059 552 2060 556
rect 2054 551 2060 552
rect 2150 556 2156 557
rect 2150 552 2151 556
rect 2155 552 2156 556
rect 2150 551 2156 552
rect 2254 556 2260 557
rect 2254 552 2255 556
rect 2259 552 2260 556
rect 2254 551 2260 552
rect 2358 556 2364 557
rect 2358 552 2359 556
rect 2363 552 2364 556
rect 2358 551 2364 552
rect 2438 556 2444 557
rect 2438 552 2439 556
rect 2443 552 2444 556
rect 2438 551 2444 552
rect 2502 553 2508 554
rect 1326 548 1332 549
rect 2502 549 2503 553
rect 2507 549 2508 553
rect 2502 548 2508 549
rect 1166 547 1172 548
rect 1326 536 1332 537
rect 2502 536 2508 537
rect 142 532 148 533
rect 110 529 116 530
rect 110 525 111 529
rect 115 525 116 529
rect 142 528 143 532
rect 147 528 148 532
rect 142 527 148 528
rect 238 532 244 533
rect 238 528 239 532
rect 243 528 244 532
rect 238 527 244 528
rect 334 532 340 533
rect 334 528 335 532
rect 339 528 340 532
rect 334 527 340 528
rect 430 532 436 533
rect 430 528 431 532
rect 435 528 436 532
rect 430 527 436 528
rect 526 532 532 533
rect 526 528 527 532
rect 531 528 532 532
rect 526 527 532 528
rect 622 532 628 533
rect 622 528 623 532
rect 627 528 628 532
rect 622 527 628 528
rect 710 532 716 533
rect 710 528 711 532
rect 715 528 716 532
rect 710 527 716 528
rect 790 532 796 533
rect 790 528 791 532
rect 795 528 796 532
rect 790 527 796 528
rect 870 532 876 533
rect 870 528 871 532
rect 875 528 876 532
rect 870 527 876 528
rect 950 532 956 533
rect 950 528 951 532
rect 955 528 956 532
rect 950 527 956 528
rect 1030 532 1036 533
rect 1030 528 1031 532
rect 1035 528 1036 532
rect 1326 532 1327 536
rect 1331 532 1332 536
rect 1326 531 1332 532
rect 1390 535 1396 536
rect 1390 531 1391 535
rect 1395 531 1396 535
rect 1390 530 1396 531
rect 1411 535 1417 536
rect 1411 531 1412 535
rect 1416 534 1417 535
rect 1450 535 1456 536
rect 1450 534 1451 535
rect 1416 532 1451 534
rect 1416 531 1417 532
rect 1411 530 1417 531
rect 1450 531 1451 532
rect 1455 531 1456 535
rect 1450 530 1456 531
rect 1470 535 1476 536
rect 1470 531 1471 535
rect 1475 531 1476 535
rect 1470 530 1476 531
rect 1478 535 1484 536
rect 1478 531 1479 535
rect 1483 534 1484 535
rect 1491 535 1497 536
rect 1491 534 1492 535
rect 1483 532 1492 534
rect 1483 531 1484 532
rect 1478 530 1484 531
rect 1491 531 1492 532
rect 1496 531 1497 535
rect 1491 530 1497 531
rect 1566 535 1572 536
rect 1566 531 1567 535
rect 1571 531 1572 535
rect 1566 530 1572 531
rect 1586 535 1593 536
rect 1586 531 1587 535
rect 1592 531 1593 535
rect 1586 530 1593 531
rect 1662 535 1668 536
rect 1662 531 1663 535
rect 1667 531 1668 535
rect 1662 530 1668 531
rect 1683 535 1689 536
rect 1683 531 1684 535
rect 1688 531 1689 535
rect 1683 530 1689 531
rect 1766 535 1772 536
rect 1766 531 1767 535
rect 1771 531 1772 535
rect 1787 535 1793 536
rect 1787 534 1788 535
rect 1766 530 1772 531
rect 1776 532 1788 534
rect 1030 527 1036 528
rect 1286 529 1292 530
rect 110 524 116 525
rect 1286 525 1287 529
rect 1291 525 1292 529
rect 1286 524 1292 525
rect 1685 522 1687 530
rect 1776 522 1778 532
rect 1787 531 1788 532
rect 1792 531 1793 535
rect 1787 530 1793 531
rect 1870 535 1876 536
rect 1870 531 1871 535
rect 1875 531 1876 535
rect 1870 530 1876 531
rect 1890 535 1897 536
rect 1890 531 1891 535
rect 1896 531 1897 535
rect 1890 530 1897 531
rect 1974 535 1980 536
rect 1974 531 1975 535
rect 1979 531 1980 535
rect 1995 535 2001 536
rect 1995 534 1996 535
rect 1974 530 1980 531
rect 1984 532 1996 534
rect 1984 522 1986 532
rect 1995 531 1996 532
rect 2000 531 2001 535
rect 1995 530 2001 531
rect 2070 535 2076 536
rect 2070 531 2071 535
rect 2075 531 2076 535
rect 2070 530 2076 531
rect 2091 535 2097 536
rect 2091 531 2092 535
rect 2096 534 2097 535
rect 2146 535 2152 536
rect 2146 534 2147 535
rect 2096 532 2147 534
rect 2096 531 2097 532
rect 2091 530 2097 531
rect 2146 531 2147 532
rect 2151 531 2152 535
rect 2146 530 2152 531
rect 2166 535 2172 536
rect 2166 531 2167 535
rect 2171 531 2172 535
rect 2166 530 2172 531
rect 2187 535 2193 536
rect 2187 531 2188 535
rect 2192 534 2193 535
rect 2250 535 2256 536
rect 2250 534 2251 535
rect 2192 532 2251 534
rect 2192 531 2193 532
rect 2187 530 2193 531
rect 2250 531 2251 532
rect 2255 531 2256 535
rect 2250 530 2256 531
rect 2270 535 2276 536
rect 2270 531 2271 535
rect 2275 531 2276 535
rect 2270 530 2276 531
rect 2278 535 2284 536
rect 2278 531 2279 535
rect 2283 534 2284 535
rect 2291 535 2297 536
rect 2291 534 2292 535
rect 2283 532 2292 534
rect 2283 531 2284 532
rect 2278 530 2284 531
rect 2291 531 2292 532
rect 2296 531 2297 535
rect 2291 530 2297 531
rect 2374 535 2380 536
rect 2374 531 2375 535
rect 2379 531 2380 535
rect 2374 530 2380 531
rect 2390 535 2401 536
rect 2390 531 2391 535
rect 2395 531 2396 535
rect 2400 531 2401 535
rect 2390 530 2401 531
rect 2454 535 2460 536
rect 2454 531 2455 535
rect 2459 531 2460 535
rect 2454 530 2460 531
rect 2470 535 2481 536
rect 2470 531 2471 535
rect 2475 531 2476 535
rect 2480 531 2481 535
rect 2502 532 2503 536
rect 2507 532 2508 536
rect 2502 531 2508 532
rect 2470 530 2481 531
rect 2214 523 2220 524
rect 2214 522 2215 523
rect 1549 520 1687 522
rect 1720 520 1778 522
rect 1852 520 1986 522
rect 2053 520 2215 522
rect 1549 518 1551 520
rect 1720 518 1722 520
rect 1852 518 1854 520
rect 2053 518 2055 520
rect 2214 519 2215 520
rect 2219 519 2220 523
rect 2214 518 2220 519
rect 1547 517 1553 518
rect 1371 515 1377 516
rect 110 512 116 513
rect 1286 512 1292 513
rect 110 508 111 512
rect 115 508 116 512
rect 110 507 116 508
rect 158 511 164 512
rect 158 507 159 511
rect 163 507 164 511
rect 158 506 164 507
rect 179 511 185 512
rect 179 507 180 511
rect 184 510 185 511
rect 234 511 240 512
rect 234 510 235 511
rect 184 508 235 510
rect 184 507 185 508
rect 179 506 185 507
rect 234 507 235 508
rect 239 507 240 511
rect 234 506 240 507
rect 254 511 260 512
rect 254 507 255 511
rect 259 507 260 511
rect 254 506 260 507
rect 275 511 281 512
rect 275 507 276 511
rect 280 510 281 511
rect 286 511 292 512
rect 286 510 287 511
rect 280 508 287 510
rect 280 507 281 508
rect 275 506 281 507
rect 286 507 287 508
rect 291 507 292 511
rect 286 506 292 507
rect 350 511 356 512
rect 350 507 351 511
rect 355 507 356 511
rect 350 506 356 507
rect 371 511 377 512
rect 371 507 372 511
rect 376 510 377 511
rect 426 511 432 512
rect 426 510 427 511
rect 376 508 427 510
rect 376 507 377 508
rect 371 506 377 507
rect 426 507 427 508
rect 431 507 432 511
rect 426 506 432 507
rect 446 511 452 512
rect 446 507 447 511
rect 451 507 452 511
rect 446 506 452 507
rect 454 511 460 512
rect 454 507 455 511
rect 459 510 460 511
rect 467 511 473 512
rect 467 510 468 511
rect 459 508 468 510
rect 459 507 460 508
rect 454 506 460 507
rect 467 507 468 508
rect 472 507 473 511
rect 467 506 473 507
rect 542 511 548 512
rect 542 507 543 511
rect 547 507 548 511
rect 563 511 569 512
rect 563 510 564 511
rect 542 506 548 507
rect 552 508 564 510
rect 552 502 554 508
rect 563 507 564 508
rect 568 507 569 511
rect 563 506 569 507
rect 638 511 644 512
rect 638 507 639 511
rect 643 507 644 511
rect 638 506 644 507
rect 659 511 665 512
rect 659 507 660 511
rect 664 510 665 511
rect 706 511 712 512
rect 706 510 707 511
rect 664 508 707 510
rect 664 507 665 508
rect 659 506 665 507
rect 706 507 707 508
rect 711 507 712 511
rect 706 506 712 507
rect 726 511 732 512
rect 726 507 727 511
rect 731 507 732 511
rect 726 506 732 507
rect 742 511 753 512
rect 742 507 743 511
rect 747 507 748 511
rect 752 507 753 511
rect 742 506 753 507
rect 806 511 812 512
rect 806 507 807 511
rect 811 507 812 511
rect 806 506 812 507
rect 826 511 833 512
rect 826 507 827 511
rect 832 507 833 511
rect 826 506 833 507
rect 886 511 892 512
rect 886 507 887 511
rect 891 507 892 511
rect 907 511 913 512
rect 907 510 908 511
rect 886 506 892 507
rect 896 508 908 510
rect 332 500 554 502
rect 332 494 334 500
rect 646 499 652 500
rect 646 498 647 499
rect 524 496 647 498
rect 524 494 526 496
rect 646 495 647 496
rect 651 495 652 499
rect 896 498 898 508
rect 907 507 908 508
rect 912 507 913 511
rect 907 506 913 507
rect 966 511 972 512
rect 966 507 967 511
rect 971 507 972 511
rect 966 506 972 507
rect 987 511 993 512
rect 987 507 988 511
rect 992 510 993 511
rect 1026 511 1032 512
rect 1026 510 1027 511
rect 992 508 1027 510
rect 992 507 993 508
rect 987 506 993 507
rect 1026 507 1027 508
rect 1031 507 1032 511
rect 1026 506 1032 507
rect 1046 511 1052 512
rect 1046 507 1047 511
rect 1051 507 1052 511
rect 1067 511 1073 512
rect 1067 510 1068 511
rect 1046 506 1052 507
rect 1056 508 1068 510
rect 1056 498 1058 508
rect 1067 507 1068 508
rect 1072 507 1073 511
rect 1286 508 1287 512
rect 1291 508 1292 512
rect 1371 511 1372 515
rect 1376 514 1377 515
rect 1398 515 1404 516
rect 1398 514 1399 515
rect 1376 512 1399 514
rect 1376 511 1377 512
rect 1371 510 1377 511
rect 1398 511 1399 512
rect 1403 511 1404 515
rect 1398 510 1404 511
rect 1450 515 1457 516
rect 1450 511 1451 515
rect 1456 511 1457 515
rect 1547 513 1548 517
rect 1552 513 1553 517
rect 1547 512 1553 513
rect 1643 517 1722 518
rect 1643 513 1644 517
rect 1648 516 1722 517
rect 1851 517 1857 518
rect 1648 513 1649 516
rect 1643 512 1649 513
rect 1747 515 1753 516
rect 1450 510 1457 511
rect 1747 511 1748 515
rect 1752 514 1753 515
rect 1826 515 1832 516
rect 1826 514 1827 515
rect 1752 512 1827 514
rect 1752 511 1753 512
rect 1747 510 1753 511
rect 1826 511 1827 512
rect 1831 511 1832 515
rect 1851 513 1852 517
rect 1856 513 1857 517
rect 2051 517 2057 518
rect 1851 512 1857 513
rect 1942 515 1948 516
rect 1826 510 1832 511
rect 1942 511 1943 515
rect 1947 514 1948 515
rect 1955 515 1961 516
rect 1955 514 1956 515
rect 1947 512 1956 514
rect 1947 511 1948 512
rect 1942 510 1948 511
rect 1955 511 1956 512
rect 1960 511 1961 515
rect 2051 513 2052 517
rect 2056 513 2057 517
rect 2051 512 2057 513
rect 2146 515 2153 516
rect 1955 510 1961 511
rect 2146 511 2147 515
rect 2152 511 2153 515
rect 2146 510 2153 511
rect 2250 515 2257 516
rect 2250 511 2251 515
rect 2256 511 2257 515
rect 2250 510 2257 511
rect 2355 515 2361 516
rect 2355 511 2356 515
rect 2360 514 2361 515
rect 2414 515 2420 516
rect 2414 514 2415 515
rect 2360 512 2415 514
rect 2360 511 2361 512
rect 2355 510 2361 511
rect 2414 511 2415 512
rect 2419 511 2420 515
rect 2414 510 2420 511
rect 2435 515 2441 516
rect 2435 511 2436 515
rect 2440 514 2441 515
rect 2462 515 2468 516
rect 2462 514 2463 515
rect 2440 512 2463 514
rect 2440 511 2441 512
rect 2435 510 2441 511
rect 2462 511 2463 512
rect 2467 511 2468 515
rect 2462 510 2468 511
rect 1286 507 1292 508
rect 2390 507 2396 508
rect 1067 506 1073 507
rect 2390 506 2391 507
rect 2188 504 2391 506
rect 2188 502 2190 504
rect 2390 503 2391 504
rect 2395 503 2396 507
rect 2390 502 2396 503
rect 2187 501 2193 502
rect 646 494 652 495
rect 789 496 898 498
rect 900 496 1058 498
rect 1347 499 1353 500
rect 789 494 791 496
rect 900 494 902 496
rect 1347 495 1348 499
rect 1352 498 1353 499
rect 1435 499 1441 500
rect 1352 496 1430 498
rect 1352 495 1353 496
rect 1347 494 1353 495
rect 331 493 337 494
rect 139 491 145 492
rect 139 487 140 491
rect 144 490 145 491
rect 170 491 176 492
rect 170 490 171 491
rect 144 488 171 490
rect 144 487 145 488
rect 139 486 145 487
rect 170 487 171 488
rect 175 487 176 491
rect 170 486 176 487
rect 234 491 241 492
rect 234 487 235 491
rect 240 487 241 491
rect 331 489 332 493
rect 336 489 337 493
rect 523 493 529 494
rect 331 488 337 489
rect 426 491 433 492
rect 234 486 241 487
rect 426 487 427 491
rect 432 487 433 491
rect 523 489 524 493
rect 528 489 529 493
rect 787 493 793 494
rect 523 488 529 489
rect 619 491 625 492
rect 426 486 433 487
rect 619 487 620 491
rect 624 490 625 491
rect 674 491 680 492
rect 674 490 675 491
rect 624 488 675 490
rect 624 487 625 488
rect 619 486 625 487
rect 674 487 675 488
rect 679 487 680 491
rect 674 486 680 487
rect 706 491 713 492
rect 706 487 707 491
rect 712 487 713 491
rect 787 489 788 493
rect 792 489 793 493
rect 787 488 793 489
rect 867 493 902 494
rect 867 489 868 493
rect 872 492 902 493
rect 872 489 873 492
rect 867 488 873 489
rect 942 491 953 492
rect 706 486 713 487
rect 942 487 943 491
rect 947 487 948 491
rect 952 487 953 491
rect 942 486 953 487
rect 1026 491 1033 492
rect 1026 487 1027 491
rect 1032 487 1033 491
rect 1026 486 1033 487
rect 1428 486 1430 496
rect 1435 495 1436 499
rect 1440 498 1441 499
rect 1478 499 1484 500
rect 1478 498 1479 499
rect 1440 496 1479 498
rect 1440 495 1441 496
rect 1435 494 1441 495
rect 1478 495 1479 496
rect 1483 495 1484 499
rect 1478 494 1484 495
rect 1555 499 1561 500
rect 1555 495 1556 499
rect 1560 498 1561 499
rect 1598 499 1604 500
rect 1560 496 1594 498
rect 1560 495 1561 496
rect 1555 494 1561 495
rect 1592 490 1594 496
rect 1598 495 1599 499
rect 1603 498 1604 499
rect 1675 499 1681 500
rect 1675 498 1676 499
rect 1603 496 1676 498
rect 1603 495 1604 496
rect 1598 494 1604 495
rect 1675 495 1676 496
rect 1680 495 1681 499
rect 1675 494 1681 495
rect 1718 499 1724 500
rect 1718 495 1719 499
rect 1723 498 1724 499
rect 1787 499 1793 500
rect 1787 498 1788 499
rect 1723 496 1788 498
rect 1723 495 1724 496
rect 1718 494 1724 495
rect 1787 495 1788 496
rect 1792 495 1793 499
rect 1787 494 1793 495
rect 1899 499 1905 500
rect 1899 495 1900 499
rect 1904 498 1905 499
rect 1962 499 1968 500
rect 1962 498 1963 499
rect 1904 496 1963 498
rect 1904 495 1905 496
rect 1899 494 1905 495
rect 1962 495 1963 496
rect 1967 495 1968 499
rect 1962 494 1968 495
rect 2003 499 2009 500
rect 2003 495 2004 499
rect 2008 498 2009 499
rect 2046 499 2052 500
rect 2008 496 2042 498
rect 2008 495 2009 496
rect 2003 494 2009 495
rect 1618 491 1624 492
rect 1618 490 1619 491
rect 1592 488 1619 490
rect 1618 487 1619 488
rect 1623 487 1624 491
rect 1618 486 1624 487
rect 2040 486 2042 496
rect 2046 495 2047 499
rect 2051 498 2052 499
rect 2099 499 2105 500
rect 2099 498 2100 499
rect 2051 496 2100 498
rect 2051 495 2052 496
rect 2046 494 2052 495
rect 2099 495 2100 496
rect 2104 495 2105 499
rect 2187 497 2188 501
rect 2192 497 2193 501
rect 2187 496 2193 497
rect 2275 499 2284 500
rect 2099 494 2105 495
rect 2275 495 2276 499
rect 2283 495 2284 499
rect 2275 494 2284 495
rect 2314 499 2320 500
rect 2314 495 2315 499
rect 2319 498 2320 499
rect 2363 499 2369 500
rect 2363 498 2364 499
rect 2319 496 2364 498
rect 2319 495 2320 496
rect 2314 494 2320 495
rect 2363 495 2364 496
rect 2368 495 2369 499
rect 2363 494 2369 495
rect 2435 499 2441 500
rect 2435 495 2436 499
rect 2440 498 2441 499
rect 2446 499 2452 500
rect 2446 498 2447 499
rect 2440 496 2447 498
rect 2440 495 2441 496
rect 2435 494 2441 495
rect 2446 495 2447 496
rect 2451 495 2452 499
rect 2446 494 2452 495
rect 2414 487 2420 488
rect 1220 484 1391 486
rect 1428 484 1478 486
rect 2040 484 2230 486
rect 578 483 584 484
rect 578 482 579 483
rect 269 480 579 482
rect 269 478 271 480
rect 578 479 579 480
rect 583 479 584 483
rect 578 478 584 479
rect 1220 478 1222 484
rect 1389 482 1391 484
rect 1476 482 1478 484
rect 2228 482 2230 484
rect 2414 483 2415 487
rect 2419 486 2420 487
rect 2419 484 2479 486
rect 2419 483 2420 484
rect 2414 482 2420 483
rect 2477 482 2479 484
rect 1366 481 1372 482
rect 1326 480 1332 481
rect 267 477 273 478
rect 131 475 137 476
rect 131 471 132 475
rect 136 471 137 475
rect 131 470 137 471
rect 187 475 193 476
rect 187 471 188 475
rect 192 471 193 475
rect 267 473 268 477
rect 272 473 273 477
rect 1219 477 1225 478
rect 267 472 273 473
rect 310 475 316 476
rect 187 470 193 471
rect 302 471 308 472
rect 302 470 303 471
rect 133 462 135 470
rect 189 468 303 470
rect 302 467 303 468
rect 307 467 308 471
rect 310 471 311 475
rect 315 474 316 475
rect 355 475 361 476
rect 355 474 356 475
rect 315 472 356 474
rect 315 471 316 472
rect 310 470 316 471
rect 355 471 356 472
rect 360 471 361 475
rect 355 470 361 471
rect 443 475 449 476
rect 443 471 444 475
rect 448 474 449 475
rect 454 475 460 476
rect 454 474 455 475
rect 448 472 455 474
rect 448 471 449 472
rect 443 470 449 471
rect 454 471 455 472
rect 459 471 460 475
rect 454 470 460 471
rect 486 475 492 476
rect 486 471 487 475
rect 491 474 492 475
rect 539 475 545 476
rect 539 474 540 475
rect 491 472 540 474
rect 491 471 492 472
rect 486 470 492 471
rect 539 471 540 472
rect 544 471 545 475
rect 539 470 545 471
rect 635 475 641 476
rect 635 471 636 475
rect 640 474 641 475
rect 731 475 737 476
rect 640 472 726 474
rect 640 471 641 472
rect 635 470 641 471
rect 302 466 308 467
rect 724 462 726 472
rect 731 471 732 475
rect 736 474 737 475
rect 742 475 748 476
rect 742 474 743 475
rect 736 472 743 474
rect 736 471 737 472
rect 731 470 737 471
rect 742 471 743 472
rect 747 471 748 475
rect 742 470 748 471
rect 826 475 833 476
rect 826 471 827 475
rect 832 471 833 475
rect 826 470 833 471
rect 870 475 876 476
rect 870 471 871 475
rect 875 474 876 475
rect 931 475 937 476
rect 931 474 932 475
rect 875 472 932 474
rect 875 471 876 472
rect 870 470 876 471
rect 931 471 932 472
rect 936 471 937 475
rect 931 470 937 471
rect 974 475 980 476
rect 974 471 975 475
rect 979 474 980 475
rect 1035 475 1041 476
rect 1035 474 1036 475
rect 979 472 1036 474
rect 979 471 980 472
rect 974 470 980 471
rect 1035 471 1036 472
rect 1040 471 1041 475
rect 1035 470 1041 471
rect 1139 475 1145 476
rect 1139 471 1140 475
rect 1144 474 1145 475
rect 1144 472 1161 474
rect 1219 473 1220 477
rect 1224 473 1225 477
rect 1326 476 1327 480
rect 1331 476 1332 480
rect 1366 477 1367 481
rect 1371 477 1372 481
rect 1366 476 1372 477
rect 1387 481 1393 482
rect 1387 477 1388 481
rect 1392 477 1393 481
rect 1387 476 1393 477
rect 1454 481 1460 482
rect 1454 477 1455 481
rect 1459 477 1460 481
rect 1454 476 1460 477
rect 1475 481 1481 482
rect 1475 477 1476 481
rect 1480 477 1481 481
rect 1475 476 1481 477
rect 1574 481 1580 482
rect 1574 477 1575 481
rect 1579 477 1580 481
rect 1694 481 1700 482
rect 1574 476 1580 477
rect 1595 479 1604 480
rect 1326 475 1332 476
rect 1595 475 1596 479
rect 1603 475 1604 479
rect 1694 477 1695 481
rect 1699 477 1700 481
rect 1806 481 1812 482
rect 1694 476 1700 477
rect 1715 479 1724 480
rect 1595 474 1604 475
rect 1715 475 1716 479
rect 1723 475 1724 479
rect 1806 477 1807 481
rect 1811 477 1812 481
rect 1918 481 1924 482
rect 1806 476 1812 477
rect 1826 479 1833 480
rect 1715 474 1724 475
rect 1826 475 1827 479
rect 1832 475 1833 479
rect 1918 477 1919 481
rect 1923 477 1924 481
rect 2022 481 2028 482
rect 1918 476 1924 477
rect 1939 479 1948 480
rect 1826 474 1833 475
rect 1939 475 1940 479
rect 1947 475 1948 479
rect 2022 477 2023 481
rect 2027 477 2028 481
rect 2118 481 2124 482
rect 2022 476 2028 477
rect 2043 479 2052 480
rect 1939 474 1948 475
rect 2043 475 2044 479
rect 2051 475 2052 479
rect 2118 477 2119 481
rect 2123 477 2124 481
rect 2206 481 2212 482
rect 2118 476 2124 477
rect 2139 479 2145 480
rect 2043 474 2052 475
rect 2139 475 2140 479
rect 2144 478 2145 479
rect 2166 479 2172 480
rect 2166 478 2167 479
rect 2144 476 2167 478
rect 2144 475 2145 476
rect 2139 474 2145 475
rect 2166 475 2167 476
rect 2171 475 2172 479
rect 2206 477 2207 481
rect 2211 477 2212 481
rect 2206 476 2212 477
rect 2227 481 2233 482
rect 2227 477 2228 481
rect 2232 477 2233 481
rect 2227 476 2233 477
rect 2294 481 2300 482
rect 2294 477 2295 481
rect 2299 477 2300 481
rect 2382 481 2388 482
rect 2294 476 2300 477
rect 2314 479 2321 480
rect 2166 474 2172 475
rect 2314 475 2315 479
rect 2320 475 2321 479
rect 2382 477 2383 481
rect 2387 477 2388 481
rect 2454 481 2460 482
rect 2382 476 2388 477
rect 2398 479 2409 480
rect 2314 474 2321 475
rect 2398 475 2399 479
rect 2403 475 2404 479
rect 2408 475 2409 479
rect 2454 477 2455 481
rect 2459 477 2460 481
rect 2454 476 2460 477
rect 2475 481 2481 482
rect 2475 477 2476 481
rect 2480 477 2481 481
rect 2475 476 2481 477
rect 2502 480 2508 481
rect 2502 476 2503 480
rect 2507 476 2508 480
rect 2502 475 2508 476
rect 2398 474 2409 475
rect 1219 472 1225 473
rect 1144 471 1145 472
rect 1139 470 1145 471
rect 838 463 844 464
rect 133 460 230 462
rect 724 460 766 462
rect 228 458 230 460
rect 764 458 766 460
rect 838 459 839 463
rect 843 462 844 463
rect 1159 462 1161 472
rect 1326 463 1332 464
rect 843 460 1079 462
rect 1159 460 1263 462
rect 843 459 844 460
rect 838 458 844 459
rect 1077 458 1079 460
rect 1261 458 1263 460
rect 1326 459 1327 463
rect 1331 459 1332 463
rect 2502 463 2508 464
rect 1326 458 1332 459
rect 1350 460 1356 461
rect 150 457 156 458
rect 110 456 116 457
rect 110 452 111 456
rect 115 452 116 456
rect 150 453 151 457
rect 155 453 156 457
rect 206 457 212 458
rect 150 452 156 453
rect 170 455 177 456
rect 110 451 116 452
rect 170 451 171 455
rect 176 451 177 455
rect 206 453 207 457
rect 211 453 212 457
rect 206 452 212 453
rect 227 457 233 458
rect 227 453 228 457
rect 232 453 233 457
rect 227 452 233 453
rect 286 457 292 458
rect 286 453 287 457
rect 291 453 292 457
rect 374 457 380 458
rect 286 452 292 453
rect 307 455 316 456
rect 170 450 177 451
rect 307 451 308 455
rect 315 451 316 455
rect 374 453 375 457
rect 379 453 380 457
rect 462 457 468 458
rect 374 452 380 453
rect 390 455 401 456
rect 307 450 316 451
rect 390 451 391 455
rect 395 451 396 455
rect 400 451 401 455
rect 462 453 463 457
rect 467 453 468 457
rect 558 457 564 458
rect 462 452 468 453
rect 483 455 492 456
rect 390 450 401 451
rect 483 451 484 455
rect 491 451 492 455
rect 558 453 559 457
rect 563 453 564 457
rect 654 457 660 458
rect 558 452 564 453
rect 578 455 585 456
rect 483 450 492 451
rect 578 451 579 455
rect 584 451 585 455
rect 654 453 655 457
rect 659 453 660 457
rect 750 457 756 458
rect 654 452 660 453
rect 674 455 681 456
rect 578 450 585 451
rect 674 451 675 455
rect 680 451 681 455
rect 750 453 751 457
rect 755 453 756 457
rect 764 457 777 458
rect 764 456 772 457
rect 750 452 756 453
rect 771 453 772 456
rect 776 453 777 457
rect 771 452 777 453
rect 846 457 852 458
rect 846 453 847 457
rect 851 453 852 457
rect 950 457 956 458
rect 846 452 852 453
rect 867 455 876 456
rect 674 450 681 451
rect 867 451 868 455
rect 875 451 876 455
rect 950 453 951 457
rect 955 453 956 457
rect 1054 457 1060 458
rect 950 452 956 453
rect 971 455 980 456
rect 867 450 876 451
rect 971 451 972 455
rect 979 451 980 455
rect 1054 453 1055 457
rect 1059 453 1060 457
rect 1054 452 1060 453
rect 1075 457 1081 458
rect 1075 453 1076 457
rect 1080 453 1081 457
rect 1075 452 1081 453
rect 1158 457 1164 458
rect 1158 453 1159 457
rect 1163 453 1164 457
rect 1238 457 1244 458
rect 1158 452 1164 453
rect 1166 455 1172 456
rect 971 450 980 451
rect 1166 451 1167 455
rect 1171 454 1172 455
rect 1179 455 1185 456
rect 1179 454 1180 455
rect 1171 452 1180 454
rect 1171 451 1172 452
rect 1166 450 1172 451
rect 1179 451 1180 452
rect 1184 451 1185 455
rect 1238 453 1239 457
rect 1243 453 1244 457
rect 1238 452 1244 453
rect 1259 457 1265 458
rect 1259 453 1260 457
rect 1264 453 1265 457
rect 1259 452 1265 453
rect 1286 456 1292 457
rect 1286 452 1287 456
rect 1291 452 1292 456
rect 1350 456 1351 460
rect 1355 456 1356 460
rect 1350 455 1356 456
rect 1438 460 1444 461
rect 1438 456 1439 460
rect 1443 456 1444 460
rect 1438 455 1444 456
rect 1558 460 1564 461
rect 1558 456 1559 460
rect 1563 456 1564 460
rect 1558 455 1564 456
rect 1678 460 1684 461
rect 1678 456 1679 460
rect 1683 456 1684 460
rect 1678 455 1684 456
rect 1790 460 1796 461
rect 1790 456 1791 460
rect 1795 456 1796 460
rect 1790 455 1796 456
rect 1902 460 1908 461
rect 1902 456 1903 460
rect 1907 456 1908 460
rect 1902 455 1908 456
rect 2006 460 2012 461
rect 2006 456 2007 460
rect 2011 456 2012 460
rect 2006 455 2012 456
rect 2102 460 2108 461
rect 2102 456 2103 460
rect 2107 456 2108 460
rect 2102 455 2108 456
rect 2190 460 2196 461
rect 2190 456 2191 460
rect 2195 456 2196 460
rect 2190 455 2196 456
rect 2278 460 2284 461
rect 2278 456 2279 460
rect 2283 456 2284 460
rect 2278 455 2284 456
rect 2366 460 2372 461
rect 2366 456 2367 460
rect 2371 456 2372 460
rect 2366 455 2372 456
rect 2438 460 2444 461
rect 2438 456 2439 460
rect 2443 456 2444 460
rect 2502 459 2503 463
rect 2507 459 2508 463
rect 2502 458 2508 459
rect 2438 455 2444 456
rect 1286 451 1292 452
rect 1179 450 1185 451
rect 110 439 116 440
rect 110 435 111 439
rect 115 435 116 439
rect 1286 439 1292 440
rect 110 434 116 435
rect 134 436 140 437
rect 134 432 135 436
rect 139 432 140 436
rect 134 431 140 432
rect 190 436 196 437
rect 190 432 191 436
rect 195 432 196 436
rect 190 431 196 432
rect 270 436 276 437
rect 270 432 271 436
rect 275 432 276 436
rect 270 431 276 432
rect 358 436 364 437
rect 358 432 359 436
rect 363 432 364 436
rect 358 431 364 432
rect 446 436 452 437
rect 446 432 447 436
rect 451 432 452 436
rect 446 431 452 432
rect 542 436 548 437
rect 542 432 543 436
rect 547 432 548 436
rect 542 431 548 432
rect 638 436 644 437
rect 638 432 639 436
rect 643 432 644 436
rect 638 431 644 432
rect 734 436 740 437
rect 734 432 735 436
rect 739 432 740 436
rect 734 431 740 432
rect 830 436 836 437
rect 830 432 831 436
rect 835 432 836 436
rect 830 431 836 432
rect 934 436 940 437
rect 934 432 935 436
rect 939 432 940 436
rect 934 431 940 432
rect 1038 436 1044 437
rect 1038 432 1039 436
rect 1043 432 1044 436
rect 1038 431 1044 432
rect 1142 436 1148 437
rect 1142 432 1143 436
rect 1147 432 1148 436
rect 1142 431 1148 432
rect 1222 436 1228 437
rect 1222 432 1223 436
rect 1227 432 1228 436
rect 1286 435 1287 439
rect 1291 435 1292 439
rect 1286 434 1292 435
rect 1582 436 1588 437
rect 1222 431 1228 432
rect 1326 433 1332 434
rect 1326 429 1327 433
rect 1331 429 1332 433
rect 1582 432 1583 436
rect 1587 432 1588 436
rect 1582 431 1588 432
rect 1638 436 1644 437
rect 1638 432 1639 436
rect 1643 432 1644 436
rect 1638 431 1644 432
rect 1694 436 1700 437
rect 1694 432 1695 436
rect 1699 432 1700 436
rect 1694 431 1700 432
rect 1758 436 1764 437
rect 1758 432 1759 436
rect 1763 432 1764 436
rect 1758 431 1764 432
rect 1830 436 1836 437
rect 1830 432 1831 436
rect 1835 432 1836 436
rect 1830 431 1836 432
rect 1910 436 1916 437
rect 1910 432 1911 436
rect 1915 432 1916 436
rect 1910 431 1916 432
rect 1990 436 1996 437
rect 1990 432 1991 436
rect 1995 432 1996 436
rect 1990 431 1996 432
rect 2078 436 2084 437
rect 2078 432 2079 436
rect 2083 432 2084 436
rect 2078 431 2084 432
rect 2174 436 2180 437
rect 2174 432 2175 436
rect 2179 432 2180 436
rect 2174 431 2180 432
rect 2270 436 2276 437
rect 2270 432 2271 436
rect 2275 432 2276 436
rect 2270 431 2276 432
rect 2366 436 2372 437
rect 2366 432 2367 436
rect 2371 432 2372 436
rect 2366 431 2372 432
rect 2438 436 2444 437
rect 2438 432 2439 436
rect 2443 432 2444 436
rect 2438 431 2444 432
rect 2502 433 2508 434
rect 1326 428 1332 429
rect 2502 429 2503 433
rect 2507 429 2508 433
rect 2502 428 2508 429
rect 134 424 140 425
rect 110 421 116 422
rect 110 417 111 421
rect 115 417 116 421
rect 134 420 135 424
rect 139 420 140 424
rect 134 419 140 420
rect 190 424 196 425
rect 190 420 191 424
rect 195 420 196 424
rect 190 419 196 420
rect 278 424 284 425
rect 278 420 279 424
rect 283 420 284 424
rect 278 419 284 420
rect 382 424 388 425
rect 382 420 383 424
rect 387 420 388 424
rect 382 419 388 420
rect 494 424 500 425
rect 494 420 495 424
rect 499 420 500 424
rect 494 419 500 420
rect 606 424 612 425
rect 606 420 607 424
rect 611 420 612 424
rect 606 419 612 420
rect 718 424 724 425
rect 718 420 719 424
rect 723 420 724 424
rect 718 419 724 420
rect 830 424 836 425
rect 830 420 831 424
rect 835 420 836 424
rect 830 419 836 420
rect 934 424 940 425
rect 934 420 935 424
rect 939 420 940 424
rect 934 419 940 420
rect 1038 424 1044 425
rect 1038 420 1039 424
rect 1043 420 1044 424
rect 1038 419 1044 420
rect 1142 424 1148 425
rect 1142 420 1143 424
rect 1147 420 1148 424
rect 1142 419 1148 420
rect 1222 424 1228 425
rect 1222 420 1223 424
rect 1227 420 1228 424
rect 1222 419 1228 420
rect 1286 421 1292 422
rect 110 416 116 417
rect 1286 417 1287 421
rect 1291 417 1292 421
rect 1286 416 1292 417
rect 1326 416 1332 417
rect 2502 416 2508 417
rect 1326 412 1327 416
rect 1331 412 1332 416
rect 1326 411 1332 412
rect 1598 415 1604 416
rect 1598 411 1599 415
rect 1603 411 1604 415
rect 1598 410 1604 411
rect 1618 415 1625 416
rect 1618 411 1619 415
rect 1624 411 1625 415
rect 1618 410 1625 411
rect 1654 415 1660 416
rect 1654 411 1655 415
rect 1659 411 1660 415
rect 1675 415 1681 416
rect 1675 414 1676 415
rect 1654 410 1660 411
rect 1664 412 1676 414
rect 1664 406 1666 412
rect 1675 411 1676 412
rect 1680 411 1681 415
rect 1675 410 1681 411
rect 1710 415 1716 416
rect 1710 411 1711 415
rect 1715 411 1716 415
rect 1731 415 1737 416
rect 1731 414 1732 415
rect 1710 410 1716 411
rect 1720 412 1732 414
rect 110 404 116 405
rect 1286 404 1292 405
rect 110 400 111 404
rect 115 400 116 404
rect 110 399 116 400
rect 150 403 156 404
rect 150 399 151 403
rect 155 399 156 403
rect 150 398 156 399
rect 171 403 177 404
rect 171 399 172 403
rect 176 402 177 403
rect 186 403 192 404
rect 186 402 187 403
rect 176 400 187 402
rect 176 399 177 400
rect 171 398 177 399
rect 186 399 187 400
rect 191 399 192 403
rect 186 398 192 399
rect 206 403 212 404
rect 206 399 207 403
rect 211 399 212 403
rect 206 398 212 399
rect 227 403 233 404
rect 227 399 228 403
rect 232 402 233 403
rect 274 403 280 404
rect 274 402 275 403
rect 232 400 275 402
rect 232 399 233 400
rect 227 398 233 399
rect 274 399 275 400
rect 279 399 280 403
rect 274 398 280 399
rect 294 403 300 404
rect 294 399 295 403
rect 299 399 300 403
rect 294 398 300 399
rect 302 403 308 404
rect 302 399 303 403
rect 307 402 308 403
rect 315 403 321 404
rect 315 402 316 403
rect 307 400 316 402
rect 307 399 308 400
rect 302 398 308 399
rect 315 399 316 400
rect 320 399 321 403
rect 315 398 321 399
rect 398 403 404 404
rect 398 399 399 403
rect 403 399 404 403
rect 398 398 404 399
rect 419 403 425 404
rect 419 399 420 403
rect 424 402 425 403
rect 490 403 496 404
rect 490 402 491 403
rect 424 400 491 402
rect 424 399 425 400
rect 419 398 425 399
rect 490 399 491 400
rect 495 399 496 403
rect 490 398 496 399
rect 510 403 516 404
rect 510 399 511 403
rect 515 399 516 403
rect 510 398 516 399
rect 531 403 537 404
rect 531 399 532 403
rect 536 402 537 403
rect 602 403 608 404
rect 602 402 603 403
rect 536 400 603 402
rect 536 399 537 400
rect 531 398 537 399
rect 602 399 603 400
rect 607 399 608 403
rect 602 398 608 399
rect 622 403 628 404
rect 622 399 623 403
rect 627 399 628 403
rect 622 398 628 399
rect 630 403 636 404
rect 630 399 631 403
rect 635 402 636 403
rect 643 403 649 404
rect 643 402 644 403
rect 635 400 644 402
rect 635 399 636 400
rect 630 398 636 399
rect 643 399 644 400
rect 648 399 649 403
rect 643 398 649 399
rect 734 403 740 404
rect 734 399 735 403
rect 739 399 740 403
rect 734 398 740 399
rect 742 403 748 404
rect 742 399 743 403
rect 747 402 748 403
rect 755 403 761 404
rect 755 402 756 403
rect 747 400 756 402
rect 747 399 748 400
rect 742 398 748 399
rect 755 399 756 400
rect 760 399 761 403
rect 755 398 761 399
rect 846 403 852 404
rect 846 399 847 403
rect 851 399 852 403
rect 846 398 852 399
rect 867 403 873 404
rect 867 399 868 403
rect 872 402 873 403
rect 930 403 936 404
rect 930 402 931 403
rect 872 400 931 402
rect 872 399 873 400
rect 867 398 873 399
rect 930 399 931 400
rect 935 399 936 403
rect 930 398 936 399
rect 950 403 956 404
rect 950 399 951 403
rect 955 399 956 403
rect 950 398 956 399
rect 971 403 977 404
rect 971 399 972 403
rect 976 402 977 403
rect 994 403 1000 404
rect 994 402 995 403
rect 976 400 995 402
rect 976 399 977 400
rect 971 398 977 399
rect 994 399 995 400
rect 999 399 1000 403
rect 994 398 1000 399
rect 1054 403 1060 404
rect 1054 399 1055 403
rect 1059 399 1060 403
rect 1054 398 1060 399
rect 1074 403 1081 404
rect 1074 399 1075 403
rect 1080 399 1081 403
rect 1074 398 1081 399
rect 1158 403 1164 404
rect 1158 399 1159 403
rect 1163 399 1164 403
rect 1158 398 1164 399
rect 1179 403 1185 404
rect 1179 399 1180 403
rect 1184 402 1185 403
rect 1218 403 1224 404
rect 1218 402 1219 403
rect 1184 400 1219 402
rect 1184 399 1185 400
rect 1179 398 1185 399
rect 1218 399 1219 400
rect 1223 399 1224 403
rect 1218 398 1224 399
rect 1238 403 1244 404
rect 1238 399 1239 403
rect 1243 399 1244 403
rect 1238 398 1244 399
rect 1259 403 1265 404
rect 1259 399 1260 403
rect 1264 399 1265 403
rect 1286 400 1287 404
rect 1291 400 1292 404
rect 1286 399 1292 400
rect 1580 404 1666 406
rect 1259 398 1265 399
rect 1580 398 1582 404
rect 1720 402 1722 412
rect 1731 411 1732 412
rect 1736 411 1737 415
rect 1731 410 1737 411
rect 1774 415 1780 416
rect 1774 411 1775 415
rect 1779 411 1780 415
rect 1795 415 1801 416
rect 1795 414 1796 415
rect 1774 410 1780 411
rect 1784 412 1796 414
rect 1784 402 1786 412
rect 1795 411 1796 412
rect 1800 411 1801 415
rect 1795 410 1801 411
rect 1846 415 1852 416
rect 1846 411 1847 415
rect 1851 411 1852 415
rect 1867 415 1873 416
rect 1867 414 1868 415
rect 1846 410 1852 411
rect 1856 412 1868 414
rect 1856 406 1858 412
rect 1867 411 1868 412
rect 1872 411 1873 415
rect 1867 410 1873 411
rect 1926 415 1932 416
rect 1926 411 1927 415
rect 1931 411 1932 415
rect 1926 410 1932 411
rect 1947 415 1953 416
rect 1947 411 1948 415
rect 1952 414 1953 415
rect 1986 415 1992 416
rect 1986 414 1987 415
rect 1952 412 1987 414
rect 1952 411 1953 412
rect 1947 410 1953 411
rect 1986 411 1987 412
rect 1991 411 1992 415
rect 1986 410 1992 411
rect 2006 415 2012 416
rect 2006 411 2007 415
rect 2011 411 2012 415
rect 2006 410 2012 411
rect 2027 415 2033 416
rect 2027 411 2028 415
rect 2032 414 2033 415
rect 2074 415 2080 416
rect 2074 414 2075 415
rect 2032 412 2075 414
rect 2032 411 2033 412
rect 2027 410 2033 411
rect 2074 411 2075 412
rect 2079 411 2080 415
rect 2074 410 2080 411
rect 2094 415 2100 416
rect 2094 411 2095 415
rect 2099 411 2100 415
rect 2094 410 2100 411
rect 2102 415 2108 416
rect 2102 411 2103 415
rect 2107 414 2108 415
rect 2115 415 2121 416
rect 2115 414 2116 415
rect 2107 412 2116 414
rect 2107 411 2108 412
rect 2102 410 2108 411
rect 2115 411 2116 412
rect 2120 411 2121 415
rect 2115 410 2121 411
rect 2190 415 2196 416
rect 2190 411 2191 415
rect 2195 411 2196 415
rect 2190 410 2196 411
rect 2211 415 2217 416
rect 2211 411 2212 415
rect 2216 414 2217 415
rect 2266 415 2272 416
rect 2266 414 2267 415
rect 2216 412 2267 414
rect 2216 411 2217 412
rect 2211 410 2217 411
rect 2266 411 2267 412
rect 2271 411 2272 415
rect 2266 410 2272 411
rect 2286 415 2292 416
rect 2286 411 2287 415
rect 2291 411 2292 415
rect 2286 410 2292 411
rect 2294 415 2300 416
rect 2294 411 2295 415
rect 2299 414 2300 415
rect 2307 415 2313 416
rect 2307 414 2308 415
rect 2299 412 2308 414
rect 2299 411 2300 412
rect 2294 410 2300 411
rect 2307 411 2308 412
rect 2312 411 2313 415
rect 2307 410 2313 411
rect 2382 415 2388 416
rect 2382 411 2383 415
rect 2387 411 2388 415
rect 2382 410 2388 411
rect 2390 415 2396 416
rect 2390 411 2391 415
rect 2395 414 2396 415
rect 2403 415 2409 416
rect 2403 414 2404 415
rect 2395 412 2404 414
rect 2395 411 2396 412
rect 2390 410 2396 411
rect 2403 411 2404 412
rect 2408 411 2409 415
rect 2403 410 2409 411
rect 2454 415 2460 416
rect 2454 411 2455 415
rect 2459 411 2460 415
rect 2454 410 2460 411
rect 2462 415 2468 416
rect 2462 411 2463 415
rect 2467 414 2468 415
rect 2475 415 2481 416
rect 2475 414 2476 415
rect 2467 412 2476 414
rect 2467 411 2468 412
rect 2462 410 2468 411
rect 2475 411 2476 412
rect 2480 411 2481 415
rect 2502 412 2503 416
rect 2507 412 2508 416
rect 2502 411 2508 412
rect 2475 410 2481 411
rect 1636 400 1722 402
rect 1728 400 1786 402
rect 1788 404 1858 406
rect 1636 398 1638 400
rect 1728 398 1730 400
rect 1788 398 1790 404
rect 1261 390 1263 398
rect 1579 397 1585 398
rect 1579 393 1580 397
rect 1584 393 1585 397
rect 1579 392 1585 393
rect 1635 397 1641 398
rect 1635 393 1636 397
rect 1640 393 1641 397
rect 1635 392 1641 393
rect 1691 397 1730 398
rect 1691 393 1692 397
rect 1696 396 1730 397
rect 1755 397 1790 398
rect 1696 393 1697 396
rect 1691 392 1697 393
rect 1755 393 1756 397
rect 1760 396 1790 397
rect 1760 393 1761 396
rect 1755 392 1761 393
rect 1827 395 1833 396
rect 1827 391 1828 395
rect 1832 394 1833 395
rect 1886 395 1892 396
rect 1886 394 1887 395
rect 1832 392 1887 394
rect 1832 391 1833 392
rect 1827 390 1833 391
rect 1886 391 1887 392
rect 1891 391 1892 395
rect 1886 390 1892 391
rect 1894 395 1900 396
rect 1894 391 1895 395
rect 1899 394 1900 395
rect 1907 395 1913 396
rect 1907 394 1908 395
rect 1899 392 1908 394
rect 1899 391 1900 392
rect 1894 390 1900 391
rect 1907 391 1908 392
rect 1912 391 1913 395
rect 1907 390 1913 391
rect 1986 395 1993 396
rect 1986 391 1987 395
rect 1992 391 1993 395
rect 1986 390 1993 391
rect 2074 395 2081 396
rect 2074 391 2075 395
rect 2080 391 2081 395
rect 2074 390 2081 391
rect 2166 395 2177 396
rect 2166 391 2167 395
rect 2171 391 2172 395
rect 2176 391 2177 395
rect 2166 390 2177 391
rect 2266 395 2273 396
rect 2266 391 2267 395
rect 2272 391 2273 395
rect 2266 390 2273 391
rect 2363 395 2369 396
rect 2363 391 2364 395
rect 2368 394 2369 395
rect 2398 395 2404 396
rect 2398 394 2399 395
rect 2368 392 2399 394
rect 2368 391 2369 392
rect 2363 390 2369 391
rect 2398 391 2399 392
rect 2403 391 2404 395
rect 2398 390 2404 391
rect 2435 395 2441 396
rect 2435 391 2436 395
rect 2440 394 2441 395
rect 2470 395 2476 396
rect 2470 394 2471 395
rect 2440 392 2471 394
rect 2440 391 2441 392
rect 2435 390 2441 391
rect 2470 391 2471 392
rect 2475 391 2476 395
rect 2470 390 2476 391
rect 1036 388 1263 390
rect 1036 386 1038 388
rect 1035 385 1041 386
rect 131 383 137 384
rect 131 379 132 383
rect 136 382 137 383
rect 170 383 176 384
rect 170 382 171 383
rect 136 380 171 382
rect 136 379 137 380
rect 131 378 137 379
rect 170 379 171 380
rect 175 379 176 383
rect 170 378 176 379
rect 186 383 193 384
rect 186 379 187 383
rect 192 379 193 383
rect 186 378 193 379
rect 274 383 281 384
rect 274 379 275 383
rect 280 379 281 383
rect 274 378 281 379
rect 379 383 385 384
rect 379 379 380 383
rect 384 382 385 383
rect 390 383 396 384
rect 390 382 391 383
rect 384 380 391 382
rect 384 379 385 380
rect 379 378 385 379
rect 390 379 391 380
rect 395 379 396 383
rect 390 378 396 379
rect 490 383 497 384
rect 490 379 491 383
rect 496 379 497 383
rect 490 378 497 379
rect 602 383 609 384
rect 602 379 603 383
rect 608 379 609 383
rect 602 378 609 379
rect 715 383 721 384
rect 715 379 716 383
rect 720 382 721 383
rect 770 383 776 384
rect 770 382 771 383
rect 720 380 771 382
rect 720 379 721 380
rect 715 378 721 379
rect 770 379 771 380
rect 775 379 776 383
rect 770 378 776 379
rect 827 383 833 384
rect 827 379 828 383
rect 832 382 833 383
rect 838 383 844 384
rect 838 382 839 383
rect 832 380 839 382
rect 832 379 833 380
rect 827 378 833 379
rect 838 379 839 380
rect 843 379 844 383
rect 838 378 844 379
rect 930 383 937 384
rect 930 379 931 383
rect 936 379 937 383
rect 1035 381 1036 385
rect 1040 381 1041 385
rect 1035 380 1041 381
rect 1139 383 1145 384
rect 930 378 937 379
rect 1139 379 1140 383
rect 1144 382 1145 383
rect 1166 383 1172 384
rect 1166 382 1167 383
rect 1144 380 1167 382
rect 1144 379 1145 380
rect 1139 378 1145 379
rect 1166 379 1167 380
rect 1171 379 1172 383
rect 1166 378 1172 379
rect 1218 383 1225 384
rect 1218 379 1219 383
rect 1224 379 1225 383
rect 1218 378 1225 379
rect 1622 379 1628 380
rect 630 375 636 376
rect 630 374 631 375
rect 319 372 631 374
rect 319 370 321 372
rect 630 371 631 372
rect 635 371 636 375
rect 1622 375 1623 379
rect 1627 378 1628 379
rect 1659 379 1665 380
rect 1659 378 1660 379
rect 1627 376 1660 378
rect 1627 375 1628 376
rect 1622 374 1628 375
rect 1659 375 1660 376
rect 1664 375 1665 379
rect 1659 374 1665 375
rect 1702 379 1708 380
rect 1702 375 1703 379
rect 1707 378 1708 379
rect 1715 379 1721 380
rect 1715 378 1716 379
rect 1707 376 1716 378
rect 1707 375 1708 376
rect 1702 374 1708 375
rect 1715 375 1716 376
rect 1720 375 1721 379
rect 1715 374 1721 375
rect 1758 379 1764 380
rect 1758 375 1759 379
rect 1763 378 1764 379
rect 1779 379 1785 380
rect 1779 378 1780 379
rect 1763 376 1780 378
rect 1763 375 1764 376
rect 1758 374 1764 375
rect 1779 375 1780 376
rect 1784 375 1785 379
rect 1779 374 1785 375
rect 1822 379 1828 380
rect 1822 375 1823 379
rect 1827 378 1828 379
rect 1851 379 1857 380
rect 1851 378 1852 379
rect 1827 376 1852 378
rect 1827 375 1828 376
rect 1822 374 1828 375
rect 1851 375 1852 376
rect 1856 375 1857 379
rect 1851 374 1857 375
rect 1878 379 1884 380
rect 1878 375 1879 379
rect 1883 378 1884 379
rect 1923 379 1929 380
rect 1923 378 1924 379
rect 1883 376 1924 378
rect 1883 375 1884 376
rect 1878 374 1884 375
rect 1923 375 1924 376
rect 1928 375 1929 379
rect 1923 374 1929 375
rect 2003 379 2009 380
rect 2003 375 2004 379
rect 2008 378 2009 379
rect 2091 379 2097 380
rect 2008 376 2086 378
rect 2008 375 2009 376
rect 2003 374 2009 375
rect 630 370 636 371
rect 315 369 321 370
rect 131 367 137 368
rect 131 363 132 367
rect 136 363 137 367
rect 131 362 137 363
rect 211 367 217 368
rect 211 363 212 367
rect 216 366 217 367
rect 250 367 256 368
rect 250 366 251 367
rect 216 364 251 366
rect 216 363 217 364
rect 211 362 217 363
rect 250 363 251 364
rect 255 363 256 367
rect 315 365 316 369
rect 320 365 321 369
rect 315 364 321 365
rect 358 367 364 368
rect 250 362 256 363
rect 358 363 359 367
rect 363 366 364 367
rect 419 367 425 368
rect 419 366 420 367
rect 363 364 420 366
rect 363 363 364 364
rect 358 362 364 363
rect 419 363 420 364
rect 424 363 425 367
rect 419 362 425 363
rect 462 367 468 368
rect 462 363 463 367
rect 467 366 468 367
rect 523 367 529 368
rect 523 366 524 367
rect 467 364 524 366
rect 467 363 468 364
rect 462 362 468 363
rect 523 363 524 364
rect 528 363 529 367
rect 523 362 529 363
rect 627 367 633 368
rect 627 363 628 367
rect 632 366 633 367
rect 662 367 668 368
rect 662 366 663 367
rect 632 364 663 366
rect 632 363 633 364
rect 627 362 633 363
rect 662 363 663 364
rect 667 363 668 367
rect 662 362 668 363
rect 670 367 676 368
rect 670 363 671 367
rect 675 366 676 367
rect 731 367 737 368
rect 731 366 732 367
rect 675 364 732 366
rect 675 363 676 364
rect 670 362 676 363
rect 731 363 732 364
rect 736 363 737 367
rect 731 362 737 363
rect 827 367 833 368
rect 827 363 828 367
rect 832 366 833 367
rect 870 367 876 368
rect 832 364 866 366
rect 832 363 833 364
rect 827 362 833 363
rect 133 354 135 362
rect 864 354 866 364
rect 870 363 871 367
rect 875 366 876 367
rect 915 367 921 368
rect 915 366 916 367
rect 875 364 916 366
rect 875 363 876 364
rect 870 362 876 363
rect 915 363 916 364
rect 920 363 921 367
rect 915 362 921 363
rect 994 367 1001 368
rect 994 363 995 367
rect 1000 363 1001 367
rect 994 362 1001 363
rect 1074 367 1081 368
rect 1074 363 1075 367
rect 1080 363 1081 367
rect 1074 362 1081 363
rect 1118 367 1124 368
rect 1118 363 1119 367
rect 1123 366 1124 367
rect 1155 367 1161 368
rect 1155 366 1156 367
rect 1123 364 1156 366
rect 1123 363 1124 364
rect 1118 362 1124 363
rect 1155 363 1156 364
rect 1160 363 1161 367
rect 1155 362 1161 363
rect 1198 367 1204 368
rect 1198 363 1199 367
rect 1203 366 1204 367
rect 1219 367 1225 368
rect 1219 366 1220 367
rect 1203 364 1220 366
rect 1203 363 1204 364
rect 1198 362 1204 363
rect 1219 363 1220 364
rect 1224 363 1225 367
rect 1219 362 1225 363
rect 1886 367 1892 368
rect 1886 363 1887 367
rect 1891 366 1892 367
rect 2084 366 2086 376
rect 2091 375 2092 379
rect 2096 378 2097 379
rect 2102 379 2108 380
rect 2102 378 2103 379
rect 2096 376 2103 378
rect 2096 375 2097 376
rect 2091 374 2097 375
rect 2102 375 2103 376
rect 2107 375 2108 379
rect 2102 374 2108 375
rect 2179 379 2185 380
rect 2179 375 2180 379
rect 2184 378 2185 379
rect 2267 379 2273 380
rect 2184 376 2262 378
rect 2184 375 2185 376
rect 2179 374 2185 375
rect 2260 366 2262 376
rect 2267 375 2268 379
rect 2272 378 2273 379
rect 2294 379 2300 380
rect 2294 378 2295 379
rect 2272 376 2295 378
rect 2272 375 2273 376
rect 2267 374 2273 375
rect 2294 375 2295 376
rect 2299 375 2300 379
rect 2294 374 2300 375
rect 2355 379 2361 380
rect 2355 375 2356 379
rect 2360 378 2361 379
rect 2390 379 2396 380
rect 2390 378 2391 379
rect 2360 376 2391 378
rect 2360 375 2361 376
rect 2355 374 2361 375
rect 2390 375 2391 376
rect 2395 375 2396 379
rect 2390 374 2396 375
rect 2435 379 2441 380
rect 2435 375 2436 379
rect 2440 378 2441 379
rect 2474 379 2480 380
rect 2474 378 2475 379
rect 2440 376 2475 378
rect 2440 375 2441 376
rect 2435 374 2441 375
rect 2474 375 2475 376
rect 2479 375 2480 379
rect 2474 374 2480 375
rect 2446 367 2452 368
rect 1891 364 2046 366
rect 2084 364 2134 366
rect 2260 364 2311 366
rect 1891 363 1892 364
rect 1886 362 1892 363
rect 2044 362 2046 364
rect 2132 362 2134 364
rect 2309 362 2311 364
rect 2446 363 2447 367
rect 2451 366 2452 367
rect 2451 364 2479 366
rect 2451 363 2452 364
rect 2446 362 2452 363
rect 2477 362 2479 364
rect 1678 361 1684 362
rect 1326 360 1332 361
rect 1326 356 1327 360
rect 1331 356 1332 360
rect 1678 357 1679 361
rect 1683 357 1684 361
rect 1734 361 1740 362
rect 1678 356 1684 357
rect 1699 359 1708 360
rect 1326 355 1332 356
rect 1699 355 1700 359
rect 1707 355 1708 359
rect 1734 357 1735 361
rect 1739 357 1740 361
rect 1798 361 1804 362
rect 1734 356 1740 357
rect 1755 359 1764 360
rect 1699 354 1708 355
rect 1755 355 1756 359
rect 1763 355 1764 359
rect 1798 357 1799 361
rect 1803 357 1804 361
rect 1870 361 1876 362
rect 1798 356 1804 357
rect 1819 359 1828 360
rect 1755 354 1764 355
rect 1819 355 1820 359
rect 1827 355 1828 359
rect 1870 357 1871 361
rect 1875 357 1876 361
rect 1942 361 1948 362
rect 1870 356 1876 357
rect 1891 359 1900 360
rect 1819 354 1828 355
rect 1891 355 1892 359
rect 1899 355 1900 359
rect 1942 357 1943 361
rect 1947 357 1948 361
rect 2022 361 2028 362
rect 1942 356 1948 357
rect 1962 359 1969 360
rect 1891 354 1900 355
rect 1962 355 1963 359
rect 1968 355 1969 359
rect 2022 357 2023 361
rect 2027 357 2028 361
rect 2022 356 2028 357
rect 2043 361 2049 362
rect 2043 357 2044 361
rect 2048 357 2049 361
rect 2043 356 2049 357
rect 2110 361 2116 362
rect 2110 357 2111 361
rect 2115 357 2116 361
rect 2110 356 2116 357
rect 2131 361 2137 362
rect 2131 357 2132 361
rect 2136 357 2137 361
rect 2131 356 2137 357
rect 2198 361 2204 362
rect 2198 357 2199 361
rect 2203 357 2204 361
rect 2286 361 2292 362
rect 2198 356 2204 357
rect 2206 359 2212 360
rect 1962 354 1969 355
rect 2206 355 2207 359
rect 2211 358 2212 359
rect 2219 359 2225 360
rect 2219 358 2220 359
rect 2211 356 2220 358
rect 2211 355 2212 356
rect 2206 354 2212 355
rect 2219 355 2220 356
rect 2224 355 2225 359
rect 2286 357 2287 361
rect 2291 357 2292 361
rect 2286 356 2292 357
rect 2307 361 2313 362
rect 2307 357 2308 361
rect 2312 357 2313 361
rect 2307 356 2313 357
rect 2374 361 2380 362
rect 2374 357 2375 361
rect 2379 357 2380 361
rect 2454 361 2460 362
rect 2374 356 2380 357
rect 2382 359 2388 360
rect 2219 354 2225 355
rect 2382 355 2383 359
rect 2387 358 2388 359
rect 2395 359 2401 360
rect 2395 358 2396 359
rect 2387 356 2396 358
rect 2387 355 2388 356
rect 2382 354 2388 355
rect 2395 355 2396 356
rect 2400 355 2401 359
rect 2454 357 2455 361
rect 2459 357 2460 361
rect 2454 356 2460 357
rect 2475 361 2481 362
rect 2475 357 2476 361
rect 2480 357 2481 361
rect 2475 356 2481 357
rect 2502 360 2508 361
rect 2502 356 2503 360
rect 2507 356 2508 360
rect 2502 355 2508 356
rect 2395 354 2401 355
rect 133 352 255 354
rect 864 352 1038 354
rect 253 350 255 352
rect 1036 350 1038 352
rect 150 349 156 350
rect 110 348 116 349
rect 110 344 111 348
rect 115 344 116 348
rect 150 345 151 349
rect 155 345 156 349
rect 230 349 236 350
rect 150 344 156 345
rect 170 347 177 348
rect 110 343 116 344
rect 170 343 171 347
rect 176 343 177 347
rect 230 345 231 349
rect 235 345 236 349
rect 230 344 236 345
rect 251 349 257 350
rect 251 345 252 349
rect 256 345 257 349
rect 251 344 257 345
rect 334 349 340 350
rect 334 345 335 349
rect 339 345 340 349
rect 438 349 444 350
rect 334 344 340 345
rect 355 347 364 348
rect 170 342 177 343
rect 355 343 356 347
rect 363 343 364 347
rect 438 345 439 349
rect 443 345 444 349
rect 542 349 548 350
rect 438 344 444 345
rect 459 347 468 348
rect 355 342 364 343
rect 459 343 460 347
rect 467 343 468 347
rect 542 345 543 349
rect 547 345 548 349
rect 646 349 652 350
rect 542 344 548 345
rect 558 347 569 348
rect 459 342 468 343
rect 558 343 559 347
rect 563 343 564 347
rect 568 343 569 347
rect 646 345 647 349
rect 651 345 652 349
rect 750 349 756 350
rect 646 344 652 345
rect 667 347 676 348
rect 558 342 569 343
rect 667 343 668 347
rect 675 343 676 347
rect 750 345 751 349
rect 755 345 756 349
rect 846 349 852 350
rect 750 344 756 345
rect 770 347 777 348
rect 667 342 676 343
rect 770 343 771 347
rect 776 343 777 347
rect 846 345 847 349
rect 851 345 852 349
rect 934 349 940 350
rect 846 344 852 345
rect 867 347 876 348
rect 770 342 777 343
rect 867 343 868 347
rect 875 343 876 347
rect 934 345 935 349
rect 939 345 940 349
rect 1014 349 1020 350
rect 934 344 940 345
rect 950 347 961 348
rect 867 342 876 343
rect 950 343 951 347
rect 955 343 956 347
rect 960 343 961 347
rect 1014 345 1015 349
rect 1019 345 1020 349
rect 1014 344 1020 345
rect 1035 349 1041 350
rect 1035 345 1036 349
rect 1040 345 1041 349
rect 1035 344 1041 345
rect 1094 349 1100 350
rect 1094 345 1095 349
rect 1099 345 1100 349
rect 1174 349 1180 350
rect 1094 344 1100 345
rect 1115 347 1124 348
rect 950 342 961 343
rect 1115 343 1116 347
rect 1123 343 1124 347
rect 1174 345 1175 349
rect 1179 345 1180 349
rect 1238 349 1244 350
rect 1174 344 1180 345
rect 1195 347 1204 348
rect 1115 342 1124 343
rect 1195 343 1196 347
rect 1203 343 1204 347
rect 1238 345 1239 349
rect 1243 345 1244 349
rect 1286 348 1292 349
rect 1238 344 1244 345
rect 1246 347 1252 348
rect 1195 342 1204 343
rect 1246 343 1247 347
rect 1251 346 1252 347
rect 1259 347 1265 348
rect 1259 346 1260 347
rect 1251 344 1260 346
rect 1251 343 1252 344
rect 1246 342 1252 343
rect 1259 343 1260 344
rect 1264 343 1265 347
rect 1286 344 1287 348
rect 1291 344 1292 348
rect 1286 343 1292 344
rect 1326 343 1332 344
rect 1259 342 1265 343
rect 1326 339 1327 343
rect 1331 339 1332 343
rect 2502 343 2508 344
rect 1326 338 1332 339
rect 1662 340 1668 341
rect 1662 336 1663 340
rect 1667 336 1668 340
rect 1662 335 1668 336
rect 1718 340 1724 341
rect 1718 336 1719 340
rect 1723 336 1724 340
rect 1718 335 1724 336
rect 1782 340 1788 341
rect 1782 336 1783 340
rect 1787 336 1788 340
rect 1782 335 1788 336
rect 1854 340 1860 341
rect 1854 336 1855 340
rect 1859 336 1860 340
rect 1854 335 1860 336
rect 1926 340 1932 341
rect 1926 336 1927 340
rect 1931 336 1932 340
rect 1926 335 1932 336
rect 2006 340 2012 341
rect 2006 336 2007 340
rect 2011 336 2012 340
rect 2006 335 2012 336
rect 2094 340 2100 341
rect 2094 336 2095 340
rect 2099 336 2100 340
rect 2094 335 2100 336
rect 2182 340 2188 341
rect 2182 336 2183 340
rect 2187 336 2188 340
rect 2182 335 2188 336
rect 2270 340 2276 341
rect 2270 336 2271 340
rect 2275 336 2276 340
rect 2270 335 2276 336
rect 2358 340 2364 341
rect 2358 336 2359 340
rect 2363 336 2364 340
rect 2358 335 2364 336
rect 2438 340 2444 341
rect 2438 336 2439 340
rect 2443 336 2444 340
rect 2502 339 2503 343
rect 2507 339 2508 343
rect 2502 338 2508 339
rect 2438 335 2444 336
rect 110 331 116 332
rect 110 327 111 331
rect 115 327 116 331
rect 1286 331 1292 332
rect 110 326 116 327
rect 134 328 140 329
rect 134 324 135 328
rect 139 324 140 328
rect 134 323 140 324
rect 214 328 220 329
rect 214 324 215 328
rect 219 324 220 328
rect 214 323 220 324
rect 318 328 324 329
rect 318 324 319 328
rect 323 324 324 328
rect 318 323 324 324
rect 422 328 428 329
rect 422 324 423 328
rect 427 324 428 328
rect 422 323 428 324
rect 526 328 532 329
rect 526 324 527 328
rect 531 324 532 328
rect 526 323 532 324
rect 630 328 636 329
rect 630 324 631 328
rect 635 324 636 328
rect 630 323 636 324
rect 734 328 740 329
rect 734 324 735 328
rect 739 324 740 328
rect 734 323 740 324
rect 830 328 836 329
rect 830 324 831 328
rect 835 324 836 328
rect 830 323 836 324
rect 918 328 924 329
rect 918 324 919 328
rect 923 324 924 328
rect 918 323 924 324
rect 998 328 1004 329
rect 998 324 999 328
rect 1003 324 1004 328
rect 998 323 1004 324
rect 1078 328 1084 329
rect 1078 324 1079 328
rect 1083 324 1084 328
rect 1078 323 1084 324
rect 1158 328 1164 329
rect 1158 324 1159 328
rect 1163 324 1164 328
rect 1158 323 1164 324
rect 1222 328 1228 329
rect 1222 324 1223 328
rect 1227 324 1228 328
rect 1286 327 1287 331
rect 1291 327 1292 331
rect 1286 326 1292 327
rect 1222 323 1228 324
rect 1350 320 1356 321
rect 1326 317 1332 318
rect 1326 313 1327 317
rect 1331 313 1332 317
rect 1350 316 1351 320
rect 1355 316 1356 320
rect 1350 315 1356 316
rect 1454 320 1460 321
rect 1454 316 1455 320
rect 1459 316 1460 320
rect 1454 315 1460 316
rect 1582 320 1588 321
rect 1582 316 1583 320
rect 1587 316 1588 320
rect 1582 315 1588 316
rect 1710 320 1716 321
rect 1710 316 1711 320
rect 1715 316 1716 320
rect 1710 315 1716 316
rect 1838 320 1844 321
rect 1838 316 1839 320
rect 1843 316 1844 320
rect 1838 315 1844 316
rect 1950 320 1956 321
rect 1950 316 1951 320
rect 1955 316 1956 320
rect 1950 315 1956 316
rect 2062 320 2068 321
rect 2062 316 2063 320
rect 2067 316 2068 320
rect 2062 315 2068 316
rect 2166 320 2172 321
rect 2166 316 2167 320
rect 2171 316 2172 320
rect 2166 315 2172 316
rect 2262 320 2268 321
rect 2262 316 2263 320
rect 2267 316 2268 320
rect 2262 315 2268 316
rect 2358 320 2364 321
rect 2358 316 2359 320
rect 2363 316 2364 320
rect 2358 315 2364 316
rect 2438 320 2444 321
rect 2438 316 2439 320
rect 2443 316 2444 320
rect 2438 315 2444 316
rect 2502 317 2508 318
rect 134 312 140 313
rect 110 309 116 310
rect 110 305 111 309
rect 115 305 116 309
rect 134 308 135 312
rect 139 308 140 312
rect 134 307 140 308
rect 214 312 220 313
rect 214 308 215 312
rect 219 308 220 312
rect 214 307 220 308
rect 318 312 324 313
rect 318 308 319 312
rect 323 308 324 312
rect 318 307 324 308
rect 422 312 428 313
rect 422 308 423 312
rect 427 308 428 312
rect 422 307 428 308
rect 534 312 540 313
rect 534 308 535 312
rect 539 308 540 312
rect 534 307 540 308
rect 638 312 644 313
rect 638 308 639 312
rect 643 308 644 312
rect 638 307 644 308
rect 742 312 748 313
rect 742 308 743 312
rect 747 308 748 312
rect 742 307 748 308
rect 846 312 852 313
rect 846 308 847 312
rect 851 308 852 312
rect 846 307 852 308
rect 942 312 948 313
rect 942 308 943 312
rect 947 308 948 312
rect 942 307 948 308
rect 1038 312 1044 313
rect 1038 308 1039 312
rect 1043 308 1044 312
rect 1038 307 1044 308
rect 1142 312 1148 313
rect 1142 308 1143 312
rect 1147 308 1148 312
rect 1142 307 1148 308
rect 1222 312 1228 313
rect 1326 312 1332 313
rect 2502 313 2503 317
rect 2507 313 2508 317
rect 2502 312 2508 313
rect 1222 308 1223 312
rect 1227 308 1228 312
rect 1222 307 1228 308
rect 1286 309 1292 310
rect 110 304 116 305
rect 1286 305 1287 309
rect 1291 305 1292 309
rect 1286 304 1292 305
rect 1326 300 1332 301
rect 2502 300 2508 301
rect 1326 296 1327 300
rect 1331 296 1332 300
rect 1326 295 1332 296
rect 1366 299 1372 300
rect 1366 295 1367 299
rect 1371 295 1372 299
rect 1366 294 1372 295
rect 1374 299 1380 300
rect 1374 295 1375 299
rect 1379 298 1380 299
rect 1387 299 1393 300
rect 1387 298 1388 299
rect 1379 296 1388 298
rect 1379 295 1380 296
rect 1374 294 1380 295
rect 1387 295 1388 296
rect 1392 295 1393 299
rect 1387 294 1393 295
rect 1470 299 1476 300
rect 1470 295 1471 299
rect 1475 295 1476 299
rect 1470 294 1476 295
rect 1491 299 1497 300
rect 1491 295 1492 299
rect 1496 298 1497 299
rect 1578 299 1584 300
rect 1578 298 1579 299
rect 1496 296 1579 298
rect 1496 295 1497 296
rect 1491 294 1497 295
rect 1578 295 1579 296
rect 1583 295 1584 299
rect 1578 294 1584 295
rect 1598 299 1604 300
rect 1598 295 1599 299
rect 1603 295 1604 299
rect 1598 294 1604 295
rect 1619 299 1628 300
rect 1619 295 1620 299
rect 1627 295 1628 299
rect 1619 294 1628 295
rect 1726 299 1732 300
rect 1726 295 1727 299
rect 1731 295 1732 299
rect 1747 299 1753 300
rect 1747 298 1748 299
rect 1726 294 1732 295
rect 1736 296 1748 298
rect 110 292 116 293
rect 1286 292 1292 293
rect 110 288 111 292
rect 115 288 116 292
rect 110 287 116 288
rect 150 291 156 292
rect 150 287 151 291
rect 155 287 156 291
rect 150 286 156 287
rect 171 291 177 292
rect 171 287 172 291
rect 176 290 177 291
rect 210 291 216 292
rect 210 290 211 291
rect 176 288 211 290
rect 176 287 177 288
rect 171 286 177 287
rect 210 287 211 288
rect 215 287 216 291
rect 210 286 216 287
rect 230 291 236 292
rect 230 287 231 291
rect 235 287 236 291
rect 230 286 236 287
rect 250 291 257 292
rect 250 287 251 291
rect 256 287 257 291
rect 250 286 257 287
rect 334 291 340 292
rect 334 287 335 291
rect 339 287 340 291
rect 334 286 340 287
rect 355 291 361 292
rect 355 287 356 291
rect 360 290 361 291
rect 402 291 408 292
rect 402 290 403 291
rect 360 288 403 290
rect 360 287 361 288
rect 355 286 361 287
rect 402 287 403 288
rect 407 287 408 291
rect 402 286 408 287
rect 438 291 444 292
rect 438 287 439 291
rect 443 287 444 291
rect 459 291 465 292
rect 459 290 460 291
rect 438 286 444 287
rect 448 288 460 290
rect 448 278 450 288
rect 459 287 460 288
rect 464 287 465 291
rect 459 286 465 287
rect 550 291 556 292
rect 550 287 551 291
rect 555 287 556 291
rect 571 291 577 292
rect 571 290 572 291
rect 550 286 556 287
rect 560 288 572 290
rect 560 278 562 288
rect 571 287 572 288
rect 576 287 577 291
rect 571 286 577 287
rect 654 291 660 292
rect 654 287 655 291
rect 659 287 660 291
rect 654 286 660 287
rect 662 291 668 292
rect 662 287 663 291
rect 667 290 668 291
rect 675 291 681 292
rect 675 290 676 291
rect 667 288 676 290
rect 667 287 668 288
rect 662 286 668 287
rect 675 287 676 288
rect 680 287 681 291
rect 675 286 681 287
rect 758 291 764 292
rect 758 287 759 291
rect 763 287 764 291
rect 779 291 785 292
rect 779 290 780 291
rect 758 286 764 287
rect 768 288 780 290
rect 768 282 770 288
rect 779 287 780 288
rect 784 287 785 291
rect 779 286 785 287
rect 862 291 868 292
rect 862 287 863 291
rect 867 287 868 291
rect 883 291 889 292
rect 883 290 884 291
rect 862 286 868 287
rect 872 288 884 290
rect 319 276 450 278
rect 452 276 562 278
rect 636 280 770 282
rect 319 274 321 276
rect 452 274 454 276
rect 636 274 638 280
rect 872 278 874 288
rect 883 287 884 288
rect 888 287 889 291
rect 883 286 889 287
rect 958 291 964 292
rect 958 287 959 291
rect 963 287 964 291
rect 958 286 964 287
rect 979 291 985 292
rect 979 287 980 291
rect 984 290 985 291
rect 1034 291 1040 292
rect 1034 290 1035 291
rect 984 288 1035 290
rect 984 287 985 288
rect 979 286 985 287
rect 1034 287 1035 288
rect 1039 287 1040 291
rect 1034 286 1040 287
rect 1054 291 1060 292
rect 1054 287 1055 291
rect 1059 287 1060 291
rect 1054 286 1060 287
rect 1075 291 1081 292
rect 1075 287 1076 291
rect 1080 290 1081 291
rect 1138 291 1144 292
rect 1138 290 1139 291
rect 1080 288 1139 290
rect 1080 287 1081 288
rect 1075 286 1081 287
rect 1138 287 1139 288
rect 1143 287 1144 291
rect 1138 286 1144 287
rect 1158 291 1164 292
rect 1158 287 1159 291
rect 1163 287 1164 291
rect 1158 286 1164 287
rect 1179 291 1185 292
rect 1179 287 1180 291
rect 1184 290 1185 291
rect 1202 291 1208 292
rect 1202 290 1203 291
rect 1184 288 1203 290
rect 1184 287 1185 288
rect 1179 286 1185 287
rect 1202 287 1203 288
rect 1207 287 1208 291
rect 1202 286 1208 287
rect 1238 291 1244 292
rect 1238 287 1239 291
rect 1243 287 1244 291
rect 1238 286 1244 287
rect 1259 291 1265 292
rect 1259 287 1260 291
rect 1264 290 1265 291
rect 1264 288 1282 290
rect 1264 287 1265 288
rect 1259 286 1265 287
rect 1280 282 1282 288
rect 1286 288 1287 292
rect 1291 288 1292 292
rect 1286 287 1292 288
rect 1736 286 1738 296
rect 1747 295 1748 296
rect 1752 295 1753 299
rect 1747 294 1753 295
rect 1854 299 1860 300
rect 1854 295 1855 299
rect 1859 295 1860 299
rect 1854 294 1860 295
rect 1875 299 1884 300
rect 1875 295 1876 299
rect 1883 295 1884 299
rect 1875 294 1884 295
rect 1966 299 1972 300
rect 1966 295 1967 299
rect 1971 295 1972 299
rect 1987 299 1993 300
rect 1987 298 1988 299
rect 1966 294 1972 295
rect 1976 296 1988 298
rect 1976 286 1978 296
rect 1987 295 1988 296
rect 1992 295 1993 299
rect 1987 294 1993 295
rect 2078 299 2084 300
rect 2078 295 2079 299
rect 2083 295 2084 299
rect 2078 294 2084 295
rect 2086 299 2092 300
rect 2086 295 2087 299
rect 2091 298 2092 299
rect 2099 299 2105 300
rect 2099 298 2100 299
rect 2091 296 2100 298
rect 2091 295 2092 296
rect 2086 294 2092 295
rect 2099 295 2100 296
rect 2104 295 2105 299
rect 2099 294 2105 295
rect 2182 299 2188 300
rect 2182 295 2183 299
rect 2187 295 2188 299
rect 2203 299 2209 300
rect 2203 298 2204 299
rect 2182 294 2188 295
rect 2192 296 2204 298
rect 2192 286 2194 296
rect 2203 295 2204 296
rect 2208 295 2209 299
rect 2203 294 2209 295
rect 2278 299 2284 300
rect 2278 295 2279 299
rect 2283 295 2284 299
rect 2278 294 2284 295
rect 2299 299 2305 300
rect 2299 295 2300 299
rect 2304 298 2305 299
rect 2354 299 2360 300
rect 2354 298 2355 299
rect 2304 296 2355 298
rect 2304 295 2305 296
rect 2299 294 2305 295
rect 2354 295 2355 296
rect 2359 295 2360 299
rect 2354 294 2360 295
rect 2374 299 2380 300
rect 2374 295 2375 299
rect 2379 295 2380 299
rect 2395 299 2401 300
rect 2395 298 2396 299
rect 2374 294 2380 295
rect 2384 296 2396 298
rect 2384 286 2386 296
rect 2395 295 2396 296
rect 2400 295 2401 299
rect 2395 294 2401 295
rect 2454 299 2460 300
rect 2454 295 2455 299
rect 2459 295 2460 299
rect 2454 294 2460 295
rect 2474 299 2481 300
rect 2474 295 2475 299
rect 2480 295 2481 299
rect 2502 296 2503 300
rect 2507 296 2508 300
rect 2502 295 2508 296
rect 2474 294 2481 295
rect 1452 284 1738 286
rect 1836 284 1978 286
rect 2060 284 2194 286
rect 2260 284 2386 286
rect 1452 282 1454 284
rect 1836 282 1838 284
rect 2060 282 2062 284
rect 2260 282 2262 284
rect 1280 281 1353 282
rect 1280 280 1348 281
rect 740 276 874 278
rect 1347 277 1348 280
rect 1352 277 1353 281
rect 1347 276 1353 277
rect 1451 281 1457 282
rect 1451 277 1452 281
rect 1456 277 1457 281
rect 1835 281 1841 282
rect 1451 276 1457 277
rect 1578 279 1585 280
rect 740 274 742 276
rect 1578 275 1579 279
rect 1584 275 1585 279
rect 1578 274 1585 275
rect 1707 279 1713 280
rect 1707 275 1708 279
rect 1712 278 1713 279
rect 1778 279 1784 280
rect 1778 278 1779 279
rect 1712 276 1779 278
rect 1712 275 1713 276
rect 1707 274 1713 275
rect 1778 275 1779 276
rect 1783 275 1784 279
rect 1835 277 1836 281
rect 1840 277 1841 281
rect 2059 281 2065 282
rect 1835 276 1841 277
rect 1947 279 1953 280
rect 1778 274 1784 275
rect 1947 275 1948 279
rect 1952 278 1953 279
rect 1986 279 1992 280
rect 1986 278 1987 279
rect 1952 276 1987 278
rect 1952 275 1953 276
rect 1947 274 1953 275
rect 1986 275 1987 276
rect 1991 275 1992 279
rect 2059 277 2060 281
rect 2064 277 2065 281
rect 2259 281 2265 282
rect 2059 276 2065 277
rect 2163 279 2169 280
rect 1986 274 1992 275
rect 2163 275 2164 279
rect 2168 278 2169 279
rect 2206 279 2212 280
rect 2206 278 2207 279
rect 2168 276 2207 278
rect 2168 275 2169 276
rect 2163 274 2169 275
rect 2206 275 2207 276
rect 2211 275 2212 279
rect 2259 277 2260 281
rect 2264 277 2265 281
rect 2259 276 2265 277
rect 2355 279 2361 280
rect 2206 274 2212 275
rect 2355 275 2356 279
rect 2360 278 2361 279
rect 2382 279 2388 280
rect 2382 278 2383 279
rect 2360 276 2383 278
rect 2360 275 2361 276
rect 2355 274 2361 275
rect 2382 275 2383 276
rect 2387 275 2388 279
rect 2382 274 2388 275
rect 2435 279 2441 280
rect 2435 275 2436 279
rect 2440 278 2441 279
rect 2462 279 2468 280
rect 2462 278 2463 279
rect 2440 276 2463 278
rect 2440 275 2441 276
rect 2435 274 2441 275
rect 2462 275 2463 276
rect 2467 275 2468 279
rect 2462 274 2468 275
rect 315 273 321 274
rect 131 271 137 272
rect 131 267 132 271
rect 136 270 137 271
rect 170 271 176 272
rect 170 270 171 271
rect 136 268 171 270
rect 136 267 137 268
rect 131 266 137 267
rect 170 267 171 268
rect 175 267 176 271
rect 170 266 176 267
rect 210 271 217 272
rect 210 267 211 271
rect 216 267 217 271
rect 315 269 316 273
rect 320 269 321 273
rect 315 268 321 269
rect 419 273 454 274
rect 419 269 420 273
rect 424 272 454 273
rect 635 273 641 274
rect 424 269 425 272
rect 419 268 425 269
rect 531 271 537 272
rect 210 266 217 267
rect 531 267 532 271
rect 536 270 537 271
rect 558 271 564 272
rect 558 270 559 271
rect 536 268 559 270
rect 536 267 537 268
rect 531 266 537 267
rect 558 267 559 268
rect 563 267 564 271
rect 635 269 636 273
rect 640 269 641 273
rect 635 268 641 269
rect 739 273 745 274
rect 739 269 740 273
rect 744 269 745 273
rect 739 268 745 269
rect 843 271 849 272
rect 558 266 564 267
rect 843 267 844 271
rect 848 270 849 271
rect 890 271 896 272
rect 890 270 891 271
rect 848 268 891 270
rect 848 267 849 268
rect 843 266 849 267
rect 890 267 891 268
rect 895 267 896 271
rect 890 266 896 267
rect 939 271 945 272
rect 939 267 940 271
rect 944 270 945 271
rect 950 271 956 272
rect 950 270 951 271
rect 944 268 951 270
rect 944 267 945 268
rect 939 266 945 267
rect 950 267 951 268
rect 955 267 956 271
rect 950 266 956 267
rect 1034 271 1041 272
rect 1034 267 1035 271
rect 1040 267 1041 271
rect 1034 266 1041 267
rect 1138 271 1145 272
rect 1138 267 1139 271
rect 1144 267 1145 271
rect 1138 266 1145 267
rect 1219 271 1225 272
rect 1219 267 1220 271
rect 1224 270 1225 271
rect 1246 271 1252 272
rect 1246 270 1247 271
rect 1224 268 1247 270
rect 1224 267 1225 268
rect 1219 266 1225 267
rect 1246 267 1247 268
rect 1251 267 1252 271
rect 1246 266 1252 267
rect 131 259 137 260
rect 131 255 132 259
rect 136 258 137 259
rect 203 259 209 260
rect 136 256 198 258
rect 136 255 137 256
rect 131 254 137 255
rect 196 246 198 256
rect 203 255 204 259
rect 208 258 209 259
rect 299 259 305 260
rect 208 256 266 258
rect 208 255 209 256
rect 203 254 209 255
rect 264 246 266 256
rect 299 255 300 259
rect 304 258 305 259
rect 310 259 316 260
rect 310 258 311 259
rect 304 256 311 258
rect 304 255 305 256
rect 299 254 305 255
rect 310 255 311 256
rect 315 255 316 259
rect 310 254 316 255
rect 402 259 409 260
rect 402 255 403 259
rect 408 255 409 259
rect 402 254 409 255
rect 446 259 452 260
rect 446 255 447 259
rect 451 258 452 259
rect 515 259 521 260
rect 515 258 516 259
rect 451 256 516 258
rect 451 255 452 256
rect 446 254 452 255
rect 515 255 516 256
rect 520 255 521 259
rect 515 254 521 255
rect 558 259 564 260
rect 558 255 559 259
rect 563 258 564 259
rect 627 259 633 260
rect 627 258 628 259
rect 563 256 628 258
rect 563 255 564 256
rect 558 254 564 255
rect 627 255 628 256
rect 632 255 633 259
rect 627 254 633 255
rect 734 259 745 260
rect 734 255 735 259
rect 739 255 740 259
rect 744 255 745 259
rect 734 254 745 255
rect 782 259 788 260
rect 782 255 783 259
rect 787 258 788 259
rect 851 259 857 260
rect 851 258 852 259
rect 787 256 852 258
rect 787 255 788 256
rect 782 254 788 255
rect 851 255 852 256
rect 856 255 857 259
rect 851 254 857 255
rect 963 259 969 260
rect 963 255 964 259
rect 968 258 969 259
rect 1083 259 1089 260
rect 968 256 1078 258
rect 968 255 969 256
rect 963 254 969 255
rect 1076 246 1078 256
rect 1083 255 1084 259
rect 1088 258 1089 259
rect 1202 259 1209 260
rect 1088 256 1161 258
rect 1088 255 1089 256
rect 1083 254 1089 255
rect 1159 246 1161 256
rect 1202 255 1203 259
rect 1208 255 1209 259
rect 1202 254 1209 255
rect 1347 259 1353 260
rect 1347 255 1348 259
rect 1352 258 1353 259
rect 1374 259 1380 260
rect 1374 258 1375 259
rect 1352 256 1375 258
rect 1352 255 1353 256
rect 1347 254 1353 255
rect 1374 255 1375 256
rect 1379 255 1380 259
rect 1374 254 1380 255
rect 1390 259 1396 260
rect 1390 255 1391 259
rect 1395 258 1396 259
rect 1427 259 1433 260
rect 1427 258 1428 259
rect 1395 256 1428 258
rect 1395 255 1396 256
rect 1390 254 1396 255
rect 1427 255 1428 256
rect 1432 255 1433 259
rect 1427 254 1433 255
rect 1531 259 1537 260
rect 1531 255 1532 259
rect 1536 258 1537 259
rect 1574 259 1580 260
rect 1536 256 1570 258
rect 1536 255 1537 256
rect 1531 254 1537 255
rect 1568 250 1570 256
rect 1574 255 1575 259
rect 1579 258 1580 259
rect 1635 259 1641 260
rect 1635 258 1636 259
rect 1579 256 1636 258
rect 1579 255 1580 256
rect 1574 254 1580 255
rect 1635 255 1636 256
rect 1640 255 1641 259
rect 1635 254 1641 255
rect 1678 259 1684 260
rect 1678 255 1679 259
rect 1683 258 1684 259
rect 1739 259 1745 260
rect 1739 258 1740 259
rect 1683 256 1740 258
rect 1683 255 1684 256
rect 1678 254 1684 255
rect 1739 255 1740 256
rect 1744 255 1745 259
rect 1739 254 1745 255
rect 1838 259 1849 260
rect 1838 255 1839 259
rect 1843 255 1844 259
rect 1848 255 1849 259
rect 1838 254 1849 255
rect 1886 259 1892 260
rect 1886 255 1887 259
rect 1891 258 1892 259
rect 1947 259 1953 260
rect 1947 258 1948 259
rect 1891 256 1948 258
rect 1891 255 1892 256
rect 1886 254 1892 255
rect 1947 255 1948 256
rect 1952 255 1953 259
rect 1947 254 1953 255
rect 2051 259 2057 260
rect 2051 255 2052 259
rect 2056 258 2057 259
rect 2086 259 2092 260
rect 2086 258 2087 259
rect 2056 256 2087 258
rect 2056 255 2057 256
rect 2051 254 2057 255
rect 2086 255 2087 256
rect 2091 255 2092 259
rect 2086 254 2092 255
rect 2094 259 2100 260
rect 2094 255 2095 259
rect 2099 258 2100 259
rect 2155 259 2161 260
rect 2155 258 2156 259
rect 2099 256 2156 258
rect 2099 255 2100 256
rect 2094 254 2100 255
rect 2155 255 2156 256
rect 2160 255 2161 259
rect 2155 254 2161 255
rect 2198 259 2204 260
rect 2198 255 2199 259
rect 2203 258 2204 259
rect 2251 259 2257 260
rect 2251 258 2252 259
rect 2203 256 2252 258
rect 2203 255 2204 256
rect 2198 254 2204 255
rect 2251 255 2252 256
rect 2256 255 2257 259
rect 2251 254 2257 255
rect 2354 259 2361 260
rect 2354 255 2355 259
rect 2360 255 2361 259
rect 2354 254 2361 255
rect 2398 259 2404 260
rect 2398 255 2399 259
rect 2403 258 2404 259
rect 2435 259 2441 260
rect 2435 258 2436 259
rect 2403 256 2436 258
rect 2403 255 2404 256
rect 2398 254 2404 255
rect 2435 255 2436 256
rect 2440 255 2441 259
rect 2435 254 2441 255
rect 1586 251 1592 252
rect 1586 250 1587 251
rect 1568 248 1587 250
rect 1586 247 1587 248
rect 1591 247 1592 251
rect 1586 246 1592 247
rect 196 244 246 246
rect 264 244 342 246
rect 1076 244 1126 246
rect 1159 244 1246 246
rect 244 242 246 244
rect 340 242 342 244
rect 1124 242 1126 244
rect 1244 242 1246 244
rect 150 241 156 242
rect 110 240 116 241
rect 110 236 111 240
rect 115 236 116 240
rect 150 237 151 241
rect 155 237 156 241
rect 222 241 228 242
rect 150 236 156 237
rect 170 239 177 240
rect 110 235 116 236
rect 170 235 171 239
rect 176 235 177 239
rect 222 237 223 241
rect 227 237 228 241
rect 222 236 228 237
rect 243 241 249 242
rect 243 237 244 241
rect 248 237 249 241
rect 243 236 249 237
rect 318 241 324 242
rect 318 237 319 241
rect 323 237 324 241
rect 318 236 324 237
rect 339 241 345 242
rect 339 237 340 241
rect 344 237 345 241
rect 339 236 345 237
rect 422 241 428 242
rect 422 237 423 241
rect 427 237 428 241
rect 534 241 540 242
rect 422 236 428 237
rect 443 239 452 240
rect 170 234 177 235
rect 443 235 444 239
rect 451 235 452 239
rect 534 237 535 241
rect 539 237 540 241
rect 646 241 652 242
rect 534 236 540 237
rect 555 239 564 240
rect 443 234 452 235
rect 555 235 556 239
rect 563 235 564 239
rect 646 237 647 241
rect 651 237 652 241
rect 758 241 764 242
rect 646 236 652 237
rect 654 239 660 240
rect 555 234 564 235
rect 654 235 655 239
rect 659 238 660 239
rect 667 239 673 240
rect 667 238 668 239
rect 659 236 668 238
rect 659 235 660 236
rect 654 234 660 235
rect 667 235 668 236
rect 672 235 673 239
rect 758 237 759 241
rect 763 237 764 241
rect 870 241 876 242
rect 758 236 764 237
rect 779 239 788 240
rect 667 234 673 235
rect 779 235 780 239
rect 787 235 788 239
rect 870 237 871 241
rect 875 237 876 241
rect 982 241 988 242
rect 870 236 876 237
rect 890 239 897 240
rect 779 234 788 235
rect 890 235 891 239
rect 896 235 897 239
rect 982 237 983 241
rect 987 237 988 241
rect 1102 241 1108 242
rect 982 236 988 237
rect 990 239 996 240
rect 890 234 897 235
rect 990 235 991 239
rect 995 238 996 239
rect 1003 239 1009 240
rect 1003 238 1004 239
rect 995 236 1004 238
rect 995 235 996 236
rect 990 234 996 235
rect 1003 235 1004 236
rect 1008 235 1009 239
rect 1102 237 1103 241
rect 1107 237 1108 241
rect 1102 236 1108 237
rect 1123 241 1129 242
rect 1123 237 1124 241
rect 1128 237 1129 241
rect 1123 236 1129 237
rect 1222 241 1228 242
rect 1222 237 1223 241
rect 1227 237 1228 241
rect 1222 236 1228 237
rect 1243 241 1249 242
rect 1366 241 1372 242
rect 1243 237 1244 241
rect 1248 237 1249 241
rect 1243 236 1249 237
rect 1286 240 1292 241
rect 1286 236 1287 240
rect 1291 236 1292 240
rect 1286 235 1292 236
rect 1326 240 1332 241
rect 1326 236 1327 240
rect 1331 236 1332 240
rect 1366 237 1367 241
rect 1371 237 1372 241
rect 1446 241 1452 242
rect 1366 236 1372 237
rect 1387 239 1396 240
rect 1326 235 1332 236
rect 1387 235 1388 239
rect 1395 235 1396 239
rect 1446 237 1447 241
rect 1451 237 1452 241
rect 1550 241 1556 242
rect 1446 236 1452 237
rect 1462 239 1473 240
rect 1003 234 1009 235
rect 1387 234 1396 235
rect 1462 235 1463 239
rect 1467 235 1468 239
rect 1472 235 1473 239
rect 1550 237 1551 241
rect 1555 237 1556 241
rect 1654 241 1660 242
rect 1550 236 1556 237
rect 1571 239 1580 240
rect 1462 234 1473 235
rect 1571 235 1572 239
rect 1579 235 1580 239
rect 1654 237 1655 241
rect 1659 237 1660 241
rect 1758 241 1764 242
rect 1654 236 1660 237
rect 1675 239 1684 240
rect 1571 234 1580 235
rect 1675 235 1676 239
rect 1683 235 1684 239
rect 1758 237 1759 241
rect 1763 237 1764 241
rect 1862 241 1868 242
rect 1758 236 1764 237
rect 1778 239 1785 240
rect 1675 234 1684 235
rect 1778 235 1779 239
rect 1784 235 1785 239
rect 1862 237 1863 241
rect 1867 237 1868 241
rect 1966 241 1972 242
rect 1862 236 1868 237
rect 1883 239 1892 240
rect 1778 234 1785 235
rect 1883 235 1884 239
rect 1891 235 1892 239
rect 1966 237 1967 241
rect 1971 237 1972 241
rect 2070 241 2076 242
rect 1966 236 1972 237
rect 1986 239 1993 240
rect 1883 234 1892 235
rect 1986 235 1987 239
rect 1992 235 1993 239
rect 2070 237 2071 241
rect 2075 237 2076 241
rect 2174 241 2180 242
rect 2070 236 2076 237
rect 2091 239 2100 240
rect 1986 234 1993 235
rect 2091 235 2092 239
rect 2099 235 2100 239
rect 2174 237 2175 241
rect 2179 237 2180 241
rect 2270 241 2276 242
rect 2174 236 2180 237
rect 2195 239 2204 240
rect 2091 234 2100 235
rect 2195 235 2196 239
rect 2203 235 2204 239
rect 2270 237 2271 241
rect 2275 237 2276 241
rect 2374 241 2380 242
rect 2270 236 2276 237
rect 2291 239 2297 240
rect 2195 234 2204 235
rect 2291 235 2292 239
rect 2296 238 2297 239
rect 2326 239 2332 240
rect 2326 238 2327 239
rect 2296 236 2327 238
rect 2296 235 2297 236
rect 2291 234 2297 235
rect 2326 235 2327 236
rect 2331 235 2332 239
rect 2374 237 2375 241
rect 2379 237 2380 241
rect 2454 241 2460 242
rect 2374 236 2380 237
rect 2395 239 2404 240
rect 2326 234 2332 235
rect 2395 235 2396 239
rect 2403 235 2404 239
rect 2454 237 2455 241
rect 2459 237 2460 241
rect 2502 240 2508 241
rect 2454 236 2460 237
rect 2470 239 2481 240
rect 2395 234 2404 235
rect 2470 235 2471 239
rect 2475 235 2476 239
rect 2480 235 2481 239
rect 2502 236 2503 240
rect 2507 236 2508 240
rect 2502 235 2508 236
rect 2470 234 2481 235
rect 110 223 116 224
rect 110 219 111 223
rect 115 219 116 223
rect 1286 223 1292 224
rect 110 218 116 219
rect 134 220 140 221
rect 134 216 135 220
rect 139 216 140 220
rect 134 215 140 216
rect 206 220 212 221
rect 206 216 207 220
rect 211 216 212 220
rect 206 215 212 216
rect 302 220 308 221
rect 302 216 303 220
rect 307 216 308 220
rect 302 215 308 216
rect 406 220 412 221
rect 406 216 407 220
rect 411 216 412 220
rect 406 215 412 216
rect 518 220 524 221
rect 518 216 519 220
rect 523 216 524 220
rect 518 215 524 216
rect 630 220 636 221
rect 630 216 631 220
rect 635 216 636 220
rect 630 215 636 216
rect 742 220 748 221
rect 742 216 743 220
rect 747 216 748 220
rect 742 215 748 216
rect 854 220 860 221
rect 854 216 855 220
rect 859 216 860 220
rect 854 215 860 216
rect 966 220 972 221
rect 966 216 967 220
rect 971 216 972 220
rect 966 215 972 216
rect 1086 220 1092 221
rect 1086 216 1087 220
rect 1091 216 1092 220
rect 1086 215 1092 216
rect 1206 220 1212 221
rect 1206 216 1207 220
rect 1211 216 1212 220
rect 1286 219 1287 223
rect 1291 219 1292 223
rect 1286 218 1292 219
rect 1326 223 1332 224
rect 1326 219 1327 223
rect 1331 219 1332 223
rect 2502 223 2508 224
rect 1326 218 1332 219
rect 1350 220 1356 221
rect 1206 215 1212 216
rect 1350 216 1351 220
rect 1355 216 1356 220
rect 1350 215 1356 216
rect 1430 220 1436 221
rect 1430 216 1431 220
rect 1435 216 1436 220
rect 1430 215 1436 216
rect 1534 220 1540 221
rect 1534 216 1535 220
rect 1539 216 1540 220
rect 1534 215 1540 216
rect 1638 220 1644 221
rect 1638 216 1639 220
rect 1643 216 1644 220
rect 1638 215 1644 216
rect 1742 220 1748 221
rect 1742 216 1743 220
rect 1747 216 1748 220
rect 1742 215 1748 216
rect 1846 220 1852 221
rect 1846 216 1847 220
rect 1851 216 1852 220
rect 1846 215 1852 216
rect 1950 220 1956 221
rect 1950 216 1951 220
rect 1955 216 1956 220
rect 1950 215 1956 216
rect 2054 220 2060 221
rect 2054 216 2055 220
rect 2059 216 2060 220
rect 2054 215 2060 216
rect 2158 220 2164 221
rect 2158 216 2159 220
rect 2163 216 2164 220
rect 2158 215 2164 216
rect 2254 220 2260 221
rect 2254 216 2255 220
rect 2259 216 2260 220
rect 2254 215 2260 216
rect 2358 220 2364 221
rect 2358 216 2359 220
rect 2363 216 2364 220
rect 2358 215 2364 216
rect 2438 220 2444 221
rect 2438 216 2439 220
rect 2443 216 2444 220
rect 2502 219 2503 223
rect 2507 219 2508 223
rect 2502 218 2508 219
rect 2438 215 2444 216
rect 182 204 188 205
rect 110 201 116 202
rect 110 197 111 201
rect 115 197 116 201
rect 182 200 183 204
rect 187 200 188 204
rect 182 199 188 200
rect 278 204 284 205
rect 278 200 279 204
rect 283 200 284 204
rect 278 199 284 200
rect 382 204 388 205
rect 382 200 383 204
rect 387 200 388 204
rect 382 199 388 200
rect 486 204 492 205
rect 486 200 487 204
rect 491 200 492 204
rect 486 199 492 200
rect 590 204 596 205
rect 590 200 591 204
rect 595 200 596 204
rect 590 199 596 200
rect 694 204 700 205
rect 694 200 695 204
rect 699 200 700 204
rect 694 199 700 200
rect 798 204 804 205
rect 798 200 799 204
rect 803 200 804 204
rect 798 199 804 200
rect 894 204 900 205
rect 894 200 895 204
rect 899 200 900 204
rect 894 199 900 200
rect 998 204 1004 205
rect 998 200 999 204
rect 1003 200 1004 204
rect 998 199 1004 200
rect 1102 204 1108 205
rect 1102 200 1103 204
rect 1107 200 1108 204
rect 1350 204 1356 205
rect 1102 199 1108 200
rect 1286 201 1292 202
rect 110 196 116 197
rect 1286 197 1287 201
rect 1291 197 1292 201
rect 1286 196 1292 197
rect 1326 201 1332 202
rect 1326 197 1327 201
rect 1331 197 1332 201
rect 1350 200 1351 204
rect 1355 200 1356 204
rect 1350 199 1356 200
rect 1406 204 1412 205
rect 1406 200 1407 204
rect 1411 200 1412 204
rect 1406 199 1412 200
rect 1470 204 1476 205
rect 1470 200 1471 204
rect 1475 200 1476 204
rect 1470 199 1476 200
rect 1550 204 1556 205
rect 1550 200 1551 204
rect 1555 200 1556 204
rect 1550 199 1556 200
rect 1638 204 1644 205
rect 1638 200 1639 204
rect 1643 200 1644 204
rect 1638 199 1644 200
rect 1718 204 1724 205
rect 1718 200 1719 204
rect 1723 200 1724 204
rect 1718 199 1724 200
rect 1806 204 1812 205
rect 1806 200 1807 204
rect 1811 200 1812 204
rect 1806 199 1812 200
rect 1894 204 1900 205
rect 1894 200 1895 204
rect 1899 200 1900 204
rect 1894 199 1900 200
rect 1990 204 1996 205
rect 1990 200 1991 204
rect 1995 200 1996 204
rect 1990 199 1996 200
rect 2102 204 2108 205
rect 2102 200 2103 204
rect 2107 200 2108 204
rect 2102 199 2108 200
rect 2214 204 2220 205
rect 2214 200 2215 204
rect 2219 200 2220 204
rect 2214 199 2220 200
rect 2334 204 2340 205
rect 2334 200 2335 204
rect 2339 200 2340 204
rect 2334 199 2340 200
rect 2438 204 2444 205
rect 2438 200 2439 204
rect 2443 200 2444 204
rect 2438 199 2444 200
rect 2502 201 2508 202
rect 1326 196 1332 197
rect 2502 197 2503 201
rect 2507 197 2508 201
rect 2502 196 2508 197
rect 110 184 116 185
rect 1286 184 1292 185
rect 110 180 111 184
rect 115 180 116 184
rect 110 179 116 180
rect 198 183 204 184
rect 198 179 199 183
rect 203 179 204 183
rect 198 178 204 179
rect 219 183 225 184
rect 219 179 220 183
rect 224 182 225 183
rect 274 183 280 184
rect 274 182 275 183
rect 224 180 275 182
rect 224 179 225 180
rect 219 178 225 179
rect 274 179 275 180
rect 279 179 280 183
rect 274 178 280 179
rect 294 183 300 184
rect 294 179 295 183
rect 299 179 300 183
rect 294 178 300 179
rect 310 183 321 184
rect 310 179 311 183
rect 315 179 316 183
rect 320 179 321 183
rect 310 178 321 179
rect 398 183 404 184
rect 398 179 399 183
rect 403 179 404 183
rect 398 178 404 179
rect 419 183 425 184
rect 419 179 420 183
rect 424 182 425 183
rect 466 183 472 184
rect 466 182 467 183
rect 424 180 467 182
rect 424 179 425 180
rect 419 178 425 179
rect 466 179 467 180
rect 471 179 472 183
rect 466 178 472 179
rect 502 183 508 184
rect 502 179 503 183
rect 507 179 508 183
rect 523 183 529 184
rect 523 182 524 183
rect 502 178 508 179
rect 512 180 524 182
rect 512 174 514 180
rect 523 179 524 180
rect 528 179 529 183
rect 523 178 529 179
rect 606 183 612 184
rect 606 179 607 183
rect 611 179 612 183
rect 627 183 633 184
rect 627 182 628 183
rect 606 178 612 179
rect 616 180 628 182
rect 380 172 514 174
rect 380 166 382 172
rect 616 170 618 180
rect 627 179 628 180
rect 632 179 633 183
rect 627 178 633 179
rect 710 183 716 184
rect 710 179 711 183
rect 715 179 716 183
rect 710 178 716 179
rect 731 183 740 184
rect 731 179 732 183
rect 739 179 740 183
rect 731 178 740 179
rect 814 183 820 184
rect 814 179 815 183
rect 819 179 820 183
rect 835 183 841 184
rect 835 182 836 183
rect 814 178 820 179
rect 824 180 836 182
rect 824 170 826 180
rect 835 179 836 180
rect 840 179 841 183
rect 835 178 841 179
rect 910 183 916 184
rect 910 179 911 183
rect 915 179 916 183
rect 910 178 916 179
rect 931 183 937 184
rect 931 179 932 183
rect 936 182 937 183
rect 994 183 1000 184
rect 994 182 995 183
rect 936 180 995 182
rect 936 179 937 180
rect 931 178 937 179
rect 994 179 995 180
rect 999 179 1000 183
rect 994 178 1000 179
rect 1014 183 1020 184
rect 1014 179 1015 183
rect 1019 179 1020 183
rect 1014 178 1020 179
rect 1035 183 1041 184
rect 1035 179 1036 183
rect 1040 182 1041 183
rect 1098 183 1104 184
rect 1098 182 1099 183
rect 1040 180 1099 182
rect 1040 179 1041 180
rect 1035 178 1041 179
rect 1098 179 1099 180
rect 1103 179 1104 183
rect 1098 178 1104 179
rect 1118 183 1124 184
rect 1118 179 1119 183
rect 1123 179 1124 183
rect 1118 178 1124 179
rect 1134 183 1145 184
rect 1134 179 1135 183
rect 1139 179 1140 183
rect 1144 179 1145 183
rect 1286 180 1287 184
rect 1291 180 1292 184
rect 1286 179 1292 180
rect 1326 184 1332 185
rect 2502 184 2508 185
rect 1326 180 1327 184
rect 1331 180 1332 184
rect 1326 179 1332 180
rect 1366 183 1372 184
rect 1366 179 1367 183
rect 1371 179 1372 183
rect 1134 178 1145 179
rect 1366 178 1372 179
rect 1374 183 1380 184
rect 1374 179 1375 183
rect 1379 182 1380 183
rect 1387 183 1393 184
rect 1387 182 1388 183
rect 1379 180 1388 182
rect 1379 179 1380 180
rect 1374 178 1380 179
rect 1387 179 1388 180
rect 1392 179 1393 183
rect 1387 178 1393 179
rect 1422 183 1428 184
rect 1422 179 1423 183
rect 1427 179 1428 183
rect 1443 183 1449 184
rect 1443 182 1444 183
rect 1422 178 1428 179
rect 1432 180 1444 182
rect 1432 170 1434 180
rect 1443 179 1444 180
rect 1448 179 1449 183
rect 1443 178 1449 179
rect 1486 183 1492 184
rect 1486 179 1487 183
rect 1491 179 1492 183
rect 1507 183 1513 184
rect 1507 182 1508 183
rect 1486 178 1492 179
rect 1496 180 1508 182
rect 1496 174 1498 180
rect 1507 179 1508 180
rect 1512 179 1513 183
rect 1507 178 1513 179
rect 1566 183 1572 184
rect 1566 179 1567 183
rect 1571 179 1572 183
rect 1566 178 1572 179
rect 1586 183 1593 184
rect 1586 179 1587 183
rect 1592 179 1593 183
rect 1586 178 1593 179
rect 1654 183 1660 184
rect 1654 179 1655 183
rect 1659 179 1660 183
rect 1675 183 1681 184
rect 1675 182 1676 183
rect 1654 178 1660 179
rect 1664 180 1676 182
rect 1664 174 1666 180
rect 1675 179 1676 180
rect 1680 179 1681 183
rect 1675 178 1681 179
rect 1734 183 1740 184
rect 1734 179 1735 183
rect 1739 179 1740 183
rect 1755 183 1761 184
rect 1755 182 1756 183
rect 1734 178 1740 179
rect 1744 180 1756 182
rect 484 168 618 170
rect 692 168 826 170
rect 1348 168 1434 170
rect 1436 172 1498 174
rect 1548 172 1666 174
rect 484 166 486 168
rect 692 166 694 168
rect 1348 166 1350 168
rect 1436 166 1438 172
rect 1548 166 1550 172
rect 1744 170 1746 180
rect 1755 179 1756 180
rect 1760 179 1761 183
rect 1755 178 1761 179
rect 1822 183 1828 184
rect 1822 179 1823 183
rect 1827 179 1828 183
rect 1822 178 1828 179
rect 1838 183 1849 184
rect 1838 179 1839 183
rect 1843 179 1844 183
rect 1848 179 1849 183
rect 1838 178 1849 179
rect 1910 183 1916 184
rect 1910 179 1911 183
rect 1915 179 1916 183
rect 1931 183 1937 184
rect 1931 182 1932 183
rect 1910 178 1916 179
rect 1920 180 1932 182
rect 1920 174 1922 180
rect 1931 179 1932 180
rect 1936 179 1937 183
rect 1931 178 1937 179
rect 2006 183 2012 184
rect 2006 179 2007 183
rect 2011 179 2012 183
rect 2027 183 2033 184
rect 2027 182 2028 183
rect 2006 178 2012 179
rect 2016 180 2028 182
rect 1636 168 1746 170
rect 1804 172 1922 174
rect 1636 166 1638 168
rect 1804 166 1806 172
rect 2016 170 2018 180
rect 2027 179 2028 180
rect 2032 179 2033 183
rect 2027 178 2033 179
rect 2118 183 2124 184
rect 2118 179 2119 183
rect 2123 179 2124 183
rect 2118 178 2124 179
rect 2126 183 2132 184
rect 2126 179 2127 183
rect 2131 182 2132 183
rect 2139 183 2145 184
rect 2139 182 2140 183
rect 2131 180 2140 182
rect 2131 179 2132 180
rect 2126 178 2132 179
rect 2139 179 2140 180
rect 2144 179 2145 183
rect 2139 178 2145 179
rect 2230 183 2236 184
rect 2230 179 2231 183
rect 2235 179 2236 183
rect 2251 183 2257 184
rect 2251 182 2252 183
rect 2230 178 2236 179
rect 2240 180 2252 182
rect 2240 170 2242 180
rect 2251 179 2252 180
rect 2256 179 2257 183
rect 2251 178 2257 179
rect 2350 183 2356 184
rect 2350 179 2351 183
rect 2355 179 2356 183
rect 2371 183 2377 184
rect 2371 182 2372 183
rect 2350 178 2356 179
rect 2360 180 2372 182
rect 2360 174 2362 180
rect 2371 179 2372 180
rect 2376 179 2377 183
rect 2371 178 2377 179
rect 2454 183 2460 184
rect 2454 179 2455 183
rect 2459 179 2460 183
rect 2454 178 2460 179
rect 2462 183 2468 184
rect 2462 179 2463 183
rect 2467 182 2468 183
rect 2475 183 2481 184
rect 2475 182 2476 183
rect 2467 180 2476 182
rect 2467 179 2468 180
rect 2462 178 2468 179
rect 2475 179 2476 180
rect 2480 179 2481 183
rect 2502 180 2503 184
rect 2507 180 2508 184
rect 2502 179 2508 180
rect 2475 178 2481 179
rect 1892 168 2018 170
rect 2100 168 2242 170
rect 2244 172 2362 174
rect 1892 166 1894 168
rect 2100 166 2102 168
rect 2244 166 2246 172
rect 379 165 385 166
rect 179 163 185 164
rect 179 159 180 163
rect 184 162 185 163
rect 226 163 232 164
rect 226 162 227 163
rect 184 160 227 162
rect 184 159 185 160
rect 179 158 185 159
rect 226 159 227 160
rect 231 159 232 163
rect 226 158 232 159
rect 274 163 281 164
rect 274 159 275 163
rect 280 159 281 163
rect 379 161 380 165
rect 384 161 385 165
rect 379 160 385 161
rect 483 165 489 166
rect 483 161 484 165
rect 488 161 489 165
rect 691 165 697 166
rect 483 160 489 161
rect 587 163 593 164
rect 274 158 281 159
rect 587 159 588 163
rect 592 162 593 163
rect 654 163 660 164
rect 654 162 655 163
rect 592 160 655 162
rect 592 159 593 160
rect 587 158 593 159
rect 654 159 655 160
rect 659 159 660 163
rect 691 161 692 165
rect 696 161 697 165
rect 1347 165 1353 166
rect 691 160 697 161
rect 790 163 801 164
rect 654 158 660 159
rect 790 159 791 163
rect 795 159 796 163
rect 800 159 801 163
rect 790 158 801 159
rect 891 163 897 164
rect 891 159 892 163
rect 896 162 897 163
rect 986 163 992 164
rect 986 162 987 163
rect 896 160 987 162
rect 896 159 897 160
rect 891 158 897 159
rect 986 159 987 160
rect 991 159 992 163
rect 986 158 992 159
rect 994 163 1001 164
rect 994 159 995 163
rect 1000 159 1001 163
rect 994 158 1001 159
rect 1098 163 1105 164
rect 1098 159 1099 163
rect 1104 159 1105 163
rect 1347 161 1348 165
rect 1352 161 1353 165
rect 1347 160 1353 161
rect 1403 165 1438 166
rect 1403 161 1404 165
rect 1408 164 1438 165
rect 1547 165 1553 166
rect 1408 161 1409 164
rect 1403 160 1409 161
rect 1462 163 1473 164
rect 1098 158 1105 159
rect 1462 159 1463 163
rect 1467 159 1468 163
rect 1472 159 1473 163
rect 1547 161 1548 165
rect 1552 161 1553 165
rect 1547 160 1553 161
rect 1635 165 1641 166
rect 1635 161 1636 165
rect 1640 161 1641 165
rect 1803 165 1809 166
rect 1635 160 1641 161
rect 1715 163 1721 164
rect 1462 158 1473 159
rect 1715 159 1716 163
rect 1720 162 1721 163
rect 1778 163 1784 164
rect 1778 162 1779 163
rect 1720 160 1779 162
rect 1720 159 1721 160
rect 1715 158 1721 159
rect 1778 159 1779 160
rect 1783 159 1784 163
rect 1803 161 1804 165
rect 1808 161 1809 165
rect 1803 160 1809 161
rect 1891 165 1897 166
rect 1891 161 1892 165
rect 1896 161 1897 165
rect 2099 165 2105 166
rect 1891 160 1897 161
rect 1966 163 1972 164
rect 1778 158 1784 159
rect 1966 159 1967 163
rect 1971 162 1972 163
rect 1987 163 1993 164
rect 1987 162 1988 163
rect 1971 160 1988 162
rect 1971 159 1972 160
rect 1966 158 1972 159
rect 1987 159 1988 160
rect 1992 159 1993 163
rect 2099 161 2100 165
rect 2104 161 2105 165
rect 2099 160 2105 161
rect 2211 165 2246 166
rect 2211 161 2212 165
rect 2216 164 2246 165
rect 2216 161 2217 164
rect 2211 160 2217 161
rect 2326 163 2337 164
rect 1987 158 1993 159
rect 2326 159 2327 163
rect 2331 159 2332 163
rect 2336 159 2337 163
rect 2326 158 2337 159
rect 2435 163 2441 164
rect 2435 159 2436 163
rect 2440 162 2441 163
rect 2470 163 2476 164
rect 2470 162 2471 163
rect 2440 160 2471 162
rect 2440 159 2441 160
rect 2435 158 2441 159
rect 2470 159 2471 160
rect 2475 159 2476 163
rect 2470 158 2476 159
rect 131 143 137 144
rect 131 139 132 143
rect 136 142 137 143
rect 174 143 180 144
rect 136 140 170 142
rect 136 139 137 140
rect 131 138 137 139
rect 168 130 170 140
rect 174 139 175 143
rect 179 142 180 143
rect 187 143 193 144
rect 187 142 188 143
rect 179 140 188 142
rect 179 139 180 140
rect 174 138 180 139
rect 187 139 188 140
rect 192 139 193 143
rect 187 138 193 139
rect 243 143 249 144
rect 243 139 244 143
rect 248 142 249 143
rect 299 143 305 144
rect 248 140 286 142
rect 248 139 249 140
rect 243 138 249 139
rect 284 130 286 140
rect 299 139 300 143
rect 304 142 305 143
rect 355 143 361 144
rect 304 140 321 142
rect 304 139 305 140
rect 299 138 305 139
rect 319 134 321 140
rect 355 139 356 143
rect 360 142 361 143
rect 411 143 417 144
rect 360 140 406 142
rect 360 139 361 140
rect 355 138 361 139
rect 319 132 398 134
rect 168 128 282 130
rect 284 128 342 130
rect 280 126 282 128
rect 340 126 342 128
rect 396 126 398 132
rect 404 130 406 140
rect 411 139 412 143
rect 416 142 417 143
rect 466 143 473 144
rect 416 140 462 142
rect 416 139 417 140
rect 411 138 417 139
rect 460 130 462 140
rect 466 139 467 143
rect 472 139 473 143
rect 466 138 473 139
rect 510 143 516 144
rect 510 139 511 143
rect 515 142 516 143
rect 523 143 529 144
rect 523 142 524 143
rect 515 140 524 142
rect 515 139 516 140
rect 510 138 516 139
rect 523 139 524 140
rect 528 139 529 143
rect 523 138 529 139
rect 566 143 572 144
rect 566 139 567 143
rect 571 142 572 143
rect 579 143 585 144
rect 579 142 580 143
rect 571 140 580 142
rect 571 139 572 140
rect 566 138 572 139
rect 579 139 580 140
rect 584 139 585 143
rect 579 138 585 139
rect 635 143 641 144
rect 635 139 636 143
rect 640 142 641 143
rect 678 143 684 144
rect 640 140 674 142
rect 640 139 641 140
rect 635 138 641 139
rect 672 130 674 140
rect 678 139 679 143
rect 683 142 684 143
rect 691 143 697 144
rect 691 142 692 143
rect 683 140 692 142
rect 683 139 684 140
rect 678 138 684 139
rect 691 139 692 140
rect 696 139 697 143
rect 691 138 697 139
rect 734 143 740 144
rect 734 139 735 143
rect 739 142 740 143
rect 747 143 753 144
rect 747 142 748 143
rect 739 140 748 142
rect 739 139 740 140
rect 734 138 740 139
rect 747 139 748 140
rect 752 139 753 143
rect 747 138 753 139
rect 811 143 817 144
rect 811 139 812 143
rect 816 142 817 143
rect 875 143 881 144
rect 816 140 870 142
rect 816 139 817 140
rect 811 138 817 139
rect 868 130 870 140
rect 875 139 876 143
rect 880 142 881 143
rect 939 143 945 144
rect 880 140 934 142
rect 880 139 881 140
rect 875 138 881 139
rect 932 130 934 140
rect 939 139 940 143
rect 944 142 945 143
rect 1003 143 1009 144
rect 944 140 998 142
rect 944 139 945 140
rect 939 138 945 139
rect 996 130 998 140
rect 1003 139 1004 143
rect 1008 142 1009 143
rect 1067 143 1073 144
rect 1008 140 1062 142
rect 1008 139 1009 140
rect 1003 138 1009 139
rect 1060 130 1062 140
rect 1067 139 1068 143
rect 1072 142 1073 143
rect 1131 143 1140 144
rect 1072 140 1126 142
rect 1072 139 1073 140
rect 1067 138 1073 139
rect 1124 134 1126 140
rect 1131 139 1132 143
rect 1139 139 1140 143
rect 1131 138 1140 139
rect 1124 132 1161 134
rect 404 128 454 130
rect 460 128 622 130
rect 672 128 854 130
rect 868 128 918 130
rect 932 128 982 130
rect 996 128 1046 130
rect 1060 128 1110 130
rect 452 126 454 128
rect 620 126 622 128
rect 852 126 854 128
rect 916 126 918 128
rect 980 126 982 128
rect 1044 126 1046 128
rect 1108 126 1110 128
rect 1159 126 1161 132
rect 1347 131 1353 132
rect 1347 127 1348 131
rect 1352 130 1353 131
rect 1374 131 1380 132
rect 1374 130 1375 131
rect 1352 128 1375 130
rect 1352 127 1353 128
rect 1347 126 1353 127
rect 1374 127 1375 128
rect 1379 127 1380 131
rect 1374 126 1380 127
rect 1390 131 1396 132
rect 1390 127 1391 131
rect 1395 130 1396 131
rect 1403 131 1409 132
rect 1403 130 1404 131
rect 1395 128 1404 130
rect 1395 127 1396 128
rect 1390 126 1396 127
rect 1403 127 1404 128
rect 1408 127 1409 131
rect 1403 126 1409 127
rect 1446 131 1452 132
rect 1446 127 1447 131
rect 1451 130 1452 131
rect 1459 131 1465 132
rect 1459 130 1460 131
rect 1451 128 1460 130
rect 1451 127 1452 128
rect 1446 126 1452 127
rect 1459 127 1460 128
rect 1464 127 1465 131
rect 1459 126 1465 127
rect 1502 131 1508 132
rect 1502 127 1503 131
rect 1507 130 1508 131
rect 1515 131 1521 132
rect 1515 130 1516 131
rect 1507 128 1516 130
rect 1507 127 1508 128
rect 1502 126 1508 127
rect 1515 127 1516 128
rect 1520 127 1521 131
rect 1515 126 1521 127
rect 1558 131 1564 132
rect 1558 127 1559 131
rect 1563 130 1564 131
rect 1571 131 1577 132
rect 1571 130 1572 131
rect 1563 128 1572 130
rect 1563 127 1564 128
rect 1558 126 1564 127
rect 1571 127 1572 128
rect 1576 127 1577 131
rect 1571 126 1577 127
rect 1614 131 1620 132
rect 1614 127 1615 131
rect 1619 130 1620 131
rect 1627 131 1633 132
rect 1627 130 1628 131
rect 1619 128 1628 130
rect 1619 127 1620 128
rect 1614 126 1620 127
rect 1627 127 1628 128
rect 1632 127 1633 131
rect 1627 126 1633 127
rect 1670 131 1676 132
rect 1670 127 1671 131
rect 1675 130 1676 131
rect 1683 131 1689 132
rect 1683 130 1684 131
rect 1675 128 1684 130
rect 1675 127 1676 128
rect 1670 126 1676 127
rect 1683 127 1684 128
rect 1688 127 1689 131
rect 1683 126 1689 127
rect 1726 131 1732 132
rect 1726 127 1727 131
rect 1731 130 1732 131
rect 1739 131 1745 132
rect 1739 130 1740 131
rect 1731 128 1740 130
rect 1731 127 1732 128
rect 1726 126 1732 127
rect 1739 127 1740 128
rect 1744 127 1745 131
rect 1739 126 1745 127
rect 1803 131 1809 132
rect 1803 127 1804 131
rect 1808 130 1809 131
rect 1846 131 1852 132
rect 1808 128 1842 130
rect 1808 127 1809 128
rect 1803 126 1809 127
rect 150 125 156 126
rect 110 124 116 125
rect 110 120 111 124
rect 115 120 116 124
rect 150 121 151 125
rect 155 121 156 125
rect 206 125 212 126
rect 150 120 156 121
rect 171 123 180 124
rect 110 119 116 120
rect 171 119 172 123
rect 179 119 180 123
rect 206 121 207 125
rect 211 121 212 125
rect 262 125 268 126
rect 206 120 212 121
rect 226 123 233 124
rect 171 118 180 119
rect 226 119 227 123
rect 232 119 233 123
rect 262 121 263 125
rect 267 121 268 125
rect 280 125 289 126
rect 280 124 284 125
rect 262 120 268 121
rect 283 121 284 124
rect 288 121 289 125
rect 283 120 289 121
rect 318 125 324 126
rect 318 121 319 125
rect 323 121 324 125
rect 318 120 324 121
rect 339 125 345 126
rect 339 121 340 125
rect 344 121 345 125
rect 339 120 345 121
rect 374 125 380 126
rect 374 121 375 125
rect 379 121 380 125
rect 374 120 380 121
rect 395 125 401 126
rect 395 121 396 125
rect 400 121 401 125
rect 395 120 401 121
rect 430 125 436 126
rect 430 121 431 125
rect 435 121 436 125
rect 430 120 436 121
rect 451 125 457 126
rect 451 121 452 125
rect 456 121 457 125
rect 451 120 457 121
rect 486 125 492 126
rect 486 121 487 125
rect 491 121 492 125
rect 542 125 548 126
rect 486 120 492 121
rect 507 123 516 124
rect 226 118 233 119
rect 507 119 508 123
rect 515 119 516 123
rect 542 121 543 125
rect 547 121 548 125
rect 598 125 604 126
rect 542 120 548 121
rect 563 123 572 124
rect 507 118 516 119
rect 563 119 564 123
rect 571 119 572 123
rect 598 121 599 125
rect 603 121 604 125
rect 598 120 604 121
rect 619 125 625 126
rect 619 121 620 125
rect 624 121 625 125
rect 619 120 625 121
rect 654 125 660 126
rect 654 121 655 125
rect 659 121 660 125
rect 710 125 716 126
rect 654 120 660 121
rect 675 123 684 124
rect 563 118 572 119
rect 675 119 676 123
rect 683 119 684 123
rect 710 121 711 125
rect 715 121 716 125
rect 766 125 772 126
rect 710 120 716 121
rect 731 123 740 124
rect 675 118 684 119
rect 731 119 732 123
rect 739 119 740 123
rect 766 121 767 125
rect 771 121 772 125
rect 830 125 836 126
rect 766 120 772 121
rect 787 123 796 124
rect 731 118 740 119
rect 787 119 788 123
rect 795 119 796 123
rect 830 121 831 125
rect 835 121 836 125
rect 830 120 836 121
rect 851 125 857 126
rect 851 121 852 125
rect 856 121 857 125
rect 851 120 857 121
rect 894 125 900 126
rect 894 121 895 125
rect 899 121 900 125
rect 894 120 900 121
rect 915 125 921 126
rect 915 121 916 125
rect 920 121 921 125
rect 915 120 921 121
rect 958 125 964 126
rect 958 121 959 125
rect 963 121 964 125
rect 958 120 964 121
rect 979 125 985 126
rect 979 121 980 125
rect 984 121 985 125
rect 979 120 985 121
rect 1022 125 1028 126
rect 1022 121 1023 125
rect 1027 121 1028 125
rect 1022 120 1028 121
rect 1043 125 1049 126
rect 1043 121 1044 125
rect 1048 121 1049 125
rect 1043 120 1049 121
rect 1086 125 1092 126
rect 1086 121 1087 125
rect 1091 121 1092 125
rect 1086 120 1092 121
rect 1107 125 1113 126
rect 1107 121 1108 125
rect 1112 121 1113 125
rect 1107 120 1113 121
rect 1150 125 1156 126
rect 1150 121 1151 125
rect 1155 121 1156 125
rect 1159 125 1177 126
rect 1159 124 1172 125
rect 1150 120 1156 121
rect 1171 121 1172 124
rect 1176 121 1177 125
rect 1171 120 1177 121
rect 1286 124 1292 125
rect 1286 120 1287 124
rect 1291 120 1292 124
rect 1286 119 1292 120
rect 787 118 796 119
rect 1840 118 1842 128
rect 1846 127 1847 131
rect 1851 130 1852 131
rect 1859 131 1865 132
rect 1859 130 1860 131
rect 1851 128 1860 130
rect 1851 127 1852 128
rect 1846 126 1852 127
rect 1859 127 1860 128
rect 1864 127 1865 131
rect 1859 126 1865 127
rect 1902 131 1908 132
rect 1902 127 1903 131
rect 1907 130 1908 131
rect 1923 131 1929 132
rect 1923 130 1924 131
rect 1907 128 1924 130
rect 1907 127 1908 128
rect 1902 126 1908 127
rect 1923 127 1924 128
rect 1928 127 1929 131
rect 1923 126 1929 127
rect 1987 131 1993 132
rect 1987 127 1988 131
rect 1992 130 1993 131
rect 2051 131 2057 132
rect 1992 128 2001 130
rect 1992 127 1993 128
rect 1987 126 1993 127
rect 1999 122 2001 128
rect 2051 127 2052 131
rect 2056 130 2057 131
rect 2123 131 2132 132
rect 2056 128 2118 130
rect 2056 127 2057 128
rect 2051 126 2057 127
rect 1999 120 2094 122
rect 1840 116 2030 118
rect 2028 114 2030 116
rect 2092 114 2094 120
rect 2116 118 2118 128
rect 2123 127 2124 131
rect 2131 127 2132 131
rect 2123 126 2132 127
rect 2166 131 2172 132
rect 2166 127 2167 131
rect 2171 130 2172 131
rect 2203 131 2209 132
rect 2203 130 2204 131
rect 2171 128 2204 130
rect 2171 127 2172 128
rect 2166 126 2172 127
rect 2203 127 2204 128
rect 2208 127 2209 131
rect 2203 126 2209 127
rect 2246 131 2252 132
rect 2246 127 2247 131
rect 2251 130 2252 131
rect 2283 131 2289 132
rect 2283 130 2284 131
rect 2251 128 2284 130
rect 2251 127 2252 128
rect 2246 126 2252 127
rect 2283 127 2284 128
rect 2288 127 2289 131
rect 2283 126 2289 127
rect 2371 131 2377 132
rect 2371 127 2372 131
rect 2376 130 2377 131
rect 2435 131 2441 132
rect 2376 128 2430 130
rect 2376 127 2377 128
rect 2371 126 2377 127
rect 2428 118 2430 128
rect 2435 127 2436 131
rect 2440 130 2441 131
rect 2462 131 2468 132
rect 2462 130 2463 131
rect 2440 128 2463 130
rect 2440 127 2441 128
rect 2435 126 2441 127
rect 2462 127 2463 128
rect 2467 127 2468 131
rect 2462 126 2468 127
rect 2116 116 2326 118
rect 2428 116 2478 118
rect 2324 114 2326 116
rect 2476 114 2478 116
rect 1366 113 1372 114
rect 1326 112 1332 113
rect 1326 108 1327 112
rect 1331 108 1332 112
rect 1366 109 1367 113
rect 1371 109 1372 113
rect 1422 113 1428 114
rect 1366 108 1372 109
rect 1387 111 1396 112
rect 110 107 116 108
rect 110 103 111 107
rect 115 103 116 107
rect 1286 107 1292 108
rect 1326 107 1332 108
rect 1387 107 1388 111
rect 1395 107 1396 111
rect 1422 109 1423 113
rect 1427 109 1428 113
rect 1478 113 1484 114
rect 1422 108 1428 109
rect 1443 111 1452 112
rect 110 102 116 103
rect 134 104 140 105
rect 134 100 135 104
rect 139 100 140 104
rect 134 99 140 100
rect 190 104 196 105
rect 190 100 191 104
rect 195 100 196 104
rect 190 99 196 100
rect 246 104 252 105
rect 246 100 247 104
rect 251 100 252 104
rect 246 99 252 100
rect 302 104 308 105
rect 302 100 303 104
rect 307 100 308 104
rect 302 99 308 100
rect 358 104 364 105
rect 358 100 359 104
rect 363 100 364 104
rect 358 99 364 100
rect 414 104 420 105
rect 414 100 415 104
rect 419 100 420 104
rect 414 99 420 100
rect 470 104 476 105
rect 470 100 471 104
rect 475 100 476 104
rect 470 99 476 100
rect 526 104 532 105
rect 526 100 527 104
rect 531 100 532 104
rect 526 99 532 100
rect 582 104 588 105
rect 582 100 583 104
rect 587 100 588 104
rect 582 99 588 100
rect 638 104 644 105
rect 638 100 639 104
rect 643 100 644 104
rect 638 99 644 100
rect 694 104 700 105
rect 694 100 695 104
rect 699 100 700 104
rect 694 99 700 100
rect 750 104 756 105
rect 750 100 751 104
rect 755 100 756 104
rect 750 99 756 100
rect 814 104 820 105
rect 814 100 815 104
rect 819 100 820 104
rect 814 99 820 100
rect 878 104 884 105
rect 878 100 879 104
rect 883 100 884 104
rect 878 99 884 100
rect 942 104 948 105
rect 942 100 943 104
rect 947 100 948 104
rect 942 99 948 100
rect 1006 104 1012 105
rect 1006 100 1007 104
rect 1011 100 1012 104
rect 1006 99 1012 100
rect 1070 104 1076 105
rect 1070 100 1071 104
rect 1075 100 1076 104
rect 1070 99 1076 100
rect 1134 104 1140 105
rect 1134 100 1135 104
rect 1139 100 1140 104
rect 1286 103 1287 107
rect 1291 103 1292 107
rect 1387 106 1396 107
rect 1443 107 1444 111
rect 1451 107 1452 111
rect 1478 109 1479 113
rect 1483 109 1484 113
rect 1534 113 1540 114
rect 1478 108 1484 109
rect 1499 111 1508 112
rect 1443 106 1452 107
rect 1499 107 1500 111
rect 1507 107 1508 111
rect 1534 109 1535 113
rect 1539 109 1540 113
rect 1590 113 1596 114
rect 1534 108 1540 109
rect 1555 111 1564 112
rect 1499 106 1508 107
rect 1555 107 1556 111
rect 1563 107 1564 111
rect 1590 109 1591 113
rect 1595 109 1596 113
rect 1646 113 1652 114
rect 1590 108 1596 109
rect 1611 111 1620 112
rect 1555 106 1564 107
rect 1611 107 1612 111
rect 1619 107 1620 111
rect 1646 109 1647 113
rect 1651 109 1652 113
rect 1702 113 1708 114
rect 1646 108 1652 109
rect 1667 111 1676 112
rect 1611 106 1620 107
rect 1667 107 1668 111
rect 1675 107 1676 111
rect 1702 109 1703 113
rect 1707 109 1708 113
rect 1758 113 1764 114
rect 1702 108 1708 109
rect 1723 111 1732 112
rect 1667 106 1676 107
rect 1723 107 1724 111
rect 1731 107 1732 111
rect 1758 109 1759 113
rect 1763 109 1764 113
rect 1822 113 1828 114
rect 1758 108 1764 109
rect 1778 111 1785 112
rect 1723 106 1732 107
rect 1778 107 1779 111
rect 1784 107 1785 111
rect 1822 109 1823 113
rect 1827 109 1828 113
rect 1878 113 1884 114
rect 1822 108 1828 109
rect 1843 111 1852 112
rect 1778 106 1785 107
rect 1843 107 1844 111
rect 1851 107 1852 111
rect 1878 109 1879 113
rect 1883 109 1884 113
rect 1942 113 1948 114
rect 1878 108 1884 109
rect 1899 111 1908 112
rect 1843 106 1852 107
rect 1899 107 1900 111
rect 1907 107 1908 111
rect 1942 109 1943 113
rect 1947 109 1948 113
rect 2006 113 2012 114
rect 1942 108 1948 109
rect 1963 111 1972 112
rect 1899 106 1908 107
rect 1963 107 1964 111
rect 1971 107 1972 111
rect 2006 109 2007 113
rect 2011 109 2012 113
rect 2006 108 2012 109
rect 2027 113 2033 114
rect 2027 109 2028 113
rect 2032 109 2033 113
rect 2027 108 2033 109
rect 2070 113 2076 114
rect 2070 109 2071 113
rect 2075 109 2076 113
rect 2070 108 2076 109
rect 2091 113 2097 114
rect 2091 109 2092 113
rect 2096 109 2097 113
rect 2091 108 2097 109
rect 2142 113 2148 114
rect 2142 109 2143 113
rect 2147 109 2148 113
rect 2222 113 2228 114
rect 2142 108 2148 109
rect 2163 111 2172 112
rect 1963 106 1972 107
rect 2163 107 2164 111
rect 2171 107 2172 111
rect 2222 109 2223 113
rect 2227 109 2228 113
rect 2302 113 2308 114
rect 2222 108 2228 109
rect 2243 111 2252 112
rect 2163 106 2172 107
rect 2243 107 2244 111
rect 2251 107 2252 111
rect 2302 109 2303 113
rect 2307 109 2308 113
rect 2302 108 2308 109
rect 2323 113 2329 114
rect 2323 109 2324 113
rect 2328 109 2329 113
rect 2323 108 2329 109
rect 2390 113 2396 114
rect 2390 109 2391 113
rect 2395 109 2396 113
rect 2390 108 2396 109
rect 2454 113 2460 114
rect 2454 109 2455 113
rect 2459 109 2460 113
rect 2454 108 2460 109
rect 2475 113 2481 114
rect 2475 109 2476 113
rect 2480 109 2481 113
rect 2475 108 2481 109
rect 2502 112 2508 113
rect 2502 108 2503 112
rect 2507 108 2508 112
rect 2502 107 2508 108
rect 2243 106 2252 107
rect 1286 102 1292 103
rect 1134 99 1140 100
rect 1326 95 1332 96
rect 1326 91 1327 95
rect 1331 91 1332 95
rect 2502 95 2508 96
rect 1326 90 1332 91
rect 1350 92 1356 93
rect 1350 88 1351 92
rect 1355 88 1356 92
rect 1350 87 1356 88
rect 1406 92 1412 93
rect 1406 88 1407 92
rect 1411 88 1412 92
rect 1406 87 1412 88
rect 1462 92 1468 93
rect 1462 88 1463 92
rect 1467 88 1468 92
rect 1462 87 1468 88
rect 1518 92 1524 93
rect 1518 88 1519 92
rect 1523 88 1524 92
rect 1518 87 1524 88
rect 1574 92 1580 93
rect 1574 88 1575 92
rect 1579 88 1580 92
rect 1574 87 1580 88
rect 1630 92 1636 93
rect 1630 88 1631 92
rect 1635 88 1636 92
rect 1630 87 1636 88
rect 1686 92 1692 93
rect 1686 88 1687 92
rect 1691 88 1692 92
rect 1686 87 1692 88
rect 1742 92 1748 93
rect 1742 88 1743 92
rect 1747 88 1748 92
rect 1742 87 1748 88
rect 1806 92 1812 93
rect 1806 88 1807 92
rect 1811 88 1812 92
rect 1806 87 1812 88
rect 1862 92 1868 93
rect 1862 88 1863 92
rect 1867 88 1868 92
rect 1862 87 1868 88
rect 1926 92 1932 93
rect 1926 88 1927 92
rect 1931 88 1932 92
rect 1926 87 1932 88
rect 1990 92 1996 93
rect 1990 88 1991 92
rect 1995 88 1996 92
rect 1990 87 1996 88
rect 2054 92 2060 93
rect 2054 88 2055 92
rect 2059 88 2060 92
rect 2054 87 2060 88
rect 2126 92 2132 93
rect 2126 88 2127 92
rect 2131 88 2132 92
rect 2126 87 2132 88
rect 2206 92 2212 93
rect 2206 88 2207 92
rect 2211 88 2212 92
rect 2206 87 2212 88
rect 2286 92 2292 93
rect 2286 88 2287 92
rect 2291 88 2292 92
rect 2286 87 2292 88
rect 2374 92 2380 93
rect 2374 88 2375 92
rect 2379 88 2380 92
rect 2374 87 2380 88
rect 2438 92 2444 93
rect 2438 88 2439 92
rect 2443 88 2444 92
rect 2502 91 2503 95
rect 2507 91 2508 95
rect 2502 90 2508 91
rect 2438 87 2444 88
<< m3c >>
rect 111 2569 115 2573
rect 135 2572 139 2576
rect 191 2572 195 2576
rect 247 2572 251 2576
rect 303 2572 307 2576
rect 359 2572 363 2576
rect 1287 2569 1291 2573
rect 111 2552 115 2556
rect 151 2551 155 2555
rect 187 2551 191 2555
rect 207 2551 211 2555
rect 243 2551 247 2555
rect 263 2551 267 2555
rect 299 2551 303 2555
rect 319 2551 323 2555
rect 355 2551 359 2555
rect 375 2551 379 2555
rect 1287 2552 1291 2556
rect 215 2543 219 2547
rect 1327 2549 1331 2553
rect 1495 2552 1499 2556
rect 1551 2552 1555 2556
rect 1607 2552 1611 2556
rect 1663 2552 1667 2556
rect 1719 2552 1723 2556
rect 1775 2552 1779 2556
rect 1831 2552 1835 2556
rect 1887 2552 1891 2556
rect 1943 2552 1947 2556
rect 1999 2552 2003 2556
rect 2055 2552 2059 2556
rect 2111 2552 2115 2556
rect 2167 2552 2171 2556
rect 2503 2549 2507 2553
rect 187 2531 188 2535
rect 188 2531 191 2535
rect 243 2531 244 2535
rect 244 2531 247 2535
rect 299 2531 300 2535
rect 300 2531 303 2535
rect 355 2531 356 2535
rect 356 2531 359 2535
rect 1327 2532 1331 2536
rect 1511 2531 1515 2535
rect 1535 2531 1536 2535
rect 1536 2531 1539 2535
rect 1567 2531 1571 2535
rect 1599 2531 1603 2535
rect 1623 2531 1627 2535
rect 1659 2531 1663 2535
rect 1679 2531 1683 2535
rect 1715 2531 1719 2535
rect 1735 2531 1739 2535
rect 1771 2531 1775 2535
rect 1791 2531 1795 2535
rect 1815 2531 1816 2535
rect 1816 2531 1819 2535
rect 1847 2531 1851 2535
rect 1883 2531 1887 2535
rect 1903 2531 1907 2535
rect 1939 2531 1943 2535
rect 1959 2531 1963 2535
rect 1995 2531 1999 2535
rect 2015 2531 2019 2535
rect 2051 2531 2055 2535
rect 2071 2531 2075 2535
rect 2103 2531 2107 2535
rect 2127 2531 2131 2535
rect 2163 2531 2167 2535
rect 2183 2531 2187 2535
rect 2191 2531 2195 2535
rect 2503 2532 2507 2536
rect 215 2519 219 2523
rect 247 2519 251 2523
rect 303 2519 307 2523
rect 367 2519 371 2523
rect 439 2519 443 2523
rect 567 2519 571 2523
rect 575 2519 579 2523
rect 639 2519 643 2523
rect 703 2519 707 2523
rect 763 2519 767 2523
rect 827 2519 831 2523
rect 891 2519 895 2523
rect 959 2519 963 2523
rect 1019 2519 1023 2523
rect 1527 2511 1531 2515
rect 1535 2511 1539 2515
rect 1599 2511 1603 2515
rect 1659 2511 1660 2515
rect 1660 2511 1663 2515
rect 1715 2511 1716 2515
rect 1716 2511 1719 2515
rect 1771 2511 1772 2515
rect 1772 2511 1775 2515
rect 1815 2511 1819 2515
rect 1883 2511 1884 2515
rect 1884 2511 1887 2515
rect 1939 2511 1940 2515
rect 1940 2511 1943 2515
rect 1995 2511 1996 2515
rect 1996 2511 1999 2515
rect 2051 2511 2052 2515
rect 2052 2511 2055 2515
rect 2103 2511 2107 2515
rect 2163 2511 2164 2515
rect 2164 2511 2167 2515
rect 111 2500 115 2504
rect 223 2501 227 2505
rect 247 2499 248 2503
rect 248 2499 251 2503
rect 279 2501 283 2505
rect 303 2499 304 2503
rect 304 2499 307 2503
rect 343 2501 347 2505
rect 367 2499 368 2503
rect 368 2499 371 2503
rect 415 2501 419 2505
rect 439 2499 440 2503
rect 440 2499 443 2503
rect 487 2501 491 2505
rect 495 2499 499 2503
rect 551 2501 555 2505
rect 575 2499 576 2503
rect 576 2499 579 2503
rect 615 2501 619 2505
rect 639 2499 640 2503
rect 640 2499 643 2503
rect 679 2501 683 2505
rect 703 2499 704 2503
rect 704 2499 707 2503
rect 743 2501 747 2505
rect 763 2499 764 2503
rect 764 2499 767 2503
rect 807 2501 811 2505
rect 827 2499 828 2503
rect 828 2499 831 2503
rect 871 2501 875 2505
rect 891 2499 892 2503
rect 892 2499 895 2503
rect 935 2501 939 2505
rect 959 2499 960 2503
rect 960 2499 963 2503
rect 999 2501 1003 2505
rect 1019 2499 1020 2503
rect 1020 2499 1023 2503
rect 1063 2501 1067 2505
rect 1071 2499 1075 2503
rect 1287 2500 1291 2504
rect 1567 2495 1571 2499
rect 1575 2499 1579 2503
rect 1631 2499 1635 2503
rect 1703 2499 1707 2503
rect 1775 2499 1779 2503
rect 1911 2499 1915 2503
rect 1919 2499 1923 2503
rect 1991 2499 1995 2503
rect 2063 2499 2067 2503
rect 2135 2499 2139 2503
rect 111 2483 115 2487
rect 207 2480 211 2484
rect 263 2480 267 2484
rect 327 2480 331 2484
rect 399 2480 403 2484
rect 471 2480 475 2484
rect 535 2480 539 2484
rect 599 2480 603 2484
rect 663 2480 667 2484
rect 727 2480 731 2484
rect 791 2480 795 2484
rect 855 2480 859 2484
rect 919 2480 923 2484
rect 983 2480 987 2484
rect 1047 2480 1051 2484
rect 1287 2483 1291 2487
rect 1327 2480 1331 2484
rect 1543 2481 1547 2485
rect 1575 2479 1579 2483
rect 1607 2481 1611 2485
rect 1631 2479 1632 2483
rect 1632 2479 1635 2483
rect 1679 2481 1683 2485
rect 1703 2479 1704 2483
rect 1704 2479 1707 2483
rect 1751 2481 1755 2485
rect 1775 2479 1776 2483
rect 1776 2479 1779 2483
rect 1823 2481 1827 2485
rect 1843 2479 1844 2483
rect 1844 2479 1847 2483
rect 1895 2481 1899 2485
rect 1919 2479 1920 2483
rect 1920 2479 1923 2483
rect 1967 2481 1971 2485
rect 1991 2479 1992 2483
rect 1992 2479 1995 2483
rect 2039 2481 2043 2485
rect 2063 2479 2064 2483
rect 2064 2479 2067 2483
rect 2111 2481 2115 2485
rect 2135 2479 2136 2483
rect 2136 2479 2139 2483
rect 2183 2481 2187 2485
rect 2191 2479 2195 2483
rect 2503 2480 2507 2484
rect 111 2457 115 2461
rect 167 2460 171 2464
rect 223 2460 227 2464
rect 279 2460 283 2464
rect 335 2460 339 2464
rect 391 2460 395 2464
rect 447 2460 451 2464
rect 503 2460 507 2464
rect 559 2460 563 2464
rect 615 2460 619 2464
rect 671 2460 675 2464
rect 727 2460 731 2464
rect 783 2460 787 2464
rect 839 2460 843 2464
rect 895 2460 899 2464
rect 951 2460 955 2464
rect 1007 2460 1011 2464
rect 1063 2460 1067 2464
rect 1327 2463 1331 2467
rect 1287 2457 1291 2461
rect 1527 2460 1531 2464
rect 1591 2460 1595 2464
rect 1663 2460 1667 2464
rect 1735 2460 1739 2464
rect 1807 2460 1811 2464
rect 1879 2460 1883 2464
rect 1951 2460 1955 2464
rect 2023 2460 2027 2464
rect 2095 2460 2099 2464
rect 2167 2460 2171 2464
rect 2503 2463 2507 2467
rect 111 2440 115 2444
rect 183 2439 187 2443
rect 219 2439 223 2443
rect 239 2439 243 2443
rect 275 2439 279 2443
rect 295 2439 299 2443
rect 331 2439 335 2443
rect 351 2439 355 2443
rect 387 2439 391 2443
rect 407 2439 411 2443
rect 443 2439 447 2443
rect 463 2439 467 2443
rect 499 2439 503 2443
rect 519 2439 523 2443
rect 555 2439 559 2443
rect 575 2439 579 2443
rect 611 2439 615 2443
rect 631 2439 635 2443
rect 667 2439 671 2443
rect 687 2439 691 2443
rect 723 2439 727 2443
rect 743 2439 747 2443
rect 779 2439 783 2443
rect 799 2439 803 2443
rect 835 2439 839 2443
rect 855 2439 859 2443
rect 875 2439 876 2443
rect 876 2439 879 2443
rect 911 2439 915 2443
rect 919 2439 923 2443
rect 967 2439 971 2443
rect 975 2439 979 2443
rect 1023 2439 1027 2443
rect 1079 2439 1083 2443
rect 1287 2440 1291 2444
rect 1327 2441 1331 2445
rect 1543 2444 1547 2448
rect 1607 2444 1611 2448
rect 1671 2444 1675 2448
rect 1743 2444 1747 2448
rect 1815 2444 1819 2448
rect 1879 2444 1883 2448
rect 1951 2444 1955 2448
rect 2023 2444 2027 2448
rect 2095 2444 2099 2448
rect 2167 2444 2171 2448
rect 2503 2441 2507 2445
rect 167 2419 168 2423
rect 168 2419 171 2423
rect 219 2419 220 2423
rect 220 2419 223 2423
rect 275 2419 276 2423
rect 276 2419 279 2423
rect 331 2419 332 2423
rect 332 2419 335 2423
rect 387 2419 388 2423
rect 388 2419 391 2423
rect 443 2419 444 2423
rect 444 2419 447 2423
rect 499 2419 500 2423
rect 500 2419 503 2423
rect 555 2419 556 2423
rect 556 2419 559 2423
rect 611 2419 612 2423
rect 612 2419 615 2423
rect 667 2419 668 2423
rect 668 2419 671 2423
rect 723 2419 724 2423
rect 724 2419 727 2423
rect 779 2419 780 2423
rect 780 2419 783 2423
rect 835 2419 836 2423
rect 836 2419 839 2423
rect 1327 2424 1331 2428
rect 975 2415 979 2419
rect 1559 2423 1563 2427
rect 1071 2419 1075 2423
rect 1567 2423 1571 2427
rect 1623 2423 1627 2427
rect 1687 2423 1691 2427
rect 1759 2423 1763 2427
rect 1831 2423 1835 2427
rect 1895 2423 1899 2427
rect 1947 2423 1951 2427
rect 1967 2423 1971 2427
rect 1975 2423 1979 2427
rect 2039 2423 2043 2427
rect 2055 2423 2059 2427
rect 2111 2423 2115 2427
rect 2183 2423 2187 2427
rect 2503 2424 2507 2428
rect 1811 2403 1812 2407
rect 1812 2403 1815 2407
rect 919 2395 923 2399
rect 1947 2403 1948 2407
rect 1948 2403 1951 2407
rect 2191 2403 2195 2407
rect 2055 2395 2059 2399
rect 1591 2387 1595 2391
rect 1647 2387 1651 2391
rect 1703 2387 1707 2391
rect 1767 2387 1771 2391
rect 111 2376 115 2380
rect 519 2377 523 2381
rect 543 2375 544 2379
rect 544 2375 547 2379
rect 575 2377 579 2381
rect 631 2377 635 2381
rect 687 2377 691 2381
rect 1287 2376 1291 2380
rect 1783 2379 1787 2383
rect 1975 2387 1979 2391
rect 2007 2387 2011 2391
rect 2071 2387 2075 2391
rect 1327 2368 1331 2372
rect 1567 2369 1571 2373
rect 1591 2367 1592 2371
rect 1592 2367 1595 2371
rect 1623 2369 1627 2373
rect 1647 2367 1648 2371
rect 1648 2367 1651 2371
rect 1679 2369 1683 2373
rect 1703 2367 1704 2371
rect 1704 2367 1707 2371
rect 1735 2369 1739 2373
rect 1767 2367 1771 2371
rect 1791 2369 1795 2373
rect 1811 2367 1812 2371
rect 1812 2367 1815 2371
rect 1855 2369 1859 2373
rect 1863 2367 1867 2371
rect 1919 2369 1923 2373
rect 1983 2369 1987 2373
rect 2007 2367 2008 2371
rect 2008 2367 2011 2371
rect 2047 2369 2051 2373
rect 2071 2367 2072 2371
rect 2072 2367 2075 2371
rect 2111 2369 2115 2373
rect 2503 2368 2507 2372
rect 111 2359 115 2363
rect 503 2356 507 2360
rect 559 2356 563 2360
rect 615 2356 619 2360
rect 671 2356 675 2360
rect 1287 2359 1291 2363
rect 1327 2351 1331 2355
rect 1551 2348 1555 2352
rect 1607 2348 1611 2352
rect 1663 2348 1667 2352
rect 1719 2348 1723 2352
rect 1775 2348 1779 2352
rect 1839 2348 1843 2352
rect 1903 2348 1907 2352
rect 1967 2348 1971 2352
rect 2031 2348 2035 2352
rect 2095 2348 2099 2352
rect 2503 2351 2507 2355
rect 111 2333 115 2337
rect 319 2336 323 2340
rect 391 2336 395 2340
rect 463 2336 467 2340
rect 535 2336 539 2340
rect 607 2336 611 2340
rect 679 2336 683 2340
rect 743 2336 747 2340
rect 807 2336 811 2340
rect 863 2336 867 2340
rect 927 2336 931 2340
rect 991 2336 995 2340
rect 1055 2336 1059 2340
rect 1111 2336 1115 2340
rect 1167 2336 1171 2340
rect 1223 2336 1227 2340
rect 1287 2333 1291 2337
rect 1327 2325 1331 2329
rect 1471 2328 1475 2332
rect 1535 2328 1539 2332
rect 1607 2328 1611 2332
rect 1687 2328 1691 2332
rect 1759 2328 1763 2332
rect 1831 2328 1835 2332
rect 1903 2328 1907 2332
rect 1983 2328 1987 2332
rect 2063 2328 2067 2332
rect 2143 2328 2147 2332
rect 2503 2325 2507 2329
rect 111 2316 115 2320
rect 335 2315 339 2319
rect 387 2315 391 2319
rect 407 2315 411 2319
rect 459 2315 463 2319
rect 479 2315 483 2319
rect 551 2315 555 2319
rect 623 2315 627 2319
rect 675 2315 679 2319
rect 695 2315 699 2319
rect 711 2315 715 2319
rect 759 2315 763 2319
rect 767 2315 771 2319
rect 823 2315 827 2319
rect 879 2315 883 2319
rect 943 2315 947 2319
rect 1007 2315 1011 2319
rect 1071 2315 1075 2319
rect 1079 2315 1083 2319
rect 1127 2315 1131 2319
rect 1183 2315 1187 2319
rect 1239 2315 1243 2319
rect 1287 2316 1291 2320
rect 1327 2308 1331 2312
rect 1487 2307 1491 2311
rect 1531 2307 1535 2311
rect 1551 2307 1555 2311
rect 1603 2307 1607 2311
rect 1623 2307 1627 2311
rect 1679 2307 1683 2311
rect 1703 2307 1707 2311
rect 1755 2307 1759 2311
rect 1775 2307 1779 2311
rect 1783 2307 1787 2311
rect 1847 2307 1851 2311
rect 1895 2307 1899 2311
rect 1919 2307 1923 2311
rect 1979 2307 1983 2311
rect 1999 2307 2003 2311
rect 2059 2307 2063 2311
rect 2079 2307 2083 2311
rect 2139 2307 2143 2311
rect 2159 2307 2163 2311
rect 387 2295 388 2299
rect 388 2295 391 2299
rect 543 2295 547 2299
rect 675 2295 676 2299
rect 676 2295 679 2299
rect 767 2287 771 2291
rect 1079 2291 1083 2295
rect 1259 2295 1263 2299
rect 1887 2299 1891 2303
rect 2503 2308 2507 2312
rect 1523 2287 1527 2291
rect 1531 2287 1532 2291
rect 1532 2287 1535 2291
rect 1603 2287 1604 2291
rect 1604 2287 1607 2291
rect 1679 2287 1683 2291
rect 1755 2287 1756 2291
rect 1756 2287 1759 2291
rect 1863 2287 1867 2291
rect 1895 2287 1899 2291
rect 1979 2287 1980 2291
rect 1980 2287 1983 2291
rect 2059 2287 2060 2291
rect 2060 2287 2063 2291
rect 2139 2287 2140 2291
rect 2140 2287 2143 2291
rect 459 2275 460 2279
rect 460 2275 463 2279
rect 503 2275 507 2279
rect 711 2275 715 2279
rect 727 2275 731 2279
rect 831 2275 835 2279
rect 1039 2275 1043 2279
rect 1151 2275 1155 2279
rect 1399 2275 1403 2279
rect 1407 2275 1411 2279
rect 1503 2275 1507 2279
rect 1607 2275 1611 2279
rect 1711 2275 1715 2279
rect 1887 2275 1888 2279
rect 1888 2275 1891 2279
rect 1927 2275 1931 2279
rect 2039 2275 2043 2279
rect 2151 2275 2155 2279
rect 1075 2267 1079 2271
rect 1523 2263 1527 2267
rect 111 2256 115 2260
rect 175 2257 179 2261
rect 183 2255 187 2259
rect 271 2257 275 2261
rect 375 2257 379 2261
rect 479 2257 483 2261
rect 503 2255 504 2259
rect 504 2255 507 2259
rect 591 2257 595 2261
rect 703 2257 707 2261
rect 727 2255 728 2259
rect 728 2255 731 2259
rect 807 2257 811 2261
rect 831 2255 832 2259
rect 832 2255 835 2259
rect 911 2257 915 2261
rect 927 2255 931 2259
rect 1015 2257 1019 2261
rect 1039 2255 1040 2259
rect 1040 2255 1043 2259
rect 1127 2257 1131 2261
rect 1151 2255 1152 2259
rect 1152 2255 1155 2259
rect 1239 2257 1243 2261
rect 1259 2255 1260 2259
rect 1260 2255 1263 2259
rect 1287 2256 1291 2260
rect 1327 2256 1331 2260
rect 1383 2257 1387 2261
rect 1407 2255 1408 2259
rect 1408 2255 1411 2259
rect 1479 2257 1483 2261
rect 1503 2255 1504 2259
rect 1504 2255 1507 2259
rect 1583 2257 1587 2261
rect 1607 2255 1608 2259
rect 1608 2255 1611 2259
rect 1687 2257 1691 2261
rect 1711 2255 1712 2259
rect 1712 2255 1715 2259
rect 1791 2257 1795 2261
rect 1903 2257 1907 2261
rect 1927 2255 1928 2259
rect 1928 2255 1931 2259
rect 2015 2257 2019 2261
rect 2039 2255 2040 2259
rect 2040 2255 2043 2259
rect 2127 2257 2131 2261
rect 2151 2255 2152 2259
rect 2152 2255 2155 2259
rect 2239 2257 2243 2261
rect 2247 2255 2251 2259
rect 2503 2256 2507 2260
rect 111 2239 115 2243
rect 159 2236 163 2240
rect 255 2236 259 2240
rect 359 2236 363 2240
rect 463 2236 467 2240
rect 575 2236 579 2240
rect 687 2236 691 2240
rect 791 2236 795 2240
rect 895 2236 899 2240
rect 999 2236 1003 2240
rect 1111 2236 1115 2240
rect 1223 2236 1227 2240
rect 1287 2239 1291 2243
rect 1327 2239 1331 2243
rect 1367 2236 1371 2240
rect 1463 2236 1467 2240
rect 1567 2236 1571 2240
rect 1671 2236 1675 2240
rect 1775 2236 1779 2240
rect 1887 2236 1891 2240
rect 1999 2236 2003 2240
rect 2111 2236 2115 2240
rect 2223 2236 2227 2240
rect 2503 2239 2507 2243
rect 111 2221 115 2225
rect 143 2224 147 2228
rect 231 2224 235 2228
rect 319 2224 323 2228
rect 415 2224 419 2228
rect 519 2224 523 2228
rect 623 2224 627 2228
rect 727 2224 731 2228
rect 831 2224 835 2228
rect 935 2224 939 2228
rect 1039 2224 1043 2228
rect 1143 2224 1147 2228
rect 1223 2224 1227 2228
rect 1287 2221 1291 2225
rect 1327 2221 1331 2225
rect 1367 2224 1371 2228
rect 1487 2224 1491 2228
rect 1607 2224 1611 2228
rect 1719 2224 1723 2228
rect 1815 2224 1819 2228
rect 1903 2224 1907 2228
rect 1983 2224 1987 2228
rect 2055 2224 2059 2228
rect 2127 2224 2131 2228
rect 2191 2224 2195 2228
rect 2255 2224 2259 2228
rect 2319 2224 2323 2228
rect 2383 2224 2387 2228
rect 2439 2224 2443 2228
rect 2503 2221 2507 2225
rect 111 2204 115 2208
rect 159 2203 163 2207
rect 227 2203 231 2207
rect 247 2203 251 2207
rect 315 2203 319 2207
rect 335 2203 339 2207
rect 411 2203 415 2207
rect 431 2203 435 2207
rect 515 2203 519 2207
rect 535 2203 539 2207
rect 239 2195 243 2199
rect 639 2203 643 2207
rect 647 2203 651 2207
rect 743 2203 747 2207
rect 751 2203 755 2207
rect 847 2203 851 2207
rect 951 2203 955 2207
rect 1055 2203 1059 2207
rect 1075 2203 1076 2207
rect 1076 2203 1079 2207
rect 1159 2203 1163 2207
rect 1219 2203 1223 2207
rect 1239 2203 1243 2207
rect 1287 2204 1291 2208
rect 1327 2204 1331 2208
rect 1383 2203 1387 2207
rect 1399 2203 1403 2207
rect 1503 2203 1507 2207
rect 1603 2203 1607 2207
rect 1623 2203 1627 2207
rect 1735 2203 1739 2207
rect 1811 2203 1815 2207
rect 1831 2203 1835 2207
rect 1899 2203 1903 2207
rect 1919 2203 1923 2207
rect 1979 2203 1983 2207
rect 1999 2203 2003 2207
rect 2051 2203 2055 2207
rect 2071 2203 2075 2207
rect 2123 2203 2127 2207
rect 2143 2203 2147 2207
rect 2187 2203 2191 2207
rect 2207 2203 2211 2207
rect 2251 2203 2255 2207
rect 2271 2203 2275 2207
rect 2315 2203 2319 2207
rect 2335 2203 2339 2207
rect 2379 2203 2383 2207
rect 2399 2203 2403 2207
rect 2435 2203 2439 2207
rect 2455 2203 2459 2207
rect 2463 2203 2467 2207
rect 2503 2204 2507 2208
rect 183 2183 187 2187
rect 227 2183 228 2187
rect 228 2183 231 2187
rect 315 2183 316 2187
rect 316 2183 319 2187
rect 411 2183 412 2187
rect 412 2183 415 2187
rect 515 2183 516 2187
rect 516 2183 519 2187
rect 751 2179 755 2183
rect 927 2183 931 2187
rect 1079 2183 1083 2187
rect 1219 2183 1220 2187
rect 1220 2183 1223 2187
rect 1431 2183 1435 2187
rect 1603 2183 1604 2187
rect 1604 2183 1607 2187
rect 1719 2183 1720 2187
rect 1720 2183 1723 2187
rect 1811 2183 1812 2187
rect 1812 2183 1815 2187
rect 1899 2183 1900 2187
rect 1900 2183 1903 2187
rect 1979 2183 1980 2187
rect 1980 2183 1983 2187
rect 2051 2183 2052 2187
rect 2052 2183 2055 2187
rect 2123 2183 2124 2187
rect 2124 2183 2127 2187
rect 2187 2183 2188 2187
rect 2188 2183 2191 2187
rect 2251 2183 2252 2187
rect 2252 2183 2255 2187
rect 2315 2183 2316 2187
rect 2316 2183 2319 2187
rect 2379 2183 2380 2187
rect 2380 2183 2383 2187
rect 2435 2183 2436 2187
rect 2436 2183 2439 2187
rect 239 2171 240 2175
rect 240 2171 243 2175
rect 279 2171 283 2175
rect 375 2171 379 2175
rect 479 2171 483 2175
rect 647 2171 648 2175
rect 648 2171 651 2175
rect 687 2171 691 2175
rect 791 2171 795 2175
rect 887 2171 891 2175
rect 1259 2171 1263 2175
rect 111 2152 115 2156
rect 255 2153 259 2157
rect 279 2151 280 2155
rect 280 2151 283 2155
rect 351 2153 355 2157
rect 375 2151 376 2155
rect 376 2151 379 2155
rect 455 2153 459 2157
rect 479 2151 480 2155
rect 480 2151 483 2155
rect 559 2153 563 2157
rect 567 2151 571 2155
rect 663 2153 667 2157
rect 687 2151 688 2155
rect 688 2151 691 2155
rect 767 2153 771 2157
rect 791 2151 792 2155
rect 792 2151 795 2155
rect 863 2153 867 2157
rect 887 2151 888 2155
rect 888 2151 891 2155
rect 959 2153 963 2157
rect 983 2151 984 2155
rect 984 2151 987 2155
rect 1055 2153 1059 2157
rect 1079 2151 1080 2155
rect 1080 2151 1083 2155
rect 1159 2153 1163 2157
rect 1239 2153 1243 2157
rect 1287 2152 1291 2156
rect 1747 2151 1751 2155
rect 1839 2151 1843 2155
rect 2463 2151 2467 2155
rect 111 2135 115 2139
rect 239 2132 243 2136
rect 335 2132 339 2136
rect 439 2132 443 2136
rect 543 2132 547 2136
rect 647 2132 651 2136
rect 751 2132 755 2136
rect 847 2132 851 2136
rect 943 2132 947 2136
rect 1039 2132 1043 2136
rect 1143 2132 1147 2136
rect 1223 2132 1227 2136
rect 1287 2135 1291 2139
rect 1327 2132 1331 2136
rect 1407 2133 1411 2137
rect 1431 2131 1432 2135
rect 1432 2131 1435 2135
rect 1623 2133 1627 2137
rect 1815 2133 1819 2137
rect 1839 2131 1840 2135
rect 1840 2131 1843 2135
rect 1991 2133 1995 2137
rect 2111 2131 2115 2135
rect 2159 2133 2163 2137
rect 2319 2133 2323 2137
rect 2455 2133 2459 2137
rect 2503 2132 2507 2136
rect 111 2117 115 2121
rect 303 2120 307 2124
rect 359 2120 363 2124
rect 423 2120 427 2124
rect 487 2120 491 2124
rect 559 2120 563 2124
rect 631 2120 635 2124
rect 711 2120 715 2124
rect 799 2120 803 2124
rect 887 2120 891 2124
rect 975 2120 979 2124
rect 1063 2120 1067 2124
rect 1151 2120 1155 2124
rect 1223 2120 1227 2124
rect 1287 2117 1291 2121
rect 1327 2115 1331 2119
rect 1391 2112 1395 2116
rect 1607 2112 1611 2116
rect 1799 2112 1803 2116
rect 1975 2112 1979 2116
rect 2143 2112 2147 2116
rect 2303 2112 2307 2116
rect 2439 2112 2443 2116
rect 2503 2115 2507 2119
rect 111 2100 115 2104
rect 319 2099 323 2103
rect 355 2099 359 2103
rect 375 2099 379 2103
rect 419 2099 423 2103
rect 439 2099 443 2103
rect 483 2099 487 2103
rect 503 2099 507 2103
rect 555 2099 559 2103
rect 575 2099 579 2103
rect 627 2099 631 2103
rect 647 2099 651 2103
rect 655 2099 659 2103
rect 727 2099 731 2103
rect 795 2099 799 2103
rect 815 2099 819 2103
rect 839 2099 840 2103
rect 840 2099 843 2103
rect 903 2099 907 2103
rect 991 2099 995 2103
rect 567 2087 571 2091
rect 1079 2099 1083 2103
rect 1147 2099 1151 2103
rect 1167 2099 1171 2103
rect 1219 2099 1223 2103
rect 1239 2099 1243 2103
rect 1259 2099 1260 2103
rect 1260 2099 1263 2103
rect 1287 2100 1291 2104
rect 1327 2097 1331 2101
rect 1383 2100 1387 2104
rect 1551 2100 1555 2104
rect 1711 2100 1715 2104
rect 1855 2100 1859 2104
rect 1991 2100 1995 2104
rect 2119 2100 2123 2104
rect 2239 2100 2243 2104
rect 2367 2100 2371 2104
rect 2503 2097 2507 2101
rect 355 2079 356 2083
rect 356 2079 359 2083
rect 419 2079 420 2083
rect 420 2079 423 2083
rect 483 2079 484 2083
rect 484 2079 487 2083
rect 555 2079 556 2083
rect 556 2079 559 2083
rect 627 2079 628 2083
rect 628 2079 631 2083
rect 795 2079 796 2083
rect 796 2079 799 2083
rect 983 2079 987 2083
rect 1111 2079 1115 2083
rect 1147 2079 1148 2083
rect 1148 2079 1151 2083
rect 1219 2079 1220 2083
rect 1220 2079 1223 2083
rect 1327 2080 1331 2084
rect 1399 2079 1403 2083
rect 1547 2079 1551 2083
rect 1567 2079 1571 2083
rect 1707 2079 1711 2083
rect 1727 2079 1731 2083
rect 1747 2079 1748 2083
rect 1748 2079 1751 2083
rect 1871 2079 1875 2083
rect 1907 2079 1911 2083
rect 2007 2079 2011 2083
rect 475 2071 479 2075
rect 2135 2079 2139 2083
rect 2235 2079 2239 2083
rect 2255 2079 2259 2083
rect 2363 2079 2367 2083
rect 2383 2079 2387 2083
rect 655 2063 659 2067
rect 839 2063 843 2067
rect 999 2063 1003 2067
rect 1127 2063 1131 2067
rect 1207 2063 1211 2067
rect 2503 2080 2507 2084
rect 1467 2059 1471 2063
rect 1547 2059 1548 2063
rect 1548 2059 1551 2063
rect 1707 2059 1708 2063
rect 1708 2059 1711 2063
rect 2111 2059 2115 2063
rect 2235 2059 2236 2063
rect 2236 2059 2239 2063
rect 2363 2059 2364 2063
rect 2364 2059 2367 2063
rect 1111 2051 1115 2055
rect 111 2044 115 2048
rect 399 2045 403 2049
rect 431 2043 435 2047
rect 455 2045 459 2049
rect 475 2043 476 2047
rect 476 2043 479 2047
rect 511 2045 515 2049
rect 575 2045 579 2049
rect 639 2045 643 2049
rect 711 2045 715 2049
rect 727 2043 731 2047
rect 791 2045 795 2049
rect 863 2045 867 2049
rect 943 2045 947 2049
rect 1023 2045 1027 2049
rect 1103 2045 1107 2049
rect 1127 2043 1128 2047
rect 1128 2043 1131 2047
rect 1183 2045 1187 2049
rect 1207 2043 1208 2047
rect 1208 2043 1211 2047
rect 1239 2045 1243 2049
rect 1287 2044 1291 2048
rect 1543 2043 1547 2047
rect 1575 2043 1579 2047
rect 1907 2043 1908 2047
rect 1908 2043 1911 2047
rect 1951 2043 1955 2047
rect 2047 2043 2051 2047
rect 111 2027 115 2031
rect 383 2024 387 2028
rect 439 2024 443 2028
rect 495 2024 499 2028
rect 559 2024 563 2028
rect 623 2024 627 2028
rect 695 2024 699 2028
rect 775 2024 779 2028
rect 847 2024 851 2028
rect 927 2024 931 2028
rect 1007 2024 1011 2028
rect 1087 2024 1091 2028
rect 1167 2024 1171 2028
rect 1223 2024 1227 2028
rect 1287 2027 1291 2031
rect 1327 2024 1331 2028
rect 1447 2025 1451 2029
rect 1467 2023 1468 2027
rect 1468 2023 1471 2027
rect 1551 2025 1555 2029
rect 1575 2023 1576 2027
rect 1576 2023 1579 2027
rect 1655 2025 1659 2029
rect 1751 2025 1755 2029
rect 1775 2023 1776 2027
rect 1776 2023 1779 2027
rect 1839 2025 1843 2029
rect 1927 2025 1931 2029
rect 1951 2023 1952 2027
rect 1952 2023 1955 2027
rect 2023 2025 2027 2029
rect 2047 2023 2048 2027
rect 2048 2023 2051 2027
rect 2119 2025 2123 2029
rect 2503 2024 2507 2028
rect 111 2005 115 2009
rect 231 2008 235 2012
rect 287 2008 291 2012
rect 359 2008 363 2012
rect 439 2008 443 2012
rect 535 2008 539 2012
rect 631 2008 635 2012
rect 735 2008 739 2012
rect 847 2008 851 2012
rect 959 2008 963 2012
rect 1079 2008 1083 2012
rect 1199 2008 1203 2012
rect 1287 2005 1291 2009
rect 1327 2007 1331 2011
rect 1431 2004 1435 2008
rect 1535 2004 1539 2008
rect 1639 2004 1643 2008
rect 1735 2004 1739 2008
rect 1823 2004 1827 2008
rect 1911 2004 1915 2008
rect 2007 2004 2011 2008
rect 2103 2004 2107 2008
rect 2503 2007 2507 2011
rect 111 1988 115 1992
rect 247 1987 251 1991
rect 283 1987 287 1991
rect 303 1987 307 1991
rect 355 1987 359 1991
rect 375 1987 379 1991
rect 419 1987 423 1991
rect 455 1987 459 1991
rect 531 1987 535 1991
rect 551 1987 555 1991
rect 627 1987 631 1991
rect 647 1987 651 1991
rect 655 1987 659 1991
rect 751 1987 755 1991
rect 843 1987 847 1991
rect 863 1987 867 1991
rect 899 1987 903 1991
rect 975 1987 979 1991
rect 999 1987 1000 1991
rect 1000 1987 1003 1991
rect 1095 1987 1099 1991
rect 1195 1987 1199 1991
rect 1215 1987 1219 1991
rect 1287 1988 1291 1992
rect 1327 1985 1331 1989
rect 1455 1988 1459 1992
rect 1511 1988 1515 1992
rect 1575 1988 1579 1992
rect 1639 1988 1643 1992
rect 1703 1988 1707 1992
rect 1767 1988 1771 1992
rect 1831 1988 1835 1992
rect 1895 1988 1899 1992
rect 1959 1988 1963 1992
rect 2031 1988 2035 1992
rect 2503 1985 2507 1989
rect 231 1967 232 1971
rect 232 1967 235 1971
rect 283 1967 284 1971
rect 284 1967 287 1971
rect 355 1967 356 1971
rect 356 1967 359 1971
rect 431 1967 435 1971
rect 531 1967 532 1971
rect 532 1967 535 1971
rect 627 1967 628 1971
rect 628 1967 631 1971
rect 727 1967 731 1971
rect 843 1967 844 1971
rect 844 1967 847 1971
rect 1115 1967 1119 1971
rect 1195 1967 1196 1971
rect 1196 1967 1199 1971
rect 1327 1968 1331 1972
rect 1471 1967 1475 1971
rect 1507 1967 1511 1971
rect 1527 1967 1531 1971
rect 1543 1967 1547 1971
rect 1591 1967 1595 1971
rect 1599 1967 1603 1971
rect 1655 1967 1659 1971
rect 1719 1967 1723 1971
rect 167 1951 171 1955
rect 175 1951 179 1955
rect 239 1951 243 1955
rect 419 1951 420 1955
rect 420 1951 423 1955
rect 463 1951 467 1955
rect 899 1951 900 1955
rect 900 1951 903 1955
rect 1055 1951 1059 1955
rect 1783 1967 1787 1971
rect 1827 1967 1831 1971
rect 1847 1967 1851 1971
rect 1891 1967 1895 1971
rect 1911 1967 1915 1971
rect 1955 1967 1959 1971
rect 1975 1967 1979 1971
rect 2027 1967 2031 1971
rect 2047 1967 2051 1971
rect 2055 1967 2059 1971
rect 2503 1968 2507 1972
rect 1507 1947 1508 1951
rect 1508 1947 1511 1951
rect 1711 1947 1715 1951
rect 1775 1947 1779 1951
rect 1827 1947 1828 1951
rect 1828 1947 1831 1951
rect 1891 1947 1892 1951
rect 1892 1947 1895 1951
rect 1955 1947 1956 1951
rect 1956 1947 1959 1951
rect 2027 1947 2028 1951
rect 2028 1947 2031 1951
rect 1599 1939 1603 1943
rect 2055 1939 2059 1943
rect 111 1932 115 1936
rect 151 1933 155 1937
rect 175 1931 176 1935
rect 176 1931 179 1935
rect 215 1933 219 1937
rect 239 1931 240 1935
rect 240 1931 243 1935
rect 319 1933 323 1937
rect 351 1931 355 1935
rect 439 1933 443 1937
rect 463 1931 464 1935
rect 464 1931 467 1935
rect 583 1933 587 1937
rect 603 1931 604 1935
rect 604 1931 607 1935
rect 743 1933 747 1937
rect 751 1931 755 1935
rect 919 1933 923 1937
rect 1095 1933 1099 1937
rect 1115 1931 1116 1935
rect 1116 1931 1119 1935
rect 1287 1932 1291 1936
rect 1599 1931 1603 1935
rect 1663 1931 1667 1935
rect 1767 1931 1771 1935
rect 1815 1931 1819 1935
rect 1943 1931 1947 1935
rect 2023 1931 2027 1935
rect 2111 1931 2115 1935
rect 2207 1931 2211 1935
rect 2399 1931 2403 1935
rect 2419 1923 2423 1927
rect 111 1915 115 1919
rect 135 1912 139 1916
rect 199 1912 203 1916
rect 303 1912 307 1916
rect 423 1912 427 1916
rect 567 1912 571 1916
rect 727 1912 731 1916
rect 903 1912 907 1916
rect 1079 1912 1083 1916
rect 1287 1915 1291 1919
rect 1327 1912 1331 1916
rect 1567 1913 1571 1917
rect 1599 1911 1603 1915
rect 1631 1913 1635 1917
rect 1663 1911 1667 1915
rect 1703 1913 1707 1917
rect 1711 1911 1715 1915
rect 1775 1913 1779 1917
rect 1815 1911 1819 1915
rect 1847 1913 1851 1917
rect 1919 1913 1923 1917
rect 1943 1911 1944 1915
rect 1944 1911 1947 1915
rect 1999 1913 2003 1917
rect 2023 1911 2024 1915
rect 2024 1911 2027 1915
rect 2087 1913 2091 1917
rect 2111 1911 2112 1915
rect 2112 1911 2115 1915
rect 2183 1913 2187 1917
rect 2207 1911 2208 1915
rect 2208 1911 2211 1915
rect 2279 1913 2283 1917
rect 2287 1911 2291 1915
rect 2375 1913 2379 1917
rect 2399 1911 2400 1915
rect 2400 1911 2403 1915
rect 2455 1913 2459 1917
rect 2471 1911 2475 1915
rect 2503 1912 2507 1916
rect 111 1889 115 1893
rect 135 1892 139 1896
rect 191 1892 195 1896
rect 271 1892 275 1896
rect 359 1892 363 1896
rect 455 1892 459 1896
rect 543 1892 547 1896
rect 631 1892 635 1896
rect 719 1892 723 1896
rect 799 1892 803 1896
rect 871 1892 875 1896
rect 943 1892 947 1896
rect 1015 1892 1019 1896
rect 1087 1892 1091 1896
rect 1159 1892 1163 1896
rect 1327 1895 1331 1899
rect 1287 1889 1291 1893
rect 1551 1892 1555 1896
rect 1615 1892 1619 1896
rect 1687 1892 1691 1896
rect 1759 1892 1763 1896
rect 1831 1892 1835 1896
rect 1903 1892 1907 1896
rect 1983 1892 1987 1896
rect 2071 1892 2075 1896
rect 2167 1892 2171 1896
rect 2263 1892 2267 1896
rect 2359 1892 2363 1896
rect 2439 1892 2443 1896
rect 2503 1895 2507 1899
rect 111 1872 115 1876
rect 151 1871 155 1875
rect 159 1871 163 1875
rect 207 1871 211 1875
rect 287 1871 291 1875
rect 375 1871 379 1875
rect 451 1871 455 1875
rect 471 1871 475 1875
rect 559 1871 563 1875
rect 575 1871 579 1875
rect 647 1871 651 1875
rect 735 1871 739 1875
rect 795 1871 799 1875
rect 815 1871 819 1875
rect 867 1871 871 1875
rect 887 1871 891 1875
rect 939 1871 943 1875
rect 959 1871 963 1875
rect 1023 1871 1027 1875
rect 1031 1871 1035 1875
rect 1055 1871 1056 1875
rect 1056 1871 1059 1875
rect 1103 1871 1107 1875
rect 1151 1871 1155 1875
rect 1175 1871 1179 1875
rect 751 1859 755 1863
rect 983 1863 987 1867
rect 1287 1872 1291 1876
rect 1327 1873 1331 1877
rect 1607 1876 1611 1880
rect 1663 1876 1667 1880
rect 1727 1876 1731 1880
rect 1799 1876 1803 1880
rect 1871 1876 1875 1880
rect 1943 1876 1947 1880
rect 2007 1876 2011 1880
rect 2071 1876 2075 1880
rect 2135 1876 2139 1880
rect 2199 1876 2203 1880
rect 2263 1876 2267 1880
rect 2327 1876 2331 1880
rect 2383 1876 2387 1880
rect 2439 1876 2443 1880
rect 2503 1873 2507 1877
rect 351 1851 355 1855
rect 451 1851 452 1855
rect 452 1851 455 1855
rect 1327 1856 1331 1860
rect 711 1851 715 1855
rect 787 1847 791 1851
rect 795 1851 796 1855
rect 796 1851 799 1855
rect 867 1851 868 1855
rect 868 1851 871 1855
rect 939 1851 940 1855
rect 940 1851 943 1855
rect 951 1851 955 1855
rect 1023 1851 1027 1855
rect 1623 1855 1627 1859
rect 1151 1851 1155 1855
rect 1659 1855 1663 1859
rect 1679 1855 1683 1859
rect 1723 1855 1727 1859
rect 1743 1855 1747 1859
rect 1767 1855 1768 1859
rect 1768 1855 1771 1859
rect 1815 1855 1819 1859
rect 1887 1855 1891 1859
rect 1895 1855 1899 1859
rect 1959 1855 1963 1859
rect 2023 1855 2027 1859
rect 2067 1855 2071 1859
rect 2087 1855 2091 1859
rect 2131 1855 2135 1859
rect 2151 1855 2155 1859
rect 2195 1855 2199 1859
rect 2215 1855 2219 1859
rect 2259 1855 2263 1859
rect 2279 1855 2283 1859
rect 2323 1855 2327 1859
rect 2343 1855 2347 1859
rect 2379 1855 2383 1859
rect 2399 1855 2403 1859
rect 2419 1855 2420 1859
rect 2420 1855 2423 1859
rect 2455 1855 2459 1859
rect 2463 1855 2467 1859
rect 2503 1856 2507 1860
rect 159 1839 163 1843
rect 175 1839 179 1843
rect 231 1839 235 1843
rect 411 1839 415 1843
rect 575 1839 576 1843
rect 576 1839 579 1843
rect 831 1839 835 1843
rect 919 1839 923 1843
rect 983 1839 984 1843
rect 984 1839 987 1843
rect 1023 1839 1027 1843
rect 1111 1839 1115 1843
rect 2287 1843 2291 1847
rect 1659 1835 1660 1839
rect 1660 1835 1663 1839
rect 1723 1835 1724 1839
rect 1724 1835 1727 1839
rect 1895 1831 1899 1835
rect 1971 1835 1975 1839
rect 2067 1835 2068 1839
rect 2068 1835 2071 1839
rect 2131 1835 2132 1839
rect 2132 1835 2135 1839
rect 2195 1835 2196 1839
rect 2196 1835 2199 1839
rect 2259 1835 2260 1839
rect 2260 1835 2263 1839
rect 2323 1835 2324 1839
rect 2324 1835 2327 1839
rect 2379 1835 2380 1839
rect 2380 1835 2383 1839
rect 2471 1835 2475 1839
rect 111 1820 115 1824
rect 151 1821 155 1825
rect 175 1819 176 1823
rect 176 1819 179 1823
rect 207 1821 211 1825
rect 231 1819 232 1823
rect 232 1819 235 1823
rect 295 1821 299 1825
rect 391 1821 395 1825
rect 411 1819 412 1823
rect 412 1819 415 1823
rect 495 1821 499 1825
rect 511 1819 515 1823
rect 591 1821 595 1825
rect 615 1819 616 1823
rect 616 1819 619 1823
rect 687 1821 691 1825
rect 711 1819 712 1823
rect 712 1819 715 1823
rect 775 1821 779 1825
rect 787 1819 791 1823
rect 855 1821 859 1825
rect 927 1821 931 1825
rect 951 1819 952 1823
rect 952 1819 955 1823
rect 999 1821 1003 1825
rect 1023 1819 1024 1823
rect 1024 1819 1027 1823
rect 1079 1821 1083 1825
rect 1111 1819 1115 1823
rect 1159 1821 1163 1825
rect 1175 1819 1179 1823
rect 1287 1820 1291 1824
rect 1655 1819 1659 1823
rect 1663 1819 1667 1823
rect 1751 1819 1755 1823
rect 111 1803 115 1807
rect 135 1800 139 1804
rect 191 1800 195 1804
rect 279 1800 283 1804
rect 375 1800 379 1804
rect 479 1800 483 1804
rect 575 1800 579 1804
rect 671 1800 675 1804
rect 759 1800 763 1804
rect 839 1800 843 1804
rect 911 1800 915 1804
rect 983 1800 987 1804
rect 1063 1800 1067 1804
rect 1143 1800 1147 1804
rect 1287 1803 1291 1807
rect 1971 1807 1975 1811
rect 2327 1819 2331 1823
rect 2463 1819 2467 1823
rect 1327 1800 1331 1804
rect 1631 1801 1635 1805
rect 1663 1799 1667 1803
rect 1719 1801 1723 1805
rect 1751 1799 1755 1803
rect 1815 1801 1819 1805
rect 1927 1801 1931 1805
rect 2055 1801 2059 1805
rect 2191 1801 2195 1805
rect 2207 1799 2211 1803
rect 2335 1801 2339 1805
rect 2455 1801 2459 1805
rect 2471 1799 2475 1803
rect 2503 1800 2507 1804
rect 1327 1783 1331 1787
rect 111 1773 115 1777
rect 135 1776 139 1780
rect 199 1776 203 1780
rect 295 1776 299 1780
rect 399 1776 403 1780
rect 503 1776 507 1780
rect 607 1776 611 1780
rect 703 1776 707 1780
rect 799 1776 803 1780
rect 887 1776 891 1780
rect 975 1776 979 1780
rect 1063 1776 1067 1780
rect 1151 1776 1155 1780
rect 1615 1780 1619 1784
rect 1703 1780 1707 1784
rect 1799 1780 1803 1784
rect 1911 1780 1915 1784
rect 2039 1780 2043 1784
rect 2175 1780 2179 1784
rect 2319 1780 2323 1784
rect 2439 1780 2443 1784
rect 2503 1783 2507 1787
rect 1287 1773 1291 1777
rect 1327 1765 1331 1769
rect 1527 1768 1531 1772
rect 1607 1768 1611 1772
rect 1695 1768 1699 1772
rect 1791 1768 1795 1772
rect 1879 1768 1883 1772
rect 1967 1768 1971 1772
rect 2055 1768 2059 1772
rect 2135 1768 2139 1772
rect 2215 1768 2219 1772
rect 2295 1768 2299 1772
rect 2375 1768 2379 1772
rect 2439 1768 2443 1772
rect 2503 1765 2507 1769
rect 111 1756 115 1760
rect 151 1755 155 1759
rect 195 1755 199 1759
rect 215 1755 219 1759
rect 291 1755 295 1759
rect 311 1755 315 1759
rect 395 1755 399 1759
rect 415 1755 419 1759
rect 423 1755 427 1759
rect 519 1755 523 1759
rect 587 1755 591 1759
rect 623 1755 627 1759
rect 719 1755 723 1759
rect 795 1755 799 1759
rect 815 1755 819 1759
rect 831 1755 835 1759
rect 903 1755 907 1759
rect 919 1755 923 1759
rect 991 1755 995 1759
rect 1027 1755 1031 1759
rect 1079 1755 1083 1759
rect 1167 1755 1171 1759
rect 1287 1756 1291 1760
rect 1327 1748 1331 1752
rect 1543 1747 1547 1751
rect 1603 1747 1607 1751
rect 1623 1747 1627 1751
rect 1691 1747 1695 1751
rect 1711 1747 1715 1751
rect 1787 1747 1791 1751
rect 1807 1747 1811 1751
rect 1875 1747 1879 1751
rect 1895 1747 1899 1751
rect 1915 1747 1916 1751
rect 1916 1747 1919 1751
rect 1983 1747 1987 1751
rect 2051 1747 2055 1751
rect 2071 1747 2075 1751
rect 2091 1747 2092 1751
rect 2092 1747 2095 1751
rect 2151 1747 2155 1751
rect 2231 1747 2235 1751
rect 135 1735 136 1739
rect 136 1735 139 1739
rect 195 1735 196 1739
rect 196 1735 199 1739
rect 291 1735 292 1739
rect 292 1735 295 1739
rect 395 1735 396 1739
rect 396 1735 399 1739
rect 615 1735 619 1739
rect 731 1735 735 1739
rect 795 1735 796 1739
rect 796 1735 799 1739
rect 955 1735 959 1739
rect 1175 1735 1179 1739
rect 2311 1747 2315 1751
rect 2327 1747 2331 1751
rect 2391 1747 2395 1751
rect 2455 1747 2459 1751
rect 2463 1747 2467 1751
rect 2503 1748 2507 1752
rect 423 1727 427 1731
rect 1595 1727 1599 1731
rect 1603 1727 1604 1731
rect 1604 1727 1607 1731
rect 1691 1727 1692 1731
rect 1692 1727 1695 1731
rect 1787 1727 1788 1731
rect 1788 1727 1791 1731
rect 1875 1727 1876 1731
rect 1876 1727 1879 1731
rect 2051 1727 2052 1731
rect 2052 1727 2055 1731
rect 2207 1727 2211 1731
rect 2403 1727 2407 1731
rect 2471 1727 2475 1731
rect 191 1719 195 1723
rect 263 1719 267 1723
rect 343 1719 347 1723
rect 431 1719 435 1723
rect 587 1719 588 1723
rect 588 1719 591 1723
rect 799 1719 803 1723
rect 911 1719 915 1723
rect 1027 1719 1028 1723
rect 1028 1719 1031 1723
rect 1071 1719 1075 1723
rect 1415 1711 1419 1715
rect 1423 1711 1427 1715
rect 1487 1711 1491 1715
rect 1567 1711 1571 1715
rect 1655 1711 1659 1715
rect 1751 1711 1755 1715
rect 111 1700 115 1704
rect 167 1701 171 1705
rect 191 1699 192 1703
rect 192 1699 195 1703
rect 239 1701 243 1705
rect 263 1699 264 1703
rect 264 1699 267 1703
rect 319 1701 323 1705
rect 343 1699 344 1703
rect 344 1699 347 1703
rect 407 1701 411 1705
rect 431 1699 432 1703
rect 432 1699 435 1703
rect 503 1701 507 1705
rect 511 1699 515 1703
rect 607 1701 611 1705
rect 615 1699 619 1703
rect 711 1701 715 1705
rect 731 1699 732 1703
rect 732 1699 735 1703
rect 823 1701 827 1705
rect 935 1701 939 1705
rect 955 1699 956 1703
rect 956 1699 959 1703
rect 1047 1701 1051 1705
rect 1071 1699 1072 1703
rect 1072 1699 1075 1703
rect 1159 1701 1163 1705
rect 1175 1699 1179 1703
rect 1287 1700 1291 1704
rect 1943 1711 1947 1715
rect 2091 1711 2092 1715
rect 2092 1711 2095 1715
rect 2135 1711 2139 1715
rect 2319 1711 2323 1715
rect 2463 1711 2467 1715
rect 2475 1703 2479 1707
rect 1327 1692 1331 1696
rect 1399 1693 1403 1697
rect 1423 1691 1424 1695
rect 1424 1691 1427 1695
rect 1463 1693 1467 1697
rect 1487 1691 1488 1695
rect 1488 1691 1491 1695
rect 1543 1693 1547 1697
rect 1567 1691 1568 1695
rect 1568 1691 1571 1695
rect 1631 1693 1635 1697
rect 1655 1691 1656 1695
rect 1656 1691 1659 1695
rect 1727 1693 1731 1697
rect 1751 1691 1752 1695
rect 1752 1691 1755 1695
rect 1823 1693 1827 1697
rect 1843 1691 1844 1695
rect 1844 1691 1847 1695
rect 1919 1693 1923 1697
rect 1943 1691 1944 1695
rect 1944 1691 1947 1695
rect 2015 1693 2019 1697
rect 2031 1691 2035 1695
rect 2111 1693 2115 1697
rect 2135 1691 2136 1695
rect 2136 1691 2139 1695
rect 2199 1693 2203 1697
rect 2287 1693 2291 1697
rect 2319 1691 2323 1695
rect 2383 1693 2387 1697
rect 2403 1691 2404 1695
rect 2404 1691 2407 1695
rect 2455 1693 2459 1697
rect 2463 1691 2467 1695
rect 2503 1692 2507 1696
rect 111 1683 115 1687
rect 151 1680 155 1684
rect 223 1680 227 1684
rect 303 1680 307 1684
rect 391 1680 395 1684
rect 487 1680 491 1684
rect 591 1680 595 1684
rect 695 1680 699 1684
rect 807 1680 811 1684
rect 919 1680 923 1684
rect 1031 1680 1035 1684
rect 1143 1680 1147 1684
rect 1287 1683 1291 1687
rect 1327 1675 1331 1679
rect 1383 1672 1387 1676
rect 1447 1672 1451 1676
rect 1527 1672 1531 1676
rect 1615 1672 1619 1676
rect 1711 1672 1715 1676
rect 1807 1672 1811 1676
rect 1903 1672 1907 1676
rect 1999 1672 2003 1676
rect 2095 1672 2099 1676
rect 2183 1672 2187 1676
rect 2271 1672 2275 1676
rect 2367 1672 2371 1676
rect 2439 1672 2443 1676
rect 2503 1675 2507 1679
rect 111 1661 115 1665
rect 255 1664 259 1668
rect 319 1664 323 1668
rect 399 1664 403 1668
rect 487 1664 491 1668
rect 575 1664 579 1668
rect 671 1664 675 1668
rect 767 1664 771 1668
rect 863 1664 867 1668
rect 959 1664 963 1668
rect 1063 1664 1067 1668
rect 1167 1664 1171 1668
rect 1287 1661 1291 1665
rect 1327 1653 1331 1657
rect 1351 1656 1355 1660
rect 1407 1656 1411 1660
rect 1495 1656 1499 1660
rect 1583 1656 1587 1660
rect 1679 1656 1683 1660
rect 1783 1656 1787 1660
rect 1895 1656 1899 1660
rect 2023 1656 2027 1660
rect 2159 1656 2163 1660
rect 2303 1656 2307 1660
rect 2439 1656 2443 1660
rect 2503 1653 2507 1657
rect 111 1644 115 1648
rect 271 1643 275 1647
rect 315 1643 319 1647
rect 335 1643 339 1647
rect 395 1643 399 1647
rect 415 1643 419 1647
rect 483 1643 487 1647
rect 503 1643 507 1647
rect 519 1643 523 1647
rect 591 1643 595 1647
rect 607 1643 611 1647
rect 687 1643 691 1647
rect 763 1643 767 1647
rect 783 1643 787 1647
rect 799 1643 803 1647
rect 879 1643 883 1647
rect 911 1643 915 1647
rect 975 1643 979 1647
rect 1059 1643 1063 1647
rect 1079 1643 1083 1647
rect 1099 1643 1100 1647
rect 1100 1643 1103 1647
rect 1183 1643 1187 1647
rect 511 1631 515 1635
rect 1287 1644 1291 1648
rect 1327 1636 1331 1640
rect 1367 1635 1371 1639
rect 1403 1635 1407 1639
rect 1423 1635 1427 1639
rect 1491 1635 1495 1639
rect 1511 1635 1515 1639
rect 1579 1635 1583 1639
rect 1599 1635 1603 1639
rect 1675 1635 1679 1639
rect 1695 1635 1699 1639
rect 1703 1635 1707 1639
rect 1799 1635 1803 1639
rect 1891 1635 1895 1639
rect 1911 1635 1915 1639
rect 1931 1635 1932 1639
rect 1932 1635 1935 1639
rect 2039 1635 2043 1639
rect 2155 1635 2159 1639
rect 2175 1635 2179 1639
rect 2299 1635 2303 1639
rect 2319 1635 2323 1639
rect 2455 1635 2459 1639
rect 2475 1635 2476 1639
rect 2476 1635 2479 1639
rect 2503 1636 2507 1640
rect 315 1623 316 1627
rect 316 1623 319 1627
rect 395 1623 396 1627
rect 396 1623 399 1627
rect 483 1623 484 1627
rect 484 1623 487 1627
rect 615 1623 619 1627
rect 755 1623 759 1627
rect 763 1623 764 1627
rect 764 1623 767 1627
rect 915 1623 919 1627
rect 1059 1623 1060 1627
rect 1060 1623 1063 1627
rect 1175 1623 1179 1627
rect 519 1615 523 1619
rect 1403 1615 1404 1619
rect 1404 1615 1407 1619
rect 1491 1615 1492 1619
rect 1492 1615 1495 1619
rect 1579 1615 1580 1619
rect 1580 1615 1583 1619
rect 1675 1615 1676 1619
rect 1676 1615 1679 1619
rect 1891 1615 1892 1619
rect 1892 1615 1895 1619
rect 2031 1619 2035 1623
rect 2155 1615 2156 1619
rect 2156 1615 2159 1619
rect 2299 1615 2300 1619
rect 2300 1615 2303 1619
rect 2463 1615 2467 1619
rect 327 1607 331 1611
rect 383 1607 387 1611
rect 607 1607 611 1611
rect 707 1607 711 1611
rect 719 1607 723 1611
rect 799 1607 803 1611
rect 255 1595 259 1599
rect 111 1588 115 1592
rect 303 1589 307 1593
rect 327 1587 328 1591
rect 328 1587 331 1591
rect 359 1589 363 1593
rect 383 1587 384 1591
rect 384 1587 387 1591
rect 431 1589 435 1593
rect 479 1587 483 1591
rect 755 1595 759 1599
rect 1099 1607 1100 1611
rect 1100 1607 1103 1611
rect 1263 1603 1267 1607
rect 1391 1603 1395 1607
rect 1447 1603 1451 1607
rect 1503 1603 1507 1607
rect 1583 1603 1587 1607
rect 503 1587 507 1591
rect 511 1589 515 1593
rect 519 1587 523 1591
rect 599 1589 603 1593
rect 695 1589 699 1593
rect 719 1587 720 1591
rect 720 1587 723 1591
rect 791 1589 795 1593
rect 895 1589 899 1593
rect 915 1587 916 1591
rect 916 1587 919 1591
rect 1007 1589 1011 1593
rect 1015 1587 1019 1591
rect 1119 1589 1123 1593
rect 1287 1588 1291 1592
rect 1931 1603 1932 1607
rect 1932 1603 1935 1607
rect 1975 1603 1979 1607
rect 1327 1584 1331 1588
rect 1367 1585 1371 1589
rect 1391 1583 1392 1587
rect 1392 1583 1395 1587
rect 1423 1585 1427 1589
rect 1447 1583 1448 1587
rect 1448 1583 1451 1587
rect 1479 1585 1483 1589
rect 1503 1583 1504 1587
rect 1504 1583 1507 1587
rect 1559 1585 1563 1589
rect 1583 1583 1584 1587
rect 1584 1583 1587 1587
rect 1639 1585 1643 1589
rect 1719 1585 1723 1589
rect 1743 1583 1744 1587
rect 1744 1583 1747 1587
rect 1791 1585 1795 1589
rect 1871 1585 1875 1589
rect 1951 1585 1955 1589
rect 1975 1583 1976 1587
rect 1976 1583 1979 1587
rect 2031 1585 2035 1589
rect 2503 1584 2507 1588
rect 111 1571 115 1575
rect 287 1568 291 1572
rect 343 1568 347 1572
rect 415 1568 419 1572
rect 495 1568 499 1572
rect 583 1568 587 1572
rect 679 1568 683 1572
rect 775 1568 779 1572
rect 879 1568 883 1572
rect 991 1568 995 1572
rect 1103 1568 1107 1572
rect 1287 1571 1291 1575
rect 1327 1567 1331 1571
rect 1351 1564 1355 1568
rect 1407 1564 1411 1568
rect 1463 1564 1467 1568
rect 1543 1564 1547 1568
rect 1623 1564 1627 1568
rect 1703 1564 1707 1568
rect 1775 1564 1779 1568
rect 1855 1564 1859 1568
rect 1935 1564 1939 1568
rect 2015 1564 2019 1568
rect 2503 1567 2507 1571
rect 111 1553 115 1557
rect 247 1556 251 1560
rect 319 1556 323 1560
rect 399 1556 403 1560
rect 487 1556 491 1560
rect 583 1556 587 1560
rect 671 1556 675 1560
rect 759 1556 763 1560
rect 847 1556 851 1560
rect 927 1556 931 1560
rect 1007 1556 1011 1560
rect 1087 1556 1091 1560
rect 1167 1556 1171 1560
rect 1223 1556 1227 1560
rect 1287 1553 1291 1557
rect 1327 1549 1331 1553
rect 1351 1552 1355 1556
rect 1471 1552 1475 1556
rect 1607 1552 1611 1556
rect 1735 1552 1739 1556
rect 1871 1552 1875 1556
rect 2007 1552 2011 1556
rect 2503 1549 2507 1553
rect 111 1536 115 1540
rect 263 1535 267 1539
rect 271 1535 275 1539
rect 335 1535 339 1539
rect 351 1535 355 1539
rect 415 1535 419 1539
rect 503 1535 507 1539
rect 579 1535 583 1539
rect 599 1535 603 1539
rect 687 1535 691 1539
rect 707 1535 708 1539
rect 708 1535 711 1539
rect 775 1535 779 1539
rect 799 1535 800 1539
rect 800 1535 803 1539
rect 863 1535 867 1539
rect 879 1535 883 1539
rect 943 1535 947 1539
rect 1023 1535 1027 1539
rect 1103 1535 1107 1539
rect 1163 1535 1167 1539
rect 1183 1535 1187 1539
rect 1219 1535 1223 1539
rect 1239 1535 1243 1539
rect 1263 1535 1264 1539
rect 1264 1535 1267 1539
rect 1287 1536 1291 1540
rect 1327 1532 1331 1536
rect 1367 1531 1371 1535
rect 1487 1531 1491 1535
rect 1603 1531 1607 1535
rect 1623 1531 1627 1535
rect 1731 1531 1735 1535
rect 1751 1531 1755 1535
rect 1863 1531 1867 1535
rect 1887 1531 1891 1535
rect 2003 1531 2007 1535
rect 2023 1531 2027 1535
rect 255 1515 259 1519
rect 479 1515 483 1519
rect 579 1515 580 1519
rect 580 1515 583 1519
rect 671 1515 672 1519
rect 672 1515 675 1519
rect 755 1515 756 1519
rect 756 1515 759 1519
rect 1015 1515 1019 1519
rect 1163 1515 1164 1519
rect 1164 1515 1167 1519
rect 1219 1515 1220 1519
rect 1220 1515 1223 1519
rect 1743 1519 1747 1523
rect 1775 1523 1779 1527
rect 2503 1532 2507 1536
rect 1387 1511 1391 1515
rect 1603 1511 1604 1515
rect 1604 1511 1607 1515
rect 1731 1511 1732 1515
rect 1732 1511 1735 1515
rect 1863 1511 1867 1515
rect 2003 1511 2004 1515
rect 2004 1511 2007 1515
rect 271 1495 275 1499
rect 351 1495 355 1499
rect 367 1495 371 1499
rect 439 1495 443 1499
rect 607 1495 611 1499
rect 851 1495 855 1499
rect 879 1495 880 1499
rect 880 1495 883 1499
rect 935 1495 939 1499
rect 999 1495 1003 1499
rect 1079 1495 1083 1499
rect 631 1487 635 1491
rect 1567 1499 1571 1503
rect 1575 1499 1579 1503
rect 1655 1499 1659 1503
rect 1775 1499 1776 1503
rect 1776 1499 1779 1503
rect 1815 1499 1819 1503
rect 1895 1499 1899 1503
rect 1975 1499 1979 1503
rect 2055 1499 2059 1503
rect 1823 1487 1827 1491
rect 111 1476 115 1480
rect 279 1477 283 1481
rect 287 1475 291 1479
rect 343 1477 347 1481
rect 367 1475 368 1479
rect 368 1475 371 1479
rect 415 1477 419 1481
rect 439 1475 440 1479
rect 440 1475 443 1479
rect 495 1477 499 1481
rect 511 1475 515 1479
rect 575 1477 579 1481
rect 607 1475 611 1479
rect 655 1477 659 1481
rect 671 1475 675 1479
rect 735 1477 739 1481
rect 755 1475 756 1479
rect 756 1475 759 1479
rect 815 1477 819 1481
rect 895 1477 899 1481
rect 935 1475 939 1479
rect 975 1477 979 1481
rect 999 1475 1000 1479
rect 1000 1475 1003 1479
rect 1055 1477 1059 1481
rect 1079 1475 1080 1479
rect 1080 1475 1083 1479
rect 1143 1477 1147 1481
rect 1151 1475 1155 1479
rect 1287 1476 1291 1480
rect 1327 1480 1331 1484
rect 1367 1481 1371 1485
rect 1387 1479 1388 1483
rect 1388 1479 1391 1483
rect 1423 1481 1427 1485
rect 1479 1481 1483 1485
rect 1551 1481 1555 1485
rect 1575 1479 1576 1483
rect 1576 1479 1579 1483
rect 1631 1481 1635 1485
rect 1655 1479 1656 1483
rect 1656 1479 1659 1483
rect 1711 1481 1715 1485
rect 1791 1481 1795 1485
rect 1815 1479 1816 1483
rect 1816 1479 1819 1483
rect 1871 1481 1875 1485
rect 1895 1479 1896 1483
rect 1896 1479 1899 1483
rect 1951 1481 1955 1485
rect 1975 1479 1976 1483
rect 1976 1479 1979 1483
rect 2031 1481 2035 1485
rect 2055 1479 2056 1483
rect 2056 1479 2059 1483
rect 2119 1481 2123 1485
rect 2503 1480 2507 1484
rect 111 1459 115 1463
rect 263 1456 267 1460
rect 327 1456 331 1460
rect 399 1456 403 1460
rect 479 1456 483 1460
rect 559 1456 563 1460
rect 639 1456 643 1460
rect 719 1456 723 1460
rect 799 1456 803 1460
rect 879 1456 883 1460
rect 959 1456 963 1460
rect 1039 1456 1043 1460
rect 1127 1456 1131 1460
rect 1287 1459 1291 1463
rect 1327 1463 1331 1467
rect 1351 1460 1355 1464
rect 1407 1460 1411 1464
rect 1463 1460 1467 1464
rect 1535 1460 1539 1464
rect 1615 1460 1619 1464
rect 1695 1460 1699 1464
rect 1775 1460 1779 1464
rect 1855 1460 1859 1464
rect 1935 1460 1939 1464
rect 2015 1460 2019 1464
rect 2103 1460 2107 1464
rect 2503 1463 2507 1467
rect 111 1437 115 1441
rect 191 1440 195 1444
rect 255 1440 259 1444
rect 327 1440 331 1444
rect 407 1440 411 1444
rect 503 1440 507 1444
rect 607 1440 611 1444
rect 711 1440 715 1444
rect 815 1440 819 1444
rect 919 1440 923 1444
rect 1023 1440 1027 1444
rect 1127 1440 1131 1444
rect 1223 1440 1227 1444
rect 1287 1437 1291 1441
rect 1327 1437 1331 1441
rect 1359 1440 1363 1444
rect 1447 1440 1451 1444
rect 1535 1440 1539 1444
rect 1631 1440 1635 1444
rect 1727 1440 1731 1444
rect 1815 1440 1819 1444
rect 1903 1440 1907 1444
rect 1991 1440 1995 1444
rect 2071 1440 2075 1444
rect 2159 1440 2163 1444
rect 2247 1440 2251 1444
rect 2503 1437 2507 1441
rect 111 1420 115 1424
rect 207 1419 211 1423
rect 215 1419 219 1423
rect 271 1419 275 1423
rect 343 1419 347 1423
rect 351 1419 355 1423
rect 423 1419 427 1423
rect 519 1419 523 1423
rect 623 1419 627 1423
rect 631 1419 635 1423
rect 727 1419 731 1423
rect 831 1419 835 1423
rect 851 1419 852 1423
rect 852 1419 855 1423
rect 935 1419 939 1423
rect 1019 1419 1023 1423
rect 1039 1419 1043 1423
rect 1123 1419 1127 1423
rect 1143 1419 1147 1423
rect 1219 1419 1223 1423
rect 1239 1419 1243 1423
rect 1247 1419 1251 1423
rect 1287 1420 1291 1424
rect 1327 1420 1331 1424
rect 1375 1419 1379 1423
rect 1443 1419 1447 1423
rect 1463 1419 1467 1423
rect 1531 1419 1535 1423
rect 1551 1419 1555 1423
rect 1567 1419 1571 1423
rect 1647 1419 1651 1423
rect 1743 1419 1747 1423
rect 1151 1407 1155 1411
rect 1831 1419 1835 1423
rect 1899 1419 1903 1423
rect 1919 1419 1923 1423
rect 1987 1419 1991 1423
rect 2007 1419 2011 1423
rect 2067 1419 2071 1423
rect 2087 1419 2091 1423
rect 2155 1419 2159 1423
rect 2175 1419 2179 1423
rect 2239 1419 2243 1423
rect 2263 1419 2267 1423
rect 2503 1420 2507 1424
rect 1995 1411 1999 1415
rect 287 1399 291 1403
rect 511 1399 515 1403
rect 687 1399 691 1403
rect 859 1399 863 1403
rect 1019 1399 1020 1403
rect 1020 1399 1023 1403
rect 1123 1399 1124 1403
rect 1124 1399 1127 1403
rect 1219 1399 1220 1403
rect 1220 1399 1223 1403
rect 1443 1399 1444 1403
rect 1444 1399 1447 1403
rect 1531 1399 1532 1403
rect 1532 1399 1535 1403
rect 1755 1399 1759 1403
rect 1823 1399 1827 1403
rect 1899 1399 1900 1403
rect 1900 1399 1903 1403
rect 1987 1399 1988 1403
rect 1988 1399 1991 1403
rect 2067 1399 2068 1403
rect 2068 1399 2071 1403
rect 2155 1399 2156 1403
rect 2156 1399 2159 1403
rect 2239 1399 2243 1403
rect 215 1391 219 1395
rect 351 1391 355 1395
rect 175 1383 179 1387
rect 383 1383 387 1387
rect 463 1383 467 1387
rect 527 1383 531 1387
rect 607 1383 611 1387
rect 655 1383 659 1387
rect 775 1383 779 1387
rect 1247 1383 1251 1387
rect 1591 1387 1595 1391
rect 1671 1387 1675 1391
rect 1931 1387 1935 1391
rect 1991 1387 1992 1391
rect 1992 1387 1995 1391
rect 2031 1387 2035 1391
rect 2119 1387 2123 1391
rect 2215 1387 2219 1391
rect 2271 1387 2275 1391
rect 2415 1387 2419 1391
rect 2423 1387 2427 1391
rect 111 1364 115 1368
rect 151 1365 155 1369
rect 175 1363 176 1367
rect 176 1363 179 1367
rect 223 1365 227 1369
rect 247 1363 248 1367
rect 248 1363 251 1367
rect 295 1365 299 1369
rect 359 1365 363 1369
rect 383 1363 384 1367
rect 384 1363 387 1367
rect 431 1365 435 1369
rect 463 1363 467 1367
rect 503 1365 507 1369
rect 527 1363 528 1367
rect 528 1363 531 1367
rect 583 1365 587 1369
rect 607 1363 608 1367
rect 608 1363 611 1367
rect 663 1365 667 1369
rect 687 1363 688 1367
rect 688 1363 691 1367
rect 751 1365 755 1369
rect 775 1363 776 1367
rect 776 1363 779 1367
rect 839 1365 843 1369
rect 859 1363 860 1367
rect 860 1363 863 1367
rect 927 1365 931 1369
rect 967 1363 971 1367
rect 1015 1365 1019 1369
rect 1103 1365 1107 1369
rect 1199 1365 1203 1369
rect 1287 1364 1291 1368
rect 1327 1368 1331 1372
rect 1567 1369 1571 1373
rect 1591 1367 1592 1371
rect 1592 1367 1595 1371
rect 1647 1369 1651 1373
rect 1671 1367 1672 1371
rect 1672 1367 1675 1371
rect 1735 1369 1739 1373
rect 1755 1367 1756 1371
rect 1756 1367 1759 1371
rect 1831 1369 1835 1373
rect 1919 1369 1923 1373
rect 2007 1369 2011 1373
rect 2031 1367 2032 1371
rect 2032 1367 2035 1371
rect 2095 1369 2099 1373
rect 2119 1367 2120 1371
rect 2120 1367 2123 1371
rect 2175 1369 2179 1373
rect 2215 1367 2219 1371
rect 2247 1369 2251 1373
rect 2271 1367 2272 1371
rect 2272 1367 2275 1371
rect 2319 1369 2323 1373
rect 2327 1367 2331 1371
rect 2399 1369 2403 1373
rect 2423 1367 2424 1371
rect 2424 1367 2427 1371
rect 2455 1369 2459 1373
rect 2463 1367 2467 1371
rect 2503 1368 2507 1372
rect 111 1347 115 1351
rect 135 1344 139 1348
rect 207 1344 211 1348
rect 279 1344 283 1348
rect 343 1344 347 1348
rect 415 1344 419 1348
rect 487 1344 491 1348
rect 567 1344 571 1348
rect 647 1344 651 1348
rect 735 1344 739 1348
rect 823 1344 827 1348
rect 911 1344 915 1348
rect 999 1344 1003 1348
rect 1087 1344 1091 1348
rect 1183 1344 1187 1348
rect 1287 1347 1291 1351
rect 1327 1351 1331 1355
rect 1551 1348 1555 1352
rect 1631 1348 1635 1352
rect 1719 1348 1723 1352
rect 1815 1348 1819 1352
rect 1903 1348 1907 1352
rect 1991 1348 1995 1352
rect 2079 1348 2083 1352
rect 2159 1348 2163 1352
rect 2231 1348 2235 1352
rect 2303 1348 2307 1352
rect 2383 1348 2387 1352
rect 2439 1348 2443 1352
rect 2503 1351 2507 1355
rect 1327 1333 1331 1337
rect 1583 1336 1587 1340
rect 1647 1336 1651 1340
rect 1727 1336 1731 1340
rect 1807 1336 1811 1340
rect 1895 1336 1899 1340
rect 1983 1336 1987 1340
rect 2063 1336 2067 1340
rect 2143 1336 2147 1340
rect 2223 1336 2227 1340
rect 2303 1336 2307 1340
rect 2383 1336 2387 1340
rect 2439 1336 2443 1340
rect 2503 1333 2507 1337
rect 111 1313 115 1317
rect 135 1316 139 1320
rect 239 1316 243 1320
rect 367 1316 371 1320
rect 479 1316 483 1320
rect 583 1316 587 1320
rect 687 1316 691 1320
rect 783 1316 787 1320
rect 879 1316 883 1320
rect 975 1316 979 1320
rect 1287 1313 1291 1317
rect 1327 1316 1331 1320
rect 1599 1315 1603 1319
rect 1643 1315 1647 1319
rect 1663 1315 1667 1319
rect 1723 1315 1727 1319
rect 1743 1315 1747 1319
rect 1779 1315 1783 1319
rect 1823 1315 1827 1319
rect 1887 1315 1891 1319
rect 1911 1315 1915 1319
rect 1931 1315 1932 1319
rect 1932 1315 1935 1319
rect 1999 1315 2003 1319
rect 2079 1315 2083 1319
rect 2139 1315 2143 1319
rect 2159 1315 2163 1319
rect 2219 1315 2223 1319
rect 2239 1315 2243 1319
rect 2299 1315 2303 1319
rect 2319 1315 2323 1319
rect 2399 1315 2403 1319
rect 2415 1315 2419 1319
rect 2455 1315 2459 1319
rect 2471 1315 2475 1319
rect 2503 1316 2507 1320
rect 111 1296 115 1300
rect 151 1295 155 1299
rect 159 1295 163 1299
rect 255 1295 259 1299
rect 363 1295 367 1299
rect 383 1295 387 1299
rect 495 1295 499 1299
rect 579 1295 583 1299
rect 599 1295 603 1299
rect 655 1295 659 1299
rect 703 1295 707 1299
rect 747 1295 751 1299
rect 799 1295 803 1299
rect 807 1295 811 1299
rect 895 1295 899 1299
rect 991 1295 995 1299
rect 1287 1296 1291 1300
rect 1583 1295 1584 1299
rect 1584 1295 1587 1299
rect 1643 1295 1644 1299
rect 1644 1295 1647 1299
rect 1723 1295 1724 1299
rect 1724 1295 1727 1299
rect 1887 1295 1891 1299
rect 2011 1295 2015 1299
rect 2139 1295 2140 1299
rect 2140 1295 2143 1299
rect 2219 1295 2220 1299
rect 2220 1295 2223 1299
rect 2327 1295 2331 1299
rect 2391 1295 2395 1299
rect 2463 1295 2467 1299
rect 247 1275 251 1279
rect 363 1275 364 1279
rect 364 1275 367 1279
rect 571 1275 575 1279
rect 579 1275 580 1279
rect 580 1275 583 1279
rect 807 1271 811 1275
rect 967 1275 971 1279
rect 1607 1283 1611 1287
rect 1779 1283 1780 1287
rect 1780 1283 1783 1287
rect 1831 1283 1835 1287
rect 2067 1283 2071 1287
rect 2299 1283 2300 1287
rect 2300 1283 2303 1287
rect 1327 1264 1331 1268
rect 1567 1265 1571 1269
rect 1583 1263 1587 1267
rect 1631 1265 1635 1269
rect 1711 1265 1715 1269
rect 1719 1263 1723 1267
rect 1799 1265 1803 1269
rect 1831 1263 1835 1267
rect 1895 1265 1899 1269
rect 1991 1265 1995 1269
rect 2011 1263 2012 1267
rect 2012 1263 2015 1267
rect 2095 1265 2099 1269
rect 2111 1263 2115 1267
rect 2207 1265 2211 1269
rect 2319 1265 2323 1269
rect 2503 1264 2507 1268
rect 159 1255 163 1259
rect 239 1255 243 1259
rect 327 1255 331 1259
rect 463 1255 467 1259
rect 503 1255 507 1259
rect 747 1255 748 1259
rect 748 1255 751 1259
rect 791 1255 795 1259
rect 863 1255 867 1259
rect 1327 1247 1331 1251
rect 1551 1244 1555 1248
rect 1615 1244 1619 1248
rect 1695 1244 1699 1248
rect 1783 1244 1787 1248
rect 1879 1244 1883 1248
rect 1975 1244 1979 1248
rect 2079 1244 2083 1248
rect 2191 1244 2195 1248
rect 2303 1244 2307 1248
rect 2503 1247 2507 1251
rect 111 1236 115 1240
rect 151 1237 155 1241
rect 215 1237 219 1241
rect 239 1235 240 1239
rect 240 1235 243 1239
rect 303 1237 307 1241
rect 327 1235 328 1239
rect 328 1235 331 1239
rect 391 1237 395 1241
rect 399 1235 403 1239
rect 471 1237 475 1241
rect 503 1235 507 1239
rect 551 1237 555 1241
rect 571 1235 572 1239
rect 572 1235 575 1239
rect 623 1237 627 1241
rect 631 1235 635 1239
rect 695 1237 699 1241
rect 767 1237 771 1241
rect 791 1235 792 1239
rect 792 1235 795 1239
rect 839 1237 843 1241
rect 863 1235 864 1239
rect 864 1235 867 1239
rect 919 1237 923 1241
rect 1287 1236 1291 1240
rect 1327 1225 1331 1229
rect 1519 1228 1523 1232
rect 1575 1228 1579 1232
rect 1631 1228 1635 1232
rect 1687 1228 1691 1232
rect 1743 1228 1747 1232
rect 1799 1228 1803 1232
rect 1855 1228 1859 1232
rect 1911 1228 1915 1232
rect 1967 1228 1971 1232
rect 2031 1228 2035 1232
rect 2103 1228 2107 1232
rect 2183 1228 2187 1232
rect 2271 1228 2275 1232
rect 2367 1228 2371 1232
rect 2439 1228 2443 1232
rect 2503 1225 2507 1229
rect 111 1219 115 1223
rect 135 1216 139 1220
rect 199 1216 203 1220
rect 287 1216 291 1220
rect 375 1216 379 1220
rect 455 1216 459 1220
rect 535 1216 539 1220
rect 607 1216 611 1220
rect 679 1216 683 1220
rect 751 1216 755 1220
rect 823 1216 827 1220
rect 903 1216 907 1220
rect 1287 1219 1291 1223
rect 1327 1208 1331 1212
rect 1535 1207 1539 1211
rect 1571 1207 1575 1211
rect 1591 1207 1595 1211
rect 1607 1207 1611 1211
rect 1647 1207 1651 1211
rect 1683 1207 1687 1211
rect 1703 1207 1707 1211
rect 1739 1207 1743 1211
rect 1759 1207 1763 1211
rect 1795 1207 1799 1211
rect 1815 1207 1819 1211
rect 1851 1207 1855 1211
rect 1871 1207 1875 1211
rect 1907 1207 1911 1211
rect 1927 1207 1931 1211
rect 1963 1207 1967 1211
rect 1983 1207 1987 1211
rect 2027 1207 2031 1211
rect 2047 1207 2051 1211
rect 2067 1207 2068 1211
rect 2068 1207 2071 1211
rect 2119 1207 2123 1211
rect 2179 1207 2183 1211
rect 2199 1207 2203 1211
rect 2267 1207 2271 1211
rect 2287 1207 2291 1211
rect 2307 1207 2308 1211
rect 2308 1207 2311 1211
rect 2383 1207 2387 1211
rect 2391 1207 2395 1211
rect 2455 1207 2459 1211
rect 2463 1207 2467 1211
rect 2503 1208 2507 1212
rect 111 1197 115 1201
rect 135 1200 139 1204
rect 191 1200 195 1204
rect 271 1200 275 1204
rect 351 1200 355 1204
rect 431 1200 435 1204
rect 511 1200 515 1204
rect 583 1200 587 1204
rect 647 1200 651 1204
rect 719 1200 723 1204
rect 791 1200 795 1204
rect 863 1200 867 1204
rect 1287 1197 1291 1201
rect 1719 1195 1723 1199
rect 111 1180 115 1184
rect 151 1179 155 1183
rect 187 1179 191 1183
rect 207 1179 211 1183
rect 267 1179 271 1183
rect 287 1179 291 1183
rect 347 1179 351 1183
rect 367 1179 371 1183
rect 383 1179 387 1183
rect 447 1179 451 1183
rect 463 1179 467 1183
rect 527 1179 531 1183
rect 599 1179 603 1183
rect 643 1179 647 1183
rect 663 1179 667 1183
rect 715 1179 719 1183
rect 735 1179 739 1183
rect 787 1179 791 1183
rect 807 1179 811 1183
rect 859 1179 863 1183
rect 879 1179 883 1183
rect 887 1179 891 1183
rect 1287 1180 1291 1184
rect 1571 1187 1572 1191
rect 1572 1187 1575 1191
rect 1683 1187 1684 1191
rect 1684 1187 1687 1191
rect 1739 1187 1740 1191
rect 1740 1187 1743 1191
rect 1795 1187 1796 1191
rect 1796 1187 1799 1191
rect 1851 1187 1852 1191
rect 1852 1187 1855 1191
rect 1907 1187 1908 1191
rect 1908 1187 1911 1191
rect 1963 1187 1964 1191
rect 1964 1187 1967 1191
rect 2027 1187 2028 1191
rect 2028 1187 2031 1191
rect 2111 1187 2115 1191
rect 2179 1187 2180 1191
rect 2180 1187 2183 1191
rect 2267 1187 2268 1191
rect 2268 1187 2271 1191
rect 1807 1179 1811 1183
rect 2471 1187 2475 1191
rect 2475 1179 2479 1183
rect 399 1167 403 1171
rect 1599 1171 1603 1175
rect 1655 1171 1659 1175
rect 1727 1171 1731 1175
rect 187 1159 188 1163
rect 188 1159 191 1163
rect 267 1159 268 1163
rect 268 1159 271 1163
rect 347 1159 348 1163
rect 348 1159 351 1163
rect 495 1159 499 1163
rect 631 1159 635 1163
rect 643 1159 644 1163
rect 644 1159 647 1163
rect 715 1159 716 1163
rect 716 1159 719 1163
rect 787 1159 788 1163
rect 788 1159 791 1163
rect 859 1159 860 1163
rect 860 1159 863 1163
rect 1783 1163 1787 1167
rect 2307 1171 2308 1175
rect 2308 1171 2311 1175
rect 2463 1171 2467 1175
rect 887 1151 891 1155
rect 1327 1152 1331 1156
rect 1567 1153 1571 1157
rect 1599 1151 1603 1155
rect 1631 1153 1635 1157
rect 1655 1151 1656 1155
rect 1656 1151 1659 1155
rect 1703 1153 1707 1157
rect 1727 1151 1728 1155
rect 1728 1151 1731 1155
rect 1791 1153 1795 1157
rect 1807 1151 1811 1155
rect 1903 1153 1907 1157
rect 1919 1151 1923 1155
rect 2031 1153 2035 1157
rect 2175 1153 2179 1157
rect 2327 1153 2331 1157
rect 2455 1153 2459 1157
rect 2463 1151 2467 1155
rect 2503 1152 2507 1156
rect 383 1143 387 1147
rect 579 1143 583 1147
rect 759 1143 763 1147
rect 827 1143 831 1147
rect 903 1143 907 1147
rect 983 1143 987 1147
rect 1327 1135 1331 1139
rect 1551 1132 1555 1136
rect 1615 1132 1619 1136
rect 1687 1132 1691 1136
rect 1775 1132 1779 1136
rect 1887 1132 1891 1136
rect 2015 1132 2019 1136
rect 2159 1132 2163 1136
rect 2311 1132 2315 1136
rect 2439 1132 2443 1136
rect 2503 1135 2507 1139
rect 111 1124 115 1128
rect 183 1125 187 1129
rect 199 1123 203 1127
rect 279 1125 283 1129
rect 375 1125 379 1129
rect 471 1125 475 1129
rect 495 1123 496 1127
rect 496 1123 499 1127
rect 567 1125 571 1129
rect 655 1125 659 1129
rect 735 1125 739 1129
rect 759 1123 760 1127
rect 760 1123 763 1127
rect 807 1125 811 1129
rect 827 1123 828 1127
rect 828 1123 831 1127
rect 879 1125 883 1129
rect 903 1123 904 1127
rect 904 1123 907 1127
rect 959 1125 963 1129
rect 983 1123 984 1127
rect 984 1123 987 1127
rect 1039 1125 1043 1129
rect 1063 1123 1064 1127
rect 1064 1123 1067 1127
rect 1287 1124 1291 1128
rect 1327 1117 1331 1121
rect 1383 1120 1387 1124
rect 1447 1120 1451 1124
rect 1519 1120 1523 1124
rect 1591 1120 1595 1124
rect 1671 1120 1675 1124
rect 1751 1120 1755 1124
rect 1831 1120 1835 1124
rect 1911 1120 1915 1124
rect 1983 1120 1987 1124
rect 2055 1120 2059 1124
rect 2135 1120 2139 1124
rect 2215 1120 2219 1124
rect 2503 1117 2507 1121
rect 111 1107 115 1111
rect 167 1104 171 1108
rect 263 1104 267 1108
rect 359 1104 363 1108
rect 455 1104 459 1108
rect 551 1104 555 1108
rect 639 1104 643 1108
rect 719 1104 723 1108
rect 791 1104 795 1108
rect 863 1104 867 1108
rect 943 1104 947 1108
rect 1023 1104 1027 1108
rect 1287 1107 1291 1111
rect 1327 1100 1331 1104
rect 1399 1099 1403 1103
rect 1443 1099 1447 1103
rect 1463 1099 1467 1103
rect 1515 1099 1519 1103
rect 1535 1099 1539 1103
rect 1587 1099 1591 1103
rect 1607 1099 1611 1103
rect 1667 1099 1671 1103
rect 1687 1099 1691 1103
rect 1747 1099 1751 1103
rect 1767 1099 1771 1103
rect 1783 1099 1787 1103
rect 1847 1099 1851 1103
rect 1907 1099 1911 1103
rect 1927 1099 1931 1103
rect 1979 1099 1983 1103
rect 1999 1099 2003 1103
rect 2051 1099 2055 1103
rect 2071 1099 2075 1103
rect 2131 1099 2135 1103
rect 2151 1099 2155 1103
rect 2211 1099 2215 1103
rect 2231 1099 2235 1103
rect 2239 1099 2243 1103
rect 2503 1100 2507 1104
rect 111 1081 115 1085
rect 207 1084 211 1088
rect 279 1084 283 1088
rect 359 1084 363 1088
rect 447 1084 451 1088
rect 543 1084 547 1088
rect 639 1084 643 1088
rect 727 1084 731 1088
rect 815 1084 819 1088
rect 895 1084 899 1088
rect 975 1084 979 1088
rect 1055 1084 1059 1088
rect 1143 1084 1147 1088
rect 1919 1087 1923 1091
rect 1287 1081 1291 1085
rect 1443 1079 1444 1083
rect 1444 1079 1447 1083
rect 1515 1079 1516 1083
rect 1516 1079 1519 1083
rect 1587 1079 1588 1083
rect 1588 1079 1591 1083
rect 1667 1079 1668 1083
rect 1668 1079 1671 1083
rect 1747 1079 1748 1083
rect 1748 1079 1751 1083
rect 1907 1079 1908 1083
rect 1908 1079 1911 1083
rect 1979 1079 1980 1083
rect 1980 1079 1983 1083
rect 2051 1079 2052 1083
rect 2052 1079 2055 1083
rect 2131 1079 2132 1083
rect 2132 1079 2135 1083
rect 2211 1079 2212 1083
rect 2212 1079 2215 1083
rect 1835 1071 1839 1075
rect 111 1064 115 1068
rect 223 1063 227 1067
rect 275 1063 279 1067
rect 295 1063 299 1067
rect 355 1063 359 1067
rect 375 1063 379 1067
rect 443 1063 447 1067
rect 463 1063 467 1067
rect 471 1063 475 1067
rect 559 1063 563 1067
rect 579 1063 580 1067
rect 580 1063 583 1067
rect 655 1063 659 1067
rect 743 1063 747 1067
rect 811 1063 815 1067
rect 831 1063 835 1067
rect 891 1063 895 1067
rect 911 1063 915 1067
rect 971 1063 975 1067
rect 991 1063 995 1067
rect 1051 1063 1055 1067
rect 1071 1063 1075 1067
rect 1139 1063 1143 1067
rect 1159 1063 1163 1067
rect 1167 1063 1171 1067
rect 1287 1064 1291 1068
rect 2239 1067 2243 1071
rect 1063 1051 1067 1055
rect 1391 1059 1395 1063
rect 1479 1059 1483 1063
rect 1599 1059 1603 1063
rect 1719 1059 1723 1063
rect 1951 1059 1955 1063
rect 2063 1059 2067 1063
rect 2175 1059 2179 1063
rect 2279 1059 2283 1063
rect 2463 1059 2467 1063
rect 1711 1051 1715 1055
rect 199 1043 203 1047
rect 275 1043 276 1047
rect 276 1043 279 1047
rect 355 1043 356 1047
rect 356 1043 359 1047
rect 443 1043 444 1047
rect 444 1043 447 1047
rect 599 1043 603 1047
rect 811 1043 812 1047
rect 812 1043 815 1047
rect 891 1043 892 1047
rect 892 1043 895 1047
rect 971 1043 972 1047
rect 972 1043 975 1047
rect 1051 1043 1052 1047
rect 1052 1043 1055 1047
rect 1139 1043 1140 1047
rect 1140 1043 1143 1047
rect 1327 1040 1331 1044
rect 1367 1041 1371 1045
rect 1391 1039 1392 1043
rect 1392 1039 1395 1043
rect 1455 1041 1459 1045
rect 1479 1039 1480 1043
rect 1480 1039 1483 1043
rect 1575 1041 1579 1045
rect 1599 1039 1600 1043
rect 1600 1039 1603 1043
rect 1695 1041 1699 1045
rect 1719 1039 1720 1043
rect 1720 1039 1723 1043
rect 1815 1041 1819 1045
rect 1835 1039 1836 1043
rect 1836 1039 1839 1043
rect 1927 1041 1931 1045
rect 1951 1039 1952 1043
rect 1952 1039 1955 1043
rect 2039 1041 2043 1045
rect 2063 1039 2064 1043
rect 2064 1039 2067 1043
rect 2151 1041 2155 1045
rect 2175 1039 2176 1043
rect 2176 1039 2179 1043
rect 2255 1041 2259 1045
rect 2279 1039 2280 1043
rect 2280 1039 2283 1043
rect 2367 1041 2371 1045
rect 2375 1039 2379 1043
rect 2455 1041 2459 1045
rect 2463 1039 2467 1043
rect 2503 1040 2507 1044
rect 1167 1031 1171 1035
rect 471 1023 475 1027
rect 691 1023 695 1027
rect 791 1023 795 1027
rect 879 1023 883 1027
rect 967 1023 971 1027
rect 1047 1023 1051 1027
rect 1207 1023 1211 1027
rect 1327 1023 1331 1027
rect 1351 1020 1355 1024
rect 1439 1020 1443 1024
rect 1559 1020 1563 1024
rect 1679 1020 1683 1024
rect 1799 1020 1803 1024
rect 1911 1020 1915 1024
rect 2023 1020 2027 1024
rect 2135 1020 2139 1024
rect 2239 1020 2243 1024
rect 2351 1020 2355 1024
rect 2439 1020 2443 1024
rect 2503 1023 2507 1027
rect 1215 1011 1219 1015
rect 111 1004 115 1008
rect 295 1005 299 1009
rect 303 1003 307 1007
rect 383 1005 387 1009
rect 479 1005 483 1009
rect 575 1005 579 1009
rect 599 1003 600 1007
rect 600 1003 603 1007
rect 671 1005 675 1009
rect 767 1005 771 1009
rect 791 1003 792 1007
rect 792 1003 795 1007
rect 855 1005 859 1009
rect 879 1003 880 1007
rect 880 1003 883 1007
rect 943 1005 947 1009
rect 967 1003 968 1007
rect 968 1003 971 1007
rect 1023 1005 1027 1009
rect 1103 1005 1107 1009
rect 1183 1005 1187 1009
rect 1207 1003 1208 1007
rect 1208 1003 1211 1007
rect 1239 1005 1243 1009
rect 1279 1003 1283 1007
rect 1287 1004 1291 1008
rect 1327 1001 1331 1005
rect 1351 1004 1355 1008
rect 1511 1004 1515 1008
rect 1679 1004 1683 1008
rect 1823 1004 1827 1008
rect 1951 1004 1955 1008
rect 2071 1004 2075 1008
rect 2175 1004 2179 1008
rect 2271 1004 2275 1008
rect 2367 1004 2371 1008
rect 2439 1004 2443 1008
rect 2503 1001 2507 1005
rect 111 987 115 991
rect 279 984 283 988
rect 367 984 371 988
rect 463 984 467 988
rect 559 984 563 988
rect 655 984 659 988
rect 751 984 755 988
rect 839 984 843 988
rect 927 984 931 988
rect 1007 984 1011 988
rect 1087 984 1091 988
rect 1167 984 1171 988
rect 1223 984 1227 988
rect 1287 987 1291 991
rect 1327 984 1331 988
rect 1367 983 1371 987
rect 1375 983 1379 987
rect 1527 983 1531 987
rect 1675 983 1679 987
rect 1695 983 1699 987
rect 1711 983 1715 987
rect 1839 983 1843 987
rect 1947 983 1951 987
rect 1967 983 1971 987
rect 2067 983 2071 987
rect 2087 983 2091 987
rect 2171 983 2175 987
rect 2191 983 2195 987
rect 2267 983 2271 987
rect 2287 983 2291 987
rect 2363 983 2367 987
rect 2383 983 2387 987
rect 2391 983 2395 987
rect 2455 983 2459 987
rect 2475 983 2476 987
rect 2476 983 2479 987
rect 2503 984 2507 988
rect 111 969 115 973
rect 271 972 275 976
rect 359 972 363 976
rect 455 972 459 976
rect 551 972 555 976
rect 655 972 659 976
rect 751 972 755 976
rect 839 972 843 976
rect 927 972 931 976
rect 1007 972 1011 976
rect 1087 972 1091 976
rect 1167 972 1171 976
rect 1223 972 1227 976
rect 1279 975 1283 979
rect 1287 969 1291 973
rect 1675 963 1676 967
rect 1676 963 1679 967
rect 1823 963 1824 967
rect 1824 963 1827 967
rect 1947 963 1948 967
rect 1948 963 1951 967
rect 2067 963 2068 967
rect 2068 963 2071 967
rect 2171 963 2172 967
rect 2172 963 2175 967
rect 2267 963 2268 967
rect 2268 963 2271 967
rect 2363 963 2364 967
rect 2364 963 2367 967
rect 2447 963 2451 967
rect 111 952 115 956
rect 287 951 291 955
rect 355 951 359 955
rect 375 951 379 955
rect 451 951 455 955
rect 471 951 475 955
rect 479 951 483 955
rect 567 951 571 955
rect 651 951 655 955
rect 671 951 675 955
rect 691 951 692 955
rect 692 951 695 955
rect 767 951 771 955
rect 835 951 839 955
rect 855 951 859 955
rect 923 951 927 955
rect 943 951 947 955
rect 1003 951 1007 955
rect 1023 951 1027 955
rect 1047 951 1048 955
rect 1048 951 1051 955
rect 1103 951 1107 955
rect 1183 951 1187 955
rect 1239 951 1243 955
rect 1287 952 1291 956
rect 1375 939 1379 943
rect 1391 939 1395 943
rect 1447 939 1451 943
rect 1535 939 1539 943
rect 1631 939 1635 943
rect 1743 939 1747 943
rect 303 931 307 935
rect 355 931 356 935
rect 356 931 359 935
rect 451 931 452 935
rect 452 931 455 935
rect 463 931 467 935
rect 651 931 652 935
rect 652 931 655 935
rect 835 931 836 935
rect 836 931 839 935
rect 923 931 924 935
rect 924 931 927 935
rect 1003 931 1004 935
rect 1004 931 1007 935
rect 1203 931 1207 935
rect 1215 931 1219 935
rect 1439 927 1443 931
rect 1959 939 1963 943
rect 2055 939 2059 943
rect 2391 939 2395 943
rect 2463 939 2467 943
rect 479 919 483 923
rect 1327 920 1331 924
rect 1367 921 1371 925
rect 1391 919 1392 923
rect 1392 919 1395 923
rect 1423 921 1427 925
rect 1447 919 1448 923
rect 1448 919 1451 923
rect 1503 921 1507 925
rect 1535 919 1539 923
rect 1607 921 1611 925
rect 1631 919 1632 923
rect 1632 919 1635 923
rect 1719 921 1723 925
rect 1743 919 1744 923
rect 1744 919 1747 923
rect 1831 921 1835 925
rect 1935 921 1939 925
rect 1959 919 1960 923
rect 1960 919 1963 923
rect 2031 921 2035 925
rect 2055 919 2056 923
rect 2056 919 2059 923
rect 2127 921 2131 925
rect 2151 919 2152 923
rect 2152 919 2155 923
rect 2215 921 2219 925
rect 2295 921 2299 925
rect 2375 921 2379 925
rect 2455 921 2459 925
rect 2463 919 2467 923
rect 2503 920 2507 924
rect 279 911 283 915
rect 295 911 299 915
rect 447 911 451 915
rect 543 911 547 915
rect 639 911 643 915
rect 831 911 835 915
rect 927 911 931 915
rect 1015 911 1019 915
rect 463 899 467 903
rect 939 903 943 907
rect 1327 903 1331 907
rect 1351 900 1355 904
rect 1407 900 1411 904
rect 1487 900 1491 904
rect 1591 900 1595 904
rect 1703 900 1707 904
rect 1815 900 1819 904
rect 1919 900 1923 904
rect 2015 900 2019 904
rect 2111 900 2115 904
rect 2199 900 2203 904
rect 2279 900 2283 904
rect 2359 900 2363 904
rect 2439 900 2443 904
rect 2503 903 2507 907
rect 111 892 115 896
rect 271 893 275 897
rect 295 891 296 895
rect 296 891 299 895
rect 343 893 347 897
rect 423 893 427 897
rect 447 891 448 895
rect 448 891 451 895
rect 519 893 523 897
rect 543 891 544 895
rect 544 891 547 895
rect 615 893 619 897
rect 639 891 640 895
rect 640 891 643 895
rect 711 893 715 897
rect 719 891 723 895
rect 807 893 811 897
rect 831 891 832 895
rect 832 891 835 895
rect 903 893 907 897
rect 927 891 928 895
rect 928 891 931 895
rect 991 893 995 897
rect 1015 891 1016 895
rect 1016 891 1019 895
rect 1087 893 1091 897
rect 1183 893 1187 897
rect 1203 891 1204 895
rect 1204 891 1207 895
rect 1287 892 1291 896
rect 1327 881 1331 885
rect 1431 884 1435 888
rect 1487 884 1491 888
rect 1551 884 1555 888
rect 1623 884 1627 888
rect 1703 884 1707 888
rect 1791 884 1795 888
rect 1895 884 1899 888
rect 2015 884 2019 888
rect 2143 884 2147 888
rect 2279 884 2283 888
rect 2423 884 2427 888
rect 2503 881 2507 885
rect 111 875 115 879
rect 255 872 259 876
rect 327 872 331 876
rect 407 872 411 876
rect 503 872 507 876
rect 599 872 603 876
rect 695 872 699 876
rect 791 872 795 876
rect 887 872 891 876
rect 975 872 979 876
rect 1071 872 1075 876
rect 1167 872 1171 876
rect 1287 875 1291 879
rect 1327 864 1331 868
rect 1447 863 1451 867
rect 1483 863 1487 867
rect 1503 863 1507 867
rect 1547 863 1551 867
rect 1567 863 1571 867
rect 1619 863 1623 867
rect 1639 863 1643 867
rect 1699 863 1703 867
rect 1719 863 1723 867
rect 1727 863 1731 867
rect 1807 863 1811 867
rect 1891 863 1895 867
rect 1911 863 1915 867
rect 1919 863 1923 867
rect 2031 863 2035 867
rect 2159 863 2163 867
rect 2275 863 2279 867
rect 2295 863 2299 867
rect 111 853 115 857
rect 247 856 251 860
rect 311 856 315 860
rect 375 856 379 860
rect 439 856 443 860
rect 503 856 507 860
rect 567 856 571 860
rect 631 856 635 860
rect 695 856 699 860
rect 759 856 763 860
rect 831 856 835 860
rect 903 856 907 860
rect 1287 853 1291 857
rect 2439 863 2443 867
rect 2447 863 2451 867
rect 2503 864 2507 868
rect 1439 843 1443 847
rect 1483 843 1484 847
rect 1484 843 1487 847
rect 1547 843 1548 847
rect 1548 843 1551 847
rect 1619 843 1620 847
rect 1620 843 1623 847
rect 1699 843 1700 847
rect 1700 843 1703 847
rect 1891 843 1892 847
rect 1892 843 1895 847
rect 2151 843 2155 847
rect 2275 843 2276 847
rect 2276 843 2279 847
rect 2407 843 2411 847
rect 111 836 115 840
rect 263 835 267 839
rect 279 835 283 839
rect 327 835 331 839
rect 391 835 395 839
rect 435 835 439 839
rect 455 835 459 839
rect 499 835 503 839
rect 519 835 523 839
rect 563 835 567 839
rect 583 835 587 839
rect 591 835 595 839
rect 647 835 651 839
rect 691 835 695 839
rect 711 835 715 839
rect 755 835 759 839
rect 775 835 779 839
rect 827 835 831 839
rect 847 835 851 839
rect 899 835 903 839
rect 919 835 923 839
rect 939 835 940 839
rect 940 835 943 839
rect 1287 836 1291 840
rect 1727 835 1731 839
rect 719 823 723 827
rect 1615 827 1619 831
rect 1671 827 1675 831
rect 1727 827 1731 831
rect 1919 827 1923 831
rect 1951 827 1955 831
rect 2039 827 2043 831
rect 2215 827 2219 831
rect 2311 827 2315 831
rect 2463 827 2467 831
rect 319 815 323 819
rect 435 815 436 819
rect 436 815 439 819
rect 499 815 500 819
rect 500 815 503 819
rect 563 815 564 819
rect 564 815 567 819
rect 683 815 687 819
rect 691 815 692 819
rect 692 815 695 819
rect 755 815 756 819
rect 756 815 759 819
rect 827 815 828 819
rect 828 815 831 819
rect 899 815 900 819
rect 900 815 903 819
rect 2375 819 2379 823
rect 591 807 595 811
rect 1327 808 1331 812
rect 1591 809 1595 813
rect 1615 807 1616 811
rect 1616 807 1619 811
rect 1647 809 1651 813
rect 1671 807 1672 811
rect 1672 807 1675 811
rect 1703 809 1707 813
rect 1727 807 1728 811
rect 1728 807 1731 811
rect 1767 809 1771 813
rect 1847 809 1851 813
rect 1855 807 1859 811
rect 1927 809 1931 813
rect 1951 807 1952 811
rect 1952 807 1955 811
rect 2015 809 2019 813
rect 2039 807 2040 811
rect 2040 807 2043 811
rect 2103 809 2107 813
rect 2127 807 2128 811
rect 2128 807 2131 811
rect 2191 809 2195 813
rect 2215 807 2216 811
rect 2216 807 2219 811
rect 2287 809 2291 813
rect 2311 807 2312 811
rect 2312 807 2315 811
rect 2383 809 2387 813
rect 2407 807 2408 811
rect 2408 807 2411 811
rect 2455 809 2459 813
rect 2471 807 2475 811
rect 2503 808 2507 812
rect 175 799 179 803
rect 239 799 243 803
rect 415 799 419 803
rect 503 799 507 803
rect 591 799 595 803
rect 655 799 659 803
rect 683 787 687 791
rect 1075 799 1079 803
rect 1327 791 1331 795
rect 1575 788 1579 792
rect 1631 788 1635 792
rect 1687 788 1691 792
rect 1751 788 1755 792
rect 1831 788 1835 792
rect 1911 788 1915 792
rect 1999 788 2003 792
rect 2087 788 2091 792
rect 2175 788 2179 792
rect 2271 788 2275 792
rect 2367 788 2371 792
rect 2439 788 2443 792
rect 2503 791 2507 795
rect 111 780 115 784
rect 215 781 219 785
rect 239 779 240 783
rect 240 779 243 783
rect 303 781 307 785
rect 319 779 323 783
rect 391 781 395 785
rect 415 779 416 783
rect 416 779 419 783
rect 479 781 483 785
rect 503 779 504 783
rect 504 779 507 783
rect 559 781 563 785
rect 591 779 595 783
rect 631 781 635 785
rect 655 779 656 783
rect 656 779 659 783
rect 703 781 707 785
rect 767 781 771 785
rect 783 779 787 783
rect 831 781 835 785
rect 895 781 899 785
rect 967 781 971 785
rect 1039 781 1043 785
rect 1287 780 1291 784
rect 1327 769 1331 773
rect 1567 772 1571 776
rect 1623 772 1627 776
rect 1687 772 1691 776
rect 1759 772 1763 776
rect 1831 772 1835 776
rect 1919 772 1923 776
rect 2015 772 2019 776
rect 2119 772 2123 776
rect 2231 772 2235 776
rect 2343 772 2347 776
rect 2439 772 2443 776
rect 2503 769 2507 773
rect 111 763 115 767
rect 199 760 203 764
rect 287 760 291 764
rect 375 760 379 764
rect 463 760 467 764
rect 543 760 547 764
rect 615 760 619 764
rect 687 760 691 764
rect 751 760 755 764
rect 815 760 819 764
rect 879 760 883 764
rect 951 760 955 764
rect 1023 760 1027 764
rect 1287 763 1291 767
rect 111 745 115 749
rect 135 748 139 752
rect 255 748 259 752
rect 391 748 395 752
rect 519 748 523 752
rect 647 748 651 752
rect 775 748 779 752
rect 903 748 907 752
rect 1039 748 1043 752
rect 1327 752 1331 756
rect 1583 751 1587 755
rect 1619 751 1623 755
rect 1639 751 1643 755
rect 1683 751 1687 755
rect 1703 751 1707 755
rect 1719 751 1723 755
rect 1775 751 1779 755
rect 1783 751 1787 755
rect 1847 751 1851 755
rect 1287 745 1291 749
rect 1603 739 1607 743
rect 1651 739 1655 743
rect 1935 751 1939 755
rect 2011 751 2015 755
rect 2031 751 2035 755
rect 2115 751 2119 755
rect 2135 751 2139 755
rect 2227 751 2231 755
rect 2247 751 2251 755
rect 2127 739 2131 743
rect 2143 743 2147 747
rect 2359 751 2363 755
rect 2375 751 2379 755
rect 2455 751 2459 755
rect 2463 751 2467 755
rect 2503 752 2507 756
rect 111 728 115 732
rect 151 727 155 731
rect 175 727 176 731
rect 176 727 179 731
rect 271 727 275 731
rect 407 727 411 731
rect 535 727 539 731
rect 643 727 647 731
rect 663 727 667 731
rect 723 727 727 731
rect 791 727 795 731
rect 919 727 923 731
rect 1035 727 1039 731
rect 1055 727 1059 731
rect 1075 727 1076 731
rect 1076 727 1079 731
rect 1287 728 1291 732
rect 1611 731 1615 735
rect 1619 731 1620 735
rect 1620 731 1623 735
rect 1683 731 1684 735
rect 1684 731 1687 735
rect 495 707 499 711
rect 643 707 644 711
rect 644 707 647 711
rect 783 707 787 711
rect 895 707 899 711
rect 1035 707 1036 711
rect 1036 707 1039 711
rect 1603 719 1607 723
rect 1623 723 1627 727
rect 1783 727 1787 731
rect 1855 731 1859 735
rect 2011 731 2012 735
rect 2012 731 2015 735
rect 2115 731 2116 735
rect 2116 731 2119 735
rect 2227 731 2228 735
rect 2228 731 2231 735
rect 2387 731 2391 735
rect 2471 731 2475 735
rect 1719 719 1720 723
rect 1720 719 1723 723
rect 1855 719 1859 723
rect 1863 719 1867 723
rect 1967 719 1971 723
rect 2143 719 2147 723
rect 2175 719 2179 723
rect 2279 719 2283 723
rect 2463 719 2467 723
rect 175 695 179 699
rect 231 695 235 699
rect 415 695 419 699
rect 287 687 291 691
rect 495 683 499 687
rect 723 695 724 699
rect 724 695 727 699
rect 975 695 979 699
rect 1327 700 1331 704
rect 1367 701 1371 705
rect 1431 701 1435 705
rect 1527 701 1531 705
rect 1631 701 1635 705
rect 1151 695 1155 699
rect 1651 699 1652 703
rect 1652 699 1655 703
rect 1735 701 1739 705
rect 1839 701 1843 705
rect 1863 699 1864 703
rect 1864 699 1867 703
rect 1943 701 1947 705
rect 1967 699 1968 703
rect 1968 699 1971 703
rect 2047 701 2051 705
rect 2063 699 2067 703
rect 2151 701 2155 705
rect 2175 699 2176 703
rect 2176 699 2179 703
rect 2255 701 2259 705
rect 2279 699 2280 703
rect 2280 699 2283 703
rect 2367 701 2371 705
rect 2387 699 2388 703
rect 2388 699 2391 703
rect 2455 701 2459 705
rect 2471 699 2475 703
rect 2503 700 2507 704
rect 1327 683 1331 687
rect 111 676 115 680
rect 151 677 155 681
rect 175 675 176 679
rect 176 675 179 679
rect 207 677 211 681
rect 231 675 232 679
rect 232 675 235 679
rect 295 677 299 681
rect 391 677 395 681
rect 415 675 416 679
rect 416 675 419 679
rect 503 677 507 681
rect 623 677 627 681
rect 647 675 648 679
rect 648 675 651 679
rect 743 677 747 681
rect 871 677 875 681
rect 895 675 896 679
rect 896 675 899 679
rect 999 677 1003 681
rect 1127 677 1131 681
rect 1151 675 1152 679
rect 1152 675 1155 679
rect 1239 677 1243 681
rect 1287 676 1291 680
rect 1351 680 1355 684
rect 1415 680 1419 684
rect 1511 680 1515 684
rect 1615 680 1619 684
rect 1719 680 1723 684
rect 1823 680 1827 684
rect 1927 680 1931 684
rect 2031 680 2035 684
rect 2135 680 2139 684
rect 2239 680 2243 684
rect 2351 680 2355 684
rect 2439 680 2443 684
rect 2503 683 2507 687
rect 1343 667 1347 671
rect 111 659 115 663
rect 135 656 139 660
rect 191 656 195 660
rect 279 656 283 660
rect 375 656 379 660
rect 487 656 491 660
rect 607 656 611 660
rect 727 656 731 660
rect 855 656 859 660
rect 983 656 987 660
rect 1111 656 1115 660
rect 1223 656 1227 660
rect 1287 659 1291 663
rect 1327 653 1331 657
rect 1351 656 1355 660
rect 1415 656 1419 660
rect 1511 656 1515 660
rect 1607 656 1611 660
rect 1711 656 1715 660
rect 1823 656 1827 660
rect 1935 656 1939 660
rect 2055 656 2059 660
rect 2183 656 2187 660
rect 2319 656 2323 660
rect 2439 656 2443 660
rect 2503 653 2507 657
rect 111 637 115 641
rect 151 640 155 644
rect 263 640 267 644
rect 367 640 371 644
rect 463 640 467 644
rect 559 640 563 644
rect 655 640 659 644
rect 751 640 755 644
rect 847 640 851 644
rect 943 640 947 644
rect 1039 640 1043 644
rect 1143 640 1147 644
rect 1223 640 1227 644
rect 1287 637 1291 641
rect 1327 636 1331 640
rect 1367 635 1371 639
rect 1411 635 1415 639
rect 1431 635 1435 639
rect 1507 635 1511 639
rect 1527 635 1531 639
rect 1535 635 1539 639
rect 1623 635 1627 639
rect 1263 627 1267 631
rect 1727 635 1731 639
rect 1839 635 1843 639
rect 1855 635 1859 639
rect 1951 635 1955 639
rect 2071 635 2075 639
rect 2179 635 2183 639
rect 2199 635 2203 639
rect 2315 635 2319 639
rect 2335 635 2339 639
rect 2351 635 2355 639
rect 2455 635 2459 639
rect 2463 635 2467 639
rect 2503 636 2507 640
rect 111 620 115 624
rect 167 619 171 623
rect 259 619 263 623
rect 279 619 283 623
rect 287 619 291 623
rect 383 619 387 623
rect 407 619 408 623
rect 408 619 411 623
rect 479 619 483 623
rect 487 619 491 623
rect 575 619 579 623
rect 671 619 675 623
rect 767 619 771 623
rect 843 619 847 623
rect 863 619 867 623
rect 939 619 943 623
rect 959 619 963 623
rect 975 619 979 623
rect 1055 619 1059 623
rect 1139 619 1143 623
rect 1159 619 1163 623
rect 1167 619 1171 623
rect 1239 619 1243 623
rect 1287 620 1291 624
rect 1343 615 1347 619
rect 1411 615 1412 619
rect 1412 615 1415 619
rect 1507 615 1508 619
rect 1508 615 1511 619
rect 1535 611 1539 615
rect 1763 615 1767 619
rect 2043 615 2047 619
rect 2063 615 2067 619
rect 2179 615 2180 619
rect 2180 615 2183 619
rect 2315 615 2316 619
rect 2316 615 2319 619
rect 2471 615 2475 619
rect 159 599 163 603
rect 259 599 260 603
rect 260 599 263 603
rect 487 595 491 599
rect 647 599 651 603
rect 835 599 839 603
rect 843 599 844 603
rect 844 599 847 603
rect 939 599 940 603
rect 940 599 943 603
rect 1019 595 1023 599
rect 1139 599 1140 603
rect 1140 599 1143 603
rect 1263 599 1267 603
rect 1575 603 1579 607
rect 1587 595 1591 599
rect 1871 603 1875 607
rect 1983 603 1987 607
rect 1891 595 1895 599
rect 287 587 291 591
rect 407 587 411 591
rect 455 587 459 591
rect 559 587 563 591
rect 743 587 747 591
rect 751 587 755 591
rect 1167 587 1168 591
rect 1168 587 1171 591
rect 2043 591 2047 595
rect 2351 603 2355 607
rect 2463 603 2467 607
rect 1327 584 1331 588
rect 1383 585 1387 589
rect 1399 583 1403 587
rect 1463 585 1467 589
rect 1551 585 1555 589
rect 1575 583 1576 587
rect 1576 583 1579 587
rect 1647 585 1651 589
rect 1743 585 1747 589
rect 1763 583 1764 587
rect 1764 583 1767 587
rect 1847 585 1851 589
rect 1871 583 1872 587
rect 1872 583 1875 587
rect 1959 585 1963 589
rect 1983 583 1984 587
rect 1984 583 1987 587
rect 2079 585 2083 589
rect 2207 585 2211 589
rect 2215 583 2219 587
rect 2343 585 2347 589
rect 2455 585 2459 589
rect 2463 583 2467 587
rect 2503 584 2507 588
rect 111 568 115 572
rect 151 569 155 573
rect 159 567 163 571
rect 239 569 243 573
rect 335 569 339 573
rect 431 569 435 573
rect 455 567 456 571
rect 456 567 459 571
rect 535 569 539 573
rect 559 567 560 571
rect 560 567 563 571
rect 631 569 635 573
rect 647 567 651 571
rect 727 569 731 573
rect 751 567 752 571
rect 752 567 755 571
rect 823 569 827 573
rect 835 567 839 571
rect 911 569 915 573
rect 943 567 947 571
rect 999 569 1003 573
rect 1019 567 1020 571
rect 1020 567 1023 571
rect 1087 569 1091 573
rect 1183 569 1187 573
rect 1287 568 1291 572
rect 1327 567 1331 571
rect 1367 564 1371 568
rect 1447 564 1451 568
rect 1535 564 1539 568
rect 1631 564 1635 568
rect 1727 564 1731 568
rect 1831 564 1835 568
rect 1943 564 1947 568
rect 2063 564 2067 568
rect 2191 564 2195 568
rect 2327 564 2331 568
rect 2439 564 2443 568
rect 2503 567 2507 571
rect 111 551 115 555
rect 135 548 139 552
rect 223 548 227 552
rect 319 548 323 552
rect 415 548 419 552
rect 519 548 523 552
rect 615 548 619 552
rect 711 548 715 552
rect 807 548 811 552
rect 895 548 899 552
rect 983 548 987 552
rect 1071 548 1075 552
rect 1167 548 1171 552
rect 1287 551 1291 555
rect 1327 549 1331 553
rect 1375 552 1379 556
rect 1455 552 1459 556
rect 1551 552 1555 556
rect 1647 552 1651 556
rect 1751 552 1755 556
rect 1855 552 1859 556
rect 1959 552 1963 556
rect 2055 552 2059 556
rect 2151 552 2155 556
rect 2255 552 2259 556
rect 2359 552 2363 556
rect 2439 552 2443 556
rect 2503 549 2507 553
rect 111 525 115 529
rect 143 528 147 532
rect 239 528 243 532
rect 335 528 339 532
rect 431 528 435 532
rect 527 528 531 532
rect 623 528 627 532
rect 711 528 715 532
rect 791 528 795 532
rect 871 528 875 532
rect 951 528 955 532
rect 1031 528 1035 532
rect 1327 532 1331 536
rect 1391 531 1395 535
rect 1451 531 1455 535
rect 1471 531 1475 535
rect 1479 531 1483 535
rect 1567 531 1571 535
rect 1587 531 1588 535
rect 1588 531 1591 535
rect 1663 531 1667 535
rect 1767 531 1771 535
rect 1287 525 1291 529
rect 1871 531 1875 535
rect 1891 531 1892 535
rect 1892 531 1895 535
rect 1975 531 1979 535
rect 2071 531 2075 535
rect 2147 531 2151 535
rect 2167 531 2171 535
rect 2251 531 2255 535
rect 2271 531 2275 535
rect 2279 531 2283 535
rect 2375 531 2379 535
rect 2391 531 2395 535
rect 2455 531 2459 535
rect 2471 531 2475 535
rect 2503 532 2507 536
rect 2215 519 2219 523
rect 111 508 115 512
rect 159 507 163 511
rect 235 507 239 511
rect 255 507 259 511
rect 287 507 291 511
rect 351 507 355 511
rect 427 507 431 511
rect 447 507 451 511
rect 455 507 459 511
rect 543 507 547 511
rect 639 507 643 511
rect 707 507 711 511
rect 727 507 731 511
rect 743 507 747 511
rect 807 507 811 511
rect 827 507 828 511
rect 828 507 831 511
rect 887 507 891 511
rect 647 495 651 499
rect 967 507 971 511
rect 1027 507 1031 511
rect 1047 507 1051 511
rect 1287 508 1291 512
rect 1399 511 1403 515
rect 1451 511 1452 515
rect 1452 511 1455 515
rect 1827 511 1831 515
rect 1943 511 1947 515
rect 2147 511 2148 515
rect 2148 511 2151 515
rect 2251 511 2252 515
rect 2252 511 2255 515
rect 2415 511 2419 515
rect 2463 511 2467 515
rect 2391 503 2395 507
rect 171 487 175 491
rect 235 487 236 491
rect 236 487 239 491
rect 427 487 428 491
rect 428 487 431 491
rect 675 487 679 491
rect 707 487 708 491
rect 708 487 711 491
rect 943 487 947 491
rect 1027 487 1028 491
rect 1028 487 1031 491
rect 1479 495 1483 499
rect 1599 495 1603 499
rect 1719 495 1723 499
rect 1963 495 1967 499
rect 1619 487 1623 491
rect 2047 495 2051 499
rect 2279 495 2280 499
rect 2280 495 2283 499
rect 2315 495 2319 499
rect 2447 495 2451 499
rect 579 479 583 483
rect 2415 483 2419 487
rect 303 467 307 471
rect 311 471 315 475
rect 455 471 459 475
rect 487 471 491 475
rect 743 471 747 475
rect 827 471 828 475
rect 828 471 831 475
rect 871 471 875 475
rect 975 471 979 475
rect 1327 476 1331 480
rect 1367 477 1371 481
rect 1455 477 1459 481
rect 1575 477 1579 481
rect 1599 475 1600 479
rect 1600 475 1603 479
rect 1695 477 1699 481
rect 1719 475 1720 479
rect 1720 475 1723 479
rect 1807 477 1811 481
rect 1827 475 1828 479
rect 1828 475 1831 479
rect 1919 477 1923 481
rect 1943 475 1944 479
rect 1944 475 1947 479
rect 2023 477 2027 481
rect 2047 475 2048 479
rect 2048 475 2051 479
rect 2119 477 2123 481
rect 2167 475 2171 479
rect 2207 477 2211 481
rect 2295 477 2299 481
rect 2315 475 2316 479
rect 2316 475 2319 479
rect 2383 477 2387 481
rect 2399 475 2403 479
rect 2455 477 2459 481
rect 2503 476 2507 480
rect 839 459 843 463
rect 1327 459 1331 463
rect 111 452 115 456
rect 151 453 155 457
rect 171 451 172 455
rect 172 451 175 455
rect 207 453 211 457
rect 287 453 291 457
rect 311 451 312 455
rect 312 451 315 455
rect 375 453 379 457
rect 391 451 395 455
rect 463 453 467 457
rect 487 451 488 455
rect 488 451 491 455
rect 559 453 563 457
rect 579 451 580 455
rect 580 451 583 455
rect 655 453 659 457
rect 675 451 676 455
rect 676 451 679 455
rect 751 453 755 457
rect 847 453 851 457
rect 871 451 872 455
rect 872 451 875 455
rect 951 453 955 457
rect 975 451 976 455
rect 976 451 979 455
rect 1055 453 1059 457
rect 1159 453 1163 457
rect 1167 451 1171 455
rect 1239 453 1243 457
rect 1287 452 1291 456
rect 1351 456 1355 460
rect 1439 456 1443 460
rect 1559 456 1563 460
rect 1679 456 1683 460
rect 1791 456 1795 460
rect 1903 456 1907 460
rect 2007 456 2011 460
rect 2103 456 2107 460
rect 2191 456 2195 460
rect 2279 456 2283 460
rect 2367 456 2371 460
rect 2439 456 2443 460
rect 2503 459 2507 463
rect 111 435 115 439
rect 135 432 139 436
rect 191 432 195 436
rect 271 432 275 436
rect 359 432 363 436
rect 447 432 451 436
rect 543 432 547 436
rect 639 432 643 436
rect 735 432 739 436
rect 831 432 835 436
rect 935 432 939 436
rect 1039 432 1043 436
rect 1143 432 1147 436
rect 1223 432 1227 436
rect 1287 435 1291 439
rect 1327 429 1331 433
rect 1583 432 1587 436
rect 1639 432 1643 436
rect 1695 432 1699 436
rect 1759 432 1763 436
rect 1831 432 1835 436
rect 1911 432 1915 436
rect 1991 432 1995 436
rect 2079 432 2083 436
rect 2175 432 2179 436
rect 2271 432 2275 436
rect 2367 432 2371 436
rect 2439 432 2443 436
rect 2503 429 2507 433
rect 111 417 115 421
rect 135 420 139 424
rect 191 420 195 424
rect 279 420 283 424
rect 383 420 387 424
rect 495 420 499 424
rect 607 420 611 424
rect 719 420 723 424
rect 831 420 835 424
rect 935 420 939 424
rect 1039 420 1043 424
rect 1143 420 1147 424
rect 1223 420 1227 424
rect 1287 417 1291 421
rect 1327 412 1331 416
rect 1599 411 1603 415
rect 1619 411 1620 415
rect 1620 411 1623 415
rect 1655 411 1659 415
rect 1711 411 1715 415
rect 111 400 115 404
rect 151 399 155 403
rect 187 399 191 403
rect 207 399 211 403
rect 275 399 279 403
rect 295 399 299 403
rect 303 399 307 403
rect 399 399 403 403
rect 491 399 495 403
rect 511 399 515 403
rect 603 399 607 403
rect 623 399 627 403
rect 631 399 635 403
rect 735 399 739 403
rect 743 399 747 403
rect 847 399 851 403
rect 931 399 935 403
rect 951 399 955 403
rect 995 399 999 403
rect 1055 399 1059 403
rect 1075 399 1076 403
rect 1076 399 1079 403
rect 1159 399 1163 403
rect 1219 399 1223 403
rect 1239 399 1243 403
rect 1287 400 1291 404
rect 1775 411 1779 415
rect 1847 411 1851 415
rect 1927 411 1931 415
rect 1987 411 1991 415
rect 2007 411 2011 415
rect 2075 411 2079 415
rect 2095 411 2099 415
rect 2103 411 2107 415
rect 2191 411 2195 415
rect 2267 411 2271 415
rect 2287 411 2291 415
rect 2295 411 2299 415
rect 2383 411 2387 415
rect 2391 411 2395 415
rect 2455 411 2459 415
rect 2463 411 2467 415
rect 2503 412 2507 416
rect 1887 391 1891 395
rect 1895 391 1899 395
rect 1987 391 1988 395
rect 1988 391 1991 395
rect 2075 391 2076 395
rect 2076 391 2079 395
rect 2167 391 2171 395
rect 2267 391 2268 395
rect 2268 391 2271 395
rect 2399 391 2403 395
rect 2471 391 2475 395
rect 171 379 175 383
rect 187 379 188 383
rect 188 379 191 383
rect 275 379 276 383
rect 276 379 279 383
rect 391 379 395 383
rect 491 379 492 383
rect 492 379 495 383
rect 603 379 604 383
rect 604 379 607 383
rect 771 379 775 383
rect 839 379 843 383
rect 931 379 932 383
rect 932 379 935 383
rect 1167 379 1171 383
rect 1219 379 1220 383
rect 1220 379 1223 383
rect 631 371 635 375
rect 1623 375 1627 379
rect 1703 375 1707 379
rect 1759 375 1763 379
rect 1823 375 1827 379
rect 1879 375 1883 379
rect 251 363 255 367
rect 359 363 363 367
rect 463 363 467 367
rect 663 363 667 367
rect 671 363 675 367
rect 871 363 875 367
rect 995 363 996 367
rect 996 363 999 367
rect 1075 363 1076 367
rect 1076 363 1079 367
rect 1119 363 1123 367
rect 1199 363 1203 367
rect 1887 363 1891 367
rect 2103 375 2107 379
rect 2295 375 2299 379
rect 2391 375 2395 379
rect 2475 375 2479 379
rect 2447 363 2451 367
rect 1327 356 1331 360
rect 1679 357 1683 361
rect 1703 355 1704 359
rect 1704 355 1707 359
rect 1735 357 1739 361
rect 1759 355 1760 359
rect 1760 355 1763 359
rect 1799 357 1803 361
rect 1823 355 1824 359
rect 1824 355 1827 359
rect 1871 357 1875 361
rect 1895 355 1896 359
rect 1896 355 1899 359
rect 1943 357 1947 361
rect 1963 355 1964 359
rect 1964 355 1967 359
rect 2023 357 2027 361
rect 2111 357 2115 361
rect 2199 357 2203 361
rect 2207 355 2211 359
rect 2287 357 2291 361
rect 2375 357 2379 361
rect 2383 355 2387 359
rect 2455 357 2459 361
rect 2503 356 2507 360
rect 111 344 115 348
rect 151 345 155 349
rect 171 343 172 347
rect 172 343 175 347
rect 231 345 235 349
rect 335 345 339 349
rect 359 343 360 347
rect 360 343 363 347
rect 439 345 443 349
rect 463 343 464 347
rect 464 343 467 347
rect 543 345 547 349
rect 559 343 563 347
rect 647 345 651 349
rect 671 343 672 347
rect 672 343 675 347
rect 751 345 755 349
rect 771 343 772 347
rect 772 343 775 347
rect 847 345 851 349
rect 871 343 872 347
rect 872 343 875 347
rect 935 345 939 349
rect 951 343 955 347
rect 1015 345 1019 349
rect 1095 345 1099 349
rect 1119 343 1120 347
rect 1120 343 1123 347
rect 1175 345 1179 349
rect 1199 343 1200 347
rect 1200 343 1203 347
rect 1239 345 1243 349
rect 1247 343 1251 347
rect 1287 344 1291 348
rect 1327 339 1331 343
rect 1663 336 1667 340
rect 1719 336 1723 340
rect 1783 336 1787 340
rect 1855 336 1859 340
rect 1927 336 1931 340
rect 2007 336 2011 340
rect 2095 336 2099 340
rect 2183 336 2187 340
rect 2271 336 2275 340
rect 2359 336 2363 340
rect 2439 336 2443 340
rect 2503 339 2507 343
rect 111 327 115 331
rect 135 324 139 328
rect 215 324 219 328
rect 319 324 323 328
rect 423 324 427 328
rect 527 324 531 328
rect 631 324 635 328
rect 735 324 739 328
rect 831 324 835 328
rect 919 324 923 328
rect 999 324 1003 328
rect 1079 324 1083 328
rect 1159 324 1163 328
rect 1223 324 1227 328
rect 1287 327 1291 331
rect 1327 313 1331 317
rect 1351 316 1355 320
rect 1455 316 1459 320
rect 1583 316 1587 320
rect 1711 316 1715 320
rect 1839 316 1843 320
rect 1951 316 1955 320
rect 2063 316 2067 320
rect 2167 316 2171 320
rect 2263 316 2267 320
rect 2359 316 2363 320
rect 2439 316 2443 320
rect 111 305 115 309
rect 135 308 139 312
rect 215 308 219 312
rect 319 308 323 312
rect 423 308 427 312
rect 535 308 539 312
rect 639 308 643 312
rect 743 308 747 312
rect 847 308 851 312
rect 943 308 947 312
rect 1039 308 1043 312
rect 1143 308 1147 312
rect 2503 313 2507 317
rect 1223 308 1227 312
rect 1287 305 1291 309
rect 1327 296 1331 300
rect 1367 295 1371 299
rect 1375 295 1379 299
rect 1471 295 1475 299
rect 1579 295 1583 299
rect 1599 295 1603 299
rect 1623 295 1624 299
rect 1624 295 1627 299
rect 1727 295 1731 299
rect 111 288 115 292
rect 151 287 155 291
rect 211 287 215 291
rect 231 287 235 291
rect 251 287 252 291
rect 252 287 255 291
rect 335 287 339 291
rect 403 287 407 291
rect 439 287 443 291
rect 551 287 555 291
rect 655 287 659 291
rect 663 287 667 291
rect 759 287 763 291
rect 863 287 867 291
rect 959 287 963 291
rect 1035 287 1039 291
rect 1055 287 1059 291
rect 1139 287 1143 291
rect 1159 287 1163 291
rect 1203 287 1207 291
rect 1239 287 1243 291
rect 1287 288 1291 292
rect 1855 295 1859 299
rect 1879 295 1880 299
rect 1880 295 1883 299
rect 1967 295 1971 299
rect 2079 295 2083 299
rect 2087 295 2091 299
rect 2183 295 2187 299
rect 2279 295 2283 299
rect 2355 295 2359 299
rect 2375 295 2379 299
rect 2455 295 2459 299
rect 2475 295 2476 299
rect 2476 295 2479 299
rect 2503 296 2507 300
rect 1579 275 1580 279
rect 1580 275 1583 279
rect 1779 275 1783 279
rect 1987 275 1991 279
rect 2207 275 2211 279
rect 2383 275 2387 279
rect 2463 275 2467 279
rect 171 267 175 271
rect 211 267 212 271
rect 212 267 215 271
rect 559 267 563 271
rect 891 267 895 271
rect 951 267 955 271
rect 1035 267 1036 271
rect 1036 267 1039 271
rect 1139 267 1140 271
rect 1140 267 1143 271
rect 1247 267 1251 271
rect 311 255 315 259
rect 403 255 404 259
rect 404 255 407 259
rect 447 255 451 259
rect 559 255 563 259
rect 735 255 739 259
rect 783 255 787 259
rect 1203 255 1204 259
rect 1204 255 1207 259
rect 1375 255 1379 259
rect 1391 255 1395 259
rect 1575 255 1579 259
rect 1679 255 1683 259
rect 1839 255 1843 259
rect 1887 255 1891 259
rect 2087 255 2091 259
rect 2095 255 2099 259
rect 2199 255 2203 259
rect 2355 255 2356 259
rect 2356 255 2359 259
rect 2399 255 2403 259
rect 1587 247 1591 251
rect 111 236 115 240
rect 151 237 155 241
rect 171 235 172 239
rect 172 235 175 239
rect 223 237 227 241
rect 319 237 323 241
rect 423 237 427 241
rect 447 235 448 239
rect 448 235 451 239
rect 535 237 539 241
rect 559 235 560 239
rect 560 235 563 239
rect 647 237 651 241
rect 655 235 659 239
rect 759 237 763 241
rect 783 235 784 239
rect 784 235 787 239
rect 871 237 875 241
rect 891 235 892 239
rect 892 235 895 239
rect 983 237 987 241
rect 991 235 995 239
rect 1103 237 1107 241
rect 1223 237 1227 241
rect 1287 236 1291 240
rect 1327 236 1331 240
rect 1367 237 1371 241
rect 1391 235 1392 239
rect 1392 235 1395 239
rect 1447 237 1451 241
rect 1463 235 1467 239
rect 1551 237 1555 241
rect 1575 235 1576 239
rect 1576 235 1579 239
rect 1655 237 1659 241
rect 1679 235 1680 239
rect 1680 235 1683 239
rect 1759 237 1763 241
rect 1779 235 1780 239
rect 1780 235 1783 239
rect 1863 237 1867 241
rect 1887 235 1888 239
rect 1888 235 1891 239
rect 1967 237 1971 241
rect 1987 235 1988 239
rect 1988 235 1991 239
rect 2071 237 2075 241
rect 2095 235 2096 239
rect 2096 235 2099 239
rect 2175 237 2179 241
rect 2199 235 2200 239
rect 2200 235 2203 239
rect 2271 237 2275 241
rect 2327 235 2331 239
rect 2375 237 2379 241
rect 2399 235 2400 239
rect 2400 235 2403 239
rect 2455 237 2459 241
rect 2471 235 2475 239
rect 2503 236 2507 240
rect 111 219 115 223
rect 135 216 139 220
rect 207 216 211 220
rect 303 216 307 220
rect 407 216 411 220
rect 519 216 523 220
rect 631 216 635 220
rect 743 216 747 220
rect 855 216 859 220
rect 967 216 971 220
rect 1087 216 1091 220
rect 1207 216 1211 220
rect 1287 219 1291 223
rect 1327 219 1331 223
rect 1351 216 1355 220
rect 1431 216 1435 220
rect 1535 216 1539 220
rect 1639 216 1643 220
rect 1743 216 1747 220
rect 1847 216 1851 220
rect 1951 216 1955 220
rect 2055 216 2059 220
rect 2159 216 2163 220
rect 2255 216 2259 220
rect 2359 216 2363 220
rect 2439 216 2443 220
rect 2503 219 2507 223
rect 111 197 115 201
rect 183 200 187 204
rect 279 200 283 204
rect 383 200 387 204
rect 487 200 491 204
rect 591 200 595 204
rect 695 200 699 204
rect 799 200 803 204
rect 895 200 899 204
rect 999 200 1003 204
rect 1103 200 1107 204
rect 1287 197 1291 201
rect 1327 197 1331 201
rect 1351 200 1355 204
rect 1407 200 1411 204
rect 1471 200 1475 204
rect 1551 200 1555 204
rect 1639 200 1643 204
rect 1719 200 1723 204
rect 1807 200 1811 204
rect 1895 200 1899 204
rect 1991 200 1995 204
rect 2103 200 2107 204
rect 2215 200 2219 204
rect 2335 200 2339 204
rect 2439 200 2443 204
rect 2503 197 2507 201
rect 111 180 115 184
rect 199 179 203 183
rect 275 179 279 183
rect 295 179 299 183
rect 311 179 315 183
rect 399 179 403 183
rect 467 179 471 183
rect 503 179 507 183
rect 607 179 611 183
rect 711 179 715 183
rect 735 179 736 183
rect 736 179 739 183
rect 815 179 819 183
rect 911 179 915 183
rect 995 179 999 183
rect 1015 179 1019 183
rect 1099 179 1103 183
rect 1119 179 1123 183
rect 1135 179 1139 183
rect 1287 180 1291 184
rect 1327 180 1331 184
rect 1367 179 1371 183
rect 1375 179 1379 183
rect 1423 179 1427 183
rect 1487 179 1491 183
rect 1567 179 1571 183
rect 1587 179 1588 183
rect 1588 179 1591 183
rect 1655 179 1659 183
rect 1735 179 1739 183
rect 1823 179 1827 183
rect 1839 179 1843 183
rect 1911 179 1915 183
rect 2007 179 2011 183
rect 2119 179 2123 183
rect 2127 179 2131 183
rect 2231 179 2235 183
rect 2351 179 2355 183
rect 2455 179 2459 183
rect 2463 179 2467 183
rect 2503 180 2507 184
rect 227 159 231 163
rect 275 159 276 163
rect 276 159 279 163
rect 655 159 659 163
rect 791 159 795 163
rect 987 159 991 163
rect 995 159 996 163
rect 996 159 999 163
rect 1099 159 1100 163
rect 1100 159 1103 163
rect 1463 159 1467 163
rect 1779 159 1783 163
rect 1967 159 1971 163
rect 2327 159 2331 163
rect 2471 159 2475 163
rect 175 139 179 143
rect 467 139 468 143
rect 468 139 471 143
rect 511 139 515 143
rect 567 139 571 143
rect 679 139 683 143
rect 735 139 739 143
rect 1135 139 1136 143
rect 1136 139 1139 143
rect 1375 127 1379 131
rect 1391 127 1395 131
rect 1447 127 1451 131
rect 1503 127 1507 131
rect 1559 127 1563 131
rect 1615 127 1619 131
rect 1671 127 1675 131
rect 1727 127 1731 131
rect 111 120 115 124
rect 151 121 155 125
rect 175 119 176 123
rect 176 119 179 123
rect 207 121 211 125
rect 227 119 228 123
rect 228 119 231 123
rect 263 121 267 125
rect 319 121 323 125
rect 375 121 379 125
rect 431 121 435 125
rect 487 121 491 125
rect 511 119 512 123
rect 512 119 515 123
rect 543 121 547 125
rect 567 119 568 123
rect 568 119 571 123
rect 599 121 603 125
rect 655 121 659 125
rect 679 119 680 123
rect 680 119 683 123
rect 711 121 715 125
rect 735 119 736 123
rect 736 119 739 123
rect 767 121 771 125
rect 791 119 792 123
rect 792 119 795 123
rect 831 121 835 125
rect 895 121 899 125
rect 959 121 963 125
rect 1023 121 1027 125
rect 1087 121 1091 125
rect 1151 121 1155 125
rect 1287 120 1291 124
rect 1847 127 1851 131
rect 1903 127 1907 131
rect 2127 127 2128 131
rect 2128 127 2131 131
rect 2167 127 2171 131
rect 2247 127 2251 131
rect 2463 127 2467 131
rect 1327 108 1331 112
rect 1367 109 1371 113
rect 111 103 115 107
rect 1391 107 1392 111
rect 1392 107 1395 111
rect 1423 109 1427 113
rect 135 100 139 104
rect 191 100 195 104
rect 247 100 251 104
rect 303 100 307 104
rect 359 100 363 104
rect 415 100 419 104
rect 471 100 475 104
rect 527 100 531 104
rect 583 100 587 104
rect 639 100 643 104
rect 695 100 699 104
rect 751 100 755 104
rect 815 100 819 104
rect 879 100 883 104
rect 943 100 947 104
rect 1007 100 1011 104
rect 1071 100 1075 104
rect 1135 100 1139 104
rect 1287 103 1291 107
rect 1447 107 1448 111
rect 1448 107 1451 111
rect 1479 109 1483 113
rect 1503 107 1504 111
rect 1504 107 1507 111
rect 1535 109 1539 113
rect 1559 107 1560 111
rect 1560 107 1563 111
rect 1591 109 1595 113
rect 1615 107 1616 111
rect 1616 107 1619 111
rect 1647 109 1651 113
rect 1671 107 1672 111
rect 1672 107 1675 111
rect 1703 109 1707 113
rect 1727 107 1728 111
rect 1728 107 1731 111
rect 1759 109 1763 113
rect 1779 107 1780 111
rect 1780 107 1783 111
rect 1823 109 1827 113
rect 1847 107 1848 111
rect 1848 107 1851 111
rect 1879 109 1883 113
rect 1903 107 1904 111
rect 1904 107 1907 111
rect 1943 109 1947 113
rect 1967 107 1968 111
rect 1968 107 1971 111
rect 2007 109 2011 113
rect 2071 109 2075 113
rect 2143 109 2147 113
rect 2167 107 2168 111
rect 2168 107 2171 111
rect 2223 109 2227 113
rect 2247 107 2248 111
rect 2248 107 2251 111
rect 2303 109 2307 113
rect 2391 109 2395 113
rect 2455 109 2459 113
rect 2503 108 2507 112
rect 1327 91 1331 95
rect 1351 88 1355 92
rect 1407 88 1411 92
rect 1463 88 1467 92
rect 1519 88 1523 92
rect 1575 88 1579 92
rect 1631 88 1635 92
rect 1687 88 1691 92
rect 1743 88 1747 92
rect 1807 88 1811 92
rect 1863 88 1867 92
rect 1927 88 1931 92
rect 1991 88 1995 92
rect 2055 88 2059 92
rect 2127 88 2131 92
rect 2207 88 2211 92
rect 2287 88 2291 92
rect 2375 88 2379 92
rect 2439 88 2443 92
rect 2503 91 2507 95
<< m3 >>
rect 111 2582 115 2583
rect 111 2577 115 2578
rect 135 2582 139 2583
rect 135 2577 139 2578
rect 191 2582 195 2583
rect 191 2577 195 2578
rect 247 2582 251 2583
rect 247 2577 251 2578
rect 303 2582 307 2583
rect 303 2577 307 2578
rect 359 2582 363 2583
rect 359 2577 363 2578
rect 1287 2582 1291 2583
rect 1287 2577 1291 2578
rect 112 2574 114 2577
rect 134 2576 140 2577
rect 110 2573 116 2574
rect 110 2569 111 2573
rect 115 2569 116 2573
rect 134 2572 135 2576
rect 139 2572 140 2576
rect 134 2571 140 2572
rect 190 2576 196 2577
rect 190 2572 191 2576
rect 195 2572 196 2576
rect 190 2571 196 2572
rect 246 2576 252 2577
rect 246 2572 247 2576
rect 251 2572 252 2576
rect 246 2571 252 2572
rect 302 2576 308 2577
rect 302 2572 303 2576
rect 307 2572 308 2576
rect 302 2571 308 2572
rect 358 2576 364 2577
rect 358 2572 359 2576
rect 363 2572 364 2576
rect 1288 2574 1290 2577
rect 358 2571 364 2572
rect 1286 2573 1292 2574
rect 110 2568 116 2569
rect 1286 2569 1287 2573
rect 1291 2569 1292 2573
rect 1286 2568 1292 2569
rect 1327 2562 1331 2563
rect 1327 2557 1331 2558
rect 1495 2562 1499 2563
rect 1495 2557 1499 2558
rect 1551 2562 1555 2563
rect 1551 2557 1555 2558
rect 1607 2562 1611 2563
rect 1607 2557 1611 2558
rect 1663 2562 1667 2563
rect 1663 2557 1667 2558
rect 1719 2562 1723 2563
rect 1719 2557 1723 2558
rect 1775 2562 1779 2563
rect 1775 2557 1779 2558
rect 1831 2562 1835 2563
rect 1831 2557 1835 2558
rect 1887 2562 1891 2563
rect 1887 2557 1891 2558
rect 1943 2562 1947 2563
rect 1943 2557 1947 2558
rect 1999 2562 2003 2563
rect 1999 2557 2003 2558
rect 2055 2562 2059 2563
rect 2055 2557 2059 2558
rect 2111 2562 2115 2563
rect 2111 2557 2115 2558
rect 2167 2562 2171 2563
rect 2167 2557 2171 2558
rect 2503 2562 2507 2563
rect 2503 2557 2507 2558
rect 110 2556 116 2557
rect 1286 2556 1292 2557
rect 110 2552 111 2556
rect 115 2552 116 2556
rect 110 2551 116 2552
rect 150 2555 156 2556
rect 150 2551 151 2555
rect 155 2551 156 2555
rect 112 2531 114 2551
rect 150 2550 156 2551
rect 186 2555 192 2556
rect 186 2551 187 2555
rect 191 2551 192 2555
rect 186 2550 192 2551
rect 206 2555 212 2556
rect 206 2551 207 2555
rect 211 2551 212 2555
rect 206 2550 212 2551
rect 242 2555 248 2556
rect 242 2551 243 2555
rect 247 2551 248 2555
rect 242 2550 248 2551
rect 262 2555 268 2556
rect 262 2551 263 2555
rect 267 2551 268 2555
rect 262 2550 268 2551
rect 298 2555 304 2556
rect 298 2551 299 2555
rect 303 2551 304 2555
rect 298 2550 304 2551
rect 318 2555 324 2556
rect 318 2551 319 2555
rect 323 2551 324 2555
rect 318 2550 324 2551
rect 354 2555 360 2556
rect 354 2551 355 2555
rect 359 2551 360 2555
rect 354 2550 360 2551
rect 374 2555 380 2556
rect 374 2551 375 2555
rect 379 2551 380 2555
rect 1286 2552 1287 2556
rect 1291 2552 1292 2556
rect 1328 2554 1330 2557
rect 1494 2556 1500 2557
rect 1286 2551 1292 2552
rect 1326 2553 1332 2554
rect 374 2550 380 2551
rect 152 2531 154 2550
rect 188 2536 190 2550
rect 186 2535 192 2536
rect 186 2531 187 2535
rect 191 2531 192 2535
rect 208 2531 210 2550
rect 214 2547 220 2548
rect 214 2543 215 2547
rect 219 2543 220 2547
rect 214 2542 220 2543
rect 111 2530 115 2531
rect 111 2525 115 2526
rect 151 2530 155 2531
rect 186 2530 192 2531
rect 207 2530 211 2531
rect 151 2525 155 2526
rect 207 2525 211 2526
rect 112 2505 114 2525
rect 216 2524 218 2542
rect 244 2536 246 2550
rect 242 2535 248 2536
rect 242 2531 243 2535
rect 247 2531 248 2535
rect 264 2531 266 2550
rect 300 2536 302 2550
rect 298 2535 304 2536
rect 298 2531 299 2535
rect 303 2531 304 2535
rect 320 2531 322 2550
rect 356 2536 358 2550
rect 354 2535 360 2536
rect 354 2531 355 2535
rect 359 2531 360 2535
rect 376 2531 378 2550
rect 1288 2531 1290 2551
rect 1326 2549 1327 2553
rect 1331 2549 1332 2553
rect 1494 2552 1495 2556
rect 1499 2552 1500 2556
rect 1494 2551 1500 2552
rect 1550 2556 1556 2557
rect 1550 2552 1551 2556
rect 1555 2552 1556 2556
rect 1550 2551 1556 2552
rect 1606 2556 1612 2557
rect 1606 2552 1607 2556
rect 1611 2552 1612 2556
rect 1606 2551 1612 2552
rect 1662 2556 1668 2557
rect 1662 2552 1663 2556
rect 1667 2552 1668 2556
rect 1662 2551 1668 2552
rect 1718 2556 1724 2557
rect 1718 2552 1719 2556
rect 1723 2552 1724 2556
rect 1718 2551 1724 2552
rect 1774 2556 1780 2557
rect 1774 2552 1775 2556
rect 1779 2552 1780 2556
rect 1774 2551 1780 2552
rect 1830 2556 1836 2557
rect 1830 2552 1831 2556
rect 1835 2552 1836 2556
rect 1830 2551 1836 2552
rect 1886 2556 1892 2557
rect 1886 2552 1887 2556
rect 1891 2552 1892 2556
rect 1886 2551 1892 2552
rect 1942 2556 1948 2557
rect 1942 2552 1943 2556
rect 1947 2552 1948 2556
rect 1942 2551 1948 2552
rect 1998 2556 2004 2557
rect 1998 2552 1999 2556
rect 2003 2552 2004 2556
rect 1998 2551 2004 2552
rect 2054 2556 2060 2557
rect 2054 2552 2055 2556
rect 2059 2552 2060 2556
rect 2054 2551 2060 2552
rect 2110 2556 2116 2557
rect 2110 2552 2111 2556
rect 2115 2552 2116 2556
rect 2110 2551 2116 2552
rect 2166 2556 2172 2557
rect 2166 2552 2167 2556
rect 2171 2552 2172 2556
rect 2504 2554 2506 2557
rect 2166 2551 2172 2552
rect 2502 2553 2508 2554
rect 1326 2548 1332 2549
rect 2502 2549 2503 2553
rect 2507 2549 2508 2553
rect 2502 2548 2508 2549
rect 1326 2536 1332 2537
rect 2502 2536 2508 2537
rect 1326 2532 1327 2536
rect 1331 2532 1332 2536
rect 1326 2531 1332 2532
rect 1510 2535 1516 2536
rect 1510 2531 1511 2535
rect 1515 2531 1516 2535
rect 223 2530 227 2531
rect 242 2530 248 2531
rect 263 2530 267 2531
rect 223 2525 227 2526
rect 263 2525 267 2526
rect 279 2530 283 2531
rect 298 2530 304 2531
rect 319 2530 323 2531
rect 279 2525 283 2526
rect 319 2525 323 2526
rect 343 2530 347 2531
rect 354 2530 360 2531
rect 375 2530 379 2531
rect 343 2525 347 2526
rect 375 2525 379 2526
rect 415 2530 419 2531
rect 415 2525 419 2526
rect 487 2530 491 2531
rect 487 2525 491 2526
rect 551 2530 555 2531
rect 551 2525 555 2526
rect 615 2530 619 2531
rect 615 2525 619 2526
rect 679 2530 683 2531
rect 679 2525 683 2526
rect 743 2530 747 2531
rect 743 2525 747 2526
rect 807 2530 811 2531
rect 807 2525 811 2526
rect 871 2530 875 2531
rect 871 2525 875 2526
rect 935 2530 939 2531
rect 935 2525 939 2526
rect 999 2530 1003 2531
rect 999 2525 1003 2526
rect 1063 2530 1067 2531
rect 1063 2525 1067 2526
rect 1287 2530 1291 2531
rect 1287 2525 1291 2526
rect 214 2523 220 2524
rect 214 2519 215 2523
rect 219 2519 220 2523
rect 214 2518 220 2519
rect 224 2506 226 2525
rect 246 2523 252 2524
rect 246 2519 247 2523
rect 251 2519 252 2523
rect 246 2518 252 2519
rect 222 2505 228 2506
rect 110 2504 116 2505
rect 110 2500 111 2504
rect 115 2500 116 2504
rect 222 2501 223 2505
rect 227 2501 228 2505
rect 248 2504 250 2518
rect 280 2506 282 2525
rect 302 2523 308 2524
rect 302 2519 303 2523
rect 307 2519 308 2523
rect 302 2518 308 2519
rect 278 2505 284 2506
rect 222 2500 228 2501
rect 246 2503 252 2504
rect 110 2499 116 2500
rect 246 2499 247 2503
rect 251 2499 252 2503
rect 278 2501 279 2505
rect 283 2501 284 2505
rect 304 2504 306 2518
rect 344 2506 346 2525
rect 366 2523 372 2524
rect 366 2519 367 2523
rect 371 2519 372 2523
rect 366 2518 372 2519
rect 342 2505 348 2506
rect 278 2500 284 2501
rect 302 2503 308 2504
rect 246 2498 252 2499
rect 302 2499 303 2503
rect 307 2499 308 2503
rect 342 2501 343 2505
rect 347 2501 348 2505
rect 368 2504 370 2518
rect 416 2506 418 2525
rect 438 2523 444 2524
rect 438 2519 439 2523
rect 443 2519 444 2523
rect 438 2518 444 2519
rect 414 2505 420 2506
rect 342 2500 348 2501
rect 366 2503 372 2504
rect 302 2498 308 2499
rect 366 2499 367 2503
rect 371 2499 372 2503
rect 414 2501 415 2505
rect 419 2501 420 2505
rect 440 2504 442 2518
rect 488 2506 490 2525
rect 552 2506 554 2525
rect 566 2523 572 2524
rect 566 2519 567 2523
rect 571 2519 572 2523
rect 566 2518 572 2519
rect 574 2523 580 2524
rect 574 2519 575 2523
rect 579 2519 580 2523
rect 574 2518 580 2519
rect 486 2505 492 2506
rect 414 2500 420 2501
rect 438 2503 444 2504
rect 366 2498 372 2499
rect 438 2499 439 2503
rect 443 2499 444 2503
rect 486 2501 487 2505
rect 491 2501 492 2505
rect 550 2505 556 2506
rect 486 2500 492 2501
rect 494 2503 500 2504
rect 438 2498 444 2499
rect 494 2499 495 2503
rect 499 2499 500 2503
rect 550 2501 551 2505
rect 555 2501 556 2505
rect 550 2500 556 2501
rect 494 2498 500 2499
rect 110 2487 116 2488
rect 110 2483 111 2487
rect 115 2483 116 2487
rect 110 2482 116 2483
rect 206 2484 212 2485
rect 112 2471 114 2482
rect 206 2480 207 2484
rect 211 2480 212 2484
rect 206 2479 212 2480
rect 262 2484 268 2485
rect 262 2480 263 2484
rect 267 2480 268 2484
rect 262 2479 268 2480
rect 326 2484 332 2485
rect 326 2480 327 2484
rect 331 2480 332 2484
rect 326 2479 332 2480
rect 398 2484 404 2485
rect 398 2480 399 2484
rect 403 2480 404 2484
rect 398 2479 404 2480
rect 470 2484 476 2485
rect 470 2480 471 2484
rect 475 2480 476 2484
rect 470 2479 476 2480
rect 208 2471 210 2479
rect 264 2471 266 2479
rect 328 2471 330 2479
rect 400 2471 402 2479
rect 472 2471 474 2479
rect 111 2470 115 2471
rect 111 2465 115 2466
rect 167 2470 171 2471
rect 167 2465 171 2466
rect 207 2470 211 2471
rect 207 2465 211 2466
rect 223 2470 227 2471
rect 223 2465 227 2466
rect 263 2470 267 2471
rect 263 2465 267 2466
rect 279 2470 283 2471
rect 279 2465 283 2466
rect 327 2470 331 2471
rect 327 2465 331 2466
rect 335 2470 339 2471
rect 335 2465 339 2466
rect 391 2470 395 2471
rect 391 2465 395 2466
rect 399 2470 403 2471
rect 399 2465 403 2466
rect 447 2470 451 2471
rect 447 2465 451 2466
rect 471 2470 475 2471
rect 471 2465 475 2466
rect 112 2462 114 2465
rect 166 2464 172 2465
rect 110 2461 116 2462
rect 110 2457 111 2461
rect 115 2457 116 2461
rect 166 2460 167 2464
rect 171 2460 172 2464
rect 166 2459 172 2460
rect 222 2464 228 2465
rect 222 2460 223 2464
rect 227 2460 228 2464
rect 222 2459 228 2460
rect 278 2464 284 2465
rect 278 2460 279 2464
rect 283 2460 284 2464
rect 278 2459 284 2460
rect 334 2464 340 2465
rect 334 2460 335 2464
rect 339 2460 340 2464
rect 334 2459 340 2460
rect 390 2464 396 2465
rect 390 2460 391 2464
rect 395 2460 396 2464
rect 390 2459 396 2460
rect 446 2464 452 2465
rect 446 2460 447 2464
rect 451 2460 452 2464
rect 446 2459 452 2460
rect 110 2456 116 2457
rect 496 2453 498 2498
rect 534 2484 540 2485
rect 534 2480 535 2484
rect 539 2480 540 2484
rect 534 2479 540 2480
rect 536 2471 538 2479
rect 503 2470 507 2471
rect 503 2465 507 2466
rect 535 2470 539 2471
rect 535 2465 539 2466
rect 559 2470 563 2471
rect 559 2465 563 2466
rect 502 2464 508 2465
rect 502 2460 503 2464
rect 507 2460 508 2464
rect 502 2459 508 2460
rect 558 2464 564 2465
rect 558 2460 559 2464
rect 563 2460 564 2464
rect 558 2459 564 2460
rect 568 2453 570 2518
rect 576 2504 578 2518
rect 616 2506 618 2525
rect 638 2523 644 2524
rect 638 2519 639 2523
rect 643 2519 644 2523
rect 638 2518 644 2519
rect 614 2505 620 2506
rect 574 2503 580 2504
rect 574 2499 575 2503
rect 579 2499 580 2503
rect 614 2501 615 2505
rect 619 2501 620 2505
rect 640 2504 642 2518
rect 680 2506 682 2525
rect 702 2523 708 2524
rect 702 2519 703 2523
rect 707 2519 708 2523
rect 702 2518 708 2519
rect 678 2505 684 2506
rect 614 2500 620 2501
rect 638 2503 644 2504
rect 574 2498 580 2499
rect 638 2499 639 2503
rect 643 2499 644 2503
rect 678 2501 679 2505
rect 683 2501 684 2505
rect 704 2504 706 2518
rect 744 2506 746 2525
rect 762 2523 768 2524
rect 762 2519 763 2523
rect 767 2519 768 2523
rect 762 2518 768 2519
rect 742 2505 748 2506
rect 678 2500 684 2501
rect 702 2503 708 2504
rect 638 2498 644 2499
rect 702 2499 703 2503
rect 707 2499 708 2503
rect 742 2501 743 2505
rect 747 2501 748 2505
rect 764 2504 766 2518
rect 808 2506 810 2525
rect 826 2523 832 2524
rect 826 2519 827 2523
rect 831 2519 832 2523
rect 826 2518 832 2519
rect 806 2505 812 2506
rect 742 2500 748 2501
rect 762 2503 768 2504
rect 702 2498 708 2499
rect 762 2499 763 2503
rect 767 2499 768 2503
rect 806 2501 807 2505
rect 811 2501 812 2505
rect 828 2504 830 2518
rect 872 2506 874 2525
rect 890 2523 896 2524
rect 890 2519 891 2523
rect 895 2519 896 2523
rect 890 2518 896 2519
rect 870 2505 876 2506
rect 806 2500 812 2501
rect 826 2503 832 2504
rect 762 2498 768 2499
rect 826 2499 827 2503
rect 831 2499 832 2503
rect 870 2501 871 2505
rect 875 2501 876 2505
rect 892 2504 894 2518
rect 936 2506 938 2525
rect 958 2523 964 2524
rect 958 2519 959 2523
rect 963 2519 964 2523
rect 958 2518 964 2519
rect 934 2505 940 2506
rect 870 2500 876 2501
rect 890 2503 896 2504
rect 826 2498 832 2499
rect 890 2499 891 2503
rect 895 2499 896 2503
rect 934 2501 935 2505
rect 939 2501 940 2505
rect 960 2504 962 2518
rect 1000 2506 1002 2525
rect 1018 2523 1024 2524
rect 1018 2519 1019 2523
rect 1023 2519 1024 2523
rect 1018 2518 1024 2519
rect 998 2505 1004 2506
rect 934 2500 940 2501
rect 958 2503 964 2504
rect 890 2498 896 2499
rect 958 2499 959 2503
rect 963 2499 964 2503
rect 998 2501 999 2505
rect 1003 2501 1004 2505
rect 1020 2504 1022 2518
rect 1064 2506 1066 2525
rect 1062 2505 1068 2506
rect 1288 2505 1290 2525
rect 1328 2511 1330 2531
rect 1510 2530 1516 2531
rect 1534 2535 1540 2536
rect 1534 2531 1535 2535
rect 1539 2531 1540 2535
rect 1534 2530 1540 2531
rect 1566 2535 1572 2536
rect 1566 2531 1567 2535
rect 1571 2531 1572 2535
rect 1566 2530 1572 2531
rect 1598 2535 1604 2536
rect 1598 2531 1599 2535
rect 1603 2531 1604 2535
rect 1598 2530 1604 2531
rect 1622 2535 1628 2536
rect 1622 2531 1623 2535
rect 1627 2531 1628 2535
rect 1622 2530 1628 2531
rect 1658 2535 1664 2536
rect 1658 2531 1659 2535
rect 1663 2531 1664 2535
rect 1658 2530 1664 2531
rect 1678 2535 1684 2536
rect 1678 2531 1679 2535
rect 1683 2531 1684 2535
rect 1678 2530 1684 2531
rect 1714 2535 1720 2536
rect 1714 2531 1715 2535
rect 1719 2531 1720 2535
rect 1714 2530 1720 2531
rect 1734 2535 1740 2536
rect 1734 2531 1735 2535
rect 1739 2531 1740 2535
rect 1734 2530 1740 2531
rect 1770 2535 1776 2536
rect 1770 2531 1771 2535
rect 1775 2531 1776 2535
rect 1770 2530 1776 2531
rect 1790 2535 1796 2536
rect 1790 2531 1791 2535
rect 1795 2531 1796 2535
rect 1790 2530 1796 2531
rect 1814 2535 1820 2536
rect 1814 2531 1815 2535
rect 1819 2531 1820 2535
rect 1814 2530 1820 2531
rect 1846 2535 1852 2536
rect 1846 2531 1847 2535
rect 1851 2531 1852 2535
rect 1846 2530 1852 2531
rect 1882 2535 1888 2536
rect 1882 2531 1883 2535
rect 1887 2531 1888 2535
rect 1882 2530 1888 2531
rect 1902 2535 1908 2536
rect 1902 2531 1903 2535
rect 1907 2531 1908 2535
rect 1902 2530 1908 2531
rect 1938 2535 1944 2536
rect 1938 2531 1939 2535
rect 1943 2531 1944 2535
rect 1938 2530 1944 2531
rect 1958 2535 1964 2536
rect 1958 2531 1959 2535
rect 1963 2531 1964 2535
rect 1958 2530 1964 2531
rect 1994 2535 2000 2536
rect 1994 2531 1995 2535
rect 1999 2531 2000 2535
rect 1994 2530 2000 2531
rect 2014 2535 2020 2536
rect 2014 2531 2015 2535
rect 2019 2531 2020 2535
rect 2014 2530 2020 2531
rect 2050 2535 2056 2536
rect 2050 2531 2051 2535
rect 2055 2531 2056 2535
rect 2050 2530 2056 2531
rect 2070 2535 2076 2536
rect 2070 2531 2071 2535
rect 2075 2531 2076 2535
rect 2070 2530 2076 2531
rect 2102 2535 2108 2536
rect 2102 2531 2103 2535
rect 2107 2531 2108 2535
rect 2102 2530 2108 2531
rect 2126 2535 2132 2536
rect 2126 2531 2127 2535
rect 2131 2531 2132 2535
rect 2126 2530 2132 2531
rect 2162 2535 2168 2536
rect 2162 2531 2163 2535
rect 2167 2531 2168 2535
rect 2162 2530 2168 2531
rect 2182 2535 2188 2536
rect 2182 2531 2183 2535
rect 2187 2531 2188 2535
rect 2182 2530 2188 2531
rect 2190 2535 2196 2536
rect 2190 2531 2191 2535
rect 2195 2531 2196 2535
rect 2502 2532 2503 2536
rect 2507 2532 2508 2536
rect 2502 2531 2508 2532
rect 2190 2530 2196 2531
rect 1512 2511 1514 2530
rect 1536 2516 1538 2530
rect 1526 2515 1532 2516
rect 1526 2511 1527 2515
rect 1531 2511 1532 2515
rect 1327 2510 1331 2511
rect 1327 2505 1331 2506
rect 1511 2510 1515 2511
rect 1526 2510 1532 2511
rect 1534 2515 1540 2516
rect 1534 2511 1535 2515
rect 1539 2511 1540 2515
rect 1568 2511 1570 2530
rect 1600 2516 1602 2530
rect 1598 2515 1604 2516
rect 1598 2511 1599 2515
rect 1603 2511 1604 2515
rect 1624 2511 1626 2530
rect 1660 2516 1662 2530
rect 1658 2515 1664 2516
rect 1658 2511 1659 2515
rect 1663 2511 1664 2515
rect 1680 2511 1682 2530
rect 1716 2516 1718 2530
rect 1714 2515 1720 2516
rect 1714 2511 1715 2515
rect 1719 2511 1720 2515
rect 1736 2511 1738 2530
rect 1772 2516 1774 2530
rect 1770 2515 1776 2516
rect 1770 2511 1771 2515
rect 1775 2511 1776 2515
rect 1792 2511 1794 2530
rect 1816 2516 1818 2530
rect 1814 2515 1820 2516
rect 1814 2511 1815 2515
rect 1819 2511 1820 2515
rect 1848 2511 1850 2530
rect 1884 2516 1886 2530
rect 1882 2515 1888 2516
rect 1882 2511 1883 2515
rect 1887 2511 1888 2515
rect 1904 2511 1906 2530
rect 1911 2524 1915 2525
rect 1911 2519 1915 2520
rect 1534 2510 1540 2511
rect 1543 2510 1547 2511
rect 1511 2505 1515 2506
rect 998 2500 1004 2501
rect 1018 2503 1024 2504
rect 958 2498 964 2499
rect 1018 2499 1019 2503
rect 1023 2499 1024 2503
rect 1062 2501 1063 2505
rect 1067 2501 1068 2505
rect 1286 2504 1292 2505
rect 1062 2500 1068 2501
rect 1070 2503 1076 2504
rect 1018 2498 1024 2499
rect 1070 2499 1071 2503
rect 1075 2499 1076 2503
rect 1286 2500 1287 2504
rect 1291 2500 1292 2504
rect 1286 2499 1292 2500
rect 1070 2498 1076 2499
rect 598 2484 604 2485
rect 598 2480 599 2484
rect 603 2480 604 2484
rect 598 2479 604 2480
rect 662 2484 668 2485
rect 662 2480 663 2484
rect 667 2480 668 2484
rect 662 2479 668 2480
rect 726 2484 732 2485
rect 726 2480 727 2484
rect 731 2480 732 2484
rect 726 2479 732 2480
rect 790 2484 796 2485
rect 790 2480 791 2484
rect 795 2480 796 2484
rect 790 2479 796 2480
rect 854 2484 860 2485
rect 854 2480 855 2484
rect 859 2480 860 2484
rect 854 2479 860 2480
rect 918 2484 924 2485
rect 918 2480 919 2484
rect 923 2480 924 2484
rect 918 2479 924 2480
rect 982 2484 988 2485
rect 982 2480 983 2484
rect 987 2480 988 2484
rect 982 2479 988 2480
rect 1046 2484 1052 2485
rect 1046 2480 1047 2484
rect 1051 2480 1052 2484
rect 1046 2479 1052 2480
rect 600 2471 602 2479
rect 664 2471 666 2479
rect 728 2471 730 2479
rect 792 2471 794 2479
rect 856 2471 858 2479
rect 920 2471 922 2479
rect 984 2471 986 2479
rect 1048 2471 1050 2479
rect 599 2470 603 2471
rect 599 2465 603 2466
rect 615 2470 619 2471
rect 615 2465 619 2466
rect 663 2470 667 2471
rect 663 2465 667 2466
rect 671 2470 675 2471
rect 671 2465 675 2466
rect 727 2470 731 2471
rect 727 2465 731 2466
rect 783 2470 787 2471
rect 783 2465 787 2466
rect 791 2470 795 2471
rect 791 2465 795 2466
rect 839 2470 843 2471
rect 839 2465 843 2466
rect 855 2470 859 2471
rect 855 2465 859 2466
rect 895 2470 899 2471
rect 895 2465 899 2466
rect 919 2470 923 2471
rect 919 2465 923 2466
rect 951 2470 955 2471
rect 951 2465 955 2466
rect 983 2470 987 2471
rect 983 2465 987 2466
rect 1007 2470 1011 2471
rect 1007 2465 1011 2466
rect 1047 2470 1051 2471
rect 1047 2465 1051 2466
rect 1063 2470 1067 2471
rect 1063 2465 1067 2466
rect 614 2464 620 2465
rect 614 2460 615 2464
rect 619 2460 620 2464
rect 614 2459 620 2460
rect 670 2464 676 2465
rect 670 2460 671 2464
rect 675 2460 676 2464
rect 670 2459 676 2460
rect 726 2464 732 2465
rect 726 2460 727 2464
rect 731 2460 732 2464
rect 726 2459 732 2460
rect 782 2464 788 2465
rect 782 2460 783 2464
rect 787 2460 788 2464
rect 782 2459 788 2460
rect 838 2464 844 2465
rect 838 2460 839 2464
rect 843 2460 844 2464
rect 838 2459 844 2460
rect 894 2464 900 2465
rect 894 2460 895 2464
rect 899 2460 900 2464
rect 894 2459 900 2460
rect 950 2464 956 2465
rect 950 2460 951 2464
rect 955 2460 956 2464
rect 950 2459 956 2460
rect 1006 2464 1012 2465
rect 1006 2460 1007 2464
rect 1011 2460 1012 2464
rect 1006 2459 1012 2460
rect 1062 2464 1068 2465
rect 1062 2460 1063 2464
rect 1067 2460 1068 2464
rect 1062 2459 1068 2460
rect 167 2452 171 2453
rect 167 2447 171 2448
rect 495 2452 499 2453
rect 495 2447 499 2448
rect 567 2452 571 2453
rect 567 2447 571 2448
rect 875 2452 879 2453
rect 875 2447 879 2448
rect 110 2444 116 2445
rect 110 2440 111 2444
rect 115 2440 116 2444
rect 110 2439 116 2440
rect 112 2407 114 2439
rect 168 2424 170 2447
rect 876 2444 878 2447
rect 182 2443 188 2444
rect 182 2439 183 2443
rect 187 2439 188 2443
rect 182 2438 188 2439
rect 218 2443 224 2444
rect 218 2439 219 2443
rect 223 2439 224 2443
rect 218 2438 224 2439
rect 238 2443 244 2444
rect 238 2439 239 2443
rect 243 2439 244 2443
rect 238 2438 244 2439
rect 274 2443 280 2444
rect 274 2439 275 2443
rect 279 2439 280 2443
rect 274 2438 280 2439
rect 294 2443 300 2444
rect 294 2439 295 2443
rect 299 2439 300 2443
rect 294 2438 300 2439
rect 330 2443 336 2444
rect 330 2439 331 2443
rect 335 2439 336 2443
rect 330 2438 336 2439
rect 350 2443 356 2444
rect 350 2439 351 2443
rect 355 2439 356 2443
rect 350 2438 356 2439
rect 386 2443 392 2444
rect 386 2439 387 2443
rect 391 2439 392 2443
rect 386 2438 392 2439
rect 406 2443 412 2444
rect 406 2439 407 2443
rect 411 2439 412 2443
rect 406 2438 412 2439
rect 442 2443 448 2444
rect 442 2439 443 2443
rect 447 2439 448 2443
rect 442 2438 448 2439
rect 462 2443 468 2444
rect 462 2439 463 2443
rect 467 2439 468 2443
rect 462 2438 468 2439
rect 498 2443 504 2444
rect 498 2439 499 2443
rect 503 2439 504 2443
rect 498 2438 504 2439
rect 518 2443 524 2444
rect 518 2439 519 2443
rect 523 2439 524 2443
rect 518 2438 524 2439
rect 554 2443 560 2444
rect 554 2439 555 2443
rect 559 2439 560 2443
rect 554 2438 560 2439
rect 574 2443 580 2444
rect 574 2439 575 2443
rect 579 2439 580 2443
rect 574 2438 580 2439
rect 610 2443 616 2444
rect 610 2439 611 2443
rect 615 2439 616 2443
rect 610 2438 616 2439
rect 630 2443 636 2444
rect 630 2439 631 2443
rect 635 2439 636 2443
rect 630 2438 636 2439
rect 666 2443 672 2444
rect 666 2439 667 2443
rect 671 2439 672 2443
rect 666 2438 672 2439
rect 686 2443 692 2444
rect 686 2439 687 2443
rect 691 2439 692 2443
rect 686 2438 692 2439
rect 722 2443 728 2444
rect 722 2439 723 2443
rect 727 2439 728 2443
rect 722 2438 728 2439
rect 742 2443 748 2444
rect 742 2439 743 2443
rect 747 2439 748 2443
rect 742 2438 748 2439
rect 778 2443 784 2444
rect 778 2439 779 2443
rect 783 2439 784 2443
rect 778 2438 784 2439
rect 798 2443 804 2444
rect 798 2439 799 2443
rect 803 2439 804 2443
rect 798 2438 804 2439
rect 834 2443 840 2444
rect 834 2439 835 2443
rect 839 2439 840 2443
rect 834 2438 840 2439
rect 854 2443 860 2444
rect 854 2439 855 2443
rect 859 2439 860 2443
rect 854 2438 860 2439
rect 874 2443 880 2444
rect 874 2439 875 2443
rect 879 2439 880 2443
rect 874 2438 880 2439
rect 910 2443 916 2444
rect 910 2439 911 2443
rect 915 2439 916 2443
rect 910 2438 916 2439
rect 918 2443 924 2444
rect 918 2439 919 2443
rect 923 2439 924 2443
rect 918 2438 924 2439
rect 966 2443 972 2444
rect 966 2439 967 2443
rect 971 2439 972 2443
rect 966 2438 972 2439
rect 974 2443 980 2444
rect 974 2439 975 2443
rect 979 2439 980 2443
rect 974 2438 980 2439
rect 1022 2443 1028 2444
rect 1022 2439 1023 2443
rect 1027 2439 1028 2443
rect 1022 2438 1028 2439
rect 166 2423 172 2424
rect 166 2419 167 2423
rect 171 2419 172 2423
rect 166 2418 172 2419
rect 184 2407 186 2438
rect 220 2424 222 2438
rect 218 2423 224 2424
rect 218 2419 219 2423
rect 223 2419 224 2423
rect 218 2418 224 2419
rect 240 2407 242 2438
rect 276 2424 278 2438
rect 274 2423 280 2424
rect 274 2419 275 2423
rect 279 2419 280 2423
rect 274 2418 280 2419
rect 296 2407 298 2438
rect 332 2424 334 2438
rect 330 2423 336 2424
rect 330 2419 331 2423
rect 335 2419 336 2423
rect 330 2418 336 2419
rect 352 2407 354 2438
rect 388 2424 390 2438
rect 386 2423 392 2424
rect 386 2419 387 2423
rect 391 2419 392 2423
rect 386 2418 392 2419
rect 408 2407 410 2438
rect 444 2424 446 2438
rect 442 2423 448 2424
rect 442 2419 443 2423
rect 447 2419 448 2423
rect 442 2418 448 2419
rect 464 2407 466 2438
rect 500 2424 502 2438
rect 498 2423 504 2424
rect 498 2419 499 2423
rect 503 2419 504 2423
rect 498 2418 504 2419
rect 520 2407 522 2438
rect 556 2424 558 2438
rect 554 2423 560 2424
rect 554 2419 555 2423
rect 559 2419 560 2423
rect 554 2418 560 2419
rect 576 2407 578 2438
rect 612 2424 614 2438
rect 610 2423 616 2424
rect 610 2419 611 2423
rect 615 2419 616 2423
rect 610 2418 616 2419
rect 632 2407 634 2438
rect 668 2424 670 2438
rect 666 2423 672 2424
rect 666 2419 667 2423
rect 671 2419 672 2423
rect 666 2418 672 2419
rect 688 2407 690 2438
rect 724 2424 726 2438
rect 722 2423 728 2424
rect 722 2419 723 2423
rect 727 2419 728 2423
rect 722 2418 728 2419
rect 744 2407 746 2438
rect 780 2424 782 2438
rect 778 2423 784 2424
rect 778 2419 779 2423
rect 783 2419 784 2423
rect 778 2418 784 2419
rect 800 2407 802 2438
rect 836 2424 838 2438
rect 834 2423 840 2424
rect 834 2419 835 2423
rect 839 2419 840 2423
rect 834 2418 840 2419
rect 856 2407 858 2438
rect 912 2407 914 2438
rect 111 2406 115 2407
rect 111 2401 115 2402
rect 183 2406 187 2407
rect 183 2401 187 2402
rect 239 2406 243 2407
rect 239 2401 243 2402
rect 295 2406 299 2407
rect 295 2401 299 2402
rect 351 2406 355 2407
rect 351 2401 355 2402
rect 407 2406 411 2407
rect 407 2401 411 2402
rect 463 2406 467 2407
rect 463 2401 467 2402
rect 519 2406 523 2407
rect 519 2401 523 2402
rect 575 2406 579 2407
rect 575 2401 579 2402
rect 631 2406 635 2407
rect 631 2401 635 2402
rect 687 2406 691 2407
rect 687 2401 691 2402
rect 743 2406 747 2407
rect 743 2401 747 2402
rect 799 2406 803 2407
rect 799 2401 803 2402
rect 855 2406 859 2407
rect 855 2401 859 2402
rect 911 2406 915 2407
rect 911 2401 915 2402
rect 112 2381 114 2401
rect 520 2382 522 2401
rect 576 2382 578 2401
rect 632 2382 634 2401
rect 688 2382 690 2401
rect 920 2400 922 2438
rect 968 2407 970 2438
rect 976 2420 978 2438
rect 974 2419 980 2420
rect 974 2415 975 2419
rect 979 2415 980 2419
rect 974 2414 980 2415
rect 1024 2407 1026 2438
rect 1072 2424 1074 2498
rect 1286 2487 1292 2488
rect 1286 2483 1287 2487
rect 1291 2483 1292 2487
rect 1328 2485 1330 2505
rect 1528 2493 1530 2510
rect 1543 2505 1547 2506
rect 1567 2510 1571 2511
rect 1598 2510 1604 2511
rect 1607 2510 1611 2511
rect 1567 2505 1571 2506
rect 1607 2505 1611 2506
rect 1623 2510 1627 2511
rect 1658 2510 1664 2511
rect 1679 2510 1683 2511
rect 1714 2510 1720 2511
rect 1735 2510 1739 2511
rect 1623 2505 1627 2506
rect 1679 2505 1683 2506
rect 1735 2505 1739 2506
rect 1751 2510 1755 2511
rect 1770 2510 1776 2511
rect 1791 2510 1795 2511
rect 1814 2510 1820 2511
rect 1823 2510 1827 2511
rect 1751 2505 1755 2506
rect 1791 2505 1795 2506
rect 1823 2505 1827 2506
rect 1847 2510 1851 2511
rect 1882 2510 1888 2511
rect 1895 2510 1899 2511
rect 1847 2505 1851 2506
rect 1895 2505 1899 2506
rect 1903 2510 1907 2511
rect 1903 2505 1907 2506
rect 1527 2492 1531 2493
rect 1527 2487 1531 2488
rect 1544 2486 1546 2505
rect 1574 2503 1580 2504
rect 1566 2499 1572 2500
rect 1566 2495 1567 2499
rect 1571 2495 1572 2499
rect 1574 2499 1575 2503
rect 1579 2499 1580 2503
rect 1574 2498 1580 2499
rect 1566 2494 1572 2495
rect 1542 2485 1548 2486
rect 1286 2482 1292 2483
rect 1326 2484 1332 2485
rect 1288 2471 1290 2482
rect 1326 2480 1327 2484
rect 1331 2480 1332 2484
rect 1542 2481 1543 2485
rect 1547 2481 1548 2485
rect 1542 2480 1548 2481
rect 1326 2479 1332 2480
rect 1287 2470 1291 2471
rect 1287 2465 1291 2466
rect 1326 2467 1332 2468
rect 1288 2462 1290 2465
rect 1326 2463 1327 2467
rect 1331 2463 1332 2467
rect 1326 2462 1332 2463
rect 1526 2464 1532 2465
rect 1286 2461 1292 2462
rect 1286 2457 1287 2461
rect 1291 2457 1292 2461
rect 1286 2456 1292 2457
rect 1328 2455 1330 2462
rect 1526 2460 1527 2464
rect 1531 2460 1532 2464
rect 1526 2459 1532 2460
rect 1528 2455 1530 2459
rect 1327 2454 1331 2455
rect 1327 2449 1331 2450
rect 1527 2454 1531 2455
rect 1527 2449 1531 2450
rect 1543 2454 1547 2455
rect 1543 2449 1547 2450
rect 1328 2446 1330 2449
rect 1542 2448 1548 2449
rect 1326 2445 1332 2446
rect 1286 2444 1292 2445
rect 1078 2443 1084 2444
rect 1078 2439 1079 2443
rect 1083 2439 1084 2443
rect 1286 2440 1287 2444
rect 1291 2440 1292 2444
rect 1326 2441 1327 2445
rect 1331 2441 1332 2445
rect 1542 2444 1543 2448
rect 1547 2444 1548 2448
rect 1542 2443 1548 2444
rect 1326 2440 1332 2441
rect 1286 2439 1292 2440
rect 1078 2438 1084 2439
rect 1070 2423 1076 2424
rect 1070 2419 1071 2423
rect 1075 2419 1076 2423
rect 1070 2418 1076 2419
rect 1080 2407 1082 2438
rect 1288 2407 1290 2439
rect 1326 2428 1332 2429
rect 1568 2428 1570 2494
rect 1576 2484 1578 2498
rect 1608 2486 1610 2505
rect 1630 2503 1636 2504
rect 1630 2499 1631 2503
rect 1635 2499 1636 2503
rect 1630 2498 1636 2499
rect 1606 2485 1612 2486
rect 1574 2483 1580 2484
rect 1574 2479 1575 2483
rect 1579 2479 1580 2483
rect 1606 2481 1607 2485
rect 1611 2481 1612 2485
rect 1632 2484 1634 2498
rect 1680 2486 1682 2505
rect 1702 2503 1708 2504
rect 1702 2499 1703 2503
rect 1707 2499 1708 2503
rect 1702 2498 1708 2499
rect 1678 2485 1684 2486
rect 1606 2480 1612 2481
rect 1630 2483 1636 2484
rect 1574 2478 1580 2479
rect 1630 2479 1631 2483
rect 1635 2479 1636 2483
rect 1678 2481 1679 2485
rect 1683 2481 1684 2485
rect 1704 2484 1706 2498
rect 1752 2486 1754 2505
rect 1774 2503 1780 2504
rect 1774 2499 1775 2503
rect 1779 2499 1780 2503
rect 1774 2498 1780 2499
rect 1750 2485 1756 2486
rect 1678 2480 1684 2481
rect 1702 2483 1708 2484
rect 1630 2478 1636 2479
rect 1702 2479 1703 2483
rect 1707 2479 1708 2483
rect 1750 2481 1751 2485
rect 1755 2481 1756 2485
rect 1776 2484 1778 2498
rect 1824 2486 1826 2505
rect 1843 2492 1847 2493
rect 1843 2487 1847 2488
rect 1822 2485 1828 2486
rect 1750 2480 1756 2481
rect 1774 2483 1780 2484
rect 1702 2478 1708 2479
rect 1774 2479 1775 2483
rect 1779 2479 1780 2483
rect 1822 2481 1823 2485
rect 1827 2481 1828 2485
rect 1844 2484 1846 2487
rect 1896 2486 1898 2505
rect 1912 2504 1914 2519
rect 1940 2516 1942 2530
rect 1938 2515 1944 2516
rect 1938 2511 1939 2515
rect 1943 2511 1944 2515
rect 1960 2511 1962 2530
rect 1996 2516 1998 2530
rect 1994 2515 2000 2516
rect 1994 2511 1995 2515
rect 1999 2511 2000 2515
rect 2016 2511 2018 2530
rect 2052 2516 2054 2530
rect 2050 2515 2056 2516
rect 2050 2511 2051 2515
rect 2055 2511 2056 2515
rect 2072 2511 2074 2530
rect 2104 2516 2106 2530
rect 2102 2515 2108 2516
rect 2102 2511 2103 2515
rect 2107 2511 2108 2515
rect 2128 2511 2130 2530
rect 2164 2516 2166 2530
rect 2162 2515 2168 2516
rect 2162 2511 2163 2515
rect 2167 2511 2168 2515
rect 2184 2511 2186 2530
rect 2192 2525 2194 2530
rect 2191 2524 2195 2525
rect 2191 2519 2195 2520
rect 2504 2511 2506 2531
rect 1938 2510 1944 2511
rect 1959 2510 1963 2511
rect 1959 2505 1963 2506
rect 1967 2510 1971 2511
rect 1994 2510 2000 2511
rect 2015 2510 2019 2511
rect 1967 2505 1971 2506
rect 2015 2505 2019 2506
rect 2039 2510 2043 2511
rect 2050 2510 2056 2511
rect 2071 2510 2075 2511
rect 2102 2510 2108 2511
rect 2111 2510 2115 2511
rect 2039 2505 2043 2506
rect 2071 2505 2075 2506
rect 2111 2505 2115 2506
rect 2127 2510 2131 2511
rect 2162 2510 2168 2511
rect 2183 2510 2187 2511
rect 2127 2505 2131 2506
rect 2183 2505 2187 2506
rect 2503 2510 2507 2511
rect 2503 2505 2507 2506
rect 1910 2503 1916 2504
rect 1910 2499 1911 2503
rect 1915 2499 1916 2503
rect 1910 2498 1916 2499
rect 1918 2503 1924 2504
rect 1918 2499 1919 2503
rect 1923 2499 1924 2503
rect 1918 2498 1924 2499
rect 1894 2485 1900 2486
rect 1822 2480 1828 2481
rect 1842 2483 1848 2484
rect 1774 2478 1780 2479
rect 1842 2479 1843 2483
rect 1847 2479 1848 2483
rect 1894 2481 1895 2485
rect 1899 2481 1900 2485
rect 1920 2484 1922 2498
rect 1968 2486 1970 2505
rect 1990 2503 1996 2504
rect 1990 2499 1991 2503
rect 1995 2499 1996 2503
rect 1990 2498 1996 2499
rect 1966 2485 1972 2486
rect 1894 2480 1900 2481
rect 1918 2483 1924 2484
rect 1842 2478 1848 2479
rect 1918 2479 1919 2483
rect 1923 2479 1924 2483
rect 1966 2481 1967 2485
rect 1971 2481 1972 2485
rect 1992 2484 1994 2498
rect 2040 2486 2042 2505
rect 2062 2503 2068 2504
rect 2062 2499 2063 2503
rect 2067 2499 2068 2503
rect 2062 2498 2068 2499
rect 2038 2485 2044 2486
rect 1966 2480 1972 2481
rect 1990 2483 1996 2484
rect 1918 2478 1924 2479
rect 1990 2479 1991 2483
rect 1995 2479 1996 2483
rect 2038 2481 2039 2485
rect 2043 2481 2044 2485
rect 2064 2484 2066 2498
rect 2112 2486 2114 2505
rect 2134 2503 2140 2504
rect 2134 2499 2135 2503
rect 2139 2499 2140 2503
rect 2134 2498 2140 2499
rect 2110 2485 2116 2486
rect 2038 2480 2044 2481
rect 2062 2483 2068 2484
rect 1990 2478 1996 2479
rect 2062 2479 2063 2483
rect 2067 2479 2068 2483
rect 2110 2481 2111 2485
rect 2115 2481 2116 2485
rect 2136 2484 2138 2498
rect 2184 2486 2186 2505
rect 2182 2485 2188 2486
rect 2504 2485 2506 2505
rect 2110 2480 2116 2481
rect 2134 2483 2140 2484
rect 2062 2478 2068 2479
rect 2134 2479 2135 2483
rect 2139 2479 2140 2483
rect 2182 2481 2183 2485
rect 2187 2481 2188 2485
rect 2502 2484 2508 2485
rect 2182 2480 2188 2481
rect 2190 2483 2196 2484
rect 2134 2478 2140 2479
rect 2190 2479 2191 2483
rect 2195 2479 2196 2483
rect 2502 2480 2503 2484
rect 2507 2480 2508 2484
rect 2502 2479 2508 2480
rect 2190 2478 2196 2479
rect 1590 2464 1596 2465
rect 1590 2460 1591 2464
rect 1595 2460 1596 2464
rect 1590 2459 1596 2460
rect 1662 2464 1668 2465
rect 1662 2460 1663 2464
rect 1667 2460 1668 2464
rect 1662 2459 1668 2460
rect 1734 2464 1740 2465
rect 1734 2460 1735 2464
rect 1739 2460 1740 2464
rect 1734 2459 1740 2460
rect 1806 2464 1812 2465
rect 1806 2460 1807 2464
rect 1811 2460 1812 2464
rect 1806 2459 1812 2460
rect 1878 2464 1884 2465
rect 1878 2460 1879 2464
rect 1883 2460 1884 2464
rect 1878 2459 1884 2460
rect 1950 2464 1956 2465
rect 1950 2460 1951 2464
rect 1955 2460 1956 2464
rect 1950 2459 1956 2460
rect 2022 2464 2028 2465
rect 2022 2460 2023 2464
rect 2027 2460 2028 2464
rect 2022 2459 2028 2460
rect 2094 2464 2100 2465
rect 2094 2460 2095 2464
rect 2099 2460 2100 2464
rect 2094 2459 2100 2460
rect 2166 2464 2172 2465
rect 2166 2460 2167 2464
rect 2171 2460 2172 2464
rect 2166 2459 2172 2460
rect 1592 2455 1594 2459
rect 1664 2455 1666 2459
rect 1736 2455 1738 2459
rect 1808 2455 1810 2459
rect 1880 2455 1882 2459
rect 1952 2455 1954 2459
rect 2024 2455 2026 2459
rect 2096 2455 2098 2459
rect 2168 2455 2170 2459
rect 1591 2454 1595 2455
rect 1591 2449 1595 2450
rect 1607 2454 1611 2455
rect 1607 2449 1611 2450
rect 1663 2454 1667 2455
rect 1663 2449 1667 2450
rect 1671 2454 1675 2455
rect 1671 2449 1675 2450
rect 1735 2454 1739 2455
rect 1735 2449 1739 2450
rect 1743 2454 1747 2455
rect 1743 2449 1747 2450
rect 1807 2454 1811 2455
rect 1807 2449 1811 2450
rect 1815 2454 1819 2455
rect 1815 2449 1819 2450
rect 1879 2454 1883 2455
rect 1879 2449 1883 2450
rect 1951 2454 1955 2455
rect 1951 2449 1955 2450
rect 2023 2454 2027 2455
rect 2023 2449 2027 2450
rect 2095 2454 2099 2455
rect 2095 2449 2099 2450
rect 2167 2454 2171 2455
rect 2167 2449 2171 2450
rect 1606 2448 1612 2449
rect 1606 2444 1607 2448
rect 1611 2444 1612 2448
rect 1606 2443 1612 2444
rect 1670 2448 1676 2449
rect 1670 2444 1671 2448
rect 1675 2444 1676 2448
rect 1670 2443 1676 2444
rect 1742 2448 1748 2449
rect 1742 2444 1743 2448
rect 1747 2444 1748 2448
rect 1742 2443 1748 2444
rect 1814 2448 1820 2449
rect 1814 2444 1815 2448
rect 1819 2444 1820 2448
rect 1814 2443 1820 2444
rect 1878 2448 1884 2449
rect 1878 2444 1879 2448
rect 1883 2444 1884 2448
rect 1878 2443 1884 2444
rect 1950 2448 1956 2449
rect 1950 2444 1951 2448
rect 1955 2444 1956 2448
rect 1950 2443 1956 2444
rect 2022 2448 2028 2449
rect 2022 2444 2023 2448
rect 2027 2444 2028 2448
rect 2022 2443 2028 2444
rect 2094 2448 2100 2449
rect 2094 2444 2095 2448
rect 2099 2444 2100 2448
rect 2094 2443 2100 2444
rect 2166 2448 2172 2449
rect 2166 2444 2167 2448
rect 2171 2444 2172 2448
rect 2166 2443 2172 2444
rect 1326 2424 1327 2428
rect 1331 2424 1332 2428
rect 1326 2423 1332 2424
rect 1558 2427 1564 2428
rect 1558 2423 1559 2427
rect 1563 2423 1564 2427
rect 967 2406 971 2407
rect 967 2401 971 2402
rect 1023 2406 1027 2407
rect 1023 2401 1027 2402
rect 1079 2406 1083 2407
rect 1079 2401 1083 2402
rect 1287 2406 1291 2407
rect 1287 2401 1291 2402
rect 918 2399 924 2400
rect 918 2395 919 2399
rect 923 2395 924 2399
rect 918 2394 924 2395
rect 518 2381 524 2382
rect 110 2380 116 2381
rect 110 2376 111 2380
rect 115 2376 116 2380
rect 518 2377 519 2381
rect 523 2377 524 2381
rect 574 2381 580 2382
rect 518 2376 524 2377
rect 542 2379 548 2380
rect 110 2375 116 2376
rect 542 2375 543 2379
rect 547 2375 548 2379
rect 574 2377 575 2381
rect 579 2377 580 2381
rect 574 2376 580 2377
rect 630 2381 636 2382
rect 630 2377 631 2381
rect 635 2377 636 2381
rect 630 2376 636 2377
rect 686 2381 692 2382
rect 1288 2381 1290 2401
rect 1328 2399 1330 2423
rect 1558 2422 1564 2423
rect 1566 2427 1572 2428
rect 1566 2423 1567 2427
rect 1571 2423 1572 2427
rect 1566 2422 1572 2423
rect 1622 2427 1628 2428
rect 1622 2423 1623 2427
rect 1627 2423 1628 2427
rect 1622 2422 1628 2423
rect 1686 2427 1692 2428
rect 1686 2423 1687 2427
rect 1691 2423 1692 2427
rect 1686 2422 1692 2423
rect 1758 2427 1764 2428
rect 1758 2423 1759 2427
rect 1763 2423 1764 2427
rect 1758 2422 1764 2423
rect 1830 2427 1836 2428
rect 1830 2423 1831 2427
rect 1835 2423 1836 2427
rect 1830 2422 1836 2423
rect 1894 2427 1900 2428
rect 1894 2423 1895 2427
rect 1899 2423 1900 2427
rect 1894 2422 1900 2423
rect 1946 2427 1952 2428
rect 1946 2423 1947 2427
rect 1951 2423 1952 2427
rect 1946 2422 1952 2423
rect 1966 2427 1972 2428
rect 1966 2423 1967 2427
rect 1971 2423 1972 2427
rect 1966 2422 1972 2423
rect 1974 2427 1980 2428
rect 1974 2423 1975 2427
rect 1979 2423 1980 2427
rect 1974 2422 1980 2423
rect 2038 2427 2044 2428
rect 2038 2423 2039 2427
rect 2043 2423 2044 2427
rect 2038 2422 2044 2423
rect 2054 2427 2060 2428
rect 2054 2423 2055 2427
rect 2059 2423 2060 2427
rect 2054 2422 2060 2423
rect 2110 2427 2116 2428
rect 2110 2423 2111 2427
rect 2115 2423 2116 2427
rect 2110 2422 2116 2423
rect 2182 2427 2188 2428
rect 2182 2423 2183 2427
rect 2187 2423 2188 2427
rect 2182 2422 2188 2423
rect 1560 2399 1562 2422
rect 1624 2399 1626 2422
rect 1688 2399 1690 2422
rect 1760 2399 1762 2422
rect 1810 2407 1816 2408
rect 1810 2403 1811 2407
rect 1815 2403 1816 2407
rect 1810 2402 1816 2403
rect 1327 2398 1331 2399
rect 1327 2393 1331 2394
rect 1559 2398 1563 2399
rect 1559 2393 1563 2394
rect 1567 2398 1571 2399
rect 1567 2393 1571 2394
rect 1623 2398 1627 2399
rect 1623 2393 1627 2394
rect 1679 2398 1683 2399
rect 1679 2393 1683 2394
rect 1687 2398 1691 2399
rect 1687 2393 1691 2394
rect 1735 2398 1739 2399
rect 1735 2393 1739 2394
rect 1759 2398 1763 2399
rect 1759 2393 1763 2394
rect 1791 2398 1795 2399
rect 1791 2393 1795 2394
rect 686 2377 687 2381
rect 691 2377 692 2381
rect 686 2376 692 2377
rect 1286 2380 1292 2381
rect 1286 2376 1287 2380
rect 1291 2376 1292 2380
rect 1286 2375 1292 2376
rect 542 2374 548 2375
rect 110 2363 116 2364
rect 110 2359 111 2363
rect 115 2359 116 2363
rect 110 2358 116 2359
rect 502 2360 508 2361
rect 112 2347 114 2358
rect 502 2356 503 2360
rect 507 2356 508 2360
rect 502 2355 508 2356
rect 504 2347 506 2355
rect 111 2346 115 2347
rect 111 2341 115 2342
rect 319 2346 323 2347
rect 319 2341 323 2342
rect 391 2346 395 2347
rect 391 2341 395 2342
rect 463 2346 467 2347
rect 463 2341 467 2342
rect 503 2346 507 2347
rect 503 2341 507 2342
rect 535 2346 539 2347
rect 535 2341 539 2342
rect 112 2338 114 2341
rect 318 2340 324 2341
rect 110 2337 116 2338
rect 110 2333 111 2337
rect 115 2333 116 2337
rect 318 2336 319 2340
rect 323 2336 324 2340
rect 318 2335 324 2336
rect 390 2340 396 2341
rect 390 2336 391 2340
rect 395 2336 396 2340
rect 390 2335 396 2336
rect 462 2340 468 2341
rect 462 2336 463 2340
rect 467 2336 468 2340
rect 462 2335 468 2336
rect 534 2340 540 2341
rect 534 2336 535 2340
rect 539 2336 540 2340
rect 534 2335 540 2336
rect 110 2332 116 2333
rect 110 2320 116 2321
rect 110 2316 111 2320
rect 115 2316 116 2320
rect 110 2315 116 2316
rect 334 2319 340 2320
rect 334 2315 335 2319
rect 339 2315 340 2319
rect 112 2287 114 2315
rect 334 2314 340 2315
rect 386 2319 392 2320
rect 386 2315 387 2319
rect 391 2315 392 2319
rect 386 2314 392 2315
rect 406 2319 412 2320
rect 406 2315 407 2319
rect 411 2315 412 2319
rect 406 2314 412 2315
rect 458 2319 464 2320
rect 458 2315 459 2319
rect 463 2315 464 2319
rect 458 2314 464 2315
rect 478 2319 484 2320
rect 478 2315 479 2319
rect 483 2315 484 2319
rect 478 2314 484 2315
rect 336 2287 338 2314
rect 388 2300 390 2314
rect 386 2299 392 2300
rect 386 2295 387 2299
rect 391 2295 392 2299
rect 386 2294 392 2295
rect 408 2287 410 2314
rect 111 2286 115 2287
rect 111 2281 115 2282
rect 175 2286 179 2287
rect 175 2281 179 2282
rect 271 2286 275 2287
rect 271 2281 275 2282
rect 335 2286 339 2287
rect 335 2281 339 2282
rect 375 2286 379 2287
rect 375 2281 379 2282
rect 407 2286 411 2287
rect 407 2281 411 2282
rect 112 2261 114 2281
rect 176 2262 178 2281
rect 272 2262 274 2281
rect 376 2262 378 2281
rect 460 2280 462 2314
rect 480 2287 482 2314
rect 544 2300 546 2374
rect 1328 2373 1330 2393
rect 1568 2374 1570 2393
rect 1590 2391 1596 2392
rect 1590 2387 1591 2391
rect 1595 2387 1596 2391
rect 1590 2386 1596 2387
rect 1566 2373 1572 2374
rect 1326 2372 1332 2373
rect 1326 2368 1327 2372
rect 1331 2368 1332 2372
rect 1566 2369 1567 2373
rect 1571 2369 1572 2373
rect 1592 2372 1594 2386
rect 1624 2374 1626 2393
rect 1646 2391 1652 2392
rect 1646 2387 1647 2391
rect 1651 2387 1652 2391
rect 1646 2386 1652 2387
rect 1622 2373 1628 2374
rect 1566 2368 1572 2369
rect 1590 2371 1596 2372
rect 1326 2367 1332 2368
rect 1590 2367 1591 2371
rect 1595 2367 1596 2371
rect 1622 2369 1623 2373
rect 1627 2369 1628 2373
rect 1648 2372 1650 2386
rect 1680 2374 1682 2393
rect 1702 2391 1708 2392
rect 1702 2387 1703 2391
rect 1707 2387 1708 2391
rect 1702 2386 1708 2387
rect 1678 2373 1684 2374
rect 1622 2368 1628 2369
rect 1646 2371 1652 2372
rect 1590 2366 1596 2367
rect 1646 2367 1647 2371
rect 1651 2367 1652 2371
rect 1678 2369 1679 2373
rect 1683 2369 1684 2373
rect 1704 2372 1706 2386
rect 1736 2374 1738 2393
rect 1766 2391 1772 2392
rect 1766 2387 1767 2391
rect 1771 2387 1772 2391
rect 1766 2386 1772 2387
rect 1734 2373 1740 2374
rect 1678 2368 1684 2369
rect 1702 2371 1708 2372
rect 1646 2366 1652 2367
rect 1702 2367 1703 2371
rect 1707 2367 1708 2371
rect 1734 2369 1735 2373
rect 1739 2369 1740 2373
rect 1768 2372 1770 2386
rect 1782 2383 1788 2384
rect 1782 2379 1783 2383
rect 1787 2379 1788 2383
rect 1782 2378 1788 2379
rect 1734 2368 1740 2369
rect 1766 2371 1772 2372
rect 1702 2366 1708 2367
rect 1766 2367 1767 2371
rect 1771 2367 1772 2371
rect 1766 2366 1772 2367
rect 1286 2363 1292 2364
rect 558 2360 564 2361
rect 558 2356 559 2360
rect 563 2356 564 2360
rect 558 2355 564 2356
rect 614 2360 620 2361
rect 614 2356 615 2360
rect 619 2356 620 2360
rect 614 2355 620 2356
rect 670 2360 676 2361
rect 670 2356 671 2360
rect 675 2356 676 2360
rect 1286 2359 1287 2363
rect 1291 2359 1292 2363
rect 1286 2358 1292 2359
rect 670 2355 676 2356
rect 560 2347 562 2355
rect 616 2347 618 2355
rect 672 2347 674 2355
rect 1288 2347 1290 2358
rect 1326 2355 1332 2356
rect 1326 2351 1327 2355
rect 1331 2351 1332 2355
rect 1326 2350 1332 2351
rect 1550 2352 1556 2353
rect 559 2346 563 2347
rect 559 2341 563 2342
rect 607 2346 611 2347
rect 607 2341 611 2342
rect 615 2346 619 2347
rect 615 2341 619 2342
rect 671 2346 675 2347
rect 671 2341 675 2342
rect 679 2346 683 2347
rect 679 2341 683 2342
rect 743 2346 747 2347
rect 743 2341 747 2342
rect 807 2346 811 2347
rect 807 2341 811 2342
rect 863 2346 867 2347
rect 863 2341 867 2342
rect 927 2346 931 2347
rect 927 2341 931 2342
rect 991 2346 995 2347
rect 991 2341 995 2342
rect 1055 2346 1059 2347
rect 1055 2341 1059 2342
rect 1111 2346 1115 2347
rect 1111 2341 1115 2342
rect 1167 2346 1171 2347
rect 1167 2341 1171 2342
rect 1223 2346 1227 2347
rect 1223 2341 1227 2342
rect 1287 2346 1291 2347
rect 1287 2341 1291 2342
rect 606 2340 612 2341
rect 606 2336 607 2340
rect 611 2336 612 2340
rect 606 2335 612 2336
rect 678 2340 684 2341
rect 678 2336 679 2340
rect 683 2336 684 2340
rect 678 2335 684 2336
rect 742 2340 748 2341
rect 742 2336 743 2340
rect 747 2336 748 2340
rect 742 2335 748 2336
rect 806 2340 812 2341
rect 806 2336 807 2340
rect 811 2336 812 2340
rect 806 2335 812 2336
rect 862 2340 868 2341
rect 862 2336 863 2340
rect 867 2336 868 2340
rect 862 2335 868 2336
rect 926 2340 932 2341
rect 926 2336 927 2340
rect 931 2336 932 2340
rect 926 2335 932 2336
rect 990 2340 996 2341
rect 990 2336 991 2340
rect 995 2336 996 2340
rect 990 2335 996 2336
rect 1054 2340 1060 2341
rect 1054 2336 1055 2340
rect 1059 2336 1060 2340
rect 1054 2335 1060 2336
rect 1110 2340 1116 2341
rect 1110 2336 1111 2340
rect 1115 2336 1116 2340
rect 1110 2335 1116 2336
rect 1166 2340 1172 2341
rect 1166 2336 1167 2340
rect 1171 2336 1172 2340
rect 1166 2335 1172 2336
rect 1222 2340 1228 2341
rect 1222 2336 1223 2340
rect 1227 2336 1228 2340
rect 1288 2338 1290 2341
rect 1328 2339 1330 2350
rect 1550 2348 1551 2352
rect 1555 2348 1556 2352
rect 1550 2347 1556 2348
rect 1606 2352 1612 2353
rect 1606 2348 1607 2352
rect 1611 2348 1612 2352
rect 1606 2347 1612 2348
rect 1662 2352 1668 2353
rect 1662 2348 1663 2352
rect 1667 2348 1668 2352
rect 1662 2347 1668 2348
rect 1718 2352 1724 2353
rect 1718 2348 1719 2352
rect 1723 2348 1724 2352
rect 1718 2347 1724 2348
rect 1774 2352 1780 2353
rect 1774 2348 1775 2352
rect 1779 2348 1780 2352
rect 1774 2347 1780 2348
rect 1552 2339 1554 2347
rect 1608 2339 1610 2347
rect 1664 2339 1666 2347
rect 1720 2339 1722 2347
rect 1776 2339 1778 2347
rect 1327 2338 1331 2339
rect 1222 2335 1228 2336
rect 1286 2337 1292 2338
rect 1286 2333 1287 2337
rect 1291 2333 1292 2337
rect 1327 2333 1331 2334
rect 1471 2338 1475 2339
rect 1471 2333 1475 2334
rect 1535 2338 1539 2339
rect 1535 2333 1539 2334
rect 1551 2338 1555 2339
rect 1551 2333 1555 2334
rect 1607 2338 1611 2339
rect 1607 2333 1611 2334
rect 1663 2338 1667 2339
rect 1663 2333 1667 2334
rect 1687 2338 1691 2339
rect 1687 2333 1691 2334
rect 1719 2338 1723 2339
rect 1719 2333 1723 2334
rect 1759 2338 1763 2339
rect 1759 2333 1763 2334
rect 1775 2338 1779 2339
rect 1775 2333 1779 2334
rect 1286 2332 1292 2333
rect 1328 2330 1330 2333
rect 1470 2332 1476 2333
rect 1326 2329 1332 2330
rect 1326 2325 1327 2329
rect 1331 2325 1332 2329
rect 1470 2328 1471 2332
rect 1475 2328 1476 2332
rect 1470 2327 1476 2328
rect 1534 2332 1540 2333
rect 1534 2328 1535 2332
rect 1539 2328 1540 2332
rect 1534 2327 1540 2328
rect 1606 2332 1612 2333
rect 1606 2328 1607 2332
rect 1611 2328 1612 2332
rect 1606 2327 1612 2328
rect 1686 2332 1692 2333
rect 1686 2328 1687 2332
rect 1691 2328 1692 2332
rect 1686 2327 1692 2328
rect 1758 2332 1764 2333
rect 1758 2328 1759 2332
rect 1763 2328 1764 2332
rect 1758 2327 1764 2328
rect 1326 2324 1332 2325
rect 1286 2320 1292 2321
rect 550 2319 556 2320
rect 550 2315 551 2319
rect 555 2315 556 2319
rect 550 2314 556 2315
rect 622 2319 628 2320
rect 622 2315 623 2319
rect 627 2315 628 2319
rect 622 2314 628 2315
rect 674 2319 680 2320
rect 674 2315 675 2319
rect 679 2315 680 2319
rect 674 2314 680 2315
rect 694 2319 700 2320
rect 694 2315 695 2319
rect 699 2315 700 2319
rect 694 2314 700 2315
rect 710 2319 716 2320
rect 710 2315 711 2319
rect 715 2315 716 2319
rect 710 2314 716 2315
rect 758 2319 764 2320
rect 758 2315 759 2319
rect 763 2315 764 2319
rect 758 2314 764 2315
rect 766 2319 772 2320
rect 766 2315 767 2319
rect 771 2315 772 2319
rect 766 2314 772 2315
rect 822 2319 828 2320
rect 822 2315 823 2319
rect 827 2315 828 2319
rect 822 2314 828 2315
rect 878 2319 884 2320
rect 878 2315 879 2319
rect 883 2315 884 2319
rect 878 2314 884 2315
rect 942 2319 948 2320
rect 942 2315 943 2319
rect 947 2315 948 2319
rect 942 2314 948 2315
rect 1006 2319 1012 2320
rect 1006 2315 1007 2319
rect 1011 2315 1012 2319
rect 1006 2314 1012 2315
rect 1070 2319 1076 2320
rect 1070 2315 1071 2319
rect 1075 2315 1076 2319
rect 1070 2314 1076 2315
rect 1078 2319 1084 2320
rect 1078 2315 1079 2319
rect 1083 2315 1084 2319
rect 1078 2314 1084 2315
rect 1126 2319 1132 2320
rect 1126 2315 1127 2319
rect 1131 2315 1132 2319
rect 1126 2314 1132 2315
rect 1182 2319 1188 2320
rect 1182 2315 1183 2319
rect 1187 2315 1188 2319
rect 1182 2314 1188 2315
rect 1238 2319 1244 2320
rect 1238 2315 1239 2319
rect 1243 2315 1244 2319
rect 1286 2316 1287 2320
rect 1291 2316 1292 2320
rect 1286 2315 1292 2316
rect 1238 2314 1244 2315
rect 542 2299 548 2300
rect 542 2295 543 2299
rect 547 2295 548 2299
rect 542 2294 548 2295
rect 552 2287 554 2314
rect 624 2287 626 2314
rect 676 2300 678 2314
rect 674 2299 680 2300
rect 674 2295 675 2299
rect 679 2295 680 2299
rect 674 2294 680 2295
rect 696 2287 698 2314
rect 479 2286 483 2287
rect 479 2281 483 2282
rect 551 2286 555 2287
rect 551 2281 555 2282
rect 591 2286 595 2287
rect 591 2281 595 2282
rect 623 2286 627 2287
rect 623 2281 627 2282
rect 695 2286 699 2287
rect 695 2281 699 2282
rect 703 2286 707 2287
rect 703 2281 707 2282
rect 458 2279 464 2280
rect 458 2275 459 2279
rect 463 2275 464 2279
rect 458 2274 464 2275
rect 480 2262 482 2281
rect 502 2279 508 2280
rect 502 2275 503 2279
rect 507 2275 508 2279
rect 502 2274 508 2275
rect 174 2261 180 2262
rect 110 2260 116 2261
rect 110 2256 111 2260
rect 115 2256 116 2260
rect 174 2257 175 2261
rect 179 2257 180 2261
rect 270 2261 276 2262
rect 174 2256 180 2257
rect 182 2259 188 2260
rect 110 2255 116 2256
rect 182 2255 183 2259
rect 187 2255 188 2259
rect 270 2257 271 2261
rect 275 2257 276 2261
rect 270 2256 276 2257
rect 374 2261 380 2262
rect 374 2257 375 2261
rect 379 2257 380 2261
rect 374 2256 380 2257
rect 478 2261 484 2262
rect 478 2257 479 2261
rect 483 2257 484 2261
rect 504 2260 506 2274
rect 592 2262 594 2281
rect 704 2262 706 2281
rect 712 2280 714 2314
rect 760 2287 762 2314
rect 768 2292 770 2314
rect 766 2291 772 2292
rect 766 2287 767 2291
rect 771 2287 772 2291
rect 824 2287 826 2314
rect 880 2287 882 2314
rect 944 2287 946 2314
rect 1008 2287 1010 2314
rect 1072 2287 1074 2314
rect 1080 2296 1082 2314
rect 1078 2295 1084 2296
rect 1078 2291 1079 2295
rect 1083 2291 1084 2295
rect 1078 2290 1084 2291
rect 1128 2287 1130 2314
rect 1184 2287 1186 2314
rect 1240 2287 1242 2314
rect 1258 2299 1264 2300
rect 1258 2295 1259 2299
rect 1263 2295 1264 2299
rect 1258 2294 1264 2295
rect 759 2286 763 2287
rect 766 2286 772 2287
rect 807 2286 811 2287
rect 759 2281 763 2282
rect 807 2281 811 2282
rect 823 2286 827 2287
rect 823 2281 827 2282
rect 879 2286 883 2287
rect 879 2281 883 2282
rect 911 2286 915 2287
rect 911 2281 915 2282
rect 943 2286 947 2287
rect 943 2281 947 2282
rect 1007 2286 1011 2287
rect 1007 2281 1011 2282
rect 1015 2286 1019 2287
rect 1015 2281 1019 2282
rect 1071 2286 1075 2287
rect 1071 2281 1075 2282
rect 1127 2286 1131 2287
rect 1127 2281 1131 2282
rect 1183 2286 1187 2287
rect 1183 2281 1187 2282
rect 1239 2286 1243 2287
rect 1239 2281 1243 2282
rect 710 2279 716 2280
rect 710 2275 711 2279
rect 715 2275 716 2279
rect 710 2274 716 2275
rect 726 2279 732 2280
rect 726 2275 727 2279
rect 731 2275 732 2279
rect 726 2274 732 2275
rect 590 2261 596 2262
rect 478 2256 484 2257
rect 502 2259 508 2260
rect 182 2254 188 2255
rect 502 2255 503 2259
rect 507 2255 508 2259
rect 590 2257 591 2261
rect 595 2257 596 2261
rect 590 2256 596 2257
rect 702 2261 708 2262
rect 702 2257 703 2261
rect 707 2257 708 2261
rect 728 2260 730 2274
rect 808 2262 810 2281
rect 830 2279 836 2280
rect 830 2275 831 2279
rect 835 2275 836 2279
rect 830 2274 836 2275
rect 806 2261 812 2262
rect 702 2256 708 2257
rect 726 2259 732 2260
rect 502 2254 508 2255
rect 726 2255 727 2259
rect 731 2255 732 2259
rect 806 2257 807 2261
rect 811 2257 812 2261
rect 832 2260 834 2274
rect 912 2262 914 2281
rect 1016 2262 1018 2281
rect 1038 2279 1044 2280
rect 1038 2275 1039 2279
rect 1043 2275 1044 2279
rect 1038 2274 1044 2275
rect 910 2261 916 2262
rect 806 2256 812 2257
rect 830 2259 836 2260
rect 726 2254 732 2255
rect 830 2255 831 2259
rect 835 2255 836 2259
rect 910 2257 911 2261
rect 915 2257 916 2261
rect 1014 2261 1020 2262
rect 910 2256 916 2257
rect 926 2259 932 2260
rect 830 2254 836 2255
rect 926 2255 927 2259
rect 931 2255 932 2259
rect 1014 2257 1015 2261
rect 1019 2257 1020 2261
rect 1040 2260 1042 2274
rect 1074 2271 1080 2272
rect 1074 2267 1075 2271
rect 1079 2267 1080 2271
rect 1074 2266 1080 2267
rect 1014 2256 1020 2257
rect 1038 2259 1044 2260
rect 926 2254 932 2255
rect 1038 2255 1039 2259
rect 1043 2255 1044 2259
rect 1038 2254 1044 2255
rect 110 2243 116 2244
rect 110 2239 111 2243
rect 115 2239 116 2243
rect 110 2238 116 2239
rect 158 2240 164 2241
rect 112 2235 114 2238
rect 158 2236 159 2240
rect 163 2236 164 2240
rect 158 2235 164 2236
rect 111 2234 115 2235
rect 111 2229 115 2230
rect 143 2234 147 2235
rect 143 2229 147 2230
rect 159 2234 163 2235
rect 159 2229 163 2230
rect 112 2226 114 2229
rect 142 2228 148 2229
rect 110 2225 116 2226
rect 110 2221 111 2225
rect 115 2221 116 2225
rect 142 2224 143 2228
rect 147 2224 148 2228
rect 142 2223 148 2224
rect 110 2220 116 2221
rect 110 2208 116 2209
rect 110 2204 111 2208
rect 115 2204 116 2208
rect 110 2203 116 2204
rect 158 2207 164 2208
rect 158 2203 159 2207
rect 163 2203 164 2207
rect 112 2183 114 2203
rect 158 2202 164 2203
rect 160 2183 162 2202
rect 184 2188 186 2254
rect 254 2240 260 2241
rect 254 2236 255 2240
rect 259 2236 260 2240
rect 254 2235 260 2236
rect 358 2240 364 2241
rect 358 2236 359 2240
rect 363 2236 364 2240
rect 358 2235 364 2236
rect 462 2240 468 2241
rect 462 2236 463 2240
rect 467 2236 468 2240
rect 462 2235 468 2236
rect 574 2240 580 2241
rect 574 2236 575 2240
rect 579 2236 580 2240
rect 574 2235 580 2236
rect 686 2240 692 2241
rect 686 2236 687 2240
rect 691 2236 692 2240
rect 686 2235 692 2236
rect 790 2240 796 2241
rect 790 2236 791 2240
rect 795 2236 796 2240
rect 790 2235 796 2236
rect 894 2240 900 2241
rect 894 2236 895 2240
rect 899 2236 900 2240
rect 894 2235 900 2236
rect 231 2234 235 2235
rect 231 2229 235 2230
rect 255 2234 259 2235
rect 255 2229 259 2230
rect 319 2234 323 2235
rect 319 2229 323 2230
rect 359 2234 363 2235
rect 359 2229 363 2230
rect 415 2234 419 2235
rect 415 2229 419 2230
rect 463 2234 467 2235
rect 463 2229 467 2230
rect 519 2234 523 2235
rect 519 2229 523 2230
rect 575 2234 579 2235
rect 575 2229 579 2230
rect 623 2234 627 2235
rect 623 2229 627 2230
rect 687 2234 691 2235
rect 687 2229 691 2230
rect 727 2234 731 2235
rect 727 2229 731 2230
rect 791 2234 795 2235
rect 791 2229 795 2230
rect 831 2234 835 2235
rect 831 2229 835 2230
rect 895 2234 899 2235
rect 895 2229 899 2230
rect 230 2228 236 2229
rect 230 2224 231 2228
rect 235 2224 236 2228
rect 230 2223 236 2224
rect 318 2228 324 2229
rect 318 2224 319 2228
rect 323 2224 324 2228
rect 318 2223 324 2224
rect 414 2228 420 2229
rect 414 2224 415 2228
rect 419 2224 420 2228
rect 414 2223 420 2224
rect 518 2228 524 2229
rect 518 2224 519 2228
rect 523 2224 524 2228
rect 518 2223 524 2224
rect 622 2228 628 2229
rect 622 2224 623 2228
rect 627 2224 628 2228
rect 622 2223 628 2224
rect 726 2228 732 2229
rect 726 2224 727 2228
rect 731 2224 732 2228
rect 726 2223 732 2224
rect 830 2228 836 2229
rect 830 2224 831 2228
rect 835 2224 836 2228
rect 830 2223 836 2224
rect 226 2207 232 2208
rect 226 2203 227 2207
rect 231 2203 232 2207
rect 226 2202 232 2203
rect 246 2207 252 2208
rect 246 2203 247 2207
rect 251 2203 252 2207
rect 246 2202 252 2203
rect 314 2207 320 2208
rect 314 2203 315 2207
rect 319 2203 320 2207
rect 314 2202 320 2203
rect 334 2207 340 2208
rect 334 2203 335 2207
rect 339 2203 340 2207
rect 334 2202 340 2203
rect 410 2207 416 2208
rect 410 2203 411 2207
rect 415 2203 416 2207
rect 410 2202 416 2203
rect 430 2207 436 2208
rect 430 2203 431 2207
rect 435 2203 436 2207
rect 430 2202 436 2203
rect 514 2207 520 2208
rect 514 2203 515 2207
rect 519 2203 520 2207
rect 514 2202 520 2203
rect 534 2207 540 2208
rect 534 2203 535 2207
rect 539 2203 540 2207
rect 534 2202 540 2203
rect 638 2207 644 2208
rect 638 2203 639 2207
rect 643 2203 644 2207
rect 638 2202 644 2203
rect 646 2207 652 2208
rect 646 2203 647 2207
rect 651 2203 652 2207
rect 646 2202 652 2203
rect 742 2207 748 2208
rect 742 2203 743 2207
rect 747 2203 748 2207
rect 742 2202 748 2203
rect 750 2207 756 2208
rect 750 2203 751 2207
rect 755 2203 756 2207
rect 750 2202 756 2203
rect 846 2207 852 2208
rect 846 2203 847 2207
rect 851 2203 852 2207
rect 846 2202 852 2203
rect 228 2188 230 2202
rect 238 2199 244 2200
rect 238 2195 239 2199
rect 243 2195 244 2199
rect 238 2194 244 2195
rect 182 2187 188 2188
rect 182 2183 183 2187
rect 187 2183 188 2187
rect 111 2182 115 2183
rect 111 2177 115 2178
rect 159 2182 163 2183
rect 182 2182 188 2183
rect 226 2187 232 2188
rect 226 2183 227 2187
rect 231 2183 232 2187
rect 226 2182 232 2183
rect 159 2177 163 2178
rect 112 2157 114 2177
rect 240 2176 242 2194
rect 248 2183 250 2202
rect 316 2188 318 2202
rect 314 2187 320 2188
rect 314 2183 315 2187
rect 319 2183 320 2187
rect 336 2183 338 2202
rect 412 2188 414 2202
rect 410 2187 416 2188
rect 410 2183 411 2187
rect 415 2183 416 2187
rect 432 2183 434 2202
rect 516 2188 518 2202
rect 514 2187 520 2188
rect 514 2183 515 2187
rect 519 2183 520 2187
rect 536 2183 538 2202
rect 640 2183 642 2202
rect 247 2182 251 2183
rect 247 2177 251 2178
rect 255 2182 259 2183
rect 314 2182 320 2183
rect 335 2182 339 2183
rect 255 2177 259 2178
rect 335 2177 339 2178
rect 351 2182 355 2183
rect 410 2182 416 2183
rect 431 2182 435 2183
rect 351 2177 355 2178
rect 431 2177 435 2178
rect 455 2182 459 2183
rect 514 2182 520 2183
rect 535 2182 539 2183
rect 455 2177 459 2178
rect 535 2177 539 2178
rect 559 2182 563 2183
rect 559 2177 563 2178
rect 639 2182 643 2183
rect 639 2177 643 2178
rect 238 2175 244 2176
rect 238 2171 239 2175
rect 243 2171 244 2175
rect 238 2170 244 2171
rect 256 2158 258 2177
rect 278 2175 284 2176
rect 278 2171 279 2175
rect 283 2171 284 2175
rect 278 2170 284 2171
rect 254 2157 260 2158
rect 110 2156 116 2157
rect 110 2152 111 2156
rect 115 2152 116 2156
rect 254 2153 255 2157
rect 259 2153 260 2157
rect 280 2156 282 2170
rect 352 2158 354 2177
rect 374 2175 380 2176
rect 374 2171 375 2175
rect 379 2171 380 2175
rect 374 2170 380 2171
rect 350 2157 356 2158
rect 254 2152 260 2153
rect 278 2155 284 2156
rect 110 2151 116 2152
rect 278 2151 279 2155
rect 283 2151 284 2155
rect 350 2153 351 2157
rect 355 2153 356 2157
rect 376 2156 378 2170
rect 456 2158 458 2177
rect 478 2175 484 2176
rect 478 2171 479 2175
rect 483 2171 484 2175
rect 478 2170 484 2171
rect 454 2157 460 2158
rect 350 2152 356 2153
rect 374 2155 380 2156
rect 278 2150 284 2151
rect 374 2151 375 2155
rect 379 2151 380 2155
rect 454 2153 455 2157
rect 459 2153 460 2157
rect 480 2156 482 2170
rect 560 2158 562 2177
rect 648 2176 650 2202
rect 744 2183 746 2202
rect 752 2184 754 2202
rect 750 2183 756 2184
rect 848 2183 850 2202
rect 928 2188 930 2254
rect 998 2240 1004 2241
rect 998 2236 999 2240
rect 1003 2236 1004 2240
rect 998 2235 1004 2236
rect 935 2234 939 2235
rect 935 2229 939 2230
rect 999 2234 1003 2235
rect 999 2229 1003 2230
rect 1039 2234 1043 2235
rect 1039 2229 1043 2230
rect 934 2228 940 2229
rect 934 2224 935 2228
rect 939 2224 940 2228
rect 934 2223 940 2224
rect 1038 2228 1044 2229
rect 1038 2224 1039 2228
rect 1043 2224 1044 2228
rect 1038 2223 1044 2224
rect 1076 2208 1078 2266
rect 1128 2262 1130 2281
rect 1150 2279 1156 2280
rect 1150 2275 1151 2279
rect 1155 2275 1156 2279
rect 1150 2274 1156 2275
rect 1126 2261 1132 2262
rect 1126 2257 1127 2261
rect 1131 2257 1132 2261
rect 1152 2260 1154 2274
rect 1240 2262 1242 2281
rect 1238 2261 1244 2262
rect 1126 2256 1132 2257
rect 1150 2259 1156 2260
rect 1150 2255 1151 2259
rect 1155 2255 1156 2259
rect 1238 2257 1239 2261
rect 1243 2257 1244 2261
rect 1260 2260 1262 2294
rect 1288 2287 1290 2315
rect 1326 2312 1332 2313
rect 1784 2312 1786 2378
rect 1792 2374 1794 2393
rect 1790 2373 1796 2374
rect 1790 2369 1791 2373
rect 1795 2369 1796 2373
rect 1812 2372 1814 2402
rect 1832 2399 1834 2422
rect 1896 2399 1898 2422
rect 1948 2408 1950 2422
rect 1946 2407 1952 2408
rect 1946 2403 1947 2407
rect 1951 2403 1952 2407
rect 1946 2402 1952 2403
rect 1968 2399 1970 2422
rect 1831 2398 1835 2399
rect 1831 2393 1835 2394
rect 1855 2398 1859 2399
rect 1855 2393 1859 2394
rect 1895 2398 1899 2399
rect 1895 2393 1899 2394
rect 1919 2398 1923 2399
rect 1919 2393 1923 2394
rect 1967 2398 1971 2399
rect 1967 2393 1971 2394
rect 1856 2374 1858 2393
rect 1920 2374 1922 2393
rect 1976 2392 1978 2422
rect 2040 2399 2042 2422
rect 2056 2400 2058 2422
rect 2054 2399 2060 2400
rect 2112 2399 2114 2422
rect 2184 2399 2186 2422
rect 2192 2408 2194 2478
rect 2502 2467 2508 2468
rect 2502 2463 2503 2467
rect 2507 2463 2508 2467
rect 2502 2462 2508 2463
rect 2504 2455 2506 2462
rect 2503 2454 2507 2455
rect 2503 2449 2507 2450
rect 2504 2446 2506 2449
rect 2502 2445 2508 2446
rect 2502 2441 2503 2445
rect 2507 2441 2508 2445
rect 2502 2440 2508 2441
rect 2502 2428 2508 2429
rect 2502 2424 2503 2428
rect 2507 2424 2508 2428
rect 2502 2423 2508 2424
rect 2190 2407 2196 2408
rect 2190 2403 2191 2407
rect 2195 2403 2196 2407
rect 2190 2402 2196 2403
rect 2504 2399 2506 2423
rect 1983 2398 1987 2399
rect 1983 2393 1987 2394
rect 2039 2398 2043 2399
rect 2039 2393 2043 2394
rect 2047 2398 2051 2399
rect 2054 2395 2055 2399
rect 2059 2395 2060 2399
rect 2054 2394 2060 2395
rect 2111 2398 2115 2399
rect 2047 2393 2051 2394
rect 2111 2393 2115 2394
rect 2183 2398 2187 2399
rect 2183 2393 2187 2394
rect 2503 2398 2507 2399
rect 2503 2393 2507 2394
rect 1974 2391 1980 2392
rect 1974 2387 1975 2391
rect 1979 2387 1980 2391
rect 1974 2386 1980 2387
rect 1984 2374 1986 2393
rect 2006 2391 2012 2392
rect 2006 2387 2007 2391
rect 2011 2387 2012 2391
rect 2006 2386 2012 2387
rect 1854 2373 1860 2374
rect 1790 2368 1796 2369
rect 1810 2371 1816 2372
rect 1810 2367 1811 2371
rect 1815 2367 1816 2371
rect 1854 2369 1855 2373
rect 1859 2369 1860 2373
rect 1918 2373 1924 2374
rect 1854 2368 1860 2369
rect 1862 2371 1868 2372
rect 1810 2366 1816 2367
rect 1862 2367 1863 2371
rect 1867 2367 1868 2371
rect 1918 2369 1919 2373
rect 1923 2369 1924 2373
rect 1918 2368 1924 2369
rect 1982 2373 1988 2374
rect 1982 2369 1983 2373
rect 1987 2369 1988 2373
rect 2008 2372 2010 2386
rect 2048 2374 2050 2393
rect 2070 2391 2076 2392
rect 2070 2387 2071 2391
rect 2075 2387 2076 2391
rect 2070 2386 2076 2387
rect 2046 2373 2052 2374
rect 1982 2368 1988 2369
rect 2006 2371 2012 2372
rect 1862 2366 1868 2367
rect 2006 2367 2007 2371
rect 2011 2367 2012 2371
rect 2046 2369 2047 2373
rect 2051 2369 2052 2373
rect 2072 2372 2074 2386
rect 2112 2374 2114 2393
rect 2110 2373 2116 2374
rect 2504 2373 2506 2393
rect 2046 2368 2052 2369
rect 2070 2371 2076 2372
rect 2006 2366 2012 2367
rect 2070 2367 2071 2371
rect 2075 2367 2076 2371
rect 2110 2369 2111 2373
rect 2115 2369 2116 2373
rect 2110 2368 2116 2369
rect 2502 2372 2508 2373
rect 2502 2368 2503 2372
rect 2507 2368 2508 2372
rect 2502 2367 2508 2368
rect 2070 2366 2076 2367
rect 1838 2352 1844 2353
rect 1838 2348 1839 2352
rect 1843 2348 1844 2352
rect 1838 2347 1844 2348
rect 1840 2339 1842 2347
rect 1831 2338 1835 2339
rect 1831 2333 1835 2334
rect 1839 2338 1843 2339
rect 1839 2333 1843 2334
rect 1830 2332 1836 2333
rect 1830 2328 1831 2332
rect 1835 2328 1836 2332
rect 1830 2327 1836 2328
rect 1326 2308 1327 2312
rect 1331 2308 1332 2312
rect 1326 2307 1332 2308
rect 1486 2311 1492 2312
rect 1486 2307 1487 2311
rect 1491 2307 1492 2311
rect 1328 2287 1330 2307
rect 1486 2306 1492 2307
rect 1530 2311 1536 2312
rect 1530 2307 1531 2311
rect 1535 2307 1536 2311
rect 1530 2306 1536 2307
rect 1550 2311 1556 2312
rect 1550 2307 1551 2311
rect 1555 2307 1556 2311
rect 1550 2306 1556 2307
rect 1602 2311 1608 2312
rect 1602 2307 1603 2311
rect 1607 2307 1608 2311
rect 1602 2306 1608 2307
rect 1622 2311 1628 2312
rect 1622 2307 1623 2311
rect 1627 2307 1628 2311
rect 1622 2306 1628 2307
rect 1678 2311 1684 2312
rect 1678 2307 1679 2311
rect 1683 2307 1684 2311
rect 1678 2306 1684 2307
rect 1702 2311 1708 2312
rect 1702 2307 1703 2311
rect 1707 2307 1708 2311
rect 1702 2306 1708 2307
rect 1754 2311 1760 2312
rect 1754 2307 1755 2311
rect 1759 2307 1760 2311
rect 1754 2306 1760 2307
rect 1774 2311 1780 2312
rect 1774 2307 1775 2311
rect 1779 2307 1780 2311
rect 1774 2306 1780 2307
rect 1782 2311 1788 2312
rect 1782 2307 1783 2311
rect 1787 2307 1788 2311
rect 1782 2306 1788 2307
rect 1846 2311 1852 2312
rect 1846 2307 1847 2311
rect 1851 2307 1852 2311
rect 1846 2306 1852 2307
rect 1488 2287 1490 2306
rect 1532 2292 1534 2306
rect 1522 2291 1528 2292
rect 1522 2287 1523 2291
rect 1527 2287 1528 2291
rect 1287 2286 1291 2287
rect 1287 2281 1291 2282
rect 1327 2286 1331 2287
rect 1327 2281 1331 2282
rect 1383 2286 1387 2287
rect 1383 2281 1387 2282
rect 1479 2286 1483 2287
rect 1479 2281 1483 2282
rect 1487 2286 1491 2287
rect 1522 2286 1528 2287
rect 1530 2291 1536 2292
rect 1530 2287 1531 2291
rect 1535 2287 1536 2291
rect 1552 2287 1554 2306
rect 1604 2292 1606 2306
rect 1602 2291 1608 2292
rect 1602 2287 1603 2291
rect 1607 2287 1608 2291
rect 1624 2287 1626 2306
rect 1680 2292 1682 2306
rect 1678 2291 1684 2292
rect 1678 2287 1679 2291
rect 1683 2287 1684 2291
rect 1704 2287 1706 2306
rect 1756 2292 1758 2306
rect 1754 2291 1760 2292
rect 1754 2287 1755 2291
rect 1759 2287 1760 2291
rect 1776 2287 1778 2306
rect 1848 2287 1850 2306
rect 1864 2292 1866 2366
rect 2502 2355 2508 2356
rect 1902 2352 1908 2353
rect 1902 2348 1903 2352
rect 1907 2348 1908 2352
rect 1902 2347 1908 2348
rect 1966 2352 1972 2353
rect 1966 2348 1967 2352
rect 1971 2348 1972 2352
rect 1966 2347 1972 2348
rect 2030 2352 2036 2353
rect 2030 2348 2031 2352
rect 2035 2348 2036 2352
rect 2030 2347 2036 2348
rect 2094 2352 2100 2353
rect 2094 2348 2095 2352
rect 2099 2348 2100 2352
rect 2502 2351 2503 2355
rect 2507 2351 2508 2355
rect 2502 2350 2508 2351
rect 2094 2347 2100 2348
rect 1904 2339 1906 2347
rect 1968 2339 1970 2347
rect 2032 2339 2034 2347
rect 2096 2339 2098 2347
rect 2504 2339 2506 2350
rect 1903 2338 1907 2339
rect 1903 2333 1907 2334
rect 1967 2338 1971 2339
rect 1967 2333 1971 2334
rect 1983 2338 1987 2339
rect 1983 2333 1987 2334
rect 2031 2338 2035 2339
rect 2031 2333 2035 2334
rect 2063 2338 2067 2339
rect 2063 2333 2067 2334
rect 2095 2338 2099 2339
rect 2095 2333 2099 2334
rect 2143 2338 2147 2339
rect 2143 2333 2147 2334
rect 2503 2338 2507 2339
rect 2503 2333 2507 2334
rect 1902 2332 1908 2333
rect 1902 2328 1903 2332
rect 1907 2328 1908 2332
rect 1902 2327 1908 2328
rect 1982 2332 1988 2333
rect 1982 2328 1983 2332
rect 1987 2328 1988 2332
rect 1982 2327 1988 2328
rect 2062 2332 2068 2333
rect 2062 2328 2063 2332
rect 2067 2328 2068 2332
rect 2062 2327 2068 2328
rect 2142 2332 2148 2333
rect 2142 2328 2143 2332
rect 2147 2328 2148 2332
rect 2504 2330 2506 2333
rect 2142 2327 2148 2328
rect 2502 2329 2508 2330
rect 2502 2325 2503 2329
rect 2507 2325 2508 2329
rect 2502 2324 2508 2325
rect 2502 2312 2508 2313
rect 1894 2311 1900 2312
rect 1894 2307 1895 2311
rect 1899 2307 1900 2311
rect 1894 2306 1900 2307
rect 1918 2311 1924 2312
rect 1918 2307 1919 2311
rect 1923 2307 1924 2311
rect 1918 2306 1924 2307
rect 1978 2311 1984 2312
rect 1978 2307 1979 2311
rect 1983 2307 1984 2311
rect 1978 2306 1984 2307
rect 1998 2311 2004 2312
rect 1998 2307 1999 2311
rect 2003 2307 2004 2311
rect 1998 2306 2004 2307
rect 2058 2311 2064 2312
rect 2058 2307 2059 2311
rect 2063 2307 2064 2311
rect 2058 2306 2064 2307
rect 2078 2311 2084 2312
rect 2078 2307 2079 2311
rect 2083 2307 2084 2311
rect 2078 2306 2084 2307
rect 2138 2311 2144 2312
rect 2138 2307 2139 2311
rect 2143 2307 2144 2311
rect 2138 2306 2144 2307
rect 2158 2311 2164 2312
rect 2158 2307 2159 2311
rect 2163 2307 2164 2311
rect 2502 2308 2503 2312
rect 2507 2308 2508 2312
rect 2502 2307 2508 2308
rect 2158 2306 2164 2307
rect 1886 2303 1892 2304
rect 1886 2299 1887 2303
rect 1891 2299 1892 2303
rect 1886 2298 1892 2299
rect 1862 2291 1868 2292
rect 1862 2287 1863 2291
rect 1867 2287 1868 2291
rect 1530 2286 1536 2287
rect 1551 2286 1555 2287
rect 1487 2281 1491 2282
rect 1288 2261 1290 2281
rect 1328 2261 1330 2281
rect 1384 2262 1386 2281
rect 1398 2279 1404 2280
rect 1398 2275 1399 2279
rect 1403 2275 1404 2279
rect 1398 2274 1404 2275
rect 1406 2279 1412 2280
rect 1406 2275 1407 2279
rect 1411 2275 1412 2279
rect 1406 2274 1412 2275
rect 1382 2261 1388 2262
rect 1286 2260 1292 2261
rect 1238 2256 1244 2257
rect 1258 2259 1264 2260
rect 1150 2254 1156 2255
rect 1258 2255 1259 2259
rect 1263 2255 1264 2259
rect 1286 2256 1287 2260
rect 1291 2256 1292 2260
rect 1286 2255 1292 2256
rect 1326 2260 1332 2261
rect 1326 2256 1327 2260
rect 1331 2256 1332 2260
rect 1382 2257 1383 2261
rect 1387 2257 1388 2261
rect 1382 2256 1388 2257
rect 1326 2255 1332 2256
rect 1258 2254 1264 2255
rect 1286 2243 1292 2244
rect 1110 2240 1116 2241
rect 1110 2236 1111 2240
rect 1115 2236 1116 2240
rect 1110 2235 1116 2236
rect 1222 2240 1228 2241
rect 1222 2236 1223 2240
rect 1227 2236 1228 2240
rect 1286 2239 1287 2243
rect 1291 2239 1292 2243
rect 1286 2238 1292 2239
rect 1326 2243 1332 2244
rect 1326 2239 1327 2243
rect 1331 2239 1332 2243
rect 1326 2238 1332 2239
rect 1366 2240 1372 2241
rect 1222 2235 1228 2236
rect 1288 2235 1290 2238
rect 1328 2235 1330 2238
rect 1366 2236 1367 2240
rect 1371 2236 1372 2240
rect 1366 2235 1372 2236
rect 1111 2234 1115 2235
rect 1111 2229 1115 2230
rect 1143 2234 1147 2235
rect 1143 2229 1147 2230
rect 1223 2234 1227 2235
rect 1223 2229 1227 2230
rect 1287 2234 1291 2235
rect 1287 2229 1291 2230
rect 1327 2234 1331 2235
rect 1327 2229 1331 2230
rect 1367 2234 1371 2235
rect 1367 2229 1371 2230
rect 1142 2228 1148 2229
rect 1142 2224 1143 2228
rect 1147 2224 1148 2228
rect 1142 2223 1148 2224
rect 1222 2228 1228 2229
rect 1222 2224 1223 2228
rect 1227 2224 1228 2228
rect 1288 2226 1290 2229
rect 1328 2226 1330 2229
rect 1366 2228 1372 2229
rect 1222 2223 1228 2224
rect 1286 2225 1292 2226
rect 1286 2221 1287 2225
rect 1291 2221 1292 2225
rect 1286 2220 1292 2221
rect 1326 2225 1332 2226
rect 1326 2221 1327 2225
rect 1331 2221 1332 2225
rect 1366 2224 1367 2228
rect 1371 2224 1372 2228
rect 1366 2223 1372 2224
rect 1326 2220 1332 2221
rect 1286 2208 1292 2209
rect 950 2207 956 2208
rect 950 2203 951 2207
rect 955 2203 956 2207
rect 950 2202 956 2203
rect 1054 2207 1060 2208
rect 1054 2203 1055 2207
rect 1059 2203 1060 2207
rect 1054 2202 1060 2203
rect 1074 2207 1080 2208
rect 1074 2203 1075 2207
rect 1079 2203 1080 2207
rect 1074 2202 1080 2203
rect 1158 2207 1164 2208
rect 1158 2203 1159 2207
rect 1163 2203 1164 2207
rect 1158 2202 1164 2203
rect 1218 2207 1224 2208
rect 1218 2203 1219 2207
rect 1223 2203 1224 2207
rect 1218 2202 1224 2203
rect 1238 2207 1244 2208
rect 1238 2203 1239 2207
rect 1243 2203 1244 2207
rect 1286 2204 1287 2208
rect 1291 2204 1292 2208
rect 1286 2203 1292 2204
rect 1326 2208 1332 2209
rect 1400 2208 1402 2274
rect 1408 2260 1410 2274
rect 1480 2262 1482 2281
rect 1502 2279 1508 2280
rect 1502 2275 1503 2279
rect 1507 2275 1508 2279
rect 1502 2274 1508 2275
rect 1478 2261 1484 2262
rect 1406 2259 1412 2260
rect 1406 2255 1407 2259
rect 1411 2255 1412 2259
rect 1478 2257 1479 2261
rect 1483 2257 1484 2261
rect 1504 2260 1506 2274
rect 1524 2268 1526 2286
rect 1551 2281 1555 2282
rect 1583 2286 1587 2287
rect 1602 2286 1608 2287
rect 1623 2286 1627 2287
rect 1678 2286 1684 2287
rect 1687 2286 1691 2287
rect 1583 2281 1587 2282
rect 1623 2281 1627 2282
rect 1687 2281 1691 2282
rect 1703 2286 1707 2287
rect 1754 2286 1760 2287
rect 1775 2286 1779 2287
rect 1703 2281 1707 2282
rect 1775 2281 1779 2282
rect 1791 2286 1795 2287
rect 1791 2281 1795 2282
rect 1847 2286 1851 2287
rect 1862 2286 1868 2287
rect 1847 2281 1851 2282
rect 1522 2267 1528 2268
rect 1522 2263 1523 2267
rect 1527 2263 1528 2267
rect 1522 2262 1528 2263
rect 1584 2262 1586 2281
rect 1606 2279 1612 2280
rect 1606 2275 1607 2279
rect 1611 2275 1612 2279
rect 1606 2274 1612 2275
rect 1582 2261 1588 2262
rect 1478 2256 1484 2257
rect 1502 2259 1508 2260
rect 1406 2254 1412 2255
rect 1502 2255 1503 2259
rect 1507 2255 1508 2259
rect 1582 2257 1583 2261
rect 1587 2257 1588 2261
rect 1608 2260 1610 2274
rect 1688 2262 1690 2281
rect 1710 2279 1716 2280
rect 1710 2275 1711 2279
rect 1715 2275 1716 2279
rect 1710 2274 1716 2275
rect 1686 2261 1692 2262
rect 1582 2256 1588 2257
rect 1606 2259 1612 2260
rect 1502 2254 1508 2255
rect 1606 2255 1607 2259
rect 1611 2255 1612 2259
rect 1686 2257 1687 2261
rect 1691 2257 1692 2261
rect 1712 2260 1714 2274
rect 1792 2262 1794 2281
rect 1888 2280 1890 2298
rect 1896 2292 1898 2306
rect 1894 2291 1900 2292
rect 1894 2287 1895 2291
rect 1899 2287 1900 2291
rect 1920 2287 1922 2306
rect 1980 2292 1982 2306
rect 1978 2291 1984 2292
rect 1978 2287 1979 2291
rect 1983 2287 1984 2291
rect 2000 2287 2002 2306
rect 2060 2292 2062 2306
rect 2058 2291 2064 2292
rect 2058 2287 2059 2291
rect 2063 2287 2064 2291
rect 2080 2287 2082 2306
rect 2140 2292 2142 2306
rect 2138 2291 2144 2292
rect 2138 2287 2139 2291
rect 2143 2287 2144 2291
rect 2160 2287 2162 2306
rect 2504 2287 2506 2307
rect 1894 2286 1900 2287
rect 1903 2286 1907 2287
rect 1903 2281 1907 2282
rect 1919 2286 1923 2287
rect 1978 2286 1984 2287
rect 1999 2286 2003 2287
rect 1919 2281 1923 2282
rect 1999 2281 2003 2282
rect 2015 2286 2019 2287
rect 2058 2286 2064 2287
rect 2079 2286 2083 2287
rect 2015 2281 2019 2282
rect 2079 2281 2083 2282
rect 2127 2286 2131 2287
rect 2138 2286 2144 2287
rect 2159 2286 2163 2287
rect 2127 2281 2131 2282
rect 2159 2281 2163 2282
rect 2239 2286 2243 2287
rect 2239 2281 2243 2282
rect 2503 2286 2507 2287
rect 2503 2281 2507 2282
rect 1886 2279 1892 2280
rect 1886 2275 1887 2279
rect 1891 2275 1892 2279
rect 1886 2274 1892 2275
rect 1904 2262 1906 2281
rect 1926 2279 1932 2280
rect 1926 2275 1927 2279
rect 1931 2275 1932 2279
rect 1926 2274 1932 2275
rect 1790 2261 1796 2262
rect 1686 2256 1692 2257
rect 1710 2259 1716 2260
rect 1606 2254 1612 2255
rect 1710 2255 1711 2259
rect 1715 2255 1716 2259
rect 1790 2257 1791 2261
rect 1795 2257 1796 2261
rect 1790 2256 1796 2257
rect 1902 2261 1908 2262
rect 1902 2257 1903 2261
rect 1907 2257 1908 2261
rect 1928 2260 1930 2274
rect 2016 2262 2018 2281
rect 2038 2279 2044 2280
rect 2038 2275 2039 2279
rect 2043 2275 2044 2279
rect 2038 2274 2044 2275
rect 2014 2261 2020 2262
rect 1902 2256 1908 2257
rect 1926 2259 1932 2260
rect 1710 2254 1716 2255
rect 1926 2255 1927 2259
rect 1931 2255 1932 2259
rect 2014 2257 2015 2261
rect 2019 2257 2020 2261
rect 2040 2260 2042 2274
rect 2128 2262 2130 2281
rect 2150 2279 2156 2280
rect 2150 2275 2151 2279
rect 2155 2275 2156 2279
rect 2150 2274 2156 2275
rect 2126 2261 2132 2262
rect 2014 2256 2020 2257
rect 2038 2259 2044 2260
rect 1926 2254 1932 2255
rect 2038 2255 2039 2259
rect 2043 2255 2044 2259
rect 2126 2257 2127 2261
rect 2131 2257 2132 2261
rect 2152 2260 2154 2274
rect 2240 2262 2242 2281
rect 2238 2261 2244 2262
rect 2504 2261 2506 2281
rect 2126 2256 2132 2257
rect 2150 2259 2156 2260
rect 2038 2254 2044 2255
rect 2150 2255 2151 2259
rect 2155 2255 2156 2259
rect 2238 2257 2239 2261
rect 2243 2257 2244 2261
rect 2502 2260 2508 2261
rect 2238 2256 2244 2257
rect 2246 2259 2252 2260
rect 2150 2254 2156 2255
rect 2246 2255 2247 2259
rect 2251 2255 2252 2259
rect 2502 2256 2503 2260
rect 2507 2256 2508 2260
rect 2502 2255 2508 2256
rect 2246 2254 2252 2255
rect 1462 2240 1468 2241
rect 1462 2236 1463 2240
rect 1467 2236 1468 2240
rect 1462 2235 1468 2236
rect 1566 2240 1572 2241
rect 1566 2236 1567 2240
rect 1571 2236 1572 2240
rect 1566 2235 1572 2236
rect 1670 2240 1676 2241
rect 1670 2236 1671 2240
rect 1675 2236 1676 2240
rect 1670 2235 1676 2236
rect 1774 2240 1780 2241
rect 1774 2236 1775 2240
rect 1779 2236 1780 2240
rect 1774 2235 1780 2236
rect 1886 2240 1892 2241
rect 1886 2236 1887 2240
rect 1891 2236 1892 2240
rect 1886 2235 1892 2236
rect 1998 2240 2004 2241
rect 1998 2236 1999 2240
rect 2003 2236 2004 2240
rect 1998 2235 2004 2236
rect 2110 2240 2116 2241
rect 2110 2236 2111 2240
rect 2115 2236 2116 2240
rect 2110 2235 2116 2236
rect 2222 2240 2228 2241
rect 2222 2236 2223 2240
rect 2227 2236 2228 2240
rect 2222 2235 2228 2236
rect 1463 2234 1467 2235
rect 1463 2229 1467 2230
rect 1487 2234 1491 2235
rect 1487 2229 1491 2230
rect 1567 2234 1571 2235
rect 1567 2229 1571 2230
rect 1607 2234 1611 2235
rect 1607 2229 1611 2230
rect 1671 2234 1675 2235
rect 1671 2229 1675 2230
rect 1719 2234 1723 2235
rect 1719 2229 1723 2230
rect 1775 2234 1779 2235
rect 1775 2229 1779 2230
rect 1815 2234 1819 2235
rect 1815 2229 1819 2230
rect 1887 2234 1891 2235
rect 1887 2229 1891 2230
rect 1903 2234 1907 2235
rect 1903 2229 1907 2230
rect 1983 2234 1987 2235
rect 1983 2229 1987 2230
rect 1999 2234 2003 2235
rect 1999 2229 2003 2230
rect 2055 2234 2059 2235
rect 2055 2229 2059 2230
rect 2111 2234 2115 2235
rect 2111 2229 2115 2230
rect 2127 2234 2131 2235
rect 2127 2229 2131 2230
rect 2191 2234 2195 2235
rect 2191 2229 2195 2230
rect 2223 2234 2227 2235
rect 2223 2229 2227 2230
rect 1486 2228 1492 2229
rect 1486 2224 1487 2228
rect 1491 2224 1492 2228
rect 1486 2223 1492 2224
rect 1606 2228 1612 2229
rect 1606 2224 1607 2228
rect 1611 2224 1612 2228
rect 1606 2223 1612 2224
rect 1718 2228 1724 2229
rect 1718 2224 1719 2228
rect 1723 2224 1724 2228
rect 1718 2223 1724 2224
rect 1814 2228 1820 2229
rect 1814 2224 1815 2228
rect 1819 2224 1820 2228
rect 1814 2223 1820 2224
rect 1902 2228 1908 2229
rect 1902 2224 1903 2228
rect 1907 2224 1908 2228
rect 1902 2223 1908 2224
rect 1982 2228 1988 2229
rect 1982 2224 1983 2228
rect 1987 2224 1988 2228
rect 1982 2223 1988 2224
rect 2054 2228 2060 2229
rect 2054 2224 2055 2228
rect 2059 2224 2060 2228
rect 2054 2223 2060 2224
rect 2126 2228 2132 2229
rect 2126 2224 2127 2228
rect 2131 2224 2132 2228
rect 2126 2223 2132 2224
rect 2190 2228 2196 2229
rect 2190 2224 2191 2228
rect 2195 2224 2196 2228
rect 2190 2223 2196 2224
rect 2248 2221 2250 2254
rect 2502 2243 2508 2244
rect 2502 2239 2503 2243
rect 2507 2239 2508 2243
rect 2502 2238 2508 2239
rect 2504 2235 2506 2238
rect 2255 2234 2259 2235
rect 2255 2229 2259 2230
rect 2319 2234 2323 2235
rect 2319 2229 2323 2230
rect 2383 2234 2387 2235
rect 2383 2229 2387 2230
rect 2439 2234 2443 2235
rect 2439 2229 2443 2230
rect 2503 2234 2507 2235
rect 2503 2229 2507 2230
rect 2254 2228 2260 2229
rect 2254 2224 2255 2228
rect 2259 2224 2260 2228
rect 2254 2223 2260 2224
rect 2318 2228 2324 2229
rect 2318 2224 2319 2228
rect 2323 2224 2324 2228
rect 2318 2223 2324 2224
rect 2382 2228 2388 2229
rect 2382 2224 2383 2228
rect 2387 2224 2388 2228
rect 2382 2223 2388 2224
rect 2438 2228 2444 2229
rect 2438 2224 2439 2228
rect 2443 2224 2444 2228
rect 2504 2226 2506 2229
rect 2438 2223 2444 2224
rect 2502 2225 2508 2226
rect 2502 2221 2503 2225
rect 2507 2221 2508 2225
rect 1719 2220 1723 2221
rect 1719 2215 1723 2216
rect 2247 2220 2251 2221
rect 2502 2220 2508 2221
rect 2247 2215 2251 2216
rect 1326 2204 1327 2208
rect 1331 2204 1332 2208
rect 1326 2203 1332 2204
rect 1382 2207 1388 2208
rect 1382 2203 1383 2207
rect 1387 2203 1388 2207
rect 1238 2202 1244 2203
rect 926 2187 932 2188
rect 926 2183 927 2187
rect 931 2183 932 2187
rect 952 2183 954 2202
rect 1056 2183 1058 2202
rect 1078 2187 1084 2188
rect 1078 2183 1079 2187
rect 1083 2183 1084 2187
rect 1160 2183 1162 2202
rect 1220 2188 1222 2202
rect 1218 2187 1224 2188
rect 1218 2183 1219 2187
rect 1223 2183 1224 2187
rect 1240 2183 1242 2202
rect 1288 2183 1290 2203
rect 663 2182 667 2183
rect 663 2177 667 2178
rect 743 2182 747 2183
rect 750 2179 751 2183
rect 755 2179 756 2183
rect 750 2178 756 2179
rect 767 2182 771 2183
rect 743 2177 747 2178
rect 767 2177 771 2178
rect 847 2182 851 2183
rect 847 2177 851 2178
rect 863 2182 867 2183
rect 926 2182 932 2183
rect 951 2182 955 2183
rect 863 2177 867 2178
rect 951 2177 955 2178
rect 959 2182 963 2183
rect 959 2177 963 2178
rect 1055 2182 1059 2183
rect 1078 2182 1084 2183
rect 1159 2182 1163 2183
rect 1218 2182 1224 2183
rect 1239 2182 1243 2183
rect 1055 2177 1059 2178
rect 646 2175 652 2176
rect 646 2171 647 2175
rect 651 2171 652 2175
rect 646 2170 652 2171
rect 664 2158 666 2177
rect 686 2175 692 2176
rect 686 2171 687 2175
rect 691 2171 692 2175
rect 686 2170 692 2171
rect 558 2157 564 2158
rect 454 2152 460 2153
rect 478 2155 484 2156
rect 374 2150 380 2151
rect 478 2151 479 2155
rect 483 2151 484 2155
rect 558 2153 559 2157
rect 563 2153 564 2157
rect 662 2157 668 2158
rect 558 2152 564 2153
rect 566 2155 572 2156
rect 478 2150 484 2151
rect 566 2151 567 2155
rect 571 2151 572 2155
rect 662 2153 663 2157
rect 667 2153 668 2157
rect 688 2156 690 2170
rect 768 2158 770 2177
rect 790 2175 796 2176
rect 790 2171 791 2175
rect 795 2171 796 2175
rect 790 2170 796 2171
rect 766 2157 772 2158
rect 662 2152 668 2153
rect 686 2155 692 2156
rect 566 2150 572 2151
rect 686 2151 687 2155
rect 691 2151 692 2155
rect 766 2153 767 2157
rect 771 2153 772 2157
rect 792 2156 794 2170
rect 864 2158 866 2177
rect 886 2175 892 2176
rect 886 2171 887 2175
rect 891 2171 892 2175
rect 886 2170 892 2171
rect 862 2157 868 2158
rect 766 2152 772 2153
rect 790 2155 796 2156
rect 686 2150 692 2151
rect 790 2151 791 2155
rect 795 2151 796 2155
rect 862 2153 863 2157
rect 867 2153 868 2157
rect 888 2156 890 2170
rect 960 2158 962 2177
rect 1056 2158 1058 2177
rect 958 2157 964 2158
rect 862 2152 868 2153
rect 886 2155 892 2156
rect 790 2150 796 2151
rect 886 2151 887 2155
rect 891 2151 892 2155
rect 958 2153 959 2157
rect 963 2153 964 2157
rect 1054 2157 1060 2158
rect 958 2152 964 2153
rect 982 2155 988 2156
rect 886 2150 892 2151
rect 982 2151 983 2155
rect 987 2151 988 2155
rect 1054 2153 1055 2157
rect 1059 2153 1060 2157
rect 1080 2156 1082 2182
rect 1159 2177 1163 2178
rect 1239 2177 1243 2178
rect 1287 2182 1291 2183
rect 1287 2177 1291 2178
rect 1160 2158 1162 2177
rect 1240 2158 1242 2177
rect 1258 2175 1264 2176
rect 1258 2171 1259 2175
rect 1263 2171 1264 2175
rect 1258 2170 1264 2171
rect 1158 2157 1164 2158
rect 1054 2152 1060 2153
rect 1078 2155 1084 2156
rect 982 2150 988 2151
rect 1078 2151 1079 2155
rect 1083 2151 1084 2155
rect 1158 2153 1159 2157
rect 1163 2153 1164 2157
rect 1158 2152 1164 2153
rect 1238 2157 1244 2158
rect 1238 2153 1239 2157
rect 1243 2153 1244 2157
rect 1238 2152 1244 2153
rect 1078 2150 1084 2151
rect 110 2139 116 2140
rect 110 2135 111 2139
rect 115 2135 116 2139
rect 110 2134 116 2135
rect 238 2136 244 2137
rect 112 2131 114 2134
rect 238 2132 239 2136
rect 243 2132 244 2136
rect 238 2131 244 2132
rect 334 2136 340 2137
rect 334 2132 335 2136
rect 339 2132 340 2136
rect 334 2131 340 2132
rect 438 2136 444 2137
rect 438 2132 439 2136
rect 443 2132 444 2136
rect 438 2131 444 2132
rect 542 2136 548 2137
rect 542 2132 543 2136
rect 547 2132 548 2136
rect 542 2131 548 2132
rect 111 2130 115 2131
rect 111 2125 115 2126
rect 239 2130 243 2131
rect 239 2125 243 2126
rect 303 2130 307 2131
rect 303 2125 307 2126
rect 335 2130 339 2131
rect 335 2125 339 2126
rect 359 2130 363 2131
rect 359 2125 363 2126
rect 423 2130 427 2131
rect 423 2125 427 2126
rect 439 2130 443 2131
rect 439 2125 443 2126
rect 487 2130 491 2131
rect 487 2125 491 2126
rect 543 2130 547 2131
rect 543 2125 547 2126
rect 559 2130 563 2131
rect 559 2125 563 2126
rect 112 2122 114 2125
rect 302 2124 308 2125
rect 110 2121 116 2122
rect 110 2117 111 2121
rect 115 2117 116 2121
rect 302 2120 303 2124
rect 307 2120 308 2124
rect 302 2119 308 2120
rect 358 2124 364 2125
rect 358 2120 359 2124
rect 363 2120 364 2124
rect 358 2119 364 2120
rect 422 2124 428 2125
rect 422 2120 423 2124
rect 427 2120 428 2124
rect 422 2119 428 2120
rect 486 2124 492 2125
rect 486 2120 487 2124
rect 491 2120 492 2124
rect 486 2119 492 2120
rect 558 2124 564 2125
rect 558 2120 559 2124
rect 563 2120 564 2124
rect 558 2119 564 2120
rect 110 2116 116 2117
rect 110 2104 116 2105
rect 110 2100 111 2104
rect 115 2100 116 2104
rect 110 2099 116 2100
rect 318 2103 324 2104
rect 318 2099 319 2103
rect 323 2099 324 2103
rect 112 2075 114 2099
rect 318 2098 324 2099
rect 354 2103 360 2104
rect 354 2099 355 2103
rect 359 2099 360 2103
rect 354 2098 360 2099
rect 374 2103 380 2104
rect 374 2099 375 2103
rect 379 2099 380 2103
rect 374 2098 380 2099
rect 418 2103 424 2104
rect 418 2099 419 2103
rect 423 2099 424 2103
rect 418 2098 424 2099
rect 438 2103 444 2104
rect 438 2099 439 2103
rect 443 2099 444 2103
rect 438 2098 444 2099
rect 482 2103 488 2104
rect 482 2099 483 2103
rect 487 2099 488 2103
rect 482 2098 488 2099
rect 502 2103 508 2104
rect 502 2099 503 2103
rect 507 2099 508 2103
rect 502 2098 508 2099
rect 554 2103 560 2104
rect 554 2099 555 2103
rect 559 2099 560 2103
rect 554 2098 560 2099
rect 320 2075 322 2098
rect 356 2084 358 2098
rect 354 2083 360 2084
rect 354 2079 355 2083
rect 359 2079 360 2083
rect 354 2078 360 2079
rect 376 2075 378 2098
rect 420 2084 422 2098
rect 418 2083 424 2084
rect 418 2079 419 2083
rect 423 2079 424 2083
rect 418 2078 424 2079
rect 440 2075 442 2098
rect 484 2084 486 2098
rect 482 2083 488 2084
rect 482 2079 483 2083
rect 487 2079 488 2083
rect 482 2078 488 2079
rect 474 2075 480 2076
rect 504 2075 506 2098
rect 556 2084 558 2098
rect 568 2092 570 2150
rect 646 2136 652 2137
rect 646 2132 647 2136
rect 651 2132 652 2136
rect 646 2131 652 2132
rect 750 2136 756 2137
rect 750 2132 751 2136
rect 755 2132 756 2136
rect 750 2131 756 2132
rect 846 2136 852 2137
rect 846 2132 847 2136
rect 851 2132 852 2136
rect 846 2131 852 2132
rect 942 2136 948 2137
rect 942 2132 943 2136
rect 947 2132 948 2136
rect 942 2131 948 2132
rect 631 2130 635 2131
rect 631 2125 635 2126
rect 647 2130 651 2131
rect 647 2125 651 2126
rect 711 2130 715 2131
rect 711 2125 715 2126
rect 751 2130 755 2131
rect 751 2125 755 2126
rect 799 2130 803 2131
rect 799 2125 803 2126
rect 847 2130 851 2131
rect 847 2125 851 2126
rect 887 2130 891 2131
rect 887 2125 891 2126
rect 943 2130 947 2131
rect 943 2125 947 2126
rect 975 2130 979 2131
rect 975 2125 979 2126
rect 630 2124 636 2125
rect 630 2120 631 2124
rect 635 2120 636 2124
rect 630 2119 636 2120
rect 710 2124 716 2125
rect 710 2120 711 2124
rect 715 2120 716 2124
rect 710 2119 716 2120
rect 798 2124 804 2125
rect 798 2120 799 2124
rect 803 2120 804 2124
rect 798 2119 804 2120
rect 886 2124 892 2125
rect 886 2120 887 2124
rect 891 2120 892 2124
rect 886 2119 892 2120
rect 974 2124 980 2125
rect 974 2120 975 2124
rect 979 2120 980 2124
rect 974 2119 980 2120
rect 574 2103 580 2104
rect 574 2099 575 2103
rect 579 2099 580 2103
rect 574 2098 580 2099
rect 626 2103 632 2104
rect 626 2099 627 2103
rect 631 2099 632 2103
rect 626 2098 632 2099
rect 646 2103 652 2104
rect 646 2099 647 2103
rect 651 2099 652 2103
rect 646 2098 652 2099
rect 654 2103 660 2104
rect 654 2099 655 2103
rect 659 2099 660 2103
rect 654 2098 660 2099
rect 726 2103 732 2104
rect 726 2099 727 2103
rect 731 2099 732 2103
rect 726 2098 732 2099
rect 794 2103 800 2104
rect 794 2099 795 2103
rect 799 2099 800 2103
rect 794 2098 800 2099
rect 814 2103 820 2104
rect 814 2099 815 2103
rect 819 2099 820 2103
rect 814 2098 820 2099
rect 838 2103 844 2104
rect 838 2099 839 2103
rect 843 2099 844 2103
rect 838 2098 844 2099
rect 902 2103 908 2104
rect 902 2099 903 2103
rect 907 2099 908 2103
rect 902 2098 908 2099
rect 566 2091 572 2092
rect 566 2087 567 2091
rect 571 2087 572 2091
rect 566 2086 572 2087
rect 554 2083 560 2084
rect 554 2079 555 2083
rect 559 2079 560 2083
rect 554 2078 560 2079
rect 576 2075 578 2098
rect 628 2084 630 2098
rect 626 2083 632 2084
rect 626 2079 627 2083
rect 631 2079 632 2083
rect 626 2078 632 2079
rect 648 2075 650 2098
rect 111 2074 115 2075
rect 111 2069 115 2070
rect 319 2074 323 2075
rect 319 2069 323 2070
rect 375 2074 379 2075
rect 375 2069 379 2070
rect 399 2074 403 2075
rect 399 2069 403 2070
rect 439 2074 443 2075
rect 439 2069 443 2070
rect 455 2074 459 2075
rect 474 2071 475 2075
rect 479 2071 480 2075
rect 474 2070 480 2071
rect 503 2074 507 2075
rect 455 2069 459 2070
rect 112 2049 114 2069
rect 400 2050 402 2069
rect 456 2050 458 2069
rect 398 2049 404 2050
rect 110 2048 116 2049
rect 110 2044 111 2048
rect 115 2044 116 2048
rect 398 2045 399 2049
rect 403 2045 404 2049
rect 454 2049 460 2050
rect 398 2044 404 2045
rect 430 2047 436 2048
rect 110 2043 116 2044
rect 430 2043 431 2047
rect 435 2043 436 2047
rect 454 2045 455 2049
rect 459 2045 460 2049
rect 476 2048 478 2070
rect 503 2069 507 2070
rect 511 2074 515 2075
rect 511 2069 515 2070
rect 575 2074 579 2075
rect 575 2069 579 2070
rect 639 2074 643 2075
rect 639 2069 643 2070
rect 647 2074 651 2075
rect 647 2069 651 2070
rect 512 2050 514 2069
rect 576 2050 578 2069
rect 640 2050 642 2069
rect 656 2068 658 2098
rect 728 2075 730 2098
rect 796 2084 798 2098
rect 794 2083 800 2084
rect 794 2079 795 2083
rect 799 2079 800 2083
rect 794 2078 800 2079
rect 816 2075 818 2098
rect 711 2074 715 2075
rect 711 2069 715 2070
rect 727 2074 731 2075
rect 727 2069 731 2070
rect 791 2074 795 2075
rect 791 2069 795 2070
rect 815 2074 819 2075
rect 815 2069 819 2070
rect 654 2067 660 2068
rect 654 2063 655 2067
rect 659 2063 660 2067
rect 654 2062 660 2063
rect 712 2050 714 2069
rect 792 2050 794 2069
rect 840 2068 842 2098
rect 904 2075 906 2098
rect 984 2084 986 2150
rect 1038 2136 1044 2137
rect 1038 2132 1039 2136
rect 1043 2132 1044 2136
rect 1038 2131 1044 2132
rect 1142 2136 1148 2137
rect 1142 2132 1143 2136
rect 1147 2132 1148 2136
rect 1142 2131 1148 2132
rect 1222 2136 1228 2137
rect 1222 2132 1223 2136
rect 1227 2132 1228 2136
rect 1222 2131 1228 2132
rect 1039 2130 1043 2131
rect 1039 2125 1043 2126
rect 1063 2130 1067 2131
rect 1063 2125 1067 2126
rect 1143 2130 1147 2131
rect 1143 2125 1147 2126
rect 1151 2130 1155 2131
rect 1151 2125 1155 2126
rect 1223 2130 1227 2131
rect 1223 2125 1227 2126
rect 1062 2124 1068 2125
rect 1062 2120 1063 2124
rect 1067 2120 1068 2124
rect 1062 2119 1068 2120
rect 1150 2124 1156 2125
rect 1150 2120 1151 2124
rect 1155 2120 1156 2124
rect 1150 2119 1156 2120
rect 1222 2124 1228 2125
rect 1222 2120 1223 2124
rect 1227 2120 1228 2124
rect 1222 2119 1228 2120
rect 1260 2104 1262 2170
rect 1288 2157 1290 2177
rect 1328 2163 1330 2203
rect 1382 2202 1388 2203
rect 1398 2207 1404 2208
rect 1398 2203 1399 2207
rect 1403 2203 1404 2207
rect 1398 2202 1404 2203
rect 1502 2207 1508 2208
rect 1502 2203 1503 2207
rect 1507 2203 1508 2207
rect 1502 2202 1508 2203
rect 1602 2207 1608 2208
rect 1602 2203 1603 2207
rect 1607 2203 1608 2207
rect 1602 2202 1608 2203
rect 1622 2207 1628 2208
rect 1622 2203 1623 2207
rect 1627 2203 1628 2207
rect 1622 2202 1628 2203
rect 1384 2163 1386 2202
rect 1430 2187 1436 2188
rect 1430 2183 1431 2187
rect 1435 2183 1436 2187
rect 1430 2182 1436 2183
rect 1327 2162 1331 2163
rect 1327 2157 1331 2158
rect 1383 2162 1387 2163
rect 1383 2157 1387 2158
rect 1407 2162 1411 2163
rect 1407 2157 1411 2158
rect 1286 2156 1292 2157
rect 1286 2152 1287 2156
rect 1291 2152 1292 2156
rect 1286 2151 1292 2152
rect 1286 2139 1292 2140
rect 1286 2135 1287 2139
rect 1291 2135 1292 2139
rect 1328 2137 1330 2157
rect 1408 2138 1410 2157
rect 1406 2137 1412 2138
rect 1286 2134 1292 2135
rect 1326 2136 1332 2137
rect 1288 2131 1290 2134
rect 1326 2132 1327 2136
rect 1331 2132 1332 2136
rect 1406 2133 1407 2137
rect 1411 2133 1412 2137
rect 1432 2136 1434 2182
rect 1504 2163 1506 2202
rect 1604 2188 1606 2202
rect 1602 2187 1608 2188
rect 1602 2183 1603 2187
rect 1607 2183 1608 2187
rect 1602 2182 1608 2183
rect 1624 2163 1626 2202
rect 1720 2188 1722 2215
rect 2502 2208 2508 2209
rect 1734 2207 1740 2208
rect 1734 2203 1735 2207
rect 1739 2203 1740 2207
rect 1734 2202 1740 2203
rect 1810 2207 1816 2208
rect 1810 2203 1811 2207
rect 1815 2203 1816 2207
rect 1810 2202 1816 2203
rect 1830 2207 1836 2208
rect 1830 2203 1831 2207
rect 1835 2203 1836 2207
rect 1830 2202 1836 2203
rect 1898 2207 1904 2208
rect 1898 2203 1899 2207
rect 1903 2203 1904 2207
rect 1898 2202 1904 2203
rect 1918 2207 1924 2208
rect 1918 2203 1919 2207
rect 1923 2203 1924 2207
rect 1918 2202 1924 2203
rect 1978 2207 1984 2208
rect 1978 2203 1979 2207
rect 1983 2203 1984 2207
rect 1978 2202 1984 2203
rect 1998 2207 2004 2208
rect 1998 2203 1999 2207
rect 2003 2203 2004 2207
rect 1998 2202 2004 2203
rect 2050 2207 2056 2208
rect 2050 2203 2051 2207
rect 2055 2203 2056 2207
rect 2050 2202 2056 2203
rect 2070 2207 2076 2208
rect 2070 2203 2071 2207
rect 2075 2203 2076 2207
rect 2070 2202 2076 2203
rect 2122 2207 2128 2208
rect 2122 2203 2123 2207
rect 2127 2203 2128 2207
rect 2122 2202 2128 2203
rect 2142 2207 2148 2208
rect 2142 2203 2143 2207
rect 2147 2203 2148 2207
rect 2142 2202 2148 2203
rect 2186 2207 2192 2208
rect 2186 2203 2187 2207
rect 2191 2203 2192 2207
rect 2186 2202 2192 2203
rect 2206 2207 2212 2208
rect 2206 2203 2207 2207
rect 2211 2203 2212 2207
rect 2206 2202 2212 2203
rect 2250 2207 2256 2208
rect 2250 2203 2251 2207
rect 2255 2203 2256 2207
rect 2250 2202 2256 2203
rect 2270 2207 2276 2208
rect 2270 2203 2271 2207
rect 2275 2203 2276 2207
rect 2270 2202 2276 2203
rect 2314 2207 2320 2208
rect 2314 2203 2315 2207
rect 2319 2203 2320 2207
rect 2314 2202 2320 2203
rect 2334 2207 2340 2208
rect 2334 2203 2335 2207
rect 2339 2203 2340 2207
rect 2334 2202 2340 2203
rect 2378 2207 2384 2208
rect 2378 2203 2379 2207
rect 2383 2203 2384 2207
rect 2378 2202 2384 2203
rect 2398 2207 2404 2208
rect 2398 2203 2399 2207
rect 2403 2203 2404 2207
rect 2398 2202 2404 2203
rect 2434 2207 2440 2208
rect 2434 2203 2435 2207
rect 2439 2203 2440 2207
rect 2434 2202 2440 2203
rect 2454 2207 2460 2208
rect 2454 2203 2455 2207
rect 2459 2203 2460 2207
rect 2454 2202 2460 2203
rect 2462 2207 2468 2208
rect 2462 2203 2463 2207
rect 2467 2203 2468 2207
rect 2502 2204 2503 2208
rect 2507 2204 2508 2208
rect 2502 2203 2508 2204
rect 2462 2202 2468 2203
rect 1718 2187 1724 2188
rect 1718 2183 1719 2187
rect 1723 2183 1724 2187
rect 1718 2182 1724 2183
rect 1736 2163 1738 2202
rect 1812 2188 1814 2202
rect 1810 2187 1816 2188
rect 1810 2183 1811 2187
rect 1815 2183 1816 2187
rect 1810 2182 1816 2183
rect 1832 2163 1834 2202
rect 1900 2188 1902 2202
rect 1898 2187 1904 2188
rect 1898 2183 1899 2187
rect 1903 2183 1904 2187
rect 1898 2182 1904 2183
rect 1920 2163 1922 2202
rect 1980 2188 1982 2202
rect 1978 2187 1984 2188
rect 1978 2183 1979 2187
rect 1983 2183 1984 2187
rect 1978 2182 1984 2183
rect 2000 2163 2002 2202
rect 2052 2188 2054 2202
rect 2050 2187 2056 2188
rect 2050 2183 2051 2187
rect 2055 2183 2056 2187
rect 2050 2182 2056 2183
rect 2072 2163 2074 2202
rect 2124 2188 2126 2202
rect 2122 2187 2128 2188
rect 2122 2183 2123 2187
rect 2127 2183 2128 2187
rect 2122 2182 2128 2183
rect 2144 2163 2146 2202
rect 2188 2188 2190 2202
rect 2186 2187 2192 2188
rect 2186 2183 2187 2187
rect 2191 2183 2192 2187
rect 2186 2182 2192 2183
rect 2208 2163 2210 2202
rect 2252 2188 2254 2202
rect 2250 2187 2256 2188
rect 2250 2183 2251 2187
rect 2255 2183 2256 2187
rect 2250 2182 2256 2183
rect 2272 2163 2274 2202
rect 2316 2188 2318 2202
rect 2314 2187 2320 2188
rect 2314 2183 2315 2187
rect 2319 2183 2320 2187
rect 2314 2182 2320 2183
rect 2336 2163 2338 2202
rect 2380 2188 2382 2202
rect 2378 2187 2384 2188
rect 2378 2183 2379 2187
rect 2383 2183 2384 2187
rect 2378 2182 2384 2183
rect 2400 2163 2402 2202
rect 2436 2188 2438 2202
rect 2434 2187 2440 2188
rect 2434 2183 2435 2187
rect 2439 2183 2440 2187
rect 2434 2182 2440 2183
rect 2456 2163 2458 2202
rect 1503 2162 1507 2163
rect 1503 2157 1507 2158
rect 1623 2162 1627 2163
rect 1623 2157 1627 2158
rect 1735 2162 1739 2163
rect 1735 2157 1739 2158
rect 1815 2162 1819 2163
rect 1815 2157 1819 2158
rect 1831 2162 1835 2163
rect 1831 2157 1835 2158
rect 1919 2162 1923 2163
rect 1919 2157 1923 2158
rect 1991 2162 1995 2163
rect 1991 2157 1995 2158
rect 1999 2162 2003 2163
rect 1999 2157 2003 2158
rect 2071 2162 2075 2163
rect 2071 2157 2075 2158
rect 2143 2162 2147 2163
rect 2143 2157 2147 2158
rect 2159 2162 2163 2163
rect 2159 2157 2163 2158
rect 2207 2162 2211 2163
rect 2207 2157 2211 2158
rect 2271 2162 2275 2163
rect 2271 2157 2275 2158
rect 2319 2162 2323 2163
rect 2319 2157 2323 2158
rect 2335 2162 2339 2163
rect 2335 2157 2339 2158
rect 2399 2162 2403 2163
rect 2399 2157 2403 2158
rect 2455 2162 2459 2163
rect 2455 2157 2459 2158
rect 1624 2138 1626 2157
rect 1746 2155 1752 2156
rect 1746 2151 1747 2155
rect 1751 2151 1752 2155
rect 1746 2150 1752 2151
rect 1622 2137 1628 2138
rect 1406 2132 1412 2133
rect 1430 2135 1436 2136
rect 1326 2131 1332 2132
rect 1430 2131 1431 2135
rect 1435 2131 1436 2135
rect 1622 2133 1623 2137
rect 1627 2133 1628 2137
rect 1622 2132 1628 2133
rect 1287 2130 1291 2131
rect 1430 2130 1436 2131
rect 1287 2125 1291 2126
rect 1288 2122 1290 2125
rect 1286 2121 1292 2122
rect 1286 2117 1287 2121
rect 1291 2117 1292 2121
rect 1286 2116 1292 2117
rect 1326 2119 1332 2120
rect 1326 2115 1327 2119
rect 1331 2115 1332 2119
rect 1326 2114 1332 2115
rect 1390 2116 1396 2117
rect 1328 2111 1330 2114
rect 1390 2112 1391 2116
rect 1395 2112 1396 2116
rect 1390 2111 1396 2112
rect 1606 2116 1612 2117
rect 1606 2112 1607 2116
rect 1611 2112 1612 2116
rect 1606 2111 1612 2112
rect 1327 2110 1331 2111
rect 1327 2105 1331 2106
rect 1383 2110 1387 2111
rect 1383 2105 1387 2106
rect 1391 2110 1395 2111
rect 1391 2105 1395 2106
rect 1551 2110 1555 2111
rect 1551 2105 1555 2106
rect 1607 2110 1611 2111
rect 1607 2105 1611 2106
rect 1711 2110 1715 2111
rect 1711 2105 1715 2106
rect 1286 2104 1292 2105
rect 990 2103 996 2104
rect 990 2099 991 2103
rect 995 2099 996 2103
rect 990 2098 996 2099
rect 1078 2103 1084 2104
rect 1078 2099 1079 2103
rect 1083 2099 1084 2103
rect 1078 2098 1084 2099
rect 1146 2103 1152 2104
rect 1146 2099 1147 2103
rect 1151 2099 1152 2103
rect 1146 2098 1152 2099
rect 1166 2103 1172 2104
rect 1166 2099 1167 2103
rect 1171 2099 1172 2103
rect 1166 2098 1172 2099
rect 1218 2103 1224 2104
rect 1218 2099 1219 2103
rect 1223 2099 1224 2103
rect 1218 2098 1224 2099
rect 1238 2103 1244 2104
rect 1238 2099 1239 2103
rect 1243 2099 1244 2103
rect 1238 2098 1244 2099
rect 1258 2103 1264 2104
rect 1258 2099 1259 2103
rect 1263 2099 1264 2103
rect 1286 2100 1287 2104
rect 1291 2100 1292 2104
rect 1328 2102 1330 2105
rect 1382 2104 1388 2105
rect 1286 2099 1292 2100
rect 1326 2101 1332 2102
rect 1258 2098 1264 2099
rect 982 2083 988 2084
rect 982 2079 983 2083
rect 987 2079 988 2083
rect 982 2078 988 2079
rect 992 2075 994 2098
rect 1080 2075 1082 2098
rect 1148 2084 1150 2098
rect 1110 2083 1116 2084
rect 1110 2079 1111 2083
rect 1115 2079 1116 2083
rect 1110 2078 1116 2079
rect 1146 2083 1152 2084
rect 1146 2079 1147 2083
rect 1151 2079 1152 2083
rect 1146 2078 1152 2079
rect 863 2074 867 2075
rect 863 2069 867 2070
rect 903 2074 907 2075
rect 903 2069 907 2070
rect 943 2074 947 2075
rect 943 2069 947 2070
rect 991 2074 995 2075
rect 991 2069 995 2070
rect 1023 2074 1027 2075
rect 1023 2069 1027 2070
rect 1079 2074 1083 2075
rect 1079 2069 1083 2070
rect 1103 2074 1107 2075
rect 1103 2069 1107 2070
rect 838 2067 844 2068
rect 838 2063 839 2067
rect 843 2063 844 2067
rect 838 2062 844 2063
rect 864 2050 866 2069
rect 944 2050 946 2069
rect 998 2067 1004 2068
rect 998 2063 999 2067
rect 1003 2063 1004 2067
rect 998 2062 1004 2063
rect 510 2049 516 2050
rect 454 2044 460 2045
rect 474 2047 480 2048
rect 430 2042 436 2043
rect 474 2043 475 2047
rect 479 2043 480 2047
rect 510 2045 511 2049
rect 515 2045 516 2049
rect 510 2044 516 2045
rect 574 2049 580 2050
rect 574 2045 575 2049
rect 579 2045 580 2049
rect 574 2044 580 2045
rect 638 2049 644 2050
rect 638 2045 639 2049
rect 643 2045 644 2049
rect 638 2044 644 2045
rect 710 2049 716 2050
rect 710 2045 711 2049
rect 715 2045 716 2049
rect 790 2049 796 2050
rect 710 2044 716 2045
rect 726 2047 732 2048
rect 474 2042 480 2043
rect 726 2043 727 2047
rect 731 2043 732 2047
rect 790 2045 791 2049
rect 795 2045 796 2049
rect 790 2044 796 2045
rect 862 2049 868 2050
rect 862 2045 863 2049
rect 867 2045 868 2049
rect 862 2044 868 2045
rect 942 2049 948 2050
rect 942 2045 943 2049
rect 947 2045 948 2049
rect 942 2044 948 2045
rect 726 2042 732 2043
rect 110 2031 116 2032
rect 110 2027 111 2031
rect 115 2027 116 2031
rect 110 2026 116 2027
rect 382 2028 388 2029
rect 112 2019 114 2026
rect 382 2024 383 2028
rect 387 2024 388 2028
rect 382 2023 388 2024
rect 384 2019 386 2023
rect 111 2018 115 2019
rect 111 2013 115 2014
rect 231 2018 235 2019
rect 231 2013 235 2014
rect 287 2018 291 2019
rect 287 2013 291 2014
rect 359 2018 363 2019
rect 359 2013 363 2014
rect 383 2018 387 2019
rect 383 2013 387 2014
rect 112 2010 114 2013
rect 230 2012 236 2013
rect 110 2009 116 2010
rect 110 2005 111 2009
rect 115 2005 116 2009
rect 230 2008 231 2012
rect 235 2008 236 2012
rect 230 2007 236 2008
rect 286 2012 292 2013
rect 286 2008 287 2012
rect 291 2008 292 2012
rect 286 2007 292 2008
rect 358 2012 364 2013
rect 358 2008 359 2012
rect 363 2008 364 2012
rect 358 2007 364 2008
rect 110 2004 116 2005
rect 110 1992 116 1993
rect 110 1988 111 1992
rect 115 1988 116 1992
rect 110 1987 116 1988
rect 246 1991 252 1992
rect 246 1987 247 1991
rect 251 1987 252 1991
rect 112 1963 114 1987
rect 246 1986 252 1987
rect 282 1991 288 1992
rect 282 1987 283 1991
rect 287 1987 288 1991
rect 282 1986 288 1987
rect 302 1991 308 1992
rect 302 1987 303 1991
rect 307 1987 308 1991
rect 302 1986 308 1987
rect 354 1991 360 1992
rect 354 1987 355 1991
rect 359 1987 360 1991
rect 354 1986 360 1987
rect 374 1991 380 1992
rect 374 1987 375 1991
rect 379 1987 380 1991
rect 374 1986 380 1987
rect 418 1991 424 1992
rect 418 1987 419 1991
rect 423 1987 424 1991
rect 418 1986 424 1987
rect 231 1980 235 1981
rect 231 1975 235 1976
rect 232 1972 234 1975
rect 230 1971 236 1972
rect 230 1967 231 1971
rect 235 1967 236 1971
rect 230 1966 236 1967
rect 248 1963 250 1986
rect 284 1972 286 1986
rect 282 1971 288 1972
rect 282 1967 283 1971
rect 287 1967 288 1971
rect 282 1966 288 1967
rect 304 1963 306 1986
rect 356 1972 358 1986
rect 354 1971 360 1972
rect 354 1967 355 1971
rect 359 1967 360 1971
rect 354 1966 360 1967
rect 376 1963 378 1986
rect 111 1962 115 1963
rect 111 1957 115 1958
rect 151 1962 155 1963
rect 151 1957 155 1958
rect 215 1962 219 1963
rect 215 1957 219 1958
rect 247 1962 251 1963
rect 247 1957 251 1958
rect 303 1962 307 1963
rect 303 1957 307 1958
rect 319 1962 323 1963
rect 319 1957 323 1958
rect 375 1962 379 1963
rect 375 1957 379 1958
rect 112 1937 114 1957
rect 152 1938 154 1957
rect 166 1955 172 1956
rect 166 1951 167 1955
rect 171 1951 172 1955
rect 166 1950 172 1951
rect 174 1955 180 1956
rect 174 1951 175 1955
rect 179 1951 180 1955
rect 174 1950 180 1951
rect 168 1941 170 1950
rect 167 1940 171 1941
rect 150 1937 156 1938
rect 110 1936 116 1937
rect 110 1932 111 1936
rect 115 1932 116 1936
rect 150 1933 151 1937
rect 155 1933 156 1937
rect 176 1936 178 1950
rect 216 1938 218 1957
rect 238 1955 244 1956
rect 238 1951 239 1955
rect 243 1951 244 1955
rect 238 1950 244 1951
rect 214 1937 220 1938
rect 167 1935 171 1936
rect 174 1935 180 1936
rect 150 1932 156 1933
rect 110 1931 116 1932
rect 174 1931 175 1935
rect 179 1931 180 1935
rect 214 1933 215 1937
rect 219 1933 220 1937
rect 240 1936 242 1950
rect 320 1938 322 1957
rect 420 1956 422 1986
rect 432 1972 434 2042
rect 438 2028 444 2029
rect 438 2024 439 2028
rect 443 2024 444 2028
rect 438 2023 444 2024
rect 494 2028 500 2029
rect 494 2024 495 2028
rect 499 2024 500 2028
rect 494 2023 500 2024
rect 558 2028 564 2029
rect 558 2024 559 2028
rect 563 2024 564 2028
rect 558 2023 564 2024
rect 622 2028 628 2029
rect 622 2024 623 2028
rect 627 2024 628 2028
rect 622 2023 628 2024
rect 694 2028 700 2029
rect 694 2024 695 2028
rect 699 2024 700 2028
rect 694 2023 700 2024
rect 440 2019 442 2023
rect 496 2019 498 2023
rect 560 2019 562 2023
rect 624 2019 626 2023
rect 696 2019 698 2023
rect 439 2018 443 2019
rect 439 2013 443 2014
rect 495 2018 499 2019
rect 495 2013 499 2014
rect 535 2018 539 2019
rect 535 2013 539 2014
rect 559 2018 563 2019
rect 559 2013 563 2014
rect 623 2018 627 2019
rect 623 2013 627 2014
rect 631 2018 635 2019
rect 631 2013 635 2014
rect 695 2018 699 2019
rect 695 2013 699 2014
rect 438 2012 444 2013
rect 438 2008 439 2012
rect 443 2008 444 2012
rect 438 2007 444 2008
rect 534 2012 540 2013
rect 534 2008 535 2012
rect 539 2008 540 2012
rect 534 2007 540 2008
rect 630 2012 636 2013
rect 630 2008 631 2012
rect 635 2008 636 2012
rect 630 2007 636 2008
rect 454 1991 460 1992
rect 454 1987 455 1991
rect 459 1987 460 1991
rect 454 1986 460 1987
rect 530 1991 536 1992
rect 530 1987 531 1991
rect 535 1987 536 1991
rect 530 1986 536 1987
rect 550 1991 556 1992
rect 550 1987 551 1991
rect 555 1987 556 1991
rect 550 1986 556 1987
rect 626 1991 632 1992
rect 626 1987 627 1991
rect 631 1987 632 1991
rect 626 1986 632 1987
rect 646 1991 652 1992
rect 646 1987 647 1991
rect 651 1987 652 1991
rect 646 1986 652 1987
rect 654 1991 660 1992
rect 654 1987 655 1991
rect 659 1987 660 1991
rect 654 1986 660 1987
rect 430 1971 436 1972
rect 430 1967 431 1971
rect 435 1967 436 1971
rect 430 1966 436 1967
rect 456 1963 458 1986
rect 532 1972 534 1986
rect 530 1971 536 1972
rect 530 1967 531 1971
rect 535 1967 536 1971
rect 530 1966 536 1967
rect 552 1963 554 1986
rect 628 1972 630 1986
rect 626 1971 632 1972
rect 626 1967 627 1971
rect 631 1967 632 1971
rect 626 1966 632 1967
rect 648 1963 650 1986
rect 656 1981 658 1986
rect 655 1980 659 1981
rect 655 1975 659 1976
rect 728 1972 730 2042
rect 774 2028 780 2029
rect 774 2024 775 2028
rect 779 2024 780 2028
rect 774 2023 780 2024
rect 846 2028 852 2029
rect 846 2024 847 2028
rect 851 2024 852 2028
rect 846 2023 852 2024
rect 926 2028 932 2029
rect 926 2024 927 2028
rect 931 2024 932 2028
rect 926 2023 932 2024
rect 776 2019 778 2023
rect 848 2019 850 2023
rect 928 2019 930 2023
rect 735 2018 739 2019
rect 735 2013 739 2014
rect 775 2018 779 2019
rect 775 2013 779 2014
rect 847 2018 851 2019
rect 847 2013 851 2014
rect 927 2018 931 2019
rect 927 2013 931 2014
rect 959 2018 963 2019
rect 959 2013 963 2014
rect 734 2012 740 2013
rect 734 2008 735 2012
rect 739 2008 740 2012
rect 734 2007 740 2008
rect 846 2012 852 2013
rect 846 2008 847 2012
rect 851 2008 852 2012
rect 846 2007 852 2008
rect 958 2012 964 2013
rect 958 2008 959 2012
rect 963 2008 964 2012
rect 958 2007 964 2008
rect 1000 1992 1002 2062
rect 1024 2050 1026 2069
rect 1104 2050 1106 2069
rect 1112 2056 1114 2078
rect 1168 2075 1170 2098
rect 1220 2084 1222 2098
rect 1218 2083 1224 2084
rect 1218 2079 1219 2083
rect 1223 2079 1224 2083
rect 1218 2078 1224 2079
rect 1240 2075 1242 2098
rect 1288 2075 1290 2099
rect 1326 2097 1327 2101
rect 1331 2097 1332 2101
rect 1382 2100 1383 2104
rect 1387 2100 1388 2104
rect 1382 2099 1388 2100
rect 1550 2104 1556 2105
rect 1550 2100 1551 2104
rect 1555 2100 1556 2104
rect 1550 2099 1556 2100
rect 1710 2104 1716 2105
rect 1710 2100 1711 2104
rect 1715 2100 1716 2104
rect 1710 2099 1716 2100
rect 1326 2096 1332 2097
rect 1326 2084 1332 2085
rect 1748 2084 1750 2150
rect 1816 2138 1818 2157
rect 1838 2155 1844 2156
rect 1838 2151 1839 2155
rect 1843 2151 1844 2155
rect 1838 2150 1844 2151
rect 1814 2137 1820 2138
rect 1814 2133 1815 2137
rect 1819 2133 1820 2137
rect 1840 2136 1842 2150
rect 1992 2138 1994 2157
rect 2160 2138 2162 2157
rect 2320 2138 2322 2157
rect 2456 2138 2458 2157
rect 2464 2156 2466 2202
rect 2504 2163 2506 2203
rect 2503 2162 2507 2163
rect 2503 2157 2507 2158
rect 2462 2155 2468 2156
rect 2462 2151 2463 2155
rect 2467 2151 2468 2155
rect 2462 2150 2468 2151
rect 1990 2137 1996 2138
rect 1814 2132 1820 2133
rect 1838 2135 1844 2136
rect 1838 2131 1839 2135
rect 1843 2131 1844 2135
rect 1990 2133 1991 2137
rect 1995 2133 1996 2137
rect 2158 2137 2164 2138
rect 1990 2132 1996 2133
rect 2110 2135 2116 2136
rect 1838 2130 1844 2131
rect 2110 2131 2111 2135
rect 2115 2131 2116 2135
rect 2158 2133 2159 2137
rect 2163 2133 2164 2137
rect 2158 2132 2164 2133
rect 2318 2137 2324 2138
rect 2318 2133 2319 2137
rect 2323 2133 2324 2137
rect 2318 2132 2324 2133
rect 2454 2137 2460 2138
rect 2504 2137 2506 2157
rect 2454 2133 2455 2137
rect 2459 2133 2460 2137
rect 2454 2132 2460 2133
rect 2502 2136 2508 2137
rect 2502 2132 2503 2136
rect 2507 2132 2508 2136
rect 2502 2131 2508 2132
rect 2110 2130 2116 2131
rect 1798 2116 1804 2117
rect 1798 2112 1799 2116
rect 1803 2112 1804 2116
rect 1798 2111 1804 2112
rect 1974 2116 1980 2117
rect 1974 2112 1975 2116
rect 1979 2112 1980 2116
rect 1974 2111 1980 2112
rect 1799 2110 1803 2111
rect 1799 2105 1803 2106
rect 1855 2110 1859 2111
rect 1855 2105 1859 2106
rect 1975 2110 1979 2111
rect 1975 2105 1979 2106
rect 1991 2110 1995 2111
rect 1991 2105 1995 2106
rect 1854 2104 1860 2105
rect 1854 2100 1855 2104
rect 1859 2100 1860 2104
rect 1854 2099 1860 2100
rect 1990 2104 1996 2105
rect 1990 2100 1991 2104
rect 1995 2100 1996 2104
rect 1990 2099 1996 2100
rect 1326 2080 1327 2084
rect 1331 2080 1332 2084
rect 1326 2079 1332 2080
rect 1398 2083 1404 2084
rect 1398 2079 1399 2083
rect 1403 2079 1404 2083
rect 1167 2074 1171 2075
rect 1167 2069 1171 2070
rect 1183 2074 1187 2075
rect 1183 2069 1187 2070
rect 1239 2074 1243 2075
rect 1239 2069 1243 2070
rect 1287 2074 1291 2075
rect 1287 2069 1291 2070
rect 1126 2067 1132 2068
rect 1126 2063 1127 2067
rect 1131 2063 1132 2067
rect 1126 2062 1132 2063
rect 1110 2055 1116 2056
rect 1110 2051 1111 2055
rect 1115 2051 1116 2055
rect 1110 2050 1116 2051
rect 1022 2049 1028 2050
rect 1022 2045 1023 2049
rect 1027 2045 1028 2049
rect 1022 2044 1028 2045
rect 1102 2049 1108 2050
rect 1102 2045 1103 2049
rect 1107 2045 1108 2049
rect 1128 2048 1130 2062
rect 1184 2050 1186 2069
rect 1206 2067 1212 2068
rect 1206 2063 1207 2067
rect 1211 2063 1212 2067
rect 1206 2062 1212 2063
rect 1182 2049 1188 2050
rect 1102 2044 1108 2045
rect 1126 2047 1132 2048
rect 1126 2043 1127 2047
rect 1131 2043 1132 2047
rect 1182 2045 1183 2049
rect 1187 2045 1188 2049
rect 1208 2048 1210 2062
rect 1240 2050 1242 2069
rect 1238 2049 1244 2050
rect 1288 2049 1290 2069
rect 1328 2055 1330 2079
rect 1398 2078 1404 2079
rect 1546 2083 1552 2084
rect 1546 2079 1547 2083
rect 1551 2079 1552 2083
rect 1546 2078 1552 2079
rect 1566 2083 1572 2084
rect 1566 2079 1567 2083
rect 1571 2079 1572 2083
rect 1566 2078 1572 2079
rect 1706 2083 1712 2084
rect 1706 2079 1707 2083
rect 1711 2079 1712 2083
rect 1706 2078 1712 2079
rect 1726 2083 1732 2084
rect 1726 2079 1727 2083
rect 1731 2079 1732 2083
rect 1726 2078 1732 2079
rect 1746 2083 1752 2084
rect 1746 2079 1747 2083
rect 1751 2079 1752 2083
rect 1746 2078 1752 2079
rect 1870 2083 1876 2084
rect 1870 2079 1871 2083
rect 1875 2079 1876 2083
rect 1870 2078 1876 2079
rect 1906 2083 1912 2084
rect 1906 2079 1907 2083
rect 1911 2079 1912 2083
rect 1906 2078 1912 2079
rect 2006 2083 2012 2084
rect 2006 2079 2007 2083
rect 2011 2079 2012 2083
rect 2006 2078 2012 2079
rect 1400 2055 1402 2078
rect 1548 2064 1550 2078
rect 1466 2063 1472 2064
rect 1466 2059 1467 2063
rect 1471 2059 1472 2063
rect 1466 2058 1472 2059
rect 1546 2063 1552 2064
rect 1546 2059 1547 2063
rect 1551 2059 1552 2063
rect 1546 2058 1552 2059
rect 1327 2054 1331 2055
rect 1327 2049 1331 2050
rect 1399 2054 1403 2055
rect 1399 2049 1403 2050
rect 1447 2054 1451 2055
rect 1447 2049 1451 2050
rect 1182 2044 1188 2045
rect 1206 2047 1212 2048
rect 1126 2042 1132 2043
rect 1206 2043 1207 2047
rect 1211 2043 1212 2047
rect 1238 2045 1239 2049
rect 1243 2045 1244 2049
rect 1238 2044 1244 2045
rect 1286 2048 1292 2049
rect 1286 2044 1287 2048
rect 1291 2044 1292 2048
rect 1286 2043 1292 2044
rect 1206 2042 1212 2043
rect 1286 2031 1292 2032
rect 1006 2028 1012 2029
rect 1006 2024 1007 2028
rect 1011 2024 1012 2028
rect 1006 2023 1012 2024
rect 1086 2028 1092 2029
rect 1086 2024 1087 2028
rect 1091 2024 1092 2028
rect 1086 2023 1092 2024
rect 1166 2028 1172 2029
rect 1166 2024 1167 2028
rect 1171 2024 1172 2028
rect 1166 2023 1172 2024
rect 1222 2028 1228 2029
rect 1222 2024 1223 2028
rect 1227 2024 1228 2028
rect 1286 2027 1287 2031
rect 1291 2027 1292 2031
rect 1328 2029 1330 2049
rect 1448 2030 1450 2049
rect 1446 2029 1452 2030
rect 1286 2026 1292 2027
rect 1326 2028 1332 2029
rect 1222 2023 1228 2024
rect 1008 2019 1010 2023
rect 1088 2019 1090 2023
rect 1168 2019 1170 2023
rect 1224 2019 1226 2023
rect 1288 2019 1290 2026
rect 1326 2024 1327 2028
rect 1331 2024 1332 2028
rect 1446 2025 1447 2029
rect 1451 2025 1452 2029
rect 1468 2028 1470 2058
rect 1568 2055 1570 2078
rect 1708 2064 1710 2078
rect 1706 2063 1712 2064
rect 1706 2059 1707 2063
rect 1711 2059 1712 2063
rect 1706 2058 1712 2059
rect 1728 2055 1730 2078
rect 1872 2055 1874 2078
rect 1551 2054 1555 2055
rect 1551 2049 1555 2050
rect 1567 2054 1571 2055
rect 1567 2049 1571 2050
rect 1655 2054 1659 2055
rect 1655 2049 1659 2050
rect 1727 2054 1731 2055
rect 1727 2049 1731 2050
rect 1751 2054 1755 2055
rect 1751 2049 1755 2050
rect 1839 2054 1843 2055
rect 1839 2049 1843 2050
rect 1871 2054 1875 2055
rect 1871 2049 1875 2050
rect 1542 2047 1548 2048
rect 1542 2043 1543 2047
rect 1547 2043 1548 2047
rect 1542 2042 1548 2043
rect 1446 2024 1452 2025
rect 1466 2027 1472 2028
rect 1326 2023 1332 2024
rect 1466 2023 1467 2027
rect 1471 2023 1472 2027
rect 1466 2022 1472 2023
rect 1007 2018 1011 2019
rect 1007 2013 1011 2014
rect 1079 2018 1083 2019
rect 1079 2013 1083 2014
rect 1087 2018 1091 2019
rect 1087 2013 1091 2014
rect 1167 2018 1171 2019
rect 1167 2013 1171 2014
rect 1199 2018 1203 2019
rect 1199 2013 1203 2014
rect 1223 2018 1227 2019
rect 1223 2013 1227 2014
rect 1287 2018 1291 2019
rect 1287 2013 1291 2014
rect 1078 2012 1084 2013
rect 1078 2008 1079 2012
rect 1083 2008 1084 2012
rect 1078 2007 1084 2008
rect 1198 2012 1204 2013
rect 1198 2008 1199 2012
rect 1203 2008 1204 2012
rect 1288 2010 1290 2013
rect 1326 2011 1332 2012
rect 1198 2007 1204 2008
rect 1286 2009 1292 2010
rect 1286 2005 1287 2009
rect 1291 2005 1292 2009
rect 1326 2007 1327 2011
rect 1331 2007 1332 2011
rect 1326 2006 1332 2007
rect 1430 2008 1436 2009
rect 1286 2004 1292 2005
rect 1328 1999 1330 2006
rect 1430 2004 1431 2008
rect 1435 2004 1436 2008
rect 1430 2003 1436 2004
rect 1534 2008 1540 2009
rect 1534 2004 1535 2008
rect 1539 2004 1540 2008
rect 1534 2003 1540 2004
rect 1432 1999 1434 2003
rect 1536 1999 1538 2003
rect 1327 1998 1331 1999
rect 1327 1993 1331 1994
rect 1431 1998 1435 1999
rect 1431 1993 1435 1994
rect 1455 1998 1459 1999
rect 1455 1993 1459 1994
rect 1511 1998 1515 1999
rect 1511 1993 1515 1994
rect 1535 1998 1539 1999
rect 1535 1993 1539 1994
rect 1286 1992 1292 1993
rect 750 1991 756 1992
rect 750 1987 751 1991
rect 755 1987 756 1991
rect 750 1986 756 1987
rect 842 1991 848 1992
rect 842 1987 843 1991
rect 847 1987 848 1991
rect 842 1986 848 1987
rect 862 1991 868 1992
rect 862 1987 863 1991
rect 867 1987 868 1991
rect 862 1986 868 1987
rect 898 1991 904 1992
rect 898 1987 899 1991
rect 903 1987 904 1991
rect 898 1986 904 1987
rect 974 1991 980 1992
rect 974 1987 975 1991
rect 979 1987 980 1991
rect 974 1986 980 1987
rect 998 1991 1004 1992
rect 998 1987 999 1991
rect 1003 1987 1004 1991
rect 998 1986 1004 1987
rect 1094 1991 1100 1992
rect 1094 1987 1095 1991
rect 1099 1987 1100 1991
rect 1094 1986 1100 1987
rect 1194 1991 1200 1992
rect 1194 1987 1195 1991
rect 1199 1987 1200 1991
rect 1194 1986 1200 1987
rect 1214 1991 1220 1992
rect 1214 1987 1215 1991
rect 1219 1987 1220 1991
rect 1286 1988 1287 1992
rect 1291 1988 1292 1992
rect 1328 1990 1330 1993
rect 1454 1992 1460 1993
rect 1286 1987 1292 1988
rect 1326 1989 1332 1990
rect 1214 1986 1220 1987
rect 726 1971 732 1972
rect 726 1967 727 1971
rect 731 1967 732 1971
rect 726 1966 732 1967
rect 752 1963 754 1986
rect 844 1972 846 1986
rect 842 1971 848 1972
rect 842 1967 843 1971
rect 847 1967 848 1971
rect 842 1966 848 1967
rect 864 1963 866 1986
rect 439 1962 443 1963
rect 439 1957 443 1958
rect 455 1962 459 1963
rect 455 1957 459 1958
rect 551 1962 555 1963
rect 551 1957 555 1958
rect 583 1962 587 1963
rect 583 1957 587 1958
rect 647 1962 651 1963
rect 647 1957 651 1958
rect 743 1962 747 1963
rect 743 1957 747 1958
rect 751 1962 755 1963
rect 751 1957 755 1958
rect 863 1962 867 1963
rect 863 1957 867 1958
rect 418 1955 424 1956
rect 418 1951 419 1955
rect 423 1951 424 1955
rect 418 1950 424 1951
rect 440 1938 442 1957
rect 462 1955 468 1956
rect 462 1951 463 1955
rect 467 1951 468 1955
rect 462 1950 468 1951
rect 318 1937 324 1938
rect 214 1932 220 1933
rect 238 1935 244 1936
rect 174 1930 180 1931
rect 238 1931 239 1935
rect 243 1931 244 1935
rect 318 1933 319 1937
rect 323 1933 324 1937
rect 438 1937 444 1938
rect 318 1932 324 1933
rect 350 1935 356 1936
rect 238 1930 244 1931
rect 350 1931 351 1935
rect 355 1931 356 1935
rect 438 1933 439 1937
rect 443 1933 444 1937
rect 464 1936 466 1950
rect 584 1938 586 1957
rect 603 1940 607 1941
rect 582 1937 588 1938
rect 438 1932 444 1933
rect 462 1935 468 1936
rect 350 1930 356 1931
rect 462 1931 463 1935
rect 467 1931 468 1935
rect 582 1933 583 1937
rect 587 1933 588 1937
rect 744 1938 746 1957
rect 900 1956 902 1986
rect 976 1963 978 1986
rect 1096 1963 1098 1986
rect 1196 1972 1198 1986
rect 1114 1971 1120 1972
rect 1114 1967 1115 1971
rect 1119 1967 1120 1971
rect 1114 1966 1120 1967
rect 1194 1971 1200 1972
rect 1194 1967 1195 1971
rect 1199 1967 1200 1971
rect 1194 1966 1200 1967
rect 919 1962 923 1963
rect 919 1957 923 1958
rect 975 1962 979 1963
rect 975 1957 979 1958
rect 1095 1962 1099 1963
rect 1095 1957 1099 1958
rect 898 1955 904 1956
rect 898 1951 899 1955
rect 903 1951 904 1955
rect 898 1950 904 1951
rect 920 1938 922 1957
rect 1054 1955 1060 1956
rect 1054 1951 1055 1955
rect 1059 1951 1060 1955
rect 1054 1950 1060 1951
rect 742 1937 748 1938
rect 582 1932 588 1933
rect 602 1935 608 1936
rect 462 1930 468 1931
rect 602 1931 603 1935
rect 607 1931 608 1935
rect 742 1933 743 1937
rect 747 1933 748 1937
rect 918 1937 924 1938
rect 742 1932 748 1933
rect 750 1935 756 1936
rect 602 1930 608 1931
rect 750 1931 751 1935
rect 755 1931 756 1935
rect 918 1933 919 1937
rect 923 1933 924 1937
rect 918 1932 924 1933
rect 750 1930 756 1931
rect 110 1919 116 1920
rect 110 1915 111 1919
rect 115 1915 116 1919
rect 110 1914 116 1915
rect 134 1916 140 1917
rect 112 1903 114 1914
rect 134 1912 135 1916
rect 139 1912 140 1916
rect 134 1911 140 1912
rect 198 1916 204 1917
rect 198 1912 199 1916
rect 203 1912 204 1916
rect 198 1911 204 1912
rect 302 1916 308 1917
rect 302 1912 303 1916
rect 307 1912 308 1916
rect 302 1911 308 1912
rect 136 1903 138 1911
rect 200 1903 202 1911
rect 304 1903 306 1911
rect 111 1902 115 1903
rect 111 1897 115 1898
rect 135 1902 139 1903
rect 135 1897 139 1898
rect 191 1902 195 1903
rect 191 1897 195 1898
rect 199 1902 203 1903
rect 199 1897 203 1898
rect 271 1902 275 1903
rect 271 1897 275 1898
rect 303 1902 307 1903
rect 303 1897 307 1898
rect 112 1894 114 1897
rect 134 1896 140 1897
rect 110 1893 116 1894
rect 110 1889 111 1893
rect 115 1889 116 1893
rect 134 1892 135 1896
rect 139 1892 140 1896
rect 134 1891 140 1892
rect 190 1896 196 1897
rect 190 1892 191 1896
rect 195 1892 196 1896
rect 190 1891 196 1892
rect 270 1896 276 1897
rect 270 1892 271 1896
rect 275 1892 276 1896
rect 270 1891 276 1892
rect 110 1888 116 1889
rect 110 1876 116 1877
rect 110 1872 111 1876
rect 115 1872 116 1876
rect 110 1871 116 1872
rect 150 1875 156 1876
rect 150 1871 151 1875
rect 155 1871 156 1875
rect 112 1851 114 1871
rect 150 1870 156 1871
rect 158 1875 164 1876
rect 158 1871 159 1875
rect 163 1871 164 1875
rect 158 1870 164 1871
rect 206 1875 212 1876
rect 206 1871 207 1875
rect 211 1871 212 1875
rect 206 1870 212 1871
rect 286 1875 292 1876
rect 286 1871 287 1875
rect 291 1871 292 1875
rect 286 1870 292 1871
rect 152 1851 154 1870
rect 111 1850 115 1851
rect 111 1845 115 1846
rect 151 1850 155 1851
rect 151 1845 155 1846
rect 112 1825 114 1845
rect 152 1826 154 1845
rect 160 1844 162 1870
rect 208 1851 210 1870
rect 288 1851 290 1870
rect 352 1856 354 1930
rect 422 1916 428 1917
rect 422 1912 423 1916
rect 427 1912 428 1916
rect 422 1911 428 1912
rect 566 1916 572 1917
rect 566 1912 567 1916
rect 571 1912 572 1916
rect 566 1911 572 1912
rect 726 1916 732 1917
rect 726 1912 727 1916
rect 731 1912 732 1916
rect 726 1911 732 1912
rect 424 1903 426 1911
rect 568 1903 570 1911
rect 728 1903 730 1911
rect 359 1902 363 1903
rect 359 1897 363 1898
rect 423 1902 427 1903
rect 423 1897 427 1898
rect 455 1902 459 1903
rect 455 1897 459 1898
rect 543 1902 547 1903
rect 543 1897 547 1898
rect 567 1902 571 1903
rect 567 1897 571 1898
rect 631 1902 635 1903
rect 631 1897 635 1898
rect 719 1902 723 1903
rect 719 1897 723 1898
rect 727 1902 731 1903
rect 727 1897 731 1898
rect 358 1896 364 1897
rect 358 1892 359 1896
rect 363 1892 364 1896
rect 358 1891 364 1892
rect 454 1896 460 1897
rect 454 1892 455 1896
rect 459 1892 460 1896
rect 454 1891 460 1892
rect 542 1896 548 1897
rect 542 1892 543 1896
rect 547 1892 548 1896
rect 542 1891 548 1892
rect 630 1896 636 1897
rect 630 1892 631 1896
rect 635 1892 636 1896
rect 630 1891 636 1892
rect 718 1896 724 1897
rect 718 1892 719 1896
rect 723 1892 724 1896
rect 718 1891 724 1892
rect 374 1875 380 1876
rect 374 1871 375 1875
rect 379 1871 380 1875
rect 374 1870 380 1871
rect 450 1875 456 1876
rect 450 1871 451 1875
rect 455 1871 456 1875
rect 450 1870 456 1871
rect 470 1875 476 1876
rect 470 1871 471 1875
rect 475 1871 476 1875
rect 470 1870 476 1871
rect 558 1875 564 1876
rect 558 1871 559 1875
rect 563 1871 564 1875
rect 558 1870 564 1871
rect 574 1875 580 1876
rect 574 1871 575 1875
rect 579 1871 580 1875
rect 574 1870 580 1871
rect 646 1875 652 1876
rect 646 1871 647 1875
rect 651 1871 652 1875
rect 646 1870 652 1871
rect 734 1875 740 1876
rect 734 1871 735 1875
rect 739 1871 740 1875
rect 734 1870 740 1871
rect 350 1855 356 1856
rect 350 1851 351 1855
rect 355 1851 356 1855
rect 376 1851 378 1870
rect 452 1856 454 1870
rect 450 1855 456 1856
rect 450 1851 451 1855
rect 455 1851 456 1855
rect 472 1851 474 1870
rect 560 1851 562 1870
rect 207 1850 211 1851
rect 207 1845 211 1846
rect 287 1850 291 1851
rect 287 1845 291 1846
rect 295 1850 299 1851
rect 350 1850 356 1851
rect 375 1850 379 1851
rect 295 1845 299 1846
rect 375 1845 379 1846
rect 391 1850 395 1851
rect 450 1850 456 1851
rect 471 1850 475 1851
rect 391 1845 395 1846
rect 471 1845 475 1846
rect 495 1850 499 1851
rect 495 1845 499 1846
rect 559 1850 563 1851
rect 559 1845 563 1846
rect 158 1843 164 1844
rect 158 1839 159 1843
rect 163 1839 164 1843
rect 158 1838 164 1839
rect 174 1843 180 1844
rect 174 1839 175 1843
rect 179 1839 180 1843
rect 174 1838 180 1839
rect 150 1825 156 1826
rect 110 1824 116 1825
rect 110 1820 111 1824
rect 115 1820 116 1824
rect 150 1821 151 1825
rect 155 1821 156 1825
rect 176 1824 178 1838
rect 208 1826 210 1845
rect 230 1843 236 1844
rect 230 1839 231 1843
rect 235 1839 236 1843
rect 230 1838 236 1839
rect 206 1825 212 1826
rect 150 1820 156 1821
rect 174 1823 180 1824
rect 110 1819 116 1820
rect 174 1819 175 1823
rect 179 1819 180 1823
rect 206 1821 207 1825
rect 211 1821 212 1825
rect 232 1824 234 1838
rect 296 1826 298 1845
rect 392 1826 394 1845
rect 410 1843 416 1844
rect 410 1839 411 1843
rect 415 1839 416 1843
rect 410 1838 416 1839
rect 294 1825 300 1826
rect 206 1820 212 1821
rect 230 1823 236 1824
rect 174 1818 180 1819
rect 230 1819 231 1823
rect 235 1819 236 1823
rect 294 1821 295 1825
rect 299 1821 300 1825
rect 294 1820 300 1821
rect 390 1825 396 1826
rect 390 1821 391 1825
rect 395 1821 396 1825
rect 412 1824 414 1838
rect 496 1826 498 1845
rect 576 1844 578 1870
rect 648 1851 650 1870
rect 710 1855 716 1856
rect 710 1851 711 1855
rect 715 1851 716 1855
rect 736 1851 738 1870
rect 752 1864 754 1930
rect 902 1916 908 1917
rect 902 1912 903 1916
rect 907 1912 908 1916
rect 902 1911 908 1912
rect 904 1903 906 1911
rect 799 1902 803 1903
rect 799 1897 803 1898
rect 871 1902 875 1903
rect 871 1897 875 1898
rect 903 1902 907 1903
rect 903 1897 907 1898
rect 943 1902 947 1903
rect 943 1897 947 1898
rect 1015 1902 1019 1903
rect 1015 1897 1019 1898
rect 798 1896 804 1897
rect 798 1892 799 1896
rect 803 1892 804 1896
rect 798 1891 804 1892
rect 870 1896 876 1897
rect 870 1892 871 1896
rect 875 1892 876 1896
rect 870 1891 876 1892
rect 942 1896 948 1897
rect 942 1892 943 1896
rect 947 1892 948 1896
rect 942 1891 948 1892
rect 1014 1896 1020 1897
rect 1014 1892 1015 1896
rect 1019 1892 1020 1896
rect 1014 1891 1020 1892
rect 1056 1876 1058 1950
rect 1096 1938 1098 1957
rect 1094 1937 1100 1938
rect 1094 1933 1095 1937
rect 1099 1933 1100 1937
rect 1116 1936 1118 1966
rect 1216 1963 1218 1986
rect 1288 1963 1290 1987
rect 1326 1985 1327 1989
rect 1331 1985 1332 1989
rect 1454 1988 1455 1992
rect 1459 1988 1460 1992
rect 1454 1987 1460 1988
rect 1510 1992 1516 1993
rect 1510 1988 1511 1992
rect 1515 1988 1516 1992
rect 1510 1987 1516 1988
rect 1326 1984 1332 1985
rect 1326 1972 1332 1973
rect 1544 1972 1546 2042
rect 1552 2030 1554 2049
rect 1574 2047 1580 2048
rect 1574 2043 1575 2047
rect 1579 2043 1580 2047
rect 1574 2042 1580 2043
rect 1550 2029 1556 2030
rect 1550 2025 1551 2029
rect 1555 2025 1556 2029
rect 1576 2028 1578 2042
rect 1656 2030 1658 2049
rect 1752 2030 1754 2049
rect 1840 2030 1842 2049
rect 1908 2048 1910 2078
rect 2008 2055 2010 2078
rect 2112 2064 2114 2130
rect 2502 2119 2508 2120
rect 2142 2116 2148 2117
rect 2142 2112 2143 2116
rect 2147 2112 2148 2116
rect 2142 2111 2148 2112
rect 2302 2116 2308 2117
rect 2302 2112 2303 2116
rect 2307 2112 2308 2116
rect 2302 2111 2308 2112
rect 2438 2116 2444 2117
rect 2438 2112 2439 2116
rect 2443 2112 2444 2116
rect 2502 2115 2503 2119
rect 2507 2115 2508 2119
rect 2502 2114 2508 2115
rect 2438 2111 2444 2112
rect 2504 2111 2506 2114
rect 2119 2110 2123 2111
rect 2119 2105 2123 2106
rect 2143 2110 2147 2111
rect 2143 2105 2147 2106
rect 2239 2110 2243 2111
rect 2239 2105 2243 2106
rect 2303 2110 2307 2111
rect 2303 2105 2307 2106
rect 2367 2110 2371 2111
rect 2367 2105 2371 2106
rect 2439 2110 2443 2111
rect 2439 2105 2443 2106
rect 2503 2110 2507 2111
rect 2503 2105 2507 2106
rect 2118 2104 2124 2105
rect 2118 2100 2119 2104
rect 2123 2100 2124 2104
rect 2118 2099 2124 2100
rect 2238 2104 2244 2105
rect 2238 2100 2239 2104
rect 2243 2100 2244 2104
rect 2238 2099 2244 2100
rect 2366 2104 2372 2105
rect 2366 2100 2367 2104
rect 2371 2100 2372 2104
rect 2504 2102 2506 2105
rect 2366 2099 2372 2100
rect 2502 2101 2508 2102
rect 2502 2097 2503 2101
rect 2507 2097 2508 2101
rect 2502 2096 2508 2097
rect 2502 2084 2508 2085
rect 2134 2083 2140 2084
rect 2134 2079 2135 2083
rect 2139 2079 2140 2083
rect 2134 2078 2140 2079
rect 2234 2083 2240 2084
rect 2234 2079 2235 2083
rect 2239 2079 2240 2083
rect 2234 2078 2240 2079
rect 2254 2083 2260 2084
rect 2254 2079 2255 2083
rect 2259 2079 2260 2083
rect 2254 2078 2260 2079
rect 2362 2083 2368 2084
rect 2362 2079 2363 2083
rect 2367 2079 2368 2083
rect 2362 2078 2368 2079
rect 2382 2083 2388 2084
rect 2382 2079 2383 2083
rect 2387 2079 2388 2083
rect 2502 2080 2503 2084
rect 2507 2080 2508 2084
rect 2502 2079 2508 2080
rect 2382 2078 2388 2079
rect 2110 2063 2116 2064
rect 2110 2059 2111 2063
rect 2115 2059 2116 2063
rect 2110 2058 2116 2059
rect 2136 2055 2138 2078
rect 2236 2064 2238 2078
rect 2234 2063 2240 2064
rect 2234 2059 2235 2063
rect 2239 2059 2240 2063
rect 2234 2058 2240 2059
rect 2256 2055 2258 2078
rect 2364 2064 2366 2078
rect 2362 2063 2368 2064
rect 2362 2059 2363 2063
rect 2367 2059 2368 2063
rect 2362 2058 2368 2059
rect 2384 2055 2386 2078
rect 2504 2055 2506 2079
rect 1927 2054 1931 2055
rect 1927 2049 1931 2050
rect 2007 2054 2011 2055
rect 2007 2049 2011 2050
rect 2023 2054 2027 2055
rect 2023 2049 2027 2050
rect 2119 2054 2123 2055
rect 2119 2049 2123 2050
rect 2135 2054 2139 2055
rect 2135 2049 2139 2050
rect 2255 2054 2259 2055
rect 2255 2049 2259 2050
rect 2383 2054 2387 2055
rect 2383 2049 2387 2050
rect 2503 2054 2507 2055
rect 2503 2049 2507 2050
rect 1906 2047 1912 2048
rect 1906 2043 1907 2047
rect 1911 2043 1912 2047
rect 1906 2042 1912 2043
rect 1928 2030 1930 2049
rect 1950 2047 1956 2048
rect 1950 2043 1951 2047
rect 1955 2043 1956 2047
rect 1950 2042 1956 2043
rect 1654 2029 1660 2030
rect 1550 2024 1556 2025
rect 1574 2027 1580 2028
rect 1574 2023 1575 2027
rect 1579 2023 1580 2027
rect 1654 2025 1655 2029
rect 1659 2025 1660 2029
rect 1654 2024 1660 2025
rect 1750 2029 1756 2030
rect 1750 2025 1751 2029
rect 1755 2025 1756 2029
rect 1838 2029 1844 2030
rect 1750 2024 1756 2025
rect 1774 2027 1780 2028
rect 1574 2022 1580 2023
rect 1774 2023 1775 2027
rect 1779 2023 1780 2027
rect 1838 2025 1839 2029
rect 1843 2025 1844 2029
rect 1838 2024 1844 2025
rect 1926 2029 1932 2030
rect 1926 2025 1927 2029
rect 1931 2025 1932 2029
rect 1952 2028 1954 2042
rect 2024 2030 2026 2049
rect 2046 2047 2052 2048
rect 2046 2043 2047 2047
rect 2051 2043 2052 2047
rect 2046 2042 2052 2043
rect 2022 2029 2028 2030
rect 1926 2024 1932 2025
rect 1950 2027 1956 2028
rect 1774 2022 1780 2023
rect 1950 2023 1951 2027
rect 1955 2023 1956 2027
rect 2022 2025 2023 2029
rect 2027 2025 2028 2029
rect 2048 2028 2050 2042
rect 2120 2030 2122 2049
rect 2118 2029 2124 2030
rect 2504 2029 2506 2049
rect 2022 2024 2028 2025
rect 2046 2027 2052 2028
rect 1950 2022 1956 2023
rect 2046 2023 2047 2027
rect 2051 2023 2052 2027
rect 2118 2025 2119 2029
rect 2123 2025 2124 2029
rect 2118 2024 2124 2025
rect 2502 2028 2508 2029
rect 2502 2024 2503 2028
rect 2507 2024 2508 2028
rect 2502 2023 2508 2024
rect 2046 2022 2052 2023
rect 1638 2008 1644 2009
rect 1638 2004 1639 2008
rect 1643 2004 1644 2008
rect 1638 2003 1644 2004
rect 1734 2008 1740 2009
rect 1734 2004 1735 2008
rect 1739 2004 1740 2008
rect 1734 2003 1740 2004
rect 1640 1999 1642 2003
rect 1736 1999 1738 2003
rect 1575 1998 1579 1999
rect 1575 1993 1579 1994
rect 1639 1998 1643 1999
rect 1639 1993 1643 1994
rect 1703 1998 1707 1999
rect 1703 1993 1707 1994
rect 1735 1998 1739 1999
rect 1735 1993 1739 1994
rect 1767 1998 1771 1999
rect 1767 1993 1771 1994
rect 1574 1992 1580 1993
rect 1574 1988 1575 1992
rect 1579 1988 1580 1992
rect 1574 1987 1580 1988
rect 1638 1992 1644 1993
rect 1638 1988 1639 1992
rect 1643 1988 1644 1992
rect 1638 1987 1644 1988
rect 1702 1992 1708 1993
rect 1702 1988 1703 1992
rect 1707 1988 1708 1992
rect 1702 1987 1708 1988
rect 1766 1992 1772 1993
rect 1766 1988 1767 1992
rect 1771 1988 1772 1992
rect 1766 1987 1772 1988
rect 1326 1968 1327 1972
rect 1331 1968 1332 1972
rect 1326 1967 1332 1968
rect 1470 1971 1476 1972
rect 1470 1967 1471 1971
rect 1475 1967 1476 1971
rect 1215 1962 1219 1963
rect 1215 1957 1219 1958
rect 1287 1962 1291 1963
rect 1287 1957 1291 1958
rect 1288 1937 1290 1957
rect 1328 1943 1330 1967
rect 1470 1966 1476 1967
rect 1506 1971 1512 1972
rect 1506 1967 1507 1971
rect 1511 1967 1512 1971
rect 1506 1966 1512 1967
rect 1526 1971 1532 1972
rect 1526 1967 1527 1971
rect 1531 1967 1532 1971
rect 1526 1966 1532 1967
rect 1542 1971 1548 1972
rect 1542 1967 1543 1971
rect 1547 1967 1548 1971
rect 1542 1966 1548 1967
rect 1590 1971 1596 1972
rect 1590 1967 1591 1971
rect 1595 1967 1596 1971
rect 1590 1966 1596 1967
rect 1598 1971 1604 1972
rect 1598 1967 1599 1971
rect 1603 1967 1604 1971
rect 1598 1966 1604 1967
rect 1654 1971 1660 1972
rect 1654 1967 1655 1971
rect 1659 1967 1660 1971
rect 1654 1966 1660 1967
rect 1718 1971 1724 1972
rect 1718 1967 1719 1971
rect 1723 1967 1724 1971
rect 1718 1966 1724 1967
rect 1472 1943 1474 1966
rect 1508 1952 1510 1966
rect 1506 1951 1512 1952
rect 1506 1947 1507 1951
rect 1511 1947 1512 1951
rect 1506 1946 1512 1947
rect 1528 1943 1530 1966
rect 1592 1943 1594 1966
rect 1600 1944 1602 1966
rect 1598 1943 1604 1944
rect 1656 1943 1658 1966
rect 1710 1951 1716 1952
rect 1710 1947 1711 1951
rect 1715 1947 1716 1951
rect 1710 1946 1716 1947
rect 1327 1942 1331 1943
rect 1327 1937 1331 1938
rect 1471 1942 1475 1943
rect 1471 1937 1475 1938
rect 1527 1942 1531 1943
rect 1527 1937 1531 1938
rect 1567 1942 1571 1943
rect 1567 1937 1571 1938
rect 1591 1942 1595 1943
rect 1598 1939 1599 1943
rect 1603 1939 1604 1943
rect 1598 1938 1604 1939
rect 1631 1942 1635 1943
rect 1591 1937 1595 1938
rect 1631 1937 1635 1938
rect 1655 1942 1659 1943
rect 1655 1937 1659 1938
rect 1703 1942 1707 1943
rect 1703 1937 1707 1938
rect 1286 1936 1292 1937
rect 1094 1932 1100 1933
rect 1114 1935 1120 1936
rect 1114 1931 1115 1935
rect 1119 1931 1120 1935
rect 1286 1932 1287 1936
rect 1291 1932 1292 1936
rect 1286 1931 1292 1932
rect 1114 1930 1120 1931
rect 1286 1919 1292 1920
rect 1078 1916 1084 1917
rect 1078 1912 1079 1916
rect 1083 1912 1084 1916
rect 1286 1915 1287 1919
rect 1291 1915 1292 1919
rect 1328 1917 1330 1937
rect 1568 1918 1570 1937
rect 1598 1935 1604 1936
rect 1598 1931 1599 1935
rect 1603 1931 1604 1935
rect 1598 1930 1604 1931
rect 1566 1917 1572 1918
rect 1286 1914 1292 1915
rect 1326 1916 1332 1917
rect 1078 1911 1084 1912
rect 1080 1903 1082 1911
rect 1288 1903 1290 1914
rect 1326 1912 1327 1916
rect 1331 1912 1332 1916
rect 1566 1913 1567 1917
rect 1571 1913 1572 1917
rect 1600 1916 1602 1930
rect 1632 1918 1634 1937
rect 1662 1935 1668 1936
rect 1662 1931 1663 1935
rect 1667 1931 1668 1935
rect 1662 1930 1668 1931
rect 1630 1917 1636 1918
rect 1566 1912 1572 1913
rect 1598 1915 1604 1916
rect 1326 1911 1332 1912
rect 1598 1911 1599 1915
rect 1603 1911 1604 1915
rect 1630 1913 1631 1917
rect 1635 1913 1636 1917
rect 1664 1916 1666 1930
rect 1704 1918 1706 1937
rect 1702 1917 1708 1918
rect 1630 1912 1636 1913
rect 1662 1915 1668 1916
rect 1598 1910 1604 1911
rect 1662 1911 1663 1915
rect 1667 1911 1668 1915
rect 1702 1913 1703 1917
rect 1707 1913 1708 1917
rect 1712 1916 1714 1946
rect 1720 1943 1722 1966
rect 1776 1952 1778 2022
rect 2502 2011 2508 2012
rect 1822 2008 1828 2009
rect 1822 2004 1823 2008
rect 1827 2004 1828 2008
rect 1822 2003 1828 2004
rect 1910 2008 1916 2009
rect 1910 2004 1911 2008
rect 1915 2004 1916 2008
rect 1910 2003 1916 2004
rect 2006 2008 2012 2009
rect 2006 2004 2007 2008
rect 2011 2004 2012 2008
rect 2006 2003 2012 2004
rect 2102 2008 2108 2009
rect 2102 2004 2103 2008
rect 2107 2004 2108 2008
rect 2502 2007 2503 2011
rect 2507 2007 2508 2011
rect 2502 2006 2508 2007
rect 2102 2003 2108 2004
rect 1824 1999 1826 2003
rect 1912 1999 1914 2003
rect 2008 1999 2010 2003
rect 2104 1999 2106 2003
rect 2504 1999 2506 2006
rect 1823 1998 1827 1999
rect 1823 1993 1827 1994
rect 1831 1998 1835 1999
rect 1831 1993 1835 1994
rect 1895 1998 1899 1999
rect 1895 1993 1899 1994
rect 1911 1998 1915 1999
rect 1911 1993 1915 1994
rect 1959 1998 1963 1999
rect 1959 1993 1963 1994
rect 2007 1998 2011 1999
rect 2007 1993 2011 1994
rect 2031 1998 2035 1999
rect 2031 1993 2035 1994
rect 2103 1998 2107 1999
rect 2103 1993 2107 1994
rect 2503 1998 2507 1999
rect 2503 1993 2507 1994
rect 1830 1992 1836 1993
rect 1830 1988 1831 1992
rect 1835 1988 1836 1992
rect 1830 1987 1836 1988
rect 1894 1992 1900 1993
rect 1894 1988 1895 1992
rect 1899 1988 1900 1992
rect 1894 1987 1900 1988
rect 1958 1992 1964 1993
rect 1958 1988 1959 1992
rect 1963 1988 1964 1992
rect 1958 1987 1964 1988
rect 2030 1992 2036 1993
rect 2030 1988 2031 1992
rect 2035 1988 2036 1992
rect 2504 1990 2506 1993
rect 2030 1987 2036 1988
rect 2502 1989 2508 1990
rect 2502 1985 2503 1989
rect 2507 1985 2508 1989
rect 2502 1984 2508 1985
rect 2502 1972 2508 1973
rect 1782 1971 1788 1972
rect 1782 1967 1783 1971
rect 1787 1967 1788 1971
rect 1782 1966 1788 1967
rect 1826 1971 1832 1972
rect 1826 1967 1827 1971
rect 1831 1967 1832 1971
rect 1826 1966 1832 1967
rect 1846 1971 1852 1972
rect 1846 1967 1847 1971
rect 1851 1967 1852 1971
rect 1846 1966 1852 1967
rect 1890 1971 1896 1972
rect 1890 1967 1891 1971
rect 1895 1967 1896 1971
rect 1890 1966 1896 1967
rect 1910 1971 1916 1972
rect 1910 1967 1911 1971
rect 1915 1967 1916 1971
rect 1910 1966 1916 1967
rect 1954 1971 1960 1972
rect 1954 1967 1955 1971
rect 1959 1967 1960 1971
rect 1954 1966 1960 1967
rect 1974 1971 1980 1972
rect 1974 1967 1975 1971
rect 1979 1967 1980 1971
rect 1974 1966 1980 1967
rect 2026 1971 2032 1972
rect 2026 1967 2027 1971
rect 2031 1967 2032 1971
rect 2026 1966 2032 1967
rect 2046 1971 2052 1972
rect 2046 1967 2047 1971
rect 2051 1967 2052 1971
rect 2046 1966 2052 1967
rect 2054 1971 2060 1972
rect 2054 1967 2055 1971
rect 2059 1967 2060 1971
rect 2502 1968 2503 1972
rect 2507 1968 2508 1972
rect 2502 1967 2508 1968
rect 2054 1966 2060 1967
rect 1774 1951 1780 1952
rect 1774 1947 1775 1951
rect 1779 1947 1780 1951
rect 1774 1946 1780 1947
rect 1784 1943 1786 1966
rect 1828 1952 1830 1966
rect 1826 1951 1832 1952
rect 1826 1947 1827 1951
rect 1831 1947 1832 1951
rect 1826 1946 1832 1947
rect 1848 1943 1850 1966
rect 1892 1952 1894 1966
rect 1890 1951 1896 1952
rect 1890 1947 1891 1951
rect 1895 1947 1896 1951
rect 1890 1946 1896 1947
rect 1912 1943 1914 1966
rect 1956 1952 1958 1966
rect 1954 1951 1960 1952
rect 1954 1947 1955 1951
rect 1959 1947 1960 1951
rect 1954 1946 1960 1947
rect 1976 1943 1978 1966
rect 2028 1952 2030 1966
rect 2026 1951 2032 1952
rect 2026 1947 2027 1951
rect 2031 1947 2032 1951
rect 2026 1946 2032 1947
rect 2048 1943 2050 1966
rect 2056 1944 2058 1966
rect 2054 1943 2060 1944
rect 2504 1943 2506 1967
rect 1719 1942 1723 1943
rect 1719 1937 1723 1938
rect 1775 1942 1779 1943
rect 1775 1937 1779 1938
rect 1783 1942 1787 1943
rect 1783 1937 1787 1938
rect 1847 1942 1851 1943
rect 1847 1937 1851 1938
rect 1911 1942 1915 1943
rect 1911 1937 1915 1938
rect 1919 1942 1923 1943
rect 1919 1937 1923 1938
rect 1975 1942 1979 1943
rect 1975 1937 1979 1938
rect 1999 1942 2003 1943
rect 1999 1937 2003 1938
rect 2047 1942 2051 1943
rect 2054 1939 2055 1943
rect 2059 1939 2060 1943
rect 2054 1938 2060 1939
rect 2087 1942 2091 1943
rect 2047 1937 2051 1938
rect 2087 1937 2091 1938
rect 2183 1942 2187 1943
rect 2183 1937 2187 1938
rect 2279 1942 2283 1943
rect 2279 1937 2283 1938
rect 2375 1942 2379 1943
rect 2375 1937 2379 1938
rect 2455 1942 2459 1943
rect 2455 1937 2459 1938
rect 2503 1942 2507 1943
rect 2503 1937 2507 1938
rect 1766 1935 1772 1936
rect 1766 1931 1767 1935
rect 1771 1931 1772 1935
rect 1766 1930 1772 1931
rect 1702 1912 1708 1913
rect 1710 1915 1716 1916
rect 1662 1910 1668 1911
rect 1710 1911 1711 1915
rect 1715 1911 1716 1915
rect 1710 1910 1716 1911
rect 1079 1902 1083 1903
rect 1079 1897 1083 1898
rect 1087 1902 1091 1903
rect 1087 1897 1091 1898
rect 1159 1902 1163 1903
rect 1159 1897 1163 1898
rect 1287 1902 1291 1903
rect 1287 1897 1291 1898
rect 1326 1899 1332 1900
rect 1086 1896 1092 1897
rect 1086 1892 1087 1896
rect 1091 1892 1092 1896
rect 1086 1891 1092 1892
rect 1158 1896 1164 1897
rect 1158 1892 1159 1896
rect 1163 1892 1164 1896
rect 1288 1894 1290 1897
rect 1326 1895 1327 1899
rect 1331 1895 1332 1899
rect 1326 1894 1332 1895
rect 1550 1896 1556 1897
rect 1158 1891 1164 1892
rect 1286 1893 1292 1894
rect 1286 1889 1287 1893
rect 1291 1889 1292 1893
rect 1286 1888 1292 1889
rect 1328 1887 1330 1894
rect 1550 1892 1551 1896
rect 1555 1892 1556 1896
rect 1550 1891 1556 1892
rect 1614 1896 1620 1897
rect 1614 1892 1615 1896
rect 1619 1892 1620 1896
rect 1614 1891 1620 1892
rect 1686 1896 1692 1897
rect 1686 1892 1687 1896
rect 1691 1892 1692 1896
rect 1686 1891 1692 1892
rect 1758 1896 1764 1897
rect 1758 1892 1759 1896
rect 1763 1892 1764 1896
rect 1758 1891 1764 1892
rect 1552 1887 1554 1891
rect 1616 1887 1618 1891
rect 1688 1887 1690 1891
rect 1760 1887 1762 1891
rect 1327 1886 1331 1887
rect 1327 1881 1331 1882
rect 1551 1886 1555 1887
rect 1551 1881 1555 1882
rect 1607 1886 1611 1887
rect 1607 1881 1611 1882
rect 1615 1886 1619 1887
rect 1615 1881 1619 1882
rect 1663 1886 1667 1887
rect 1663 1881 1667 1882
rect 1687 1886 1691 1887
rect 1687 1881 1691 1882
rect 1727 1886 1731 1887
rect 1727 1881 1731 1882
rect 1759 1886 1763 1887
rect 1759 1881 1763 1882
rect 1328 1878 1330 1881
rect 1606 1880 1612 1881
rect 1326 1877 1332 1878
rect 1286 1876 1292 1877
rect 794 1875 800 1876
rect 794 1871 795 1875
rect 799 1871 800 1875
rect 794 1870 800 1871
rect 814 1875 820 1876
rect 814 1871 815 1875
rect 819 1871 820 1875
rect 814 1870 820 1871
rect 866 1875 872 1876
rect 866 1871 867 1875
rect 871 1871 872 1875
rect 866 1870 872 1871
rect 886 1875 892 1876
rect 886 1871 887 1875
rect 891 1871 892 1875
rect 886 1870 892 1871
rect 938 1875 944 1876
rect 938 1871 939 1875
rect 943 1871 944 1875
rect 938 1870 944 1871
rect 958 1875 964 1876
rect 958 1871 959 1875
rect 963 1871 964 1875
rect 958 1870 964 1871
rect 1022 1875 1028 1876
rect 1022 1871 1023 1875
rect 1027 1871 1028 1875
rect 1022 1870 1028 1871
rect 1030 1875 1036 1876
rect 1030 1871 1031 1875
rect 1035 1871 1036 1875
rect 1030 1870 1036 1871
rect 1054 1875 1060 1876
rect 1054 1871 1055 1875
rect 1059 1871 1060 1875
rect 1054 1870 1060 1871
rect 1102 1875 1108 1876
rect 1102 1871 1103 1875
rect 1107 1871 1108 1875
rect 1102 1870 1108 1871
rect 1150 1875 1156 1876
rect 1150 1871 1151 1875
rect 1155 1871 1156 1875
rect 1150 1870 1156 1871
rect 1174 1875 1180 1876
rect 1174 1871 1175 1875
rect 1179 1871 1180 1875
rect 1286 1872 1287 1876
rect 1291 1872 1292 1876
rect 1326 1873 1327 1877
rect 1331 1873 1332 1877
rect 1606 1876 1607 1880
rect 1611 1876 1612 1880
rect 1606 1875 1612 1876
rect 1662 1880 1668 1881
rect 1662 1876 1663 1880
rect 1667 1876 1668 1880
rect 1662 1875 1668 1876
rect 1726 1880 1732 1881
rect 1726 1876 1727 1880
rect 1731 1876 1732 1880
rect 1726 1875 1732 1876
rect 1326 1872 1332 1873
rect 1286 1871 1292 1872
rect 1174 1870 1180 1871
rect 750 1863 756 1864
rect 750 1859 751 1863
rect 755 1859 756 1863
rect 750 1858 756 1859
rect 796 1856 798 1870
rect 794 1855 800 1856
rect 786 1851 792 1852
rect 591 1850 595 1851
rect 591 1845 595 1846
rect 647 1850 651 1851
rect 647 1845 651 1846
rect 687 1850 691 1851
rect 710 1850 716 1851
rect 735 1850 739 1851
rect 687 1845 691 1846
rect 574 1843 580 1844
rect 574 1839 575 1843
rect 579 1839 580 1843
rect 574 1838 580 1839
rect 592 1826 594 1845
rect 688 1826 690 1845
rect 494 1825 500 1826
rect 390 1820 396 1821
rect 410 1823 416 1824
rect 230 1818 236 1819
rect 410 1819 411 1823
rect 415 1819 416 1823
rect 494 1821 495 1825
rect 499 1821 500 1825
rect 590 1825 596 1826
rect 494 1820 500 1821
rect 510 1823 516 1824
rect 410 1818 416 1819
rect 510 1819 511 1823
rect 515 1819 516 1823
rect 590 1821 591 1825
rect 595 1821 596 1825
rect 686 1825 692 1826
rect 590 1820 596 1821
rect 614 1823 620 1824
rect 510 1818 516 1819
rect 614 1819 615 1823
rect 619 1819 620 1823
rect 686 1821 687 1825
rect 691 1821 692 1825
rect 712 1824 714 1850
rect 735 1845 739 1846
rect 775 1850 779 1851
rect 786 1847 787 1851
rect 791 1847 792 1851
rect 794 1851 795 1855
rect 799 1851 800 1855
rect 816 1851 818 1870
rect 868 1856 870 1870
rect 866 1855 872 1856
rect 866 1851 867 1855
rect 871 1851 872 1855
rect 888 1851 890 1870
rect 940 1856 942 1870
rect 938 1855 944 1856
rect 938 1851 939 1855
rect 943 1851 944 1855
rect 794 1850 800 1851
rect 815 1850 819 1851
rect 786 1846 792 1847
rect 775 1845 779 1846
rect 776 1826 778 1845
rect 774 1825 780 1826
rect 686 1820 692 1821
rect 710 1823 716 1824
rect 614 1818 620 1819
rect 710 1819 711 1823
rect 715 1819 716 1823
rect 774 1821 775 1825
rect 779 1821 780 1825
rect 788 1824 790 1846
rect 815 1845 819 1846
rect 855 1850 859 1851
rect 866 1850 872 1851
rect 887 1850 891 1851
rect 855 1845 859 1846
rect 887 1845 891 1846
rect 927 1850 931 1851
rect 938 1850 944 1851
rect 950 1855 956 1856
rect 950 1851 951 1855
rect 955 1851 956 1855
rect 960 1851 962 1870
rect 982 1867 988 1868
rect 982 1863 983 1867
rect 987 1863 988 1867
rect 982 1862 988 1863
rect 950 1850 956 1851
rect 959 1850 963 1851
rect 927 1845 931 1846
rect 830 1843 836 1844
rect 830 1839 831 1843
rect 835 1839 836 1843
rect 830 1838 836 1839
rect 774 1820 780 1821
rect 786 1823 792 1824
rect 710 1818 716 1819
rect 786 1819 787 1823
rect 791 1819 792 1823
rect 786 1818 792 1819
rect 110 1807 116 1808
rect 110 1803 111 1807
rect 115 1803 116 1807
rect 110 1802 116 1803
rect 134 1804 140 1805
rect 112 1787 114 1802
rect 134 1800 135 1804
rect 139 1800 140 1804
rect 134 1799 140 1800
rect 190 1804 196 1805
rect 190 1800 191 1804
rect 195 1800 196 1804
rect 190 1799 196 1800
rect 278 1804 284 1805
rect 278 1800 279 1804
rect 283 1800 284 1804
rect 278 1799 284 1800
rect 374 1804 380 1805
rect 374 1800 375 1804
rect 379 1800 380 1804
rect 374 1799 380 1800
rect 478 1804 484 1805
rect 478 1800 479 1804
rect 483 1800 484 1804
rect 478 1799 484 1800
rect 136 1787 138 1799
rect 192 1787 194 1799
rect 280 1787 282 1799
rect 376 1787 378 1799
rect 480 1787 482 1799
rect 111 1786 115 1787
rect 111 1781 115 1782
rect 135 1786 139 1787
rect 135 1781 139 1782
rect 191 1786 195 1787
rect 191 1781 195 1782
rect 199 1786 203 1787
rect 199 1781 203 1782
rect 279 1786 283 1787
rect 279 1781 283 1782
rect 295 1786 299 1787
rect 295 1781 299 1782
rect 375 1786 379 1787
rect 375 1781 379 1782
rect 399 1786 403 1787
rect 399 1781 403 1782
rect 479 1786 483 1787
rect 479 1781 483 1782
rect 503 1786 507 1787
rect 503 1781 507 1782
rect 112 1778 114 1781
rect 134 1780 140 1781
rect 110 1777 116 1778
rect 110 1773 111 1777
rect 115 1773 116 1777
rect 134 1776 135 1780
rect 139 1776 140 1780
rect 134 1775 140 1776
rect 198 1780 204 1781
rect 198 1776 199 1780
rect 203 1776 204 1780
rect 198 1775 204 1776
rect 294 1780 300 1781
rect 294 1776 295 1780
rect 299 1776 300 1780
rect 294 1775 300 1776
rect 398 1780 404 1781
rect 398 1776 399 1780
rect 403 1776 404 1780
rect 398 1775 404 1776
rect 502 1780 508 1781
rect 502 1776 503 1780
rect 507 1776 508 1780
rect 502 1775 508 1776
rect 512 1773 514 1818
rect 574 1804 580 1805
rect 574 1800 575 1804
rect 579 1800 580 1804
rect 574 1799 580 1800
rect 576 1787 578 1799
rect 575 1786 579 1787
rect 575 1781 579 1782
rect 607 1786 611 1787
rect 607 1781 611 1782
rect 606 1780 612 1781
rect 606 1776 607 1780
rect 611 1776 612 1780
rect 606 1775 612 1776
rect 110 1772 116 1773
rect 135 1772 139 1773
rect 135 1767 139 1768
rect 511 1772 515 1773
rect 511 1767 515 1768
rect 110 1760 116 1761
rect 110 1756 111 1760
rect 115 1756 116 1760
rect 110 1755 116 1756
rect 112 1731 114 1755
rect 136 1740 138 1767
rect 150 1759 156 1760
rect 150 1755 151 1759
rect 155 1755 156 1759
rect 150 1754 156 1755
rect 194 1759 200 1760
rect 194 1755 195 1759
rect 199 1755 200 1759
rect 194 1754 200 1755
rect 214 1759 220 1760
rect 214 1755 215 1759
rect 219 1755 220 1759
rect 214 1754 220 1755
rect 290 1759 296 1760
rect 290 1755 291 1759
rect 295 1755 296 1759
rect 290 1754 296 1755
rect 310 1759 316 1760
rect 310 1755 311 1759
rect 315 1755 316 1759
rect 310 1754 316 1755
rect 394 1759 400 1760
rect 394 1755 395 1759
rect 399 1755 400 1759
rect 394 1754 400 1755
rect 414 1759 420 1760
rect 414 1755 415 1759
rect 419 1755 420 1759
rect 414 1754 420 1755
rect 422 1759 428 1760
rect 422 1755 423 1759
rect 427 1755 428 1759
rect 422 1754 428 1755
rect 518 1759 524 1760
rect 518 1755 519 1759
rect 523 1755 524 1759
rect 518 1754 524 1755
rect 586 1759 592 1760
rect 586 1755 587 1759
rect 591 1755 592 1759
rect 586 1754 592 1755
rect 134 1739 140 1740
rect 134 1735 135 1739
rect 139 1735 140 1739
rect 134 1734 140 1735
rect 152 1731 154 1754
rect 196 1740 198 1754
rect 194 1739 200 1740
rect 194 1735 195 1739
rect 199 1735 200 1739
rect 194 1734 200 1735
rect 216 1731 218 1754
rect 292 1740 294 1754
rect 290 1739 296 1740
rect 290 1735 291 1739
rect 295 1735 296 1739
rect 290 1734 296 1735
rect 312 1731 314 1754
rect 396 1740 398 1754
rect 394 1739 400 1740
rect 394 1735 395 1739
rect 399 1735 400 1739
rect 394 1734 400 1735
rect 416 1731 418 1754
rect 424 1732 426 1754
rect 422 1731 428 1732
rect 520 1731 522 1754
rect 111 1730 115 1731
rect 111 1725 115 1726
rect 151 1730 155 1731
rect 151 1725 155 1726
rect 167 1730 171 1731
rect 167 1725 171 1726
rect 215 1730 219 1731
rect 215 1725 219 1726
rect 239 1730 243 1731
rect 239 1725 243 1726
rect 311 1730 315 1731
rect 311 1725 315 1726
rect 319 1730 323 1731
rect 319 1725 323 1726
rect 407 1730 411 1731
rect 407 1725 411 1726
rect 415 1730 419 1731
rect 422 1727 423 1731
rect 427 1727 428 1731
rect 422 1726 428 1727
rect 503 1730 507 1731
rect 415 1725 419 1726
rect 503 1725 507 1726
rect 519 1730 523 1731
rect 519 1725 523 1726
rect 112 1705 114 1725
rect 168 1706 170 1725
rect 190 1723 196 1724
rect 190 1719 191 1723
rect 195 1719 196 1723
rect 190 1718 196 1719
rect 166 1705 172 1706
rect 110 1704 116 1705
rect 110 1700 111 1704
rect 115 1700 116 1704
rect 166 1701 167 1705
rect 171 1701 172 1705
rect 192 1704 194 1718
rect 240 1706 242 1725
rect 262 1723 268 1724
rect 262 1719 263 1723
rect 267 1719 268 1723
rect 262 1718 268 1719
rect 238 1705 244 1706
rect 166 1700 172 1701
rect 190 1703 196 1704
rect 110 1699 116 1700
rect 190 1699 191 1703
rect 195 1699 196 1703
rect 238 1701 239 1705
rect 243 1701 244 1705
rect 264 1704 266 1718
rect 320 1706 322 1725
rect 342 1723 348 1724
rect 342 1719 343 1723
rect 347 1719 348 1723
rect 342 1718 348 1719
rect 318 1705 324 1706
rect 238 1700 244 1701
rect 262 1703 268 1704
rect 190 1698 196 1699
rect 262 1699 263 1703
rect 267 1699 268 1703
rect 318 1701 319 1705
rect 323 1701 324 1705
rect 344 1704 346 1718
rect 408 1706 410 1725
rect 430 1723 436 1724
rect 430 1719 431 1723
rect 435 1719 436 1723
rect 430 1718 436 1719
rect 406 1705 412 1706
rect 318 1700 324 1701
rect 342 1703 348 1704
rect 262 1698 268 1699
rect 342 1699 343 1703
rect 347 1699 348 1703
rect 406 1701 407 1705
rect 411 1701 412 1705
rect 432 1704 434 1718
rect 504 1706 506 1725
rect 588 1724 590 1754
rect 616 1740 618 1818
rect 670 1804 676 1805
rect 670 1800 671 1804
rect 675 1800 676 1804
rect 670 1799 676 1800
rect 758 1804 764 1805
rect 758 1800 759 1804
rect 763 1800 764 1804
rect 758 1799 764 1800
rect 672 1787 674 1799
rect 760 1787 762 1799
rect 671 1786 675 1787
rect 671 1781 675 1782
rect 703 1786 707 1787
rect 703 1781 707 1782
rect 759 1786 763 1787
rect 759 1781 763 1782
rect 799 1786 803 1787
rect 799 1781 803 1782
rect 702 1780 708 1781
rect 702 1776 703 1780
rect 707 1776 708 1780
rect 702 1775 708 1776
rect 798 1780 804 1781
rect 798 1776 799 1780
rect 803 1776 804 1780
rect 798 1775 804 1776
rect 832 1760 834 1838
rect 856 1826 858 1845
rect 918 1843 924 1844
rect 918 1839 919 1843
rect 923 1839 924 1843
rect 918 1838 924 1839
rect 854 1825 860 1826
rect 854 1821 855 1825
rect 859 1821 860 1825
rect 854 1820 860 1821
rect 838 1804 844 1805
rect 838 1800 839 1804
rect 843 1800 844 1804
rect 838 1799 844 1800
rect 910 1804 916 1805
rect 910 1800 911 1804
rect 915 1800 916 1804
rect 910 1799 916 1800
rect 840 1787 842 1799
rect 912 1787 914 1799
rect 839 1786 843 1787
rect 839 1781 843 1782
rect 887 1786 891 1787
rect 887 1781 891 1782
rect 911 1786 915 1787
rect 911 1781 915 1782
rect 886 1780 892 1781
rect 886 1776 887 1780
rect 891 1776 892 1780
rect 886 1775 892 1776
rect 920 1760 922 1838
rect 928 1826 930 1845
rect 926 1825 932 1826
rect 926 1821 927 1825
rect 931 1821 932 1825
rect 952 1824 954 1850
rect 959 1845 963 1846
rect 984 1844 986 1862
rect 1024 1856 1026 1870
rect 1022 1855 1028 1856
rect 1022 1851 1023 1855
rect 1027 1851 1028 1855
rect 1032 1851 1034 1870
rect 1104 1851 1106 1870
rect 1152 1856 1154 1870
rect 1150 1855 1156 1856
rect 1150 1851 1151 1855
rect 1155 1851 1156 1855
rect 1176 1851 1178 1870
rect 1288 1851 1290 1871
rect 1326 1860 1332 1861
rect 1768 1860 1770 1930
rect 1776 1918 1778 1937
rect 1814 1935 1820 1936
rect 1814 1931 1815 1935
rect 1819 1931 1820 1935
rect 1814 1930 1820 1931
rect 1774 1917 1780 1918
rect 1774 1913 1775 1917
rect 1779 1913 1780 1917
rect 1816 1916 1818 1930
rect 1848 1918 1850 1937
rect 1920 1918 1922 1937
rect 1942 1935 1948 1936
rect 1942 1931 1943 1935
rect 1947 1931 1948 1935
rect 1942 1930 1948 1931
rect 1846 1917 1852 1918
rect 1774 1912 1780 1913
rect 1814 1915 1820 1916
rect 1814 1911 1815 1915
rect 1819 1911 1820 1915
rect 1846 1913 1847 1917
rect 1851 1913 1852 1917
rect 1846 1912 1852 1913
rect 1918 1917 1924 1918
rect 1918 1913 1919 1917
rect 1923 1913 1924 1917
rect 1944 1916 1946 1930
rect 2000 1918 2002 1937
rect 2022 1935 2028 1936
rect 2022 1931 2023 1935
rect 2027 1931 2028 1935
rect 2022 1930 2028 1931
rect 1998 1917 2004 1918
rect 1918 1912 1924 1913
rect 1942 1915 1948 1916
rect 1814 1910 1820 1911
rect 1942 1911 1943 1915
rect 1947 1911 1948 1915
rect 1998 1913 1999 1917
rect 2003 1913 2004 1917
rect 2024 1916 2026 1930
rect 2088 1918 2090 1937
rect 2110 1935 2116 1936
rect 2110 1931 2111 1935
rect 2115 1931 2116 1935
rect 2110 1930 2116 1931
rect 2086 1917 2092 1918
rect 1998 1912 2004 1913
rect 2022 1915 2028 1916
rect 1942 1910 1948 1911
rect 2022 1911 2023 1915
rect 2027 1911 2028 1915
rect 2086 1913 2087 1917
rect 2091 1913 2092 1917
rect 2112 1916 2114 1930
rect 2184 1918 2186 1937
rect 2206 1935 2212 1936
rect 2206 1931 2207 1935
rect 2211 1931 2212 1935
rect 2206 1930 2212 1931
rect 2182 1917 2188 1918
rect 2086 1912 2092 1913
rect 2110 1915 2116 1916
rect 2022 1910 2028 1911
rect 2110 1911 2111 1915
rect 2115 1911 2116 1915
rect 2182 1913 2183 1917
rect 2187 1913 2188 1917
rect 2208 1916 2210 1930
rect 2280 1918 2282 1937
rect 2376 1918 2378 1937
rect 2398 1935 2404 1936
rect 2398 1931 2399 1935
rect 2403 1931 2404 1935
rect 2398 1930 2404 1931
rect 2278 1917 2284 1918
rect 2182 1912 2188 1913
rect 2206 1915 2212 1916
rect 2110 1910 2116 1911
rect 2206 1911 2207 1915
rect 2211 1911 2212 1915
rect 2278 1913 2279 1917
rect 2283 1913 2284 1917
rect 2374 1917 2380 1918
rect 2278 1912 2284 1913
rect 2286 1915 2292 1916
rect 2206 1910 2212 1911
rect 2286 1911 2287 1915
rect 2291 1911 2292 1915
rect 2374 1913 2375 1917
rect 2379 1913 2380 1917
rect 2400 1916 2402 1930
rect 2418 1927 2424 1928
rect 2418 1923 2419 1927
rect 2423 1923 2424 1927
rect 2418 1922 2424 1923
rect 2374 1912 2380 1913
rect 2398 1915 2404 1916
rect 2286 1910 2292 1911
rect 2398 1911 2399 1915
rect 2403 1911 2404 1915
rect 2398 1910 2404 1911
rect 1830 1896 1836 1897
rect 1830 1892 1831 1896
rect 1835 1892 1836 1896
rect 1830 1891 1836 1892
rect 1902 1896 1908 1897
rect 1902 1892 1903 1896
rect 1907 1892 1908 1896
rect 1902 1891 1908 1892
rect 1982 1896 1988 1897
rect 1982 1892 1983 1896
rect 1987 1892 1988 1896
rect 1982 1891 1988 1892
rect 2070 1896 2076 1897
rect 2070 1892 2071 1896
rect 2075 1892 2076 1896
rect 2070 1891 2076 1892
rect 2166 1896 2172 1897
rect 2166 1892 2167 1896
rect 2171 1892 2172 1896
rect 2166 1891 2172 1892
rect 2262 1896 2268 1897
rect 2262 1892 2263 1896
rect 2267 1892 2268 1896
rect 2262 1891 2268 1892
rect 1832 1887 1834 1891
rect 1904 1887 1906 1891
rect 1984 1887 1986 1891
rect 2072 1887 2074 1891
rect 2168 1887 2170 1891
rect 2264 1887 2266 1891
rect 1799 1886 1803 1887
rect 1799 1881 1803 1882
rect 1831 1886 1835 1887
rect 1831 1881 1835 1882
rect 1871 1886 1875 1887
rect 1871 1881 1875 1882
rect 1903 1886 1907 1887
rect 1903 1881 1907 1882
rect 1943 1886 1947 1887
rect 1943 1881 1947 1882
rect 1983 1886 1987 1887
rect 1983 1881 1987 1882
rect 2007 1886 2011 1887
rect 2007 1881 2011 1882
rect 2071 1886 2075 1887
rect 2071 1881 2075 1882
rect 2135 1886 2139 1887
rect 2135 1881 2139 1882
rect 2167 1886 2171 1887
rect 2167 1881 2171 1882
rect 2199 1886 2203 1887
rect 2199 1881 2203 1882
rect 2263 1886 2267 1887
rect 2263 1881 2267 1882
rect 1798 1880 1804 1881
rect 1798 1876 1799 1880
rect 1803 1876 1804 1880
rect 1798 1875 1804 1876
rect 1870 1880 1876 1881
rect 1870 1876 1871 1880
rect 1875 1876 1876 1880
rect 1870 1875 1876 1876
rect 1942 1880 1948 1881
rect 1942 1876 1943 1880
rect 1947 1876 1948 1880
rect 1942 1875 1948 1876
rect 2006 1880 2012 1881
rect 2006 1876 2007 1880
rect 2011 1876 2012 1880
rect 2006 1875 2012 1876
rect 2070 1880 2076 1881
rect 2070 1876 2071 1880
rect 2075 1876 2076 1880
rect 2070 1875 2076 1876
rect 2134 1880 2140 1881
rect 2134 1876 2135 1880
rect 2139 1876 2140 1880
rect 2134 1875 2140 1876
rect 2198 1880 2204 1881
rect 2198 1876 2199 1880
rect 2203 1876 2204 1880
rect 2198 1875 2204 1876
rect 2262 1880 2268 1881
rect 2262 1876 2263 1880
rect 2267 1876 2268 1880
rect 2262 1875 2268 1876
rect 1326 1856 1327 1860
rect 1331 1856 1332 1860
rect 1326 1855 1332 1856
rect 1622 1859 1628 1860
rect 1622 1855 1623 1859
rect 1627 1855 1628 1859
rect 999 1850 1003 1851
rect 1022 1850 1028 1851
rect 1031 1850 1035 1851
rect 999 1845 1003 1846
rect 1031 1845 1035 1846
rect 1079 1850 1083 1851
rect 1079 1845 1083 1846
rect 1103 1850 1107 1851
rect 1150 1850 1156 1851
rect 1159 1850 1163 1851
rect 1103 1845 1107 1846
rect 1159 1845 1163 1846
rect 1175 1850 1179 1851
rect 1175 1845 1179 1846
rect 1287 1850 1291 1851
rect 1287 1845 1291 1846
rect 982 1843 988 1844
rect 982 1839 983 1843
rect 987 1839 988 1843
rect 982 1838 988 1839
rect 1000 1826 1002 1845
rect 1022 1843 1028 1844
rect 1022 1839 1023 1843
rect 1027 1839 1028 1843
rect 1022 1838 1028 1839
rect 998 1825 1004 1826
rect 926 1820 932 1821
rect 950 1823 956 1824
rect 950 1819 951 1823
rect 955 1819 956 1823
rect 998 1821 999 1825
rect 1003 1821 1004 1825
rect 1024 1824 1026 1838
rect 1080 1826 1082 1845
rect 1110 1843 1116 1844
rect 1110 1839 1111 1843
rect 1115 1839 1116 1843
rect 1110 1838 1116 1839
rect 1078 1825 1084 1826
rect 998 1820 1004 1821
rect 1022 1823 1028 1824
rect 950 1818 956 1819
rect 1022 1819 1023 1823
rect 1027 1819 1028 1823
rect 1078 1821 1079 1825
rect 1083 1821 1084 1825
rect 1112 1824 1114 1838
rect 1160 1826 1162 1845
rect 1158 1825 1164 1826
rect 1288 1825 1290 1845
rect 1328 1831 1330 1855
rect 1622 1854 1628 1855
rect 1658 1859 1664 1860
rect 1658 1855 1659 1859
rect 1663 1855 1664 1859
rect 1658 1854 1664 1855
rect 1678 1859 1684 1860
rect 1678 1855 1679 1859
rect 1683 1855 1684 1859
rect 1678 1854 1684 1855
rect 1722 1859 1728 1860
rect 1722 1855 1723 1859
rect 1727 1855 1728 1859
rect 1722 1854 1728 1855
rect 1742 1859 1748 1860
rect 1742 1855 1743 1859
rect 1747 1855 1748 1859
rect 1742 1854 1748 1855
rect 1766 1859 1772 1860
rect 1766 1855 1767 1859
rect 1771 1855 1772 1859
rect 1766 1854 1772 1855
rect 1814 1859 1820 1860
rect 1814 1855 1815 1859
rect 1819 1855 1820 1859
rect 1814 1854 1820 1855
rect 1886 1859 1892 1860
rect 1886 1855 1887 1859
rect 1891 1855 1892 1859
rect 1886 1854 1892 1855
rect 1894 1859 1900 1860
rect 1894 1855 1895 1859
rect 1899 1855 1900 1859
rect 1894 1854 1900 1855
rect 1958 1859 1964 1860
rect 1958 1855 1959 1859
rect 1963 1855 1964 1859
rect 1958 1854 1964 1855
rect 2022 1859 2028 1860
rect 2022 1855 2023 1859
rect 2027 1855 2028 1859
rect 2022 1854 2028 1855
rect 2066 1859 2072 1860
rect 2066 1855 2067 1859
rect 2071 1855 2072 1859
rect 2066 1854 2072 1855
rect 2086 1859 2092 1860
rect 2086 1855 2087 1859
rect 2091 1855 2092 1859
rect 2086 1854 2092 1855
rect 2130 1859 2136 1860
rect 2130 1855 2131 1859
rect 2135 1855 2136 1859
rect 2130 1854 2136 1855
rect 2150 1859 2156 1860
rect 2150 1855 2151 1859
rect 2155 1855 2156 1859
rect 2150 1854 2156 1855
rect 2194 1859 2200 1860
rect 2194 1855 2195 1859
rect 2199 1855 2200 1859
rect 2194 1854 2200 1855
rect 2214 1859 2220 1860
rect 2214 1855 2215 1859
rect 2219 1855 2220 1859
rect 2214 1854 2220 1855
rect 2258 1859 2264 1860
rect 2258 1855 2259 1859
rect 2263 1855 2264 1859
rect 2258 1854 2264 1855
rect 2278 1859 2284 1860
rect 2278 1855 2279 1859
rect 2283 1855 2284 1859
rect 2278 1854 2284 1855
rect 1624 1831 1626 1854
rect 1660 1840 1662 1854
rect 1658 1839 1664 1840
rect 1658 1835 1659 1839
rect 1663 1835 1664 1839
rect 1658 1834 1664 1835
rect 1680 1831 1682 1854
rect 1724 1840 1726 1854
rect 1722 1839 1728 1840
rect 1722 1835 1723 1839
rect 1727 1835 1728 1839
rect 1722 1834 1728 1835
rect 1744 1831 1746 1854
rect 1816 1831 1818 1854
rect 1888 1831 1890 1854
rect 1896 1836 1898 1854
rect 1894 1835 1900 1836
rect 1894 1831 1895 1835
rect 1899 1831 1900 1835
rect 1960 1831 1962 1854
rect 1970 1839 1976 1840
rect 1970 1835 1971 1839
rect 1975 1835 1976 1839
rect 1970 1834 1976 1835
rect 1327 1830 1331 1831
rect 1327 1825 1331 1826
rect 1623 1830 1627 1831
rect 1623 1825 1627 1826
rect 1631 1830 1635 1831
rect 1631 1825 1635 1826
rect 1679 1830 1683 1831
rect 1679 1825 1683 1826
rect 1719 1830 1723 1831
rect 1719 1825 1723 1826
rect 1743 1830 1747 1831
rect 1743 1825 1747 1826
rect 1815 1830 1819 1831
rect 1815 1825 1819 1826
rect 1887 1830 1891 1831
rect 1894 1830 1900 1831
rect 1927 1830 1931 1831
rect 1887 1825 1891 1826
rect 1927 1825 1931 1826
rect 1959 1830 1963 1831
rect 1959 1825 1963 1826
rect 1078 1820 1084 1821
rect 1110 1823 1116 1824
rect 1022 1818 1028 1819
rect 1110 1819 1111 1823
rect 1115 1819 1116 1823
rect 1158 1821 1159 1825
rect 1163 1821 1164 1825
rect 1286 1824 1292 1825
rect 1158 1820 1164 1821
rect 1174 1823 1180 1824
rect 1110 1818 1116 1819
rect 1174 1819 1175 1823
rect 1179 1819 1180 1823
rect 1286 1820 1287 1824
rect 1291 1820 1292 1824
rect 1286 1819 1292 1820
rect 1174 1818 1180 1819
rect 982 1804 988 1805
rect 982 1800 983 1804
rect 987 1800 988 1804
rect 982 1799 988 1800
rect 1062 1804 1068 1805
rect 1062 1800 1063 1804
rect 1067 1800 1068 1804
rect 1062 1799 1068 1800
rect 1142 1804 1148 1805
rect 1142 1800 1143 1804
rect 1147 1800 1148 1804
rect 1142 1799 1148 1800
rect 984 1787 986 1799
rect 1064 1787 1066 1799
rect 1144 1787 1146 1799
rect 975 1786 979 1787
rect 975 1781 979 1782
rect 983 1786 987 1787
rect 983 1781 987 1782
rect 1063 1786 1067 1787
rect 1063 1781 1067 1782
rect 1143 1786 1147 1787
rect 1143 1781 1147 1782
rect 1151 1786 1155 1787
rect 1151 1781 1155 1782
rect 974 1780 980 1781
rect 974 1776 975 1780
rect 979 1776 980 1780
rect 974 1775 980 1776
rect 1062 1780 1068 1781
rect 1062 1776 1063 1780
rect 1067 1776 1068 1780
rect 1062 1775 1068 1776
rect 1150 1780 1156 1781
rect 1150 1776 1151 1780
rect 1155 1776 1156 1780
rect 1150 1775 1156 1776
rect 622 1759 628 1760
rect 622 1755 623 1759
rect 627 1755 628 1759
rect 622 1754 628 1755
rect 718 1759 724 1760
rect 718 1755 719 1759
rect 723 1755 724 1759
rect 718 1754 724 1755
rect 794 1759 800 1760
rect 794 1755 795 1759
rect 799 1755 800 1759
rect 794 1754 800 1755
rect 814 1759 820 1760
rect 814 1755 815 1759
rect 819 1755 820 1759
rect 814 1754 820 1755
rect 830 1759 836 1760
rect 830 1755 831 1759
rect 835 1755 836 1759
rect 830 1754 836 1755
rect 902 1759 908 1760
rect 902 1755 903 1759
rect 907 1755 908 1759
rect 902 1754 908 1755
rect 918 1759 924 1760
rect 918 1755 919 1759
rect 923 1755 924 1759
rect 918 1754 924 1755
rect 990 1759 996 1760
rect 990 1755 991 1759
rect 995 1755 996 1759
rect 990 1754 996 1755
rect 1026 1759 1032 1760
rect 1026 1755 1027 1759
rect 1031 1755 1032 1759
rect 1026 1754 1032 1755
rect 1078 1759 1084 1760
rect 1078 1755 1079 1759
rect 1083 1755 1084 1759
rect 1078 1754 1084 1755
rect 1166 1759 1172 1760
rect 1166 1755 1167 1759
rect 1171 1755 1172 1759
rect 1166 1754 1172 1755
rect 614 1739 620 1740
rect 614 1735 615 1739
rect 619 1735 620 1739
rect 614 1734 620 1735
rect 624 1731 626 1754
rect 720 1731 722 1754
rect 796 1740 798 1754
rect 730 1739 736 1740
rect 730 1735 731 1739
rect 735 1735 736 1739
rect 730 1734 736 1735
rect 794 1739 800 1740
rect 794 1735 795 1739
rect 799 1735 800 1739
rect 794 1734 800 1735
rect 607 1730 611 1731
rect 607 1725 611 1726
rect 623 1730 627 1731
rect 623 1725 627 1726
rect 711 1730 715 1731
rect 711 1725 715 1726
rect 719 1730 723 1731
rect 719 1725 723 1726
rect 586 1723 592 1724
rect 586 1719 587 1723
rect 591 1719 592 1723
rect 586 1718 592 1719
rect 608 1706 610 1725
rect 712 1706 714 1725
rect 502 1705 508 1706
rect 406 1700 412 1701
rect 430 1703 436 1704
rect 342 1698 348 1699
rect 430 1699 431 1703
rect 435 1699 436 1703
rect 502 1701 503 1705
rect 507 1701 508 1705
rect 606 1705 612 1706
rect 502 1700 508 1701
rect 510 1703 516 1704
rect 430 1698 436 1699
rect 510 1699 511 1703
rect 515 1699 516 1703
rect 606 1701 607 1705
rect 611 1701 612 1705
rect 710 1705 716 1706
rect 606 1700 612 1701
rect 614 1703 620 1704
rect 510 1698 516 1699
rect 614 1699 615 1703
rect 619 1699 620 1703
rect 710 1701 711 1705
rect 715 1701 716 1705
rect 732 1704 734 1734
rect 816 1731 818 1754
rect 904 1731 906 1754
rect 954 1739 960 1740
rect 954 1735 955 1739
rect 959 1735 960 1739
rect 954 1734 960 1735
rect 815 1730 819 1731
rect 815 1725 819 1726
rect 823 1730 827 1731
rect 823 1725 827 1726
rect 903 1730 907 1731
rect 903 1725 907 1726
rect 935 1730 939 1731
rect 935 1725 939 1726
rect 798 1723 804 1724
rect 798 1719 799 1723
rect 803 1719 804 1723
rect 798 1718 804 1719
rect 710 1700 716 1701
rect 730 1703 736 1704
rect 614 1698 620 1699
rect 730 1699 731 1703
rect 735 1699 736 1703
rect 730 1698 736 1699
rect 110 1687 116 1688
rect 110 1683 111 1687
rect 115 1683 116 1687
rect 110 1682 116 1683
rect 150 1684 156 1685
rect 112 1675 114 1682
rect 150 1680 151 1684
rect 155 1680 156 1684
rect 150 1679 156 1680
rect 222 1684 228 1685
rect 222 1680 223 1684
rect 227 1680 228 1684
rect 222 1679 228 1680
rect 302 1684 308 1685
rect 302 1680 303 1684
rect 307 1680 308 1684
rect 302 1679 308 1680
rect 390 1684 396 1685
rect 390 1680 391 1684
rect 395 1680 396 1684
rect 390 1679 396 1680
rect 486 1684 492 1685
rect 486 1680 487 1684
rect 491 1680 492 1684
rect 486 1679 492 1680
rect 152 1675 154 1679
rect 224 1675 226 1679
rect 304 1675 306 1679
rect 392 1675 394 1679
rect 488 1675 490 1679
rect 111 1674 115 1675
rect 111 1669 115 1670
rect 151 1674 155 1675
rect 151 1669 155 1670
rect 223 1674 227 1675
rect 223 1669 227 1670
rect 255 1674 259 1675
rect 255 1669 259 1670
rect 303 1674 307 1675
rect 303 1669 307 1670
rect 319 1674 323 1675
rect 319 1669 323 1670
rect 391 1674 395 1675
rect 391 1669 395 1670
rect 399 1674 403 1675
rect 399 1669 403 1670
rect 487 1674 491 1675
rect 487 1669 491 1670
rect 112 1666 114 1669
rect 254 1668 260 1669
rect 110 1665 116 1666
rect 110 1661 111 1665
rect 115 1661 116 1665
rect 254 1664 255 1668
rect 259 1664 260 1668
rect 254 1663 260 1664
rect 318 1668 324 1669
rect 318 1664 319 1668
rect 323 1664 324 1668
rect 318 1663 324 1664
rect 398 1668 404 1669
rect 398 1664 399 1668
rect 403 1664 404 1668
rect 398 1663 404 1664
rect 486 1668 492 1669
rect 486 1664 487 1668
rect 491 1664 492 1668
rect 486 1663 492 1664
rect 110 1660 116 1661
rect 110 1648 116 1649
rect 110 1644 111 1648
rect 115 1644 116 1648
rect 110 1643 116 1644
rect 270 1647 276 1648
rect 270 1643 271 1647
rect 275 1643 276 1647
rect 112 1619 114 1643
rect 270 1642 276 1643
rect 314 1647 320 1648
rect 314 1643 315 1647
rect 319 1643 320 1647
rect 314 1642 320 1643
rect 334 1647 340 1648
rect 334 1643 335 1647
rect 339 1643 340 1647
rect 334 1642 340 1643
rect 394 1647 400 1648
rect 394 1643 395 1647
rect 399 1643 400 1647
rect 394 1642 400 1643
rect 414 1647 420 1648
rect 414 1643 415 1647
rect 419 1643 420 1647
rect 414 1642 420 1643
rect 482 1647 488 1648
rect 482 1643 483 1647
rect 487 1643 488 1647
rect 482 1642 488 1643
rect 502 1647 508 1648
rect 502 1643 503 1647
rect 507 1643 508 1647
rect 502 1642 508 1643
rect 272 1619 274 1642
rect 316 1628 318 1642
rect 314 1627 320 1628
rect 314 1623 315 1627
rect 319 1623 320 1627
rect 314 1622 320 1623
rect 336 1619 338 1642
rect 396 1628 398 1642
rect 394 1627 400 1628
rect 394 1623 395 1627
rect 399 1623 400 1627
rect 394 1622 400 1623
rect 416 1619 418 1642
rect 484 1628 486 1642
rect 482 1627 488 1628
rect 482 1623 483 1627
rect 487 1623 488 1627
rect 482 1622 488 1623
rect 504 1619 506 1642
rect 512 1636 514 1698
rect 590 1684 596 1685
rect 590 1680 591 1684
rect 595 1680 596 1684
rect 590 1679 596 1680
rect 592 1675 594 1679
rect 575 1674 579 1675
rect 575 1669 579 1670
rect 591 1674 595 1675
rect 591 1669 595 1670
rect 574 1668 580 1669
rect 574 1664 575 1668
rect 579 1664 580 1668
rect 574 1663 580 1664
rect 518 1647 524 1648
rect 518 1643 519 1647
rect 523 1643 524 1647
rect 518 1642 524 1643
rect 590 1647 596 1648
rect 590 1643 591 1647
rect 595 1643 596 1647
rect 590 1642 596 1643
rect 606 1647 612 1648
rect 606 1643 607 1647
rect 611 1643 612 1647
rect 606 1642 612 1643
rect 510 1635 516 1636
rect 510 1631 511 1635
rect 515 1631 516 1635
rect 510 1630 516 1631
rect 520 1620 522 1642
rect 518 1619 524 1620
rect 592 1619 594 1642
rect 111 1618 115 1619
rect 111 1613 115 1614
rect 271 1618 275 1619
rect 271 1613 275 1614
rect 303 1618 307 1619
rect 303 1613 307 1614
rect 335 1618 339 1619
rect 335 1613 339 1614
rect 359 1618 363 1619
rect 359 1613 363 1614
rect 415 1618 419 1619
rect 415 1613 419 1614
rect 431 1618 435 1619
rect 431 1613 435 1614
rect 503 1618 507 1619
rect 503 1613 507 1614
rect 511 1618 515 1619
rect 518 1615 519 1619
rect 523 1615 524 1619
rect 518 1614 524 1615
rect 591 1618 595 1619
rect 511 1613 515 1614
rect 591 1613 595 1614
rect 599 1618 603 1619
rect 599 1613 603 1614
rect 112 1593 114 1613
rect 254 1599 260 1600
rect 254 1595 255 1599
rect 259 1595 260 1599
rect 254 1594 260 1595
rect 304 1594 306 1613
rect 326 1611 332 1612
rect 326 1607 327 1611
rect 331 1607 332 1611
rect 326 1606 332 1607
rect 110 1592 116 1593
rect 110 1588 111 1592
rect 115 1588 116 1592
rect 110 1587 116 1588
rect 110 1575 116 1576
rect 110 1571 111 1575
rect 115 1571 116 1575
rect 110 1570 116 1571
rect 112 1567 114 1570
rect 111 1566 115 1567
rect 111 1561 115 1562
rect 247 1566 251 1567
rect 247 1561 251 1562
rect 112 1558 114 1561
rect 246 1560 252 1561
rect 110 1557 116 1558
rect 110 1553 111 1557
rect 115 1553 116 1557
rect 246 1556 247 1560
rect 251 1556 252 1560
rect 246 1555 252 1556
rect 110 1552 116 1553
rect 110 1540 116 1541
rect 110 1536 111 1540
rect 115 1536 116 1540
rect 110 1535 116 1536
rect 112 1507 114 1535
rect 256 1520 258 1594
rect 302 1593 308 1594
rect 302 1589 303 1593
rect 307 1589 308 1593
rect 328 1592 330 1606
rect 360 1594 362 1613
rect 382 1611 388 1612
rect 382 1607 383 1611
rect 387 1607 388 1611
rect 382 1606 388 1607
rect 358 1593 364 1594
rect 302 1588 308 1589
rect 326 1591 332 1592
rect 326 1587 327 1591
rect 331 1587 332 1591
rect 358 1589 359 1593
rect 363 1589 364 1593
rect 384 1592 386 1606
rect 432 1594 434 1613
rect 512 1594 514 1613
rect 600 1594 602 1613
rect 608 1612 610 1642
rect 616 1628 618 1698
rect 694 1684 700 1685
rect 694 1680 695 1684
rect 699 1680 700 1684
rect 694 1679 700 1680
rect 696 1675 698 1679
rect 671 1674 675 1675
rect 671 1669 675 1670
rect 695 1674 699 1675
rect 695 1669 699 1670
rect 767 1674 771 1675
rect 767 1669 771 1670
rect 670 1668 676 1669
rect 670 1664 671 1668
rect 675 1664 676 1668
rect 670 1663 676 1664
rect 766 1668 772 1669
rect 766 1664 767 1668
rect 771 1664 772 1668
rect 766 1663 772 1664
rect 800 1648 802 1718
rect 824 1706 826 1725
rect 910 1723 916 1724
rect 910 1719 911 1723
rect 915 1719 916 1723
rect 910 1718 916 1719
rect 822 1705 828 1706
rect 822 1701 823 1705
rect 827 1701 828 1705
rect 822 1700 828 1701
rect 806 1684 812 1685
rect 806 1680 807 1684
rect 811 1680 812 1684
rect 806 1679 812 1680
rect 808 1675 810 1679
rect 807 1674 811 1675
rect 807 1669 811 1670
rect 863 1674 867 1675
rect 863 1669 867 1670
rect 862 1668 868 1669
rect 862 1664 863 1668
rect 867 1664 868 1668
rect 862 1663 868 1664
rect 912 1648 914 1718
rect 936 1706 938 1725
rect 934 1705 940 1706
rect 934 1701 935 1705
rect 939 1701 940 1705
rect 956 1704 958 1734
rect 992 1731 994 1754
rect 991 1730 995 1731
rect 991 1725 995 1726
rect 1028 1724 1030 1754
rect 1080 1731 1082 1754
rect 1168 1731 1170 1754
rect 1176 1740 1178 1818
rect 1286 1807 1292 1808
rect 1286 1803 1287 1807
rect 1291 1803 1292 1807
rect 1328 1805 1330 1825
rect 1632 1806 1634 1825
rect 1654 1823 1660 1824
rect 1654 1819 1655 1823
rect 1659 1819 1660 1823
rect 1654 1818 1660 1819
rect 1662 1823 1668 1824
rect 1662 1819 1663 1823
rect 1667 1819 1668 1823
rect 1662 1818 1668 1819
rect 1630 1805 1636 1806
rect 1286 1802 1292 1803
rect 1326 1804 1332 1805
rect 1288 1787 1290 1802
rect 1326 1800 1327 1804
rect 1331 1800 1332 1804
rect 1630 1801 1631 1805
rect 1635 1801 1636 1805
rect 1630 1800 1636 1801
rect 1326 1799 1332 1800
rect 1326 1787 1332 1788
rect 1287 1786 1291 1787
rect 1326 1783 1327 1787
rect 1331 1783 1332 1787
rect 1326 1782 1332 1783
rect 1614 1784 1620 1785
rect 1287 1781 1291 1782
rect 1288 1778 1290 1781
rect 1328 1779 1330 1782
rect 1614 1780 1615 1784
rect 1619 1780 1620 1784
rect 1614 1779 1620 1780
rect 1327 1778 1331 1779
rect 1286 1777 1292 1778
rect 1286 1773 1287 1777
rect 1291 1773 1292 1777
rect 1327 1773 1331 1774
rect 1527 1778 1531 1779
rect 1527 1773 1531 1774
rect 1607 1778 1611 1779
rect 1607 1773 1611 1774
rect 1615 1778 1619 1779
rect 1615 1773 1619 1774
rect 1286 1772 1292 1773
rect 1328 1770 1330 1773
rect 1526 1772 1532 1773
rect 1326 1769 1332 1770
rect 1326 1765 1327 1769
rect 1331 1765 1332 1769
rect 1526 1768 1527 1772
rect 1531 1768 1532 1772
rect 1526 1767 1532 1768
rect 1606 1772 1612 1773
rect 1606 1768 1607 1772
rect 1611 1768 1612 1772
rect 1606 1767 1612 1768
rect 1326 1764 1332 1765
rect 1286 1760 1292 1761
rect 1286 1756 1287 1760
rect 1291 1756 1292 1760
rect 1656 1757 1658 1818
rect 1664 1804 1666 1818
rect 1720 1806 1722 1825
rect 1750 1823 1756 1824
rect 1750 1819 1751 1823
rect 1755 1819 1756 1823
rect 1750 1818 1756 1819
rect 1718 1805 1724 1806
rect 1662 1803 1668 1804
rect 1662 1799 1663 1803
rect 1667 1799 1668 1803
rect 1718 1801 1719 1805
rect 1723 1801 1724 1805
rect 1752 1804 1754 1818
rect 1816 1806 1818 1825
rect 1928 1806 1930 1825
rect 1972 1812 1974 1834
rect 2024 1831 2026 1854
rect 2068 1840 2070 1854
rect 2066 1839 2072 1840
rect 2066 1835 2067 1839
rect 2071 1835 2072 1839
rect 2066 1834 2072 1835
rect 2088 1831 2090 1854
rect 2132 1840 2134 1854
rect 2130 1839 2136 1840
rect 2130 1835 2131 1839
rect 2135 1835 2136 1839
rect 2130 1834 2136 1835
rect 2152 1831 2154 1854
rect 2196 1840 2198 1854
rect 2194 1839 2200 1840
rect 2194 1835 2195 1839
rect 2199 1835 2200 1839
rect 2194 1834 2200 1835
rect 2216 1831 2218 1854
rect 2260 1840 2262 1854
rect 2258 1839 2264 1840
rect 2258 1835 2259 1839
rect 2263 1835 2264 1839
rect 2258 1834 2264 1835
rect 2280 1831 2282 1854
rect 2288 1848 2290 1910
rect 2358 1896 2364 1897
rect 2358 1892 2359 1896
rect 2363 1892 2364 1896
rect 2358 1891 2364 1892
rect 2360 1887 2362 1891
rect 2327 1886 2331 1887
rect 2327 1881 2331 1882
rect 2359 1886 2363 1887
rect 2359 1881 2363 1882
rect 2383 1886 2387 1887
rect 2383 1881 2387 1882
rect 2326 1880 2332 1881
rect 2326 1876 2327 1880
rect 2331 1876 2332 1880
rect 2326 1875 2332 1876
rect 2382 1880 2388 1881
rect 2382 1876 2383 1880
rect 2387 1876 2388 1880
rect 2382 1875 2388 1876
rect 2420 1860 2422 1922
rect 2456 1918 2458 1937
rect 2454 1917 2460 1918
rect 2504 1917 2506 1937
rect 2454 1913 2455 1917
rect 2459 1913 2460 1917
rect 2502 1916 2508 1917
rect 2454 1912 2460 1913
rect 2470 1915 2476 1916
rect 2470 1911 2471 1915
rect 2475 1911 2476 1915
rect 2502 1912 2503 1916
rect 2507 1912 2508 1916
rect 2502 1911 2508 1912
rect 2470 1910 2476 1911
rect 2438 1896 2444 1897
rect 2438 1892 2439 1896
rect 2443 1892 2444 1896
rect 2438 1891 2444 1892
rect 2440 1887 2442 1891
rect 2439 1886 2443 1887
rect 2439 1881 2443 1882
rect 2438 1880 2444 1881
rect 2438 1876 2439 1880
rect 2443 1876 2444 1880
rect 2438 1875 2444 1876
rect 2322 1859 2328 1860
rect 2322 1855 2323 1859
rect 2327 1855 2328 1859
rect 2322 1854 2328 1855
rect 2342 1859 2348 1860
rect 2342 1855 2343 1859
rect 2347 1855 2348 1859
rect 2342 1854 2348 1855
rect 2378 1859 2384 1860
rect 2378 1855 2379 1859
rect 2383 1855 2384 1859
rect 2378 1854 2384 1855
rect 2398 1859 2404 1860
rect 2398 1855 2399 1859
rect 2403 1855 2404 1859
rect 2398 1854 2404 1855
rect 2418 1859 2424 1860
rect 2418 1855 2419 1859
rect 2423 1855 2424 1859
rect 2418 1854 2424 1855
rect 2454 1859 2460 1860
rect 2454 1855 2455 1859
rect 2459 1855 2460 1859
rect 2454 1854 2460 1855
rect 2462 1859 2468 1860
rect 2462 1855 2463 1859
rect 2467 1855 2468 1859
rect 2462 1854 2468 1855
rect 2286 1847 2292 1848
rect 2286 1843 2287 1847
rect 2291 1843 2292 1847
rect 2286 1842 2292 1843
rect 2324 1840 2326 1854
rect 2322 1839 2328 1840
rect 2322 1835 2323 1839
rect 2327 1835 2328 1839
rect 2322 1834 2328 1835
rect 2344 1831 2346 1854
rect 2380 1840 2382 1854
rect 2378 1839 2384 1840
rect 2378 1835 2379 1839
rect 2383 1835 2384 1839
rect 2378 1834 2384 1835
rect 2400 1831 2402 1854
rect 2456 1831 2458 1854
rect 2023 1830 2027 1831
rect 2023 1825 2027 1826
rect 2055 1830 2059 1831
rect 2055 1825 2059 1826
rect 2087 1830 2091 1831
rect 2087 1825 2091 1826
rect 2151 1830 2155 1831
rect 2151 1825 2155 1826
rect 2191 1830 2195 1831
rect 2191 1825 2195 1826
rect 2215 1830 2219 1831
rect 2215 1825 2219 1826
rect 2279 1830 2283 1831
rect 2279 1825 2283 1826
rect 2335 1830 2339 1831
rect 2335 1825 2339 1826
rect 2343 1830 2347 1831
rect 2343 1825 2347 1826
rect 2399 1830 2403 1831
rect 2399 1825 2403 1826
rect 2455 1830 2459 1831
rect 2455 1825 2459 1826
rect 1970 1811 1976 1812
rect 1970 1807 1971 1811
rect 1975 1807 1976 1811
rect 1970 1806 1976 1807
rect 2056 1806 2058 1825
rect 2192 1806 2194 1825
rect 2326 1823 2332 1824
rect 2326 1819 2327 1823
rect 2331 1819 2332 1823
rect 2326 1818 2332 1819
rect 1814 1805 1820 1806
rect 1718 1800 1724 1801
rect 1750 1803 1756 1804
rect 1662 1798 1668 1799
rect 1750 1799 1751 1803
rect 1755 1799 1756 1803
rect 1814 1801 1815 1805
rect 1819 1801 1820 1805
rect 1814 1800 1820 1801
rect 1926 1805 1932 1806
rect 1926 1801 1927 1805
rect 1931 1801 1932 1805
rect 1926 1800 1932 1801
rect 2054 1805 2060 1806
rect 2054 1801 2055 1805
rect 2059 1801 2060 1805
rect 2054 1800 2060 1801
rect 2190 1805 2196 1806
rect 2190 1801 2191 1805
rect 2195 1801 2196 1805
rect 2190 1800 2196 1801
rect 2206 1803 2212 1804
rect 1750 1798 1756 1799
rect 2206 1799 2207 1803
rect 2211 1799 2212 1803
rect 2206 1798 2212 1799
rect 1702 1784 1708 1785
rect 1702 1780 1703 1784
rect 1707 1780 1708 1784
rect 1702 1779 1708 1780
rect 1798 1784 1804 1785
rect 1798 1780 1799 1784
rect 1803 1780 1804 1784
rect 1798 1779 1804 1780
rect 1910 1784 1916 1785
rect 1910 1780 1911 1784
rect 1915 1780 1916 1784
rect 1910 1779 1916 1780
rect 2038 1784 2044 1785
rect 2038 1780 2039 1784
rect 2043 1780 2044 1784
rect 2038 1779 2044 1780
rect 2174 1784 2180 1785
rect 2174 1780 2175 1784
rect 2179 1780 2180 1784
rect 2174 1779 2180 1780
rect 1695 1778 1699 1779
rect 1695 1773 1699 1774
rect 1703 1778 1707 1779
rect 1703 1773 1707 1774
rect 1791 1778 1795 1779
rect 1791 1773 1795 1774
rect 1799 1778 1803 1779
rect 1799 1773 1803 1774
rect 1879 1778 1883 1779
rect 1879 1773 1883 1774
rect 1911 1778 1915 1779
rect 1911 1773 1915 1774
rect 1967 1778 1971 1779
rect 1967 1773 1971 1774
rect 2039 1778 2043 1779
rect 2039 1773 2043 1774
rect 2055 1778 2059 1779
rect 2055 1773 2059 1774
rect 2135 1778 2139 1779
rect 2135 1773 2139 1774
rect 2175 1778 2179 1779
rect 2175 1773 2179 1774
rect 1694 1772 1700 1773
rect 1694 1768 1695 1772
rect 1699 1768 1700 1772
rect 1694 1767 1700 1768
rect 1790 1772 1796 1773
rect 1790 1768 1791 1772
rect 1795 1768 1796 1772
rect 1790 1767 1796 1768
rect 1878 1772 1884 1773
rect 1878 1768 1879 1772
rect 1883 1768 1884 1772
rect 1878 1767 1884 1768
rect 1966 1772 1972 1773
rect 1966 1768 1967 1772
rect 1971 1768 1972 1772
rect 1966 1767 1972 1768
rect 2054 1772 2060 1773
rect 2054 1768 2055 1772
rect 2059 1768 2060 1772
rect 2054 1767 2060 1768
rect 2134 1772 2140 1773
rect 2134 1768 2135 1772
rect 2139 1768 2140 1772
rect 2134 1767 2140 1768
rect 1286 1755 1292 1756
rect 1655 1756 1659 1757
rect 1174 1739 1180 1740
rect 1174 1735 1175 1739
rect 1179 1735 1180 1739
rect 1174 1734 1180 1735
rect 1288 1731 1290 1755
rect 1326 1752 1332 1753
rect 1915 1756 1919 1757
rect 1326 1748 1327 1752
rect 1331 1748 1332 1752
rect 1326 1747 1332 1748
rect 1542 1751 1548 1752
rect 1542 1747 1543 1751
rect 1547 1747 1548 1751
rect 1047 1730 1051 1731
rect 1047 1725 1051 1726
rect 1079 1730 1083 1731
rect 1079 1725 1083 1726
rect 1159 1730 1163 1731
rect 1159 1725 1163 1726
rect 1167 1730 1171 1731
rect 1167 1725 1171 1726
rect 1287 1730 1291 1731
rect 1287 1725 1291 1726
rect 1026 1723 1032 1724
rect 1026 1719 1027 1723
rect 1031 1719 1032 1723
rect 1026 1718 1032 1719
rect 1048 1706 1050 1725
rect 1070 1723 1076 1724
rect 1070 1719 1071 1723
rect 1075 1719 1076 1723
rect 1070 1718 1076 1719
rect 1046 1705 1052 1706
rect 934 1700 940 1701
rect 954 1703 960 1704
rect 954 1699 955 1703
rect 959 1699 960 1703
rect 1046 1701 1047 1705
rect 1051 1701 1052 1705
rect 1072 1704 1074 1718
rect 1160 1706 1162 1725
rect 1158 1705 1164 1706
rect 1288 1705 1290 1725
rect 1328 1723 1330 1747
rect 1542 1746 1548 1747
rect 1602 1751 1608 1752
rect 1602 1747 1603 1751
rect 1607 1747 1608 1751
rect 1602 1746 1608 1747
rect 1622 1751 1628 1752
rect 1655 1751 1659 1752
rect 1690 1751 1696 1752
rect 1622 1747 1623 1751
rect 1627 1747 1628 1751
rect 1622 1746 1628 1747
rect 1690 1747 1691 1751
rect 1695 1747 1696 1751
rect 1690 1746 1696 1747
rect 1710 1751 1716 1752
rect 1710 1747 1711 1751
rect 1715 1747 1716 1751
rect 1710 1746 1716 1747
rect 1786 1751 1792 1752
rect 1786 1747 1787 1751
rect 1791 1747 1792 1751
rect 1786 1746 1792 1747
rect 1806 1751 1812 1752
rect 1806 1747 1807 1751
rect 1811 1747 1812 1751
rect 1806 1746 1812 1747
rect 1874 1751 1880 1752
rect 1874 1747 1875 1751
rect 1879 1747 1880 1751
rect 1874 1746 1880 1747
rect 1894 1751 1900 1752
rect 1894 1747 1895 1751
rect 1899 1747 1900 1751
rect 1894 1746 1900 1747
rect 1914 1751 1920 1752
rect 1914 1747 1915 1751
rect 1919 1747 1920 1751
rect 1914 1746 1920 1747
rect 1982 1751 1988 1752
rect 1982 1747 1983 1751
rect 1987 1747 1988 1751
rect 1982 1746 1988 1747
rect 2050 1751 2056 1752
rect 2050 1747 2051 1751
rect 2055 1747 2056 1751
rect 2050 1746 2056 1747
rect 2070 1751 2076 1752
rect 2070 1747 2071 1751
rect 2075 1747 2076 1751
rect 2070 1746 2076 1747
rect 2090 1751 2096 1752
rect 2090 1747 2091 1751
rect 2095 1747 2096 1751
rect 2090 1746 2096 1747
rect 2150 1751 2156 1752
rect 2150 1747 2151 1751
rect 2155 1747 2156 1751
rect 2150 1746 2156 1747
rect 1544 1723 1546 1746
rect 1604 1732 1606 1746
rect 1594 1731 1600 1732
rect 1594 1727 1595 1731
rect 1599 1727 1600 1731
rect 1594 1726 1600 1727
rect 1602 1731 1608 1732
rect 1602 1727 1603 1731
rect 1607 1727 1608 1731
rect 1602 1726 1608 1727
rect 1327 1722 1331 1723
rect 1327 1717 1331 1718
rect 1399 1722 1403 1723
rect 1399 1717 1403 1718
rect 1463 1722 1467 1723
rect 1463 1717 1467 1718
rect 1543 1722 1547 1723
rect 1543 1717 1547 1718
rect 1046 1700 1052 1701
rect 1070 1703 1076 1704
rect 954 1698 960 1699
rect 1070 1699 1071 1703
rect 1075 1699 1076 1703
rect 1158 1701 1159 1705
rect 1163 1701 1164 1705
rect 1286 1704 1292 1705
rect 1158 1700 1164 1701
rect 1174 1703 1180 1704
rect 1070 1698 1076 1699
rect 1174 1699 1175 1703
rect 1179 1699 1180 1703
rect 1286 1700 1287 1704
rect 1291 1700 1292 1704
rect 1286 1699 1292 1700
rect 1174 1698 1180 1699
rect 918 1684 924 1685
rect 918 1680 919 1684
rect 923 1680 924 1684
rect 918 1679 924 1680
rect 1030 1684 1036 1685
rect 1030 1680 1031 1684
rect 1035 1680 1036 1684
rect 1030 1679 1036 1680
rect 1142 1684 1148 1685
rect 1142 1680 1143 1684
rect 1147 1680 1148 1684
rect 1142 1679 1148 1680
rect 920 1675 922 1679
rect 1032 1675 1034 1679
rect 1144 1675 1146 1679
rect 919 1674 923 1675
rect 919 1669 923 1670
rect 959 1674 963 1675
rect 959 1669 963 1670
rect 1031 1674 1035 1675
rect 1031 1669 1035 1670
rect 1063 1674 1067 1675
rect 1063 1669 1067 1670
rect 1143 1674 1147 1675
rect 1143 1669 1147 1670
rect 1167 1674 1171 1675
rect 1167 1669 1171 1670
rect 958 1668 964 1669
rect 958 1664 959 1668
rect 963 1664 964 1668
rect 958 1663 964 1664
rect 1062 1668 1068 1669
rect 1062 1664 1063 1668
rect 1067 1664 1068 1668
rect 1062 1663 1068 1664
rect 1166 1668 1172 1669
rect 1166 1664 1167 1668
rect 1171 1664 1172 1668
rect 1166 1663 1172 1664
rect 686 1647 692 1648
rect 686 1643 687 1647
rect 691 1643 692 1647
rect 686 1642 692 1643
rect 762 1647 768 1648
rect 762 1643 763 1647
rect 767 1643 768 1647
rect 762 1642 768 1643
rect 782 1647 788 1648
rect 782 1643 783 1647
rect 787 1643 788 1647
rect 782 1642 788 1643
rect 798 1647 804 1648
rect 798 1643 799 1647
rect 803 1643 804 1647
rect 798 1642 804 1643
rect 878 1647 884 1648
rect 878 1643 879 1647
rect 883 1643 884 1647
rect 878 1642 884 1643
rect 910 1647 916 1648
rect 910 1643 911 1647
rect 915 1643 916 1647
rect 910 1642 916 1643
rect 974 1647 980 1648
rect 974 1643 975 1647
rect 979 1643 980 1647
rect 974 1642 980 1643
rect 1058 1647 1064 1648
rect 1058 1643 1059 1647
rect 1063 1643 1064 1647
rect 1058 1642 1064 1643
rect 1078 1647 1084 1648
rect 1078 1643 1079 1647
rect 1083 1643 1084 1647
rect 1078 1642 1084 1643
rect 1098 1647 1104 1648
rect 1098 1643 1099 1647
rect 1103 1643 1104 1647
rect 1098 1642 1104 1643
rect 614 1627 620 1628
rect 614 1623 615 1627
rect 619 1623 620 1627
rect 614 1622 620 1623
rect 688 1619 690 1642
rect 764 1628 766 1642
rect 754 1627 760 1628
rect 754 1623 755 1627
rect 759 1623 760 1627
rect 754 1622 760 1623
rect 762 1627 768 1628
rect 762 1623 763 1627
rect 767 1623 768 1627
rect 762 1622 768 1623
rect 687 1618 691 1619
rect 687 1613 691 1614
rect 695 1618 699 1619
rect 695 1613 699 1614
rect 606 1611 612 1612
rect 606 1607 607 1611
rect 611 1607 612 1611
rect 606 1606 612 1607
rect 696 1594 698 1613
rect 706 1611 712 1612
rect 706 1607 707 1611
rect 711 1607 712 1611
rect 706 1606 712 1607
rect 718 1611 724 1612
rect 718 1607 719 1611
rect 723 1607 724 1611
rect 718 1606 724 1607
rect 430 1593 436 1594
rect 358 1588 364 1589
rect 382 1591 388 1592
rect 326 1586 332 1587
rect 382 1587 383 1591
rect 387 1587 388 1591
rect 430 1589 431 1593
rect 435 1589 436 1593
rect 510 1593 516 1594
rect 430 1588 436 1589
rect 478 1591 484 1592
rect 382 1586 388 1587
rect 478 1587 479 1591
rect 483 1587 484 1591
rect 478 1586 484 1587
rect 502 1591 508 1592
rect 502 1587 503 1591
rect 507 1587 508 1591
rect 510 1589 511 1593
rect 515 1589 516 1593
rect 598 1593 604 1594
rect 510 1588 516 1589
rect 518 1591 524 1592
rect 502 1586 508 1587
rect 518 1587 519 1591
rect 523 1587 524 1591
rect 598 1589 599 1593
rect 603 1589 604 1593
rect 598 1588 604 1589
rect 694 1593 700 1594
rect 694 1589 695 1593
rect 699 1589 700 1593
rect 694 1588 700 1589
rect 518 1586 524 1587
rect 286 1572 292 1573
rect 286 1568 287 1572
rect 291 1568 292 1572
rect 286 1567 292 1568
rect 342 1572 348 1573
rect 342 1568 343 1572
rect 347 1568 348 1572
rect 342 1567 348 1568
rect 414 1572 420 1573
rect 414 1568 415 1572
rect 419 1568 420 1572
rect 414 1567 420 1568
rect 287 1566 291 1567
rect 287 1561 291 1562
rect 319 1566 323 1567
rect 319 1561 323 1562
rect 343 1566 347 1567
rect 343 1561 347 1562
rect 399 1566 403 1567
rect 399 1561 403 1562
rect 415 1566 419 1567
rect 415 1561 419 1562
rect 318 1560 324 1561
rect 318 1556 319 1560
rect 323 1556 324 1560
rect 318 1555 324 1556
rect 398 1560 404 1561
rect 398 1556 399 1560
rect 403 1556 404 1560
rect 398 1555 404 1556
rect 262 1539 268 1540
rect 262 1535 263 1539
rect 267 1535 268 1539
rect 262 1534 268 1535
rect 270 1539 276 1540
rect 270 1535 271 1539
rect 275 1535 276 1539
rect 270 1534 276 1535
rect 334 1539 340 1540
rect 334 1535 335 1539
rect 339 1535 340 1539
rect 334 1534 340 1535
rect 350 1539 356 1540
rect 350 1535 351 1539
rect 355 1535 356 1539
rect 350 1534 356 1535
rect 414 1539 420 1540
rect 414 1535 415 1539
rect 419 1535 420 1539
rect 414 1534 420 1535
rect 254 1519 260 1520
rect 254 1515 255 1519
rect 259 1515 260 1519
rect 254 1514 260 1515
rect 264 1507 266 1534
rect 111 1506 115 1507
rect 111 1501 115 1502
rect 263 1506 267 1507
rect 263 1501 267 1502
rect 112 1481 114 1501
rect 272 1500 274 1534
rect 336 1507 338 1534
rect 279 1506 283 1507
rect 279 1501 283 1502
rect 335 1506 339 1507
rect 335 1501 339 1502
rect 343 1506 347 1507
rect 343 1501 347 1502
rect 270 1499 276 1500
rect 270 1495 271 1499
rect 275 1495 276 1499
rect 270 1494 276 1495
rect 280 1482 282 1501
rect 344 1482 346 1501
rect 352 1500 354 1534
rect 416 1507 418 1534
rect 480 1520 482 1586
rect 504 1579 506 1586
rect 520 1579 522 1586
rect 504 1577 522 1579
rect 494 1572 500 1573
rect 494 1568 495 1572
rect 499 1568 500 1572
rect 494 1567 500 1568
rect 582 1572 588 1573
rect 582 1568 583 1572
rect 587 1568 588 1572
rect 582 1567 588 1568
rect 678 1572 684 1573
rect 678 1568 679 1572
rect 683 1568 684 1572
rect 678 1567 684 1568
rect 487 1566 491 1567
rect 487 1561 491 1562
rect 495 1566 499 1567
rect 495 1561 499 1562
rect 583 1566 587 1567
rect 583 1561 587 1562
rect 671 1566 675 1567
rect 671 1561 675 1562
rect 679 1566 683 1567
rect 679 1561 683 1562
rect 486 1560 492 1561
rect 486 1556 487 1560
rect 491 1556 492 1560
rect 486 1555 492 1556
rect 582 1560 588 1561
rect 582 1556 583 1560
rect 587 1556 588 1560
rect 582 1555 588 1556
rect 670 1560 676 1561
rect 670 1556 671 1560
rect 675 1556 676 1560
rect 670 1555 676 1556
rect 708 1540 710 1606
rect 720 1592 722 1606
rect 756 1600 758 1622
rect 784 1619 786 1642
rect 880 1619 882 1642
rect 914 1627 920 1628
rect 914 1623 915 1627
rect 919 1623 920 1627
rect 914 1622 920 1623
rect 783 1618 787 1619
rect 783 1613 787 1614
rect 791 1618 795 1619
rect 791 1613 795 1614
rect 879 1618 883 1619
rect 879 1613 883 1614
rect 895 1618 899 1619
rect 895 1613 899 1614
rect 754 1599 760 1600
rect 754 1595 755 1599
rect 759 1595 760 1599
rect 754 1594 760 1595
rect 792 1594 794 1613
rect 798 1611 804 1612
rect 798 1607 799 1611
rect 803 1607 804 1611
rect 798 1606 804 1607
rect 790 1593 796 1594
rect 718 1591 724 1592
rect 718 1587 719 1591
rect 723 1587 724 1591
rect 790 1589 791 1593
rect 795 1589 796 1593
rect 790 1588 796 1589
rect 718 1586 724 1587
rect 774 1572 780 1573
rect 774 1568 775 1572
rect 779 1568 780 1572
rect 774 1567 780 1568
rect 759 1566 763 1567
rect 759 1561 763 1562
rect 775 1566 779 1567
rect 775 1561 779 1562
rect 758 1560 764 1561
rect 758 1556 759 1560
rect 763 1556 764 1560
rect 758 1555 764 1556
rect 800 1540 802 1606
rect 896 1594 898 1613
rect 894 1593 900 1594
rect 894 1589 895 1593
rect 899 1589 900 1593
rect 916 1592 918 1622
rect 976 1619 978 1642
rect 1060 1628 1062 1642
rect 1058 1627 1064 1628
rect 1058 1623 1059 1627
rect 1063 1623 1064 1627
rect 1058 1622 1064 1623
rect 1080 1619 1082 1642
rect 975 1618 979 1619
rect 975 1613 979 1614
rect 1007 1618 1011 1619
rect 1007 1613 1011 1614
rect 1079 1618 1083 1619
rect 1079 1613 1083 1614
rect 1008 1594 1010 1613
rect 1100 1612 1102 1642
rect 1176 1628 1178 1698
rect 1328 1697 1330 1717
rect 1400 1698 1402 1717
rect 1414 1715 1420 1716
rect 1414 1711 1415 1715
rect 1419 1711 1420 1715
rect 1414 1710 1420 1711
rect 1422 1715 1428 1716
rect 1422 1711 1423 1715
rect 1427 1711 1428 1715
rect 1422 1710 1428 1711
rect 1398 1697 1404 1698
rect 1326 1696 1332 1697
rect 1326 1692 1327 1696
rect 1331 1692 1332 1696
rect 1398 1693 1399 1697
rect 1403 1693 1404 1697
rect 1398 1692 1404 1693
rect 1326 1691 1332 1692
rect 1286 1687 1292 1688
rect 1286 1683 1287 1687
rect 1291 1683 1292 1687
rect 1286 1682 1292 1683
rect 1288 1675 1290 1682
rect 1326 1679 1332 1680
rect 1326 1675 1327 1679
rect 1331 1675 1332 1679
rect 1287 1674 1291 1675
rect 1326 1674 1332 1675
rect 1382 1676 1388 1677
rect 1287 1669 1291 1670
rect 1288 1666 1290 1669
rect 1328 1667 1330 1674
rect 1382 1672 1383 1676
rect 1387 1672 1388 1676
rect 1382 1671 1388 1672
rect 1384 1667 1386 1671
rect 1327 1666 1331 1667
rect 1286 1665 1292 1666
rect 1286 1661 1287 1665
rect 1291 1661 1292 1665
rect 1327 1661 1331 1662
rect 1351 1666 1355 1667
rect 1351 1661 1355 1662
rect 1383 1666 1387 1667
rect 1383 1661 1387 1662
rect 1407 1666 1411 1667
rect 1407 1661 1411 1662
rect 1286 1660 1292 1661
rect 1328 1658 1330 1661
rect 1350 1660 1356 1661
rect 1326 1657 1332 1658
rect 1326 1653 1327 1657
rect 1331 1653 1332 1657
rect 1350 1656 1351 1660
rect 1355 1656 1356 1660
rect 1350 1655 1356 1656
rect 1406 1660 1412 1661
rect 1406 1656 1407 1660
rect 1411 1656 1412 1660
rect 1406 1655 1412 1656
rect 1326 1652 1332 1653
rect 1286 1648 1292 1649
rect 1182 1647 1188 1648
rect 1182 1643 1183 1647
rect 1187 1643 1188 1647
rect 1286 1644 1287 1648
rect 1291 1644 1292 1648
rect 1416 1645 1418 1710
rect 1424 1696 1426 1710
rect 1464 1698 1466 1717
rect 1486 1715 1492 1716
rect 1486 1711 1487 1715
rect 1491 1711 1492 1715
rect 1486 1710 1492 1711
rect 1462 1697 1468 1698
rect 1422 1695 1428 1696
rect 1422 1691 1423 1695
rect 1427 1691 1428 1695
rect 1462 1693 1463 1697
rect 1467 1693 1468 1697
rect 1488 1696 1490 1710
rect 1544 1698 1546 1717
rect 1566 1715 1572 1716
rect 1566 1711 1567 1715
rect 1571 1711 1572 1715
rect 1566 1710 1572 1711
rect 1542 1697 1548 1698
rect 1462 1692 1468 1693
rect 1486 1695 1492 1696
rect 1422 1690 1428 1691
rect 1486 1691 1487 1695
rect 1491 1691 1492 1695
rect 1542 1693 1543 1697
rect 1547 1693 1548 1697
rect 1568 1696 1570 1710
rect 1596 1701 1598 1726
rect 1624 1723 1626 1746
rect 1692 1732 1694 1746
rect 1690 1731 1696 1732
rect 1690 1727 1691 1731
rect 1695 1727 1696 1731
rect 1690 1726 1696 1727
rect 1712 1723 1714 1746
rect 1788 1732 1790 1746
rect 1786 1731 1792 1732
rect 1786 1727 1787 1731
rect 1791 1727 1792 1731
rect 1786 1726 1792 1727
rect 1808 1723 1810 1746
rect 1876 1732 1878 1746
rect 1874 1731 1880 1732
rect 1874 1727 1875 1731
rect 1879 1727 1880 1731
rect 1874 1726 1880 1727
rect 1896 1723 1898 1746
rect 1984 1723 1986 1746
rect 2052 1732 2054 1746
rect 2050 1731 2056 1732
rect 2050 1727 2051 1731
rect 2055 1727 2056 1731
rect 2050 1726 2056 1727
rect 2072 1723 2074 1746
rect 1623 1722 1627 1723
rect 1623 1717 1627 1718
rect 1631 1722 1635 1723
rect 1631 1717 1635 1718
rect 1711 1722 1715 1723
rect 1711 1717 1715 1718
rect 1727 1722 1731 1723
rect 1727 1717 1731 1718
rect 1807 1722 1811 1723
rect 1807 1717 1811 1718
rect 1823 1722 1827 1723
rect 1823 1717 1827 1718
rect 1895 1722 1899 1723
rect 1895 1717 1899 1718
rect 1919 1722 1923 1723
rect 1919 1717 1923 1718
rect 1983 1722 1987 1723
rect 1983 1717 1987 1718
rect 2015 1722 2019 1723
rect 2015 1717 2019 1718
rect 2071 1722 2075 1723
rect 2071 1717 2075 1718
rect 1595 1700 1599 1701
rect 1632 1698 1634 1717
rect 1654 1715 1660 1716
rect 1654 1711 1655 1715
rect 1659 1711 1660 1715
rect 1654 1710 1660 1711
rect 1542 1692 1548 1693
rect 1566 1695 1572 1696
rect 1595 1695 1599 1696
rect 1630 1697 1636 1698
rect 1486 1690 1492 1691
rect 1566 1691 1567 1695
rect 1571 1691 1572 1695
rect 1630 1693 1631 1697
rect 1635 1693 1636 1697
rect 1656 1696 1658 1710
rect 1728 1698 1730 1717
rect 1750 1715 1756 1716
rect 1750 1711 1751 1715
rect 1755 1711 1756 1715
rect 1750 1710 1756 1711
rect 1726 1697 1732 1698
rect 1630 1692 1636 1693
rect 1654 1695 1660 1696
rect 1566 1690 1572 1691
rect 1654 1691 1655 1695
rect 1659 1691 1660 1695
rect 1726 1693 1727 1697
rect 1731 1693 1732 1697
rect 1752 1696 1754 1710
rect 1824 1698 1826 1717
rect 1843 1700 1847 1701
rect 1822 1697 1828 1698
rect 1726 1692 1732 1693
rect 1750 1695 1756 1696
rect 1654 1690 1660 1691
rect 1750 1691 1751 1695
rect 1755 1691 1756 1695
rect 1822 1693 1823 1697
rect 1827 1693 1828 1697
rect 1920 1698 1922 1717
rect 1942 1715 1948 1716
rect 1942 1711 1943 1715
rect 1947 1711 1948 1715
rect 1942 1710 1948 1711
rect 1918 1697 1924 1698
rect 1822 1692 1828 1693
rect 1842 1695 1848 1696
rect 1750 1690 1756 1691
rect 1842 1691 1843 1695
rect 1847 1691 1848 1695
rect 1918 1693 1919 1697
rect 1923 1693 1924 1697
rect 1944 1696 1946 1710
rect 2016 1698 2018 1717
rect 2092 1716 2094 1746
rect 2152 1723 2154 1746
rect 2208 1732 2210 1798
rect 2318 1784 2324 1785
rect 2318 1780 2319 1784
rect 2323 1780 2324 1784
rect 2318 1779 2324 1780
rect 2215 1778 2219 1779
rect 2215 1773 2219 1774
rect 2295 1778 2299 1779
rect 2295 1773 2299 1774
rect 2319 1778 2323 1779
rect 2319 1773 2323 1774
rect 2214 1772 2220 1773
rect 2214 1768 2215 1772
rect 2219 1768 2220 1772
rect 2214 1767 2220 1768
rect 2294 1772 2300 1773
rect 2294 1768 2295 1772
rect 2299 1768 2300 1772
rect 2294 1767 2300 1768
rect 2328 1752 2330 1818
rect 2336 1806 2338 1825
rect 2456 1806 2458 1825
rect 2464 1824 2466 1854
rect 2472 1840 2474 1910
rect 2502 1899 2508 1900
rect 2502 1895 2503 1899
rect 2507 1895 2508 1899
rect 2502 1894 2508 1895
rect 2504 1887 2506 1894
rect 2503 1886 2507 1887
rect 2503 1881 2507 1882
rect 2504 1878 2506 1881
rect 2502 1877 2508 1878
rect 2502 1873 2503 1877
rect 2507 1873 2508 1877
rect 2502 1872 2508 1873
rect 2502 1860 2508 1861
rect 2502 1856 2503 1860
rect 2507 1856 2508 1860
rect 2502 1855 2508 1856
rect 2470 1839 2476 1840
rect 2470 1835 2471 1839
rect 2475 1835 2476 1839
rect 2470 1834 2476 1835
rect 2504 1831 2506 1855
rect 2503 1830 2507 1831
rect 2503 1825 2507 1826
rect 2462 1823 2468 1824
rect 2462 1819 2463 1823
rect 2467 1819 2468 1823
rect 2462 1818 2468 1819
rect 2334 1805 2340 1806
rect 2334 1801 2335 1805
rect 2339 1801 2340 1805
rect 2334 1800 2340 1801
rect 2454 1805 2460 1806
rect 2504 1805 2506 1825
rect 2454 1801 2455 1805
rect 2459 1801 2460 1805
rect 2502 1804 2508 1805
rect 2454 1800 2460 1801
rect 2470 1803 2476 1804
rect 2470 1799 2471 1803
rect 2475 1799 2476 1803
rect 2502 1800 2503 1804
rect 2507 1800 2508 1804
rect 2502 1799 2508 1800
rect 2470 1798 2476 1799
rect 2438 1784 2444 1785
rect 2438 1780 2439 1784
rect 2443 1780 2444 1784
rect 2438 1779 2444 1780
rect 2375 1778 2379 1779
rect 2375 1773 2379 1774
rect 2439 1778 2443 1779
rect 2439 1773 2443 1774
rect 2374 1772 2380 1773
rect 2374 1768 2375 1772
rect 2379 1768 2380 1772
rect 2374 1767 2380 1768
rect 2438 1772 2444 1773
rect 2438 1768 2439 1772
rect 2443 1768 2444 1772
rect 2438 1767 2444 1768
rect 2230 1751 2236 1752
rect 2230 1747 2231 1751
rect 2235 1747 2236 1751
rect 2230 1746 2236 1747
rect 2310 1751 2316 1752
rect 2310 1747 2311 1751
rect 2315 1747 2316 1751
rect 2310 1746 2316 1747
rect 2326 1751 2332 1752
rect 2326 1747 2327 1751
rect 2331 1747 2332 1751
rect 2326 1746 2332 1747
rect 2390 1751 2396 1752
rect 2390 1747 2391 1751
rect 2395 1747 2396 1751
rect 2390 1746 2396 1747
rect 2454 1751 2460 1752
rect 2454 1747 2455 1751
rect 2459 1747 2460 1751
rect 2454 1746 2460 1747
rect 2462 1751 2468 1752
rect 2462 1747 2463 1751
rect 2467 1747 2468 1751
rect 2462 1746 2468 1747
rect 2206 1731 2212 1732
rect 2206 1727 2207 1731
rect 2211 1727 2212 1731
rect 2206 1726 2212 1727
rect 2232 1723 2234 1746
rect 2312 1723 2314 1746
rect 2392 1723 2394 1746
rect 2402 1731 2408 1732
rect 2402 1727 2403 1731
rect 2407 1727 2408 1731
rect 2402 1726 2408 1727
rect 2111 1722 2115 1723
rect 2111 1717 2115 1718
rect 2151 1722 2155 1723
rect 2151 1717 2155 1718
rect 2199 1722 2203 1723
rect 2199 1717 2203 1718
rect 2231 1722 2235 1723
rect 2231 1717 2235 1718
rect 2287 1722 2291 1723
rect 2287 1717 2291 1718
rect 2311 1722 2315 1723
rect 2311 1717 2315 1718
rect 2383 1722 2387 1723
rect 2383 1717 2387 1718
rect 2391 1722 2395 1723
rect 2391 1717 2395 1718
rect 2090 1715 2096 1716
rect 2090 1711 2091 1715
rect 2095 1711 2096 1715
rect 2090 1710 2096 1711
rect 2112 1698 2114 1717
rect 2134 1715 2140 1716
rect 2134 1711 2135 1715
rect 2139 1711 2140 1715
rect 2134 1710 2140 1711
rect 2014 1697 2020 1698
rect 1918 1692 1924 1693
rect 1942 1695 1948 1696
rect 1842 1690 1848 1691
rect 1942 1691 1943 1695
rect 1947 1691 1948 1695
rect 2014 1693 2015 1697
rect 2019 1693 2020 1697
rect 2110 1697 2116 1698
rect 2014 1692 2020 1693
rect 2030 1695 2036 1696
rect 1942 1690 1948 1691
rect 2030 1691 2031 1695
rect 2035 1691 2036 1695
rect 2110 1693 2111 1697
rect 2115 1693 2116 1697
rect 2136 1696 2138 1710
rect 2200 1698 2202 1717
rect 2288 1698 2290 1717
rect 2318 1715 2324 1716
rect 2318 1711 2319 1715
rect 2323 1711 2324 1715
rect 2318 1710 2324 1711
rect 2198 1697 2204 1698
rect 2110 1692 2116 1693
rect 2134 1695 2140 1696
rect 2030 1690 2036 1691
rect 2134 1691 2135 1695
rect 2139 1691 2140 1695
rect 2198 1693 2199 1697
rect 2203 1693 2204 1697
rect 2198 1692 2204 1693
rect 2286 1697 2292 1698
rect 2286 1693 2287 1697
rect 2291 1693 2292 1697
rect 2320 1696 2322 1710
rect 2384 1698 2386 1717
rect 2382 1697 2388 1698
rect 2286 1692 2292 1693
rect 2318 1695 2324 1696
rect 2134 1690 2140 1691
rect 2318 1691 2319 1695
rect 2323 1691 2324 1695
rect 2382 1693 2383 1697
rect 2387 1693 2388 1697
rect 2404 1696 2406 1726
rect 2456 1723 2458 1746
rect 2455 1722 2459 1723
rect 2455 1717 2459 1718
rect 2456 1698 2458 1717
rect 2464 1716 2466 1746
rect 2472 1732 2474 1798
rect 2502 1787 2508 1788
rect 2502 1783 2503 1787
rect 2507 1783 2508 1787
rect 2502 1782 2508 1783
rect 2504 1779 2506 1782
rect 2503 1778 2507 1779
rect 2503 1773 2507 1774
rect 2504 1770 2506 1773
rect 2502 1769 2508 1770
rect 2502 1765 2503 1769
rect 2507 1765 2508 1769
rect 2502 1764 2508 1765
rect 2502 1752 2508 1753
rect 2502 1748 2503 1752
rect 2507 1748 2508 1752
rect 2502 1747 2508 1748
rect 2470 1731 2476 1732
rect 2470 1727 2471 1731
rect 2475 1727 2476 1731
rect 2470 1726 2476 1727
rect 2504 1723 2506 1747
rect 2503 1722 2507 1723
rect 2503 1717 2507 1718
rect 2462 1715 2468 1716
rect 2462 1711 2463 1715
rect 2467 1711 2468 1715
rect 2462 1710 2468 1711
rect 2474 1707 2480 1708
rect 2474 1703 2475 1707
rect 2479 1703 2480 1707
rect 2474 1702 2480 1703
rect 2454 1697 2460 1698
rect 2382 1692 2388 1693
rect 2402 1695 2408 1696
rect 2318 1690 2324 1691
rect 2402 1691 2403 1695
rect 2407 1691 2408 1695
rect 2454 1693 2455 1697
rect 2459 1693 2460 1697
rect 2454 1692 2460 1693
rect 2462 1695 2468 1696
rect 2402 1690 2408 1691
rect 2462 1691 2463 1695
rect 2467 1691 2468 1695
rect 2462 1690 2468 1691
rect 1446 1676 1452 1677
rect 1446 1672 1447 1676
rect 1451 1672 1452 1676
rect 1446 1671 1452 1672
rect 1526 1676 1532 1677
rect 1526 1672 1527 1676
rect 1531 1672 1532 1676
rect 1526 1671 1532 1672
rect 1614 1676 1620 1677
rect 1614 1672 1615 1676
rect 1619 1672 1620 1676
rect 1614 1671 1620 1672
rect 1710 1676 1716 1677
rect 1710 1672 1711 1676
rect 1715 1672 1716 1676
rect 1710 1671 1716 1672
rect 1806 1676 1812 1677
rect 1806 1672 1807 1676
rect 1811 1672 1812 1676
rect 1806 1671 1812 1672
rect 1902 1676 1908 1677
rect 1902 1672 1903 1676
rect 1907 1672 1908 1676
rect 1902 1671 1908 1672
rect 1998 1676 2004 1677
rect 1998 1672 1999 1676
rect 2003 1672 2004 1676
rect 1998 1671 2004 1672
rect 1448 1667 1450 1671
rect 1528 1667 1530 1671
rect 1616 1667 1618 1671
rect 1712 1667 1714 1671
rect 1808 1667 1810 1671
rect 1904 1667 1906 1671
rect 2000 1667 2002 1671
rect 1447 1666 1451 1667
rect 1447 1661 1451 1662
rect 1495 1666 1499 1667
rect 1495 1661 1499 1662
rect 1527 1666 1531 1667
rect 1527 1661 1531 1662
rect 1583 1666 1587 1667
rect 1583 1661 1587 1662
rect 1615 1666 1619 1667
rect 1615 1661 1619 1662
rect 1679 1666 1683 1667
rect 1679 1661 1683 1662
rect 1711 1666 1715 1667
rect 1711 1661 1715 1662
rect 1783 1666 1787 1667
rect 1783 1661 1787 1662
rect 1807 1666 1811 1667
rect 1807 1661 1811 1662
rect 1895 1666 1899 1667
rect 1895 1661 1899 1662
rect 1903 1666 1907 1667
rect 1903 1661 1907 1662
rect 1999 1666 2003 1667
rect 1999 1661 2003 1662
rect 2023 1666 2027 1667
rect 2023 1661 2027 1662
rect 1494 1660 1500 1661
rect 1494 1656 1495 1660
rect 1499 1656 1500 1660
rect 1494 1655 1500 1656
rect 1582 1660 1588 1661
rect 1582 1656 1583 1660
rect 1587 1656 1588 1660
rect 1582 1655 1588 1656
rect 1678 1660 1684 1661
rect 1678 1656 1679 1660
rect 1683 1656 1684 1660
rect 1678 1655 1684 1656
rect 1782 1660 1788 1661
rect 1782 1656 1783 1660
rect 1787 1656 1788 1660
rect 1782 1655 1788 1656
rect 1894 1660 1900 1661
rect 1894 1656 1895 1660
rect 1899 1656 1900 1660
rect 1894 1655 1900 1656
rect 2022 1660 2028 1661
rect 2022 1656 2023 1660
rect 2027 1656 2028 1660
rect 2022 1655 2028 1656
rect 1286 1643 1292 1644
rect 1415 1644 1419 1645
rect 1182 1642 1188 1643
rect 1174 1627 1180 1628
rect 1174 1623 1175 1627
rect 1179 1623 1180 1627
rect 1174 1622 1180 1623
rect 1184 1619 1186 1642
rect 1288 1619 1290 1643
rect 1326 1640 1332 1641
rect 1703 1644 1707 1645
rect 1326 1636 1327 1640
rect 1331 1636 1332 1640
rect 1326 1635 1332 1636
rect 1366 1639 1372 1640
rect 1366 1635 1367 1639
rect 1371 1635 1372 1639
rect 1119 1618 1123 1619
rect 1119 1613 1123 1614
rect 1183 1618 1187 1619
rect 1183 1613 1187 1614
rect 1287 1618 1291 1619
rect 1328 1615 1330 1635
rect 1366 1634 1372 1635
rect 1402 1639 1408 1640
rect 1415 1639 1419 1640
rect 1422 1639 1428 1640
rect 1402 1635 1403 1639
rect 1407 1635 1408 1639
rect 1402 1634 1408 1635
rect 1422 1635 1423 1639
rect 1427 1635 1428 1639
rect 1422 1634 1428 1635
rect 1490 1639 1496 1640
rect 1490 1635 1491 1639
rect 1495 1635 1496 1639
rect 1490 1634 1496 1635
rect 1510 1639 1516 1640
rect 1510 1635 1511 1639
rect 1515 1635 1516 1639
rect 1510 1634 1516 1635
rect 1578 1639 1584 1640
rect 1578 1635 1579 1639
rect 1583 1635 1584 1639
rect 1578 1634 1584 1635
rect 1598 1639 1604 1640
rect 1598 1635 1599 1639
rect 1603 1635 1604 1639
rect 1598 1634 1604 1635
rect 1674 1639 1680 1640
rect 1674 1635 1675 1639
rect 1679 1635 1680 1639
rect 1674 1634 1680 1635
rect 1694 1639 1700 1640
rect 1694 1635 1695 1639
rect 1699 1635 1700 1639
rect 1694 1634 1700 1635
rect 1702 1639 1708 1640
rect 1702 1635 1703 1639
rect 1707 1635 1708 1639
rect 1702 1634 1708 1635
rect 1798 1639 1804 1640
rect 1798 1635 1799 1639
rect 1803 1635 1804 1639
rect 1798 1634 1804 1635
rect 1890 1639 1896 1640
rect 1890 1635 1891 1639
rect 1895 1635 1896 1639
rect 1890 1634 1896 1635
rect 1910 1639 1916 1640
rect 1910 1635 1911 1639
rect 1915 1635 1916 1639
rect 1910 1634 1916 1635
rect 1930 1639 1936 1640
rect 1930 1635 1931 1639
rect 1935 1635 1936 1639
rect 1930 1634 1936 1635
rect 1368 1615 1370 1634
rect 1404 1620 1406 1634
rect 1402 1619 1408 1620
rect 1402 1615 1403 1619
rect 1407 1615 1408 1619
rect 1424 1615 1426 1634
rect 1492 1620 1494 1634
rect 1490 1619 1496 1620
rect 1490 1615 1491 1619
rect 1495 1615 1496 1619
rect 1512 1615 1514 1634
rect 1580 1620 1582 1634
rect 1578 1619 1584 1620
rect 1578 1615 1579 1619
rect 1583 1615 1584 1619
rect 1600 1615 1602 1634
rect 1676 1620 1678 1634
rect 1674 1619 1680 1620
rect 1674 1615 1675 1619
rect 1679 1615 1680 1619
rect 1696 1615 1698 1634
rect 1800 1615 1802 1634
rect 1892 1620 1894 1634
rect 1890 1619 1896 1620
rect 1890 1615 1891 1619
rect 1895 1615 1896 1619
rect 1912 1615 1914 1634
rect 1287 1613 1291 1614
rect 1327 1614 1331 1615
rect 1098 1611 1104 1612
rect 1098 1607 1099 1611
rect 1103 1607 1104 1611
rect 1098 1606 1104 1607
rect 1120 1594 1122 1613
rect 1262 1607 1268 1608
rect 1262 1603 1263 1607
rect 1267 1603 1268 1607
rect 1262 1602 1268 1603
rect 1006 1593 1012 1594
rect 894 1588 900 1589
rect 914 1591 920 1592
rect 914 1587 915 1591
rect 919 1587 920 1591
rect 1006 1589 1007 1593
rect 1011 1589 1012 1593
rect 1118 1593 1124 1594
rect 1006 1588 1012 1589
rect 1014 1591 1020 1592
rect 914 1586 920 1587
rect 1014 1587 1015 1591
rect 1019 1587 1020 1591
rect 1118 1589 1119 1593
rect 1123 1589 1124 1593
rect 1118 1588 1124 1589
rect 1014 1586 1020 1587
rect 878 1572 884 1573
rect 878 1568 879 1572
rect 883 1568 884 1572
rect 878 1567 884 1568
rect 990 1572 996 1573
rect 990 1568 991 1572
rect 995 1568 996 1572
rect 990 1567 996 1568
rect 847 1566 851 1567
rect 847 1561 851 1562
rect 879 1566 883 1567
rect 879 1561 883 1562
rect 927 1566 931 1567
rect 927 1561 931 1562
rect 991 1566 995 1567
rect 991 1561 995 1562
rect 1007 1566 1011 1567
rect 1007 1561 1011 1562
rect 846 1560 852 1561
rect 846 1556 847 1560
rect 851 1556 852 1560
rect 846 1555 852 1556
rect 926 1560 932 1561
rect 926 1556 927 1560
rect 931 1556 932 1560
rect 926 1555 932 1556
rect 1006 1560 1012 1561
rect 1006 1556 1007 1560
rect 1011 1556 1012 1560
rect 1006 1555 1012 1556
rect 502 1539 508 1540
rect 502 1535 503 1539
rect 507 1535 508 1539
rect 502 1534 508 1535
rect 578 1539 584 1540
rect 578 1535 579 1539
rect 583 1535 584 1539
rect 578 1534 584 1535
rect 598 1539 604 1540
rect 598 1535 599 1539
rect 603 1535 604 1539
rect 598 1534 604 1535
rect 686 1539 692 1540
rect 686 1535 687 1539
rect 691 1535 692 1539
rect 686 1534 692 1535
rect 706 1539 712 1540
rect 706 1535 707 1539
rect 711 1535 712 1539
rect 706 1534 712 1535
rect 774 1539 780 1540
rect 774 1535 775 1539
rect 779 1535 780 1539
rect 774 1534 780 1535
rect 798 1539 804 1540
rect 798 1535 799 1539
rect 803 1535 804 1539
rect 798 1534 804 1535
rect 862 1539 868 1540
rect 862 1535 863 1539
rect 867 1535 868 1539
rect 862 1534 868 1535
rect 878 1539 884 1540
rect 878 1535 879 1539
rect 883 1535 884 1539
rect 878 1534 884 1535
rect 942 1539 948 1540
rect 942 1535 943 1539
rect 947 1535 948 1539
rect 942 1534 948 1535
rect 478 1519 484 1520
rect 478 1515 479 1519
rect 483 1515 484 1519
rect 478 1514 484 1515
rect 504 1507 506 1534
rect 580 1520 582 1534
rect 578 1519 584 1520
rect 578 1515 579 1519
rect 583 1515 584 1519
rect 578 1514 584 1515
rect 600 1507 602 1534
rect 670 1519 676 1520
rect 670 1515 671 1519
rect 675 1515 676 1519
rect 670 1514 676 1515
rect 415 1506 419 1507
rect 415 1501 419 1502
rect 495 1506 499 1507
rect 495 1501 499 1502
rect 503 1506 507 1507
rect 503 1501 507 1502
rect 575 1506 579 1507
rect 575 1501 579 1502
rect 599 1506 603 1507
rect 599 1501 603 1502
rect 655 1506 659 1507
rect 655 1501 659 1502
rect 350 1499 356 1500
rect 350 1495 351 1499
rect 355 1495 356 1499
rect 350 1494 356 1495
rect 366 1499 372 1500
rect 366 1495 367 1499
rect 371 1495 372 1499
rect 366 1494 372 1495
rect 278 1481 284 1482
rect 110 1480 116 1481
rect 110 1476 111 1480
rect 115 1476 116 1480
rect 278 1477 279 1481
rect 283 1477 284 1481
rect 342 1481 348 1482
rect 278 1476 284 1477
rect 286 1479 292 1480
rect 110 1475 116 1476
rect 286 1475 287 1479
rect 291 1475 292 1479
rect 342 1477 343 1481
rect 347 1477 348 1481
rect 368 1480 370 1494
rect 416 1482 418 1501
rect 438 1499 444 1500
rect 438 1495 439 1499
rect 443 1495 444 1499
rect 438 1494 444 1495
rect 414 1481 420 1482
rect 342 1476 348 1477
rect 366 1479 372 1480
rect 286 1474 292 1475
rect 366 1475 367 1479
rect 371 1475 372 1479
rect 414 1477 415 1481
rect 419 1477 420 1481
rect 440 1480 442 1494
rect 496 1482 498 1501
rect 576 1482 578 1501
rect 606 1499 612 1500
rect 606 1495 607 1499
rect 611 1495 612 1499
rect 606 1494 612 1495
rect 494 1481 500 1482
rect 414 1476 420 1477
rect 438 1479 444 1480
rect 366 1474 372 1475
rect 438 1475 439 1479
rect 443 1475 444 1479
rect 494 1477 495 1481
rect 499 1477 500 1481
rect 574 1481 580 1482
rect 494 1476 500 1477
rect 510 1479 516 1480
rect 438 1474 444 1475
rect 510 1475 511 1479
rect 515 1475 516 1479
rect 574 1477 575 1481
rect 579 1477 580 1481
rect 608 1480 610 1494
rect 630 1491 636 1492
rect 630 1487 631 1491
rect 635 1487 636 1491
rect 630 1486 636 1487
rect 574 1476 580 1477
rect 606 1479 612 1480
rect 510 1474 516 1475
rect 606 1475 607 1479
rect 611 1475 612 1479
rect 606 1474 612 1475
rect 110 1463 116 1464
rect 110 1459 111 1463
rect 115 1459 116 1463
rect 110 1458 116 1459
rect 262 1460 268 1461
rect 112 1451 114 1458
rect 262 1456 263 1460
rect 267 1456 268 1460
rect 262 1455 268 1456
rect 264 1451 266 1455
rect 111 1450 115 1451
rect 111 1445 115 1446
rect 191 1450 195 1451
rect 191 1445 195 1446
rect 255 1450 259 1451
rect 255 1445 259 1446
rect 263 1450 267 1451
rect 263 1445 267 1446
rect 112 1442 114 1445
rect 190 1444 196 1445
rect 110 1441 116 1442
rect 110 1437 111 1441
rect 115 1437 116 1441
rect 190 1440 191 1444
rect 195 1440 196 1444
rect 190 1439 196 1440
rect 254 1444 260 1445
rect 254 1440 255 1444
rect 259 1440 260 1444
rect 254 1439 260 1440
rect 110 1436 116 1437
rect 110 1424 116 1425
rect 110 1420 111 1424
rect 115 1420 116 1424
rect 110 1419 116 1420
rect 206 1423 212 1424
rect 206 1419 207 1423
rect 211 1419 212 1423
rect 112 1395 114 1419
rect 206 1418 212 1419
rect 214 1423 220 1424
rect 214 1419 215 1423
rect 219 1419 220 1423
rect 214 1418 220 1419
rect 270 1423 276 1424
rect 270 1419 271 1423
rect 275 1419 276 1423
rect 270 1418 276 1419
rect 208 1395 210 1418
rect 216 1396 218 1418
rect 214 1395 220 1396
rect 272 1395 274 1418
rect 288 1404 290 1474
rect 326 1460 332 1461
rect 326 1456 327 1460
rect 331 1456 332 1460
rect 326 1455 332 1456
rect 398 1460 404 1461
rect 398 1456 399 1460
rect 403 1456 404 1460
rect 398 1455 404 1456
rect 478 1460 484 1461
rect 478 1456 479 1460
rect 483 1456 484 1460
rect 478 1455 484 1456
rect 328 1451 330 1455
rect 400 1451 402 1455
rect 480 1451 482 1455
rect 327 1450 331 1451
rect 327 1445 331 1446
rect 399 1450 403 1451
rect 399 1445 403 1446
rect 407 1450 411 1451
rect 407 1445 411 1446
rect 479 1450 483 1451
rect 479 1445 483 1446
rect 503 1450 507 1451
rect 503 1445 507 1446
rect 326 1444 332 1445
rect 326 1440 327 1444
rect 331 1440 332 1444
rect 326 1439 332 1440
rect 406 1444 412 1445
rect 406 1440 407 1444
rect 411 1440 412 1444
rect 406 1439 412 1440
rect 502 1444 508 1445
rect 502 1440 503 1444
rect 507 1440 508 1444
rect 502 1439 508 1440
rect 342 1423 348 1424
rect 342 1419 343 1423
rect 347 1419 348 1423
rect 342 1418 348 1419
rect 350 1423 356 1424
rect 350 1419 351 1423
rect 355 1419 356 1423
rect 350 1418 356 1419
rect 422 1423 428 1424
rect 422 1419 423 1423
rect 427 1419 428 1423
rect 422 1418 428 1419
rect 286 1403 292 1404
rect 286 1399 287 1403
rect 291 1399 292 1403
rect 286 1398 292 1399
rect 344 1395 346 1418
rect 352 1396 354 1418
rect 350 1395 356 1396
rect 424 1395 426 1418
rect 512 1404 514 1474
rect 558 1460 564 1461
rect 558 1456 559 1460
rect 563 1456 564 1460
rect 558 1455 564 1456
rect 560 1451 562 1455
rect 559 1450 563 1451
rect 559 1445 563 1446
rect 607 1450 611 1451
rect 607 1445 611 1446
rect 606 1444 612 1445
rect 606 1440 607 1444
rect 611 1440 612 1444
rect 606 1439 612 1440
rect 632 1424 634 1486
rect 656 1482 658 1501
rect 654 1481 660 1482
rect 654 1477 655 1481
rect 659 1477 660 1481
rect 672 1480 674 1514
rect 688 1507 690 1534
rect 754 1519 760 1520
rect 754 1515 755 1519
rect 759 1515 760 1519
rect 754 1514 760 1515
rect 687 1506 691 1507
rect 687 1501 691 1502
rect 735 1506 739 1507
rect 735 1501 739 1502
rect 736 1482 738 1501
rect 734 1481 740 1482
rect 654 1476 660 1477
rect 670 1479 676 1480
rect 670 1475 671 1479
rect 675 1475 676 1479
rect 734 1477 735 1481
rect 739 1477 740 1481
rect 756 1480 758 1514
rect 776 1507 778 1534
rect 864 1507 866 1534
rect 775 1506 779 1507
rect 775 1501 779 1502
rect 815 1506 819 1507
rect 815 1501 819 1502
rect 863 1506 867 1507
rect 863 1501 867 1502
rect 816 1482 818 1501
rect 880 1500 882 1534
rect 944 1507 946 1534
rect 1016 1520 1018 1586
rect 1102 1572 1108 1573
rect 1102 1568 1103 1572
rect 1107 1568 1108 1572
rect 1102 1567 1108 1568
rect 1087 1566 1091 1567
rect 1087 1561 1091 1562
rect 1103 1566 1107 1567
rect 1103 1561 1107 1562
rect 1167 1566 1171 1567
rect 1167 1561 1171 1562
rect 1223 1566 1227 1567
rect 1223 1561 1227 1562
rect 1086 1560 1092 1561
rect 1086 1556 1087 1560
rect 1091 1556 1092 1560
rect 1086 1555 1092 1556
rect 1166 1560 1172 1561
rect 1166 1556 1167 1560
rect 1171 1556 1172 1560
rect 1166 1555 1172 1556
rect 1222 1560 1228 1561
rect 1222 1556 1223 1560
rect 1227 1556 1228 1560
rect 1222 1555 1228 1556
rect 1264 1540 1266 1602
rect 1288 1593 1290 1613
rect 1327 1609 1331 1610
rect 1367 1614 1371 1615
rect 1402 1614 1408 1615
rect 1423 1614 1427 1615
rect 1367 1609 1371 1610
rect 1423 1609 1427 1610
rect 1479 1614 1483 1615
rect 1490 1614 1496 1615
rect 1511 1614 1515 1615
rect 1479 1609 1483 1610
rect 1511 1609 1515 1610
rect 1559 1614 1563 1615
rect 1578 1614 1584 1615
rect 1599 1614 1603 1615
rect 1559 1609 1563 1610
rect 1599 1609 1603 1610
rect 1639 1614 1643 1615
rect 1674 1614 1680 1615
rect 1695 1614 1699 1615
rect 1639 1609 1643 1610
rect 1695 1609 1699 1610
rect 1719 1614 1723 1615
rect 1719 1609 1723 1610
rect 1791 1614 1795 1615
rect 1791 1609 1795 1610
rect 1799 1614 1803 1615
rect 1799 1609 1803 1610
rect 1871 1614 1875 1615
rect 1890 1614 1896 1615
rect 1911 1614 1915 1615
rect 1871 1609 1875 1610
rect 1911 1609 1915 1610
rect 1286 1592 1292 1593
rect 1286 1588 1287 1592
rect 1291 1588 1292 1592
rect 1328 1589 1330 1609
rect 1368 1590 1370 1609
rect 1390 1607 1396 1608
rect 1390 1603 1391 1607
rect 1395 1603 1396 1607
rect 1390 1602 1396 1603
rect 1366 1589 1372 1590
rect 1286 1587 1292 1588
rect 1326 1588 1332 1589
rect 1326 1584 1327 1588
rect 1331 1584 1332 1588
rect 1366 1585 1367 1589
rect 1371 1585 1372 1589
rect 1392 1588 1394 1602
rect 1424 1590 1426 1609
rect 1446 1607 1452 1608
rect 1446 1603 1447 1607
rect 1451 1603 1452 1607
rect 1446 1602 1452 1603
rect 1422 1589 1428 1590
rect 1366 1584 1372 1585
rect 1390 1587 1396 1588
rect 1326 1583 1332 1584
rect 1390 1583 1391 1587
rect 1395 1583 1396 1587
rect 1422 1585 1423 1589
rect 1427 1585 1428 1589
rect 1448 1588 1450 1602
rect 1480 1590 1482 1609
rect 1502 1607 1508 1608
rect 1502 1603 1503 1607
rect 1507 1603 1508 1607
rect 1502 1602 1508 1603
rect 1478 1589 1484 1590
rect 1422 1584 1428 1585
rect 1446 1587 1452 1588
rect 1390 1582 1396 1583
rect 1446 1583 1447 1587
rect 1451 1583 1452 1587
rect 1478 1585 1479 1589
rect 1483 1585 1484 1589
rect 1504 1588 1506 1602
rect 1560 1590 1562 1609
rect 1582 1607 1588 1608
rect 1582 1603 1583 1607
rect 1587 1603 1588 1607
rect 1582 1602 1588 1603
rect 1558 1589 1564 1590
rect 1478 1584 1484 1585
rect 1502 1587 1508 1588
rect 1446 1582 1452 1583
rect 1502 1583 1503 1587
rect 1507 1583 1508 1587
rect 1558 1585 1559 1589
rect 1563 1585 1564 1589
rect 1584 1588 1586 1602
rect 1640 1590 1642 1609
rect 1720 1590 1722 1609
rect 1792 1590 1794 1609
rect 1872 1590 1874 1609
rect 1932 1608 1934 1634
rect 2032 1624 2034 1690
rect 2094 1676 2100 1677
rect 2094 1672 2095 1676
rect 2099 1672 2100 1676
rect 2094 1671 2100 1672
rect 2182 1676 2188 1677
rect 2182 1672 2183 1676
rect 2187 1672 2188 1676
rect 2182 1671 2188 1672
rect 2270 1676 2276 1677
rect 2270 1672 2271 1676
rect 2275 1672 2276 1676
rect 2270 1671 2276 1672
rect 2366 1676 2372 1677
rect 2366 1672 2367 1676
rect 2371 1672 2372 1676
rect 2366 1671 2372 1672
rect 2438 1676 2444 1677
rect 2438 1672 2439 1676
rect 2443 1672 2444 1676
rect 2438 1671 2444 1672
rect 2096 1667 2098 1671
rect 2184 1667 2186 1671
rect 2272 1667 2274 1671
rect 2368 1667 2370 1671
rect 2440 1667 2442 1671
rect 2095 1666 2099 1667
rect 2095 1661 2099 1662
rect 2159 1666 2163 1667
rect 2159 1661 2163 1662
rect 2183 1666 2187 1667
rect 2183 1661 2187 1662
rect 2271 1666 2275 1667
rect 2271 1661 2275 1662
rect 2303 1666 2307 1667
rect 2303 1661 2307 1662
rect 2367 1666 2371 1667
rect 2367 1661 2371 1662
rect 2439 1666 2443 1667
rect 2439 1661 2443 1662
rect 2158 1660 2164 1661
rect 2158 1656 2159 1660
rect 2163 1656 2164 1660
rect 2158 1655 2164 1656
rect 2302 1660 2308 1661
rect 2302 1656 2303 1660
rect 2307 1656 2308 1660
rect 2302 1655 2308 1656
rect 2438 1660 2444 1661
rect 2438 1656 2439 1660
rect 2443 1656 2444 1660
rect 2438 1655 2444 1656
rect 2038 1639 2044 1640
rect 2038 1635 2039 1639
rect 2043 1635 2044 1639
rect 2038 1634 2044 1635
rect 2154 1639 2160 1640
rect 2154 1635 2155 1639
rect 2159 1635 2160 1639
rect 2154 1634 2160 1635
rect 2174 1639 2180 1640
rect 2174 1635 2175 1639
rect 2179 1635 2180 1639
rect 2174 1634 2180 1635
rect 2298 1639 2304 1640
rect 2298 1635 2299 1639
rect 2303 1635 2304 1639
rect 2298 1634 2304 1635
rect 2318 1639 2324 1640
rect 2318 1635 2319 1639
rect 2323 1635 2324 1639
rect 2318 1634 2324 1635
rect 2454 1639 2460 1640
rect 2454 1635 2455 1639
rect 2459 1635 2460 1639
rect 2454 1634 2460 1635
rect 2030 1623 2036 1624
rect 2030 1619 2031 1623
rect 2035 1619 2036 1623
rect 2030 1618 2036 1619
rect 2040 1615 2042 1634
rect 2156 1620 2158 1634
rect 2154 1619 2160 1620
rect 2154 1615 2155 1619
rect 2159 1615 2160 1619
rect 2176 1615 2178 1634
rect 2300 1620 2302 1634
rect 2298 1619 2304 1620
rect 2298 1615 2299 1619
rect 2303 1615 2304 1619
rect 2320 1615 2322 1634
rect 2456 1615 2458 1634
rect 2464 1620 2466 1690
rect 2476 1640 2478 1702
rect 2504 1697 2506 1717
rect 2502 1696 2508 1697
rect 2502 1692 2503 1696
rect 2507 1692 2508 1696
rect 2502 1691 2508 1692
rect 2502 1679 2508 1680
rect 2502 1675 2503 1679
rect 2507 1675 2508 1679
rect 2502 1674 2508 1675
rect 2504 1667 2506 1674
rect 2503 1666 2507 1667
rect 2503 1661 2507 1662
rect 2504 1658 2506 1661
rect 2502 1657 2508 1658
rect 2502 1653 2503 1657
rect 2507 1653 2508 1657
rect 2502 1652 2508 1653
rect 2502 1640 2508 1641
rect 2474 1639 2480 1640
rect 2474 1635 2475 1639
rect 2479 1635 2480 1639
rect 2502 1636 2503 1640
rect 2507 1636 2508 1640
rect 2502 1635 2508 1636
rect 2474 1634 2480 1635
rect 2462 1619 2468 1620
rect 2462 1615 2463 1619
rect 2467 1615 2468 1619
rect 2504 1615 2506 1635
rect 1951 1614 1955 1615
rect 1951 1609 1955 1610
rect 2031 1614 2035 1615
rect 2031 1609 2035 1610
rect 2039 1614 2043 1615
rect 2154 1614 2160 1615
rect 2175 1614 2179 1615
rect 2298 1614 2304 1615
rect 2319 1614 2323 1615
rect 2039 1609 2043 1610
rect 2175 1609 2179 1610
rect 2319 1609 2323 1610
rect 2455 1614 2459 1615
rect 2462 1614 2468 1615
rect 2503 1614 2507 1615
rect 2455 1609 2459 1610
rect 2503 1609 2507 1610
rect 1930 1607 1936 1608
rect 1930 1603 1931 1607
rect 1935 1603 1936 1607
rect 1930 1602 1936 1603
rect 1952 1590 1954 1609
rect 1974 1607 1980 1608
rect 1974 1603 1975 1607
rect 1979 1603 1980 1607
rect 1974 1602 1980 1603
rect 1638 1589 1644 1590
rect 1558 1584 1564 1585
rect 1582 1587 1588 1588
rect 1502 1582 1508 1583
rect 1582 1583 1583 1587
rect 1587 1583 1588 1587
rect 1638 1585 1639 1589
rect 1643 1585 1644 1589
rect 1638 1584 1644 1585
rect 1718 1589 1724 1590
rect 1718 1585 1719 1589
rect 1723 1585 1724 1589
rect 1790 1589 1796 1590
rect 1718 1584 1724 1585
rect 1742 1587 1748 1588
rect 1582 1582 1588 1583
rect 1742 1583 1743 1587
rect 1747 1583 1748 1587
rect 1790 1585 1791 1589
rect 1795 1585 1796 1589
rect 1790 1584 1796 1585
rect 1870 1589 1876 1590
rect 1870 1585 1871 1589
rect 1875 1585 1876 1589
rect 1870 1584 1876 1585
rect 1950 1589 1956 1590
rect 1950 1585 1951 1589
rect 1955 1585 1956 1589
rect 1976 1588 1978 1602
rect 2032 1590 2034 1609
rect 2030 1589 2036 1590
rect 2504 1589 2506 1609
rect 1950 1584 1956 1585
rect 1974 1587 1980 1588
rect 1742 1582 1748 1583
rect 1974 1583 1975 1587
rect 1979 1583 1980 1587
rect 2030 1585 2031 1589
rect 2035 1585 2036 1589
rect 2030 1584 2036 1585
rect 2502 1588 2508 1589
rect 2502 1584 2503 1588
rect 2507 1584 2508 1588
rect 2502 1583 2508 1584
rect 1974 1582 1980 1583
rect 1286 1575 1292 1576
rect 1286 1571 1287 1575
rect 1291 1571 1292 1575
rect 1286 1570 1292 1571
rect 1326 1571 1332 1572
rect 1288 1567 1290 1570
rect 1326 1567 1327 1571
rect 1331 1567 1332 1571
rect 1287 1566 1291 1567
rect 1326 1566 1332 1567
rect 1350 1568 1356 1569
rect 1328 1563 1330 1566
rect 1350 1564 1351 1568
rect 1355 1564 1356 1568
rect 1350 1563 1356 1564
rect 1406 1568 1412 1569
rect 1406 1564 1407 1568
rect 1411 1564 1412 1568
rect 1406 1563 1412 1564
rect 1462 1568 1468 1569
rect 1462 1564 1463 1568
rect 1467 1564 1468 1568
rect 1462 1563 1468 1564
rect 1542 1568 1548 1569
rect 1542 1564 1543 1568
rect 1547 1564 1548 1568
rect 1542 1563 1548 1564
rect 1622 1568 1628 1569
rect 1622 1564 1623 1568
rect 1627 1564 1628 1568
rect 1622 1563 1628 1564
rect 1702 1568 1708 1569
rect 1702 1564 1703 1568
rect 1707 1564 1708 1568
rect 1702 1563 1708 1564
rect 1287 1561 1291 1562
rect 1327 1562 1331 1563
rect 1288 1558 1290 1561
rect 1286 1557 1292 1558
rect 1327 1557 1331 1558
rect 1351 1562 1355 1563
rect 1351 1557 1355 1558
rect 1407 1562 1411 1563
rect 1407 1557 1411 1558
rect 1463 1562 1467 1563
rect 1463 1557 1467 1558
rect 1471 1562 1475 1563
rect 1471 1557 1475 1558
rect 1543 1562 1547 1563
rect 1543 1557 1547 1558
rect 1607 1562 1611 1563
rect 1607 1557 1611 1558
rect 1623 1562 1627 1563
rect 1623 1557 1627 1558
rect 1703 1562 1707 1563
rect 1703 1557 1707 1558
rect 1735 1562 1739 1563
rect 1735 1557 1739 1558
rect 1286 1553 1287 1557
rect 1291 1553 1292 1557
rect 1328 1554 1330 1557
rect 1350 1556 1356 1557
rect 1286 1552 1292 1553
rect 1326 1553 1332 1554
rect 1326 1549 1327 1553
rect 1331 1549 1332 1553
rect 1350 1552 1351 1556
rect 1355 1552 1356 1556
rect 1350 1551 1356 1552
rect 1470 1556 1476 1557
rect 1470 1552 1471 1556
rect 1475 1552 1476 1556
rect 1470 1551 1476 1552
rect 1606 1556 1612 1557
rect 1606 1552 1607 1556
rect 1611 1552 1612 1556
rect 1606 1551 1612 1552
rect 1734 1556 1740 1557
rect 1734 1552 1735 1556
rect 1739 1552 1740 1556
rect 1734 1551 1740 1552
rect 1326 1548 1332 1549
rect 1286 1540 1292 1541
rect 1022 1539 1028 1540
rect 1022 1535 1023 1539
rect 1027 1535 1028 1539
rect 1022 1534 1028 1535
rect 1102 1539 1108 1540
rect 1102 1535 1103 1539
rect 1107 1535 1108 1539
rect 1102 1534 1108 1535
rect 1162 1539 1168 1540
rect 1162 1535 1163 1539
rect 1167 1535 1168 1539
rect 1162 1534 1168 1535
rect 1182 1539 1188 1540
rect 1182 1535 1183 1539
rect 1187 1535 1188 1539
rect 1182 1534 1188 1535
rect 1218 1539 1224 1540
rect 1218 1535 1219 1539
rect 1223 1535 1224 1539
rect 1218 1534 1224 1535
rect 1238 1539 1244 1540
rect 1238 1535 1239 1539
rect 1243 1535 1244 1539
rect 1238 1534 1244 1535
rect 1262 1539 1268 1540
rect 1262 1535 1263 1539
rect 1267 1535 1268 1539
rect 1286 1536 1287 1540
rect 1291 1536 1292 1540
rect 1286 1535 1292 1536
rect 1326 1536 1332 1537
rect 1262 1534 1268 1535
rect 1014 1519 1020 1520
rect 1014 1515 1015 1519
rect 1019 1515 1020 1519
rect 1014 1514 1020 1515
rect 1024 1507 1026 1534
rect 1104 1507 1106 1534
rect 1164 1520 1166 1534
rect 1162 1519 1168 1520
rect 1162 1515 1163 1519
rect 1167 1515 1168 1519
rect 1162 1514 1168 1515
rect 1184 1507 1186 1534
rect 1220 1520 1222 1534
rect 1218 1519 1224 1520
rect 1218 1515 1219 1519
rect 1223 1515 1224 1519
rect 1218 1514 1224 1515
rect 1240 1507 1242 1534
rect 1288 1507 1290 1535
rect 1326 1532 1327 1536
rect 1331 1532 1332 1536
rect 1326 1531 1332 1532
rect 1366 1535 1372 1536
rect 1366 1531 1367 1535
rect 1371 1531 1372 1535
rect 1328 1511 1330 1531
rect 1366 1530 1372 1531
rect 1486 1535 1492 1536
rect 1486 1531 1487 1535
rect 1491 1531 1492 1535
rect 1486 1530 1492 1531
rect 1602 1535 1608 1536
rect 1602 1531 1603 1535
rect 1607 1531 1608 1535
rect 1602 1530 1608 1531
rect 1622 1535 1628 1536
rect 1622 1531 1623 1535
rect 1627 1531 1628 1535
rect 1622 1530 1628 1531
rect 1730 1535 1736 1536
rect 1730 1531 1731 1535
rect 1735 1531 1736 1535
rect 1730 1530 1736 1531
rect 1368 1511 1370 1530
rect 1386 1515 1392 1516
rect 1386 1511 1387 1515
rect 1391 1511 1392 1515
rect 1488 1511 1490 1530
rect 1604 1516 1606 1530
rect 1602 1515 1608 1516
rect 1602 1511 1603 1515
rect 1607 1511 1608 1515
rect 1624 1511 1626 1530
rect 1732 1516 1734 1530
rect 1744 1524 1746 1582
rect 2502 1571 2508 1572
rect 1774 1568 1780 1569
rect 1774 1564 1775 1568
rect 1779 1564 1780 1568
rect 1774 1563 1780 1564
rect 1854 1568 1860 1569
rect 1854 1564 1855 1568
rect 1859 1564 1860 1568
rect 1854 1563 1860 1564
rect 1934 1568 1940 1569
rect 1934 1564 1935 1568
rect 1939 1564 1940 1568
rect 1934 1563 1940 1564
rect 2014 1568 2020 1569
rect 2014 1564 2015 1568
rect 2019 1564 2020 1568
rect 2502 1567 2503 1571
rect 2507 1567 2508 1571
rect 2502 1566 2508 1567
rect 2014 1563 2020 1564
rect 2504 1563 2506 1566
rect 1775 1562 1779 1563
rect 1775 1557 1779 1558
rect 1855 1562 1859 1563
rect 1855 1557 1859 1558
rect 1871 1562 1875 1563
rect 1871 1557 1875 1558
rect 1935 1562 1939 1563
rect 1935 1557 1939 1558
rect 2007 1562 2011 1563
rect 2007 1557 2011 1558
rect 2015 1562 2019 1563
rect 2015 1557 2019 1558
rect 2503 1562 2507 1563
rect 2503 1557 2507 1558
rect 1870 1556 1876 1557
rect 1870 1552 1871 1556
rect 1875 1552 1876 1556
rect 1870 1551 1876 1552
rect 2006 1556 2012 1557
rect 2006 1552 2007 1556
rect 2011 1552 2012 1556
rect 2504 1554 2506 1557
rect 2006 1551 2012 1552
rect 2502 1553 2508 1554
rect 2502 1549 2503 1553
rect 2507 1549 2508 1553
rect 2502 1548 2508 1549
rect 2502 1536 2508 1537
rect 1750 1535 1756 1536
rect 1750 1531 1751 1535
rect 1755 1531 1756 1535
rect 1750 1530 1756 1531
rect 1862 1535 1868 1536
rect 1862 1531 1863 1535
rect 1867 1531 1868 1535
rect 1862 1530 1868 1531
rect 1886 1535 1892 1536
rect 1886 1531 1887 1535
rect 1891 1531 1892 1535
rect 1886 1530 1892 1531
rect 2002 1535 2008 1536
rect 2002 1531 2003 1535
rect 2007 1531 2008 1535
rect 2002 1530 2008 1531
rect 2022 1535 2028 1536
rect 2022 1531 2023 1535
rect 2027 1531 2028 1535
rect 2502 1532 2503 1536
rect 2507 1532 2508 1536
rect 2502 1531 2508 1532
rect 2022 1530 2028 1531
rect 1742 1523 1748 1524
rect 1742 1519 1743 1523
rect 1747 1519 1748 1523
rect 1742 1518 1748 1519
rect 1730 1515 1736 1516
rect 1730 1511 1731 1515
rect 1735 1511 1736 1515
rect 1752 1511 1754 1530
rect 1774 1527 1780 1528
rect 1774 1523 1775 1527
rect 1779 1523 1780 1527
rect 1774 1522 1780 1523
rect 1327 1510 1331 1511
rect 895 1506 899 1507
rect 895 1501 899 1502
rect 943 1506 947 1507
rect 943 1501 947 1502
rect 975 1506 979 1507
rect 975 1501 979 1502
rect 1023 1506 1027 1507
rect 1023 1501 1027 1502
rect 1055 1506 1059 1507
rect 1055 1501 1059 1502
rect 1103 1506 1107 1507
rect 1103 1501 1107 1502
rect 1143 1506 1147 1507
rect 1143 1501 1147 1502
rect 1183 1506 1187 1507
rect 1183 1501 1187 1502
rect 1239 1506 1243 1507
rect 1239 1501 1243 1502
rect 1287 1506 1291 1507
rect 1327 1505 1331 1506
rect 1367 1510 1371 1511
rect 1386 1510 1392 1511
rect 1423 1510 1427 1511
rect 1367 1505 1371 1506
rect 1287 1501 1291 1502
rect 850 1499 856 1500
rect 850 1495 851 1499
rect 855 1495 856 1499
rect 850 1494 856 1495
rect 878 1499 884 1500
rect 878 1495 879 1499
rect 883 1495 884 1499
rect 878 1494 884 1495
rect 814 1481 820 1482
rect 734 1476 740 1477
rect 754 1479 760 1480
rect 670 1474 676 1475
rect 754 1475 755 1479
rect 759 1475 760 1479
rect 814 1477 815 1481
rect 819 1477 820 1481
rect 814 1476 820 1477
rect 754 1474 760 1475
rect 638 1460 644 1461
rect 638 1456 639 1460
rect 643 1456 644 1460
rect 638 1455 644 1456
rect 718 1460 724 1461
rect 718 1456 719 1460
rect 723 1456 724 1460
rect 718 1455 724 1456
rect 798 1460 804 1461
rect 798 1456 799 1460
rect 803 1456 804 1460
rect 798 1455 804 1456
rect 640 1451 642 1455
rect 720 1451 722 1455
rect 800 1451 802 1455
rect 639 1450 643 1451
rect 639 1445 643 1446
rect 711 1450 715 1451
rect 711 1445 715 1446
rect 719 1450 723 1451
rect 719 1445 723 1446
rect 799 1450 803 1451
rect 799 1445 803 1446
rect 815 1450 819 1451
rect 815 1445 819 1446
rect 710 1444 716 1445
rect 710 1440 711 1444
rect 715 1440 716 1444
rect 710 1439 716 1440
rect 814 1444 820 1445
rect 814 1440 815 1444
rect 819 1440 820 1444
rect 814 1439 820 1440
rect 852 1424 854 1494
rect 896 1482 898 1501
rect 934 1499 940 1500
rect 934 1495 935 1499
rect 939 1495 940 1499
rect 934 1494 940 1495
rect 894 1481 900 1482
rect 894 1477 895 1481
rect 899 1477 900 1481
rect 936 1480 938 1494
rect 976 1482 978 1501
rect 998 1499 1004 1500
rect 998 1495 999 1499
rect 1003 1495 1004 1499
rect 998 1494 1004 1495
rect 974 1481 980 1482
rect 894 1476 900 1477
rect 934 1479 940 1480
rect 934 1475 935 1479
rect 939 1475 940 1479
rect 974 1477 975 1481
rect 979 1477 980 1481
rect 1000 1480 1002 1494
rect 1056 1482 1058 1501
rect 1078 1499 1084 1500
rect 1078 1495 1079 1499
rect 1083 1495 1084 1499
rect 1078 1494 1084 1495
rect 1054 1481 1060 1482
rect 974 1476 980 1477
rect 998 1479 1004 1480
rect 934 1474 940 1475
rect 998 1475 999 1479
rect 1003 1475 1004 1479
rect 1054 1477 1055 1481
rect 1059 1477 1060 1481
rect 1080 1480 1082 1494
rect 1144 1482 1146 1501
rect 1142 1481 1148 1482
rect 1288 1481 1290 1501
rect 1328 1485 1330 1505
rect 1368 1486 1370 1505
rect 1366 1485 1372 1486
rect 1326 1484 1332 1485
rect 1054 1476 1060 1477
rect 1078 1479 1084 1480
rect 998 1474 1004 1475
rect 1078 1475 1079 1479
rect 1083 1475 1084 1479
rect 1142 1477 1143 1481
rect 1147 1477 1148 1481
rect 1286 1480 1292 1481
rect 1142 1476 1148 1477
rect 1150 1479 1156 1480
rect 1078 1474 1084 1475
rect 1150 1475 1151 1479
rect 1155 1475 1156 1479
rect 1286 1476 1287 1480
rect 1291 1476 1292 1480
rect 1326 1480 1327 1484
rect 1331 1480 1332 1484
rect 1366 1481 1367 1485
rect 1371 1481 1372 1485
rect 1388 1484 1390 1510
rect 1423 1505 1427 1506
rect 1479 1510 1483 1511
rect 1479 1505 1483 1506
rect 1487 1510 1491 1511
rect 1487 1505 1491 1506
rect 1551 1510 1555 1511
rect 1602 1510 1608 1511
rect 1623 1510 1627 1511
rect 1551 1505 1555 1506
rect 1623 1505 1627 1506
rect 1631 1510 1635 1511
rect 1631 1505 1635 1506
rect 1711 1510 1715 1511
rect 1730 1510 1736 1511
rect 1751 1510 1755 1511
rect 1711 1505 1715 1506
rect 1751 1505 1755 1506
rect 1424 1486 1426 1505
rect 1480 1486 1482 1505
rect 1552 1486 1554 1505
rect 1566 1503 1572 1504
rect 1566 1499 1567 1503
rect 1571 1499 1572 1503
rect 1566 1498 1572 1499
rect 1574 1503 1580 1504
rect 1574 1499 1575 1503
rect 1579 1499 1580 1503
rect 1574 1498 1580 1499
rect 1422 1485 1428 1486
rect 1366 1480 1372 1481
rect 1386 1483 1392 1484
rect 1326 1479 1332 1480
rect 1386 1479 1387 1483
rect 1391 1479 1392 1483
rect 1422 1481 1423 1485
rect 1427 1481 1428 1485
rect 1422 1480 1428 1481
rect 1478 1485 1484 1486
rect 1478 1481 1479 1485
rect 1483 1481 1484 1485
rect 1478 1480 1484 1481
rect 1550 1485 1556 1486
rect 1550 1481 1551 1485
rect 1555 1481 1556 1485
rect 1550 1480 1556 1481
rect 1386 1478 1392 1479
rect 1286 1475 1292 1476
rect 1150 1474 1156 1475
rect 878 1460 884 1461
rect 878 1456 879 1460
rect 883 1456 884 1460
rect 878 1455 884 1456
rect 958 1460 964 1461
rect 958 1456 959 1460
rect 963 1456 964 1460
rect 958 1455 964 1456
rect 1038 1460 1044 1461
rect 1038 1456 1039 1460
rect 1043 1456 1044 1460
rect 1038 1455 1044 1456
rect 1126 1460 1132 1461
rect 1126 1456 1127 1460
rect 1131 1456 1132 1460
rect 1126 1455 1132 1456
rect 880 1451 882 1455
rect 960 1451 962 1455
rect 1040 1451 1042 1455
rect 1128 1451 1130 1455
rect 879 1450 883 1451
rect 879 1445 883 1446
rect 919 1450 923 1451
rect 919 1445 923 1446
rect 959 1450 963 1451
rect 959 1445 963 1446
rect 1023 1450 1027 1451
rect 1023 1445 1027 1446
rect 1039 1450 1043 1451
rect 1039 1445 1043 1446
rect 1127 1450 1131 1451
rect 1127 1445 1131 1446
rect 918 1444 924 1445
rect 918 1440 919 1444
rect 923 1440 924 1444
rect 918 1439 924 1440
rect 1022 1444 1028 1445
rect 1022 1440 1023 1444
rect 1027 1440 1028 1444
rect 1022 1439 1028 1440
rect 1126 1444 1132 1445
rect 1126 1440 1127 1444
rect 1131 1440 1132 1444
rect 1126 1439 1132 1440
rect 518 1423 524 1424
rect 518 1419 519 1423
rect 523 1419 524 1423
rect 518 1418 524 1419
rect 622 1423 628 1424
rect 622 1419 623 1423
rect 627 1419 628 1423
rect 622 1418 628 1419
rect 630 1423 636 1424
rect 630 1419 631 1423
rect 635 1419 636 1423
rect 630 1418 636 1419
rect 726 1423 732 1424
rect 726 1419 727 1423
rect 731 1419 732 1423
rect 726 1418 732 1419
rect 830 1423 836 1424
rect 830 1419 831 1423
rect 835 1419 836 1423
rect 830 1418 836 1419
rect 850 1423 856 1424
rect 850 1419 851 1423
rect 855 1419 856 1423
rect 850 1418 856 1419
rect 934 1423 940 1424
rect 934 1419 935 1423
rect 939 1419 940 1423
rect 934 1418 940 1419
rect 1018 1423 1024 1424
rect 1018 1419 1019 1423
rect 1023 1419 1024 1423
rect 1018 1418 1024 1419
rect 1038 1423 1044 1424
rect 1038 1419 1039 1423
rect 1043 1419 1044 1423
rect 1038 1418 1044 1419
rect 1122 1423 1128 1424
rect 1122 1419 1123 1423
rect 1127 1419 1128 1423
rect 1122 1418 1128 1419
rect 1142 1423 1148 1424
rect 1142 1419 1143 1423
rect 1147 1419 1148 1423
rect 1142 1418 1148 1419
rect 510 1403 516 1404
rect 510 1399 511 1403
rect 515 1399 516 1403
rect 510 1398 516 1399
rect 520 1395 522 1418
rect 624 1395 626 1418
rect 686 1403 692 1404
rect 686 1399 687 1403
rect 691 1399 692 1403
rect 686 1398 692 1399
rect 111 1394 115 1395
rect 111 1389 115 1390
rect 151 1394 155 1395
rect 151 1389 155 1390
rect 207 1394 211 1395
rect 214 1391 215 1395
rect 219 1391 220 1395
rect 214 1390 220 1391
rect 223 1394 227 1395
rect 207 1389 211 1390
rect 223 1389 227 1390
rect 271 1394 275 1395
rect 271 1389 275 1390
rect 295 1394 299 1395
rect 295 1389 299 1390
rect 343 1394 347 1395
rect 350 1391 351 1395
rect 355 1391 356 1395
rect 350 1390 356 1391
rect 359 1394 363 1395
rect 343 1389 347 1390
rect 359 1389 363 1390
rect 423 1394 427 1395
rect 423 1389 427 1390
rect 431 1394 435 1395
rect 431 1389 435 1390
rect 503 1394 507 1395
rect 503 1389 507 1390
rect 519 1394 523 1395
rect 519 1389 523 1390
rect 583 1394 587 1395
rect 583 1389 587 1390
rect 623 1394 627 1395
rect 623 1389 627 1390
rect 663 1394 667 1395
rect 663 1389 667 1390
rect 112 1369 114 1389
rect 152 1370 154 1389
rect 174 1387 180 1388
rect 174 1383 175 1387
rect 179 1383 180 1387
rect 174 1382 180 1383
rect 150 1369 156 1370
rect 110 1368 116 1369
rect 110 1364 111 1368
rect 115 1364 116 1368
rect 150 1365 151 1369
rect 155 1365 156 1369
rect 176 1368 178 1382
rect 224 1370 226 1389
rect 296 1370 298 1389
rect 360 1370 362 1389
rect 382 1387 388 1388
rect 382 1383 383 1387
rect 387 1383 388 1387
rect 382 1382 388 1383
rect 222 1369 228 1370
rect 150 1364 156 1365
rect 174 1367 180 1368
rect 110 1363 116 1364
rect 174 1363 175 1367
rect 179 1363 180 1367
rect 222 1365 223 1369
rect 227 1365 228 1369
rect 294 1369 300 1370
rect 222 1364 228 1365
rect 246 1367 252 1368
rect 174 1362 180 1363
rect 246 1363 247 1367
rect 251 1363 252 1367
rect 294 1365 295 1369
rect 299 1365 300 1369
rect 294 1364 300 1365
rect 358 1369 364 1370
rect 358 1365 359 1369
rect 363 1365 364 1369
rect 384 1368 386 1382
rect 432 1370 434 1389
rect 462 1387 468 1388
rect 462 1383 463 1387
rect 467 1383 468 1387
rect 462 1382 468 1383
rect 430 1369 436 1370
rect 358 1364 364 1365
rect 382 1367 388 1368
rect 246 1362 252 1363
rect 382 1363 383 1367
rect 387 1363 388 1367
rect 430 1365 431 1369
rect 435 1365 436 1369
rect 464 1368 466 1382
rect 504 1370 506 1389
rect 526 1387 532 1388
rect 526 1383 527 1387
rect 531 1383 532 1387
rect 526 1382 532 1383
rect 502 1369 508 1370
rect 430 1364 436 1365
rect 462 1367 468 1368
rect 382 1362 388 1363
rect 462 1363 463 1367
rect 467 1363 468 1367
rect 502 1365 503 1369
rect 507 1365 508 1369
rect 528 1368 530 1382
rect 584 1370 586 1389
rect 606 1387 612 1388
rect 606 1383 607 1387
rect 611 1383 612 1387
rect 606 1382 612 1383
rect 654 1387 660 1388
rect 654 1383 655 1387
rect 659 1383 660 1387
rect 654 1382 660 1383
rect 582 1369 588 1370
rect 502 1364 508 1365
rect 526 1367 532 1368
rect 462 1362 468 1363
rect 526 1363 527 1367
rect 531 1363 532 1367
rect 582 1365 583 1369
rect 587 1365 588 1369
rect 608 1368 610 1382
rect 582 1364 588 1365
rect 606 1367 612 1368
rect 526 1362 532 1363
rect 606 1363 607 1367
rect 611 1363 612 1367
rect 606 1362 612 1363
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 110 1346 116 1347
rect 134 1348 140 1349
rect 112 1327 114 1346
rect 134 1344 135 1348
rect 139 1344 140 1348
rect 134 1343 140 1344
rect 206 1348 212 1349
rect 206 1344 207 1348
rect 211 1344 212 1348
rect 206 1343 212 1344
rect 136 1327 138 1343
rect 208 1327 210 1343
rect 111 1326 115 1327
rect 111 1321 115 1322
rect 135 1326 139 1327
rect 135 1321 139 1322
rect 207 1326 211 1327
rect 207 1321 211 1322
rect 239 1326 243 1327
rect 239 1321 243 1322
rect 112 1318 114 1321
rect 134 1320 140 1321
rect 110 1317 116 1318
rect 110 1313 111 1317
rect 115 1313 116 1317
rect 134 1316 135 1320
rect 139 1316 140 1320
rect 134 1315 140 1316
rect 238 1320 244 1321
rect 238 1316 239 1320
rect 243 1316 244 1320
rect 238 1315 244 1316
rect 110 1312 116 1313
rect 110 1300 116 1301
rect 110 1296 111 1300
rect 115 1296 116 1300
rect 110 1295 116 1296
rect 150 1299 156 1300
rect 150 1295 151 1299
rect 155 1295 156 1299
rect 112 1267 114 1295
rect 150 1294 156 1295
rect 158 1299 164 1300
rect 158 1295 159 1299
rect 163 1295 164 1299
rect 158 1294 164 1295
rect 152 1267 154 1294
rect 111 1266 115 1267
rect 111 1261 115 1262
rect 151 1266 155 1267
rect 151 1261 155 1262
rect 112 1241 114 1261
rect 152 1242 154 1261
rect 160 1260 162 1294
rect 248 1280 250 1362
rect 278 1348 284 1349
rect 278 1344 279 1348
rect 283 1344 284 1348
rect 278 1343 284 1344
rect 342 1348 348 1349
rect 342 1344 343 1348
rect 347 1344 348 1348
rect 342 1343 348 1344
rect 414 1348 420 1349
rect 414 1344 415 1348
rect 419 1344 420 1348
rect 414 1343 420 1344
rect 486 1348 492 1349
rect 486 1344 487 1348
rect 491 1344 492 1348
rect 486 1343 492 1344
rect 566 1348 572 1349
rect 566 1344 567 1348
rect 571 1344 572 1348
rect 566 1343 572 1344
rect 646 1348 652 1349
rect 646 1344 647 1348
rect 651 1344 652 1348
rect 646 1343 652 1344
rect 280 1327 282 1343
rect 344 1327 346 1343
rect 416 1327 418 1343
rect 488 1327 490 1343
rect 568 1327 570 1343
rect 648 1327 650 1343
rect 279 1326 283 1327
rect 279 1321 283 1322
rect 343 1326 347 1327
rect 343 1321 347 1322
rect 367 1326 371 1327
rect 367 1321 371 1322
rect 415 1326 419 1327
rect 415 1321 419 1322
rect 479 1326 483 1327
rect 479 1321 483 1322
rect 487 1326 491 1327
rect 487 1321 491 1322
rect 567 1326 571 1327
rect 567 1321 571 1322
rect 583 1326 587 1327
rect 583 1321 587 1322
rect 647 1326 651 1327
rect 647 1321 651 1322
rect 366 1320 372 1321
rect 366 1316 367 1320
rect 371 1316 372 1320
rect 366 1315 372 1316
rect 478 1320 484 1321
rect 478 1316 479 1320
rect 483 1316 484 1320
rect 478 1315 484 1316
rect 582 1320 588 1321
rect 582 1316 583 1320
rect 587 1316 588 1320
rect 582 1315 588 1316
rect 656 1300 658 1382
rect 664 1370 666 1389
rect 662 1369 668 1370
rect 662 1365 663 1369
rect 667 1365 668 1369
rect 688 1368 690 1398
rect 728 1395 730 1418
rect 832 1395 834 1418
rect 858 1403 864 1404
rect 858 1399 859 1403
rect 863 1399 864 1403
rect 858 1398 864 1399
rect 727 1394 731 1395
rect 727 1389 731 1390
rect 751 1394 755 1395
rect 751 1389 755 1390
rect 831 1394 835 1395
rect 831 1389 835 1390
rect 839 1394 843 1395
rect 839 1389 843 1390
rect 752 1370 754 1389
rect 774 1387 780 1388
rect 774 1383 775 1387
rect 779 1383 780 1387
rect 774 1382 780 1383
rect 750 1369 756 1370
rect 662 1364 668 1365
rect 686 1367 692 1368
rect 686 1363 687 1367
rect 691 1363 692 1367
rect 750 1365 751 1369
rect 755 1365 756 1369
rect 776 1368 778 1382
rect 840 1370 842 1389
rect 838 1369 844 1370
rect 750 1364 756 1365
rect 774 1367 780 1368
rect 686 1362 692 1363
rect 774 1363 775 1367
rect 779 1363 780 1367
rect 838 1365 839 1369
rect 843 1365 844 1369
rect 860 1368 862 1398
rect 936 1395 938 1418
rect 1020 1404 1022 1418
rect 1018 1403 1024 1404
rect 1018 1399 1019 1403
rect 1023 1399 1024 1403
rect 1018 1398 1024 1399
rect 1040 1395 1042 1418
rect 1124 1404 1126 1418
rect 1122 1403 1128 1404
rect 1122 1399 1123 1403
rect 1127 1399 1128 1403
rect 1122 1398 1128 1399
rect 1144 1395 1146 1418
rect 1152 1412 1154 1474
rect 1326 1467 1332 1468
rect 1286 1463 1292 1464
rect 1286 1459 1287 1463
rect 1291 1459 1292 1463
rect 1326 1463 1327 1467
rect 1331 1463 1332 1467
rect 1326 1462 1332 1463
rect 1350 1464 1356 1465
rect 1286 1458 1292 1459
rect 1288 1451 1290 1458
rect 1328 1451 1330 1462
rect 1350 1460 1351 1464
rect 1355 1460 1356 1464
rect 1350 1459 1356 1460
rect 1406 1464 1412 1465
rect 1406 1460 1407 1464
rect 1411 1460 1412 1464
rect 1406 1459 1412 1460
rect 1462 1464 1468 1465
rect 1462 1460 1463 1464
rect 1467 1460 1468 1464
rect 1462 1459 1468 1460
rect 1534 1464 1540 1465
rect 1534 1460 1535 1464
rect 1539 1460 1540 1464
rect 1534 1459 1540 1460
rect 1352 1451 1354 1459
rect 1408 1451 1410 1459
rect 1464 1451 1466 1459
rect 1536 1451 1538 1459
rect 1223 1450 1227 1451
rect 1223 1445 1227 1446
rect 1287 1450 1291 1451
rect 1287 1445 1291 1446
rect 1327 1450 1331 1451
rect 1327 1445 1331 1446
rect 1351 1450 1355 1451
rect 1351 1445 1355 1446
rect 1359 1450 1363 1451
rect 1359 1445 1363 1446
rect 1407 1450 1411 1451
rect 1407 1445 1411 1446
rect 1447 1450 1451 1451
rect 1447 1445 1451 1446
rect 1463 1450 1467 1451
rect 1463 1445 1467 1446
rect 1535 1450 1539 1451
rect 1535 1445 1539 1446
rect 1222 1444 1228 1445
rect 1222 1440 1223 1444
rect 1227 1440 1228 1444
rect 1288 1442 1290 1445
rect 1328 1442 1330 1445
rect 1358 1444 1364 1445
rect 1222 1439 1228 1440
rect 1286 1441 1292 1442
rect 1286 1437 1287 1441
rect 1291 1437 1292 1441
rect 1286 1436 1292 1437
rect 1326 1441 1332 1442
rect 1326 1437 1327 1441
rect 1331 1437 1332 1441
rect 1358 1440 1359 1444
rect 1363 1440 1364 1444
rect 1358 1439 1364 1440
rect 1446 1444 1452 1445
rect 1446 1440 1447 1444
rect 1451 1440 1452 1444
rect 1446 1439 1452 1440
rect 1534 1444 1540 1445
rect 1534 1440 1535 1444
rect 1539 1440 1540 1444
rect 1534 1439 1540 1440
rect 1326 1436 1332 1437
rect 1286 1424 1292 1425
rect 1218 1423 1224 1424
rect 1218 1419 1219 1423
rect 1223 1419 1224 1423
rect 1218 1418 1224 1419
rect 1238 1423 1244 1424
rect 1238 1419 1239 1423
rect 1243 1419 1244 1423
rect 1238 1418 1244 1419
rect 1246 1423 1252 1424
rect 1246 1419 1247 1423
rect 1251 1419 1252 1423
rect 1286 1420 1287 1424
rect 1291 1420 1292 1424
rect 1286 1419 1292 1420
rect 1326 1424 1332 1425
rect 1568 1424 1570 1498
rect 1576 1484 1578 1498
rect 1632 1486 1634 1505
rect 1654 1503 1660 1504
rect 1654 1499 1655 1503
rect 1659 1499 1660 1503
rect 1654 1498 1660 1499
rect 1630 1485 1636 1486
rect 1574 1483 1580 1484
rect 1574 1479 1575 1483
rect 1579 1479 1580 1483
rect 1630 1481 1631 1485
rect 1635 1481 1636 1485
rect 1656 1484 1658 1498
rect 1712 1486 1714 1505
rect 1776 1504 1778 1522
rect 1864 1516 1866 1530
rect 1862 1515 1868 1516
rect 1862 1511 1863 1515
rect 1867 1511 1868 1515
rect 1888 1511 1890 1530
rect 2004 1516 2006 1530
rect 2002 1515 2008 1516
rect 2002 1511 2003 1515
rect 2007 1511 2008 1515
rect 2024 1511 2026 1530
rect 2504 1511 2506 1531
rect 1791 1510 1795 1511
rect 1862 1510 1868 1511
rect 1871 1510 1875 1511
rect 1791 1505 1795 1506
rect 1871 1505 1875 1506
rect 1887 1510 1891 1511
rect 1887 1505 1891 1506
rect 1951 1510 1955 1511
rect 2002 1510 2008 1511
rect 2023 1510 2027 1511
rect 1951 1505 1955 1506
rect 2023 1505 2027 1506
rect 2031 1510 2035 1511
rect 2031 1505 2035 1506
rect 2119 1510 2123 1511
rect 2119 1505 2123 1506
rect 2503 1510 2507 1511
rect 2503 1505 2507 1506
rect 1774 1503 1780 1504
rect 1774 1499 1775 1503
rect 1779 1499 1780 1503
rect 1774 1498 1780 1499
rect 1792 1486 1794 1505
rect 1814 1503 1820 1504
rect 1814 1499 1815 1503
rect 1819 1499 1820 1503
rect 1814 1498 1820 1499
rect 1710 1485 1716 1486
rect 1630 1480 1636 1481
rect 1654 1483 1660 1484
rect 1574 1478 1580 1479
rect 1654 1479 1655 1483
rect 1659 1479 1660 1483
rect 1710 1481 1711 1485
rect 1715 1481 1716 1485
rect 1710 1480 1716 1481
rect 1790 1485 1796 1486
rect 1790 1481 1791 1485
rect 1795 1481 1796 1485
rect 1816 1484 1818 1498
rect 1822 1491 1828 1492
rect 1822 1487 1823 1491
rect 1827 1487 1828 1491
rect 1822 1486 1828 1487
rect 1872 1486 1874 1505
rect 1894 1503 1900 1504
rect 1894 1499 1895 1503
rect 1899 1499 1900 1503
rect 1894 1498 1900 1499
rect 1790 1480 1796 1481
rect 1814 1483 1820 1484
rect 1654 1478 1660 1479
rect 1814 1479 1815 1483
rect 1819 1479 1820 1483
rect 1814 1478 1820 1479
rect 1614 1464 1620 1465
rect 1614 1460 1615 1464
rect 1619 1460 1620 1464
rect 1614 1459 1620 1460
rect 1694 1464 1700 1465
rect 1694 1460 1695 1464
rect 1699 1460 1700 1464
rect 1694 1459 1700 1460
rect 1774 1464 1780 1465
rect 1774 1460 1775 1464
rect 1779 1460 1780 1464
rect 1774 1459 1780 1460
rect 1616 1451 1618 1459
rect 1696 1451 1698 1459
rect 1776 1451 1778 1459
rect 1615 1450 1619 1451
rect 1615 1445 1619 1446
rect 1631 1450 1635 1451
rect 1631 1445 1635 1446
rect 1695 1450 1699 1451
rect 1695 1445 1699 1446
rect 1727 1450 1731 1451
rect 1727 1445 1731 1446
rect 1775 1450 1779 1451
rect 1775 1445 1779 1446
rect 1815 1450 1819 1451
rect 1815 1445 1819 1446
rect 1630 1444 1636 1445
rect 1630 1440 1631 1444
rect 1635 1440 1636 1444
rect 1630 1439 1636 1440
rect 1726 1444 1732 1445
rect 1726 1440 1727 1444
rect 1731 1440 1732 1444
rect 1726 1439 1732 1440
rect 1814 1444 1820 1445
rect 1814 1440 1815 1444
rect 1819 1440 1820 1444
rect 1814 1439 1820 1440
rect 1326 1420 1327 1424
rect 1331 1420 1332 1424
rect 1326 1419 1332 1420
rect 1374 1423 1380 1424
rect 1374 1419 1375 1423
rect 1379 1419 1380 1423
rect 1246 1418 1252 1419
rect 1150 1411 1156 1412
rect 1150 1407 1151 1411
rect 1155 1407 1156 1411
rect 1150 1406 1156 1407
rect 1220 1404 1222 1418
rect 1218 1403 1224 1404
rect 1218 1399 1219 1403
rect 1223 1399 1224 1403
rect 1218 1398 1224 1399
rect 1240 1395 1242 1418
rect 927 1394 931 1395
rect 927 1389 931 1390
rect 935 1394 939 1395
rect 935 1389 939 1390
rect 1015 1394 1019 1395
rect 1015 1389 1019 1390
rect 1039 1394 1043 1395
rect 1039 1389 1043 1390
rect 1103 1394 1107 1395
rect 1103 1389 1107 1390
rect 1143 1394 1147 1395
rect 1143 1389 1147 1390
rect 1199 1394 1203 1395
rect 1199 1389 1203 1390
rect 1239 1394 1243 1395
rect 1239 1389 1243 1390
rect 928 1370 930 1389
rect 1016 1370 1018 1389
rect 1104 1370 1106 1389
rect 1200 1370 1202 1389
rect 1248 1388 1250 1418
rect 1288 1395 1290 1419
rect 1328 1399 1330 1419
rect 1374 1418 1380 1419
rect 1442 1423 1448 1424
rect 1442 1419 1443 1423
rect 1447 1419 1448 1423
rect 1442 1418 1448 1419
rect 1462 1423 1468 1424
rect 1462 1419 1463 1423
rect 1467 1419 1468 1423
rect 1462 1418 1468 1419
rect 1530 1423 1536 1424
rect 1530 1419 1531 1423
rect 1535 1419 1536 1423
rect 1530 1418 1536 1419
rect 1550 1423 1556 1424
rect 1550 1419 1551 1423
rect 1555 1419 1556 1423
rect 1550 1418 1556 1419
rect 1566 1423 1572 1424
rect 1566 1419 1567 1423
rect 1571 1419 1572 1423
rect 1566 1418 1572 1419
rect 1646 1423 1652 1424
rect 1646 1419 1647 1423
rect 1651 1419 1652 1423
rect 1646 1418 1652 1419
rect 1742 1423 1748 1424
rect 1742 1419 1743 1423
rect 1747 1419 1748 1423
rect 1742 1418 1748 1419
rect 1376 1399 1378 1418
rect 1444 1404 1446 1418
rect 1442 1403 1448 1404
rect 1442 1399 1443 1403
rect 1447 1399 1448 1403
rect 1464 1399 1466 1418
rect 1532 1404 1534 1418
rect 1530 1403 1536 1404
rect 1530 1399 1531 1403
rect 1535 1399 1536 1403
rect 1552 1399 1554 1418
rect 1648 1399 1650 1418
rect 1744 1399 1746 1418
rect 1824 1404 1826 1486
rect 1870 1485 1876 1486
rect 1870 1481 1871 1485
rect 1875 1481 1876 1485
rect 1896 1484 1898 1498
rect 1952 1486 1954 1505
rect 1974 1503 1980 1504
rect 1974 1499 1975 1503
rect 1979 1499 1980 1503
rect 1974 1498 1980 1499
rect 1950 1485 1956 1486
rect 1870 1480 1876 1481
rect 1894 1483 1900 1484
rect 1894 1479 1895 1483
rect 1899 1479 1900 1483
rect 1950 1481 1951 1485
rect 1955 1481 1956 1485
rect 1976 1484 1978 1498
rect 2032 1486 2034 1505
rect 2054 1503 2060 1504
rect 2054 1499 2055 1503
rect 2059 1499 2060 1503
rect 2054 1498 2060 1499
rect 2030 1485 2036 1486
rect 1950 1480 1956 1481
rect 1974 1483 1980 1484
rect 1894 1478 1900 1479
rect 1974 1479 1975 1483
rect 1979 1479 1980 1483
rect 2030 1481 2031 1485
rect 2035 1481 2036 1485
rect 2056 1484 2058 1498
rect 2120 1486 2122 1505
rect 2118 1485 2124 1486
rect 2504 1485 2506 1505
rect 2030 1480 2036 1481
rect 2054 1483 2060 1484
rect 1974 1478 1980 1479
rect 2054 1479 2055 1483
rect 2059 1479 2060 1483
rect 2118 1481 2119 1485
rect 2123 1481 2124 1485
rect 2118 1480 2124 1481
rect 2502 1484 2508 1485
rect 2502 1480 2503 1484
rect 2507 1480 2508 1484
rect 2502 1479 2508 1480
rect 2054 1478 2060 1479
rect 2502 1467 2508 1468
rect 1854 1464 1860 1465
rect 1854 1460 1855 1464
rect 1859 1460 1860 1464
rect 1854 1459 1860 1460
rect 1934 1464 1940 1465
rect 1934 1460 1935 1464
rect 1939 1460 1940 1464
rect 1934 1459 1940 1460
rect 2014 1464 2020 1465
rect 2014 1460 2015 1464
rect 2019 1460 2020 1464
rect 2014 1459 2020 1460
rect 2102 1464 2108 1465
rect 2102 1460 2103 1464
rect 2107 1460 2108 1464
rect 2502 1463 2503 1467
rect 2507 1463 2508 1467
rect 2502 1462 2508 1463
rect 2102 1459 2108 1460
rect 1856 1451 1858 1459
rect 1936 1451 1938 1459
rect 2016 1451 2018 1459
rect 2104 1451 2106 1459
rect 2504 1451 2506 1462
rect 1855 1450 1859 1451
rect 1855 1445 1859 1446
rect 1903 1450 1907 1451
rect 1903 1445 1907 1446
rect 1935 1450 1939 1451
rect 1935 1445 1939 1446
rect 1991 1450 1995 1451
rect 1991 1445 1995 1446
rect 2015 1450 2019 1451
rect 2015 1445 2019 1446
rect 2071 1450 2075 1451
rect 2071 1445 2075 1446
rect 2103 1450 2107 1451
rect 2103 1445 2107 1446
rect 2159 1450 2163 1451
rect 2159 1445 2163 1446
rect 2247 1450 2251 1451
rect 2247 1445 2251 1446
rect 2503 1450 2507 1451
rect 2503 1445 2507 1446
rect 1902 1444 1908 1445
rect 1902 1440 1903 1444
rect 1907 1440 1908 1444
rect 1902 1439 1908 1440
rect 1990 1444 1996 1445
rect 1990 1440 1991 1444
rect 1995 1440 1996 1444
rect 1990 1439 1996 1440
rect 2070 1444 2076 1445
rect 2070 1440 2071 1444
rect 2075 1440 2076 1444
rect 2070 1439 2076 1440
rect 2158 1444 2164 1445
rect 2158 1440 2159 1444
rect 2163 1440 2164 1444
rect 2158 1439 2164 1440
rect 2246 1444 2252 1445
rect 2246 1440 2247 1444
rect 2251 1440 2252 1444
rect 2504 1442 2506 1445
rect 2246 1439 2252 1440
rect 2502 1441 2508 1442
rect 2502 1437 2503 1441
rect 2507 1437 2508 1441
rect 2502 1436 2508 1437
rect 2502 1424 2508 1425
rect 1830 1423 1836 1424
rect 1830 1419 1831 1423
rect 1835 1419 1836 1423
rect 1830 1418 1836 1419
rect 1898 1423 1904 1424
rect 1898 1419 1899 1423
rect 1903 1419 1904 1423
rect 1898 1418 1904 1419
rect 1918 1423 1924 1424
rect 1918 1419 1919 1423
rect 1923 1419 1924 1423
rect 1918 1418 1924 1419
rect 1986 1423 1992 1424
rect 1986 1419 1987 1423
rect 1991 1419 1992 1423
rect 1986 1418 1992 1419
rect 2006 1423 2012 1424
rect 2006 1419 2007 1423
rect 2011 1419 2012 1423
rect 2006 1418 2012 1419
rect 2066 1423 2072 1424
rect 2066 1419 2067 1423
rect 2071 1419 2072 1423
rect 2066 1418 2072 1419
rect 2086 1423 2092 1424
rect 2086 1419 2087 1423
rect 2091 1419 2092 1423
rect 2086 1418 2092 1419
rect 2154 1423 2160 1424
rect 2154 1419 2155 1423
rect 2159 1419 2160 1423
rect 2154 1418 2160 1419
rect 2174 1423 2180 1424
rect 2174 1419 2175 1423
rect 2179 1419 2180 1423
rect 2174 1418 2180 1419
rect 2238 1423 2244 1424
rect 2238 1419 2239 1423
rect 2243 1419 2244 1423
rect 2238 1418 2244 1419
rect 2262 1423 2268 1424
rect 2262 1419 2263 1423
rect 2267 1419 2268 1423
rect 2502 1420 2503 1424
rect 2507 1420 2508 1424
rect 2502 1419 2508 1420
rect 2262 1418 2268 1419
rect 1754 1403 1760 1404
rect 1754 1399 1755 1403
rect 1759 1399 1760 1403
rect 1327 1398 1331 1399
rect 1287 1394 1291 1395
rect 1327 1393 1331 1394
rect 1375 1398 1379 1399
rect 1442 1398 1448 1399
rect 1463 1398 1467 1399
rect 1530 1398 1536 1399
rect 1551 1398 1555 1399
rect 1375 1393 1379 1394
rect 1463 1393 1467 1394
rect 1551 1393 1555 1394
rect 1567 1398 1571 1399
rect 1567 1393 1571 1394
rect 1647 1398 1651 1399
rect 1647 1393 1651 1394
rect 1735 1398 1739 1399
rect 1735 1393 1739 1394
rect 1743 1398 1747 1399
rect 1754 1398 1760 1399
rect 1822 1403 1828 1404
rect 1822 1399 1823 1403
rect 1827 1399 1828 1403
rect 1832 1399 1834 1418
rect 1900 1404 1902 1418
rect 1898 1403 1904 1404
rect 1898 1399 1899 1403
rect 1903 1399 1904 1403
rect 1920 1399 1922 1418
rect 1988 1404 1990 1418
rect 1994 1415 2000 1416
rect 1994 1411 1995 1415
rect 1999 1411 2000 1415
rect 1994 1410 2000 1411
rect 1986 1403 1992 1404
rect 1986 1399 1987 1403
rect 1991 1399 1992 1403
rect 1822 1398 1828 1399
rect 1831 1398 1835 1399
rect 1898 1398 1904 1399
rect 1919 1398 1923 1399
rect 1986 1398 1992 1399
rect 1743 1393 1747 1394
rect 1287 1389 1291 1390
rect 1246 1387 1252 1388
rect 1246 1383 1247 1387
rect 1251 1383 1252 1387
rect 1246 1382 1252 1383
rect 926 1369 932 1370
rect 838 1364 844 1365
rect 858 1367 864 1368
rect 774 1362 780 1363
rect 858 1363 859 1367
rect 863 1363 864 1367
rect 926 1365 927 1369
rect 931 1365 932 1369
rect 1014 1369 1020 1370
rect 926 1364 932 1365
rect 966 1367 972 1368
rect 858 1362 864 1363
rect 966 1363 967 1367
rect 971 1363 972 1367
rect 1014 1365 1015 1369
rect 1019 1365 1020 1369
rect 1014 1364 1020 1365
rect 1102 1369 1108 1370
rect 1102 1365 1103 1369
rect 1107 1365 1108 1369
rect 1102 1364 1108 1365
rect 1198 1369 1204 1370
rect 1288 1369 1290 1389
rect 1328 1373 1330 1393
rect 1568 1374 1570 1393
rect 1590 1391 1596 1392
rect 1590 1387 1591 1391
rect 1595 1387 1596 1391
rect 1590 1386 1596 1387
rect 1566 1373 1572 1374
rect 1326 1372 1332 1373
rect 1198 1365 1199 1369
rect 1203 1365 1204 1369
rect 1198 1364 1204 1365
rect 1286 1368 1292 1369
rect 1286 1364 1287 1368
rect 1291 1364 1292 1368
rect 1326 1368 1327 1372
rect 1331 1368 1332 1372
rect 1566 1369 1567 1373
rect 1571 1369 1572 1373
rect 1592 1372 1594 1386
rect 1648 1374 1650 1393
rect 1670 1391 1676 1392
rect 1670 1387 1671 1391
rect 1675 1387 1676 1391
rect 1670 1386 1676 1387
rect 1646 1373 1652 1374
rect 1566 1368 1572 1369
rect 1590 1371 1596 1372
rect 1326 1367 1332 1368
rect 1590 1367 1591 1371
rect 1595 1367 1596 1371
rect 1646 1369 1647 1373
rect 1651 1369 1652 1373
rect 1672 1372 1674 1386
rect 1736 1374 1738 1393
rect 1734 1373 1740 1374
rect 1646 1368 1652 1369
rect 1670 1371 1676 1372
rect 1590 1366 1596 1367
rect 1670 1367 1671 1371
rect 1675 1367 1676 1371
rect 1734 1369 1735 1373
rect 1739 1369 1740 1373
rect 1756 1372 1758 1398
rect 1831 1393 1835 1394
rect 1919 1393 1923 1394
rect 1832 1374 1834 1393
rect 1920 1374 1922 1393
rect 1996 1392 1998 1410
rect 2008 1399 2010 1418
rect 2068 1404 2070 1418
rect 2066 1403 2072 1404
rect 2066 1399 2067 1403
rect 2071 1399 2072 1403
rect 2088 1399 2090 1418
rect 2156 1404 2158 1418
rect 2154 1403 2160 1404
rect 2154 1399 2155 1403
rect 2159 1399 2160 1403
rect 2176 1399 2178 1418
rect 2240 1404 2242 1418
rect 2238 1403 2244 1404
rect 2238 1399 2239 1403
rect 2243 1399 2244 1403
rect 2264 1399 2266 1418
rect 2504 1399 2506 1419
rect 2007 1398 2011 1399
rect 2066 1398 2072 1399
rect 2087 1398 2091 1399
rect 2007 1393 2011 1394
rect 2087 1393 2091 1394
rect 2095 1398 2099 1399
rect 2154 1398 2160 1399
rect 2175 1398 2179 1399
rect 2238 1398 2244 1399
rect 2247 1398 2251 1399
rect 2095 1393 2099 1394
rect 2175 1393 2179 1394
rect 2247 1393 2251 1394
rect 2263 1398 2267 1399
rect 2263 1393 2267 1394
rect 2319 1398 2323 1399
rect 2319 1393 2323 1394
rect 2399 1398 2403 1399
rect 2399 1393 2403 1394
rect 2455 1398 2459 1399
rect 2455 1393 2459 1394
rect 2503 1398 2507 1399
rect 2503 1393 2507 1394
rect 1930 1391 1936 1392
rect 1930 1387 1931 1391
rect 1935 1387 1936 1391
rect 1930 1386 1936 1387
rect 1990 1391 1998 1392
rect 1990 1387 1991 1391
rect 1995 1388 1998 1391
rect 1995 1387 1996 1388
rect 1990 1386 1996 1387
rect 1830 1373 1836 1374
rect 1734 1368 1740 1369
rect 1754 1371 1760 1372
rect 1670 1366 1676 1367
rect 1754 1367 1755 1371
rect 1759 1367 1760 1371
rect 1830 1369 1831 1373
rect 1835 1369 1836 1373
rect 1830 1368 1836 1369
rect 1918 1373 1924 1374
rect 1918 1369 1919 1373
rect 1923 1369 1924 1373
rect 1918 1368 1924 1369
rect 1754 1366 1760 1367
rect 1286 1363 1292 1364
rect 966 1362 972 1363
rect 734 1348 740 1349
rect 734 1344 735 1348
rect 739 1344 740 1348
rect 734 1343 740 1344
rect 822 1348 828 1349
rect 822 1344 823 1348
rect 827 1344 828 1348
rect 822 1343 828 1344
rect 910 1348 916 1349
rect 910 1344 911 1348
rect 915 1344 916 1348
rect 910 1343 916 1344
rect 736 1327 738 1343
rect 824 1327 826 1343
rect 912 1327 914 1343
rect 687 1326 691 1327
rect 687 1321 691 1322
rect 735 1326 739 1327
rect 735 1321 739 1322
rect 783 1326 787 1327
rect 783 1321 787 1322
rect 823 1326 827 1327
rect 823 1321 827 1322
rect 879 1326 883 1327
rect 879 1321 883 1322
rect 911 1326 915 1327
rect 911 1321 915 1322
rect 686 1320 692 1321
rect 686 1316 687 1320
rect 691 1316 692 1320
rect 686 1315 692 1316
rect 782 1320 788 1321
rect 782 1316 783 1320
rect 787 1316 788 1320
rect 782 1315 788 1316
rect 878 1320 884 1321
rect 878 1316 879 1320
rect 883 1316 884 1320
rect 878 1315 884 1316
rect 254 1299 260 1300
rect 254 1295 255 1299
rect 259 1295 260 1299
rect 254 1294 260 1295
rect 362 1299 368 1300
rect 362 1295 363 1299
rect 367 1295 368 1299
rect 362 1294 368 1295
rect 382 1299 388 1300
rect 382 1295 383 1299
rect 387 1295 388 1299
rect 382 1294 388 1295
rect 494 1299 500 1300
rect 494 1295 495 1299
rect 499 1295 500 1299
rect 494 1294 500 1295
rect 578 1299 584 1300
rect 578 1295 579 1299
rect 583 1295 584 1299
rect 578 1294 584 1295
rect 598 1299 604 1300
rect 598 1295 599 1299
rect 603 1295 604 1299
rect 598 1294 604 1295
rect 654 1299 660 1300
rect 654 1295 655 1299
rect 659 1295 660 1299
rect 654 1294 660 1295
rect 702 1299 708 1300
rect 702 1295 703 1299
rect 707 1295 708 1299
rect 702 1294 708 1295
rect 746 1299 752 1300
rect 746 1295 747 1299
rect 751 1295 752 1299
rect 746 1294 752 1295
rect 798 1299 804 1300
rect 798 1295 799 1299
rect 803 1295 804 1299
rect 798 1294 804 1295
rect 806 1299 812 1300
rect 806 1295 807 1299
rect 811 1295 812 1299
rect 806 1294 812 1295
rect 894 1299 900 1300
rect 894 1295 895 1299
rect 899 1295 900 1299
rect 894 1294 900 1295
rect 246 1279 252 1280
rect 246 1275 247 1279
rect 251 1275 252 1279
rect 246 1274 252 1275
rect 256 1267 258 1294
rect 364 1280 366 1294
rect 362 1279 368 1280
rect 362 1275 363 1279
rect 367 1275 368 1279
rect 362 1274 368 1275
rect 384 1267 386 1294
rect 496 1267 498 1294
rect 580 1280 582 1294
rect 570 1279 576 1280
rect 570 1275 571 1279
rect 575 1275 576 1279
rect 570 1274 576 1275
rect 578 1279 584 1280
rect 578 1275 579 1279
rect 583 1275 584 1279
rect 578 1274 584 1275
rect 215 1266 219 1267
rect 215 1261 219 1262
rect 255 1266 259 1267
rect 255 1261 259 1262
rect 303 1266 307 1267
rect 303 1261 307 1262
rect 383 1266 387 1267
rect 383 1261 387 1262
rect 391 1266 395 1267
rect 391 1261 395 1262
rect 471 1266 475 1267
rect 471 1261 475 1262
rect 495 1266 499 1267
rect 495 1261 499 1262
rect 551 1266 555 1267
rect 551 1261 555 1262
rect 158 1259 164 1260
rect 158 1255 159 1259
rect 163 1255 164 1259
rect 158 1254 164 1255
rect 216 1242 218 1261
rect 238 1259 244 1260
rect 238 1255 239 1259
rect 243 1255 244 1259
rect 238 1254 244 1255
rect 150 1241 156 1242
rect 110 1240 116 1241
rect 110 1236 111 1240
rect 115 1236 116 1240
rect 150 1237 151 1241
rect 155 1237 156 1241
rect 150 1236 156 1237
rect 214 1241 220 1242
rect 214 1237 215 1241
rect 219 1237 220 1241
rect 240 1240 242 1254
rect 304 1242 306 1261
rect 326 1259 332 1260
rect 326 1255 327 1259
rect 331 1255 332 1259
rect 326 1254 332 1255
rect 302 1241 308 1242
rect 214 1236 220 1237
rect 238 1239 244 1240
rect 110 1235 116 1236
rect 238 1235 239 1239
rect 243 1235 244 1239
rect 302 1237 303 1241
rect 307 1237 308 1241
rect 328 1240 330 1254
rect 392 1242 394 1261
rect 462 1259 468 1260
rect 462 1255 463 1259
rect 467 1255 468 1259
rect 462 1254 468 1255
rect 390 1241 396 1242
rect 302 1236 308 1237
rect 326 1239 332 1240
rect 238 1234 244 1235
rect 326 1235 327 1239
rect 331 1235 332 1239
rect 390 1237 391 1241
rect 395 1237 396 1241
rect 390 1236 396 1237
rect 398 1239 404 1240
rect 326 1234 332 1235
rect 398 1235 399 1239
rect 403 1235 404 1239
rect 398 1234 404 1235
rect 110 1223 116 1224
rect 110 1219 111 1223
rect 115 1219 116 1223
rect 110 1218 116 1219
rect 134 1220 140 1221
rect 112 1211 114 1218
rect 134 1216 135 1220
rect 139 1216 140 1220
rect 134 1215 140 1216
rect 198 1220 204 1221
rect 198 1216 199 1220
rect 203 1216 204 1220
rect 198 1215 204 1216
rect 286 1220 292 1221
rect 286 1216 287 1220
rect 291 1216 292 1220
rect 286 1215 292 1216
rect 374 1220 380 1221
rect 374 1216 375 1220
rect 379 1216 380 1220
rect 374 1215 380 1216
rect 136 1211 138 1215
rect 200 1211 202 1215
rect 288 1211 290 1215
rect 376 1211 378 1215
rect 111 1210 115 1211
rect 111 1205 115 1206
rect 135 1210 139 1211
rect 135 1205 139 1206
rect 191 1210 195 1211
rect 191 1205 195 1206
rect 199 1210 203 1211
rect 199 1205 203 1206
rect 271 1210 275 1211
rect 271 1205 275 1206
rect 287 1210 291 1211
rect 287 1205 291 1206
rect 351 1210 355 1211
rect 351 1205 355 1206
rect 375 1210 379 1211
rect 375 1205 379 1206
rect 112 1202 114 1205
rect 134 1204 140 1205
rect 110 1201 116 1202
rect 110 1197 111 1201
rect 115 1197 116 1201
rect 134 1200 135 1204
rect 139 1200 140 1204
rect 134 1199 140 1200
rect 190 1204 196 1205
rect 190 1200 191 1204
rect 195 1200 196 1204
rect 190 1199 196 1200
rect 270 1204 276 1205
rect 270 1200 271 1204
rect 275 1200 276 1204
rect 270 1199 276 1200
rect 350 1204 356 1205
rect 350 1200 351 1204
rect 355 1200 356 1204
rect 350 1199 356 1200
rect 110 1196 116 1197
rect 110 1184 116 1185
rect 110 1180 111 1184
rect 115 1180 116 1184
rect 110 1179 116 1180
rect 150 1183 156 1184
rect 150 1179 151 1183
rect 155 1179 156 1183
rect 112 1155 114 1179
rect 150 1178 156 1179
rect 186 1183 192 1184
rect 186 1179 187 1183
rect 191 1179 192 1183
rect 186 1178 192 1179
rect 206 1183 212 1184
rect 206 1179 207 1183
rect 211 1179 212 1183
rect 206 1178 212 1179
rect 266 1183 272 1184
rect 266 1179 267 1183
rect 271 1179 272 1183
rect 266 1178 272 1179
rect 286 1183 292 1184
rect 286 1179 287 1183
rect 291 1179 292 1183
rect 286 1178 292 1179
rect 346 1183 352 1184
rect 346 1179 347 1183
rect 351 1179 352 1183
rect 346 1178 352 1179
rect 366 1183 372 1184
rect 366 1179 367 1183
rect 371 1179 372 1183
rect 366 1178 372 1179
rect 382 1183 388 1184
rect 382 1179 383 1183
rect 387 1179 388 1183
rect 382 1178 388 1179
rect 152 1155 154 1178
rect 188 1164 190 1178
rect 186 1163 192 1164
rect 186 1159 187 1163
rect 191 1159 192 1163
rect 186 1158 192 1159
rect 208 1155 210 1178
rect 268 1164 270 1178
rect 266 1163 272 1164
rect 266 1159 267 1163
rect 271 1159 272 1163
rect 266 1158 272 1159
rect 288 1155 290 1178
rect 348 1164 350 1178
rect 346 1163 352 1164
rect 346 1159 347 1163
rect 351 1159 352 1163
rect 346 1158 352 1159
rect 368 1155 370 1178
rect 111 1154 115 1155
rect 111 1149 115 1150
rect 151 1154 155 1155
rect 151 1149 155 1150
rect 183 1154 187 1155
rect 183 1149 187 1150
rect 207 1154 211 1155
rect 207 1149 211 1150
rect 279 1154 283 1155
rect 279 1149 283 1150
rect 287 1154 291 1155
rect 287 1149 291 1150
rect 367 1154 371 1155
rect 367 1149 371 1150
rect 375 1154 379 1155
rect 375 1149 379 1150
rect 112 1129 114 1149
rect 184 1130 186 1149
rect 280 1130 282 1149
rect 376 1130 378 1149
rect 384 1148 386 1178
rect 400 1172 402 1234
rect 454 1220 460 1221
rect 454 1216 455 1220
rect 459 1216 460 1220
rect 454 1215 460 1216
rect 456 1211 458 1215
rect 431 1210 435 1211
rect 431 1205 435 1206
rect 455 1210 459 1211
rect 455 1205 459 1206
rect 430 1204 436 1205
rect 430 1200 431 1204
rect 435 1200 436 1204
rect 430 1199 436 1200
rect 464 1184 466 1254
rect 472 1242 474 1261
rect 502 1259 508 1260
rect 502 1255 503 1259
rect 507 1255 508 1259
rect 502 1254 508 1255
rect 470 1241 476 1242
rect 470 1237 471 1241
rect 475 1237 476 1241
rect 504 1240 506 1254
rect 552 1242 554 1261
rect 550 1241 556 1242
rect 470 1236 476 1237
rect 502 1239 508 1240
rect 502 1235 503 1239
rect 507 1235 508 1239
rect 550 1237 551 1241
rect 555 1237 556 1241
rect 572 1240 574 1274
rect 600 1267 602 1294
rect 704 1267 706 1294
rect 599 1266 603 1267
rect 599 1261 603 1262
rect 623 1266 627 1267
rect 623 1261 627 1262
rect 695 1266 699 1267
rect 695 1261 699 1262
rect 703 1266 707 1267
rect 703 1261 707 1262
rect 624 1242 626 1261
rect 696 1242 698 1261
rect 748 1260 750 1294
rect 800 1267 802 1294
rect 808 1276 810 1294
rect 806 1275 812 1276
rect 806 1271 807 1275
rect 811 1271 812 1275
rect 806 1270 812 1271
rect 896 1267 898 1294
rect 968 1280 970 1362
rect 1326 1355 1332 1356
rect 1286 1351 1292 1352
rect 998 1348 1004 1349
rect 998 1344 999 1348
rect 1003 1344 1004 1348
rect 998 1343 1004 1344
rect 1086 1348 1092 1349
rect 1086 1344 1087 1348
rect 1091 1344 1092 1348
rect 1086 1343 1092 1344
rect 1182 1348 1188 1349
rect 1182 1344 1183 1348
rect 1187 1344 1188 1348
rect 1286 1347 1287 1351
rect 1291 1347 1292 1351
rect 1326 1351 1327 1355
rect 1331 1351 1332 1355
rect 1326 1350 1332 1351
rect 1550 1352 1556 1353
rect 1328 1347 1330 1350
rect 1550 1348 1551 1352
rect 1555 1348 1556 1352
rect 1550 1347 1556 1348
rect 1630 1352 1636 1353
rect 1630 1348 1631 1352
rect 1635 1348 1636 1352
rect 1630 1347 1636 1348
rect 1718 1352 1724 1353
rect 1718 1348 1719 1352
rect 1723 1348 1724 1352
rect 1718 1347 1724 1348
rect 1814 1352 1820 1353
rect 1814 1348 1815 1352
rect 1819 1348 1820 1352
rect 1814 1347 1820 1348
rect 1902 1352 1908 1353
rect 1902 1348 1903 1352
rect 1907 1348 1908 1352
rect 1902 1347 1908 1348
rect 1286 1346 1292 1347
rect 1327 1346 1331 1347
rect 1182 1343 1188 1344
rect 1000 1327 1002 1343
rect 1088 1327 1090 1343
rect 1184 1327 1186 1343
rect 1288 1327 1290 1346
rect 1327 1341 1331 1342
rect 1551 1346 1555 1347
rect 1551 1341 1555 1342
rect 1583 1346 1587 1347
rect 1583 1341 1587 1342
rect 1631 1346 1635 1347
rect 1631 1341 1635 1342
rect 1647 1346 1651 1347
rect 1647 1341 1651 1342
rect 1719 1346 1723 1347
rect 1719 1341 1723 1342
rect 1727 1346 1731 1347
rect 1727 1341 1731 1342
rect 1807 1346 1811 1347
rect 1807 1341 1811 1342
rect 1815 1346 1819 1347
rect 1815 1341 1819 1342
rect 1895 1346 1899 1347
rect 1895 1341 1899 1342
rect 1903 1346 1907 1347
rect 1903 1341 1907 1342
rect 1328 1338 1330 1341
rect 1582 1340 1588 1341
rect 1326 1337 1332 1338
rect 1326 1333 1327 1337
rect 1331 1333 1332 1337
rect 1582 1336 1583 1340
rect 1587 1336 1588 1340
rect 1582 1335 1588 1336
rect 1646 1340 1652 1341
rect 1646 1336 1647 1340
rect 1651 1336 1652 1340
rect 1646 1335 1652 1336
rect 1726 1340 1732 1341
rect 1726 1336 1727 1340
rect 1731 1336 1732 1340
rect 1726 1335 1732 1336
rect 1806 1340 1812 1341
rect 1806 1336 1807 1340
rect 1811 1336 1812 1340
rect 1806 1335 1812 1336
rect 1894 1340 1900 1341
rect 1894 1336 1895 1340
rect 1899 1336 1900 1340
rect 1894 1335 1900 1336
rect 1326 1332 1332 1333
rect 975 1326 979 1327
rect 975 1321 979 1322
rect 999 1326 1003 1327
rect 999 1321 1003 1322
rect 1087 1326 1091 1327
rect 1087 1321 1091 1322
rect 1183 1326 1187 1327
rect 1183 1321 1187 1322
rect 1287 1326 1291 1327
rect 1287 1321 1291 1322
rect 974 1320 980 1321
rect 974 1316 975 1320
rect 979 1316 980 1320
rect 1288 1318 1290 1321
rect 1326 1320 1332 1321
rect 1932 1320 1934 1386
rect 2008 1374 2010 1393
rect 2030 1391 2036 1392
rect 2030 1387 2031 1391
rect 2035 1387 2036 1391
rect 2030 1386 2036 1387
rect 2006 1373 2012 1374
rect 2006 1369 2007 1373
rect 2011 1369 2012 1373
rect 2032 1372 2034 1386
rect 2096 1374 2098 1393
rect 2118 1391 2124 1392
rect 2118 1387 2119 1391
rect 2123 1387 2124 1391
rect 2118 1386 2124 1387
rect 2094 1373 2100 1374
rect 2006 1368 2012 1369
rect 2030 1371 2036 1372
rect 2030 1367 2031 1371
rect 2035 1367 2036 1371
rect 2094 1369 2095 1373
rect 2099 1369 2100 1373
rect 2120 1372 2122 1386
rect 2176 1374 2178 1393
rect 2214 1391 2220 1392
rect 2214 1387 2215 1391
rect 2219 1387 2220 1391
rect 2214 1386 2220 1387
rect 2174 1373 2180 1374
rect 2094 1368 2100 1369
rect 2118 1371 2124 1372
rect 2030 1366 2036 1367
rect 2118 1367 2119 1371
rect 2123 1367 2124 1371
rect 2174 1369 2175 1373
rect 2179 1369 2180 1373
rect 2216 1372 2218 1386
rect 2248 1374 2250 1393
rect 2270 1391 2276 1392
rect 2270 1387 2271 1391
rect 2275 1387 2276 1391
rect 2270 1386 2276 1387
rect 2246 1373 2252 1374
rect 2174 1368 2180 1369
rect 2214 1371 2220 1372
rect 2118 1366 2124 1367
rect 2214 1367 2215 1371
rect 2219 1367 2220 1371
rect 2246 1369 2247 1373
rect 2251 1369 2252 1373
rect 2272 1372 2274 1386
rect 2320 1374 2322 1393
rect 2400 1374 2402 1393
rect 2414 1391 2420 1392
rect 2414 1387 2415 1391
rect 2419 1387 2420 1391
rect 2414 1386 2420 1387
rect 2422 1391 2428 1392
rect 2422 1387 2423 1391
rect 2427 1387 2428 1391
rect 2422 1386 2428 1387
rect 2318 1373 2324 1374
rect 2246 1368 2252 1369
rect 2270 1371 2276 1372
rect 2214 1366 2220 1367
rect 2270 1367 2271 1371
rect 2275 1367 2276 1371
rect 2318 1369 2319 1373
rect 2323 1369 2324 1373
rect 2398 1373 2404 1374
rect 2318 1368 2324 1369
rect 2326 1371 2332 1372
rect 2270 1366 2276 1367
rect 2326 1367 2327 1371
rect 2331 1367 2332 1371
rect 2398 1369 2399 1373
rect 2403 1369 2404 1373
rect 2398 1368 2404 1369
rect 2326 1366 2332 1367
rect 1990 1352 1996 1353
rect 1990 1348 1991 1352
rect 1995 1348 1996 1352
rect 1990 1347 1996 1348
rect 2078 1352 2084 1353
rect 2078 1348 2079 1352
rect 2083 1348 2084 1352
rect 2078 1347 2084 1348
rect 2158 1352 2164 1353
rect 2158 1348 2159 1352
rect 2163 1348 2164 1352
rect 2158 1347 2164 1348
rect 2230 1352 2236 1353
rect 2230 1348 2231 1352
rect 2235 1348 2236 1352
rect 2230 1347 2236 1348
rect 2302 1352 2308 1353
rect 2302 1348 2303 1352
rect 2307 1348 2308 1352
rect 2302 1347 2308 1348
rect 1983 1346 1987 1347
rect 1983 1341 1987 1342
rect 1991 1346 1995 1347
rect 1991 1341 1995 1342
rect 2063 1346 2067 1347
rect 2063 1341 2067 1342
rect 2079 1346 2083 1347
rect 2079 1341 2083 1342
rect 2143 1346 2147 1347
rect 2143 1341 2147 1342
rect 2159 1346 2163 1347
rect 2159 1341 2163 1342
rect 2223 1346 2227 1347
rect 2223 1341 2227 1342
rect 2231 1346 2235 1347
rect 2231 1341 2235 1342
rect 2303 1346 2307 1347
rect 2303 1341 2307 1342
rect 1982 1340 1988 1341
rect 1982 1336 1983 1340
rect 1987 1336 1988 1340
rect 1982 1335 1988 1336
rect 2062 1340 2068 1341
rect 2062 1336 2063 1340
rect 2067 1336 2068 1340
rect 2062 1335 2068 1336
rect 2142 1340 2148 1341
rect 2142 1336 2143 1340
rect 2147 1336 2148 1340
rect 2142 1335 2148 1336
rect 2222 1340 2228 1341
rect 2222 1336 2223 1340
rect 2227 1336 2228 1340
rect 2222 1335 2228 1336
rect 2302 1340 2308 1341
rect 2302 1336 2303 1340
rect 2307 1336 2308 1340
rect 2302 1335 2308 1336
rect 974 1315 980 1316
rect 1286 1317 1292 1318
rect 1286 1313 1287 1317
rect 1291 1313 1292 1317
rect 1326 1316 1327 1320
rect 1331 1316 1332 1320
rect 1326 1315 1332 1316
rect 1598 1319 1604 1320
rect 1598 1315 1599 1319
rect 1603 1315 1604 1319
rect 1286 1312 1292 1313
rect 1286 1300 1292 1301
rect 990 1299 996 1300
rect 990 1295 991 1299
rect 995 1295 996 1299
rect 1286 1296 1287 1300
rect 1291 1296 1292 1300
rect 1286 1295 1292 1296
rect 1328 1295 1330 1315
rect 1598 1314 1604 1315
rect 1642 1319 1648 1320
rect 1642 1315 1643 1319
rect 1647 1315 1648 1319
rect 1642 1314 1648 1315
rect 1662 1319 1668 1320
rect 1662 1315 1663 1319
rect 1667 1315 1668 1319
rect 1662 1314 1668 1315
rect 1722 1319 1728 1320
rect 1722 1315 1723 1319
rect 1727 1315 1728 1319
rect 1722 1314 1728 1315
rect 1742 1319 1748 1320
rect 1742 1315 1743 1319
rect 1747 1315 1748 1319
rect 1742 1314 1748 1315
rect 1778 1319 1784 1320
rect 1778 1315 1779 1319
rect 1783 1315 1784 1319
rect 1778 1314 1784 1315
rect 1822 1319 1828 1320
rect 1822 1315 1823 1319
rect 1827 1315 1828 1319
rect 1822 1314 1828 1315
rect 1886 1319 1892 1320
rect 1886 1315 1887 1319
rect 1891 1315 1892 1319
rect 1886 1314 1892 1315
rect 1910 1319 1916 1320
rect 1910 1315 1911 1319
rect 1915 1315 1916 1319
rect 1910 1314 1916 1315
rect 1930 1319 1936 1320
rect 1930 1315 1931 1319
rect 1935 1315 1936 1319
rect 1930 1314 1936 1315
rect 1998 1319 2004 1320
rect 1998 1315 1999 1319
rect 2003 1315 2004 1319
rect 1998 1314 2004 1315
rect 2078 1319 2084 1320
rect 2078 1315 2079 1319
rect 2083 1315 2084 1319
rect 2078 1314 2084 1315
rect 2138 1319 2144 1320
rect 2138 1315 2139 1319
rect 2143 1315 2144 1319
rect 2138 1314 2144 1315
rect 2158 1319 2164 1320
rect 2158 1315 2159 1319
rect 2163 1315 2164 1319
rect 2158 1314 2164 1315
rect 2218 1319 2224 1320
rect 2218 1315 2219 1319
rect 2223 1315 2224 1319
rect 2218 1314 2224 1315
rect 2238 1319 2244 1320
rect 2238 1315 2239 1319
rect 2243 1315 2244 1319
rect 2238 1314 2244 1315
rect 2298 1319 2304 1320
rect 2298 1315 2299 1319
rect 2303 1315 2304 1319
rect 2298 1314 2304 1315
rect 2318 1319 2324 1320
rect 2318 1315 2319 1319
rect 2323 1315 2324 1319
rect 2318 1314 2324 1315
rect 1582 1299 1588 1300
rect 1582 1295 1583 1299
rect 1587 1295 1588 1299
rect 1600 1295 1602 1314
rect 1644 1300 1646 1314
rect 1642 1299 1648 1300
rect 1642 1295 1643 1299
rect 1647 1295 1648 1299
rect 1664 1295 1666 1314
rect 1724 1300 1726 1314
rect 1722 1299 1728 1300
rect 1722 1295 1723 1299
rect 1727 1295 1728 1299
rect 1744 1295 1746 1314
rect 990 1294 996 1295
rect 966 1279 972 1280
rect 966 1275 967 1279
rect 971 1275 972 1279
rect 966 1274 972 1275
rect 992 1267 994 1294
rect 1288 1267 1290 1295
rect 1327 1294 1331 1295
rect 1327 1289 1331 1290
rect 1567 1294 1571 1295
rect 1582 1294 1588 1295
rect 1599 1294 1603 1295
rect 1567 1289 1571 1290
rect 1328 1269 1330 1289
rect 1568 1270 1570 1289
rect 1566 1269 1572 1270
rect 1326 1268 1332 1269
rect 767 1266 771 1267
rect 767 1261 771 1262
rect 799 1266 803 1267
rect 799 1261 803 1262
rect 839 1266 843 1267
rect 839 1261 843 1262
rect 895 1266 899 1267
rect 895 1261 899 1262
rect 919 1266 923 1267
rect 919 1261 923 1262
rect 991 1266 995 1267
rect 991 1261 995 1262
rect 1287 1266 1291 1267
rect 1326 1264 1327 1268
rect 1331 1264 1332 1268
rect 1566 1265 1567 1269
rect 1571 1265 1572 1269
rect 1584 1268 1586 1294
rect 1599 1289 1603 1290
rect 1631 1294 1635 1295
rect 1642 1294 1648 1295
rect 1663 1294 1667 1295
rect 1631 1289 1635 1290
rect 1663 1289 1667 1290
rect 1711 1294 1715 1295
rect 1722 1294 1728 1295
rect 1743 1294 1747 1295
rect 1711 1289 1715 1290
rect 1743 1289 1747 1290
rect 1606 1287 1612 1288
rect 1606 1283 1607 1287
rect 1611 1283 1612 1287
rect 1606 1282 1612 1283
rect 1566 1264 1572 1265
rect 1582 1267 1588 1268
rect 1326 1263 1332 1264
rect 1582 1263 1583 1267
rect 1587 1263 1588 1267
rect 1582 1262 1588 1263
rect 1287 1261 1291 1262
rect 746 1259 752 1260
rect 746 1255 747 1259
rect 751 1255 752 1259
rect 746 1254 752 1255
rect 768 1242 770 1261
rect 790 1259 796 1260
rect 790 1255 791 1259
rect 795 1255 796 1259
rect 790 1254 796 1255
rect 622 1241 628 1242
rect 550 1236 556 1237
rect 570 1239 576 1240
rect 502 1234 508 1235
rect 570 1235 571 1239
rect 575 1235 576 1239
rect 622 1237 623 1241
rect 627 1237 628 1241
rect 694 1241 700 1242
rect 622 1236 628 1237
rect 630 1239 636 1240
rect 570 1234 576 1235
rect 630 1235 631 1239
rect 635 1235 636 1239
rect 694 1237 695 1241
rect 699 1237 700 1241
rect 694 1236 700 1237
rect 766 1241 772 1242
rect 766 1237 767 1241
rect 771 1237 772 1241
rect 792 1240 794 1254
rect 840 1242 842 1261
rect 862 1259 868 1260
rect 862 1255 863 1259
rect 867 1255 868 1259
rect 862 1254 868 1255
rect 838 1241 844 1242
rect 766 1236 772 1237
rect 790 1239 796 1240
rect 630 1234 636 1235
rect 790 1235 791 1239
rect 795 1235 796 1239
rect 838 1237 839 1241
rect 843 1237 844 1241
rect 864 1240 866 1254
rect 920 1242 922 1261
rect 918 1241 924 1242
rect 1288 1241 1290 1261
rect 1326 1251 1332 1252
rect 1326 1247 1327 1251
rect 1331 1247 1332 1251
rect 1326 1246 1332 1247
rect 1550 1248 1556 1249
rect 838 1236 844 1237
rect 862 1239 868 1240
rect 790 1234 796 1235
rect 862 1235 863 1239
rect 867 1235 868 1239
rect 918 1237 919 1241
rect 923 1237 924 1241
rect 918 1236 924 1237
rect 1286 1240 1292 1241
rect 1286 1236 1287 1240
rect 1291 1236 1292 1240
rect 1328 1239 1330 1246
rect 1550 1244 1551 1248
rect 1555 1244 1556 1248
rect 1550 1243 1556 1244
rect 1552 1239 1554 1243
rect 1286 1235 1292 1236
rect 1327 1238 1331 1239
rect 862 1234 868 1235
rect 534 1220 540 1221
rect 534 1216 535 1220
rect 539 1216 540 1220
rect 534 1215 540 1216
rect 606 1220 612 1221
rect 606 1216 607 1220
rect 611 1216 612 1220
rect 606 1215 612 1216
rect 536 1211 538 1215
rect 608 1211 610 1215
rect 511 1210 515 1211
rect 511 1205 515 1206
rect 535 1210 539 1211
rect 535 1205 539 1206
rect 583 1210 587 1211
rect 583 1205 587 1206
rect 607 1210 611 1211
rect 607 1205 611 1206
rect 510 1204 516 1205
rect 510 1200 511 1204
rect 515 1200 516 1204
rect 510 1199 516 1200
rect 582 1204 588 1205
rect 582 1200 583 1204
rect 587 1200 588 1204
rect 582 1199 588 1200
rect 446 1183 452 1184
rect 446 1179 447 1183
rect 451 1179 452 1183
rect 446 1178 452 1179
rect 462 1183 468 1184
rect 462 1179 463 1183
rect 467 1179 468 1183
rect 462 1178 468 1179
rect 526 1183 532 1184
rect 526 1179 527 1183
rect 531 1179 532 1183
rect 526 1178 532 1179
rect 598 1183 604 1184
rect 598 1179 599 1183
rect 603 1179 604 1183
rect 598 1178 604 1179
rect 398 1171 404 1172
rect 398 1167 399 1171
rect 403 1167 404 1171
rect 398 1166 404 1167
rect 448 1155 450 1178
rect 494 1163 500 1164
rect 494 1159 495 1163
rect 499 1159 500 1163
rect 494 1158 500 1159
rect 447 1154 451 1155
rect 447 1149 451 1150
rect 471 1154 475 1155
rect 471 1149 475 1150
rect 382 1147 388 1148
rect 382 1143 383 1147
rect 387 1143 388 1147
rect 382 1142 388 1143
rect 472 1130 474 1149
rect 182 1129 188 1130
rect 110 1128 116 1129
rect 110 1124 111 1128
rect 115 1124 116 1128
rect 182 1125 183 1129
rect 187 1125 188 1129
rect 278 1129 284 1130
rect 182 1124 188 1125
rect 198 1127 204 1128
rect 110 1123 116 1124
rect 198 1123 199 1127
rect 203 1123 204 1127
rect 278 1125 279 1129
rect 283 1125 284 1129
rect 278 1124 284 1125
rect 374 1129 380 1130
rect 374 1125 375 1129
rect 379 1125 380 1129
rect 374 1124 380 1125
rect 470 1129 476 1130
rect 470 1125 471 1129
rect 475 1125 476 1129
rect 496 1128 498 1158
rect 528 1155 530 1178
rect 600 1155 602 1178
rect 632 1164 634 1234
rect 1327 1233 1331 1234
rect 1519 1238 1523 1239
rect 1519 1233 1523 1234
rect 1551 1238 1555 1239
rect 1551 1233 1555 1234
rect 1575 1238 1579 1239
rect 1575 1233 1579 1234
rect 1328 1230 1330 1233
rect 1518 1232 1524 1233
rect 1326 1229 1332 1230
rect 1326 1225 1327 1229
rect 1331 1225 1332 1229
rect 1518 1228 1519 1232
rect 1523 1228 1524 1232
rect 1518 1227 1524 1228
rect 1574 1232 1580 1233
rect 1574 1228 1575 1232
rect 1579 1228 1580 1232
rect 1574 1227 1580 1228
rect 1326 1224 1332 1225
rect 1286 1223 1292 1224
rect 678 1220 684 1221
rect 678 1216 679 1220
rect 683 1216 684 1220
rect 678 1215 684 1216
rect 750 1220 756 1221
rect 750 1216 751 1220
rect 755 1216 756 1220
rect 750 1215 756 1216
rect 822 1220 828 1221
rect 822 1216 823 1220
rect 827 1216 828 1220
rect 822 1215 828 1216
rect 902 1220 908 1221
rect 902 1216 903 1220
rect 907 1216 908 1220
rect 1286 1219 1287 1223
rect 1291 1219 1292 1223
rect 1286 1218 1292 1219
rect 902 1215 908 1216
rect 680 1211 682 1215
rect 752 1211 754 1215
rect 824 1211 826 1215
rect 904 1211 906 1215
rect 1288 1211 1290 1218
rect 1326 1212 1332 1213
rect 1608 1212 1610 1282
rect 1632 1270 1634 1289
rect 1712 1270 1714 1289
rect 1780 1288 1782 1314
rect 1824 1295 1826 1314
rect 1888 1300 1890 1314
rect 1886 1299 1892 1300
rect 1886 1295 1887 1299
rect 1891 1295 1892 1299
rect 1912 1295 1914 1314
rect 2000 1295 2002 1314
rect 2010 1299 2016 1300
rect 2010 1295 2011 1299
rect 2015 1295 2016 1299
rect 2080 1295 2082 1314
rect 2140 1300 2142 1314
rect 2138 1299 2144 1300
rect 2138 1295 2139 1299
rect 2143 1295 2144 1299
rect 2160 1295 2162 1314
rect 2220 1300 2222 1314
rect 2218 1299 2224 1300
rect 2218 1295 2219 1299
rect 2223 1295 2224 1299
rect 2240 1295 2242 1314
rect 1799 1294 1803 1295
rect 1799 1289 1803 1290
rect 1823 1294 1827 1295
rect 1886 1294 1892 1295
rect 1895 1294 1899 1295
rect 1823 1289 1827 1290
rect 1895 1289 1899 1290
rect 1911 1294 1915 1295
rect 1911 1289 1915 1290
rect 1991 1294 1995 1295
rect 1991 1289 1995 1290
rect 1999 1294 2003 1295
rect 2010 1294 2016 1295
rect 2079 1294 2083 1295
rect 1999 1289 2003 1290
rect 1778 1287 1784 1288
rect 1778 1283 1779 1287
rect 1783 1283 1784 1287
rect 1778 1282 1784 1283
rect 1800 1270 1802 1289
rect 1830 1287 1836 1288
rect 1830 1283 1831 1287
rect 1835 1283 1836 1287
rect 1830 1282 1836 1283
rect 1630 1269 1636 1270
rect 1630 1265 1631 1269
rect 1635 1265 1636 1269
rect 1630 1264 1636 1265
rect 1710 1269 1716 1270
rect 1710 1265 1711 1269
rect 1715 1265 1716 1269
rect 1798 1269 1804 1270
rect 1710 1264 1716 1265
rect 1718 1267 1724 1268
rect 1718 1263 1719 1267
rect 1723 1263 1724 1267
rect 1798 1265 1799 1269
rect 1803 1265 1804 1269
rect 1832 1268 1834 1282
rect 1896 1270 1898 1289
rect 1992 1270 1994 1289
rect 1894 1269 1900 1270
rect 1798 1264 1804 1265
rect 1830 1267 1836 1268
rect 1718 1262 1724 1263
rect 1830 1263 1831 1267
rect 1835 1263 1836 1267
rect 1894 1265 1895 1269
rect 1899 1265 1900 1269
rect 1894 1264 1900 1265
rect 1990 1269 1996 1270
rect 1990 1265 1991 1269
rect 1995 1265 1996 1269
rect 2012 1268 2014 1294
rect 2079 1289 2083 1290
rect 2095 1294 2099 1295
rect 2138 1294 2144 1295
rect 2159 1294 2163 1295
rect 2095 1289 2099 1290
rect 2159 1289 2163 1290
rect 2207 1294 2211 1295
rect 2218 1294 2224 1295
rect 2239 1294 2243 1295
rect 2207 1289 2211 1290
rect 2239 1289 2243 1290
rect 2066 1287 2072 1288
rect 2066 1283 2067 1287
rect 2071 1283 2072 1287
rect 2066 1282 2072 1283
rect 1990 1264 1996 1265
rect 2010 1267 2016 1268
rect 1830 1262 1836 1263
rect 2010 1263 2011 1267
rect 2015 1263 2016 1267
rect 2010 1262 2016 1263
rect 1614 1248 1620 1249
rect 1614 1244 1615 1248
rect 1619 1244 1620 1248
rect 1614 1243 1620 1244
rect 1694 1248 1700 1249
rect 1694 1244 1695 1248
rect 1699 1244 1700 1248
rect 1694 1243 1700 1244
rect 1616 1239 1618 1243
rect 1696 1239 1698 1243
rect 1615 1238 1619 1239
rect 1615 1233 1619 1234
rect 1631 1238 1635 1239
rect 1631 1233 1635 1234
rect 1687 1238 1691 1239
rect 1687 1233 1691 1234
rect 1695 1238 1699 1239
rect 1695 1233 1699 1234
rect 1630 1232 1636 1233
rect 1630 1228 1631 1232
rect 1635 1228 1636 1232
rect 1630 1227 1636 1228
rect 1686 1232 1692 1233
rect 1686 1228 1687 1232
rect 1691 1228 1692 1232
rect 1686 1227 1692 1228
rect 647 1210 651 1211
rect 647 1205 651 1206
rect 679 1210 683 1211
rect 679 1205 683 1206
rect 719 1210 723 1211
rect 719 1205 723 1206
rect 751 1210 755 1211
rect 751 1205 755 1206
rect 791 1210 795 1211
rect 791 1205 795 1206
rect 823 1210 827 1211
rect 823 1205 827 1206
rect 863 1210 867 1211
rect 863 1205 867 1206
rect 903 1210 907 1211
rect 903 1205 907 1206
rect 1287 1210 1291 1211
rect 1326 1208 1327 1212
rect 1331 1208 1332 1212
rect 1326 1207 1332 1208
rect 1534 1211 1540 1212
rect 1534 1207 1535 1211
rect 1539 1207 1540 1211
rect 1287 1205 1291 1206
rect 646 1204 652 1205
rect 646 1200 647 1204
rect 651 1200 652 1204
rect 646 1199 652 1200
rect 718 1204 724 1205
rect 718 1200 719 1204
rect 723 1200 724 1204
rect 718 1199 724 1200
rect 790 1204 796 1205
rect 790 1200 791 1204
rect 795 1200 796 1204
rect 790 1199 796 1200
rect 862 1204 868 1205
rect 862 1200 863 1204
rect 867 1200 868 1204
rect 1288 1202 1290 1205
rect 862 1199 868 1200
rect 1286 1201 1292 1202
rect 1286 1197 1287 1201
rect 1291 1197 1292 1201
rect 1286 1196 1292 1197
rect 1286 1184 1292 1185
rect 642 1183 648 1184
rect 642 1179 643 1183
rect 647 1179 648 1183
rect 642 1178 648 1179
rect 662 1183 668 1184
rect 662 1179 663 1183
rect 667 1179 668 1183
rect 662 1178 668 1179
rect 714 1183 720 1184
rect 714 1179 715 1183
rect 719 1179 720 1183
rect 714 1178 720 1179
rect 734 1183 740 1184
rect 734 1179 735 1183
rect 739 1179 740 1183
rect 734 1178 740 1179
rect 786 1183 792 1184
rect 786 1179 787 1183
rect 791 1179 792 1183
rect 786 1178 792 1179
rect 806 1183 812 1184
rect 806 1179 807 1183
rect 811 1179 812 1183
rect 806 1178 812 1179
rect 858 1183 864 1184
rect 858 1179 859 1183
rect 863 1179 864 1183
rect 858 1178 864 1179
rect 878 1183 884 1184
rect 878 1179 879 1183
rect 883 1179 884 1183
rect 878 1178 884 1179
rect 886 1183 892 1184
rect 886 1179 887 1183
rect 891 1179 892 1183
rect 1286 1180 1287 1184
rect 1291 1180 1292 1184
rect 1328 1183 1330 1207
rect 1534 1206 1540 1207
rect 1570 1211 1576 1212
rect 1570 1207 1571 1211
rect 1575 1207 1576 1211
rect 1570 1206 1576 1207
rect 1590 1211 1596 1212
rect 1590 1207 1591 1211
rect 1595 1207 1596 1211
rect 1590 1206 1596 1207
rect 1606 1211 1612 1212
rect 1606 1207 1607 1211
rect 1611 1207 1612 1211
rect 1606 1206 1612 1207
rect 1646 1211 1652 1212
rect 1646 1207 1647 1211
rect 1651 1207 1652 1211
rect 1646 1206 1652 1207
rect 1682 1211 1688 1212
rect 1682 1207 1683 1211
rect 1687 1207 1688 1211
rect 1682 1206 1688 1207
rect 1702 1211 1708 1212
rect 1702 1207 1703 1211
rect 1707 1207 1708 1211
rect 1702 1206 1708 1207
rect 1536 1183 1538 1206
rect 1572 1192 1574 1206
rect 1570 1191 1576 1192
rect 1570 1187 1571 1191
rect 1575 1187 1576 1191
rect 1570 1186 1576 1187
rect 1592 1183 1594 1206
rect 1648 1183 1650 1206
rect 1684 1192 1686 1206
rect 1682 1191 1688 1192
rect 1682 1187 1683 1191
rect 1687 1187 1688 1191
rect 1682 1186 1688 1187
rect 1704 1183 1706 1206
rect 1720 1200 1722 1262
rect 1782 1248 1788 1249
rect 1782 1244 1783 1248
rect 1787 1244 1788 1248
rect 1782 1243 1788 1244
rect 1878 1248 1884 1249
rect 1878 1244 1879 1248
rect 1883 1244 1884 1248
rect 1878 1243 1884 1244
rect 1974 1248 1980 1249
rect 1974 1244 1975 1248
rect 1979 1244 1980 1248
rect 1974 1243 1980 1244
rect 1784 1239 1786 1243
rect 1880 1239 1882 1243
rect 1976 1239 1978 1243
rect 1743 1238 1747 1239
rect 1743 1233 1747 1234
rect 1783 1238 1787 1239
rect 1783 1233 1787 1234
rect 1799 1238 1803 1239
rect 1799 1233 1803 1234
rect 1855 1238 1859 1239
rect 1855 1233 1859 1234
rect 1879 1238 1883 1239
rect 1879 1233 1883 1234
rect 1911 1238 1915 1239
rect 1911 1233 1915 1234
rect 1967 1238 1971 1239
rect 1967 1233 1971 1234
rect 1975 1238 1979 1239
rect 1975 1233 1979 1234
rect 2031 1238 2035 1239
rect 2031 1233 2035 1234
rect 1742 1232 1748 1233
rect 1742 1228 1743 1232
rect 1747 1228 1748 1232
rect 1742 1227 1748 1228
rect 1798 1232 1804 1233
rect 1798 1228 1799 1232
rect 1803 1228 1804 1232
rect 1798 1227 1804 1228
rect 1854 1232 1860 1233
rect 1854 1228 1855 1232
rect 1859 1228 1860 1232
rect 1854 1227 1860 1228
rect 1910 1232 1916 1233
rect 1910 1228 1911 1232
rect 1915 1228 1916 1232
rect 1910 1227 1916 1228
rect 1966 1232 1972 1233
rect 1966 1228 1967 1232
rect 1971 1228 1972 1232
rect 1966 1227 1972 1228
rect 2030 1232 2036 1233
rect 2030 1228 2031 1232
rect 2035 1228 2036 1232
rect 2030 1227 2036 1228
rect 2068 1212 2070 1282
rect 2096 1270 2098 1289
rect 2208 1270 2210 1289
rect 2300 1288 2302 1314
rect 2320 1295 2322 1314
rect 2328 1300 2330 1366
rect 2382 1352 2388 1353
rect 2382 1348 2383 1352
rect 2387 1348 2388 1352
rect 2382 1347 2388 1348
rect 2383 1346 2387 1347
rect 2383 1341 2387 1342
rect 2382 1340 2388 1341
rect 2382 1336 2383 1340
rect 2387 1336 2388 1340
rect 2382 1335 2388 1336
rect 2416 1320 2418 1386
rect 2424 1372 2426 1386
rect 2456 1374 2458 1393
rect 2454 1373 2460 1374
rect 2504 1373 2506 1393
rect 2422 1371 2428 1372
rect 2422 1367 2423 1371
rect 2427 1367 2428 1371
rect 2454 1369 2455 1373
rect 2459 1369 2460 1373
rect 2502 1372 2508 1373
rect 2454 1368 2460 1369
rect 2462 1371 2468 1372
rect 2422 1366 2428 1367
rect 2462 1367 2463 1371
rect 2467 1367 2468 1371
rect 2502 1368 2503 1372
rect 2507 1368 2508 1372
rect 2502 1367 2508 1368
rect 2462 1366 2468 1367
rect 2438 1352 2444 1353
rect 2438 1348 2439 1352
rect 2443 1348 2444 1352
rect 2438 1347 2444 1348
rect 2439 1346 2443 1347
rect 2439 1341 2443 1342
rect 2438 1340 2444 1341
rect 2438 1336 2439 1340
rect 2443 1336 2444 1340
rect 2438 1335 2444 1336
rect 2398 1319 2404 1320
rect 2398 1315 2399 1319
rect 2403 1315 2404 1319
rect 2398 1314 2404 1315
rect 2414 1319 2420 1320
rect 2414 1315 2415 1319
rect 2419 1315 2420 1319
rect 2414 1314 2420 1315
rect 2454 1319 2460 1320
rect 2454 1315 2455 1319
rect 2459 1315 2460 1319
rect 2454 1314 2460 1315
rect 2326 1299 2332 1300
rect 2326 1295 2327 1299
rect 2331 1295 2332 1299
rect 2319 1294 2323 1295
rect 2326 1294 2332 1295
rect 2390 1299 2396 1300
rect 2390 1295 2391 1299
rect 2395 1295 2396 1299
rect 2400 1295 2402 1314
rect 2456 1295 2458 1314
rect 2464 1300 2466 1366
rect 2502 1355 2508 1356
rect 2502 1351 2503 1355
rect 2507 1351 2508 1355
rect 2502 1350 2508 1351
rect 2504 1347 2506 1350
rect 2503 1346 2507 1347
rect 2503 1341 2507 1342
rect 2504 1338 2506 1341
rect 2502 1337 2508 1338
rect 2502 1333 2503 1337
rect 2507 1333 2508 1337
rect 2502 1332 2508 1333
rect 2502 1320 2508 1321
rect 2470 1319 2476 1320
rect 2470 1315 2471 1319
rect 2475 1315 2476 1319
rect 2502 1316 2503 1320
rect 2507 1316 2508 1320
rect 2502 1315 2508 1316
rect 2470 1314 2476 1315
rect 2462 1299 2468 1300
rect 2462 1295 2463 1299
rect 2467 1295 2468 1299
rect 2390 1294 2396 1295
rect 2399 1294 2403 1295
rect 2319 1289 2323 1290
rect 2298 1287 2304 1288
rect 2298 1283 2299 1287
rect 2303 1283 2304 1287
rect 2298 1282 2304 1283
rect 2320 1270 2322 1289
rect 2094 1269 2100 1270
rect 2094 1265 2095 1269
rect 2099 1265 2100 1269
rect 2206 1269 2212 1270
rect 2094 1264 2100 1265
rect 2110 1267 2116 1268
rect 2110 1263 2111 1267
rect 2115 1263 2116 1267
rect 2206 1265 2207 1269
rect 2211 1265 2212 1269
rect 2206 1264 2212 1265
rect 2318 1269 2324 1270
rect 2318 1265 2319 1269
rect 2323 1265 2324 1269
rect 2318 1264 2324 1265
rect 2110 1262 2116 1263
rect 2078 1248 2084 1249
rect 2078 1244 2079 1248
rect 2083 1244 2084 1248
rect 2078 1243 2084 1244
rect 2080 1239 2082 1243
rect 2079 1238 2083 1239
rect 2079 1233 2083 1234
rect 2103 1238 2107 1239
rect 2103 1233 2107 1234
rect 2102 1232 2108 1233
rect 2102 1228 2103 1232
rect 2107 1228 2108 1232
rect 2102 1227 2108 1228
rect 1738 1211 1744 1212
rect 1738 1207 1739 1211
rect 1743 1207 1744 1211
rect 1738 1206 1744 1207
rect 1758 1211 1764 1212
rect 1758 1207 1759 1211
rect 1763 1207 1764 1211
rect 1758 1206 1764 1207
rect 1794 1211 1800 1212
rect 1794 1207 1795 1211
rect 1799 1207 1800 1211
rect 1794 1206 1800 1207
rect 1814 1211 1820 1212
rect 1814 1207 1815 1211
rect 1819 1207 1820 1211
rect 1814 1206 1820 1207
rect 1850 1211 1856 1212
rect 1850 1207 1851 1211
rect 1855 1207 1856 1211
rect 1850 1206 1856 1207
rect 1870 1211 1876 1212
rect 1870 1207 1871 1211
rect 1875 1207 1876 1211
rect 1870 1206 1876 1207
rect 1906 1211 1912 1212
rect 1906 1207 1907 1211
rect 1911 1207 1912 1211
rect 1906 1206 1912 1207
rect 1926 1211 1932 1212
rect 1926 1207 1927 1211
rect 1931 1207 1932 1211
rect 1926 1206 1932 1207
rect 1962 1211 1968 1212
rect 1962 1207 1963 1211
rect 1967 1207 1968 1211
rect 1962 1206 1968 1207
rect 1982 1211 1988 1212
rect 1982 1207 1983 1211
rect 1987 1207 1988 1211
rect 1982 1206 1988 1207
rect 2026 1211 2032 1212
rect 2026 1207 2027 1211
rect 2031 1207 2032 1211
rect 2026 1206 2032 1207
rect 2046 1211 2052 1212
rect 2046 1207 2047 1211
rect 2051 1207 2052 1211
rect 2046 1206 2052 1207
rect 2066 1211 2072 1212
rect 2066 1207 2067 1211
rect 2071 1207 2072 1211
rect 2066 1206 2072 1207
rect 1718 1199 1724 1200
rect 1718 1195 1719 1199
rect 1723 1195 1724 1199
rect 1718 1194 1724 1195
rect 1740 1192 1742 1206
rect 1738 1191 1744 1192
rect 1738 1187 1739 1191
rect 1743 1187 1744 1191
rect 1738 1186 1744 1187
rect 1760 1183 1762 1206
rect 1796 1192 1798 1206
rect 1794 1191 1800 1192
rect 1794 1187 1795 1191
rect 1799 1187 1800 1191
rect 1794 1186 1800 1187
rect 1806 1183 1812 1184
rect 1816 1183 1818 1206
rect 1852 1192 1854 1206
rect 1850 1191 1856 1192
rect 1850 1187 1851 1191
rect 1855 1187 1856 1191
rect 1850 1186 1856 1187
rect 1872 1183 1874 1206
rect 1908 1192 1910 1206
rect 1906 1191 1912 1192
rect 1906 1187 1907 1191
rect 1911 1187 1912 1191
rect 1906 1186 1912 1187
rect 1928 1183 1930 1206
rect 1964 1192 1966 1206
rect 1962 1191 1968 1192
rect 1962 1187 1963 1191
rect 1967 1187 1968 1191
rect 1962 1186 1968 1187
rect 1984 1183 1986 1206
rect 2028 1192 2030 1206
rect 2026 1191 2032 1192
rect 2026 1187 2027 1191
rect 2031 1187 2032 1191
rect 2026 1186 2032 1187
rect 2048 1183 2050 1206
rect 2112 1192 2114 1262
rect 2190 1248 2196 1249
rect 2190 1244 2191 1248
rect 2195 1244 2196 1248
rect 2190 1243 2196 1244
rect 2302 1248 2308 1249
rect 2302 1244 2303 1248
rect 2307 1244 2308 1248
rect 2302 1243 2308 1244
rect 2192 1239 2194 1243
rect 2304 1239 2306 1243
rect 2183 1238 2187 1239
rect 2183 1233 2187 1234
rect 2191 1238 2195 1239
rect 2191 1233 2195 1234
rect 2271 1238 2275 1239
rect 2271 1233 2275 1234
rect 2303 1238 2307 1239
rect 2303 1233 2307 1234
rect 2367 1238 2371 1239
rect 2367 1233 2371 1234
rect 2182 1232 2188 1233
rect 2182 1228 2183 1232
rect 2187 1228 2188 1232
rect 2182 1227 2188 1228
rect 2270 1232 2276 1233
rect 2270 1228 2271 1232
rect 2275 1228 2276 1232
rect 2270 1227 2276 1228
rect 2366 1232 2372 1233
rect 2366 1228 2367 1232
rect 2371 1228 2372 1232
rect 2366 1227 2372 1228
rect 2392 1212 2394 1294
rect 2399 1289 2403 1290
rect 2455 1294 2459 1295
rect 2462 1294 2468 1295
rect 2455 1289 2459 1290
rect 2439 1238 2443 1239
rect 2439 1233 2443 1234
rect 2438 1232 2444 1233
rect 2438 1228 2439 1232
rect 2443 1228 2444 1232
rect 2438 1227 2444 1228
rect 2118 1211 2124 1212
rect 2118 1207 2119 1211
rect 2123 1207 2124 1211
rect 2118 1206 2124 1207
rect 2178 1211 2184 1212
rect 2178 1207 2179 1211
rect 2183 1207 2184 1211
rect 2178 1206 2184 1207
rect 2198 1211 2204 1212
rect 2198 1207 2199 1211
rect 2203 1207 2204 1211
rect 2198 1206 2204 1207
rect 2266 1211 2272 1212
rect 2266 1207 2267 1211
rect 2271 1207 2272 1211
rect 2266 1206 2272 1207
rect 2286 1211 2292 1212
rect 2286 1207 2287 1211
rect 2291 1207 2292 1211
rect 2286 1206 2292 1207
rect 2306 1211 2312 1212
rect 2306 1207 2307 1211
rect 2311 1207 2312 1211
rect 2306 1206 2312 1207
rect 2382 1211 2388 1212
rect 2382 1207 2383 1211
rect 2387 1207 2388 1211
rect 2382 1206 2388 1207
rect 2390 1211 2396 1212
rect 2390 1207 2391 1211
rect 2395 1207 2396 1211
rect 2390 1206 2396 1207
rect 2454 1211 2460 1212
rect 2454 1207 2455 1211
rect 2459 1207 2460 1211
rect 2454 1206 2460 1207
rect 2462 1211 2468 1212
rect 2462 1207 2463 1211
rect 2467 1207 2468 1211
rect 2462 1206 2468 1207
rect 2110 1191 2116 1192
rect 2110 1187 2111 1191
rect 2115 1187 2116 1191
rect 2110 1186 2116 1187
rect 2120 1183 2122 1206
rect 2180 1192 2182 1206
rect 2178 1191 2184 1192
rect 2178 1187 2179 1191
rect 2183 1187 2184 1191
rect 2178 1186 2184 1187
rect 2200 1183 2202 1206
rect 2268 1192 2270 1206
rect 2266 1191 2272 1192
rect 2266 1187 2267 1191
rect 2271 1187 2272 1191
rect 2266 1186 2272 1187
rect 2288 1183 2290 1206
rect 1286 1179 1292 1180
rect 1327 1182 1331 1183
rect 886 1178 892 1179
rect 644 1164 646 1178
rect 630 1163 636 1164
rect 630 1159 631 1163
rect 635 1159 636 1163
rect 630 1158 636 1159
rect 642 1163 648 1164
rect 642 1159 643 1163
rect 647 1159 648 1163
rect 642 1158 648 1159
rect 664 1155 666 1178
rect 716 1164 718 1178
rect 714 1163 720 1164
rect 714 1159 715 1163
rect 719 1159 720 1163
rect 714 1158 720 1159
rect 736 1155 738 1178
rect 788 1164 790 1178
rect 786 1163 792 1164
rect 786 1159 787 1163
rect 791 1159 792 1163
rect 786 1158 792 1159
rect 808 1155 810 1178
rect 860 1164 862 1178
rect 858 1163 864 1164
rect 858 1159 859 1163
rect 863 1159 864 1163
rect 858 1158 864 1159
rect 880 1155 882 1178
rect 888 1156 890 1178
rect 886 1155 892 1156
rect 1288 1155 1290 1179
rect 1327 1177 1331 1178
rect 1535 1182 1539 1183
rect 1535 1177 1539 1178
rect 1567 1182 1571 1183
rect 1567 1177 1571 1178
rect 1591 1182 1595 1183
rect 1591 1177 1595 1178
rect 1631 1182 1635 1183
rect 1631 1177 1635 1178
rect 1647 1182 1651 1183
rect 1647 1177 1651 1178
rect 1703 1182 1707 1183
rect 1703 1177 1707 1178
rect 1759 1182 1763 1183
rect 1759 1177 1763 1178
rect 1791 1182 1795 1183
rect 1806 1179 1807 1183
rect 1811 1179 1812 1183
rect 1806 1178 1812 1179
rect 1815 1182 1819 1183
rect 1791 1177 1795 1178
rect 1328 1157 1330 1177
rect 1568 1158 1570 1177
rect 1598 1175 1604 1176
rect 1598 1171 1599 1175
rect 1603 1171 1604 1175
rect 1598 1170 1604 1171
rect 1566 1157 1572 1158
rect 1326 1156 1332 1157
rect 527 1154 531 1155
rect 527 1149 531 1150
rect 567 1154 571 1155
rect 567 1149 571 1150
rect 599 1154 603 1155
rect 599 1149 603 1150
rect 655 1154 659 1155
rect 655 1149 659 1150
rect 663 1154 667 1155
rect 663 1149 667 1150
rect 735 1154 739 1155
rect 735 1149 739 1150
rect 807 1154 811 1155
rect 807 1149 811 1150
rect 879 1154 883 1155
rect 886 1151 887 1155
rect 891 1151 892 1155
rect 886 1150 892 1151
rect 959 1154 963 1155
rect 879 1149 883 1150
rect 959 1149 963 1150
rect 1039 1154 1043 1155
rect 1039 1149 1043 1150
rect 1287 1154 1291 1155
rect 1326 1152 1327 1156
rect 1331 1152 1332 1156
rect 1566 1153 1567 1157
rect 1571 1153 1572 1157
rect 1600 1156 1602 1170
rect 1632 1158 1634 1177
rect 1654 1175 1660 1176
rect 1654 1171 1655 1175
rect 1659 1171 1660 1175
rect 1654 1170 1660 1171
rect 1630 1157 1636 1158
rect 1566 1152 1572 1153
rect 1598 1155 1604 1156
rect 1326 1151 1332 1152
rect 1598 1151 1599 1155
rect 1603 1151 1604 1155
rect 1630 1153 1631 1157
rect 1635 1153 1636 1157
rect 1656 1156 1658 1170
rect 1704 1158 1706 1177
rect 1726 1175 1732 1176
rect 1726 1171 1727 1175
rect 1731 1171 1732 1175
rect 1726 1170 1732 1171
rect 1702 1157 1708 1158
rect 1630 1152 1636 1153
rect 1654 1155 1660 1156
rect 1598 1150 1604 1151
rect 1654 1151 1655 1155
rect 1659 1151 1660 1155
rect 1702 1153 1703 1157
rect 1707 1153 1708 1157
rect 1728 1156 1730 1170
rect 1782 1167 1788 1168
rect 1782 1163 1783 1167
rect 1787 1163 1788 1167
rect 1782 1162 1788 1163
rect 1702 1152 1708 1153
rect 1726 1155 1732 1156
rect 1654 1150 1660 1151
rect 1726 1151 1727 1155
rect 1731 1151 1732 1155
rect 1726 1150 1732 1151
rect 1287 1149 1291 1150
rect 568 1130 570 1149
rect 578 1147 584 1148
rect 578 1143 579 1147
rect 583 1143 584 1147
rect 578 1142 584 1143
rect 566 1129 572 1130
rect 470 1124 476 1125
rect 494 1127 500 1128
rect 198 1122 204 1123
rect 494 1123 495 1127
rect 499 1123 500 1127
rect 566 1125 567 1129
rect 571 1125 572 1129
rect 566 1124 572 1125
rect 494 1122 500 1123
rect 110 1111 116 1112
rect 110 1107 111 1111
rect 115 1107 116 1111
rect 110 1106 116 1107
rect 166 1108 172 1109
rect 112 1095 114 1106
rect 166 1104 167 1108
rect 171 1104 172 1108
rect 166 1103 172 1104
rect 168 1095 170 1103
rect 111 1094 115 1095
rect 111 1089 115 1090
rect 167 1094 171 1095
rect 167 1089 171 1090
rect 112 1086 114 1089
rect 110 1085 116 1086
rect 110 1081 111 1085
rect 115 1081 116 1085
rect 110 1080 116 1081
rect 110 1068 116 1069
rect 110 1064 111 1068
rect 115 1064 116 1068
rect 110 1063 116 1064
rect 112 1035 114 1063
rect 200 1048 202 1122
rect 262 1108 268 1109
rect 262 1104 263 1108
rect 267 1104 268 1108
rect 262 1103 268 1104
rect 358 1108 364 1109
rect 358 1104 359 1108
rect 363 1104 364 1108
rect 358 1103 364 1104
rect 454 1108 460 1109
rect 454 1104 455 1108
rect 459 1104 460 1108
rect 454 1103 460 1104
rect 550 1108 556 1109
rect 550 1104 551 1108
rect 555 1104 556 1108
rect 550 1103 556 1104
rect 264 1095 266 1103
rect 360 1095 362 1103
rect 456 1095 458 1103
rect 552 1095 554 1103
rect 207 1094 211 1095
rect 207 1089 211 1090
rect 263 1094 267 1095
rect 263 1089 267 1090
rect 279 1094 283 1095
rect 279 1089 283 1090
rect 359 1094 363 1095
rect 359 1089 363 1090
rect 447 1094 451 1095
rect 447 1089 451 1090
rect 455 1094 459 1095
rect 455 1089 459 1090
rect 543 1094 547 1095
rect 543 1089 547 1090
rect 551 1094 555 1095
rect 551 1089 555 1090
rect 206 1088 212 1089
rect 206 1084 207 1088
rect 211 1084 212 1088
rect 206 1083 212 1084
rect 278 1088 284 1089
rect 278 1084 279 1088
rect 283 1084 284 1088
rect 278 1083 284 1084
rect 358 1088 364 1089
rect 358 1084 359 1088
rect 363 1084 364 1088
rect 358 1083 364 1084
rect 446 1088 452 1089
rect 446 1084 447 1088
rect 451 1084 452 1088
rect 446 1083 452 1084
rect 542 1088 548 1089
rect 542 1084 543 1088
rect 547 1084 548 1088
rect 542 1083 548 1084
rect 580 1068 582 1142
rect 656 1130 658 1149
rect 736 1130 738 1149
rect 758 1147 764 1148
rect 758 1143 759 1147
rect 763 1143 764 1147
rect 758 1142 764 1143
rect 654 1129 660 1130
rect 654 1125 655 1129
rect 659 1125 660 1129
rect 654 1124 660 1125
rect 734 1129 740 1130
rect 734 1125 735 1129
rect 739 1125 740 1129
rect 760 1128 762 1142
rect 808 1130 810 1149
rect 826 1147 832 1148
rect 826 1143 827 1147
rect 831 1143 832 1147
rect 826 1142 832 1143
rect 806 1129 812 1130
rect 734 1124 740 1125
rect 758 1127 764 1128
rect 758 1123 759 1127
rect 763 1123 764 1127
rect 806 1125 807 1129
rect 811 1125 812 1129
rect 828 1128 830 1142
rect 880 1130 882 1149
rect 902 1147 908 1148
rect 902 1143 903 1147
rect 907 1143 908 1147
rect 902 1142 908 1143
rect 878 1129 884 1130
rect 806 1124 812 1125
rect 826 1127 832 1128
rect 758 1122 764 1123
rect 826 1123 827 1127
rect 831 1123 832 1127
rect 878 1125 879 1129
rect 883 1125 884 1129
rect 904 1128 906 1142
rect 960 1130 962 1149
rect 982 1147 988 1148
rect 982 1143 983 1147
rect 987 1143 988 1147
rect 982 1142 988 1143
rect 958 1129 964 1130
rect 878 1124 884 1125
rect 902 1127 908 1128
rect 826 1122 832 1123
rect 902 1123 903 1127
rect 907 1123 908 1127
rect 958 1125 959 1129
rect 963 1125 964 1129
rect 984 1128 986 1142
rect 1040 1130 1042 1149
rect 1038 1129 1044 1130
rect 1288 1129 1290 1149
rect 1326 1139 1332 1140
rect 1326 1135 1327 1139
rect 1331 1135 1332 1139
rect 1326 1134 1332 1135
rect 1550 1136 1556 1137
rect 1328 1131 1330 1134
rect 1550 1132 1551 1136
rect 1555 1132 1556 1136
rect 1550 1131 1556 1132
rect 1614 1136 1620 1137
rect 1614 1132 1615 1136
rect 1619 1132 1620 1136
rect 1614 1131 1620 1132
rect 1686 1136 1692 1137
rect 1686 1132 1687 1136
rect 1691 1132 1692 1136
rect 1686 1131 1692 1132
rect 1774 1136 1780 1137
rect 1774 1132 1775 1136
rect 1779 1132 1780 1136
rect 1774 1131 1780 1132
rect 1327 1130 1331 1131
rect 958 1124 964 1125
rect 982 1127 988 1128
rect 902 1122 908 1123
rect 982 1123 983 1127
rect 987 1123 988 1127
rect 1038 1125 1039 1129
rect 1043 1125 1044 1129
rect 1286 1128 1292 1129
rect 1038 1124 1044 1125
rect 1062 1127 1068 1128
rect 982 1122 988 1123
rect 1062 1123 1063 1127
rect 1067 1123 1068 1127
rect 1286 1124 1287 1128
rect 1291 1124 1292 1128
rect 1327 1125 1331 1126
rect 1383 1130 1387 1131
rect 1383 1125 1387 1126
rect 1447 1130 1451 1131
rect 1447 1125 1451 1126
rect 1519 1130 1523 1131
rect 1519 1125 1523 1126
rect 1551 1130 1555 1131
rect 1551 1125 1555 1126
rect 1591 1130 1595 1131
rect 1591 1125 1595 1126
rect 1615 1130 1619 1131
rect 1615 1125 1619 1126
rect 1671 1130 1675 1131
rect 1671 1125 1675 1126
rect 1687 1130 1691 1131
rect 1687 1125 1691 1126
rect 1751 1130 1755 1131
rect 1751 1125 1755 1126
rect 1775 1130 1779 1131
rect 1775 1125 1779 1126
rect 1286 1123 1292 1124
rect 1062 1122 1068 1123
rect 1328 1122 1330 1125
rect 1382 1124 1388 1125
rect 638 1108 644 1109
rect 638 1104 639 1108
rect 643 1104 644 1108
rect 638 1103 644 1104
rect 718 1108 724 1109
rect 718 1104 719 1108
rect 723 1104 724 1108
rect 718 1103 724 1104
rect 790 1108 796 1109
rect 790 1104 791 1108
rect 795 1104 796 1108
rect 790 1103 796 1104
rect 862 1108 868 1109
rect 862 1104 863 1108
rect 867 1104 868 1108
rect 862 1103 868 1104
rect 942 1108 948 1109
rect 942 1104 943 1108
rect 947 1104 948 1108
rect 942 1103 948 1104
rect 1022 1108 1028 1109
rect 1022 1104 1023 1108
rect 1027 1104 1028 1108
rect 1022 1103 1028 1104
rect 640 1095 642 1103
rect 720 1095 722 1103
rect 792 1095 794 1103
rect 864 1095 866 1103
rect 944 1095 946 1103
rect 1024 1095 1026 1103
rect 639 1094 643 1095
rect 639 1089 643 1090
rect 719 1094 723 1095
rect 719 1089 723 1090
rect 727 1094 731 1095
rect 727 1089 731 1090
rect 791 1094 795 1095
rect 791 1089 795 1090
rect 815 1094 819 1095
rect 815 1089 819 1090
rect 863 1094 867 1095
rect 863 1089 867 1090
rect 895 1094 899 1095
rect 895 1089 899 1090
rect 943 1094 947 1095
rect 943 1089 947 1090
rect 975 1094 979 1095
rect 975 1089 979 1090
rect 1023 1094 1027 1095
rect 1023 1089 1027 1090
rect 1055 1094 1059 1095
rect 1055 1089 1059 1090
rect 638 1088 644 1089
rect 638 1084 639 1088
rect 643 1084 644 1088
rect 638 1083 644 1084
rect 726 1088 732 1089
rect 726 1084 727 1088
rect 731 1084 732 1088
rect 726 1083 732 1084
rect 814 1088 820 1089
rect 814 1084 815 1088
rect 819 1084 820 1088
rect 814 1083 820 1084
rect 894 1088 900 1089
rect 894 1084 895 1088
rect 899 1084 900 1088
rect 894 1083 900 1084
rect 974 1088 980 1089
rect 974 1084 975 1088
rect 979 1084 980 1088
rect 974 1083 980 1084
rect 1054 1088 1060 1089
rect 1054 1084 1055 1088
rect 1059 1084 1060 1088
rect 1054 1083 1060 1084
rect 222 1067 228 1068
rect 222 1063 223 1067
rect 227 1063 228 1067
rect 222 1062 228 1063
rect 274 1067 280 1068
rect 274 1063 275 1067
rect 279 1063 280 1067
rect 274 1062 280 1063
rect 294 1067 300 1068
rect 294 1063 295 1067
rect 299 1063 300 1067
rect 294 1062 300 1063
rect 354 1067 360 1068
rect 354 1063 355 1067
rect 359 1063 360 1067
rect 354 1062 360 1063
rect 374 1067 380 1068
rect 374 1063 375 1067
rect 379 1063 380 1067
rect 374 1062 380 1063
rect 442 1067 448 1068
rect 442 1063 443 1067
rect 447 1063 448 1067
rect 442 1062 448 1063
rect 462 1067 468 1068
rect 462 1063 463 1067
rect 467 1063 468 1067
rect 462 1062 468 1063
rect 470 1067 476 1068
rect 470 1063 471 1067
rect 475 1063 476 1067
rect 470 1062 476 1063
rect 558 1067 564 1068
rect 558 1063 559 1067
rect 563 1063 564 1067
rect 558 1062 564 1063
rect 578 1067 584 1068
rect 578 1063 579 1067
rect 583 1063 584 1067
rect 578 1062 584 1063
rect 654 1067 660 1068
rect 654 1063 655 1067
rect 659 1063 660 1067
rect 654 1062 660 1063
rect 742 1067 748 1068
rect 742 1063 743 1067
rect 747 1063 748 1067
rect 742 1062 748 1063
rect 810 1067 816 1068
rect 810 1063 811 1067
rect 815 1063 816 1067
rect 810 1062 816 1063
rect 830 1067 836 1068
rect 830 1063 831 1067
rect 835 1063 836 1067
rect 830 1062 836 1063
rect 890 1067 896 1068
rect 890 1063 891 1067
rect 895 1063 896 1067
rect 890 1062 896 1063
rect 910 1067 916 1068
rect 910 1063 911 1067
rect 915 1063 916 1067
rect 910 1062 916 1063
rect 970 1067 976 1068
rect 970 1063 971 1067
rect 975 1063 976 1067
rect 970 1062 976 1063
rect 990 1067 996 1068
rect 990 1063 991 1067
rect 995 1063 996 1067
rect 990 1062 996 1063
rect 1050 1067 1056 1068
rect 1050 1063 1051 1067
rect 1055 1063 1056 1067
rect 1050 1062 1056 1063
rect 198 1047 204 1048
rect 198 1043 199 1047
rect 203 1043 204 1047
rect 198 1042 204 1043
rect 224 1035 226 1062
rect 276 1048 278 1062
rect 274 1047 280 1048
rect 274 1043 275 1047
rect 279 1043 280 1047
rect 274 1042 280 1043
rect 296 1035 298 1062
rect 356 1048 358 1062
rect 354 1047 360 1048
rect 354 1043 355 1047
rect 359 1043 360 1047
rect 354 1042 360 1043
rect 376 1035 378 1062
rect 444 1048 446 1062
rect 442 1047 448 1048
rect 442 1043 443 1047
rect 447 1043 448 1047
rect 442 1042 448 1043
rect 464 1035 466 1062
rect 111 1034 115 1035
rect 111 1029 115 1030
rect 223 1034 227 1035
rect 223 1029 227 1030
rect 295 1034 299 1035
rect 295 1029 299 1030
rect 375 1034 379 1035
rect 375 1029 379 1030
rect 383 1034 387 1035
rect 383 1029 387 1030
rect 463 1034 467 1035
rect 463 1029 467 1030
rect 112 1009 114 1029
rect 296 1010 298 1029
rect 384 1010 386 1029
rect 472 1028 474 1062
rect 560 1035 562 1062
rect 598 1047 604 1048
rect 598 1043 599 1047
rect 603 1043 604 1047
rect 598 1042 604 1043
rect 479 1034 483 1035
rect 479 1029 483 1030
rect 559 1034 563 1035
rect 559 1029 563 1030
rect 575 1034 579 1035
rect 575 1029 579 1030
rect 470 1027 476 1028
rect 470 1023 471 1027
rect 475 1023 476 1027
rect 470 1022 476 1023
rect 480 1010 482 1029
rect 576 1010 578 1029
rect 294 1009 300 1010
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 294 1005 295 1009
rect 299 1005 300 1009
rect 382 1009 388 1010
rect 294 1004 300 1005
rect 302 1007 308 1008
rect 110 1003 116 1004
rect 302 1003 303 1007
rect 307 1003 308 1007
rect 382 1005 383 1009
rect 387 1005 388 1009
rect 382 1004 388 1005
rect 478 1009 484 1010
rect 478 1005 479 1009
rect 483 1005 484 1009
rect 478 1004 484 1005
rect 574 1009 580 1010
rect 574 1005 575 1009
rect 579 1005 580 1009
rect 600 1008 602 1042
rect 656 1035 658 1062
rect 744 1035 746 1062
rect 812 1048 814 1062
rect 810 1047 816 1048
rect 810 1043 811 1047
rect 815 1043 816 1047
rect 810 1042 816 1043
rect 832 1035 834 1062
rect 892 1048 894 1062
rect 890 1047 896 1048
rect 890 1043 891 1047
rect 895 1043 896 1047
rect 890 1042 896 1043
rect 912 1035 914 1062
rect 972 1048 974 1062
rect 970 1047 976 1048
rect 970 1043 971 1047
rect 975 1043 976 1047
rect 970 1042 976 1043
rect 992 1035 994 1062
rect 1052 1048 1054 1062
rect 1064 1056 1066 1122
rect 1326 1121 1332 1122
rect 1326 1117 1327 1121
rect 1331 1117 1332 1121
rect 1382 1120 1383 1124
rect 1387 1120 1388 1124
rect 1382 1119 1388 1120
rect 1446 1124 1452 1125
rect 1446 1120 1447 1124
rect 1451 1120 1452 1124
rect 1446 1119 1452 1120
rect 1518 1124 1524 1125
rect 1518 1120 1519 1124
rect 1523 1120 1524 1124
rect 1518 1119 1524 1120
rect 1590 1124 1596 1125
rect 1590 1120 1591 1124
rect 1595 1120 1596 1124
rect 1590 1119 1596 1120
rect 1670 1124 1676 1125
rect 1670 1120 1671 1124
rect 1675 1120 1676 1124
rect 1670 1119 1676 1120
rect 1750 1124 1756 1125
rect 1750 1120 1751 1124
rect 1755 1120 1756 1124
rect 1750 1119 1756 1120
rect 1326 1116 1332 1117
rect 1286 1111 1292 1112
rect 1286 1107 1287 1111
rect 1291 1107 1292 1111
rect 1286 1106 1292 1107
rect 1288 1095 1290 1106
rect 1326 1104 1332 1105
rect 1784 1104 1786 1162
rect 1792 1158 1794 1177
rect 1790 1157 1796 1158
rect 1790 1153 1791 1157
rect 1795 1153 1796 1157
rect 1808 1156 1810 1178
rect 1815 1177 1819 1178
rect 1871 1182 1875 1183
rect 1871 1177 1875 1178
rect 1903 1182 1907 1183
rect 1903 1177 1907 1178
rect 1927 1182 1931 1183
rect 1927 1177 1931 1178
rect 1983 1182 1987 1183
rect 1983 1177 1987 1178
rect 2031 1182 2035 1183
rect 2031 1177 2035 1178
rect 2047 1182 2051 1183
rect 2047 1177 2051 1178
rect 2119 1182 2123 1183
rect 2119 1177 2123 1178
rect 2175 1182 2179 1183
rect 2175 1177 2179 1178
rect 2199 1182 2203 1183
rect 2199 1177 2203 1178
rect 2287 1182 2291 1183
rect 2287 1177 2291 1178
rect 1904 1158 1906 1177
rect 2032 1158 2034 1177
rect 2176 1158 2178 1177
rect 2308 1176 2310 1206
rect 2384 1183 2386 1206
rect 2456 1183 2458 1206
rect 2327 1182 2331 1183
rect 2327 1177 2331 1178
rect 2383 1182 2387 1183
rect 2383 1177 2387 1178
rect 2455 1182 2459 1183
rect 2455 1177 2459 1178
rect 2306 1175 2312 1176
rect 2306 1171 2307 1175
rect 2311 1171 2312 1175
rect 2306 1170 2312 1171
rect 2328 1158 2330 1177
rect 2456 1158 2458 1177
rect 2464 1176 2466 1206
rect 2472 1192 2474 1314
rect 2504 1295 2506 1315
rect 2503 1294 2507 1295
rect 2503 1289 2507 1290
rect 2504 1269 2506 1289
rect 2502 1268 2508 1269
rect 2502 1264 2503 1268
rect 2507 1264 2508 1268
rect 2502 1263 2508 1264
rect 2502 1251 2508 1252
rect 2502 1247 2503 1251
rect 2507 1247 2508 1251
rect 2502 1246 2508 1247
rect 2504 1239 2506 1246
rect 2503 1238 2507 1239
rect 2503 1233 2507 1234
rect 2504 1230 2506 1233
rect 2502 1229 2508 1230
rect 2502 1225 2503 1229
rect 2507 1225 2508 1229
rect 2502 1224 2508 1225
rect 2502 1212 2508 1213
rect 2502 1208 2503 1212
rect 2507 1208 2508 1212
rect 2502 1207 2508 1208
rect 2470 1191 2476 1192
rect 2470 1187 2471 1191
rect 2475 1187 2476 1191
rect 2470 1186 2476 1187
rect 2474 1183 2480 1184
rect 2504 1183 2506 1207
rect 2474 1179 2475 1183
rect 2479 1179 2480 1183
rect 2474 1178 2480 1179
rect 2503 1182 2507 1183
rect 2462 1175 2468 1176
rect 2462 1171 2463 1175
rect 2467 1171 2468 1175
rect 2462 1170 2468 1171
rect 1902 1157 1908 1158
rect 1790 1152 1796 1153
rect 1806 1155 1812 1156
rect 1806 1151 1807 1155
rect 1811 1151 1812 1155
rect 1902 1153 1903 1157
rect 1907 1153 1908 1157
rect 2030 1157 2036 1158
rect 1902 1152 1908 1153
rect 1918 1155 1924 1156
rect 1806 1150 1812 1151
rect 1918 1151 1919 1155
rect 1923 1151 1924 1155
rect 2030 1153 2031 1157
rect 2035 1153 2036 1157
rect 2030 1152 2036 1153
rect 2174 1157 2180 1158
rect 2174 1153 2175 1157
rect 2179 1153 2180 1157
rect 2174 1152 2180 1153
rect 2326 1157 2332 1158
rect 2326 1153 2327 1157
rect 2331 1153 2332 1157
rect 2326 1152 2332 1153
rect 2454 1157 2460 1158
rect 2454 1153 2455 1157
rect 2459 1153 2460 1157
rect 2454 1152 2460 1153
rect 2462 1155 2468 1156
rect 1918 1150 1924 1151
rect 2462 1151 2463 1155
rect 2467 1151 2468 1155
rect 2462 1150 2468 1151
rect 1886 1136 1892 1137
rect 1886 1132 1887 1136
rect 1891 1132 1892 1136
rect 1886 1131 1892 1132
rect 1831 1130 1835 1131
rect 1831 1125 1835 1126
rect 1887 1130 1891 1131
rect 1887 1125 1891 1126
rect 1911 1130 1915 1131
rect 1911 1125 1915 1126
rect 1830 1124 1836 1125
rect 1830 1120 1831 1124
rect 1835 1120 1836 1124
rect 1830 1119 1836 1120
rect 1910 1124 1916 1125
rect 1910 1120 1911 1124
rect 1915 1120 1916 1124
rect 1910 1119 1916 1120
rect 1326 1100 1327 1104
rect 1331 1100 1332 1104
rect 1326 1099 1332 1100
rect 1398 1103 1404 1104
rect 1398 1099 1399 1103
rect 1403 1099 1404 1103
rect 1143 1094 1147 1095
rect 1143 1089 1147 1090
rect 1287 1094 1291 1095
rect 1287 1089 1291 1090
rect 1142 1088 1148 1089
rect 1142 1084 1143 1088
rect 1147 1084 1148 1088
rect 1288 1086 1290 1089
rect 1142 1083 1148 1084
rect 1286 1085 1292 1086
rect 1286 1081 1287 1085
rect 1291 1081 1292 1085
rect 1286 1080 1292 1081
rect 1328 1071 1330 1099
rect 1398 1098 1404 1099
rect 1442 1103 1448 1104
rect 1442 1099 1443 1103
rect 1447 1099 1448 1103
rect 1442 1098 1448 1099
rect 1462 1103 1468 1104
rect 1462 1099 1463 1103
rect 1467 1099 1468 1103
rect 1462 1098 1468 1099
rect 1514 1103 1520 1104
rect 1514 1099 1515 1103
rect 1519 1099 1520 1103
rect 1514 1098 1520 1099
rect 1534 1103 1540 1104
rect 1534 1099 1535 1103
rect 1539 1099 1540 1103
rect 1534 1098 1540 1099
rect 1586 1103 1592 1104
rect 1586 1099 1587 1103
rect 1591 1099 1592 1103
rect 1586 1098 1592 1099
rect 1606 1103 1612 1104
rect 1606 1099 1607 1103
rect 1611 1099 1612 1103
rect 1606 1098 1612 1099
rect 1666 1103 1672 1104
rect 1666 1099 1667 1103
rect 1671 1099 1672 1103
rect 1666 1098 1672 1099
rect 1686 1103 1692 1104
rect 1686 1099 1687 1103
rect 1691 1099 1692 1103
rect 1686 1098 1692 1099
rect 1746 1103 1752 1104
rect 1746 1099 1747 1103
rect 1751 1099 1752 1103
rect 1746 1098 1752 1099
rect 1766 1103 1772 1104
rect 1766 1099 1767 1103
rect 1771 1099 1772 1103
rect 1766 1098 1772 1099
rect 1782 1103 1788 1104
rect 1782 1099 1783 1103
rect 1787 1099 1788 1103
rect 1782 1098 1788 1099
rect 1846 1103 1852 1104
rect 1846 1099 1847 1103
rect 1851 1099 1852 1103
rect 1846 1098 1852 1099
rect 1906 1103 1912 1104
rect 1906 1099 1907 1103
rect 1911 1099 1912 1103
rect 1906 1098 1912 1099
rect 1400 1071 1402 1098
rect 1444 1084 1446 1098
rect 1442 1083 1448 1084
rect 1442 1079 1443 1083
rect 1447 1079 1448 1083
rect 1442 1078 1448 1079
rect 1464 1071 1466 1098
rect 1516 1084 1518 1098
rect 1514 1083 1520 1084
rect 1514 1079 1515 1083
rect 1519 1079 1520 1083
rect 1514 1078 1520 1079
rect 1536 1071 1538 1098
rect 1588 1084 1590 1098
rect 1586 1083 1592 1084
rect 1586 1079 1587 1083
rect 1591 1079 1592 1083
rect 1586 1078 1592 1079
rect 1608 1071 1610 1098
rect 1668 1084 1670 1098
rect 1666 1083 1672 1084
rect 1666 1079 1667 1083
rect 1671 1079 1672 1083
rect 1666 1078 1672 1079
rect 1688 1071 1690 1098
rect 1748 1084 1750 1098
rect 1746 1083 1752 1084
rect 1746 1079 1747 1083
rect 1751 1079 1752 1083
rect 1746 1078 1752 1079
rect 1768 1071 1770 1098
rect 1834 1075 1840 1076
rect 1834 1071 1835 1075
rect 1839 1071 1840 1075
rect 1848 1071 1850 1098
rect 1908 1084 1910 1098
rect 1920 1092 1922 1150
rect 2014 1136 2020 1137
rect 2014 1132 2015 1136
rect 2019 1132 2020 1136
rect 2014 1131 2020 1132
rect 2158 1136 2164 1137
rect 2158 1132 2159 1136
rect 2163 1132 2164 1136
rect 2158 1131 2164 1132
rect 2310 1136 2316 1137
rect 2310 1132 2311 1136
rect 2315 1132 2316 1136
rect 2310 1131 2316 1132
rect 2438 1136 2444 1137
rect 2438 1132 2439 1136
rect 2443 1132 2444 1136
rect 2438 1131 2444 1132
rect 1983 1130 1987 1131
rect 1983 1125 1987 1126
rect 2015 1130 2019 1131
rect 2015 1125 2019 1126
rect 2055 1130 2059 1131
rect 2055 1125 2059 1126
rect 2135 1130 2139 1131
rect 2135 1125 2139 1126
rect 2159 1130 2163 1131
rect 2159 1125 2163 1126
rect 2215 1130 2219 1131
rect 2215 1125 2219 1126
rect 2311 1130 2315 1131
rect 2311 1125 2315 1126
rect 2439 1130 2443 1131
rect 2439 1125 2443 1126
rect 1982 1124 1988 1125
rect 1982 1120 1983 1124
rect 1987 1120 1988 1124
rect 1982 1119 1988 1120
rect 2054 1124 2060 1125
rect 2054 1120 2055 1124
rect 2059 1120 2060 1124
rect 2054 1119 2060 1120
rect 2134 1124 2140 1125
rect 2134 1120 2135 1124
rect 2139 1120 2140 1124
rect 2134 1119 2140 1120
rect 2214 1124 2220 1125
rect 2214 1120 2215 1124
rect 2219 1120 2220 1124
rect 2214 1119 2220 1120
rect 1926 1103 1932 1104
rect 1926 1099 1927 1103
rect 1931 1099 1932 1103
rect 1926 1098 1932 1099
rect 1978 1103 1984 1104
rect 1978 1099 1979 1103
rect 1983 1099 1984 1103
rect 1978 1098 1984 1099
rect 1998 1103 2004 1104
rect 1998 1099 1999 1103
rect 2003 1099 2004 1103
rect 1998 1098 2004 1099
rect 2050 1103 2056 1104
rect 2050 1099 2051 1103
rect 2055 1099 2056 1103
rect 2050 1098 2056 1099
rect 2070 1103 2076 1104
rect 2070 1099 2071 1103
rect 2075 1099 2076 1103
rect 2070 1098 2076 1099
rect 2130 1103 2136 1104
rect 2130 1099 2131 1103
rect 2135 1099 2136 1103
rect 2130 1098 2136 1099
rect 2150 1103 2156 1104
rect 2150 1099 2151 1103
rect 2155 1099 2156 1103
rect 2150 1098 2156 1099
rect 2210 1103 2216 1104
rect 2210 1099 2211 1103
rect 2215 1099 2216 1103
rect 2210 1098 2216 1099
rect 2230 1103 2236 1104
rect 2230 1099 2231 1103
rect 2235 1099 2236 1103
rect 2230 1098 2236 1099
rect 2238 1103 2244 1104
rect 2238 1099 2239 1103
rect 2243 1099 2244 1103
rect 2238 1098 2244 1099
rect 1918 1091 1924 1092
rect 1918 1087 1919 1091
rect 1923 1087 1924 1091
rect 1918 1086 1924 1087
rect 1906 1083 1912 1084
rect 1906 1079 1907 1083
rect 1911 1079 1912 1083
rect 1906 1078 1912 1079
rect 1928 1071 1930 1098
rect 1980 1084 1982 1098
rect 1978 1083 1984 1084
rect 1978 1079 1979 1083
rect 1983 1079 1984 1083
rect 1978 1078 1984 1079
rect 2000 1071 2002 1098
rect 2052 1084 2054 1098
rect 2050 1083 2056 1084
rect 2050 1079 2051 1083
rect 2055 1079 2056 1083
rect 2050 1078 2056 1079
rect 2072 1071 2074 1098
rect 2132 1084 2134 1098
rect 2130 1083 2136 1084
rect 2130 1079 2131 1083
rect 2135 1079 2136 1083
rect 2130 1078 2136 1079
rect 2152 1071 2154 1098
rect 2212 1084 2214 1098
rect 2210 1083 2216 1084
rect 2210 1079 2211 1083
rect 2215 1079 2216 1083
rect 2210 1078 2216 1079
rect 2232 1071 2234 1098
rect 2240 1072 2242 1098
rect 2238 1071 2244 1072
rect 1327 1070 1331 1071
rect 1286 1068 1292 1069
rect 1070 1067 1076 1068
rect 1070 1063 1071 1067
rect 1075 1063 1076 1067
rect 1070 1062 1076 1063
rect 1138 1067 1144 1068
rect 1138 1063 1139 1067
rect 1143 1063 1144 1067
rect 1138 1062 1144 1063
rect 1158 1067 1164 1068
rect 1158 1063 1159 1067
rect 1163 1063 1164 1067
rect 1158 1062 1164 1063
rect 1166 1067 1172 1068
rect 1166 1063 1167 1067
rect 1171 1063 1172 1067
rect 1286 1064 1287 1068
rect 1291 1064 1292 1068
rect 1327 1065 1331 1066
rect 1367 1070 1371 1071
rect 1367 1065 1371 1066
rect 1399 1070 1403 1071
rect 1399 1065 1403 1066
rect 1455 1070 1459 1071
rect 1455 1065 1459 1066
rect 1463 1070 1467 1071
rect 1463 1065 1467 1066
rect 1535 1070 1539 1071
rect 1535 1065 1539 1066
rect 1575 1070 1579 1071
rect 1575 1065 1579 1066
rect 1607 1070 1611 1071
rect 1607 1065 1611 1066
rect 1687 1070 1691 1071
rect 1687 1065 1691 1066
rect 1695 1070 1699 1071
rect 1695 1065 1699 1066
rect 1767 1070 1771 1071
rect 1767 1065 1771 1066
rect 1815 1070 1819 1071
rect 1834 1070 1840 1071
rect 1847 1070 1851 1071
rect 1815 1065 1819 1066
rect 1286 1063 1292 1064
rect 1166 1062 1172 1063
rect 1062 1055 1068 1056
rect 1062 1051 1063 1055
rect 1067 1051 1068 1055
rect 1062 1050 1068 1051
rect 1050 1047 1056 1048
rect 1050 1043 1051 1047
rect 1055 1043 1056 1047
rect 1050 1042 1056 1043
rect 1072 1035 1074 1062
rect 1140 1048 1142 1062
rect 1138 1047 1144 1048
rect 1138 1043 1139 1047
rect 1143 1043 1144 1047
rect 1138 1042 1144 1043
rect 1160 1035 1162 1062
rect 1168 1036 1170 1062
rect 1166 1035 1172 1036
rect 1288 1035 1290 1063
rect 1328 1045 1330 1065
rect 1368 1046 1370 1065
rect 1390 1063 1396 1064
rect 1390 1059 1391 1063
rect 1395 1059 1396 1063
rect 1390 1058 1396 1059
rect 1366 1045 1372 1046
rect 1326 1044 1332 1045
rect 1326 1040 1327 1044
rect 1331 1040 1332 1044
rect 1366 1041 1367 1045
rect 1371 1041 1372 1045
rect 1392 1044 1394 1058
rect 1456 1046 1458 1065
rect 1478 1063 1484 1064
rect 1478 1059 1479 1063
rect 1483 1059 1484 1063
rect 1478 1058 1484 1059
rect 1454 1045 1460 1046
rect 1366 1040 1372 1041
rect 1390 1043 1396 1044
rect 1326 1039 1332 1040
rect 1390 1039 1391 1043
rect 1395 1039 1396 1043
rect 1454 1041 1455 1045
rect 1459 1041 1460 1045
rect 1480 1044 1482 1058
rect 1576 1046 1578 1065
rect 1598 1063 1604 1064
rect 1598 1059 1599 1063
rect 1603 1059 1604 1063
rect 1598 1058 1604 1059
rect 1574 1045 1580 1046
rect 1454 1040 1460 1041
rect 1478 1043 1484 1044
rect 1390 1038 1396 1039
rect 1478 1039 1479 1043
rect 1483 1039 1484 1043
rect 1574 1041 1575 1045
rect 1579 1041 1580 1045
rect 1600 1044 1602 1058
rect 1696 1046 1698 1065
rect 1718 1063 1724 1064
rect 1718 1059 1719 1063
rect 1723 1059 1724 1063
rect 1718 1058 1724 1059
rect 1710 1055 1716 1056
rect 1710 1051 1711 1055
rect 1715 1051 1716 1055
rect 1710 1050 1716 1051
rect 1694 1045 1700 1046
rect 1574 1040 1580 1041
rect 1598 1043 1604 1044
rect 1478 1038 1484 1039
rect 1598 1039 1599 1043
rect 1603 1039 1604 1043
rect 1694 1041 1695 1045
rect 1699 1041 1700 1045
rect 1694 1040 1700 1041
rect 1598 1038 1604 1039
rect 655 1034 659 1035
rect 655 1029 659 1030
rect 671 1034 675 1035
rect 671 1029 675 1030
rect 743 1034 747 1035
rect 743 1029 747 1030
rect 767 1034 771 1035
rect 767 1029 771 1030
rect 831 1034 835 1035
rect 831 1029 835 1030
rect 855 1034 859 1035
rect 855 1029 859 1030
rect 911 1034 915 1035
rect 911 1029 915 1030
rect 943 1034 947 1035
rect 943 1029 947 1030
rect 991 1034 995 1035
rect 991 1029 995 1030
rect 1023 1034 1027 1035
rect 1023 1029 1027 1030
rect 1071 1034 1075 1035
rect 1071 1029 1075 1030
rect 1103 1034 1107 1035
rect 1103 1029 1107 1030
rect 1159 1034 1163 1035
rect 1166 1031 1167 1035
rect 1171 1031 1172 1035
rect 1166 1030 1172 1031
rect 1183 1034 1187 1035
rect 1159 1029 1163 1030
rect 1183 1029 1187 1030
rect 1239 1034 1243 1035
rect 1239 1029 1243 1030
rect 1287 1034 1291 1035
rect 1287 1029 1291 1030
rect 672 1010 674 1029
rect 690 1027 696 1028
rect 690 1023 691 1027
rect 695 1023 696 1027
rect 690 1022 696 1023
rect 670 1009 676 1010
rect 574 1004 580 1005
rect 598 1007 604 1008
rect 302 1002 308 1003
rect 598 1003 599 1007
rect 603 1003 604 1007
rect 670 1005 671 1009
rect 675 1005 676 1009
rect 670 1004 676 1005
rect 598 1002 604 1003
rect 110 991 116 992
rect 110 987 111 991
rect 115 987 116 991
rect 110 986 116 987
rect 278 988 284 989
rect 112 983 114 986
rect 278 984 279 988
rect 283 984 284 988
rect 278 983 284 984
rect 111 982 115 983
rect 111 977 115 978
rect 271 982 275 983
rect 271 977 275 978
rect 279 982 283 983
rect 279 977 283 978
rect 112 974 114 977
rect 270 976 276 977
rect 110 973 116 974
rect 110 969 111 973
rect 115 969 116 973
rect 270 972 271 976
rect 275 972 276 976
rect 270 971 276 972
rect 110 968 116 969
rect 110 956 116 957
rect 110 952 111 956
rect 115 952 116 956
rect 110 951 116 952
rect 286 955 292 956
rect 286 951 287 955
rect 291 951 292 955
rect 112 923 114 951
rect 286 950 292 951
rect 288 923 290 950
rect 304 936 306 1002
rect 366 988 372 989
rect 366 984 367 988
rect 371 984 372 988
rect 366 983 372 984
rect 462 988 468 989
rect 462 984 463 988
rect 467 984 468 988
rect 462 983 468 984
rect 558 988 564 989
rect 558 984 559 988
rect 563 984 564 988
rect 558 983 564 984
rect 654 988 660 989
rect 654 984 655 988
rect 659 984 660 988
rect 654 983 660 984
rect 359 982 363 983
rect 359 977 363 978
rect 367 982 371 983
rect 367 977 371 978
rect 455 982 459 983
rect 455 977 459 978
rect 463 982 467 983
rect 463 977 467 978
rect 551 982 555 983
rect 551 977 555 978
rect 559 982 563 983
rect 559 977 563 978
rect 655 982 659 983
rect 655 977 659 978
rect 358 976 364 977
rect 358 972 359 976
rect 363 972 364 976
rect 358 971 364 972
rect 454 976 460 977
rect 454 972 455 976
rect 459 972 460 976
rect 454 971 460 972
rect 550 976 556 977
rect 550 972 551 976
rect 555 972 556 976
rect 550 971 556 972
rect 654 976 660 977
rect 654 972 655 976
rect 659 972 660 976
rect 654 971 660 972
rect 692 956 694 1022
rect 768 1010 770 1029
rect 790 1027 796 1028
rect 790 1023 791 1027
rect 795 1023 796 1027
rect 790 1022 796 1023
rect 766 1009 772 1010
rect 766 1005 767 1009
rect 771 1005 772 1009
rect 792 1008 794 1022
rect 856 1010 858 1029
rect 878 1027 884 1028
rect 878 1023 879 1027
rect 883 1023 884 1027
rect 878 1022 884 1023
rect 854 1009 860 1010
rect 766 1004 772 1005
rect 790 1007 796 1008
rect 790 1003 791 1007
rect 795 1003 796 1007
rect 854 1005 855 1009
rect 859 1005 860 1009
rect 880 1008 882 1022
rect 944 1010 946 1029
rect 966 1027 972 1028
rect 966 1023 967 1027
rect 971 1023 972 1027
rect 966 1022 972 1023
rect 942 1009 948 1010
rect 854 1004 860 1005
rect 878 1007 884 1008
rect 790 1002 796 1003
rect 878 1003 879 1007
rect 883 1003 884 1007
rect 942 1005 943 1009
rect 947 1005 948 1009
rect 968 1008 970 1022
rect 1024 1010 1026 1029
rect 1046 1027 1052 1028
rect 1046 1023 1047 1027
rect 1051 1023 1052 1027
rect 1046 1022 1052 1023
rect 1022 1009 1028 1010
rect 942 1004 948 1005
rect 966 1007 972 1008
rect 878 1002 884 1003
rect 966 1003 967 1007
rect 971 1003 972 1007
rect 1022 1005 1023 1009
rect 1027 1005 1028 1009
rect 1022 1004 1028 1005
rect 966 1002 972 1003
rect 750 988 756 989
rect 750 984 751 988
rect 755 984 756 988
rect 750 983 756 984
rect 838 988 844 989
rect 838 984 839 988
rect 843 984 844 988
rect 838 983 844 984
rect 926 988 932 989
rect 926 984 927 988
rect 931 984 932 988
rect 926 983 932 984
rect 1006 988 1012 989
rect 1006 984 1007 988
rect 1011 984 1012 988
rect 1006 983 1012 984
rect 751 982 755 983
rect 751 977 755 978
rect 839 982 843 983
rect 839 977 843 978
rect 927 982 931 983
rect 927 977 931 978
rect 1007 982 1011 983
rect 1007 977 1011 978
rect 750 976 756 977
rect 750 972 751 976
rect 755 972 756 976
rect 750 971 756 972
rect 838 976 844 977
rect 838 972 839 976
rect 843 972 844 976
rect 838 971 844 972
rect 926 976 932 977
rect 926 972 927 976
rect 931 972 932 976
rect 926 971 932 972
rect 1006 976 1012 977
rect 1006 972 1007 976
rect 1011 972 1012 976
rect 1006 971 1012 972
rect 1048 956 1050 1022
rect 1104 1010 1106 1029
rect 1184 1010 1186 1029
rect 1206 1027 1212 1028
rect 1206 1023 1207 1027
rect 1211 1023 1212 1027
rect 1206 1022 1212 1023
rect 1102 1009 1108 1010
rect 1102 1005 1103 1009
rect 1107 1005 1108 1009
rect 1102 1004 1108 1005
rect 1182 1009 1188 1010
rect 1182 1005 1183 1009
rect 1187 1005 1188 1009
rect 1208 1008 1210 1022
rect 1214 1015 1220 1016
rect 1214 1011 1215 1015
rect 1219 1011 1220 1015
rect 1214 1010 1220 1011
rect 1240 1010 1242 1029
rect 1182 1004 1188 1005
rect 1206 1007 1212 1008
rect 1206 1003 1207 1007
rect 1211 1003 1212 1007
rect 1206 1002 1212 1003
rect 1086 988 1092 989
rect 1086 984 1087 988
rect 1091 984 1092 988
rect 1086 983 1092 984
rect 1166 988 1172 989
rect 1166 984 1167 988
rect 1171 984 1172 988
rect 1166 983 1172 984
rect 1087 982 1091 983
rect 1087 977 1091 978
rect 1167 982 1171 983
rect 1167 977 1171 978
rect 1086 976 1092 977
rect 1086 972 1087 976
rect 1091 972 1092 976
rect 1086 971 1092 972
rect 1166 976 1172 977
rect 1166 972 1167 976
rect 1171 972 1172 976
rect 1166 971 1172 972
rect 354 955 360 956
rect 354 951 355 955
rect 359 951 360 955
rect 354 950 360 951
rect 374 955 380 956
rect 374 951 375 955
rect 379 951 380 955
rect 374 950 380 951
rect 450 955 456 956
rect 450 951 451 955
rect 455 951 456 955
rect 450 950 456 951
rect 470 955 476 956
rect 470 951 471 955
rect 475 951 476 955
rect 470 950 476 951
rect 478 955 484 956
rect 478 951 479 955
rect 483 951 484 955
rect 478 950 484 951
rect 566 955 572 956
rect 566 951 567 955
rect 571 951 572 955
rect 566 950 572 951
rect 650 955 656 956
rect 650 951 651 955
rect 655 951 656 955
rect 650 950 656 951
rect 670 955 676 956
rect 670 951 671 955
rect 675 951 676 955
rect 670 950 676 951
rect 690 955 696 956
rect 690 951 691 955
rect 695 951 696 955
rect 690 950 696 951
rect 766 955 772 956
rect 766 951 767 955
rect 771 951 772 955
rect 766 950 772 951
rect 834 955 840 956
rect 834 951 835 955
rect 839 951 840 955
rect 834 950 840 951
rect 854 955 860 956
rect 854 951 855 955
rect 859 951 860 955
rect 854 950 860 951
rect 922 955 928 956
rect 922 951 923 955
rect 927 951 928 955
rect 922 950 928 951
rect 942 955 948 956
rect 942 951 943 955
rect 947 951 948 955
rect 942 950 948 951
rect 1002 955 1008 956
rect 1002 951 1003 955
rect 1007 951 1008 955
rect 1002 950 1008 951
rect 1022 955 1028 956
rect 1022 951 1023 955
rect 1027 951 1028 955
rect 1022 950 1028 951
rect 1046 955 1052 956
rect 1046 951 1047 955
rect 1051 951 1052 955
rect 1046 950 1052 951
rect 1102 955 1108 956
rect 1102 951 1103 955
rect 1107 951 1108 955
rect 1102 950 1108 951
rect 1182 955 1188 956
rect 1182 951 1183 955
rect 1187 951 1188 955
rect 1182 950 1188 951
rect 356 936 358 950
rect 302 935 308 936
rect 302 931 303 935
rect 307 931 308 935
rect 302 930 308 931
rect 354 935 360 936
rect 354 931 355 935
rect 359 931 360 935
rect 354 930 360 931
rect 376 923 378 950
rect 452 936 454 950
rect 450 935 456 936
rect 450 931 451 935
rect 455 931 456 935
rect 450 930 456 931
rect 462 935 468 936
rect 462 931 463 935
rect 467 931 468 935
rect 462 930 468 931
rect 111 922 115 923
rect 111 917 115 918
rect 271 922 275 923
rect 271 917 275 918
rect 287 922 291 923
rect 287 917 291 918
rect 343 922 347 923
rect 343 917 347 918
rect 375 922 379 923
rect 375 917 379 918
rect 423 922 427 923
rect 423 917 427 918
rect 112 897 114 917
rect 272 898 274 917
rect 278 915 284 916
rect 278 911 279 915
rect 283 911 284 915
rect 278 910 284 911
rect 294 915 300 916
rect 294 911 295 915
rect 299 911 300 915
rect 294 910 300 911
rect 270 897 276 898
rect 110 896 116 897
rect 110 892 111 896
rect 115 892 116 896
rect 270 893 271 897
rect 275 893 276 897
rect 270 892 276 893
rect 110 891 116 892
rect 110 879 116 880
rect 110 875 111 879
rect 115 875 116 879
rect 110 874 116 875
rect 254 876 260 877
rect 112 867 114 874
rect 254 872 255 876
rect 259 872 260 876
rect 254 871 260 872
rect 256 867 258 871
rect 111 866 115 867
rect 111 861 115 862
rect 247 866 251 867
rect 247 861 251 862
rect 255 866 259 867
rect 255 861 259 862
rect 112 858 114 861
rect 246 860 252 861
rect 110 857 116 858
rect 110 853 111 857
rect 115 853 116 857
rect 246 856 247 860
rect 251 856 252 860
rect 246 855 252 856
rect 110 852 116 853
rect 110 840 116 841
rect 280 840 282 910
rect 296 896 298 910
rect 344 898 346 917
rect 424 898 426 917
rect 446 915 452 916
rect 446 911 447 915
rect 451 911 452 915
rect 446 910 452 911
rect 342 897 348 898
rect 294 895 300 896
rect 294 891 295 895
rect 299 891 300 895
rect 342 893 343 897
rect 347 893 348 897
rect 342 892 348 893
rect 422 897 428 898
rect 422 893 423 897
rect 427 893 428 897
rect 448 896 450 910
rect 464 904 466 930
rect 472 923 474 950
rect 480 924 482 950
rect 478 923 484 924
rect 568 923 570 950
rect 652 936 654 950
rect 650 935 656 936
rect 650 931 651 935
rect 655 931 656 935
rect 650 930 656 931
rect 672 923 674 950
rect 768 923 770 950
rect 836 936 838 950
rect 834 935 840 936
rect 834 931 835 935
rect 839 931 840 935
rect 834 930 840 931
rect 856 923 858 950
rect 924 936 926 950
rect 922 935 928 936
rect 922 931 923 935
rect 927 931 928 935
rect 922 930 928 931
rect 944 923 946 950
rect 1004 936 1006 950
rect 1002 935 1008 936
rect 1002 931 1003 935
rect 1007 931 1008 935
rect 1002 930 1008 931
rect 1024 923 1026 950
rect 1104 923 1106 950
rect 1184 923 1186 950
rect 1216 936 1218 1010
rect 1238 1009 1244 1010
rect 1288 1009 1290 1029
rect 1326 1027 1332 1028
rect 1326 1023 1327 1027
rect 1331 1023 1332 1027
rect 1326 1022 1332 1023
rect 1350 1024 1356 1025
rect 1328 1015 1330 1022
rect 1350 1020 1351 1024
rect 1355 1020 1356 1024
rect 1350 1019 1356 1020
rect 1438 1024 1444 1025
rect 1438 1020 1439 1024
rect 1443 1020 1444 1024
rect 1438 1019 1444 1020
rect 1558 1024 1564 1025
rect 1558 1020 1559 1024
rect 1563 1020 1564 1024
rect 1558 1019 1564 1020
rect 1678 1024 1684 1025
rect 1678 1020 1679 1024
rect 1683 1020 1684 1024
rect 1678 1019 1684 1020
rect 1352 1015 1354 1019
rect 1440 1015 1442 1019
rect 1560 1015 1562 1019
rect 1680 1015 1682 1019
rect 1327 1014 1331 1015
rect 1327 1009 1331 1010
rect 1351 1014 1355 1015
rect 1351 1009 1355 1010
rect 1439 1014 1443 1015
rect 1439 1009 1443 1010
rect 1511 1014 1515 1015
rect 1511 1009 1515 1010
rect 1559 1014 1563 1015
rect 1559 1009 1563 1010
rect 1679 1014 1683 1015
rect 1679 1009 1683 1010
rect 1238 1005 1239 1009
rect 1243 1005 1244 1009
rect 1286 1008 1292 1009
rect 1238 1004 1244 1005
rect 1278 1007 1284 1008
rect 1278 1003 1279 1007
rect 1283 1003 1284 1007
rect 1286 1004 1287 1008
rect 1291 1004 1292 1008
rect 1328 1006 1330 1009
rect 1350 1008 1356 1009
rect 1286 1003 1292 1004
rect 1326 1005 1332 1006
rect 1278 1002 1284 1003
rect 1222 988 1228 989
rect 1222 984 1223 988
rect 1227 984 1228 988
rect 1222 983 1228 984
rect 1223 982 1227 983
rect 1280 980 1282 1002
rect 1326 1001 1327 1005
rect 1331 1001 1332 1005
rect 1350 1004 1351 1008
rect 1355 1004 1356 1008
rect 1350 1003 1356 1004
rect 1510 1008 1516 1009
rect 1510 1004 1511 1008
rect 1515 1004 1516 1008
rect 1510 1003 1516 1004
rect 1678 1008 1684 1009
rect 1678 1004 1679 1008
rect 1683 1004 1684 1008
rect 1678 1003 1684 1004
rect 1326 1000 1332 1001
rect 1286 991 1292 992
rect 1286 987 1287 991
rect 1291 987 1292 991
rect 1286 986 1292 987
rect 1326 988 1332 989
rect 1712 988 1714 1050
rect 1720 1044 1722 1058
rect 1816 1046 1818 1065
rect 1814 1045 1820 1046
rect 1718 1043 1724 1044
rect 1718 1039 1719 1043
rect 1723 1039 1724 1043
rect 1814 1041 1815 1045
rect 1819 1041 1820 1045
rect 1836 1044 1838 1070
rect 1847 1065 1851 1066
rect 1927 1070 1931 1071
rect 1927 1065 1931 1066
rect 1999 1070 2003 1071
rect 1999 1065 2003 1066
rect 2039 1070 2043 1071
rect 2039 1065 2043 1066
rect 2071 1070 2075 1071
rect 2071 1065 2075 1066
rect 2151 1070 2155 1071
rect 2151 1065 2155 1066
rect 2231 1070 2235 1071
rect 2238 1067 2239 1071
rect 2243 1067 2244 1071
rect 2238 1066 2244 1067
rect 2255 1070 2259 1071
rect 2231 1065 2235 1066
rect 2255 1065 2259 1066
rect 2367 1070 2371 1071
rect 2367 1065 2371 1066
rect 2455 1070 2459 1071
rect 2455 1065 2459 1066
rect 1928 1046 1930 1065
rect 1950 1063 1956 1064
rect 1950 1059 1951 1063
rect 1955 1059 1956 1063
rect 1950 1058 1956 1059
rect 1926 1045 1932 1046
rect 1814 1040 1820 1041
rect 1834 1043 1840 1044
rect 1718 1038 1724 1039
rect 1834 1039 1835 1043
rect 1839 1039 1840 1043
rect 1926 1041 1927 1045
rect 1931 1041 1932 1045
rect 1952 1044 1954 1058
rect 2040 1046 2042 1065
rect 2062 1063 2068 1064
rect 2062 1059 2063 1063
rect 2067 1059 2068 1063
rect 2062 1058 2068 1059
rect 2038 1045 2044 1046
rect 1926 1040 1932 1041
rect 1950 1043 1956 1044
rect 1834 1038 1840 1039
rect 1950 1039 1951 1043
rect 1955 1039 1956 1043
rect 2038 1041 2039 1045
rect 2043 1041 2044 1045
rect 2064 1044 2066 1058
rect 2152 1046 2154 1065
rect 2174 1063 2180 1064
rect 2174 1059 2175 1063
rect 2179 1059 2180 1063
rect 2174 1058 2180 1059
rect 2150 1045 2156 1046
rect 2038 1040 2044 1041
rect 2062 1043 2068 1044
rect 1950 1038 1956 1039
rect 2062 1039 2063 1043
rect 2067 1039 2068 1043
rect 2150 1041 2151 1045
rect 2155 1041 2156 1045
rect 2176 1044 2178 1058
rect 2256 1046 2258 1065
rect 2278 1063 2284 1064
rect 2278 1059 2279 1063
rect 2283 1059 2284 1063
rect 2278 1058 2284 1059
rect 2254 1045 2260 1046
rect 2150 1040 2156 1041
rect 2174 1043 2180 1044
rect 2062 1038 2068 1039
rect 2174 1039 2175 1043
rect 2179 1039 2180 1043
rect 2254 1041 2255 1045
rect 2259 1041 2260 1045
rect 2280 1044 2282 1058
rect 2368 1046 2370 1065
rect 2456 1046 2458 1065
rect 2464 1064 2466 1150
rect 2462 1063 2468 1064
rect 2462 1059 2463 1063
rect 2467 1059 2468 1063
rect 2462 1058 2468 1059
rect 2366 1045 2372 1046
rect 2254 1040 2260 1041
rect 2278 1043 2284 1044
rect 2174 1038 2180 1039
rect 2278 1039 2279 1043
rect 2283 1039 2284 1043
rect 2366 1041 2367 1045
rect 2371 1041 2372 1045
rect 2454 1045 2460 1046
rect 2366 1040 2372 1041
rect 2374 1043 2380 1044
rect 2278 1038 2284 1039
rect 2374 1039 2375 1043
rect 2379 1039 2380 1043
rect 2454 1041 2455 1045
rect 2459 1041 2460 1045
rect 2454 1040 2460 1041
rect 2462 1043 2468 1044
rect 2374 1038 2380 1039
rect 2462 1039 2463 1043
rect 2467 1039 2468 1043
rect 2462 1038 2468 1039
rect 1798 1024 1804 1025
rect 1798 1020 1799 1024
rect 1803 1020 1804 1024
rect 1798 1019 1804 1020
rect 1910 1024 1916 1025
rect 1910 1020 1911 1024
rect 1915 1020 1916 1024
rect 1910 1019 1916 1020
rect 2022 1024 2028 1025
rect 2022 1020 2023 1024
rect 2027 1020 2028 1024
rect 2022 1019 2028 1020
rect 2134 1024 2140 1025
rect 2134 1020 2135 1024
rect 2139 1020 2140 1024
rect 2134 1019 2140 1020
rect 2238 1024 2244 1025
rect 2238 1020 2239 1024
rect 2243 1020 2244 1024
rect 2238 1019 2244 1020
rect 2350 1024 2356 1025
rect 2350 1020 2351 1024
rect 2355 1020 2356 1024
rect 2350 1019 2356 1020
rect 1800 1015 1802 1019
rect 1912 1015 1914 1019
rect 2024 1015 2026 1019
rect 2136 1015 2138 1019
rect 2240 1015 2242 1019
rect 2352 1015 2354 1019
rect 1799 1014 1803 1015
rect 1799 1009 1803 1010
rect 1823 1014 1827 1015
rect 1823 1009 1827 1010
rect 1911 1014 1915 1015
rect 1911 1009 1915 1010
rect 1951 1014 1955 1015
rect 1951 1009 1955 1010
rect 2023 1014 2027 1015
rect 2023 1009 2027 1010
rect 2071 1014 2075 1015
rect 2071 1009 2075 1010
rect 2135 1014 2139 1015
rect 2135 1009 2139 1010
rect 2175 1014 2179 1015
rect 2175 1009 2179 1010
rect 2239 1014 2243 1015
rect 2239 1009 2243 1010
rect 2271 1014 2275 1015
rect 2271 1009 2275 1010
rect 2351 1014 2355 1015
rect 2351 1009 2355 1010
rect 2367 1014 2371 1015
rect 2367 1009 2371 1010
rect 1822 1008 1828 1009
rect 1822 1004 1823 1008
rect 1827 1004 1828 1008
rect 1822 1003 1828 1004
rect 1950 1008 1956 1009
rect 1950 1004 1951 1008
rect 1955 1004 1956 1008
rect 1950 1003 1956 1004
rect 2070 1008 2076 1009
rect 2070 1004 2071 1008
rect 2075 1004 2076 1008
rect 2070 1003 2076 1004
rect 2174 1008 2180 1009
rect 2174 1004 2175 1008
rect 2179 1004 2180 1008
rect 2174 1003 2180 1004
rect 2270 1008 2276 1009
rect 2270 1004 2271 1008
rect 2275 1004 2276 1008
rect 2270 1003 2276 1004
rect 2366 1008 2372 1009
rect 2366 1004 2367 1008
rect 2371 1004 2372 1008
rect 2366 1003 2372 1004
rect 1288 983 1290 986
rect 1326 984 1327 988
rect 1331 984 1332 988
rect 1326 983 1332 984
rect 1366 987 1372 988
rect 1366 983 1367 987
rect 1371 983 1372 987
rect 1287 982 1291 983
rect 1223 977 1227 978
rect 1278 979 1284 980
rect 1222 976 1228 977
rect 1222 972 1223 976
rect 1227 972 1228 976
rect 1278 975 1279 979
rect 1283 975 1284 979
rect 1287 977 1291 978
rect 1278 974 1284 975
rect 1288 974 1290 977
rect 1222 971 1228 972
rect 1286 973 1292 974
rect 1286 969 1287 973
rect 1291 969 1292 973
rect 1286 968 1292 969
rect 1286 956 1292 957
rect 1238 955 1244 956
rect 1238 951 1239 955
rect 1243 951 1244 955
rect 1286 952 1287 956
rect 1291 952 1292 956
rect 1286 951 1292 952
rect 1328 951 1330 983
rect 1366 982 1372 983
rect 1374 987 1380 988
rect 1374 983 1375 987
rect 1379 983 1380 987
rect 1374 982 1380 983
rect 1526 987 1532 988
rect 1526 983 1527 987
rect 1531 983 1532 987
rect 1526 982 1532 983
rect 1674 987 1680 988
rect 1674 983 1675 987
rect 1679 983 1680 987
rect 1674 982 1680 983
rect 1694 987 1700 988
rect 1694 983 1695 987
rect 1699 983 1700 987
rect 1694 982 1700 983
rect 1710 987 1716 988
rect 1710 983 1711 987
rect 1715 983 1716 987
rect 1710 982 1716 983
rect 1838 987 1844 988
rect 1838 983 1839 987
rect 1843 983 1844 987
rect 1838 982 1844 983
rect 1946 987 1952 988
rect 1946 983 1947 987
rect 1951 983 1952 987
rect 1946 982 1952 983
rect 1966 987 1972 988
rect 1966 983 1967 987
rect 1971 983 1972 987
rect 1966 982 1972 983
rect 2066 987 2072 988
rect 2066 983 2067 987
rect 2071 983 2072 987
rect 2066 982 2072 983
rect 2086 987 2092 988
rect 2086 983 2087 987
rect 2091 983 2092 987
rect 2086 982 2092 983
rect 2170 987 2176 988
rect 2170 983 2171 987
rect 2175 983 2176 987
rect 2170 982 2176 983
rect 2190 987 2196 988
rect 2190 983 2191 987
rect 2195 983 2196 987
rect 2190 982 2196 983
rect 2266 987 2272 988
rect 2266 983 2267 987
rect 2271 983 2272 987
rect 2266 982 2272 983
rect 2286 987 2292 988
rect 2286 983 2287 987
rect 2291 983 2292 987
rect 2286 982 2292 983
rect 2362 987 2368 988
rect 2362 983 2363 987
rect 2367 983 2368 987
rect 2362 982 2368 983
rect 1368 951 1370 982
rect 1238 950 1244 951
rect 1202 935 1208 936
rect 1202 931 1203 935
rect 1207 931 1208 935
rect 1202 930 1208 931
rect 1214 935 1220 936
rect 1214 931 1215 935
rect 1219 931 1220 935
rect 1214 930 1220 931
rect 471 922 475 923
rect 478 919 479 923
rect 483 919 484 923
rect 478 918 484 919
rect 519 922 523 923
rect 471 917 475 918
rect 519 917 523 918
rect 567 922 571 923
rect 567 917 571 918
rect 615 922 619 923
rect 615 917 619 918
rect 671 922 675 923
rect 671 917 675 918
rect 711 922 715 923
rect 711 917 715 918
rect 767 922 771 923
rect 767 917 771 918
rect 807 922 811 923
rect 807 917 811 918
rect 855 922 859 923
rect 855 917 859 918
rect 903 922 907 923
rect 903 917 907 918
rect 943 922 947 923
rect 943 917 947 918
rect 991 922 995 923
rect 991 917 995 918
rect 1023 922 1027 923
rect 1023 917 1027 918
rect 1087 922 1091 923
rect 1087 917 1091 918
rect 1103 922 1107 923
rect 1103 917 1107 918
rect 1183 922 1187 923
rect 1183 917 1187 918
rect 462 903 468 904
rect 462 899 463 903
rect 467 899 468 903
rect 462 898 468 899
rect 520 898 522 917
rect 542 915 548 916
rect 542 911 543 915
rect 547 911 548 915
rect 542 910 548 911
rect 518 897 524 898
rect 422 892 428 893
rect 446 895 452 896
rect 294 890 300 891
rect 446 891 447 895
rect 451 891 452 895
rect 518 893 519 897
rect 523 893 524 897
rect 544 896 546 910
rect 616 898 618 917
rect 638 915 644 916
rect 638 911 639 915
rect 643 911 644 915
rect 638 910 644 911
rect 614 897 620 898
rect 518 892 524 893
rect 542 895 548 896
rect 446 890 452 891
rect 542 891 543 895
rect 547 891 548 895
rect 614 893 615 897
rect 619 893 620 897
rect 640 896 642 910
rect 712 898 714 917
rect 808 898 810 917
rect 830 915 836 916
rect 830 911 831 915
rect 835 911 836 915
rect 830 910 836 911
rect 710 897 716 898
rect 614 892 620 893
rect 638 895 644 896
rect 542 890 548 891
rect 638 891 639 895
rect 643 891 644 895
rect 710 893 711 897
rect 715 893 716 897
rect 806 897 812 898
rect 710 892 716 893
rect 718 895 724 896
rect 638 890 644 891
rect 718 891 719 895
rect 723 891 724 895
rect 806 893 807 897
rect 811 893 812 897
rect 832 896 834 910
rect 904 898 906 917
rect 926 915 932 916
rect 926 911 927 915
rect 931 911 932 915
rect 926 910 932 911
rect 902 897 908 898
rect 806 892 812 893
rect 830 895 836 896
rect 718 890 724 891
rect 830 891 831 895
rect 835 891 836 895
rect 902 893 903 897
rect 907 893 908 897
rect 928 896 930 910
rect 938 907 944 908
rect 938 903 939 907
rect 943 903 944 907
rect 938 902 944 903
rect 902 892 908 893
rect 926 895 932 896
rect 830 890 836 891
rect 926 891 927 895
rect 931 891 932 895
rect 926 890 932 891
rect 326 876 332 877
rect 326 872 327 876
rect 331 872 332 876
rect 326 871 332 872
rect 406 876 412 877
rect 406 872 407 876
rect 411 872 412 876
rect 406 871 412 872
rect 502 876 508 877
rect 502 872 503 876
rect 507 872 508 876
rect 502 871 508 872
rect 598 876 604 877
rect 598 872 599 876
rect 603 872 604 876
rect 598 871 604 872
rect 694 876 700 877
rect 694 872 695 876
rect 699 872 700 876
rect 694 871 700 872
rect 328 867 330 871
rect 408 867 410 871
rect 504 867 506 871
rect 600 867 602 871
rect 696 867 698 871
rect 311 866 315 867
rect 311 861 315 862
rect 327 866 331 867
rect 327 861 331 862
rect 375 866 379 867
rect 375 861 379 862
rect 407 866 411 867
rect 407 861 411 862
rect 439 866 443 867
rect 439 861 443 862
rect 503 866 507 867
rect 503 861 507 862
rect 567 866 571 867
rect 567 861 571 862
rect 599 866 603 867
rect 599 861 603 862
rect 631 866 635 867
rect 631 861 635 862
rect 695 866 699 867
rect 695 861 699 862
rect 310 860 316 861
rect 310 856 311 860
rect 315 856 316 860
rect 310 855 316 856
rect 374 860 380 861
rect 374 856 375 860
rect 379 856 380 860
rect 374 855 380 856
rect 438 860 444 861
rect 438 856 439 860
rect 443 856 444 860
rect 438 855 444 856
rect 502 860 508 861
rect 502 856 503 860
rect 507 856 508 860
rect 502 855 508 856
rect 566 860 572 861
rect 566 856 567 860
rect 571 856 572 860
rect 566 855 572 856
rect 630 860 636 861
rect 630 856 631 860
rect 635 856 636 860
rect 630 855 636 856
rect 694 860 700 861
rect 694 856 695 860
rect 699 856 700 860
rect 694 855 700 856
rect 110 836 111 840
rect 115 836 116 840
rect 110 835 116 836
rect 262 839 268 840
rect 262 835 263 839
rect 267 835 268 839
rect 112 811 114 835
rect 262 834 268 835
rect 278 839 284 840
rect 278 835 279 839
rect 283 835 284 839
rect 278 834 284 835
rect 326 839 332 840
rect 326 835 327 839
rect 331 835 332 839
rect 326 834 332 835
rect 390 839 396 840
rect 390 835 391 839
rect 395 835 396 839
rect 390 834 396 835
rect 434 839 440 840
rect 434 835 435 839
rect 439 835 440 839
rect 434 834 440 835
rect 454 839 460 840
rect 454 835 455 839
rect 459 835 460 839
rect 454 834 460 835
rect 498 839 504 840
rect 498 835 499 839
rect 503 835 504 839
rect 498 834 504 835
rect 518 839 524 840
rect 518 835 519 839
rect 523 835 524 839
rect 518 834 524 835
rect 562 839 568 840
rect 562 835 563 839
rect 567 835 568 839
rect 562 834 568 835
rect 582 839 588 840
rect 582 835 583 839
rect 587 835 588 839
rect 582 834 588 835
rect 590 839 596 840
rect 590 835 591 839
rect 595 835 596 839
rect 590 834 596 835
rect 646 839 652 840
rect 646 835 647 839
rect 651 835 652 839
rect 646 834 652 835
rect 690 839 696 840
rect 690 835 691 839
rect 695 835 696 839
rect 690 834 696 835
rect 710 839 716 840
rect 710 835 711 839
rect 715 835 716 839
rect 710 834 716 835
rect 264 811 266 834
rect 318 819 324 820
rect 318 815 319 819
rect 323 815 324 819
rect 318 814 324 815
rect 111 810 115 811
rect 111 805 115 806
rect 215 810 219 811
rect 215 805 219 806
rect 263 810 267 811
rect 263 805 267 806
rect 303 810 307 811
rect 303 805 307 806
rect 112 785 114 805
rect 174 803 180 804
rect 174 799 175 803
rect 179 799 180 803
rect 174 798 180 799
rect 110 784 116 785
rect 110 780 111 784
rect 115 780 116 784
rect 110 779 116 780
rect 110 767 116 768
rect 110 763 111 767
rect 115 763 116 767
rect 110 762 116 763
rect 112 759 114 762
rect 111 758 115 759
rect 111 753 115 754
rect 135 758 139 759
rect 135 753 139 754
rect 112 750 114 753
rect 134 752 140 753
rect 110 749 116 750
rect 110 745 111 749
rect 115 745 116 749
rect 134 748 135 752
rect 139 748 140 752
rect 134 747 140 748
rect 110 744 116 745
rect 110 732 116 733
rect 176 732 178 798
rect 216 786 218 805
rect 238 803 244 804
rect 238 799 239 803
rect 243 799 244 803
rect 238 798 244 799
rect 214 785 220 786
rect 214 781 215 785
rect 219 781 220 785
rect 240 784 242 798
rect 304 786 306 805
rect 302 785 308 786
rect 214 780 220 781
rect 238 783 244 784
rect 238 779 239 783
rect 243 779 244 783
rect 302 781 303 785
rect 307 781 308 785
rect 320 784 322 814
rect 328 811 330 834
rect 392 811 394 834
rect 436 820 438 834
rect 434 819 440 820
rect 434 815 435 819
rect 439 815 440 819
rect 434 814 440 815
rect 456 811 458 834
rect 500 820 502 834
rect 498 819 504 820
rect 498 815 499 819
rect 503 815 504 819
rect 498 814 504 815
rect 520 811 522 834
rect 564 820 566 834
rect 562 819 568 820
rect 562 815 563 819
rect 567 815 568 819
rect 562 814 568 815
rect 584 811 586 834
rect 592 812 594 834
rect 590 811 596 812
rect 648 811 650 834
rect 692 820 694 834
rect 682 819 688 820
rect 682 815 683 819
rect 687 815 688 819
rect 682 814 688 815
rect 690 819 696 820
rect 690 815 691 819
rect 695 815 696 819
rect 690 814 696 815
rect 327 810 331 811
rect 327 805 331 806
rect 391 810 395 811
rect 391 805 395 806
rect 455 810 459 811
rect 455 805 459 806
rect 479 810 483 811
rect 479 805 483 806
rect 519 810 523 811
rect 519 805 523 806
rect 559 810 563 811
rect 559 805 563 806
rect 583 810 587 811
rect 590 807 591 811
rect 595 807 596 811
rect 590 806 596 807
rect 631 810 635 811
rect 583 805 587 806
rect 631 805 635 806
rect 647 810 651 811
rect 647 805 651 806
rect 392 786 394 805
rect 414 803 420 804
rect 414 799 415 803
rect 419 799 420 803
rect 414 798 420 799
rect 390 785 396 786
rect 302 780 308 781
rect 318 783 324 784
rect 238 778 244 779
rect 318 779 319 783
rect 323 779 324 783
rect 390 781 391 785
rect 395 781 396 785
rect 416 784 418 798
rect 480 786 482 805
rect 502 803 508 804
rect 502 799 503 803
rect 507 799 508 803
rect 502 798 508 799
rect 478 785 484 786
rect 390 780 396 781
rect 414 783 420 784
rect 318 778 324 779
rect 414 779 415 783
rect 419 779 420 783
rect 478 781 479 785
rect 483 781 484 785
rect 504 784 506 798
rect 560 786 562 805
rect 590 803 596 804
rect 590 799 591 803
rect 595 799 596 803
rect 590 798 596 799
rect 558 785 564 786
rect 478 780 484 781
rect 502 783 508 784
rect 414 778 420 779
rect 502 779 503 783
rect 507 779 508 783
rect 558 781 559 785
rect 563 781 564 785
rect 592 784 594 798
rect 632 786 634 805
rect 654 803 660 804
rect 654 799 655 803
rect 659 799 660 803
rect 654 798 660 799
rect 630 785 636 786
rect 558 780 564 781
rect 590 783 596 784
rect 502 778 508 779
rect 590 779 591 783
rect 595 779 596 783
rect 630 781 631 785
rect 635 781 636 785
rect 656 784 658 798
rect 684 792 686 814
rect 712 811 714 834
rect 720 828 722 890
rect 790 876 796 877
rect 790 872 791 876
rect 795 872 796 876
rect 790 871 796 872
rect 886 876 892 877
rect 886 872 887 876
rect 891 872 892 876
rect 886 871 892 872
rect 792 867 794 871
rect 888 867 890 871
rect 759 866 763 867
rect 759 861 763 862
rect 791 866 795 867
rect 791 861 795 862
rect 831 866 835 867
rect 831 861 835 862
rect 887 866 891 867
rect 887 861 891 862
rect 903 866 907 867
rect 903 861 907 862
rect 758 860 764 861
rect 758 856 759 860
rect 763 856 764 860
rect 758 855 764 856
rect 830 860 836 861
rect 830 856 831 860
rect 835 856 836 860
rect 830 855 836 856
rect 902 860 908 861
rect 902 856 903 860
rect 907 856 908 860
rect 902 855 908 856
rect 940 840 942 902
rect 992 898 994 917
rect 1014 915 1020 916
rect 1014 911 1015 915
rect 1019 911 1020 915
rect 1014 910 1020 911
rect 990 897 996 898
rect 990 893 991 897
rect 995 893 996 897
rect 1016 896 1018 910
rect 1088 898 1090 917
rect 1184 898 1186 917
rect 1086 897 1092 898
rect 990 892 996 893
rect 1014 895 1020 896
rect 1014 891 1015 895
rect 1019 891 1020 895
rect 1086 893 1087 897
rect 1091 893 1092 897
rect 1086 892 1092 893
rect 1182 897 1188 898
rect 1182 893 1183 897
rect 1187 893 1188 897
rect 1204 896 1206 930
rect 1240 923 1242 950
rect 1288 923 1290 951
rect 1327 950 1331 951
rect 1327 945 1331 946
rect 1367 950 1371 951
rect 1367 945 1371 946
rect 1328 925 1330 945
rect 1368 926 1370 945
rect 1376 944 1378 982
rect 1528 951 1530 982
rect 1676 968 1678 982
rect 1674 967 1680 968
rect 1674 963 1675 967
rect 1679 963 1680 967
rect 1674 962 1680 963
rect 1696 951 1698 982
rect 1823 972 1827 973
rect 1822 967 1828 968
rect 1822 963 1823 967
rect 1827 963 1828 967
rect 1822 962 1828 963
rect 1840 951 1842 982
rect 1948 968 1950 982
rect 1946 967 1952 968
rect 1946 963 1947 967
rect 1951 963 1952 967
rect 1946 962 1952 963
rect 1968 951 1970 982
rect 2068 968 2070 982
rect 2066 967 2072 968
rect 2066 963 2067 967
rect 2071 963 2072 967
rect 2066 962 2072 963
rect 2088 951 2090 982
rect 2172 968 2174 982
rect 2170 967 2176 968
rect 2170 963 2171 967
rect 2175 963 2176 967
rect 2170 962 2176 963
rect 2192 951 2194 982
rect 2268 968 2270 982
rect 2266 967 2272 968
rect 2266 963 2267 967
rect 2271 963 2272 967
rect 2266 962 2272 963
rect 2288 951 2290 982
rect 2364 968 2366 982
rect 2376 973 2378 1038
rect 2438 1024 2444 1025
rect 2438 1020 2439 1024
rect 2443 1020 2444 1024
rect 2438 1019 2444 1020
rect 2440 1015 2442 1019
rect 2439 1014 2443 1015
rect 2439 1009 2443 1010
rect 2438 1008 2444 1009
rect 2438 1004 2439 1008
rect 2443 1004 2444 1008
rect 2438 1003 2444 1004
rect 2382 987 2388 988
rect 2382 983 2383 987
rect 2387 983 2388 987
rect 2382 982 2388 983
rect 2390 987 2396 988
rect 2390 983 2391 987
rect 2395 983 2396 987
rect 2390 982 2396 983
rect 2454 987 2460 988
rect 2454 983 2455 987
rect 2459 983 2460 987
rect 2454 982 2460 983
rect 2375 972 2379 973
rect 2362 967 2368 968
rect 2375 967 2379 968
rect 2362 963 2363 967
rect 2367 963 2368 967
rect 2362 962 2368 963
rect 2384 951 2386 982
rect 1423 950 1427 951
rect 1423 945 1427 946
rect 1503 950 1507 951
rect 1503 945 1507 946
rect 1527 950 1531 951
rect 1527 945 1531 946
rect 1607 950 1611 951
rect 1607 945 1611 946
rect 1695 950 1699 951
rect 1695 945 1699 946
rect 1719 950 1723 951
rect 1719 945 1723 946
rect 1831 950 1835 951
rect 1831 945 1835 946
rect 1839 950 1843 951
rect 1839 945 1843 946
rect 1935 950 1939 951
rect 1935 945 1939 946
rect 1967 950 1971 951
rect 1967 945 1971 946
rect 2031 950 2035 951
rect 2031 945 2035 946
rect 2087 950 2091 951
rect 2087 945 2091 946
rect 2127 950 2131 951
rect 2127 945 2131 946
rect 2191 950 2195 951
rect 2191 945 2195 946
rect 2215 950 2219 951
rect 2215 945 2219 946
rect 2287 950 2291 951
rect 2287 945 2291 946
rect 2295 950 2299 951
rect 2295 945 2299 946
rect 2375 950 2379 951
rect 2375 945 2379 946
rect 2383 950 2387 951
rect 2383 945 2387 946
rect 1374 943 1380 944
rect 1374 939 1375 943
rect 1379 939 1380 943
rect 1374 938 1380 939
rect 1390 943 1396 944
rect 1390 939 1391 943
rect 1395 939 1396 943
rect 1390 938 1396 939
rect 1366 925 1372 926
rect 1326 924 1332 925
rect 1239 922 1243 923
rect 1239 917 1243 918
rect 1287 922 1291 923
rect 1326 920 1327 924
rect 1331 920 1332 924
rect 1366 921 1367 925
rect 1371 921 1372 925
rect 1392 924 1394 938
rect 1424 926 1426 945
rect 1446 943 1452 944
rect 1446 939 1447 943
rect 1451 939 1452 943
rect 1446 938 1452 939
rect 1438 931 1444 932
rect 1438 927 1439 931
rect 1443 927 1444 931
rect 1438 926 1444 927
rect 1422 925 1428 926
rect 1366 920 1372 921
rect 1390 923 1396 924
rect 1326 919 1332 920
rect 1390 919 1391 923
rect 1395 919 1396 923
rect 1422 921 1423 925
rect 1427 921 1428 925
rect 1422 920 1428 921
rect 1390 918 1396 919
rect 1287 917 1291 918
rect 1288 897 1290 917
rect 1326 907 1332 908
rect 1326 903 1327 907
rect 1331 903 1332 907
rect 1326 902 1332 903
rect 1350 904 1356 905
rect 1286 896 1292 897
rect 1182 892 1188 893
rect 1202 895 1208 896
rect 1014 890 1020 891
rect 1202 891 1203 895
rect 1207 891 1208 895
rect 1286 892 1287 896
rect 1291 892 1292 896
rect 1328 895 1330 902
rect 1350 900 1351 904
rect 1355 900 1356 904
rect 1350 899 1356 900
rect 1406 904 1412 905
rect 1406 900 1407 904
rect 1411 900 1412 904
rect 1406 899 1412 900
rect 1352 895 1354 899
rect 1408 895 1410 899
rect 1286 891 1292 892
rect 1327 894 1331 895
rect 1202 890 1208 891
rect 1327 889 1331 890
rect 1351 894 1355 895
rect 1351 889 1355 890
rect 1407 894 1411 895
rect 1407 889 1411 890
rect 1431 894 1435 895
rect 1431 889 1435 890
rect 1328 886 1330 889
rect 1430 888 1436 889
rect 1326 885 1332 886
rect 1326 881 1327 885
rect 1331 881 1332 885
rect 1430 884 1431 888
rect 1435 884 1436 888
rect 1430 883 1436 884
rect 1326 880 1332 881
rect 1286 879 1292 880
rect 974 876 980 877
rect 974 872 975 876
rect 979 872 980 876
rect 974 871 980 872
rect 1070 876 1076 877
rect 1070 872 1071 876
rect 1075 872 1076 876
rect 1070 871 1076 872
rect 1166 876 1172 877
rect 1166 872 1167 876
rect 1171 872 1172 876
rect 1286 875 1287 879
rect 1291 875 1292 879
rect 1286 874 1292 875
rect 1166 871 1172 872
rect 976 867 978 871
rect 1072 867 1074 871
rect 1168 867 1170 871
rect 1288 867 1290 874
rect 1326 868 1332 869
rect 975 866 979 867
rect 975 861 979 862
rect 1071 866 1075 867
rect 1071 861 1075 862
rect 1167 866 1171 867
rect 1167 861 1171 862
rect 1287 866 1291 867
rect 1326 864 1327 868
rect 1331 864 1332 868
rect 1326 863 1332 864
rect 1287 861 1291 862
rect 1288 858 1290 861
rect 1286 857 1292 858
rect 1286 853 1287 857
rect 1291 853 1292 857
rect 1286 852 1292 853
rect 1286 840 1292 841
rect 754 839 760 840
rect 754 835 755 839
rect 759 835 760 839
rect 754 834 760 835
rect 774 839 780 840
rect 774 835 775 839
rect 779 835 780 839
rect 774 834 780 835
rect 826 839 832 840
rect 826 835 827 839
rect 831 835 832 839
rect 826 834 832 835
rect 846 839 852 840
rect 846 835 847 839
rect 851 835 852 839
rect 846 834 852 835
rect 898 839 904 840
rect 898 835 899 839
rect 903 835 904 839
rect 898 834 904 835
rect 918 839 924 840
rect 918 835 919 839
rect 923 835 924 839
rect 918 834 924 835
rect 938 839 944 840
rect 938 835 939 839
rect 943 835 944 839
rect 1286 836 1287 840
rect 1291 836 1292 840
rect 1328 839 1330 863
rect 1440 848 1442 926
rect 1448 924 1450 938
rect 1504 926 1506 945
rect 1534 943 1540 944
rect 1534 939 1535 943
rect 1539 939 1540 943
rect 1534 938 1540 939
rect 1502 925 1508 926
rect 1446 923 1452 924
rect 1446 919 1447 923
rect 1451 919 1452 923
rect 1502 921 1503 925
rect 1507 921 1508 925
rect 1536 924 1538 938
rect 1608 926 1610 945
rect 1630 943 1636 944
rect 1630 939 1631 943
rect 1635 939 1636 943
rect 1630 938 1636 939
rect 1606 925 1612 926
rect 1502 920 1508 921
rect 1534 923 1540 924
rect 1446 918 1452 919
rect 1534 919 1535 923
rect 1539 919 1540 923
rect 1606 921 1607 925
rect 1611 921 1612 925
rect 1632 924 1634 938
rect 1720 926 1722 945
rect 1742 943 1748 944
rect 1742 939 1743 943
rect 1747 939 1748 943
rect 1742 938 1748 939
rect 1718 925 1724 926
rect 1606 920 1612 921
rect 1630 923 1636 924
rect 1534 918 1540 919
rect 1630 919 1631 923
rect 1635 919 1636 923
rect 1718 921 1719 925
rect 1723 921 1724 925
rect 1744 924 1746 938
rect 1832 926 1834 945
rect 1936 926 1938 945
rect 1958 943 1964 944
rect 1958 939 1959 943
rect 1963 939 1964 943
rect 1958 938 1964 939
rect 1830 925 1836 926
rect 1718 920 1724 921
rect 1742 923 1748 924
rect 1630 918 1636 919
rect 1742 919 1743 923
rect 1747 919 1748 923
rect 1830 921 1831 925
rect 1835 921 1836 925
rect 1830 920 1836 921
rect 1934 925 1940 926
rect 1934 921 1935 925
rect 1939 921 1940 925
rect 1960 924 1962 938
rect 2032 926 2034 945
rect 2054 943 2060 944
rect 2054 939 2055 943
rect 2059 939 2060 943
rect 2054 938 2060 939
rect 2030 925 2036 926
rect 1934 920 1940 921
rect 1958 923 1964 924
rect 1742 918 1748 919
rect 1958 919 1959 923
rect 1963 919 1964 923
rect 2030 921 2031 925
rect 2035 921 2036 925
rect 2056 924 2058 938
rect 2128 926 2130 945
rect 2216 926 2218 945
rect 2296 926 2298 945
rect 2376 926 2378 945
rect 2392 944 2394 982
rect 2446 967 2452 968
rect 2446 963 2447 967
rect 2451 963 2452 967
rect 2446 962 2452 963
rect 2390 943 2396 944
rect 2390 939 2391 943
rect 2395 939 2396 943
rect 2390 938 2396 939
rect 2126 925 2132 926
rect 2030 920 2036 921
rect 2054 923 2060 924
rect 1958 918 1964 919
rect 2054 919 2055 923
rect 2059 919 2060 923
rect 2126 921 2127 925
rect 2131 921 2132 925
rect 2214 925 2220 926
rect 2126 920 2132 921
rect 2150 923 2156 924
rect 2054 918 2060 919
rect 2150 919 2151 923
rect 2155 919 2156 923
rect 2214 921 2215 925
rect 2219 921 2220 925
rect 2214 920 2220 921
rect 2294 925 2300 926
rect 2294 921 2295 925
rect 2299 921 2300 925
rect 2294 920 2300 921
rect 2374 925 2380 926
rect 2374 921 2375 925
rect 2379 921 2380 925
rect 2374 920 2380 921
rect 2150 918 2156 919
rect 1486 904 1492 905
rect 1486 900 1487 904
rect 1491 900 1492 904
rect 1486 899 1492 900
rect 1590 904 1596 905
rect 1590 900 1591 904
rect 1595 900 1596 904
rect 1590 899 1596 900
rect 1702 904 1708 905
rect 1702 900 1703 904
rect 1707 900 1708 904
rect 1702 899 1708 900
rect 1814 904 1820 905
rect 1814 900 1815 904
rect 1819 900 1820 904
rect 1814 899 1820 900
rect 1918 904 1924 905
rect 1918 900 1919 904
rect 1923 900 1924 904
rect 1918 899 1924 900
rect 2014 904 2020 905
rect 2014 900 2015 904
rect 2019 900 2020 904
rect 2014 899 2020 900
rect 2110 904 2116 905
rect 2110 900 2111 904
rect 2115 900 2116 904
rect 2110 899 2116 900
rect 1488 895 1490 899
rect 1592 895 1594 899
rect 1704 895 1706 899
rect 1816 895 1818 899
rect 1920 895 1922 899
rect 2016 895 2018 899
rect 2112 895 2114 899
rect 1487 894 1491 895
rect 1487 889 1491 890
rect 1551 894 1555 895
rect 1551 889 1555 890
rect 1591 894 1595 895
rect 1591 889 1595 890
rect 1623 894 1627 895
rect 1623 889 1627 890
rect 1703 894 1707 895
rect 1703 889 1707 890
rect 1791 894 1795 895
rect 1791 889 1795 890
rect 1815 894 1819 895
rect 1815 889 1819 890
rect 1895 894 1899 895
rect 1895 889 1899 890
rect 1919 894 1923 895
rect 1919 889 1923 890
rect 2015 894 2019 895
rect 2015 889 2019 890
rect 2111 894 2115 895
rect 2111 889 2115 890
rect 2143 894 2147 895
rect 2143 889 2147 890
rect 1486 888 1492 889
rect 1486 884 1487 888
rect 1491 884 1492 888
rect 1486 883 1492 884
rect 1550 888 1556 889
rect 1550 884 1551 888
rect 1555 884 1556 888
rect 1550 883 1556 884
rect 1622 888 1628 889
rect 1622 884 1623 888
rect 1627 884 1628 888
rect 1622 883 1628 884
rect 1702 888 1708 889
rect 1702 884 1703 888
rect 1707 884 1708 888
rect 1702 883 1708 884
rect 1790 888 1796 889
rect 1790 884 1791 888
rect 1795 884 1796 888
rect 1790 883 1796 884
rect 1894 888 1900 889
rect 1894 884 1895 888
rect 1899 884 1900 888
rect 1894 883 1900 884
rect 2014 888 2020 889
rect 2014 884 2015 888
rect 2019 884 2020 888
rect 2014 883 2020 884
rect 2142 888 2148 889
rect 2142 884 2143 888
rect 2147 884 2148 888
rect 2142 883 2148 884
rect 1446 867 1452 868
rect 1446 863 1447 867
rect 1451 863 1452 867
rect 1446 862 1452 863
rect 1482 867 1488 868
rect 1482 863 1483 867
rect 1487 863 1488 867
rect 1482 862 1488 863
rect 1502 867 1508 868
rect 1502 863 1503 867
rect 1507 863 1508 867
rect 1502 862 1508 863
rect 1546 867 1552 868
rect 1546 863 1547 867
rect 1551 863 1552 867
rect 1546 862 1552 863
rect 1566 867 1572 868
rect 1566 863 1567 867
rect 1571 863 1572 867
rect 1566 862 1572 863
rect 1618 867 1624 868
rect 1618 863 1619 867
rect 1623 863 1624 867
rect 1618 862 1624 863
rect 1638 867 1644 868
rect 1638 863 1639 867
rect 1643 863 1644 867
rect 1638 862 1644 863
rect 1698 867 1704 868
rect 1698 863 1699 867
rect 1703 863 1704 867
rect 1698 862 1704 863
rect 1718 867 1724 868
rect 1718 863 1719 867
rect 1723 863 1724 867
rect 1718 862 1724 863
rect 1726 867 1732 868
rect 1726 863 1727 867
rect 1731 863 1732 867
rect 1726 862 1732 863
rect 1806 867 1812 868
rect 1806 863 1807 867
rect 1811 863 1812 867
rect 1806 862 1812 863
rect 1890 867 1896 868
rect 1890 863 1891 867
rect 1895 863 1896 867
rect 1890 862 1896 863
rect 1910 867 1916 868
rect 1910 863 1911 867
rect 1915 863 1916 867
rect 1910 862 1916 863
rect 1918 867 1924 868
rect 1918 863 1919 867
rect 1923 863 1924 867
rect 1918 862 1924 863
rect 2030 867 2036 868
rect 2030 863 2031 867
rect 2035 863 2036 867
rect 2030 862 2036 863
rect 1438 847 1444 848
rect 1438 843 1439 847
rect 1443 843 1444 847
rect 1438 842 1444 843
rect 1448 839 1450 862
rect 1484 848 1486 862
rect 1482 847 1488 848
rect 1482 843 1483 847
rect 1487 843 1488 847
rect 1482 842 1488 843
rect 1504 839 1506 862
rect 1548 848 1550 862
rect 1546 847 1552 848
rect 1546 843 1547 847
rect 1551 843 1552 847
rect 1546 842 1552 843
rect 1568 839 1570 862
rect 1620 848 1622 862
rect 1618 847 1624 848
rect 1618 843 1619 847
rect 1623 843 1624 847
rect 1618 842 1624 843
rect 1640 839 1642 862
rect 1700 848 1702 862
rect 1698 847 1704 848
rect 1698 843 1699 847
rect 1703 843 1704 847
rect 1698 842 1704 843
rect 1720 839 1722 862
rect 1728 840 1730 862
rect 1726 839 1732 840
rect 1808 839 1810 862
rect 1892 848 1894 862
rect 1890 847 1896 848
rect 1890 843 1891 847
rect 1895 843 1896 847
rect 1890 842 1896 843
rect 1912 839 1914 862
rect 1286 835 1292 836
rect 1327 838 1331 839
rect 938 834 944 835
rect 718 827 724 828
rect 718 823 719 827
rect 723 823 724 827
rect 718 822 724 823
rect 756 820 758 834
rect 754 819 760 820
rect 754 815 755 819
rect 759 815 760 819
rect 754 814 760 815
rect 776 811 778 834
rect 828 820 830 834
rect 826 819 832 820
rect 826 815 827 819
rect 831 815 832 819
rect 826 814 832 815
rect 848 811 850 834
rect 900 820 902 834
rect 898 819 904 820
rect 898 815 899 819
rect 903 815 904 819
rect 898 814 904 815
rect 920 811 922 834
rect 1288 811 1290 835
rect 1327 833 1331 834
rect 1447 838 1451 839
rect 1447 833 1451 834
rect 1503 838 1507 839
rect 1503 833 1507 834
rect 1567 838 1571 839
rect 1567 833 1571 834
rect 1591 838 1595 839
rect 1591 833 1595 834
rect 1639 838 1643 839
rect 1639 833 1643 834
rect 1647 838 1651 839
rect 1647 833 1651 834
rect 1703 838 1707 839
rect 1703 833 1707 834
rect 1719 838 1723 839
rect 1726 835 1727 839
rect 1731 835 1732 839
rect 1726 834 1732 835
rect 1767 838 1771 839
rect 1719 833 1723 834
rect 1767 833 1771 834
rect 1807 838 1811 839
rect 1807 833 1811 834
rect 1847 838 1851 839
rect 1847 833 1851 834
rect 1911 838 1915 839
rect 1911 833 1915 834
rect 1328 813 1330 833
rect 1592 814 1594 833
rect 1614 831 1620 832
rect 1614 827 1615 831
rect 1619 827 1620 831
rect 1614 826 1620 827
rect 1590 813 1596 814
rect 1326 812 1332 813
rect 703 810 707 811
rect 703 805 707 806
rect 711 810 715 811
rect 711 805 715 806
rect 767 810 771 811
rect 767 805 771 806
rect 775 810 779 811
rect 775 805 779 806
rect 831 810 835 811
rect 831 805 835 806
rect 847 810 851 811
rect 847 805 851 806
rect 895 810 899 811
rect 895 805 899 806
rect 919 810 923 811
rect 919 805 923 806
rect 967 810 971 811
rect 967 805 971 806
rect 1039 810 1043 811
rect 1039 805 1043 806
rect 1287 810 1291 811
rect 1326 808 1327 812
rect 1331 808 1332 812
rect 1590 809 1591 813
rect 1595 809 1596 813
rect 1616 812 1618 826
rect 1648 814 1650 833
rect 1670 831 1676 832
rect 1670 827 1671 831
rect 1675 827 1676 831
rect 1670 826 1676 827
rect 1646 813 1652 814
rect 1590 808 1596 809
rect 1614 811 1620 812
rect 1326 807 1332 808
rect 1614 807 1615 811
rect 1619 807 1620 811
rect 1646 809 1647 813
rect 1651 809 1652 813
rect 1672 812 1674 826
rect 1704 814 1706 833
rect 1726 831 1732 832
rect 1726 827 1727 831
rect 1731 827 1732 831
rect 1726 826 1732 827
rect 1702 813 1708 814
rect 1646 808 1652 809
rect 1670 811 1676 812
rect 1614 806 1620 807
rect 1670 807 1671 811
rect 1675 807 1676 811
rect 1702 809 1703 813
rect 1707 809 1708 813
rect 1728 812 1730 826
rect 1768 814 1770 833
rect 1848 814 1850 833
rect 1920 832 1922 862
rect 2032 839 2034 862
rect 2152 848 2154 918
rect 2198 904 2204 905
rect 2198 900 2199 904
rect 2203 900 2204 904
rect 2198 899 2204 900
rect 2278 904 2284 905
rect 2278 900 2279 904
rect 2283 900 2284 904
rect 2278 899 2284 900
rect 2358 904 2364 905
rect 2358 900 2359 904
rect 2363 900 2364 904
rect 2358 899 2364 900
rect 2438 904 2444 905
rect 2438 900 2439 904
rect 2443 900 2444 904
rect 2438 899 2444 900
rect 2200 895 2202 899
rect 2280 895 2282 899
rect 2360 895 2362 899
rect 2440 895 2442 899
rect 2199 894 2203 895
rect 2199 889 2203 890
rect 2279 894 2283 895
rect 2279 889 2283 890
rect 2359 894 2363 895
rect 2359 889 2363 890
rect 2423 894 2427 895
rect 2423 889 2427 890
rect 2439 894 2443 895
rect 2439 889 2443 890
rect 2278 888 2284 889
rect 2278 884 2279 888
rect 2283 884 2284 888
rect 2278 883 2284 884
rect 2422 888 2428 889
rect 2422 884 2423 888
rect 2427 884 2428 888
rect 2422 883 2428 884
rect 2448 868 2450 962
rect 2456 951 2458 982
rect 2455 950 2459 951
rect 2455 945 2459 946
rect 2456 926 2458 945
rect 2464 944 2466 1038
rect 2476 988 2478 1178
rect 2503 1177 2507 1178
rect 2504 1157 2506 1177
rect 2502 1156 2508 1157
rect 2502 1152 2503 1156
rect 2507 1152 2508 1156
rect 2502 1151 2508 1152
rect 2502 1139 2508 1140
rect 2502 1135 2503 1139
rect 2507 1135 2508 1139
rect 2502 1134 2508 1135
rect 2504 1131 2506 1134
rect 2503 1130 2507 1131
rect 2503 1125 2507 1126
rect 2504 1122 2506 1125
rect 2502 1121 2508 1122
rect 2502 1117 2503 1121
rect 2507 1117 2508 1121
rect 2502 1116 2508 1117
rect 2502 1104 2508 1105
rect 2502 1100 2503 1104
rect 2507 1100 2508 1104
rect 2502 1099 2508 1100
rect 2504 1071 2506 1099
rect 2503 1070 2507 1071
rect 2503 1065 2507 1066
rect 2504 1045 2506 1065
rect 2502 1044 2508 1045
rect 2502 1040 2503 1044
rect 2507 1040 2508 1044
rect 2502 1039 2508 1040
rect 2502 1027 2508 1028
rect 2502 1023 2503 1027
rect 2507 1023 2508 1027
rect 2502 1022 2508 1023
rect 2504 1015 2506 1022
rect 2503 1014 2507 1015
rect 2503 1009 2507 1010
rect 2504 1006 2506 1009
rect 2502 1005 2508 1006
rect 2502 1001 2503 1005
rect 2507 1001 2508 1005
rect 2502 1000 2508 1001
rect 2502 988 2508 989
rect 2474 987 2480 988
rect 2474 983 2475 987
rect 2479 983 2480 987
rect 2502 984 2503 988
rect 2507 984 2508 988
rect 2502 983 2508 984
rect 2474 982 2480 983
rect 2504 951 2506 983
rect 2503 950 2507 951
rect 2503 945 2507 946
rect 2462 943 2468 944
rect 2462 939 2463 943
rect 2467 939 2468 943
rect 2462 938 2468 939
rect 2454 925 2460 926
rect 2504 925 2506 945
rect 2454 921 2455 925
rect 2459 921 2460 925
rect 2502 924 2508 925
rect 2454 920 2460 921
rect 2462 923 2468 924
rect 2462 919 2463 923
rect 2467 919 2468 923
rect 2502 920 2503 924
rect 2507 920 2508 924
rect 2502 919 2508 920
rect 2462 918 2468 919
rect 2158 867 2164 868
rect 2158 863 2159 867
rect 2163 863 2164 867
rect 2158 862 2164 863
rect 2274 867 2280 868
rect 2274 863 2275 867
rect 2279 863 2280 867
rect 2274 862 2280 863
rect 2294 867 2300 868
rect 2294 863 2295 867
rect 2299 863 2300 867
rect 2294 862 2300 863
rect 2438 867 2444 868
rect 2438 863 2439 867
rect 2443 863 2444 867
rect 2438 862 2444 863
rect 2446 867 2452 868
rect 2446 863 2447 867
rect 2451 863 2452 867
rect 2446 862 2452 863
rect 2150 847 2156 848
rect 2150 843 2151 847
rect 2155 843 2156 847
rect 2150 842 2156 843
rect 2160 839 2162 862
rect 2276 848 2278 862
rect 2274 847 2280 848
rect 2274 843 2275 847
rect 2279 843 2280 847
rect 2274 842 2280 843
rect 2296 839 2298 862
rect 2406 847 2412 848
rect 2406 843 2407 847
rect 2411 843 2412 847
rect 2406 842 2412 843
rect 1927 838 1931 839
rect 1927 833 1931 834
rect 2015 838 2019 839
rect 2015 833 2019 834
rect 2031 838 2035 839
rect 2031 833 2035 834
rect 2103 838 2107 839
rect 2103 833 2107 834
rect 2159 838 2163 839
rect 2159 833 2163 834
rect 2191 838 2195 839
rect 2191 833 2195 834
rect 2287 838 2291 839
rect 2287 833 2291 834
rect 2295 838 2299 839
rect 2295 833 2299 834
rect 2383 838 2387 839
rect 2383 833 2387 834
rect 1918 831 1924 832
rect 1918 827 1919 831
rect 1923 827 1924 831
rect 1918 826 1924 827
rect 1928 814 1930 833
rect 1950 831 1956 832
rect 1950 827 1951 831
rect 1955 827 1956 831
rect 1950 826 1956 827
rect 1766 813 1772 814
rect 1702 808 1708 809
rect 1726 811 1732 812
rect 1670 806 1676 807
rect 1726 807 1727 811
rect 1731 807 1732 811
rect 1766 809 1767 813
rect 1771 809 1772 813
rect 1766 808 1772 809
rect 1846 813 1852 814
rect 1846 809 1847 813
rect 1851 809 1852 813
rect 1926 813 1932 814
rect 1846 808 1852 809
rect 1854 811 1860 812
rect 1726 806 1732 807
rect 1854 807 1855 811
rect 1859 807 1860 811
rect 1926 809 1927 813
rect 1931 809 1932 813
rect 1952 812 1954 826
rect 2016 814 2018 833
rect 2038 831 2044 832
rect 2038 827 2039 831
rect 2043 827 2044 831
rect 2038 826 2044 827
rect 2014 813 2020 814
rect 1926 808 1932 809
rect 1950 811 1956 812
rect 1854 806 1860 807
rect 1950 807 1951 811
rect 1955 807 1956 811
rect 2014 809 2015 813
rect 2019 809 2020 813
rect 2040 812 2042 826
rect 2104 814 2106 833
rect 2192 814 2194 833
rect 2214 831 2220 832
rect 2214 827 2215 831
rect 2219 827 2220 831
rect 2214 826 2220 827
rect 2102 813 2108 814
rect 2014 808 2020 809
rect 2038 811 2044 812
rect 1950 806 1956 807
rect 2038 807 2039 811
rect 2043 807 2044 811
rect 2102 809 2103 813
rect 2107 809 2108 813
rect 2190 813 2196 814
rect 2102 808 2108 809
rect 2126 811 2132 812
rect 2038 806 2044 807
rect 2126 807 2127 811
rect 2131 807 2132 811
rect 2190 809 2191 813
rect 2195 809 2196 813
rect 2216 812 2218 826
rect 2288 814 2290 833
rect 2310 831 2316 832
rect 2310 827 2311 831
rect 2315 827 2316 831
rect 2310 826 2316 827
rect 2286 813 2292 814
rect 2190 808 2196 809
rect 2214 811 2220 812
rect 2126 806 2132 807
rect 2214 807 2215 811
rect 2219 807 2220 811
rect 2286 809 2287 813
rect 2291 809 2292 813
rect 2312 812 2314 826
rect 2374 823 2380 824
rect 2374 819 2375 823
rect 2379 819 2380 823
rect 2374 818 2380 819
rect 2286 808 2292 809
rect 2310 811 2316 812
rect 2214 806 2220 807
rect 2310 807 2311 811
rect 2315 807 2316 811
rect 2310 806 2316 807
rect 1287 805 1291 806
rect 682 791 688 792
rect 682 787 683 791
rect 687 787 688 791
rect 682 786 688 787
rect 704 786 706 805
rect 768 786 770 805
rect 832 786 834 805
rect 896 786 898 805
rect 968 786 970 805
rect 1040 786 1042 805
rect 1074 803 1080 804
rect 1074 799 1075 803
rect 1079 799 1080 803
rect 1074 798 1080 799
rect 702 785 708 786
rect 630 780 636 781
rect 654 783 660 784
rect 590 778 596 779
rect 654 779 655 783
rect 659 779 660 783
rect 702 781 703 785
rect 707 781 708 785
rect 702 780 708 781
rect 766 785 772 786
rect 766 781 767 785
rect 771 781 772 785
rect 830 785 836 786
rect 766 780 772 781
rect 782 783 788 784
rect 654 778 660 779
rect 782 779 783 783
rect 787 779 788 783
rect 830 781 831 785
rect 835 781 836 785
rect 830 780 836 781
rect 894 785 900 786
rect 894 781 895 785
rect 899 781 900 785
rect 894 780 900 781
rect 966 785 972 786
rect 966 781 967 785
rect 971 781 972 785
rect 966 780 972 781
rect 1038 785 1044 786
rect 1038 781 1039 785
rect 1043 781 1044 785
rect 1038 780 1044 781
rect 782 778 788 779
rect 198 764 204 765
rect 198 760 199 764
rect 203 760 204 764
rect 198 759 204 760
rect 286 764 292 765
rect 286 760 287 764
rect 291 760 292 764
rect 286 759 292 760
rect 374 764 380 765
rect 374 760 375 764
rect 379 760 380 764
rect 374 759 380 760
rect 462 764 468 765
rect 462 760 463 764
rect 467 760 468 764
rect 462 759 468 760
rect 542 764 548 765
rect 542 760 543 764
rect 547 760 548 764
rect 542 759 548 760
rect 614 764 620 765
rect 614 760 615 764
rect 619 760 620 764
rect 614 759 620 760
rect 686 764 692 765
rect 686 760 687 764
rect 691 760 692 764
rect 686 759 692 760
rect 750 764 756 765
rect 750 760 751 764
rect 755 760 756 764
rect 750 759 756 760
rect 199 758 203 759
rect 199 753 203 754
rect 255 758 259 759
rect 255 753 259 754
rect 287 758 291 759
rect 287 753 291 754
rect 375 758 379 759
rect 375 753 379 754
rect 391 758 395 759
rect 391 753 395 754
rect 463 758 467 759
rect 463 753 467 754
rect 519 758 523 759
rect 519 753 523 754
rect 543 758 547 759
rect 543 753 547 754
rect 615 758 619 759
rect 615 753 619 754
rect 647 758 651 759
rect 647 753 651 754
rect 687 758 691 759
rect 687 753 691 754
rect 751 758 755 759
rect 751 753 755 754
rect 775 758 779 759
rect 775 753 779 754
rect 254 752 260 753
rect 254 748 255 752
rect 259 748 260 752
rect 254 747 260 748
rect 390 752 396 753
rect 390 748 391 752
rect 395 748 396 752
rect 390 747 396 748
rect 518 752 524 753
rect 518 748 519 752
rect 523 748 524 752
rect 518 747 524 748
rect 646 752 652 753
rect 646 748 647 752
rect 651 748 652 752
rect 646 747 652 748
rect 774 752 780 753
rect 774 748 775 752
rect 779 748 780 752
rect 774 747 780 748
rect 110 728 111 732
rect 115 728 116 732
rect 110 727 116 728
rect 150 731 156 732
rect 150 727 151 731
rect 155 727 156 731
rect 112 707 114 727
rect 150 726 156 727
rect 174 731 180 732
rect 174 727 175 731
rect 179 727 180 731
rect 174 726 180 727
rect 270 731 276 732
rect 270 727 271 731
rect 275 727 276 731
rect 270 726 276 727
rect 406 731 412 732
rect 406 727 407 731
rect 411 727 412 731
rect 406 726 412 727
rect 534 731 540 732
rect 534 727 535 731
rect 539 727 540 731
rect 534 726 540 727
rect 642 731 648 732
rect 642 727 643 731
rect 647 727 648 731
rect 642 726 648 727
rect 662 731 668 732
rect 662 727 663 731
rect 667 727 668 731
rect 662 726 668 727
rect 722 731 728 732
rect 722 727 723 731
rect 727 727 728 731
rect 722 726 728 727
rect 152 707 154 726
rect 272 707 274 726
rect 408 707 410 726
rect 494 711 500 712
rect 494 707 495 711
rect 499 707 500 711
rect 536 707 538 726
rect 644 712 646 726
rect 642 711 648 712
rect 642 707 643 711
rect 647 707 648 711
rect 664 707 666 726
rect 111 706 115 707
rect 111 701 115 702
rect 151 706 155 707
rect 151 701 155 702
rect 207 706 211 707
rect 207 701 211 702
rect 271 706 275 707
rect 271 701 275 702
rect 295 706 299 707
rect 295 701 299 702
rect 391 706 395 707
rect 391 701 395 702
rect 407 706 411 707
rect 494 706 500 707
rect 503 706 507 707
rect 407 701 411 702
rect 112 681 114 701
rect 152 682 154 701
rect 174 699 180 700
rect 174 695 175 699
rect 179 695 180 699
rect 174 694 180 695
rect 150 681 156 682
rect 110 680 116 681
rect 110 676 111 680
rect 115 676 116 680
rect 150 677 151 681
rect 155 677 156 681
rect 176 680 178 694
rect 208 682 210 701
rect 230 699 236 700
rect 230 695 231 699
rect 235 695 236 699
rect 230 694 236 695
rect 206 681 212 682
rect 150 676 156 677
rect 174 679 180 680
rect 110 675 116 676
rect 174 675 175 679
rect 179 675 180 679
rect 206 677 207 681
rect 211 677 212 681
rect 232 680 234 694
rect 286 691 292 692
rect 286 687 287 691
rect 291 687 292 691
rect 286 686 292 687
rect 206 676 212 677
rect 230 679 236 680
rect 174 674 180 675
rect 230 675 231 679
rect 235 675 236 679
rect 230 674 236 675
rect 110 663 116 664
rect 110 659 111 663
rect 115 659 116 663
rect 110 658 116 659
rect 134 660 140 661
rect 112 651 114 658
rect 134 656 135 660
rect 139 656 140 660
rect 134 655 140 656
rect 190 660 196 661
rect 190 656 191 660
rect 195 656 196 660
rect 190 655 196 656
rect 278 660 284 661
rect 278 656 279 660
rect 283 656 284 660
rect 278 655 284 656
rect 136 651 138 655
rect 192 651 194 655
rect 280 651 282 655
rect 111 650 115 651
rect 111 645 115 646
rect 135 650 139 651
rect 135 645 139 646
rect 151 650 155 651
rect 151 645 155 646
rect 191 650 195 651
rect 191 645 195 646
rect 263 650 267 651
rect 263 645 267 646
rect 279 650 283 651
rect 279 645 283 646
rect 112 642 114 645
rect 150 644 156 645
rect 110 641 116 642
rect 110 637 111 641
rect 115 637 116 641
rect 150 640 151 644
rect 155 640 156 644
rect 150 639 156 640
rect 262 644 268 645
rect 262 640 263 644
rect 267 640 268 644
rect 262 639 268 640
rect 110 636 116 637
rect 110 624 116 625
rect 288 624 290 686
rect 296 682 298 701
rect 392 682 394 701
rect 414 699 420 700
rect 414 695 415 699
rect 419 695 420 699
rect 414 694 420 695
rect 294 681 300 682
rect 294 677 295 681
rect 299 677 300 681
rect 294 676 300 677
rect 390 681 396 682
rect 390 677 391 681
rect 395 677 396 681
rect 416 680 418 694
rect 496 688 498 706
rect 503 701 507 702
rect 535 706 539 707
rect 535 701 539 702
rect 623 706 627 707
rect 642 706 648 707
rect 663 706 667 707
rect 623 701 627 702
rect 663 701 667 702
rect 494 687 500 688
rect 494 683 495 687
rect 499 683 500 687
rect 494 682 500 683
rect 504 682 506 701
rect 624 682 626 701
rect 724 700 726 726
rect 784 712 786 778
rect 814 764 820 765
rect 814 760 815 764
rect 819 760 820 764
rect 814 759 820 760
rect 878 764 884 765
rect 878 760 879 764
rect 883 760 884 764
rect 878 759 884 760
rect 950 764 956 765
rect 950 760 951 764
rect 955 760 956 764
rect 950 759 956 760
rect 1022 764 1028 765
rect 1022 760 1023 764
rect 1027 760 1028 764
rect 1022 759 1028 760
rect 815 758 819 759
rect 815 753 819 754
rect 879 758 883 759
rect 879 753 883 754
rect 903 758 907 759
rect 903 753 907 754
rect 951 758 955 759
rect 951 753 955 754
rect 1023 758 1027 759
rect 1023 753 1027 754
rect 1039 758 1043 759
rect 1039 753 1043 754
rect 902 752 908 753
rect 902 748 903 752
rect 907 748 908 752
rect 902 747 908 748
rect 1038 752 1044 753
rect 1038 748 1039 752
rect 1043 748 1044 752
rect 1038 747 1044 748
rect 1076 732 1078 798
rect 1288 785 1290 805
rect 1326 795 1332 796
rect 1326 791 1327 795
rect 1331 791 1332 795
rect 1326 790 1332 791
rect 1574 792 1580 793
rect 1286 784 1292 785
rect 1286 780 1287 784
rect 1291 780 1292 784
rect 1328 783 1330 790
rect 1574 788 1575 792
rect 1579 788 1580 792
rect 1574 787 1580 788
rect 1630 792 1636 793
rect 1630 788 1631 792
rect 1635 788 1636 792
rect 1630 787 1636 788
rect 1686 792 1692 793
rect 1686 788 1687 792
rect 1691 788 1692 792
rect 1686 787 1692 788
rect 1750 792 1756 793
rect 1750 788 1751 792
rect 1755 788 1756 792
rect 1750 787 1756 788
rect 1830 792 1836 793
rect 1830 788 1831 792
rect 1835 788 1836 792
rect 1830 787 1836 788
rect 1576 783 1578 787
rect 1632 783 1634 787
rect 1688 783 1690 787
rect 1752 783 1754 787
rect 1832 783 1834 787
rect 1286 779 1292 780
rect 1327 782 1331 783
rect 1327 777 1331 778
rect 1567 782 1571 783
rect 1567 777 1571 778
rect 1575 782 1579 783
rect 1575 777 1579 778
rect 1623 782 1627 783
rect 1623 777 1627 778
rect 1631 782 1635 783
rect 1631 777 1635 778
rect 1687 782 1691 783
rect 1687 777 1691 778
rect 1751 782 1755 783
rect 1751 777 1755 778
rect 1759 782 1763 783
rect 1759 777 1763 778
rect 1831 782 1835 783
rect 1831 777 1835 778
rect 1328 774 1330 777
rect 1566 776 1572 777
rect 1326 773 1332 774
rect 1326 769 1327 773
rect 1331 769 1332 773
rect 1566 772 1567 776
rect 1571 772 1572 776
rect 1566 771 1572 772
rect 1622 776 1628 777
rect 1622 772 1623 776
rect 1627 772 1628 776
rect 1622 771 1628 772
rect 1686 776 1692 777
rect 1686 772 1687 776
rect 1691 772 1692 776
rect 1686 771 1692 772
rect 1758 776 1764 777
rect 1758 772 1759 776
rect 1763 772 1764 776
rect 1758 771 1764 772
rect 1830 776 1836 777
rect 1830 772 1831 776
rect 1835 772 1836 776
rect 1830 771 1836 772
rect 1326 768 1332 769
rect 1286 767 1292 768
rect 1286 763 1287 767
rect 1291 763 1292 767
rect 1286 762 1292 763
rect 1288 759 1290 762
rect 1287 758 1291 759
rect 1287 753 1291 754
rect 1326 756 1332 757
rect 1288 750 1290 753
rect 1326 752 1327 756
rect 1331 752 1332 756
rect 1326 751 1332 752
rect 1582 755 1588 756
rect 1582 751 1583 755
rect 1587 751 1588 755
rect 1286 749 1292 750
rect 1286 745 1287 749
rect 1291 745 1292 749
rect 1286 744 1292 745
rect 1286 732 1292 733
rect 790 731 796 732
rect 790 727 791 731
rect 795 727 796 731
rect 790 726 796 727
rect 918 731 924 732
rect 918 727 919 731
rect 923 727 924 731
rect 918 726 924 727
rect 1034 731 1040 732
rect 1034 727 1035 731
rect 1039 727 1040 731
rect 1034 726 1040 727
rect 1054 731 1060 732
rect 1054 727 1055 731
rect 1059 727 1060 731
rect 1054 726 1060 727
rect 1074 731 1080 732
rect 1074 727 1075 731
rect 1079 727 1080 731
rect 1286 728 1287 732
rect 1291 728 1292 732
rect 1328 731 1330 751
rect 1582 750 1588 751
rect 1618 755 1624 756
rect 1618 751 1619 755
rect 1623 751 1624 755
rect 1618 750 1624 751
rect 1638 755 1644 756
rect 1638 751 1639 755
rect 1643 751 1644 755
rect 1638 750 1644 751
rect 1682 755 1688 756
rect 1682 751 1683 755
rect 1687 751 1688 755
rect 1682 750 1688 751
rect 1702 755 1708 756
rect 1702 751 1703 755
rect 1707 751 1708 755
rect 1702 750 1708 751
rect 1718 755 1724 756
rect 1718 751 1719 755
rect 1723 751 1724 755
rect 1718 750 1724 751
rect 1774 755 1780 756
rect 1774 751 1775 755
rect 1779 751 1780 755
rect 1774 750 1780 751
rect 1782 755 1788 756
rect 1782 751 1783 755
rect 1787 751 1788 755
rect 1782 750 1788 751
rect 1846 755 1852 756
rect 1846 751 1847 755
rect 1851 751 1852 755
rect 1846 750 1852 751
rect 1584 731 1586 750
rect 1602 743 1608 744
rect 1602 739 1603 743
rect 1607 739 1608 743
rect 1602 738 1608 739
rect 1286 727 1292 728
rect 1327 730 1331 731
rect 1074 726 1080 727
rect 782 711 788 712
rect 782 707 783 711
rect 787 707 788 711
rect 792 707 794 726
rect 894 711 900 712
rect 894 707 895 711
rect 899 707 900 711
rect 920 707 922 726
rect 1036 712 1038 726
rect 1034 711 1040 712
rect 1034 707 1035 711
rect 1039 707 1040 711
rect 1056 707 1058 726
rect 1288 707 1290 727
rect 1327 725 1331 726
rect 1367 730 1371 731
rect 1367 725 1371 726
rect 1431 730 1435 731
rect 1431 725 1435 726
rect 1527 730 1531 731
rect 1527 725 1531 726
rect 1583 730 1587 731
rect 1583 725 1587 726
rect 743 706 747 707
rect 782 706 788 707
rect 791 706 795 707
rect 743 701 747 702
rect 791 701 795 702
rect 871 706 875 707
rect 894 706 900 707
rect 919 706 923 707
rect 871 701 875 702
rect 722 699 728 700
rect 722 695 723 699
rect 727 695 728 699
rect 722 694 728 695
rect 744 682 746 701
rect 872 682 874 701
rect 502 681 508 682
rect 390 676 396 677
rect 414 679 420 680
rect 414 675 415 679
rect 419 675 420 679
rect 502 677 503 681
rect 507 677 508 681
rect 502 676 508 677
rect 622 681 628 682
rect 622 677 623 681
rect 627 677 628 681
rect 742 681 748 682
rect 622 676 628 677
rect 646 679 652 680
rect 414 674 420 675
rect 646 675 647 679
rect 651 675 652 679
rect 742 677 743 681
rect 747 677 748 681
rect 742 676 748 677
rect 870 681 876 682
rect 870 677 871 681
rect 875 677 876 681
rect 896 680 898 706
rect 919 701 923 702
rect 999 706 1003 707
rect 1034 706 1040 707
rect 1055 706 1059 707
rect 999 701 1003 702
rect 1055 701 1059 702
rect 1127 706 1131 707
rect 1127 701 1131 702
rect 1239 706 1243 707
rect 1239 701 1243 702
rect 1287 706 1291 707
rect 1328 705 1330 725
rect 1368 706 1370 725
rect 1432 706 1434 725
rect 1528 706 1530 725
rect 1604 724 1606 738
rect 1620 736 1622 750
rect 1610 735 1616 736
rect 1610 731 1611 735
rect 1615 731 1616 735
rect 1610 730 1616 731
rect 1618 735 1624 736
rect 1618 731 1619 735
rect 1623 731 1624 735
rect 1640 731 1642 750
rect 1650 743 1656 744
rect 1650 739 1651 743
rect 1655 739 1656 743
rect 1650 738 1656 739
rect 1618 730 1624 731
rect 1631 730 1635 731
rect 1602 723 1608 724
rect 1602 719 1603 723
rect 1607 719 1608 723
rect 1612 723 1614 730
rect 1622 727 1628 728
rect 1622 723 1623 727
rect 1627 723 1628 727
rect 1631 725 1635 726
rect 1639 730 1643 731
rect 1639 725 1643 726
rect 1612 722 1628 723
rect 1612 721 1626 722
rect 1602 718 1608 719
rect 1632 706 1634 725
rect 1366 705 1372 706
rect 1287 701 1291 702
rect 1326 704 1332 705
rect 974 699 980 700
rect 974 695 975 699
rect 979 695 980 699
rect 974 694 980 695
rect 870 676 876 677
rect 894 679 900 680
rect 646 674 652 675
rect 894 675 895 679
rect 899 675 900 679
rect 894 674 900 675
rect 374 660 380 661
rect 374 656 375 660
rect 379 656 380 660
rect 374 655 380 656
rect 486 660 492 661
rect 486 656 487 660
rect 491 656 492 660
rect 486 655 492 656
rect 606 660 612 661
rect 606 656 607 660
rect 611 656 612 660
rect 606 655 612 656
rect 376 651 378 655
rect 488 651 490 655
rect 608 651 610 655
rect 367 650 371 651
rect 367 645 371 646
rect 375 650 379 651
rect 375 645 379 646
rect 463 650 467 651
rect 463 645 467 646
rect 487 650 491 651
rect 487 645 491 646
rect 559 650 563 651
rect 559 645 563 646
rect 607 650 611 651
rect 607 645 611 646
rect 366 644 372 645
rect 366 640 367 644
rect 371 640 372 644
rect 366 639 372 640
rect 462 644 468 645
rect 462 640 463 644
rect 467 640 468 644
rect 462 639 468 640
rect 558 644 564 645
rect 558 640 559 644
rect 563 640 564 644
rect 558 639 564 640
rect 110 620 111 624
rect 115 620 116 624
rect 110 619 116 620
rect 166 623 172 624
rect 166 619 167 623
rect 171 619 172 623
rect 112 599 114 619
rect 166 618 172 619
rect 258 623 264 624
rect 258 619 259 623
rect 263 619 264 623
rect 258 618 264 619
rect 278 623 284 624
rect 278 619 279 623
rect 283 619 284 623
rect 278 618 284 619
rect 286 623 292 624
rect 286 619 287 623
rect 291 619 292 623
rect 286 618 292 619
rect 382 623 388 624
rect 382 619 383 623
rect 387 619 388 623
rect 382 618 388 619
rect 406 623 412 624
rect 406 619 407 623
rect 411 619 412 623
rect 406 618 412 619
rect 478 623 484 624
rect 478 619 479 623
rect 483 619 484 623
rect 478 618 484 619
rect 486 623 492 624
rect 486 619 487 623
rect 491 619 492 623
rect 486 618 492 619
rect 574 623 580 624
rect 574 619 575 623
rect 579 619 580 623
rect 574 618 580 619
rect 158 603 164 604
rect 158 599 159 603
rect 163 599 164 603
rect 168 599 170 618
rect 260 604 262 618
rect 258 603 264 604
rect 258 599 259 603
rect 263 599 264 603
rect 280 599 282 618
rect 384 599 386 618
rect 111 598 115 599
rect 111 593 115 594
rect 151 598 155 599
rect 158 598 164 599
rect 167 598 171 599
rect 151 593 155 594
rect 112 573 114 593
rect 152 574 154 593
rect 150 573 156 574
rect 110 572 116 573
rect 110 568 111 572
rect 115 568 116 572
rect 150 569 151 573
rect 155 569 156 573
rect 160 572 162 598
rect 167 593 171 594
rect 239 598 243 599
rect 258 598 264 599
rect 279 598 283 599
rect 239 593 243 594
rect 279 593 283 594
rect 335 598 339 599
rect 335 593 339 594
rect 383 598 387 599
rect 383 593 387 594
rect 240 574 242 593
rect 286 591 292 592
rect 286 587 287 591
rect 291 587 292 591
rect 286 586 292 587
rect 238 573 244 574
rect 150 568 156 569
rect 158 571 164 572
rect 110 567 116 568
rect 158 567 159 571
rect 163 567 164 571
rect 238 569 239 573
rect 243 569 244 573
rect 238 568 244 569
rect 158 566 164 567
rect 110 555 116 556
rect 110 551 111 555
rect 115 551 116 555
rect 110 550 116 551
rect 134 552 140 553
rect 112 539 114 550
rect 134 548 135 552
rect 139 548 140 552
rect 134 547 140 548
rect 222 552 228 553
rect 222 548 223 552
rect 227 548 228 552
rect 222 547 228 548
rect 136 539 138 547
rect 224 539 226 547
rect 111 538 115 539
rect 111 533 115 534
rect 135 538 139 539
rect 135 533 139 534
rect 143 538 147 539
rect 143 533 147 534
rect 223 538 227 539
rect 223 533 227 534
rect 239 538 243 539
rect 239 533 243 534
rect 112 530 114 533
rect 142 532 148 533
rect 110 529 116 530
rect 110 525 111 529
rect 115 525 116 529
rect 142 528 143 532
rect 147 528 148 532
rect 142 527 148 528
rect 238 532 244 533
rect 238 528 239 532
rect 243 528 244 532
rect 238 527 244 528
rect 110 524 116 525
rect 110 512 116 513
rect 288 512 290 586
rect 336 574 338 593
rect 408 592 410 618
rect 480 599 482 618
rect 488 600 490 618
rect 486 599 492 600
rect 576 599 578 618
rect 648 604 650 674
rect 726 660 732 661
rect 726 656 727 660
rect 731 656 732 660
rect 726 655 732 656
rect 854 660 860 661
rect 854 656 855 660
rect 859 656 860 660
rect 854 655 860 656
rect 728 651 730 655
rect 856 651 858 655
rect 655 650 659 651
rect 655 645 659 646
rect 727 650 731 651
rect 727 645 731 646
rect 751 650 755 651
rect 751 645 755 646
rect 847 650 851 651
rect 847 645 851 646
rect 855 650 859 651
rect 855 645 859 646
rect 943 650 947 651
rect 943 645 947 646
rect 654 644 660 645
rect 654 640 655 644
rect 659 640 660 644
rect 654 639 660 640
rect 750 644 756 645
rect 750 640 751 644
rect 755 640 756 644
rect 750 639 756 640
rect 846 644 852 645
rect 846 640 847 644
rect 851 640 852 644
rect 846 639 852 640
rect 942 644 948 645
rect 942 640 943 644
rect 947 640 948 644
rect 942 639 948 640
rect 976 624 978 694
rect 1000 682 1002 701
rect 1128 682 1130 701
rect 1150 699 1156 700
rect 1150 695 1151 699
rect 1155 695 1156 699
rect 1150 694 1156 695
rect 998 681 1004 682
rect 998 677 999 681
rect 1003 677 1004 681
rect 998 676 1004 677
rect 1126 681 1132 682
rect 1126 677 1127 681
rect 1131 677 1132 681
rect 1152 680 1154 694
rect 1240 682 1242 701
rect 1238 681 1244 682
rect 1288 681 1290 701
rect 1326 700 1327 704
rect 1331 700 1332 704
rect 1366 701 1367 705
rect 1371 701 1372 705
rect 1366 700 1372 701
rect 1430 705 1436 706
rect 1430 701 1431 705
rect 1435 701 1436 705
rect 1430 700 1436 701
rect 1526 705 1532 706
rect 1526 701 1527 705
rect 1531 701 1532 705
rect 1526 700 1532 701
rect 1630 705 1636 706
rect 1630 701 1631 705
rect 1635 701 1636 705
rect 1652 704 1654 738
rect 1684 736 1686 750
rect 1682 735 1688 736
rect 1682 731 1683 735
rect 1687 731 1688 735
rect 1704 731 1706 750
rect 1682 730 1688 731
rect 1703 730 1707 731
rect 1703 725 1707 726
rect 1720 724 1722 750
rect 1776 731 1778 750
rect 1784 732 1786 750
rect 1782 731 1788 732
rect 1848 731 1850 750
rect 1856 736 1858 806
rect 1910 792 1916 793
rect 1910 788 1911 792
rect 1915 788 1916 792
rect 1910 787 1916 788
rect 1998 792 2004 793
rect 1998 788 1999 792
rect 2003 788 2004 792
rect 1998 787 2004 788
rect 2086 792 2092 793
rect 2086 788 2087 792
rect 2091 788 2092 792
rect 2086 787 2092 788
rect 1912 783 1914 787
rect 2000 783 2002 787
rect 2088 783 2090 787
rect 1911 782 1915 783
rect 1911 777 1915 778
rect 1919 782 1923 783
rect 1919 777 1923 778
rect 1999 782 2003 783
rect 1999 777 2003 778
rect 2015 782 2019 783
rect 2015 777 2019 778
rect 2087 782 2091 783
rect 2087 777 2091 778
rect 2119 782 2123 783
rect 2119 777 2123 778
rect 1918 776 1924 777
rect 1918 772 1919 776
rect 1923 772 1924 776
rect 1918 771 1924 772
rect 2014 776 2020 777
rect 2014 772 2015 776
rect 2019 772 2020 776
rect 2014 771 2020 772
rect 2118 776 2124 777
rect 2118 772 2119 776
rect 2123 772 2124 776
rect 2118 771 2124 772
rect 1934 755 1940 756
rect 1934 751 1935 755
rect 1939 751 1940 755
rect 1934 750 1940 751
rect 2010 755 2016 756
rect 2010 751 2011 755
rect 2015 751 2016 755
rect 2010 750 2016 751
rect 2030 755 2036 756
rect 2030 751 2031 755
rect 2035 751 2036 755
rect 2030 750 2036 751
rect 2114 755 2120 756
rect 2114 751 2115 755
rect 2119 751 2120 755
rect 2114 750 2120 751
rect 1854 735 1860 736
rect 1854 731 1855 735
rect 1859 731 1860 735
rect 1936 731 1938 750
rect 2012 736 2014 750
rect 2010 735 2016 736
rect 2010 731 2011 735
rect 2015 731 2016 735
rect 2032 731 2034 750
rect 2116 736 2118 750
rect 2128 744 2130 806
rect 2174 792 2180 793
rect 2174 788 2175 792
rect 2179 788 2180 792
rect 2174 787 2180 788
rect 2270 792 2276 793
rect 2270 788 2271 792
rect 2275 788 2276 792
rect 2270 787 2276 788
rect 2366 792 2372 793
rect 2366 788 2367 792
rect 2371 788 2372 792
rect 2366 787 2372 788
rect 2176 783 2178 787
rect 2272 783 2274 787
rect 2368 783 2370 787
rect 2175 782 2179 783
rect 2175 777 2179 778
rect 2231 782 2235 783
rect 2231 777 2235 778
rect 2271 782 2275 783
rect 2271 777 2275 778
rect 2343 782 2347 783
rect 2343 777 2347 778
rect 2367 782 2371 783
rect 2367 777 2371 778
rect 2230 776 2236 777
rect 2230 772 2231 776
rect 2235 772 2236 776
rect 2230 771 2236 772
rect 2342 776 2348 777
rect 2342 772 2343 776
rect 2347 772 2348 776
rect 2342 771 2348 772
rect 2376 756 2378 818
rect 2384 814 2386 833
rect 2382 813 2388 814
rect 2382 809 2383 813
rect 2387 809 2388 813
rect 2408 812 2410 842
rect 2440 839 2442 862
rect 2439 838 2443 839
rect 2439 833 2443 834
rect 2455 838 2459 839
rect 2455 833 2459 834
rect 2456 814 2458 833
rect 2464 832 2466 918
rect 2502 907 2508 908
rect 2502 903 2503 907
rect 2507 903 2508 907
rect 2502 902 2508 903
rect 2504 895 2506 902
rect 2503 894 2507 895
rect 2503 889 2507 890
rect 2504 886 2506 889
rect 2502 885 2508 886
rect 2502 881 2503 885
rect 2507 881 2508 885
rect 2502 880 2508 881
rect 2502 868 2508 869
rect 2502 864 2503 868
rect 2507 864 2508 868
rect 2502 863 2508 864
rect 2504 839 2506 863
rect 2503 838 2507 839
rect 2503 833 2507 834
rect 2462 831 2468 832
rect 2462 827 2463 831
rect 2467 827 2468 831
rect 2462 826 2468 827
rect 2454 813 2460 814
rect 2504 813 2506 833
rect 2382 808 2388 809
rect 2406 811 2412 812
rect 2406 807 2407 811
rect 2411 807 2412 811
rect 2454 809 2455 813
rect 2459 809 2460 813
rect 2502 812 2508 813
rect 2454 808 2460 809
rect 2470 811 2476 812
rect 2406 806 2412 807
rect 2470 807 2471 811
rect 2475 807 2476 811
rect 2502 808 2503 812
rect 2507 808 2508 812
rect 2502 807 2508 808
rect 2470 806 2476 807
rect 2438 792 2444 793
rect 2438 788 2439 792
rect 2443 788 2444 792
rect 2438 787 2444 788
rect 2440 783 2442 787
rect 2439 782 2443 783
rect 2439 777 2443 778
rect 2438 776 2444 777
rect 2438 772 2439 776
rect 2443 772 2444 776
rect 2438 771 2444 772
rect 2134 755 2140 756
rect 2134 751 2135 755
rect 2139 751 2140 755
rect 2134 750 2140 751
rect 2226 755 2232 756
rect 2226 751 2227 755
rect 2231 751 2232 755
rect 2226 750 2232 751
rect 2246 755 2252 756
rect 2246 751 2247 755
rect 2251 751 2252 755
rect 2246 750 2252 751
rect 2358 755 2364 756
rect 2358 751 2359 755
rect 2363 751 2364 755
rect 2358 750 2364 751
rect 2374 755 2380 756
rect 2374 751 2375 755
rect 2379 751 2380 755
rect 2374 750 2380 751
rect 2454 755 2460 756
rect 2454 751 2455 755
rect 2459 751 2460 755
rect 2454 750 2460 751
rect 2462 755 2468 756
rect 2462 751 2463 755
rect 2467 751 2468 755
rect 2462 750 2468 751
rect 2126 743 2132 744
rect 2126 739 2127 743
rect 2131 739 2132 743
rect 2126 738 2132 739
rect 2114 735 2120 736
rect 2114 731 2115 735
rect 2119 731 2120 735
rect 2136 731 2138 750
rect 2142 747 2148 748
rect 2142 743 2143 747
rect 2147 743 2148 747
rect 2142 742 2148 743
rect 1735 730 1739 731
rect 1735 725 1739 726
rect 1775 730 1779 731
rect 1782 727 1783 731
rect 1787 727 1788 731
rect 1782 726 1788 727
rect 1839 730 1843 731
rect 1775 725 1779 726
rect 1839 725 1843 726
rect 1847 730 1851 731
rect 1854 730 1860 731
rect 1935 730 1939 731
rect 1847 725 1851 726
rect 1935 725 1939 726
rect 1943 730 1947 731
rect 2010 730 2016 731
rect 2031 730 2035 731
rect 1943 725 1947 726
rect 2031 725 2035 726
rect 2047 730 2051 731
rect 2114 730 2120 731
rect 2135 730 2139 731
rect 2047 725 2051 726
rect 2135 725 2139 726
rect 1718 723 1724 724
rect 1718 719 1719 723
rect 1723 719 1724 723
rect 1718 718 1724 719
rect 1736 706 1738 725
rect 1840 706 1842 725
rect 1854 723 1860 724
rect 1854 719 1855 723
rect 1859 719 1860 723
rect 1854 718 1860 719
rect 1862 723 1868 724
rect 1862 719 1863 723
rect 1867 719 1868 723
rect 1862 718 1868 719
rect 1734 705 1740 706
rect 1630 700 1636 701
rect 1650 703 1656 704
rect 1326 699 1332 700
rect 1650 699 1651 703
rect 1655 699 1656 703
rect 1734 701 1735 705
rect 1739 701 1740 705
rect 1734 700 1740 701
rect 1838 705 1844 706
rect 1838 701 1839 705
rect 1843 701 1844 705
rect 1838 700 1844 701
rect 1650 698 1656 699
rect 1326 687 1332 688
rect 1326 683 1327 687
rect 1331 683 1332 687
rect 1326 682 1332 683
rect 1350 684 1356 685
rect 1126 676 1132 677
rect 1150 679 1156 680
rect 1150 675 1151 679
rect 1155 675 1156 679
rect 1238 677 1239 681
rect 1243 677 1244 681
rect 1238 676 1244 677
rect 1286 680 1292 681
rect 1286 676 1287 680
rect 1291 676 1292 680
rect 1286 675 1292 676
rect 1150 674 1156 675
rect 1328 667 1330 682
rect 1350 680 1351 684
rect 1355 680 1356 684
rect 1350 679 1356 680
rect 1414 684 1420 685
rect 1414 680 1415 684
rect 1419 680 1420 684
rect 1414 679 1420 680
rect 1510 684 1516 685
rect 1510 680 1511 684
rect 1515 680 1516 684
rect 1510 679 1516 680
rect 1614 684 1620 685
rect 1614 680 1615 684
rect 1619 680 1620 684
rect 1614 679 1620 680
rect 1718 684 1724 685
rect 1718 680 1719 684
rect 1723 680 1724 684
rect 1718 679 1724 680
rect 1822 684 1828 685
rect 1822 680 1823 684
rect 1827 680 1828 684
rect 1822 679 1828 680
rect 1342 671 1348 672
rect 1342 667 1343 671
rect 1347 667 1348 671
rect 1352 667 1354 679
rect 1416 667 1418 679
rect 1512 667 1514 679
rect 1616 667 1618 679
rect 1720 667 1722 679
rect 1824 667 1826 679
rect 1327 666 1331 667
rect 1342 666 1348 667
rect 1351 666 1355 667
rect 1286 663 1292 664
rect 982 660 988 661
rect 982 656 983 660
rect 987 656 988 660
rect 982 655 988 656
rect 1110 660 1116 661
rect 1110 656 1111 660
rect 1115 656 1116 660
rect 1110 655 1116 656
rect 1222 660 1228 661
rect 1222 656 1223 660
rect 1227 656 1228 660
rect 1286 659 1287 663
rect 1291 659 1292 663
rect 1327 661 1331 662
rect 1286 658 1292 659
rect 1328 658 1330 661
rect 1222 655 1228 656
rect 984 651 986 655
rect 1112 651 1114 655
rect 1224 651 1226 655
rect 1288 651 1290 658
rect 1326 657 1332 658
rect 1326 653 1327 657
rect 1331 653 1332 657
rect 1326 652 1332 653
rect 983 650 987 651
rect 983 645 987 646
rect 1039 650 1043 651
rect 1039 645 1043 646
rect 1111 650 1115 651
rect 1111 645 1115 646
rect 1143 650 1147 651
rect 1143 645 1147 646
rect 1223 650 1227 651
rect 1223 645 1227 646
rect 1287 650 1291 651
rect 1287 645 1291 646
rect 1038 644 1044 645
rect 1038 640 1039 644
rect 1043 640 1044 644
rect 1038 639 1044 640
rect 1142 644 1148 645
rect 1142 640 1143 644
rect 1147 640 1148 644
rect 1142 639 1148 640
rect 1222 644 1228 645
rect 1222 640 1223 644
rect 1227 640 1228 644
rect 1288 642 1290 645
rect 1222 639 1228 640
rect 1286 641 1292 642
rect 1286 637 1287 641
rect 1291 637 1292 641
rect 1286 636 1292 637
rect 1326 640 1332 641
rect 1326 636 1327 640
rect 1331 636 1332 640
rect 1326 635 1332 636
rect 1262 631 1268 632
rect 1262 627 1263 631
rect 1267 627 1268 631
rect 1262 626 1268 627
rect 670 623 676 624
rect 670 619 671 623
rect 675 619 676 623
rect 670 618 676 619
rect 766 623 772 624
rect 766 619 767 623
rect 771 619 772 623
rect 766 618 772 619
rect 842 623 848 624
rect 842 619 843 623
rect 847 619 848 623
rect 842 618 848 619
rect 862 623 868 624
rect 862 619 863 623
rect 867 619 868 623
rect 862 618 868 619
rect 938 623 944 624
rect 938 619 939 623
rect 943 619 944 623
rect 938 618 944 619
rect 958 623 964 624
rect 958 619 959 623
rect 963 619 964 623
rect 958 618 964 619
rect 974 623 980 624
rect 974 619 975 623
rect 979 619 980 623
rect 974 618 980 619
rect 1054 623 1060 624
rect 1054 619 1055 623
rect 1059 619 1060 623
rect 1054 618 1060 619
rect 1138 623 1144 624
rect 1138 619 1139 623
rect 1143 619 1144 623
rect 1138 618 1144 619
rect 1158 623 1164 624
rect 1158 619 1159 623
rect 1163 619 1164 623
rect 1158 618 1164 619
rect 1166 623 1172 624
rect 1166 619 1167 623
rect 1171 619 1172 623
rect 1166 618 1172 619
rect 1238 623 1244 624
rect 1238 619 1239 623
rect 1243 619 1244 623
rect 1238 618 1244 619
rect 646 603 652 604
rect 646 599 647 603
rect 651 599 652 603
rect 672 599 674 618
rect 768 599 770 618
rect 844 604 846 618
rect 834 603 840 604
rect 834 599 835 603
rect 839 599 840 603
rect 431 598 435 599
rect 431 593 435 594
rect 479 598 483 599
rect 486 595 487 599
rect 491 595 492 599
rect 486 594 492 595
rect 535 598 539 599
rect 479 593 483 594
rect 535 593 539 594
rect 575 598 579 599
rect 575 593 579 594
rect 631 598 635 599
rect 646 598 652 599
rect 671 598 675 599
rect 631 593 635 594
rect 671 593 675 594
rect 727 598 731 599
rect 727 593 731 594
rect 767 598 771 599
rect 767 593 771 594
rect 823 598 827 599
rect 834 598 840 599
rect 842 603 848 604
rect 842 599 843 603
rect 847 599 848 603
rect 864 599 866 618
rect 940 604 942 618
rect 938 603 944 604
rect 938 599 939 603
rect 943 599 944 603
rect 960 599 962 618
rect 1018 599 1024 600
rect 1056 599 1058 618
rect 1140 604 1142 618
rect 1138 603 1144 604
rect 1138 599 1139 603
rect 1143 599 1144 603
rect 1160 599 1162 618
rect 842 598 848 599
rect 863 598 867 599
rect 823 593 827 594
rect 406 591 412 592
rect 406 587 407 591
rect 411 587 412 591
rect 406 586 412 587
rect 432 574 434 593
rect 454 591 460 592
rect 454 587 455 591
rect 459 587 460 591
rect 454 586 460 587
rect 334 573 340 574
rect 334 569 335 573
rect 339 569 340 573
rect 334 568 340 569
rect 430 573 436 574
rect 430 569 431 573
rect 435 569 436 573
rect 456 572 458 586
rect 536 574 538 593
rect 558 591 564 592
rect 558 587 559 591
rect 563 587 564 591
rect 558 586 564 587
rect 534 573 540 574
rect 430 568 436 569
rect 454 571 460 572
rect 454 567 455 571
rect 459 567 460 571
rect 534 569 535 573
rect 539 569 540 573
rect 560 572 562 586
rect 632 574 634 593
rect 728 574 730 593
rect 742 591 748 592
rect 742 587 743 591
rect 747 587 748 591
rect 742 586 748 587
rect 750 591 756 592
rect 750 587 751 591
rect 755 587 756 591
rect 750 586 756 587
rect 630 573 636 574
rect 534 568 540 569
rect 558 571 564 572
rect 454 566 460 567
rect 558 567 559 571
rect 563 567 564 571
rect 630 569 631 573
rect 635 569 636 573
rect 726 573 732 574
rect 630 568 636 569
rect 646 571 652 572
rect 558 566 564 567
rect 646 567 647 571
rect 651 567 652 571
rect 726 569 727 573
rect 731 569 732 573
rect 726 568 732 569
rect 646 566 652 567
rect 318 552 324 553
rect 318 548 319 552
rect 323 548 324 552
rect 318 547 324 548
rect 414 552 420 553
rect 414 548 415 552
rect 419 548 420 552
rect 414 547 420 548
rect 518 552 524 553
rect 518 548 519 552
rect 523 548 524 552
rect 518 547 524 548
rect 614 552 620 553
rect 614 548 615 552
rect 619 548 620 552
rect 614 547 620 548
rect 320 539 322 547
rect 416 539 418 547
rect 520 539 522 547
rect 616 539 618 547
rect 319 538 323 539
rect 319 533 323 534
rect 335 538 339 539
rect 335 533 339 534
rect 415 538 419 539
rect 415 533 419 534
rect 431 538 435 539
rect 431 533 435 534
rect 519 538 523 539
rect 519 533 523 534
rect 527 538 531 539
rect 527 533 531 534
rect 615 538 619 539
rect 615 533 619 534
rect 623 538 627 539
rect 623 533 627 534
rect 334 532 340 533
rect 334 528 335 532
rect 339 528 340 532
rect 334 527 340 528
rect 430 532 436 533
rect 430 528 431 532
rect 435 528 436 532
rect 430 527 436 528
rect 526 532 532 533
rect 526 528 527 532
rect 531 528 532 532
rect 526 527 532 528
rect 622 532 628 533
rect 622 528 623 532
rect 627 528 628 532
rect 622 527 628 528
rect 110 508 111 512
rect 115 508 116 512
rect 110 507 116 508
rect 158 511 164 512
rect 158 507 159 511
rect 163 507 164 511
rect 112 483 114 507
rect 158 506 164 507
rect 234 511 240 512
rect 234 507 235 511
rect 239 507 240 511
rect 234 506 240 507
rect 254 511 260 512
rect 254 507 255 511
rect 259 507 260 511
rect 254 506 260 507
rect 286 511 292 512
rect 286 507 287 511
rect 291 507 292 511
rect 286 506 292 507
rect 350 511 356 512
rect 350 507 351 511
rect 355 507 356 511
rect 350 506 356 507
rect 426 511 432 512
rect 426 507 427 511
rect 431 507 432 511
rect 426 506 432 507
rect 446 511 452 512
rect 446 507 447 511
rect 451 507 452 511
rect 446 506 452 507
rect 454 511 460 512
rect 454 507 455 511
rect 459 507 460 511
rect 454 506 460 507
rect 542 511 548 512
rect 542 507 543 511
rect 547 507 548 511
rect 542 506 548 507
rect 638 511 644 512
rect 638 507 639 511
rect 643 507 644 511
rect 638 506 644 507
rect 160 483 162 506
rect 236 492 238 506
rect 170 491 176 492
rect 170 487 171 491
rect 175 487 176 491
rect 170 486 176 487
rect 234 491 240 492
rect 234 487 235 491
rect 239 487 240 491
rect 234 486 240 487
rect 111 482 115 483
rect 111 477 115 478
rect 151 482 155 483
rect 151 477 155 478
rect 159 482 163 483
rect 159 477 163 478
rect 112 457 114 477
rect 152 458 154 477
rect 150 457 156 458
rect 110 456 116 457
rect 110 452 111 456
rect 115 452 116 456
rect 150 453 151 457
rect 155 453 156 457
rect 172 456 174 486
rect 256 483 258 506
rect 352 483 354 506
rect 428 492 430 506
rect 426 491 432 492
rect 426 487 427 491
rect 431 487 432 491
rect 426 486 432 487
rect 448 483 450 506
rect 207 482 211 483
rect 207 477 211 478
rect 255 482 259 483
rect 255 477 259 478
rect 287 482 291 483
rect 287 477 291 478
rect 351 482 355 483
rect 351 477 355 478
rect 375 482 379 483
rect 375 477 379 478
rect 447 482 451 483
rect 447 477 451 478
rect 208 458 210 477
rect 288 458 290 477
rect 310 475 316 476
rect 302 471 308 472
rect 302 467 303 471
rect 307 467 308 471
rect 310 471 311 475
rect 315 471 316 475
rect 310 470 316 471
rect 302 466 308 467
rect 206 457 212 458
rect 150 452 156 453
rect 170 455 176 456
rect 110 451 116 452
rect 170 451 171 455
rect 175 451 176 455
rect 206 453 207 457
rect 211 453 212 457
rect 206 452 212 453
rect 286 457 292 458
rect 286 453 287 457
rect 291 453 292 457
rect 286 452 292 453
rect 170 450 176 451
rect 110 439 116 440
rect 110 435 111 439
rect 115 435 116 439
rect 110 434 116 435
rect 134 436 140 437
rect 112 431 114 434
rect 134 432 135 436
rect 139 432 140 436
rect 134 431 140 432
rect 190 436 196 437
rect 190 432 191 436
rect 195 432 196 436
rect 190 431 196 432
rect 270 436 276 437
rect 270 432 271 436
rect 275 432 276 436
rect 270 431 276 432
rect 111 430 115 431
rect 111 425 115 426
rect 135 430 139 431
rect 135 425 139 426
rect 191 430 195 431
rect 191 425 195 426
rect 271 430 275 431
rect 271 425 275 426
rect 279 430 283 431
rect 279 425 283 426
rect 112 422 114 425
rect 134 424 140 425
rect 110 421 116 422
rect 110 417 111 421
rect 115 417 116 421
rect 134 420 135 424
rect 139 420 140 424
rect 134 419 140 420
rect 190 424 196 425
rect 190 420 191 424
rect 195 420 196 424
rect 190 419 196 420
rect 278 424 284 425
rect 278 420 279 424
rect 283 420 284 424
rect 278 419 284 420
rect 110 416 116 417
rect 110 404 116 405
rect 304 404 306 466
rect 312 456 314 470
rect 376 458 378 477
rect 456 476 458 506
rect 544 483 546 506
rect 578 483 584 484
rect 640 483 642 506
rect 648 500 650 566
rect 710 552 716 553
rect 710 548 711 552
rect 715 548 716 552
rect 710 547 716 548
rect 712 539 714 547
rect 711 538 715 539
rect 711 533 715 534
rect 710 532 716 533
rect 710 528 711 532
rect 715 528 716 532
rect 710 527 716 528
rect 744 512 746 586
rect 752 572 754 586
rect 824 574 826 593
rect 822 573 828 574
rect 750 571 756 572
rect 750 567 751 571
rect 755 567 756 571
rect 822 569 823 573
rect 827 569 828 573
rect 836 572 838 598
rect 863 593 867 594
rect 911 598 915 599
rect 938 598 944 599
rect 959 598 963 599
rect 911 593 915 594
rect 959 593 963 594
rect 999 598 1003 599
rect 1018 595 1019 599
rect 1023 595 1024 599
rect 1018 594 1024 595
rect 1055 598 1059 599
rect 999 593 1003 594
rect 912 574 914 593
rect 1000 574 1002 593
rect 910 573 916 574
rect 822 568 828 569
rect 834 571 840 572
rect 750 566 756 567
rect 834 567 835 571
rect 839 567 840 571
rect 910 569 911 573
rect 915 569 916 573
rect 998 573 1004 574
rect 910 568 916 569
rect 942 571 948 572
rect 834 566 840 567
rect 942 567 943 571
rect 947 567 948 571
rect 998 569 999 573
rect 1003 569 1004 573
rect 1020 572 1022 594
rect 1055 593 1059 594
rect 1087 598 1091 599
rect 1138 598 1144 599
rect 1159 598 1163 599
rect 1087 593 1091 594
rect 1159 593 1163 594
rect 1088 574 1090 593
rect 1168 592 1170 618
rect 1240 599 1242 618
rect 1264 604 1266 626
rect 1286 624 1292 625
rect 1286 620 1287 624
rect 1291 620 1292 624
rect 1286 619 1292 620
rect 1262 603 1268 604
rect 1262 599 1263 603
rect 1267 599 1268 603
rect 1288 599 1290 619
rect 1328 615 1330 635
rect 1344 620 1346 666
rect 1351 661 1355 662
rect 1415 666 1419 667
rect 1415 661 1419 662
rect 1511 666 1515 667
rect 1511 661 1515 662
rect 1607 666 1611 667
rect 1607 661 1611 662
rect 1615 666 1619 667
rect 1615 661 1619 662
rect 1711 666 1715 667
rect 1711 661 1715 662
rect 1719 666 1723 667
rect 1719 661 1723 662
rect 1823 666 1827 667
rect 1823 661 1827 662
rect 1350 660 1356 661
rect 1350 656 1351 660
rect 1355 656 1356 660
rect 1350 655 1356 656
rect 1414 660 1420 661
rect 1414 656 1415 660
rect 1419 656 1420 660
rect 1414 655 1420 656
rect 1510 660 1516 661
rect 1510 656 1511 660
rect 1515 656 1516 660
rect 1510 655 1516 656
rect 1606 660 1612 661
rect 1606 656 1607 660
rect 1611 656 1612 660
rect 1606 655 1612 656
rect 1710 660 1716 661
rect 1710 656 1711 660
rect 1715 656 1716 660
rect 1710 655 1716 656
rect 1822 660 1828 661
rect 1822 656 1823 660
rect 1827 656 1828 660
rect 1822 655 1828 656
rect 1856 640 1858 718
rect 1864 704 1866 718
rect 1944 706 1946 725
rect 1966 723 1972 724
rect 1966 719 1967 723
rect 1971 719 1972 723
rect 1966 718 1972 719
rect 1942 705 1948 706
rect 1862 703 1868 704
rect 1862 699 1863 703
rect 1867 699 1868 703
rect 1942 701 1943 705
rect 1947 701 1948 705
rect 1968 704 1970 718
rect 2048 706 2050 725
rect 2144 724 2146 742
rect 2228 736 2230 750
rect 2226 735 2232 736
rect 2226 731 2227 735
rect 2231 731 2232 735
rect 2248 731 2250 750
rect 2360 731 2362 750
rect 2386 735 2392 736
rect 2386 731 2387 735
rect 2391 731 2392 735
rect 2456 731 2458 750
rect 2151 730 2155 731
rect 2226 730 2232 731
rect 2247 730 2251 731
rect 2151 725 2155 726
rect 2247 725 2251 726
rect 2255 730 2259 731
rect 2255 725 2259 726
rect 2359 730 2363 731
rect 2359 725 2363 726
rect 2367 730 2371 731
rect 2386 730 2392 731
rect 2455 730 2459 731
rect 2367 725 2371 726
rect 2142 723 2148 724
rect 2142 719 2143 723
rect 2147 719 2148 723
rect 2142 718 2148 719
rect 2152 706 2154 725
rect 2174 723 2180 724
rect 2174 719 2175 723
rect 2179 719 2180 723
rect 2174 718 2180 719
rect 2046 705 2052 706
rect 1942 700 1948 701
rect 1966 703 1972 704
rect 1862 698 1868 699
rect 1966 699 1967 703
rect 1971 699 1972 703
rect 2046 701 2047 705
rect 2051 701 2052 705
rect 2150 705 2156 706
rect 2046 700 2052 701
rect 2062 703 2068 704
rect 1966 698 1972 699
rect 2062 699 2063 703
rect 2067 699 2068 703
rect 2150 701 2151 705
rect 2155 701 2156 705
rect 2176 704 2178 718
rect 2256 706 2258 725
rect 2278 723 2284 724
rect 2278 719 2279 723
rect 2283 719 2284 723
rect 2278 718 2284 719
rect 2254 705 2260 706
rect 2150 700 2156 701
rect 2174 703 2180 704
rect 2062 698 2068 699
rect 2174 699 2175 703
rect 2179 699 2180 703
rect 2254 701 2255 705
rect 2259 701 2260 705
rect 2280 704 2282 718
rect 2368 706 2370 725
rect 2366 705 2372 706
rect 2254 700 2260 701
rect 2278 703 2284 704
rect 2174 698 2180 699
rect 2278 699 2279 703
rect 2283 699 2284 703
rect 2366 701 2367 705
rect 2371 701 2372 705
rect 2388 704 2390 730
rect 2455 725 2459 726
rect 2456 706 2458 725
rect 2464 724 2466 750
rect 2472 736 2474 806
rect 2502 795 2508 796
rect 2502 791 2503 795
rect 2507 791 2508 795
rect 2502 790 2508 791
rect 2504 783 2506 790
rect 2503 782 2507 783
rect 2503 777 2507 778
rect 2504 774 2506 777
rect 2502 773 2508 774
rect 2502 769 2503 773
rect 2507 769 2508 773
rect 2502 768 2508 769
rect 2502 756 2508 757
rect 2502 752 2503 756
rect 2507 752 2508 756
rect 2502 751 2508 752
rect 2470 735 2476 736
rect 2470 731 2471 735
rect 2475 731 2476 735
rect 2504 731 2506 751
rect 2470 730 2476 731
rect 2503 730 2507 731
rect 2503 725 2507 726
rect 2462 723 2468 724
rect 2462 719 2463 723
rect 2467 719 2468 723
rect 2462 718 2468 719
rect 2454 705 2460 706
rect 2504 705 2506 725
rect 2366 700 2372 701
rect 2386 703 2392 704
rect 2278 698 2284 699
rect 2386 699 2387 703
rect 2391 699 2392 703
rect 2454 701 2455 705
rect 2459 701 2460 705
rect 2502 704 2508 705
rect 2454 700 2460 701
rect 2470 703 2476 704
rect 2386 698 2392 699
rect 2470 699 2471 703
rect 2475 699 2476 703
rect 2502 700 2503 704
rect 2507 700 2508 704
rect 2502 699 2508 700
rect 2470 698 2476 699
rect 1926 684 1932 685
rect 1926 680 1927 684
rect 1931 680 1932 684
rect 1926 679 1932 680
rect 2030 684 2036 685
rect 2030 680 2031 684
rect 2035 680 2036 684
rect 2030 679 2036 680
rect 1928 667 1930 679
rect 2032 667 2034 679
rect 1927 666 1931 667
rect 1927 661 1931 662
rect 1935 666 1939 667
rect 1935 661 1939 662
rect 2031 666 2035 667
rect 2031 661 2035 662
rect 2055 666 2059 667
rect 2055 661 2059 662
rect 1934 660 1940 661
rect 1934 656 1935 660
rect 1939 656 1940 660
rect 1934 655 1940 656
rect 2054 660 2060 661
rect 2054 656 2055 660
rect 2059 656 2060 660
rect 2054 655 2060 656
rect 1366 639 1372 640
rect 1366 635 1367 639
rect 1371 635 1372 639
rect 1366 634 1372 635
rect 1410 639 1416 640
rect 1410 635 1411 639
rect 1415 635 1416 639
rect 1410 634 1416 635
rect 1430 639 1436 640
rect 1430 635 1431 639
rect 1435 635 1436 639
rect 1430 634 1436 635
rect 1506 639 1512 640
rect 1506 635 1507 639
rect 1511 635 1512 639
rect 1506 634 1512 635
rect 1526 639 1532 640
rect 1526 635 1527 639
rect 1531 635 1532 639
rect 1526 634 1532 635
rect 1534 639 1540 640
rect 1534 635 1535 639
rect 1539 635 1540 639
rect 1534 634 1540 635
rect 1622 639 1628 640
rect 1622 635 1623 639
rect 1627 635 1628 639
rect 1622 634 1628 635
rect 1726 639 1732 640
rect 1726 635 1727 639
rect 1731 635 1732 639
rect 1726 634 1732 635
rect 1838 639 1844 640
rect 1838 635 1839 639
rect 1843 635 1844 639
rect 1838 634 1844 635
rect 1854 639 1860 640
rect 1854 635 1855 639
rect 1859 635 1860 639
rect 1854 634 1860 635
rect 1950 639 1956 640
rect 1950 635 1951 639
rect 1955 635 1956 639
rect 1950 634 1956 635
rect 1342 619 1348 620
rect 1342 615 1343 619
rect 1347 615 1348 619
rect 1368 615 1370 634
rect 1412 620 1414 634
rect 1410 619 1416 620
rect 1410 615 1411 619
rect 1415 615 1416 619
rect 1432 615 1434 634
rect 1508 620 1510 634
rect 1506 619 1512 620
rect 1506 615 1507 619
rect 1511 615 1512 619
rect 1528 615 1530 634
rect 1536 616 1538 634
rect 1534 615 1540 616
rect 1624 615 1626 634
rect 1728 615 1730 634
rect 1762 619 1768 620
rect 1762 615 1763 619
rect 1767 615 1768 619
rect 1840 615 1842 634
rect 1952 615 1954 634
rect 2064 620 2066 698
rect 2134 684 2140 685
rect 2134 680 2135 684
rect 2139 680 2140 684
rect 2134 679 2140 680
rect 2238 684 2244 685
rect 2238 680 2239 684
rect 2243 680 2244 684
rect 2238 679 2244 680
rect 2350 684 2356 685
rect 2350 680 2351 684
rect 2355 680 2356 684
rect 2350 679 2356 680
rect 2438 684 2444 685
rect 2438 680 2439 684
rect 2443 680 2444 684
rect 2438 679 2444 680
rect 2136 667 2138 679
rect 2240 667 2242 679
rect 2352 667 2354 679
rect 2440 667 2442 679
rect 2135 666 2139 667
rect 2135 661 2139 662
rect 2183 666 2187 667
rect 2183 661 2187 662
rect 2239 666 2243 667
rect 2239 661 2243 662
rect 2319 666 2323 667
rect 2319 661 2323 662
rect 2351 666 2355 667
rect 2351 661 2355 662
rect 2439 666 2443 667
rect 2439 661 2443 662
rect 2182 660 2188 661
rect 2182 656 2183 660
rect 2187 656 2188 660
rect 2182 655 2188 656
rect 2318 660 2324 661
rect 2318 656 2319 660
rect 2323 656 2324 660
rect 2318 655 2324 656
rect 2438 660 2444 661
rect 2438 656 2439 660
rect 2443 656 2444 660
rect 2438 655 2444 656
rect 2070 639 2076 640
rect 2070 635 2071 639
rect 2075 635 2076 639
rect 2070 634 2076 635
rect 2178 639 2184 640
rect 2178 635 2179 639
rect 2183 635 2184 639
rect 2178 634 2184 635
rect 2198 639 2204 640
rect 2198 635 2199 639
rect 2203 635 2204 639
rect 2198 634 2204 635
rect 2314 639 2320 640
rect 2314 635 2315 639
rect 2319 635 2320 639
rect 2314 634 2320 635
rect 2334 639 2340 640
rect 2334 635 2335 639
rect 2339 635 2340 639
rect 2334 634 2340 635
rect 2350 639 2356 640
rect 2350 635 2351 639
rect 2355 635 2356 639
rect 2350 634 2356 635
rect 2454 639 2460 640
rect 2454 635 2455 639
rect 2459 635 2460 639
rect 2454 634 2460 635
rect 2462 639 2468 640
rect 2462 635 2463 639
rect 2467 635 2468 639
rect 2462 634 2468 635
rect 2042 619 2048 620
rect 2042 615 2043 619
rect 2047 615 2048 619
rect 1327 614 1331 615
rect 1342 614 1348 615
rect 1367 614 1371 615
rect 1327 609 1331 610
rect 1367 609 1371 610
rect 1383 614 1387 615
rect 1410 614 1416 615
rect 1431 614 1435 615
rect 1383 609 1387 610
rect 1431 609 1435 610
rect 1463 614 1467 615
rect 1506 614 1512 615
rect 1527 614 1531 615
rect 1463 609 1467 610
rect 1534 611 1535 615
rect 1539 611 1540 615
rect 1534 610 1540 611
rect 1551 614 1555 615
rect 1527 609 1531 610
rect 1551 609 1555 610
rect 1623 614 1627 615
rect 1623 609 1627 610
rect 1647 614 1651 615
rect 1647 609 1651 610
rect 1727 614 1731 615
rect 1727 609 1731 610
rect 1743 614 1747 615
rect 1762 614 1768 615
rect 1839 614 1843 615
rect 1743 609 1747 610
rect 1183 598 1187 599
rect 1183 593 1187 594
rect 1239 598 1243 599
rect 1262 598 1268 599
rect 1287 598 1291 599
rect 1239 593 1243 594
rect 1287 593 1291 594
rect 1166 591 1172 592
rect 1166 587 1167 591
rect 1171 587 1172 591
rect 1166 586 1172 587
rect 1184 574 1186 593
rect 1086 573 1092 574
rect 998 568 1004 569
rect 1018 571 1024 572
rect 942 566 948 567
rect 1018 567 1019 571
rect 1023 567 1024 571
rect 1086 569 1087 573
rect 1091 569 1092 573
rect 1086 568 1092 569
rect 1182 573 1188 574
rect 1288 573 1290 593
rect 1328 589 1330 609
rect 1384 590 1386 609
rect 1464 590 1466 609
rect 1552 590 1554 609
rect 1574 607 1580 608
rect 1574 603 1575 607
rect 1579 603 1580 607
rect 1574 602 1580 603
rect 1382 589 1388 590
rect 1326 588 1332 589
rect 1326 584 1327 588
rect 1331 584 1332 588
rect 1382 585 1383 589
rect 1387 585 1388 589
rect 1462 589 1468 590
rect 1382 584 1388 585
rect 1398 587 1404 588
rect 1326 583 1332 584
rect 1398 583 1399 587
rect 1403 583 1404 587
rect 1462 585 1463 589
rect 1467 585 1468 589
rect 1462 584 1468 585
rect 1550 589 1556 590
rect 1550 585 1551 589
rect 1555 585 1556 589
rect 1576 588 1578 602
rect 1586 599 1592 600
rect 1586 595 1587 599
rect 1591 595 1592 599
rect 1586 594 1592 595
rect 1550 584 1556 585
rect 1574 587 1580 588
rect 1398 582 1404 583
rect 1574 583 1575 587
rect 1579 583 1580 587
rect 1574 582 1580 583
rect 1182 569 1183 573
rect 1187 569 1188 573
rect 1182 568 1188 569
rect 1286 572 1292 573
rect 1286 568 1287 572
rect 1291 568 1292 572
rect 1286 567 1292 568
rect 1326 571 1332 572
rect 1326 567 1327 571
rect 1331 567 1332 571
rect 1018 566 1024 567
rect 1326 566 1332 567
rect 1366 568 1372 569
rect 806 552 812 553
rect 806 548 807 552
rect 811 548 812 552
rect 806 547 812 548
rect 894 552 900 553
rect 894 548 895 552
rect 899 548 900 552
rect 894 547 900 548
rect 808 539 810 547
rect 896 539 898 547
rect 791 538 795 539
rect 791 533 795 534
rect 807 538 811 539
rect 807 533 811 534
rect 871 538 875 539
rect 871 533 875 534
rect 895 538 899 539
rect 895 533 899 534
rect 790 532 796 533
rect 790 528 791 532
rect 795 528 796 532
rect 790 527 796 528
rect 870 532 876 533
rect 870 528 871 532
rect 875 528 876 532
rect 870 527 876 528
rect 706 511 712 512
rect 706 507 707 511
rect 711 507 712 511
rect 706 506 712 507
rect 726 511 732 512
rect 726 507 727 511
rect 731 507 732 511
rect 726 506 732 507
rect 742 511 748 512
rect 742 507 743 511
rect 747 507 748 511
rect 742 506 748 507
rect 806 511 812 512
rect 806 507 807 511
rect 811 507 812 511
rect 806 506 812 507
rect 826 511 832 512
rect 826 507 827 511
rect 831 507 832 511
rect 826 506 832 507
rect 886 511 892 512
rect 886 507 887 511
rect 891 507 892 511
rect 886 506 892 507
rect 646 499 652 500
rect 646 495 647 499
rect 651 495 652 499
rect 646 494 652 495
rect 708 492 710 506
rect 674 491 680 492
rect 674 487 675 491
rect 679 487 680 491
rect 674 486 680 487
rect 706 491 712 492
rect 706 487 707 491
rect 711 487 712 491
rect 706 486 712 487
rect 463 482 467 483
rect 463 477 467 478
rect 543 482 547 483
rect 543 477 547 478
rect 559 482 563 483
rect 578 479 579 483
rect 583 479 584 483
rect 578 478 584 479
rect 639 482 643 483
rect 559 477 563 478
rect 454 475 460 476
rect 454 471 455 475
rect 459 471 460 475
rect 454 470 460 471
rect 464 458 466 477
rect 486 475 492 476
rect 486 471 487 475
rect 491 471 492 475
rect 486 470 492 471
rect 374 457 380 458
rect 310 455 316 456
rect 310 451 311 455
rect 315 451 316 455
rect 374 453 375 457
rect 379 453 380 457
rect 462 457 468 458
rect 374 452 380 453
rect 390 455 396 456
rect 310 450 316 451
rect 390 451 391 455
rect 395 451 396 455
rect 462 453 463 457
rect 467 453 468 457
rect 488 456 490 470
rect 560 458 562 477
rect 558 457 564 458
rect 462 452 468 453
rect 486 455 492 456
rect 390 450 396 451
rect 486 451 487 455
rect 491 451 492 455
rect 558 453 559 457
rect 563 453 564 457
rect 580 456 582 478
rect 639 477 643 478
rect 655 482 659 483
rect 655 477 659 478
rect 656 458 658 477
rect 654 457 660 458
rect 558 452 564 453
rect 578 455 584 456
rect 486 450 492 451
rect 578 451 579 455
rect 583 451 584 455
rect 654 453 655 457
rect 659 453 660 457
rect 676 456 678 486
rect 728 483 730 506
rect 808 483 810 506
rect 727 482 731 483
rect 727 477 731 478
rect 751 482 755 483
rect 751 477 755 478
rect 807 482 811 483
rect 807 477 811 478
rect 742 475 748 476
rect 742 471 743 475
rect 747 471 748 475
rect 742 470 748 471
rect 654 452 660 453
rect 674 455 680 456
rect 578 450 584 451
rect 674 451 675 455
rect 679 451 680 455
rect 674 450 680 451
rect 358 436 364 437
rect 358 432 359 436
rect 363 432 364 436
rect 358 431 364 432
rect 359 430 363 431
rect 359 425 363 426
rect 383 430 387 431
rect 383 425 387 426
rect 382 424 388 425
rect 382 420 383 424
rect 387 420 388 424
rect 382 419 388 420
rect 110 400 111 404
rect 115 400 116 404
rect 110 399 116 400
rect 150 403 156 404
rect 150 399 151 403
rect 155 399 156 403
rect 112 375 114 399
rect 150 398 156 399
rect 186 403 192 404
rect 186 399 187 403
rect 191 399 192 403
rect 186 398 192 399
rect 206 403 212 404
rect 206 399 207 403
rect 211 399 212 403
rect 206 398 212 399
rect 274 403 280 404
rect 274 399 275 403
rect 279 399 280 403
rect 274 398 280 399
rect 294 403 300 404
rect 294 399 295 403
rect 299 399 300 403
rect 294 398 300 399
rect 302 403 308 404
rect 302 399 303 403
rect 307 399 308 403
rect 302 398 308 399
rect 152 375 154 398
rect 188 384 190 398
rect 170 383 176 384
rect 170 379 171 383
rect 175 379 176 383
rect 170 378 176 379
rect 186 383 192 384
rect 186 379 187 383
rect 191 379 192 383
rect 186 378 192 379
rect 111 374 115 375
rect 111 369 115 370
rect 151 374 155 375
rect 151 369 155 370
rect 112 349 114 369
rect 152 350 154 369
rect 150 349 156 350
rect 110 348 116 349
rect 110 344 111 348
rect 115 344 116 348
rect 150 345 151 349
rect 155 345 156 349
rect 172 348 174 378
rect 208 375 210 398
rect 276 384 278 398
rect 274 383 280 384
rect 274 379 275 383
rect 279 379 280 383
rect 274 378 280 379
rect 296 375 298 398
rect 392 384 394 450
rect 446 436 452 437
rect 446 432 447 436
rect 451 432 452 436
rect 446 431 452 432
rect 542 436 548 437
rect 542 432 543 436
rect 547 432 548 436
rect 542 431 548 432
rect 638 436 644 437
rect 638 432 639 436
rect 643 432 644 436
rect 638 431 644 432
rect 734 436 740 437
rect 734 432 735 436
rect 739 432 740 436
rect 734 431 740 432
rect 447 430 451 431
rect 447 425 451 426
rect 495 430 499 431
rect 495 425 499 426
rect 543 430 547 431
rect 543 425 547 426
rect 607 430 611 431
rect 607 425 611 426
rect 639 430 643 431
rect 639 425 643 426
rect 719 430 723 431
rect 719 425 723 426
rect 735 430 739 431
rect 735 425 739 426
rect 494 424 500 425
rect 494 420 495 424
rect 499 420 500 424
rect 494 419 500 420
rect 606 424 612 425
rect 606 420 607 424
rect 611 420 612 424
rect 606 419 612 420
rect 718 424 724 425
rect 718 420 719 424
rect 723 420 724 424
rect 718 419 724 420
rect 744 404 746 470
rect 752 458 754 477
rect 828 476 830 506
rect 888 483 890 506
rect 944 492 946 566
rect 1328 563 1330 566
rect 1366 564 1367 568
rect 1371 564 1372 568
rect 1366 563 1372 564
rect 1327 562 1331 563
rect 1327 557 1331 558
rect 1367 562 1371 563
rect 1367 557 1371 558
rect 1375 562 1379 563
rect 1375 557 1379 558
rect 1286 555 1292 556
rect 982 552 988 553
rect 982 548 983 552
rect 987 548 988 552
rect 982 547 988 548
rect 1070 552 1076 553
rect 1070 548 1071 552
rect 1075 548 1076 552
rect 1070 547 1076 548
rect 1166 552 1172 553
rect 1166 548 1167 552
rect 1171 548 1172 552
rect 1286 551 1287 555
rect 1291 551 1292 555
rect 1328 554 1330 557
rect 1374 556 1380 557
rect 1286 550 1292 551
rect 1326 553 1332 554
rect 1166 547 1172 548
rect 984 539 986 547
rect 1072 539 1074 547
rect 1168 539 1170 547
rect 1288 539 1290 550
rect 1326 549 1327 553
rect 1331 549 1332 553
rect 1374 552 1375 556
rect 1379 552 1380 556
rect 1374 551 1380 552
rect 1326 548 1332 549
rect 951 538 955 539
rect 951 533 955 534
rect 983 538 987 539
rect 983 533 987 534
rect 1031 538 1035 539
rect 1031 533 1035 534
rect 1071 538 1075 539
rect 1071 533 1075 534
rect 1167 538 1171 539
rect 1167 533 1171 534
rect 1287 538 1291 539
rect 1287 533 1291 534
rect 1326 536 1332 537
rect 950 532 956 533
rect 950 528 951 532
rect 955 528 956 532
rect 950 527 956 528
rect 1030 532 1036 533
rect 1030 528 1031 532
rect 1035 528 1036 532
rect 1288 530 1290 533
rect 1326 532 1327 536
rect 1331 532 1332 536
rect 1326 531 1332 532
rect 1390 535 1396 536
rect 1390 531 1391 535
rect 1395 531 1396 535
rect 1030 527 1036 528
rect 1286 529 1292 530
rect 1286 525 1287 529
rect 1291 525 1292 529
rect 1286 524 1292 525
rect 1286 512 1292 513
rect 966 511 972 512
rect 966 507 967 511
rect 971 507 972 511
rect 966 506 972 507
rect 1026 511 1032 512
rect 1026 507 1027 511
rect 1031 507 1032 511
rect 1026 506 1032 507
rect 1046 511 1052 512
rect 1046 507 1047 511
rect 1051 507 1052 511
rect 1286 508 1287 512
rect 1291 508 1292 512
rect 1286 507 1292 508
rect 1328 507 1330 531
rect 1390 530 1396 531
rect 1392 507 1394 530
rect 1400 516 1402 582
rect 1446 568 1452 569
rect 1446 564 1447 568
rect 1451 564 1452 568
rect 1446 563 1452 564
rect 1534 568 1540 569
rect 1534 564 1535 568
rect 1539 564 1540 568
rect 1534 563 1540 564
rect 1447 562 1451 563
rect 1447 557 1451 558
rect 1455 562 1459 563
rect 1455 557 1459 558
rect 1535 562 1539 563
rect 1535 557 1539 558
rect 1551 562 1555 563
rect 1551 557 1555 558
rect 1454 556 1460 557
rect 1454 552 1455 556
rect 1459 552 1460 556
rect 1454 551 1460 552
rect 1550 556 1556 557
rect 1550 552 1551 556
rect 1555 552 1556 556
rect 1550 551 1556 552
rect 1588 536 1590 594
rect 1648 590 1650 609
rect 1744 590 1746 609
rect 1646 589 1652 590
rect 1646 585 1647 589
rect 1651 585 1652 589
rect 1646 584 1652 585
rect 1742 589 1748 590
rect 1742 585 1743 589
rect 1747 585 1748 589
rect 1764 588 1766 614
rect 1839 609 1843 610
rect 1847 614 1851 615
rect 1847 609 1851 610
rect 1951 614 1955 615
rect 1951 609 1955 610
rect 1959 614 1963 615
rect 2042 614 2048 615
rect 2062 619 2068 620
rect 2062 615 2063 619
rect 2067 615 2068 619
rect 2072 615 2074 634
rect 2180 620 2182 634
rect 2178 619 2184 620
rect 2178 615 2179 619
rect 2183 615 2184 619
rect 2200 615 2202 634
rect 2316 620 2318 634
rect 2314 619 2320 620
rect 2314 615 2315 619
rect 2319 615 2320 619
rect 2336 615 2338 634
rect 2062 614 2068 615
rect 2071 614 2075 615
rect 1959 609 1963 610
rect 1848 590 1850 609
rect 1870 607 1876 608
rect 1870 603 1871 607
rect 1875 603 1876 607
rect 1870 602 1876 603
rect 1846 589 1852 590
rect 1742 584 1748 585
rect 1762 587 1768 588
rect 1762 583 1763 587
rect 1767 583 1768 587
rect 1846 585 1847 589
rect 1851 585 1852 589
rect 1872 588 1874 602
rect 1890 599 1896 600
rect 1890 595 1891 599
rect 1895 595 1896 599
rect 1890 594 1896 595
rect 1846 584 1852 585
rect 1870 587 1876 588
rect 1762 582 1768 583
rect 1870 583 1871 587
rect 1875 583 1876 587
rect 1870 582 1876 583
rect 1630 568 1636 569
rect 1630 564 1631 568
rect 1635 564 1636 568
rect 1630 563 1636 564
rect 1726 568 1732 569
rect 1726 564 1727 568
rect 1731 564 1732 568
rect 1726 563 1732 564
rect 1830 568 1836 569
rect 1830 564 1831 568
rect 1835 564 1836 568
rect 1830 563 1836 564
rect 1631 562 1635 563
rect 1631 557 1635 558
rect 1647 562 1651 563
rect 1647 557 1651 558
rect 1727 562 1731 563
rect 1727 557 1731 558
rect 1751 562 1755 563
rect 1751 557 1755 558
rect 1831 562 1835 563
rect 1831 557 1835 558
rect 1855 562 1859 563
rect 1855 557 1859 558
rect 1646 556 1652 557
rect 1646 552 1647 556
rect 1651 552 1652 556
rect 1646 551 1652 552
rect 1750 556 1756 557
rect 1750 552 1751 556
rect 1755 552 1756 556
rect 1750 551 1756 552
rect 1854 556 1860 557
rect 1854 552 1855 556
rect 1859 552 1860 556
rect 1854 551 1860 552
rect 1892 536 1894 594
rect 1960 590 1962 609
rect 1982 607 1988 608
rect 1982 603 1983 607
rect 1987 603 1988 607
rect 1982 602 1988 603
rect 1958 589 1964 590
rect 1958 585 1959 589
rect 1963 585 1964 589
rect 1984 588 1986 602
rect 2044 596 2046 614
rect 2071 609 2075 610
rect 2079 614 2083 615
rect 2178 614 2184 615
rect 2199 614 2203 615
rect 2079 609 2083 610
rect 2199 609 2203 610
rect 2207 614 2211 615
rect 2314 614 2320 615
rect 2335 614 2339 615
rect 2207 609 2211 610
rect 2335 609 2339 610
rect 2343 614 2347 615
rect 2343 609 2347 610
rect 2042 595 2048 596
rect 2042 591 2043 595
rect 2047 591 2048 595
rect 2042 590 2048 591
rect 2080 590 2082 609
rect 2208 590 2210 609
rect 2344 590 2346 609
rect 2352 608 2354 634
rect 2456 615 2458 634
rect 2455 614 2459 615
rect 2455 609 2459 610
rect 2350 607 2356 608
rect 2350 603 2351 607
rect 2355 603 2356 607
rect 2350 602 2356 603
rect 2456 590 2458 609
rect 2464 608 2466 634
rect 2472 620 2474 698
rect 2502 687 2508 688
rect 2502 683 2503 687
rect 2507 683 2508 687
rect 2502 682 2508 683
rect 2504 667 2506 682
rect 2503 666 2507 667
rect 2503 661 2507 662
rect 2504 658 2506 661
rect 2502 657 2508 658
rect 2502 653 2503 657
rect 2507 653 2508 657
rect 2502 652 2508 653
rect 2502 640 2508 641
rect 2502 636 2503 640
rect 2507 636 2508 640
rect 2502 635 2508 636
rect 2470 619 2476 620
rect 2470 615 2471 619
rect 2475 615 2476 619
rect 2504 615 2506 635
rect 2470 614 2476 615
rect 2503 614 2507 615
rect 2503 609 2507 610
rect 2462 607 2468 608
rect 2462 603 2463 607
rect 2467 603 2468 607
rect 2462 602 2468 603
rect 2078 589 2084 590
rect 1958 584 1964 585
rect 1982 587 1988 588
rect 1982 583 1983 587
rect 1987 583 1988 587
rect 2078 585 2079 589
rect 2083 585 2084 589
rect 2078 584 2084 585
rect 2206 589 2212 590
rect 2206 585 2207 589
rect 2211 585 2212 589
rect 2342 589 2348 590
rect 2206 584 2212 585
rect 2214 587 2220 588
rect 1982 582 1988 583
rect 2214 583 2215 587
rect 2219 583 2220 587
rect 2342 585 2343 589
rect 2347 585 2348 589
rect 2342 584 2348 585
rect 2454 589 2460 590
rect 2504 589 2506 609
rect 2454 585 2455 589
rect 2459 585 2460 589
rect 2502 588 2508 589
rect 2454 584 2460 585
rect 2462 587 2468 588
rect 2214 582 2220 583
rect 2462 583 2463 587
rect 2467 583 2468 587
rect 2502 584 2503 588
rect 2507 584 2508 588
rect 2502 583 2508 584
rect 2462 582 2468 583
rect 1942 568 1948 569
rect 1942 564 1943 568
rect 1947 564 1948 568
rect 1942 563 1948 564
rect 2062 568 2068 569
rect 2062 564 2063 568
rect 2067 564 2068 568
rect 2062 563 2068 564
rect 2190 568 2196 569
rect 2190 564 2191 568
rect 2195 564 2196 568
rect 2190 563 2196 564
rect 1943 562 1947 563
rect 1943 557 1947 558
rect 1959 562 1963 563
rect 1959 557 1963 558
rect 2055 562 2059 563
rect 2055 557 2059 558
rect 2063 562 2067 563
rect 2063 557 2067 558
rect 2151 562 2155 563
rect 2151 557 2155 558
rect 2191 562 2195 563
rect 2191 557 2195 558
rect 1958 556 1964 557
rect 1958 552 1959 556
rect 1963 552 1964 556
rect 1958 551 1964 552
rect 2054 556 2060 557
rect 2054 552 2055 556
rect 2059 552 2060 556
rect 2054 551 2060 552
rect 2150 556 2156 557
rect 2150 552 2151 556
rect 2155 552 2156 556
rect 2150 551 2156 552
rect 1450 535 1456 536
rect 1450 531 1451 535
rect 1455 531 1456 535
rect 1450 530 1456 531
rect 1470 535 1476 536
rect 1470 531 1471 535
rect 1475 531 1476 535
rect 1470 530 1476 531
rect 1478 535 1484 536
rect 1478 531 1479 535
rect 1483 531 1484 535
rect 1478 530 1484 531
rect 1566 535 1572 536
rect 1566 531 1567 535
rect 1571 531 1572 535
rect 1566 530 1572 531
rect 1586 535 1592 536
rect 1586 531 1587 535
rect 1591 531 1592 535
rect 1586 530 1592 531
rect 1662 535 1668 536
rect 1662 531 1663 535
rect 1667 531 1668 535
rect 1662 530 1668 531
rect 1766 535 1772 536
rect 1766 531 1767 535
rect 1771 531 1772 535
rect 1766 530 1772 531
rect 1870 535 1876 536
rect 1870 531 1871 535
rect 1875 531 1876 535
rect 1870 530 1876 531
rect 1890 535 1896 536
rect 1890 531 1891 535
rect 1895 531 1896 535
rect 1890 530 1896 531
rect 1974 535 1980 536
rect 1974 531 1975 535
rect 1979 531 1980 535
rect 1974 530 1980 531
rect 2070 535 2076 536
rect 2070 531 2071 535
rect 2075 531 2076 535
rect 2070 530 2076 531
rect 2146 535 2152 536
rect 2146 531 2147 535
rect 2151 531 2152 535
rect 2146 530 2152 531
rect 2166 535 2172 536
rect 2166 531 2167 535
rect 2171 531 2172 535
rect 2166 530 2172 531
rect 1452 516 1454 530
rect 1398 515 1404 516
rect 1398 511 1399 515
rect 1403 511 1404 515
rect 1398 510 1404 511
rect 1450 515 1456 516
rect 1450 511 1451 515
rect 1455 511 1456 515
rect 1450 510 1456 511
rect 1472 507 1474 530
rect 1046 506 1052 507
rect 942 491 948 492
rect 942 487 943 491
rect 947 487 948 491
rect 942 486 948 487
rect 968 483 970 506
rect 1028 492 1030 506
rect 1026 491 1032 492
rect 1026 487 1027 491
rect 1031 487 1032 491
rect 1026 486 1032 487
rect 1048 483 1050 506
rect 1288 483 1290 507
rect 1327 506 1331 507
rect 1327 501 1331 502
rect 1367 506 1371 507
rect 1367 501 1371 502
rect 1391 506 1395 507
rect 1391 501 1395 502
rect 1455 506 1459 507
rect 1455 501 1459 502
rect 1471 506 1475 507
rect 1471 501 1475 502
rect 847 482 851 483
rect 847 477 851 478
rect 887 482 891 483
rect 887 477 891 478
rect 951 482 955 483
rect 951 477 955 478
rect 967 482 971 483
rect 967 477 971 478
rect 1047 482 1051 483
rect 1047 477 1051 478
rect 1055 482 1059 483
rect 1055 477 1059 478
rect 1159 482 1163 483
rect 1159 477 1163 478
rect 1239 482 1243 483
rect 1239 477 1243 478
rect 1287 482 1291 483
rect 1328 481 1330 501
rect 1368 482 1370 501
rect 1456 482 1458 501
rect 1480 500 1482 530
rect 1568 507 1570 530
rect 1664 507 1666 530
rect 1768 507 1770 530
rect 1826 515 1832 516
rect 1826 511 1827 515
rect 1831 511 1832 515
rect 1826 510 1832 511
rect 1567 506 1571 507
rect 1567 501 1571 502
rect 1575 506 1579 507
rect 1575 501 1579 502
rect 1663 506 1667 507
rect 1663 501 1667 502
rect 1695 506 1699 507
rect 1695 501 1699 502
rect 1767 506 1771 507
rect 1767 501 1771 502
rect 1807 506 1811 507
rect 1807 501 1811 502
rect 1478 499 1484 500
rect 1478 495 1479 499
rect 1483 495 1484 499
rect 1478 494 1484 495
rect 1576 482 1578 501
rect 1598 499 1604 500
rect 1598 495 1599 499
rect 1603 495 1604 499
rect 1598 494 1604 495
rect 1366 481 1372 482
rect 1287 477 1291 478
rect 1326 480 1332 481
rect 826 475 832 476
rect 826 471 827 475
rect 831 471 832 475
rect 826 470 832 471
rect 838 463 844 464
rect 838 459 839 463
rect 843 459 844 463
rect 838 458 844 459
rect 848 458 850 477
rect 870 475 876 476
rect 870 471 871 475
rect 875 471 876 475
rect 870 470 876 471
rect 750 457 756 458
rect 750 453 751 457
rect 755 453 756 457
rect 750 452 756 453
rect 830 436 836 437
rect 830 432 831 436
rect 835 432 836 436
rect 830 431 836 432
rect 831 430 835 431
rect 831 425 835 426
rect 830 424 836 425
rect 830 420 831 424
rect 835 420 836 424
rect 830 419 836 420
rect 398 403 404 404
rect 398 399 399 403
rect 403 399 404 403
rect 398 398 404 399
rect 490 403 496 404
rect 490 399 491 403
rect 495 399 496 403
rect 490 398 496 399
rect 510 403 516 404
rect 510 399 511 403
rect 515 399 516 403
rect 510 398 516 399
rect 602 403 608 404
rect 602 399 603 403
rect 607 399 608 403
rect 602 398 608 399
rect 622 403 628 404
rect 622 399 623 403
rect 627 399 628 403
rect 622 398 628 399
rect 630 403 636 404
rect 630 399 631 403
rect 635 399 636 403
rect 630 398 636 399
rect 734 403 740 404
rect 734 399 735 403
rect 739 399 740 403
rect 734 398 740 399
rect 742 403 748 404
rect 742 399 743 403
rect 747 399 748 403
rect 742 398 748 399
rect 390 383 396 384
rect 390 379 391 383
rect 395 379 396 383
rect 390 378 396 379
rect 400 375 402 398
rect 492 384 494 398
rect 490 383 496 384
rect 490 379 491 383
rect 495 379 496 383
rect 490 378 496 379
rect 512 375 514 398
rect 604 384 606 398
rect 602 383 608 384
rect 602 379 603 383
rect 607 379 608 383
rect 602 378 608 379
rect 624 375 626 398
rect 632 376 634 398
rect 630 375 636 376
rect 736 375 738 398
rect 840 384 842 458
rect 846 457 852 458
rect 846 453 847 457
rect 851 453 852 457
rect 872 456 874 470
rect 952 458 954 477
rect 974 475 980 476
rect 974 471 975 475
rect 979 471 980 475
rect 974 470 980 471
rect 950 457 956 458
rect 846 452 852 453
rect 870 455 876 456
rect 870 451 871 455
rect 875 451 876 455
rect 950 453 951 457
rect 955 453 956 457
rect 976 456 978 470
rect 1056 458 1058 477
rect 1160 458 1162 477
rect 1240 458 1242 477
rect 1054 457 1060 458
rect 950 452 956 453
rect 974 455 980 456
rect 870 450 876 451
rect 974 451 975 455
rect 979 451 980 455
rect 1054 453 1055 457
rect 1059 453 1060 457
rect 1054 452 1060 453
rect 1158 457 1164 458
rect 1158 453 1159 457
rect 1163 453 1164 457
rect 1238 457 1244 458
rect 1288 457 1290 477
rect 1326 476 1327 480
rect 1331 476 1332 480
rect 1366 477 1367 481
rect 1371 477 1372 481
rect 1366 476 1372 477
rect 1454 481 1460 482
rect 1454 477 1455 481
rect 1459 477 1460 481
rect 1454 476 1460 477
rect 1574 481 1580 482
rect 1574 477 1575 481
rect 1579 477 1580 481
rect 1600 480 1602 494
rect 1618 491 1624 492
rect 1618 487 1619 491
rect 1623 487 1624 491
rect 1618 486 1624 487
rect 1574 476 1580 477
rect 1598 479 1604 480
rect 1326 475 1332 476
rect 1598 475 1599 479
rect 1603 475 1604 479
rect 1598 474 1604 475
rect 1326 463 1332 464
rect 1326 459 1327 463
rect 1331 459 1332 463
rect 1326 458 1332 459
rect 1350 460 1356 461
rect 1158 452 1164 453
rect 1166 455 1172 456
rect 974 450 980 451
rect 1166 451 1167 455
rect 1171 451 1172 455
rect 1238 453 1239 457
rect 1243 453 1244 457
rect 1238 452 1244 453
rect 1286 456 1292 457
rect 1286 452 1287 456
rect 1291 452 1292 456
rect 1286 451 1292 452
rect 1166 450 1172 451
rect 934 436 940 437
rect 934 432 935 436
rect 939 432 940 436
rect 934 431 940 432
rect 1038 436 1044 437
rect 1038 432 1039 436
rect 1043 432 1044 436
rect 1038 431 1044 432
rect 1142 436 1148 437
rect 1142 432 1143 436
rect 1147 432 1148 436
rect 1142 431 1148 432
rect 935 430 939 431
rect 935 425 939 426
rect 1039 430 1043 431
rect 1039 425 1043 426
rect 1143 430 1147 431
rect 1143 425 1147 426
rect 934 424 940 425
rect 934 420 935 424
rect 939 420 940 424
rect 934 419 940 420
rect 1038 424 1044 425
rect 1038 420 1039 424
rect 1043 420 1044 424
rect 1038 419 1044 420
rect 1142 424 1148 425
rect 1142 420 1143 424
rect 1147 420 1148 424
rect 1142 419 1148 420
rect 846 403 852 404
rect 846 399 847 403
rect 851 399 852 403
rect 846 398 852 399
rect 930 403 936 404
rect 930 399 931 403
rect 935 399 936 403
rect 930 398 936 399
rect 950 403 956 404
rect 950 399 951 403
rect 955 399 956 403
rect 950 398 956 399
rect 994 403 1000 404
rect 994 399 995 403
rect 999 399 1000 403
rect 994 398 1000 399
rect 1054 403 1060 404
rect 1054 399 1055 403
rect 1059 399 1060 403
rect 1054 398 1060 399
rect 1074 403 1080 404
rect 1074 399 1075 403
rect 1079 399 1080 403
rect 1074 398 1080 399
rect 1158 403 1164 404
rect 1158 399 1159 403
rect 1163 399 1164 403
rect 1158 398 1164 399
rect 770 383 776 384
rect 770 379 771 383
rect 775 379 776 383
rect 770 378 776 379
rect 838 383 844 384
rect 838 379 839 383
rect 843 379 844 383
rect 838 378 844 379
rect 207 374 211 375
rect 207 369 211 370
rect 231 374 235 375
rect 231 369 235 370
rect 295 374 299 375
rect 295 369 299 370
rect 335 374 339 375
rect 335 369 339 370
rect 399 374 403 375
rect 399 369 403 370
rect 439 374 443 375
rect 439 369 443 370
rect 511 374 515 375
rect 511 369 515 370
rect 543 374 547 375
rect 543 369 547 370
rect 623 374 627 375
rect 630 371 631 375
rect 635 371 636 375
rect 630 370 636 371
rect 647 374 651 375
rect 623 369 627 370
rect 647 369 651 370
rect 735 374 739 375
rect 735 369 739 370
rect 751 374 755 375
rect 751 369 755 370
rect 232 350 234 369
rect 250 367 256 368
rect 250 363 251 367
rect 255 363 256 367
rect 250 362 256 363
rect 230 349 236 350
rect 150 344 156 345
rect 170 347 176 348
rect 110 343 116 344
rect 170 343 171 347
rect 175 343 176 347
rect 230 345 231 349
rect 235 345 236 349
rect 230 344 236 345
rect 170 342 176 343
rect 110 331 116 332
rect 110 327 111 331
rect 115 327 116 331
rect 110 326 116 327
rect 134 328 140 329
rect 112 319 114 326
rect 134 324 135 328
rect 139 324 140 328
rect 134 323 140 324
rect 214 328 220 329
rect 214 324 215 328
rect 219 324 220 328
rect 214 323 220 324
rect 136 319 138 323
rect 216 319 218 323
rect 111 318 115 319
rect 111 313 115 314
rect 135 318 139 319
rect 135 313 139 314
rect 215 318 219 319
rect 215 313 219 314
rect 112 310 114 313
rect 134 312 140 313
rect 110 309 116 310
rect 110 305 111 309
rect 115 305 116 309
rect 134 308 135 312
rect 139 308 140 312
rect 134 307 140 308
rect 214 312 220 313
rect 214 308 215 312
rect 219 308 220 312
rect 214 307 220 308
rect 110 304 116 305
rect 110 292 116 293
rect 252 292 254 362
rect 336 350 338 369
rect 358 367 364 368
rect 358 363 359 367
rect 363 363 364 367
rect 358 362 364 363
rect 334 349 340 350
rect 334 345 335 349
rect 339 345 340 349
rect 360 348 362 362
rect 440 350 442 369
rect 462 367 468 368
rect 462 363 463 367
rect 467 363 468 367
rect 462 362 468 363
rect 438 349 444 350
rect 334 344 340 345
rect 358 347 364 348
rect 358 343 359 347
rect 363 343 364 347
rect 438 345 439 349
rect 443 345 444 349
rect 464 348 466 362
rect 544 350 546 369
rect 648 350 650 369
rect 662 367 668 368
rect 662 363 663 367
rect 667 363 668 367
rect 662 362 668 363
rect 670 367 676 368
rect 670 363 671 367
rect 675 363 676 367
rect 670 362 676 363
rect 542 349 548 350
rect 438 344 444 345
rect 462 347 468 348
rect 358 342 364 343
rect 462 343 463 347
rect 467 343 468 347
rect 542 345 543 349
rect 547 345 548 349
rect 646 349 652 350
rect 542 344 548 345
rect 558 347 564 348
rect 462 342 468 343
rect 558 343 559 347
rect 563 343 564 347
rect 646 345 647 349
rect 651 345 652 349
rect 646 344 652 345
rect 558 342 564 343
rect 318 328 324 329
rect 318 324 319 328
rect 323 324 324 328
rect 318 323 324 324
rect 422 328 428 329
rect 422 324 423 328
rect 427 324 428 328
rect 422 323 428 324
rect 526 328 532 329
rect 526 324 527 328
rect 531 324 532 328
rect 526 323 532 324
rect 320 319 322 323
rect 424 319 426 323
rect 528 319 530 323
rect 319 318 323 319
rect 319 313 323 314
rect 423 318 427 319
rect 423 313 427 314
rect 527 318 531 319
rect 527 313 531 314
rect 535 318 539 319
rect 535 313 539 314
rect 318 312 324 313
rect 318 308 319 312
rect 323 308 324 312
rect 318 307 324 308
rect 422 312 428 313
rect 422 308 423 312
rect 427 308 428 312
rect 422 307 428 308
rect 534 312 540 313
rect 534 308 535 312
rect 539 308 540 312
rect 534 307 540 308
rect 110 288 111 292
rect 115 288 116 292
rect 110 287 116 288
rect 150 291 156 292
rect 150 287 151 291
rect 155 287 156 291
rect 112 267 114 287
rect 150 286 156 287
rect 210 291 216 292
rect 210 287 211 291
rect 215 287 216 291
rect 210 286 216 287
rect 230 291 236 292
rect 230 287 231 291
rect 235 287 236 291
rect 230 286 236 287
rect 250 291 256 292
rect 250 287 251 291
rect 255 287 256 291
rect 250 286 256 287
rect 334 291 340 292
rect 334 287 335 291
rect 339 287 340 291
rect 334 286 340 287
rect 402 291 408 292
rect 402 287 403 291
rect 407 287 408 291
rect 402 286 408 287
rect 438 291 444 292
rect 438 287 439 291
rect 443 287 444 291
rect 438 286 444 287
rect 550 291 556 292
rect 550 287 551 291
rect 555 287 556 291
rect 550 286 556 287
rect 152 267 154 286
rect 212 272 214 286
rect 170 271 176 272
rect 170 267 171 271
rect 175 267 176 271
rect 111 266 115 267
rect 111 261 115 262
rect 151 266 155 267
rect 170 266 176 267
rect 210 271 216 272
rect 210 267 211 271
rect 215 267 216 271
rect 232 267 234 286
rect 336 267 338 286
rect 210 266 216 267
rect 223 266 227 267
rect 151 261 155 262
rect 112 241 114 261
rect 152 242 154 261
rect 150 241 156 242
rect 110 240 116 241
rect 110 236 111 240
rect 115 236 116 240
rect 150 237 151 241
rect 155 237 156 241
rect 172 240 174 266
rect 223 261 227 262
rect 231 266 235 267
rect 231 261 235 262
rect 319 266 323 267
rect 319 261 323 262
rect 335 266 339 267
rect 335 261 339 262
rect 224 242 226 261
rect 310 259 316 260
rect 310 255 311 259
rect 315 255 316 259
rect 310 254 316 255
rect 222 241 228 242
rect 150 236 156 237
rect 170 239 176 240
rect 110 235 116 236
rect 170 235 171 239
rect 175 235 176 239
rect 222 237 223 241
rect 227 237 228 241
rect 222 236 228 237
rect 170 234 176 235
rect 110 223 116 224
rect 110 219 111 223
rect 115 219 116 223
rect 110 218 116 219
rect 134 220 140 221
rect 112 211 114 218
rect 134 216 135 220
rect 139 216 140 220
rect 134 215 140 216
rect 206 220 212 221
rect 206 216 207 220
rect 211 216 212 220
rect 206 215 212 216
rect 302 220 308 221
rect 302 216 303 220
rect 307 216 308 220
rect 302 215 308 216
rect 136 211 138 215
rect 208 211 210 215
rect 304 211 306 215
rect 111 210 115 211
rect 111 205 115 206
rect 135 210 139 211
rect 135 205 139 206
rect 183 210 187 211
rect 183 205 187 206
rect 207 210 211 211
rect 207 205 211 206
rect 279 210 283 211
rect 279 205 283 206
rect 303 210 307 211
rect 303 205 307 206
rect 112 202 114 205
rect 182 204 188 205
rect 110 201 116 202
rect 110 197 111 201
rect 115 197 116 201
rect 182 200 183 204
rect 187 200 188 204
rect 182 199 188 200
rect 278 204 284 205
rect 278 200 279 204
rect 283 200 284 204
rect 278 199 284 200
rect 110 196 116 197
rect 110 184 116 185
rect 312 184 314 254
rect 320 242 322 261
rect 404 260 406 286
rect 440 267 442 286
rect 552 267 554 286
rect 560 272 562 342
rect 630 328 636 329
rect 630 324 631 328
rect 635 324 636 328
rect 630 323 636 324
rect 632 319 634 323
rect 631 318 635 319
rect 631 313 635 314
rect 639 318 643 319
rect 639 313 643 314
rect 638 312 644 313
rect 638 308 639 312
rect 643 308 644 312
rect 638 307 644 308
rect 664 292 666 362
rect 672 348 674 362
rect 752 350 754 369
rect 750 349 756 350
rect 670 347 676 348
rect 670 343 671 347
rect 675 343 676 347
rect 750 345 751 349
rect 755 345 756 349
rect 772 348 774 378
rect 848 375 850 398
rect 932 384 934 398
rect 930 383 936 384
rect 930 379 931 383
rect 935 379 936 383
rect 930 378 936 379
rect 952 375 954 398
rect 847 374 851 375
rect 847 369 851 370
rect 935 374 939 375
rect 935 369 939 370
rect 951 374 955 375
rect 951 369 955 370
rect 848 350 850 369
rect 870 367 876 368
rect 870 363 871 367
rect 875 363 876 367
rect 870 362 876 363
rect 846 349 852 350
rect 750 344 756 345
rect 770 347 776 348
rect 670 342 676 343
rect 770 343 771 347
rect 775 343 776 347
rect 846 345 847 349
rect 851 345 852 349
rect 872 348 874 362
rect 936 350 938 369
rect 996 368 998 398
rect 1056 375 1058 398
rect 1015 374 1019 375
rect 1015 369 1019 370
rect 1055 374 1059 375
rect 1055 369 1059 370
rect 994 367 1000 368
rect 994 363 995 367
rect 999 363 1000 367
rect 994 362 1000 363
rect 1016 350 1018 369
rect 1076 368 1078 398
rect 1160 375 1162 398
rect 1168 384 1170 450
rect 1328 443 1330 458
rect 1350 456 1351 460
rect 1355 456 1356 460
rect 1350 455 1356 456
rect 1438 460 1444 461
rect 1438 456 1439 460
rect 1443 456 1444 460
rect 1438 455 1444 456
rect 1558 460 1564 461
rect 1558 456 1559 460
rect 1563 456 1564 460
rect 1558 455 1564 456
rect 1352 443 1354 455
rect 1440 443 1442 455
rect 1560 443 1562 455
rect 1327 442 1331 443
rect 1286 439 1292 440
rect 1222 436 1228 437
rect 1222 432 1223 436
rect 1227 432 1228 436
rect 1286 435 1287 439
rect 1291 435 1292 439
rect 1327 437 1331 438
rect 1351 442 1355 443
rect 1351 437 1355 438
rect 1439 442 1443 443
rect 1439 437 1443 438
rect 1559 442 1563 443
rect 1559 437 1563 438
rect 1583 442 1587 443
rect 1583 437 1587 438
rect 1286 434 1292 435
rect 1328 434 1330 437
rect 1582 436 1588 437
rect 1222 431 1228 432
rect 1288 431 1290 434
rect 1326 433 1332 434
rect 1223 430 1227 431
rect 1223 425 1227 426
rect 1287 430 1291 431
rect 1326 429 1327 433
rect 1331 429 1332 433
rect 1582 432 1583 436
rect 1587 432 1588 436
rect 1582 431 1588 432
rect 1326 428 1332 429
rect 1287 425 1291 426
rect 1222 424 1228 425
rect 1222 420 1223 424
rect 1227 420 1228 424
rect 1288 422 1290 425
rect 1222 419 1228 420
rect 1286 421 1292 422
rect 1286 417 1287 421
rect 1291 417 1292 421
rect 1286 416 1292 417
rect 1326 416 1332 417
rect 1620 416 1622 486
rect 1696 482 1698 501
rect 1718 499 1724 500
rect 1718 495 1719 499
rect 1723 495 1724 499
rect 1718 494 1724 495
rect 1694 481 1700 482
rect 1694 477 1695 481
rect 1699 477 1700 481
rect 1720 480 1722 494
rect 1808 482 1810 501
rect 1806 481 1812 482
rect 1694 476 1700 477
rect 1718 479 1724 480
rect 1718 475 1719 479
rect 1723 475 1724 479
rect 1806 477 1807 481
rect 1811 477 1812 481
rect 1828 480 1830 510
rect 1872 507 1874 530
rect 1942 515 1948 516
rect 1942 511 1943 515
rect 1947 511 1948 515
rect 1942 510 1948 511
rect 1871 506 1875 507
rect 1871 501 1875 502
rect 1919 506 1923 507
rect 1919 501 1923 502
rect 1920 482 1922 501
rect 1918 481 1924 482
rect 1806 476 1812 477
rect 1826 479 1832 480
rect 1718 474 1724 475
rect 1826 475 1827 479
rect 1831 475 1832 479
rect 1918 477 1919 481
rect 1923 477 1924 481
rect 1944 480 1946 510
rect 1976 507 1978 530
rect 2072 507 2074 530
rect 2148 516 2150 530
rect 2146 515 2152 516
rect 2146 511 2147 515
rect 2151 511 2152 515
rect 2146 510 2152 511
rect 2168 507 2170 530
rect 2216 524 2218 582
rect 2326 568 2332 569
rect 2326 564 2327 568
rect 2331 564 2332 568
rect 2326 563 2332 564
rect 2438 568 2444 569
rect 2438 564 2439 568
rect 2443 564 2444 568
rect 2438 563 2444 564
rect 2255 562 2259 563
rect 2255 557 2259 558
rect 2327 562 2331 563
rect 2327 557 2331 558
rect 2359 562 2363 563
rect 2359 557 2363 558
rect 2439 562 2443 563
rect 2439 557 2443 558
rect 2254 556 2260 557
rect 2254 552 2255 556
rect 2259 552 2260 556
rect 2254 551 2260 552
rect 2358 556 2364 557
rect 2358 552 2359 556
rect 2363 552 2364 556
rect 2358 551 2364 552
rect 2438 556 2444 557
rect 2438 552 2439 556
rect 2443 552 2444 556
rect 2438 551 2444 552
rect 2250 535 2256 536
rect 2250 531 2251 535
rect 2255 531 2256 535
rect 2250 530 2256 531
rect 2270 535 2276 536
rect 2270 531 2271 535
rect 2275 531 2276 535
rect 2270 530 2276 531
rect 2278 535 2284 536
rect 2278 531 2279 535
rect 2283 531 2284 535
rect 2278 530 2284 531
rect 2374 535 2380 536
rect 2374 531 2375 535
rect 2379 531 2380 535
rect 2374 530 2380 531
rect 2390 535 2396 536
rect 2390 531 2391 535
rect 2395 531 2396 535
rect 2390 530 2396 531
rect 2454 535 2460 536
rect 2454 531 2455 535
rect 2459 531 2460 535
rect 2454 530 2460 531
rect 2214 523 2220 524
rect 2214 519 2215 523
rect 2219 519 2220 523
rect 2214 518 2220 519
rect 2252 516 2254 530
rect 2250 515 2256 516
rect 2250 511 2251 515
rect 2255 511 2256 515
rect 2250 510 2256 511
rect 2272 507 2274 530
rect 1975 506 1979 507
rect 1975 501 1979 502
rect 2023 506 2027 507
rect 2023 501 2027 502
rect 2071 506 2075 507
rect 2071 501 2075 502
rect 2119 506 2123 507
rect 2119 501 2123 502
rect 2167 506 2171 507
rect 2167 501 2171 502
rect 2207 506 2211 507
rect 2207 501 2211 502
rect 2271 506 2275 507
rect 2271 501 2275 502
rect 1962 499 1968 500
rect 1962 495 1963 499
rect 1967 495 1968 499
rect 1962 494 1968 495
rect 1918 476 1924 477
rect 1942 479 1948 480
rect 1826 474 1832 475
rect 1942 475 1943 479
rect 1947 475 1948 479
rect 1942 474 1948 475
rect 1678 460 1684 461
rect 1678 456 1679 460
rect 1683 456 1684 460
rect 1678 455 1684 456
rect 1790 460 1796 461
rect 1790 456 1791 460
rect 1795 456 1796 460
rect 1790 455 1796 456
rect 1902 460 1908 461
rect 1902 456 1903 460
rect 1907 456 1908 460
rect 1902 455 1908 456
rect 1680 443 1682 455
rect 1792 443 1794 455
rect 1904 443 1906 455
rect 1639 442 1643 443
rect 1639 437 1643 438
rect 1679 442 1683 443
rect 1679 437 1683 438
rect 1695 442 1699 443
rect 1695 437 1699 438
rect 1759 442 1763 443
rect 1759 437 1763 438
rect 1791 442 1795 443
rect 1791 437 1795 438
rect 1831 442 1835 443
rect 1831 437 1835 438
rect 1903 442 1907 443
rect 1903 437 1907 438
rect 1911 442 1915 443
rect 1911 437 1915 438
rect 1638 436 1644 437
rect 1638 432 1639 436
rect 1643 432 1644 436
rect 1638 431 1644 432
rect 1694 436 1700 437
rect 1694 432 1695 436
rect 1699 432 1700 436
rect 1694 431 1700 432
rect 1758 436 1764 437
rect 1758 432 1759 436
rect 1763 432 1764 436
rect 1758 431 1764 432
rect 1830 436 1836 437
rect 1830 432 1831 436
rect 1835 432 1836 436
rect 1830 431 1836 432
rect 1910 436 1916 437
rect 1910 432 1911 436
rect 1915 432 1916 436
rect 1910 431 1916 432
rect 1326 412 1327 416
rect 1331 412 1332 416
rect 1326 411 1332 412
rect 1598 415 1604 416
rect 1598 411 1599 415
rect 1603 411 1604 415
rect 1286 404 1292 405
rect 1218 403 1224 404
rect 1218 399 1219 403
rect 1223 399 1224 403
rect 1218 398 1224 399
rect 1238 403 1244 404
rect 1238 399 1239 403
rect 1243 399 1244 403
rect 1286 400 1287 404
rect 1291 400 1292 404
rect 1286 399 1292 400
rect 1238 398 1244 399
rect 1220 384 1222 398
rect 1166 383 1172 384
rect 1166 379 1167 383
rect 1171 379 1172 383
rect 1166 378 1172 379
rect 1218 383 1224 384
rect 1218 379 1219 383
rect 1223 379 1224 383
rect 1218 378 1224 379
rect 1240 375 1242 398
rect 1288 375 1290 399
rect 1328 387 1330 411
rect 1598 410 1604 411
rect 1618 415 1624 416
rect 1618 411 1619 415
rect 1623 411 1624 415
rect 1618 410 1624 411
rect 1654 415 1660 416
rect 1654 411 1655 415
rect 1659 411 1660 415
rect 1654 410 1660 411
rect 1710 415 1716 416
rect 1710 411 1711 415
rect 1715 411 1716 415
rect 1710 410 1716 411
rect 1774 415 1780 416
rect 1774 411 1775 415
rect 1779 411 1780 415
rect 1774 410 1780 411
rect 1846 415 1852 416
rect 1846 411 1847 415
rect 1851 411 1852 415
rect 1846 410 1852 411
rect 1926 415 1932 416
rect 1926 411 1927 415
rect 1931 411 1932 415
rect 1926 410 1932 411
rect 1600 387 1602 410
rect 1656 387 1658 410
rect 1712 387 1714 410
rect 1776 387 1778 410
rect 1848 387 1850 410
rect 1886 395 1892 396
rect 1886 391 1887 395
rect 1891 391 1892 395
rect 1886 390 1892 391
rect 1894 395 1900 396
rect 1894 391 1895 395
rect 1899 391 1900 395
rect 1894 390 1900 391
rect 1327 386 1331 387
rect 1327 381 1331 382
rect 1599 386 1603 387
rect 1599 381 1603 382
rect 1655 386 1659 387
rect 1655 381 1659 382
rect 1679 386 1683 387
rect 1679 381 1683 382
rect 1711 386 1715 387
rect 1711 381 1715 382
rect 1735 386 1739 387
rect 1735 381 1739 382
rect 1775 386 1779 387
rect 1775 381 1779 382
rect 1799 386 1803 387
rect 1799 381 1803 382
rect 1847 386 1851 387
rect 1847 381 1851 382
rect 1871 386 1875 387
rect 1871 381 1875 382
rect 1095 374 1099 375
rect 1095 369 1099 370
rect 1159 374 1163 375
rect 1159 369 1163 370
rect 1175 374 1179 375
rect 1175 369 1179 370
rect 1239 374 1243 375
rect 1239 369 1243 370
rect 1287 374 1291 375
rect 1287 369 1291 370
rect 1074 367 1080 368
rect 1074 363 1075 367
rect 1079 363 1080 367
rect 1074 362 1080 363
rect 1096 350 1098 369
rect 1118 367 1124 368
rect 1118 363 1119 367
rect 1123 363 1124 367
rect 1118 362 1124 363
rect 934 349 940 350
rect 846 344 852 345
rect 870 347 876 348
rect 770 342 776 343
rect 870 343 871 347
rect 875 343 876 347
rect 934 345 935 349
rect 939 345 940 349
rect 1014 349 1020 350
rect 934 344 940 345
rect 950 347 956 348
rect 870 342 876 343
rect 950 343 951 347
rect 955 343 956 347
rect 1014 345 1015 349
rect 1019 345 1020 349
rect 1014 344 1020 345
rect 1094 349 1100 350
rect 1094 345 1095 349
rect 1099 345 1100 349
rect 1120 348 1122 362
rect 1176 350 1178 369
rect 1198 367 1204 368
rect 1198 363 1199 367
rect 1203 363 1204 367
rect 1198 362 1204 363
rect 1174 349 1180 350
rect 1094 344 1100 345
rect 1118 347 1124 348
rect 950 342 956 343
rect 1118 343 1119 347
rect 1123 343 1124 347
rect 1174 345 1175 349
rect 1179 345 1180 349
rect 1200 348 1202 362
rect 1240 350 1242 369
rect 1238 349 1244 350
rect 1288 349 1290 369
rect 1328 361 1330 381
rect 1622 379 1628 380
rect 1622 375 1623 379
rect 1627 375 1628 379
rect 1622 374 1628 375
rect 1326 360 1332 361
rect 1326 356 1327 360
rect 1331 356 1332 360
rect 1326 355 1332 356
rect 1174 344 1180 345
rect 1198 347 1204 348
rect 1118 342 1124 343
rect 1198 343 1199 347
rect 1203 343 1204 347
rect 1238 345 1239 349
rect 1243 345 1244 349
rect 1286 348 1292 349
rect 1238 344 1244 345
rect 1246 347 1252 348
rect 1198 342 1204 343
rect 1246 343 1247 347
rect 1251 343 1252 347
rect 1286 344 1287 348
rect 1291 344 1292 348
rect 1286 343 1292 344
rect 1326 343 1332 344
rect 1246 342 1252 343
rect 734 328 740 329
rect 734 324 735 328
rect 739 324 740 328
rect 734 323 740 324
rect 830 328 836 329
rect 830 324 831 328
rect 835 324 836 328
rect 830 323 836 324
rect 918 328 924 329
rect 918 324 919 328
rect 923 324 924 328
rect 918 323 924 324
rect 736 319 738 323
rect 832 319 834 323
rect 920 319 922 323
rect 735 318 739 319
rect 735 313 739 314
rect 743 318 747 319
rect 743 313 747 314
rect 831 318 835 319
rect 831 313 835 314
rect 847 318 851 319
rect 847 313 851 314
rect 919 318 923 319
rect 919 313 923 314
rect 943 318 947 319
rect 943 313 947 314
rect 742 312 748 313
rect 742 308 743 312
rect 747 308 748 312
rect 742 307 748 308
rect 846 312 852 313
rect 846 308 847 312
rect 851 308 852 312
rect 846 307 852 308
rect 942 312 948 313
rect 942 308 943 312
rect 947 308 948 312
rect 942 307 948 308
rect 654 291 660 292
rect 654 287 655 291
rect 659 287 660 291
rect 654 286 660 287
rect 662 291 668 292
rect 662 287 663 291
rect 667 287 668 291
rect 662 286 668 287
rect 758 291 764 292
rect 758 287 759 291
rect 763 287 764 291
rect 758 286 764 287
rect 862 291 868 292
rect 862 287 863 291
rect 867 287 868 291
rect 862 286 868 287
rect 558 271 564 272
rect 558 267 559 271
rect 563 267 564 271
rect 656 267 658 286
rect 760 267 762 286
rect 864 267 866 286
rect 952 272 954 342
rect 998 328 1004 329
rect 998 324 999 328
rect 1003 324 1004 328
rect 998 323 1004 324
rect 1078 328 1084 329
rect 1078 324 1079 328
rect 1083 324 1084 328
rect 1078 323 1084 324
rect 1158 328 1164 329
rect 1158 324 1159 328
rect 1163 324 1164 328
rect 1158 323 1164 324
rect 1222 328 1228 329
rect 1222 324 1223 328
rect 1227 324 1228 328
rect 1222 323 1228 324
rect 1000 319 1002 323
rect 1080 319 1082 323
rect 1160 319 1162 323
rect 1224 319 1226 323
rect 999 318 1003 319
rect 999 313 1003 314
rect 1039 318 1043 319
rect 1039 313 1043 314
rect 1079 318 1083 319
rect 1079 313 1083 314
rect 1143 318 1147 319
rect 1143 313 1147 314
rect 1159 318 1163 319
rect 1159 313 1163 314
rect 1223 318 1227 319
rect 1223 313 1227 314
rect 1038 312 1044 313
rect 1038 308 1039 312
rect 1043 308 1044 312
rect 1038 307 1044 308
rect 1142 312 1148 313
rect 1142 308 1143 312
rect 1147 308 1148 312
rect 1142 307 1148 308
rect 1222 312 1228 313
rect 1222 308 1223 312
rect 1227 308 1228 312
rect 1222 307 1228 308
rect 958 291 964 292
rect 958 287 959 291
rect 963 287 964 291
rect 958 286 964 287
rect 1034 291 1040 292
rect 1034 287 1035 291
rect 1039 287 1040 291
rect 1034 286 1040 287
rect 1054 291 1060 292
rect 1054 287 1055 291
rect 1059 287 1060 291
rect 1054 286 1060 287
rect 1138 291 1144 292
rect 1138 287 1139 291
rect 1143 287 1144 291
rect 1138 286 1144 287
rect 1158 291 1164 292
rect 1158 287 1159 291
rect 1163 287 1164 291
rect 1158 286 1164 287
rect 1202 291 1208 292
rect 1202 287 1203 291
rect 1207 287 1208 291
rect 1202 286 1208 287
rect 1238 291 1244 292
rect 1238 287 1239 291
rect 1243 287 1244 291
rect 1238 286 1244 287
rect 890 271 896 272
rect 890 267 891 271
rect 895 267 896 271
rect 423 266 427 267
rect 423 261 427 262
rect 439 266 443 267
rect 439 261 443 262
rect 535 266 539 267
rect 535 261 539 262
rect 551 266 555 267
rect 558 266 564 267
rect 647 266 651 267
rect 551 261 555 262
rect 647 261 651 262
rect 655 266 659 267
rect 655 261 659 262
rect 759 266 763 267
rect 759 261 763 262
rect 863 266 867 267
rect 863 261 867 262
rect 871 266 875 267
rect 890 266 896 267
rect 950 271 956 272
rect 950 267 951 271
rect 955 267 956 271
rect 960 267 962 286
rect 1036 272 1038 286
rect 1034 271 1040 272
rect 1034 267 1035 271
rect 1039 267 1040 271
rect 1056 267 1058 286
rect 1140 272 1142 286
rect 1138 271 1144 272
rect 1138 267 1139 271
rect 1143 267 1144 271
rect 1160 267 1162 286
rect 950 266 956 267
rect 959 266 963 267
rect 871 261 875 262
rect 402 259 408 260
rect 402 255 403 259
rect 407 255 408 259
rect 402 254 408 255
rect 424 242 426 261
rect 446 259 452 260
rect 446 255 447 259
rect 451 255 452 259
rect 446 254 452 255
rect 318 241 324 242
rect 318 237 319 241
rect 323 237 324 241
rect 318 236 324 237
rect 422 241 428 242
rect 422 237 423 241
rect 427 237 428 241
rect 448 240 450 254
rect 536 242 538 261
rect 558 259 564 260
rect 558 255 559 259
rect 563 255 564 259
rect 558 254 564 255
rect 534 241 540 242
rect 422 236 428 237
rect 446 239 452 240
rect 446 235 447 239
rect 451 235 452 239
rect 534 237 535 241
rect 539 237 540 241
rect 560 240 562 254
rect 648 242 650 261
rect 734 259 740 260
rect 734 255 735 259
rect 739 255 740 259
rect 734 254 740 255
rect 646 241 652 242
rect 534 236 540 237
rect 558 239 564 240
rect 446 234 452 235
rect 558 235 559 239
rect 563 235 564 239
rect 646 237 647 241
rect 651 237 652 241
rect 646 236 652 237
rect 654 239 660 240
rect 558 234 564 235
rect 654 235 655 239
rect 659 235 660 239
rect 654 234 660 235
rect 406 220 412 221
rect 406 216 407 220
rect 411 216 412 220
rect 406 215 412 216
rect 518 220 524 221
rect 518 216 519 220
rect 523 216 524 220
rect 518 215 524 216
rect 630 220 636 221
rect 630 216 631 220
rect 635 216 636 220
rect 630 215 636 216
rect 408 211 410 215
rect 520 211 522 215
rect 632 211 634 215
rect 383 210 387 211
rect 383 205 387 206
rect 407 210 411 211
rect 407 205 411 206
rect 487 210 491 211
rect 487 205 491 206
rect 519 210 523 211
rect 519 205 523 206
rect 591 210 595 211
rect 591 205 595 206
rect 631 210 635 211
rect 631 205 635 206
rect 382 204 388 205
rect 382 200 383 204
rect 387 200 388 204
rect 382 199 388 200
rect 486 204 492 205
rect 486 200 487 204
rect 491 200 492 204
rect 486 199 492 200
rect 590 204 596 205
rect 590 200 591 204
rect 595 200 596 204
rect 590 199 596 200
rect 110 180 111 184
rect 115 180 116 184
rect 110 179 116 180
rect 198 183 204 184
rect 198 179 199 183
rect 203 179 204 183
rect 112 151 114 179
rect 198 178 204 179
rect 274 183 280 184
rect 274 179 275 183
rect 279 179 280 183
rect 274 178 280 179
rect 294 183 300 184
rect 294 179 295 183
rect 299 179 300 183
rect 294 178 300 179
rect 310 183 316 184
rect 310 179 311 183
rect 315 179 316 183
rect 310 178 316 179
rect 398 183 404 184
rect 398 179 399 183
rect 403 179 404 183
rect 398 178 404 179
rect 466 183 472 184
rect 466 179 467 183
rect 471 179 472 183
rect 466 178 472 179
rect 502 183 508 184
rect 502 179 503 183
rect 507 179 508 183
rect 502 178 508 179
rect 606 183 612 184
rect 606 179 607 183
rect 611 179 612 183
rect 606 178 612 179
rect 200 151 202 178
rect 276 164 278 178
rect 226 163 232 164
rect 226 159 227 163
rect 231 159 232 163
rect 226 158 232 159
rect 274 163 280 164
rect 274 159 275 163
rect 279 159 280 163
rect 274 158 280 159
rect 111 150 115 151
rect 111 145 115 146
rect 151 150 155 151
rect 151 145 155 146
rect 199 150 203 151
rect 199 145 203 146
rect 207 150 211 151
rect 207 145 211 146
rect 112 125 114 145
rect 152 126 154 145
rect 174 143 180 144
rect 174 139 175 143
rect 179 139 180 143
rect 174 138 180 139
rect 150 125 156 126
rect 110 124 116 125
rect 110 120 111 124
rect 115 120 116 124
rect 150 121 151 125
rect 155 121 156 125
rect 176 124 178 138
rect 208 126 210 145
rect 206 125 212 126
rect 150 120 156 121
rect 174 123 180 124
rect 110 119 116 120
rect 174 119 175 123
rect 179 119 180 123
rect 206 121 207 125
rect 211 121 212 125
rect 228 124 230 158
rect 296 151 298 178
rect 400 151 402 178
rect 263 150 267 151
rect 263 145 267 146
rect 295 150 299 151
rect 295 145 299 146
rect 319 150 323 151
rect 319 145 323 146
rect 375 150 379 151
rect 375 145 379 146
rect 399 150 403 151
rect 399 145 403 146
rect 431 150 435 151
rect 431 145 435 146
rect 264 126 266 145
rect 320 126 322 145
rect 376 126 378 145
rect 432 126 434 145
rect 468 144 470 178
rect 504 151 506 178
rect 608 151 610 178
rect 656 164 658 234
rect 695 210 699 211
rect 695 205 699 206
rect 694 204 700 205
rect 694 200 695 204
rect 699 200 700 204
rect 694 199 700 200
rect 736 184 738 254
rect 760 242 762 261
rect 782 259 788 260
rect 782 255 783 259
rect 787 255 788 259
rect 782 254 788 255
rect 758 241 764 242
rect 758 237 759 241
rect 763 237 764 241
rect 784 240 786 254
rect 872 242 874 261
rect 870 241 876 242
rect 758 236 764 237
rect 782 239 788 240
rect 782 235 783 239
rect 787 235 788 239
rect 870 237 871 241
rect 875 237 876 241
rect 892 240 894 266
rect 959 261 963 262
rect 983 266 987 267
rect 1034 266 1040 267
rect 1055 266 1059 267
rect 983 261 987 262
rect 1055 261 1059 262
rect 1103 266 1107 267
rect 1138 266 1144 267
rect 1159 266 1163 267
rect 1103 261 1107 262
rect 1159 261 1163 262
rect 984 242 986 261
rect 1104 242 1106 261
rect 1204 260 1206 286
rect 1240 267 1242 286
rect 1248 272 1250 342
rect 1326 339 1327 343
rect 1331 339 1332 343
rect 1326 338 1332 339
rect 1286 331 1292 332
rect 1286 327 1287 331
rect 1291 327 1292 331
rect 1328 327 1330 338
rect 1286 326 1292 327
rect 1327 326 1331 327
rect 1288 319 1290 326
rect 1327 321 1331 322
rect 1351 326 1355 327
rect 1351 321 1355 322
rect 1455 326 1459 327
rect 1455 321 1459 322
rect 1583 326 1587 327
rect 1583 321 1587 322
rect 1287 318 1291 319
rect 1328 318 1330 321
rect 1350 320 1356 321
rect 1287 313 1291 314
rect 1326 317 1332 318
rect 1326 313 1327 317
rect 1331 313 1332 317
rect 1350 316 1351 320
rect 1355 316 1356 320
rect 1350 315 1356 316
rect 1454 320 1460 321
rect 1454 316 1455 320
rect 1459 316 1460 320
rect 1454 315 1460 316
rect 1582 320 1588 321
rect 1582 316 1583 320
rect 1587 316 1588 320
rect 1582 315 1588 316
rect 1288 310 1290 313
rect 1326 312 1332 313
rect 1286 309 1292 310
rect 1286 305 1287 309
rect 1291 305 1292 309
rect 1286 304 1292 305
rect 1326 300 1332 301
rect 1624 300 1626 374
rect 1680 362 1682 381
rect 1702 379 1708 380
rect 1702 375 1703 379
rect 1707 375 1708 379
rect 1702 374 1708 375
rect 1678 361 1684 362
rect 1678 357 1679 361
rect 1683 357 1684 361
rect 1704 360 1706 374
rect 1736 362 1738 381
rect 1758 379 1764 380
rect 1758 375 1759 379
rect 1763 375 1764 379
rect 1758 374 1764 375
rect 1734 361 1740 362
rect 1678 356 1684 357
rect 1702 359 1708 360
rect 1702 355 1703 359
rect 1707 355 1708 359
rect 1734 357 1735 361
rect 1739 357 1740 361
rect 1760 360 1762 374
rect 1800 362 1802 381
rect 1822 379 1828 380
rect 1822 375 1823 379
rect 1827 375 1828 379
rect 1822 374 1828 375
rect 1798 361 1804 362
rect 1734 356 1740 357
rect 1758 359 1764 360
rect 1702 354 1708 355
rect 1758 355 1759 359
rect 1763 355 1764 359
rect 1798 357 1799 361
rect 1803 357 1804 361
rect 1824 360 1826 374
rect 1872 362 1874 381
rect 1878 379 1884 380
rect 1878 375 1879 379
rect 1883 375 1884 379
rect 1878 374 1884 375
rect 1870 361 1876 362
rect 1798 356 1804 357
rect 1822 359 1828 360
rect 1758 354 1764 355
rect 1822 355 1823 359
rect 1827 355 1828 359
rect 1870 357 1871 361
rect 1875 357 1876 361
rect 1870 356 1876 357
rect 1822 354 1828 355
rect 1662 340 1668 341
rect 1662 336 1663 340
rect 1667 336 1668 340
rect 1662 335 1668 336
rect 1718 340 1724 341
rect 1718 336 1719 340
rect 1723 336 1724 340
rect 1718 335 1724 336
rect 1782 340 1788 341
rect 1782 336 1783 340
rect 1787 336 1788 340
rect 1782 335 1788 336
rect 1854 340 1860 341
rect 1854 336 1855 340
rect 1859 336 1860 340
rect 1854 335 1860 336
rect 1664 327 1666 335
rect 1720 327 1722 335
rect 1784 327 1786 335
rect 1856 327 1858 335
rect 1663 326 1667 327
rect 1663 321 1667 322
rect 1711 326 1715 327
rect 1711 321 1715 322
rect 1719 326 1723 327
rect 1719 321 1723 322
rect 1783 326 1787 327
rect 1783 321 1787 322
rect 1839 326 1843 327
rect 1839 321 1843 322
rect 1855 326 1859 327
rect 1855 321 1859 322
rect 1710 320 1716 321
rect 1710 316 1711 320
rect 1715 316 1716 320
rect 1710 315 1716 316
rect 1838 320 1844 321
rect 1838 316 1839 320
rect 1843 316 1844 320
rect 1838 315 1844 316
rect 1880 300 1882 374
rect 1888 368 1890 390
rect 1886 367 1892 368
rect 1886 363 1887 367
rect 1891 363 1892 367
rect 1886 362 1892 363
rect 1896 360 1898 390
rect 1928 387 1930 410
rect 1927 386 1931 387
rect 1927 381 1931 382
rect 1943 386 1947 387
rect 1943 381 1947 382
rect 1944 362 1946 381
rect 1942 361 1948 362
rect 1894 359 1900 360
rect 1894 355 1895 359
rect 1899 355 1900 359
rect 1942 357 1943 361
rect 1947 357 1948 361
rect 1964 360 1966 494
rect 2024 482 2026 501
rect 2046 499 2052 500
rect 2046 495 2047 499
rect 2051 495 2052 499
rect 2046 494 2052 495
rect 2022 481 2028 482
rect 2022 477 2023 481
rect 2027 477 2028 481
rect 2048 480 2050 494
rect 2120 482 2122 501
rect 2208 482 2210 501
rect 2280 500 2282 530
rect 2376 507 2378 530
rect 2392 508 2394 530
rect 2414 515 2420 516
rect 2414 511 2415 515
rect 2419 511 2420 515
rect 2414 510 2420 511
rect 2390 507 2396 508
rect 2295 506 2299 507
rect 2295 501 2299 502
rect 2375 506 2379 507
rect 2375 501 2379 502
rect 2383 506 2387 507
rect 2390 503 2391 507
rect 2395 503 2396 507
rect 2390 502 2396 503
rect 2383 501 2387 502
rect 2278 499 2284 500
rect 2278 495 2279 499
rect 2283 495 2284 499
rect 2278 494 2284 495
rect 2296 482 2298 501
rect 2314 499 2320 500
rect 2314 495 2315 499
rect 2319 495 2320 499
rect 2314 494 2320 495
rect 2118 481 2124 482
rect 2022 476 2028 477
rect 2046 479 2052 480
rect 2046 475 2047 479
rect 2051 475 2052 479
rect 2118 477 2119 481
rect 2123 477 2124 481
rect 2206 481 2212 482
rect 2118 476 2124 477
rect 2166 479 2172 480
rect 2046 474 2052 475
rect 2166 475 2167 479
rect 2171 475 2172 479
rect 2206 477 2207 481
rect 2211 477 2212 481
rect 2206 476 2212 477
rect 2294 481 2300 482
rect 2294 477 2295 481
rect 2299 477 2300 481
rect 2316 480 2318 494
rect 2384 482 2386 501
rect 2416 488 2418 510
rect 2456 507 2458 530
rect 2464 516 2466 582
rect 2502 571 2508 572
rect 2502 567 2503 571
rect 2507 567 2508 571
rect 2502 566 2508 567
rect 2504 563 2506 566
rect 2503 562 2507 563
rect 2503 557 2507 558
rect 2504 554 2506 557
rect 2502 553 2508 554
rect 2502 549 2503 553
rect 2507 549 2508 553
rect 2502 548 2508 549
rect 2502 536 2508 537
rect 2470 535 2476 536
rect 2470 531 2471 535
rect 2475 531 2476 535
rect 2502 532 2503 536
rect 2507 532 2508 536
rect 2502 531 2508 532
rect 2470 530 2476 531
rect 2462 515 2468 516
rect 2462 511 2463 515
rect 2467 511 2468 515
rect 2462 510 2468 511
rect 2455 506 2459 507
rect 2455 501 2459 502
rect 2446 499 2452 500
rect 2446 495 2447 499
rect 2451 495 2452 499
rect 2446 494 2452 495
rect 2414 487 2420 488
rect 2414 483 2415 487
rect 2419 483 2420 487
rect 2414 482 2420 483
rect 2382 481 2388 482
rect 2294 476 2300 477
rect 2314 479 2320 480
rect 2166 474 2172 475
rect 2314 475 2315 479
rect 2319 475 2320 479
rect 2382 477 2383 481
rect 2387 477 2388 481
rect 2382 476 2388 477
rect 2398 479 2404 480
rect 2314 474 2320 475
rect 2398 475 2399 479
rect 2403 475 2404 479
rect 2398 474 2404 475
rect 2006 460 2012 461
rect 2006 456 2007 460
rect 2011 456 2012 460
rect 2006 455 2012 456
rect 2102 460 2108 461
rect 2102 456 2103 460
rect 2107 456 2108 460
rect 2102 455 2108 456
rect 2008 443 2010 455
rect 2104 443 2106 455
rect 1991 442 1995 443
rect 1991 437 1995 438
rect 2007 442 2011 443
rect 2007 437 2011 438
rect 2079 442 2083 443
rect 2079 437 2083 438
rect 2103 442 2107 443
rect 2103 437 2107 438
rect 1990 436 1996 437
rect 1990 432 1991 436
rect 1995 432 1996 436
rect 1990 431 1996 432
rect 2078 436 2084 437
rect 2078 432 2079 436
rect 2083 432 2084 436
rect 2078 431 2084 432
rect 1986 415 1992 416
rect 1986 411 1987 415
rect 1991 411 1992 415
rect 1986 410 1992 411
rect 2006 415 2012 416
rect 2006 411 2007 415
rect 2011 411 2012 415
rect 2006 410 2012 411
rect 2074 415 2080 416
rect 2074 411 2075 415
rect 2079 411 2080 415
rect 2074 410 2080 411
rect 2094 415 2100 416
rect 2094 411 2095 415
rect 2099 411 2100 415
rect 2094 410 2100 411
rect 2102 415 2108 416
rect 2102 411 2103 415
rect 2107 411 2108 415
rect 2102 410 2108 411
rect 1988 396 1990 410
rect 1986 395 1992 396
rect 1986 391 1987 395
rect 1991 391 1992 395
rect 1986 390 1992 391
rect 2008 387 2010 410
rect 2076 396 2078 410
rect 2074 395 2080 396
rect 2074 391 2075 395
rect 2079 391 2080 395
rect 2074 390 2080 391
rect 2096 387 2098 410
rect 2007 386 2011 387
rect 2007 381 2011 382
rect 2023 386 2027 387
rect 2023 381 2027 382
rect 2095 386 2099 387
rect 2095 381 2099 382
rect 2024 362 2026 381
rect 2104 380 2106 410
rect 2168 396 2170 474
rect 2190 460 2196 461
rect 2190 456 2191 460
rect 2195 456 2196 460
rect 2190 455 2196 456
rect 2278 460 2284 461
rect 2278 456 2279 460
rect 2283 456 2284 460
rect 2278 455 2284 456
rect 2366 460 2372 461
rect 2366 456 2367 460
rect 2371 456 2372 460
rect 2366 455 2372 456
rect 2192 443 2194 455
rect 2280 443 2282 455
rect 2368 443 2370 455
rect 2175 442 2179 443
rect 2175 437 2179 438
rect 2191 442 2195 443
rect 2191 437 2195 438
rect 2271 442 2275 443
rect 2271 437 2275 438
rect 2279 442 2283 443
rect 2279 437 2283 438
rect 2367 442 2371 443
rect 2367 437 2371 438
rect 2174 436 2180 437
rect 2174 432 2175 436
rect 2179 432 2180 436
rect 2174 431 2180 432
rect 2270 436 2276 437
rect 2270 432 2271 436
rect 2275 432 2276 436
rect 2270 431 2276 432
rect 2366 436 2372 437
rect 2366 432 2367 436
rect 2371 432 2372 436
rect 2366 431 2372 432
rect 2190 415 2196 416
rect 2190 411 2191 415
rect 2195 411 2196 415
rect 2190 410 2196 411
rect 2266 415 2272 416
rect 2266 411 2267 415
rect 2271 411 2272 415
rect 2266 410 2272 411
rect 2286 415 2292 416
rect 2286 411 2287 415
rect 2291 411 2292 415
rect 2286 410 2292 411
rect 2294 415 2300 416
rect 2294 411 2295 415
rect 2299 411 2300 415
rect 2294 410 2300 411
rect 2382 415 2388 416
rect 2382 411 2383 415
rect 2387 411 2388 415
rect 2382 410 2388 411
rect 2390 415 2396 416
rect 2390 411 2391 415
rect 2395 411 2396 415
rect 2390 410 2396 411
rect 2166 395 2172 396
rect 2166 391 2167 395
rect 2171 391 2172 395
rect 2166 390 2172 391
rect 2192 387 2194 410
rect 2268 396 2270 410
rect 2266 395 2272 396
rect 2266 391 2267 395
rect 2271 391 2272 395
rect 2266 390 2272 391
rect 2288 387 2290 410
rect 2111 386 2115 387
rect 2111 381 2115 382
rect 2191 386 2195 387
rect 2191 381 2195 382
rect 2199 386 2203 387
rect 2199 381 2203 382
rect 2287 386 2291 387
rect 2287 381 2291 382
rect 2102 379 2108 380
rect 2102 375 2103 379
rect 2107 375 2108 379
rect 2102 374 2108 375
rect 2112 362 2114 381
rect 2200 362 2202 381
rect 2288 362 2290 381
rect 2296 380 2298 410
rect 2384 387 2386 410
rect 2375 386 2379 387
rect 2375 381 2379 382
rect 2383 386 2387 387
rect 2383 381 2387 382
rect 2294 379 2300 380
rect 2294 375 2295 379
rect 2299 375 2300 379
rect 2294 374 2300 375
rect 2376 362 2378 381
rect 2392 380 2394 410
rect 2400 396 2402 474
rect 2438 460 2444 461
rect 2438 456 2439 460
rect 2443 456 2444 460
rect 2438 455 2444 456
rect 2440 443 2442 455
rect 2439 442 2443 443
rect 2439 437 2443 438
rect 2438 436 2444 437
rect 2438 432 2439 436
rect 2443 432 2444 436
rect 2438 431 2444 432
rect 2398 395 2404 396
rect 2398 391 2399 395
rect 2403 391 2404 395
rect 2398 390 2404 391
rect 2390 379 2396 380
rect 2390 375 2391 379
rect 2395 375 2396 379
rect 2390 374 2396 375
rect 2448 368 2450 494
rect 2456 482 2458 501
rect 2454 481 2460 482
rect 2454 477 2455 481
rect 2459 477 2460 481
rect 2454 476 2460 477
rect 2454 415 2460 416
rect 2454 411 2455 415
rect 2459 411 2460 415
rect 2454 410 2460 411
rect 2462 415 2468 416
rect 2462 411 2463 415
rect 2467 411 2468 415
rect 2462 410 2468 411
rect 2456 387 2458 410
rect 2455 386 2459 387
rect 2455 381 2459 382
rect 2446 367 2452 368
rect 2446 363 2447 367
rect 2451 363 2452 367
rect 2446 362 2452 363
rect 2456 362 2458 381
rect 2022 361 2028 362
rect 1942 356 1948 357
rect 1962 359 1968 360
rect 1894 354 1900 355
rect 1962 355 1963 359
rect 1967 355 1968 359
rect 2022 357 2023 361
rect 2027 357 2028 361
rect 2022 356 2028 357
rect 2110 361 2116 362
rect 2110 357 2111 361
rect 2115 357 2116 361
rect 2110 356 2116 357
rect 2198 361 2204 362
rect 2198 357 2199 361
rect 2203 357 2204 361
rect 2286 361 2292 362
rect 2198 356 2204 357
rect 2206 359 2212 360
rect 1962 354 1968 355
rect 2206 355 2207 359
rect 2211 355 2212 359
rect 2286 357 2287 361
rect 2291 357 2292 361
rect 2286 356 2292 357
rect 2374 361 2380 362
rect 2374 357 2375 361
rect 2379 357 2380 361
rect 2454 361 2460 362
rect 2374 356 2380 357
rect 2382 359 2388 360
rect 2206 354 2212 355
rect 2382 355 2383 359
rect 2387 355 2388 359
rect 2454 357 2455 361
rect 2459 357 2460 361
rect 2454 356 2460 357
rect 2382 354 2388 355
rect 1926 340 1932 341
rect 1926 336 1927 340
rect 1931 336 1932 340
rect 1926 335 1932 336
rect 2006 340 2012 341
rect 2006 336 2007 340
rect 2011 336 2012 340
rect 2006 335 2012 336
rect 2094 340 2100 341
rect 2094 336 2095 340
rect 2099 336 2100 340
rect 2094 335 2100 336
rect 2182 340 2188 341
rect 2182 336 2183 340
rect 2187 336 2188 340
rect 2182 335 2188 336
rect 1928 327 1930 335
rect 2008 327 2010 335
rect 2096 327 2098 335
rect 2184 327 2186 335
rect 1927 326 1931 327
rect 1927 321 1931 322
rect 1951 326 1955 327
rect 1951 321 1955 322
rect 2007 326 2011 327
rect 2007 321 2011 322
rect 2063 326 2067 327
rect 2063 321 2067 322
rect 2095 326 2099 327
rect 2095 321 2099 322
rect 2167 326 2171 327
rect 2167 321 2171 322
rect 2183 326 2187 327
rect 2183 321 2187 322
rect 1950 320 1956 321
rect 1950 316 1951 320
rect 1955 316 1956 320
rect 1950 315 1956 316
rect 2062 320 2068 321
rect 2062 316 2063 320
rect 2067 316 2068 320
rect 2062 315 2068 316
rect 2166 320 2172 321
rect 2166 316 2167 320
rect 2171 316 2172 320
rect 2166 315 2172 316
rect 1326 296 1327 300
rect 1331 296 1332 300
rect 1326 295 1332 296
rect 1366 299 1372 300
rect 1366 295 1367 299
rect 1371 295 1372 299
rect 1286 292 1292 293
rect 1286 288 1287 292
rect 1291 288 1292 292
rect 1286 287 1292 288
rect 1246 271 1252 272
rect 1246 267 1247 271
rect 1251 267 1252 271
rect 1288 267 1290 287
rect 1328 267 1330 295
rect 1366 294 1372 295
rect 1374 299 1380 300
rect 1374 295 1375 299
rect 1379 295 1380 299
rect 1374 294 1380 295
rect 1470 299 1476 300
rect 1470 295 1471 299
rect 1475 295 1476 299
rect 1470 294 1476 295
rect 1578 299 1584 300
rect 1578 295 1579 299
rect 1583 295 1584 299
rect 1578 294 1584 295
rect 1598 299 1604 300
rect 1598 295 1599 299
rect 1603 295 1604 299
rect 1598 294 1604 295
rect 1622 299 1628 300
rect 1622 295 1623 299
rect 1627 295 1628 299
rect 1622 294 1628 295
rect 1726 299 1732 300
rect 1726 295 1727 299
rect 1731 295 1732 299
rect 1726 294 1732 295
rect 1854 299 1860 300
rect 1854 295 1855 299
rect 1859 295 1860 299
rect 1854 294 1860 295
rect 1878 299 1884 300
rect 1878 295 1879 299
rect 1883 295 1884 299
rect 1878 294 1884 295
rect 1966 299 1972 300
rect 1966 295 1967 299
rect 1971 295 1972 299
rect 1966 294 1972 295
rect 2078 299 2084 300
rect 2078 295 2079 299
rect 2083 295 2084 299
rect 2078 294 2084 295
rect 2086 299 2092 300
rect 2086 295 2087 299
rect 2091 295 2092 299
rect 2086 294 2092 295
rect 2182 299 2188 300
rect 2182 295 2183 299
rect 2187 295 2188 299
rect 2182 294 2188 295
rect 1368 267 1370 294
rect 1223 266 1227 267
rect 1223 261 1227 262
rect 1239 266 1243 267
rect 1246 266 1252 267
rect 1287 266 1291 267
rect 1239 261 1243 262
rect 1287 261 1291 262
rect 1327 266 1331 267
rect 1327 261 1331 262
rect 1367 266 1371 267
rect 1367 261 1371 262
rect 1202 259 1208 260
rect 1202 255 1203 259
rect 1207 255 1208 259
rect 1202 254 1208 255
rect 1224 242 1226 261
rect 982 241 988 242
rect 870 236 876 237
rect 890 239 896 240
rect 782 234 788 235
rect 890 235 891 239
rect 895 235 896 239
rect 982 237 983 241
rect 987 237 988 241
rect 1102 241 1108 242
rect 982 236 988 237
rect 990 239 996 240
rect 890 234 896 235
rect 990 235 991 239
rect 995 235 996 239
rect 1102 237 1103 241
rect 1107 237 1108 241
rect 1102 236 1108 237
rect 1222 241 1228 242
rect 1288 241 1290 261
rect 1328 241 1330 261
rect 1368 242 1370 261
rect 1376 260 1378 294
rect 1472 267 1474 294
rect 1580 280 1582 294
rect 1578 279 1584 280
rect 1578 275 1579 279
rect 1583 275 1584 279
rect 1578 274 1584 275
rect 1600 267 1602 294
rect 1728 267 1730 294
rect 1778 279 1784 280
rect 1778 275 1779 279
rect 1783 275 1784 279
rect 1778 274 1784 275
rect 1447 266 1451 267
rect 1447 261 1451 262
rect 1471 266 1475 267
rect 1471 261 1475 262
rect 1551 266 1555 267
rect 1551 261 1555 262
rect 1599 266 1603 267
rect 1599 261 1603 262
rect 1655 266 1659 267
rect 1655 261 1659 262
rect 1727 266 1731 267
rect 1727 261 1731 262
rect 1759 266 1763 267
rect 1759 261 1763 262
rect 1374 259 1380 260
rect 1374 255 1375 259
rect 1379 255 1380 259
rect 1374 254 1380 255
rect 1390 259 1396 260
rect 1390 255 1391 259
rect 1395 255 1396 259
rect 1390 254 1396 255
rect 1366 241 1372 242
rect 1222 237 1223 241
rect 1227 237 1228 241
rect 1222 236 1228 237
rect 1286 240 1292 241
rect 1286 236 1287 240
rect 1291 236 1292 240
rect 1286 235 1292 236
rect 1326 240 1332 241
rect 1326 236 1327 240
rect 1331 236 1332 240
rect 1366 237 1367 241
rect 1371 237 1372 241
rect 1392 240 1394 254
rect 1448 242 1450 261
rect 1552 242 1554 261
rect 1574 259 1580 260
rect 1574 255 1575 259
rect 1579 255 1580 259
rect 1574 254 1580 255
rect 1446 241 1452 242
rect 1366 236 1372 237
rect 1390 239 1396 240
rect 1326 235 1332 236
rect 1390 235 1391 239
rect 1395 235 1396 239
rect 1446 237 1447 241
rect 1451 237 1452 241
rect 1550 241 1556 242
rect 1446 236 1452 237
rect 1462 239 1468 240
rect 990 234 996 235
rect 1390 234 1396 235
rect 1462 235 1463 239
rect 1467 235 1468 239
rect 1550 237 1551 241
rect 1555 237 1556 241
rect 1576 240 1578 254
rect 1586 251 1592 252
rect 1586 247 1587 251
rect 1591 247 1592 251
rect 1586 246 1592 247
rect 1550 236 1556 237
rect 1574 239 1580 240
rect 1462 234 1468 235
rect 1574 235 1575 239
rect 1579 235 1580 239
rect 1574 234 1580 235
rect 742 220 748 221
rect 742 216 743 220
rect 747 216 748 220
rect 742 215 748 216
rect 854 220 860 221
rect 854 216 855 220
rect 859 216 860 220
rect 854 215 860 216
rect 966 220 972 221
rect 966 216 967 220
rect 971 216 972 220
rect 966 215 972 216
rect 744 211 746 215
rect 856 211 858 215
rect 968 211 970 215
rect 743 210 747 211
rect 743 205 747 206
rect 799 210 803 211
rect 799 205 803 206
rect 855 210 859 211
rect 855 205 859 206
rect 895 210 899 211
rect 895 205 899 206
rect 967 210 971 211
rect 967 205 971 206
rect 798 204 804 205
rect 798 200 799 204
rect 803 200 804 204
rect 798 199 804 200
rect 894 204 900 205
rect 894 200 895 204
rect 899 200 900 204
rect 894 199 900 200
rect 992 195 994 234
rect 1286 223 1292 224
rect 1086 220 1092 221
rect 1086 216 1087 220
rect 1091 216 1092 220
rect 1086 215 1092 216
rect 1206 220 1212 221
rect 1206 216 1207 220
rect 1211 216 1212 220
rect 1286 219 1287 223
rect 1291 219 1292 223
rect 1286 218 1292 219
rect 1326 223 1332 224
rect 1326 219 1327 223
rect 1331 219 1332 223
rect 1326 218 1332 219
rect 1350 220 1356 221
rect 1206 215 1212 216
rect 1088 211 1090 215
rect 1208 211 1210 215
rect 1288 211 1290 218
rect 1328 211 1330 218
rect 1350 216 1351 220
rect 1355 216 1356 220
rect 1350 215 1356 216
rect 1430 220 1436 221
rect 1430 216 1431 220
rect 1435 216 1436 220
rect 1430 215 1436 216
rect 1352 211 1354 215
rect 1432 211 1434 215
rect 999 210 1003 211
rect 999 205 1003 206
rect 1087 210 1091 211
rect 1087 205 1091 206
rect 1103 210 1107 211
rect 1103 205 1107 206
rect 1207 210 1211 211
rect 1207 205 1211 206
rect 1287 210 1291 211
rect 1287 205 1291 206
rect 1327 210 1331 211
rect 1327 205 1331 206
rect 1351 210 1355 211
rect 1351 205 1355 206
rect 1407 210 1411 211
rect 1407 205 1411 206
rect 1431 210 1435 211
rect 1431 205 1435 206
rect 998 204 1004 205
rect 998 200 999 204
rect 1003 200 1004 204
rect 998 199 1004 200
rect 1102 204 1108 205
rect 1102 200 1103 204
rect 1107 200 1108 204
rect 1288 202 1290 205
rect 1328 202 1330 205
rect 1350 204 1356 205
rect 1102 199 1108 200
rect 1286 201 1292 202
rect 1286 197 1287 201
rect 1291 197 1292 201
rect 1286 196 1292 197
rect 1326 201 1332 202
rect 1326 197 1327 201
rect 1331 197 1332 201
rect 1350 200 1351 204
rect 1355 200 1356 204
rect 1350 199 1356 200
rect 1406 204 1412 205
rect 1406 200 1407 204
rect 1411 200 1412 204
rect 1406 199 1412 200
rect 1326 196 1332 197
rect 988 193 994 195
rect 710 183 716 184
rect 710 179 711 183
rect 715 179 716 183
rect 710 178 716 179
rect 734 183 740 184
rect 734 179 735 183
rect 739 179 740 183
rect 734 178 740 179
rect 814 183 820 184
rect 814 179 815 183
rect 819 179 820 183
rect 814 178 820 179
rect 910 183 916 184
rect 910 179 911 183
rect 915 179 916 183
rect 910 178 916 179
rect 654 163 660 164
rect 654 159 655 163
rect 659 159 660 163
rect 654 158 660 159
rect 712 151 714 178
rect 790 163 796 164
rect 790 159 791 163
rect 795 159 796 163
rect 790 158 796 159
rect 487 150 491 151
rect 487 145 491 146
rect 503 150 507 151
rect 503 145 507 146
rect 543 150 547 151
rect 543 145 547 146
rect 599 150 603 151
rect 599 145 603 146
rect 607 150 611 151
rect 607 145 611 146
rect 655 150 659 151
rect 655 145 659 146
rect 711 150 715 151
rect 711 145 715 146
rect 767 150 771 151
rect 767 145 771 146
rect 466 143 472 144
rect 466 139 467 143
rect 471 139 472 143
rect 466 138 472 139
rect 488 126 490 145
rect 510 143 516 144
rect 510 139 511 143
rect 515 139 516 143
rect 510 138 516 139
rect 262 125 268 126
rect 206 120 212 121
rect 226 123 232 124
rect 174 118 180 119
rect 226 119 227 123
rect 231 119 232 123
rect 262 121 263 125
rect 267 121 268 125
rect 262 120 268 121
rect 318 125 324 126
rect 318 121 319 125
rect 323 121 324 125
rect 318 120 324 121
rect 374 125 380 126
rect 374 121 375 125
rect 379 121 380 125
rect 374 120 380 121
rect 430 125 436 126
rect 430 121 431 125
rect 435 121 436 125
rect 430 120 436 121
rect 486 125 492 126
rect 486 121 487 125
rect 491 121 492 125
rect 512 124 514 138
rect 544 126 546 145
rect 566 143 572 144
rect 566 139 567 143
rect 571 139 572 143
rect 566 138 572 139
rect 542 125 548 126
rect 486 120 492 121
rect 510 123 516 124
rect 226 118 232 119
rect 510 119 511 123
rect 515 119 516 123
rect 542 121 543 125
rect 547 121 548 125
rect 568 124 570 138
rect 600 126 602 145
rect 656 126 658 145
rect 678 143 684 144
rect 678 139 679 143
rect 683 139 684 143
rect 678 138 684 139
rect 598 125 604 126
rect 542 120 548 121
rect 566 123 572 124
rect 510 118 516 119
rect 566 119 567 123
rect 571 119 572 123
rect 598 121 599 125
rect 603 121 604 125
rect 598 120 604 121
rect 654 125 660 126
rect 654 121 655 125
rect 659 121 660 125
rect 680 124 682 138
rect 712 126 714 145
rect 734 143 740 144
rect 734 139 735 143
rect 739 139 740 143
rect 734 138 740 139
rect 710 125 716 126
rect 654 120 660 121
rect 678 123 684 124
rect 566 118 572 119
rect 678 119 679 123
rect 683 119 684 123
rect 710 121 711 125
rect 715 121 716 125
rect 736 124 738 138
rect 768 126 770 145
rect 766 125 772 126
rect 710 120 716 121
rect 734 123 740 124
rect 678 118 684 119
rect 734 119 735 123
rect 739 119 740 123
rect 766 121 767 125
rect 771 121 772 125
rect 792 124 794 158
rect 816 151 818 178
rect 912 151 914 178
rect 988 164 990 193
rect 1286 184 1292 185
rect 994 183 1000 184
rect 994 179 995 183
rect 999 179 1000 183
rect 994 178 1000 179
rect 1014 183 1020 184
rect 1014 179 1015 183
rect 1019 179 1020 183
rect 1014 178 1020 179
rect 1098 183 1104 184
rect 1098 179 1099 183
rect 1103 179 1104 183
rect 1098 178 1104 179
rect 1118 183 1124 184
rect 1118 179 1119 183
rect 1123 179 1124 183
rect 1118 178 1124 179
rect 1134 183 1140 184
rect 1134 179 1135 183
rect 1139 179 1140 183
rect 1286 180 1287 184
rect 1291 180 1292 184
rect 1286 179 1292 180
rect 1326 184 1332 185
rect 1326 180 1327 184
rect 1331 180 1332 184
rect 1326 179 1332 180
rect 1366 183 1372 184
rect 1366 179 1367 183
rect 1371 179 1372 183
rect 1134 178 1140 179
rect 996 164 998 178
rect 986 163 992 164
rect 986 159 987 163
rect 991 159 992 163
rect 986 158 992 159
rect 994 163 1000 164
rect 994 159 995 163
rect 999 159 1000 163
rect 994 158 1000 159
rect 1016 151 1018 178
rect 1100 164 1102 178
rect 1098 163 1104 164
rect 1098 159 1099 163
rect 1103 159 1104 163
rect 1098 158 1104 159
rect 1120 151 1122 178
rect 815 150 819 151
rect 815 145 819 146
rect 831 150 835 151
rect 831 145 835 146
rect 895 150 899 151
rect 895 145 899 146
rect 911 150 915 151
rect 911 145 915 146
rect 959 150 963 151
rect 959 145 963 146
rect 1015 150 1019 151
rect 1015 145 1019 146
rect 1023 150 1027 151
rect 1023 145 1027 146
rect 1087 150 1091 151
rect 1087 145 1091 146
rect 1119 150 1123 151
rect 1119 145 1123 146
rect 832 126 834 145
rect 896 126 898 145
rect 960 126 962 145
rect 1024 126 1026 145
rect 1088 126 1090 145
rect 1136 144 1138 178
rect 1288 151 1290 179
rect 1151 150 1155 151
rect 1151 145 1155 146
rect 1287 150 1291 151
rect 1287 145 1291 146
rect 1134 143 1140 144
rect 1134 139 1135 143
rect 1139 139 1140 143
rect 1134 138 1140 139
rect 1152 126 1154 145
rect 830 125 836 126
rect 766 120 772 121
rect 790 123 796 124
rect 734 118 740 119
rect 790 119 791 123
rect 795 119 796 123
rect 830 121 831 125
rect 835 121 836 125
rect 830 120 836 121
rect 894 125 900 126
rect 894 121 895 125
rect 899 121 900 125
rect 894 120 900 121
rect 958 125 964 126
rect 958 121 959 125
rect 963 121 964 125
rect 958 120 964 121
rect 1022 125 1028 126
rect 1022 121 1023 125
rect 1027 121 1028 125
rect 1022 120 1028 121
rect 1086 125 1092 126
rect 1086 121 1087 125
rect 1091 121 1092 125
rect 1086 120 1092 121
rect 1150 125 1156 126
rect 1288 125 1290 145
rect 1328 139 1330 179
rect 1366 178 1372 179
rect 1374 183 1380 184
rect 1374 179 1375 183
rect 1379 179 1380 183
rect 1374 178 1380 179
rect 1422 183 1428 184
rect 1422 179 1423 183
rect 1427 179 1428 183
rect 1422 178 1428 179
rect 1368 139 1370 178
rect 1327 138 1331 139
rect 1327 133 1331 134
rect 1367 138 1371 139
rect 1367 133 1371 134
rect 1150 121 1151 125
rect 1155 121 1156 125
rect 1150 120 1156 121
rect 1286 124 1292 125
rect 1286 120 1287 124
rect 1291 120 1292 124
rect 1286 119 1292 120
rect 790 118 796 119
rect 1328 113 1330 133
rect 1368 114 1370 133
rect 1376 132 1378 178
rect 1424 139 1426 178
rect 1464 164 1466 234
rect 1534 220 1540 221
rect 1534 216 1535 220
rect 1539 216 1540 220
rect 1534 215 1540 216
rect 1536 211 1538 215
rect 1471 210 1475 211
rect 1471 205 1475 206
rect 1535 210 1539 211
rect 1535 205 1539 206
rect 1551 210 1555 211
rect 1551 205 1555 206
rect 1470 204 1476 205
rect 1470 200 1471 204
rect 1475 200 1476 204
rect 1470 199 1476 200
rect 1550 204 1556 205
rect 1550 200 1551 204
rect 1555 200 1556 204
rect 1550 199 1556 200
rect 1588 184 1590 246
rect 1656 242 1658 261
rect 1678 259 1684 260
rect 1678 255 1679 259
rect 1683 255 1684 259
rect 1678 254 1684 255
rect 1654 241 1660 242
rect 1654 237 1655 241
rect 1659 237 1660 241
rect 1680 240 1682 254
rect 1760 242 1762 261
rect 1758 241 1764 242
rect 1654 236 1660 237
rect 1678 239 1684 240
rect 1678 235 1679 239
rect 1683 235 1684 239
rect 1758 237 1759 241
rect 1763 237 1764 241
rect 1780 240 1782 274
rect 1856 267 1858 294
rect 1968 267 1970 294
rect 1986 279 1992 280
rect 1986 275 1987 279
rect 1991 275 1992 279
rect 1986 274 1992 275
rect 1855 266 1859 267
rect 1855 261 1859 262
rect 1863 266 1867 267
rect 1863 261 1867 262
rect 1967 266 1971 267
rect 1967 261 1971 262
rect 1838 259 1844 260
rect 1838 255 1839 259
rect 1843 255 1844 259
rect 1838 254 1844 255
rect 1758 236 1764 237
rect 1778 239 1784 240
rect 1678 234 1684 235
rect 1778 235 1779 239
rect 1783 235 1784 239
rect 1778 234 1784 235
rect 1638 220 1644 221
rect 1638 216 1639 220
rect 1643 216 1644 220
rect 1638 215 1644 216
rect 1742 220 1748 221
rect 1742 216 1743 220
rect 1747 216 1748 220
rect 1742 215 1748 216
rect 1640 211 1642 215
rect 1744 211 1746 215
rect 1639 210 1643 211
rect 1639 205 1643 206
rect 1719 210 1723 211
rect 1719 205 1723 206
rect 1743 210 1747 211
rect 1743 205 1747 206
rect 1807 210 1811 211
rect 1807 205 1811 206
rect 1638 204 1644 205
rect 1638 200 1639 204
rect 1643 200 1644 204
rect 1638 199 1644 200
rect 1718 204 1724 205
rect 1718 200 1719 204
rect 1723 200 1724 204
rect 1718 199 1724 200
rect 1806 204 1812 205
rect 1806 200 1807 204
rect 1811 200 1812 204
rect 1806 199 1812 200
rect 1840 184 1842 254
rect 1864 242 1866 261
rect 1886 259 1892 260
rect 1886 255 1887 259
rect 1891 255 1892 259
rect 1886 254 1892 255
rect 1862 241 1868 242
rect 1862 237 1863 241
rect 1867 237 1868 241
rect 1888 240 1890 254
rect 1968 242 1970 261
rect 1966 241 1972 242
rect 1862 236 1868 237
rect 1886 239 1892 240
rect 1886 235 1887 239
rect 1891 235 1892 239
rect 1966 237 1967 241
rect 1971 237 1972 241
rect 1988 240 1990 274
rect 2080 267 2082 294
rect 2071 266 2075 267
rect 2071 261 2075 262
rect 2079 266 2083 267
rect 2079 261 2083 262
rect 2072 242 2074 261
rect 2088 260 2090 294
rect 2184 267 2186 294
rect 2208 280 2210 354
rect 2270 340 2276 341
rect 2270 336 2271 340
rect 2275 336 2276 340
rect 2270 335 2276 336
rect 2358 340 2364 341
rect 2358 336 2359 340
rect 2363 336 2364 340
rect 2358 335 2364 336
rect 2272 327 2274 335
rect 2360 327 2362 335
rect 2263 326 2267 327
rect 2263 321 2267 322
rect 2271 326 2275 327
rect 2271 321 2275 322
rect 2359 326 2363 327
rect 2359 321 2363 322
rect 2262 320 2268 321
rect 2262 316 2263 320
rect 2267 316 2268 320
rect 2262 315 2268 316
rect 2358 320 2364 321
rect 2358 316 2359 320
rect 2363 316 2364 320
rect 2358 315 2364 316
rect 2278 299 2284 300
rect 2278 295 2279 299
rect 2283 295 2284 299
rect 2278 294 2284 295
rect 2354 299 2360 300
rect 2354 295 2355 299
rect 2359 295 2360 299
rect 2354 294 2360 295
rect 2374 299 2380 300
rect 2374 295 2375 299
rect 2379 295 2380 299
rect 2374 294 2380 295
rect 2206 279 2212 280
rect 2206 275 2207 279
rect 2211 275 2212 279
rect 2206 274 2212 275
rect 2280 267 2282 294
rect 2175 266 2179 267
rect 2175 261 2179 262
rect 2183 266 2187 267
rect 2183 261 2187 262
rect 2271 266 2275 267
rect 2271 261 2275 262
rect 2279 266 2283 267
rect 2279 261 2283 262
rect 2086 259 2092 260
rect 2086 255 2087 259
rect 2091 255 2092 259
rect 2086 254 2092 255
rect 2094 259 2100 260
rect 2094 255 2095 259
rect 2099 255 2100 259
rect 2094 254 2100 255
rect 2070 241 2076 242
rect 1966 236 1972 237
rect 1986 239 1992 240
rect 1886 234 1892 235
rect 1986 235 1987 239
rect 1991 235 1992 239
rect 2070 237 2071 241
rect 2075 237 2076 241
rect 2096 240 2098 254
rect 2176 242 2178 261
rect 2198 259 2204 260
rect 2198 255 2199 259
rect 2203 255 2204 259
rect 2198 254 2204 255
rect 2174 241 2180 242
rect 2070 236 2076 237
rect 2094 239 2100 240
rect 1986 234 1992 235
rect 2094 235 2095 239
rect 2099 235 2100 239
rect 2174 237 2175 241
rect 2179 237 2180 241
rect 2200 240 2202 254
rect 2272 242 2274 261
rect 2356 260 2358 294
rect 2376 267 2378 294
rect 2384 280 2386 354
rect 2438 340 2444 341
rect 2438 336 2439 340
rect 2443 336 2444 340
rect 2438 335 2444 336
rect 2440 327 2442 335
rect 2439 326 2443 327
rect 2439 321 2443 322
rect 2438 320 2444 321
rect 2438 316 2439 320
rect 2443 316 2444 320
rect 2438 315 2444 316
rect 2454 299 2460 300
rect 2454 295 2455 299
rect 2459 295 2460 299
rect 2454 294 2460 295
rect 2382 279 2388 280
rect 2382 275 2383 279
rect 2387 275 2388 279
rect 2382 274 2388 275
rect 2456 267 2458 294
rect 2464 280 2466 410
rect 2472 396 2474 530
rect 2504 507 2506 531
rect 2503 506 2507 507
rect 2503 501 2507 502
rect 2504 481 2506 501
rect 2502 480 2508 481
rect 2502 476 2503 480
rect 2507 476 2508 480
rect 2502 475 2508 476
rect 2502 463 2508 464
rect 2502 459 2503 463
rect 2507 459 2508 463
rect 2502 458 2508 459
rect 2504 443 2506 458
rect 2503 442 2507 443
rect 2503 437 2507 438
rect 2504 434 2506 437
rect 2502 433 2508 434
rect 2502 429 2503 433
rect 2507 429 2508 433
rect 2502 428 2508 429
rect 2502 416 2508 417
rect 2502 412 2503 416
rect 2507 412 2508 416
rect 2502 411 2508 412
rect 2470 395 2476 396
rect 2470 391 2471 395
rect 2475 391 2476 395
rect 2470 390 2476 391
rect 2504 387 2506 411
rect 2503 386 2507 387
rect 2503 381 2507 382
rect 2474 379 2480 380
rect 2474 375 2475 379
rect 2479 375 2480 379
rect 2474 374 2480 375
rect 2476 300 2478 374
rect 2504 361 2506 381
rect 2502 360 2508 361
rect 2502 356 2503 360
rect 2507 356 2508 360
rect 2502 355 2508 356
rect 2502 343 2508 344
rect 2502 339 2503 343
rect 2507 339 2508 343
rect 2502 338 2508 339
rect 2504 327 2506 338
rect 2503 326 2507 327
rect 2503 321 2507 322
rect 2504 318 2506 321
rect 2502 317 2508 318
rect 2502 313 2503 317
rect 2507 313 2508 317
rect 2502 312 2508 313
rect 2502 300 2508 301
rect 2474 299 2480 300
rect 2474 295 2475 299
rect 2479 295 2480 299
rect 2502 296 2503 300
rect 2507 296 2508 300
rect 2502 295 2508 296
rect 2474 294 2480 295
rect 2462 279 2468 280
rect 2462 275 2463 279
rect 2467 275 2468 279
rect 2462 274 2468 275
rect 2504 267 2506 295
rect 2375 266 2379 267
rect 2375 261 2379 262
rect 2455 266 2459 267
rect 2455 261 2459 262
rect 2503 266 2507 267
rect 2503 261 2507 262
rect 2354 259 2360 260
rect 2354 255 2355 259
rect 2359 255 2360 259
rect 2354 254 2360 255
rect 2376 242 2378 261
rect 2398 259 2404 260
rect 2398 255 2399 259
rect 2403 255 2404 259
rect 2398 254 2404 255
rect 2270 241 2276 242
rect 2174 236 2180 237
rect 2198 239 2204 240
rect 2094 234 2100 235
rect 2198 235 2199 239
rect 2203 235 2204 239
rect 2270 237 2271 241
rect 2275 237 2276 241
rect 2374 241 2380 242
rect 2270 236 2276 237
rect 2326 239 2332 240
rect 2198 234 2204 235
rect 2326 235 2327 239
rect 2331 235 2332 239
rect 2374 237 2375 241
rect 2379 237 2380 241
rect 2400 240 2402 254
rect 2456 242 2458 261
rect 2454 241 2460 242
rect 2504 241 2506 261
rect 2374 236 2380 237
rect 2398 239 2404 240
rect 2326 234 2332 235
rect 2398 235 2399 239
rect 2403 235 2404 239
rect 2454 237 2455 241
rect 2459 237 2460 241
rect 2502 240 2508 241
rect 2454 236 2460 237
rect 2470 239 2476 240
rect 2398 234 2404 235
rect 2470 235 2471 239
rect 2475 235 2476 239
rect 2502 236 2503 240
rect 2507 236 2508 240
rect 2502 235 2508 236
rect 2470 234 2476 235
rect 1846 220 1852 221
rect 1846 216 1847 220
rect 1851 216 1852 220
rect 1846 215 1852 216
rect 1950 220 1956 221
rect 1950 216 1951 220
rect 1955 216 1956 220
rect 1950 215 1956 216
rect 2054 220 2060 221
rect 2054 216 2055 220
rect 2059 216 2060 220
rect 2054 215 2060 216
rect 2158 220 2164 221
rect 2158 216 2159 220
rect 2163 216 2164 220
rect 2158 215 2164 216
rect 2254 220 2260 221
rect 2254 216 2255 220
rect 2259 216 2260 220
rect 2254 215 2260 216
rect 1848 211 1850 215
rect 1952 211 1954 215
rect 2056 211 2058 215
rect 2160 211 2162 215
rect 2256 211 2258 215
rect 1847 210 1851 211
rect 1847 205 1851 206
rect 1895 210 1899 211
rect 1895 205 1899 206
rect 1951 210 1955 211
rect 1951 205 1955 206
rect 1991 210 1995 211
rect 1991 205 1995 206
rect 2055 210 2059 211
rect 2055 205 2059 206
rect 2103 210 2107 211
rect 2103 205 2107 206
rect 2159 210 2163 211
rect 2159 205 2163 206
rect 2215 210 2219 211
rect 2215 205 2219 206
rect 2255 210 2259 211
rect 2255 205 2259 206
rect 1894 204 1900 205
rect 1894 200 1895 204
rect 1899 200 1900 204
rect 1894 199 1900 200
rect 1990 204 1996 205
rect 1990 200 1991 204
rect 1995 200 1996 204
rect 1990 199 1996 200
rect 2102 204 2108 205
rect 2102 200 2103 204
rect 2107 200 2108 204
rect 2102 199 2108 200
rect 2214 204 2220 205
rect 2214 200 2215 204
rect 2219 200 2220 204
rect 2214 199 2220 200
rect 1486 183 1492 184
rect 1486 179 1487 183
rect 1491 179 1492 183
rect 1486 178 1492 179
rect 1566 183 1572 184
rect 1566 179 1567 183
rect 1571 179 1572 183
rect 1566 178 1572 179
rect 1586 183 1592 184
rect 1586 179 1587 183
rect 1591 179 1592 183
rect 1586 178 1592 179
rect 1654 183 1660 184
rect 1654 179 1655 183
rect 1659 179 1660 183
rect 1654 178 1660 179
rect 1734 183 1740 184
rect 1734 179 1735 183
rect 1739 179 1740 183
rect 1734 178 1740 179
rect 1822 183 1828 184
rect 1822 179 1823 183
rect 1827 179 1828 183
rect 1822 178 1828 179
rect 1838 183 1844 184
rect 1838 179 1839 183
rect 1843 179 1844 183
rect 1838 178 1844 179
rect 1910 183 1916 184
rect 1910 179 1911 183
rect 1915 179 1916 183
rect 1910 178 1916 179
rect 2006 183 2012 184
rect 2006 179 2007 183
rect 2011 179 2012 183
rect 2006 178 2012 179
rect 2118 183 2124 184
rect 2118 179 2119 183
rect 2123 179 2124 183
rect 2118 178 2124 179
rect 2126 183 2132 184
rect 2126 179 2127 183
rect 2131 179 2132 183
rect 2126 178 2132 179
rect 2230 183 2236 184
rect 2230 179 2231 183
rect 2235 179 2236 183
rect 2230 178 2236 179
rect 1462 163 1468 164
rect 1462 159 1463 163
rect 1467 159 1468 163
rect 1462 158 1468 159
rect 1488 139 1490 178
rect 1568 139 1570 178
rect 1656 139 1658 178
rect 1736 139 1738 178
rect 1778 163 1784 164
rect 1778 159 1779 163
rect 1783 159 1784 163
rect 1778 158 1784 159
rect 1423 138 1427 139
rect 1423 133 1427 134
rect 1479 138 1483 139
rect 1479 133 1483 134
rect 1487 138 1491 139
rect 1487 133 1491 134
rect 1535 138 1539 139
rect 1535 133 1539 134
rect 1567 138 1571 139
rect 1567 133 1571 134
rect 1591 138 1595 139
rect 1591 133 1595 134
rect 1647 138 1651 139
rect 1647 133 1651 134
rect 1655 138 1659 139
rect 1655 133 1659 134
rect 1703 138 1707 139
rect 1703 133 1707 134
rect 1735 138 1739 139
rect 1735 133 1739 134
rect 1759 138 1763 139
rect 1759 133 1763 134
rect 1374 131 1380 132
rect 1374 127 1375 131
rect 1379 127 1380 131
rect 1374 126 1380 127
rect 1390 131 1396 132
rect 1390 127 1391 131
rect 1395 127 1396 131
rect 1390 126 1396 127
rect 1366 113 1372 114
rect 1326 112 1332 113
rect 1326 108 1327 112
rect 1331 108 1332 112
rect 1366 109 1367 113
rect 1371 109 1372 113
rect 1392 112 1394 126
rect 1424 114 1426 133
rect 1446 131 1452 132
rect 1446 127 1447 131
rect 1451 127 1452 131
rect 1446 126 1452 127
rect 1422 113 1428 114
rect 1366 108 1372 109
rect 1390 111 1396 112
rect 110 107 116 108
rect 110 103 111 107
rect 115 103 116 107
rect 1286 107 1292 108
rect 1326 107 1332 108
rect 1390 107 1391 111
rect 1395 107 1396 111
rect 1422 109 1423 113
rect 1427 109 1428 113
rect 1448 112 1450 126
rect 1480 114 1482 133
rect 1502 131 1508 132
rect 1502 127 1503 131
rect 1507 127 1508 131
rect 1502 126 1508 127
rect 1478 113 1484 114
rect 1422 108 1428 109
rect 1446 111 1452 112
rect 110 102 116 103
rect 134 104 140 105
rect 112 99 114 102
rect 134 100 135 104
rect 139 100 140 104
rect 134 99 140 100
rect 190 104 196 105
rect 190 100 191 104
rect 195 100 196 104
rect 190 99 196 100
rect 246 104 252 105
rect 246 100 247 104
rect 251 100 252 104
rect 246 99 252 100
rect 302 104 308 105
rect 302 100 303 104
rect 307 100 308 104
rect 302 99 308 100
rect 358 104 364 105
rect 358 100 359 104
rect 363 100 364 104
rect 358 99 364 100
rect 414 104 420 105
rect 414 100 415 104
rect 419 100 420 104
rect 414 99 420 100
rect 470 104 476 105
rect 470 100 471 104
rect 475 100 476 104
rect 470 99 476 100
rect 526 104 532 105
rect 526 100 527 104
rect 531 100 532 104
rect 526 99 532 100
rect 582 104 588 105
rect 582 100 583 104
rect 587 100 588 104
rect 582 99 588 100
rect 638 104 644 105
rect 638 100 639 104
rect 643 100 644 104
rect 638 99 644 100
rect 694 104 700 105
rect 694 100 695 104
rect 699 100 700 104
rect 694 99 700 100
rect 750 104 756 105
rect 750 100 751 104
rect 755 100 756 104
rect 750 99 756 100
rect 814 104 820 105
rect 814 100 815 104
rect 819 100 820 104
rect 814 99 820 100
rect 878 104 884 105
rect 878 100 879 104
rect 883 100 884 104
rect 878 99 884 100
rect 942 104 948 105
rect 942 100 943 104
rect 947 100 948 104
rect 942 99 948 100
rect 1006 104 1012 105
rect 1006 100 1007 104
rect 1011 100 1012 104
rect 1006 99 1012 100
rect 1070 104 1076 105
rect 1070 100 1071 104
rect 1075 100 1076 104
rect 1070 99 1076 100
rect 1134 104 1140 105
rect 1134 100 1135 104
rect 1139 100 1140 104
rect 1286 103 1287 107
rect 1291 103 1292 107
rect 1390 106 1396 107
rect 1446 107 1447 111
rect 1451 107 1452 111
rect 1478 109 1479 113
rect 1483 109 1484 113
rect 1504 112 1506 126
rect 1536 114 1538 133
rect 1558 131 1564 132
rect 1558 127 1559 131
rect 1563 127 1564 131
rect 1558 126 1564 127
rect 1534 113 1540 114
rect 1478 108 1484 109
rect 1502 111 1508 112
rect 1446 106 1452 107
rect 1502 107 1503 111
rect 1507 107 1508 111
rect 1534 109 1535 113
rect 1539 109 1540 113
rect 1560 112 1562 126
rect 1592 114 1594 133
rect 1614 131 1620 132
rect 1614 127 1615 131
rect 1619 127 1620 131
rect 1614 126 1620 127
rect 1590 113 1596 114
rect 1534 108 1540 109
rect 1558 111 1564 112
rect 1502 106 1508 107
rect 1558 107 1559 111
rect 1563 107 1564 111
rect 1590 109 1591 113
rect 1595 109 1596 113
rect 1616 112 1618 126
rect 1648 114 1650 133
rect 1670 131 1676 132
rect 1670 127 1671 131
rect 1675 127 1676 131
rect 1670 126 1676 127
rect 1646 113 1652 114
rect 1590 108 1596 109
rect 1614 111 1620 112
rect 1558 106 1564 107
rect 1614 107 1615 111
rect 1619 107 1620 111
rect 1646 109 1647 113
rect 1651 109 1652 113
rect 1672 112 1674 126
rect 1704 114 1706 133
rect 1726 131 1732 132
rect 1726 127 1727 131
rect 1731 127 1732 131
rect 1726 126 1732 127
rect 1702 113 1708 114
rect 1646 108 1652 109
rect 1670 111 1676 112
rect 1614 106 1620 107
rect 1670 107 1671 111
rect 1675 107 1676 111
rect 1702 109 1703 113
rect 1707 109 1708 113
rect 1728 112 1730 126
rect 1760 114 1762 133
rect 1758 113 1764 114
rect 1702 108 1708 109
rect 1726 111 1732 112
rect 1670 106 1676 107
rect 1726 107 1727 111
rect 1731 107 1732 111
rect 1758 109 1759 113
rect 1763 109 1764 113
rect 1780 112 1782 158
rect 1824 139 1826 178
rect 1912 139 1914 178
rect 1966 163 1972 164
rect 1966 159 1967 163
rect 1971 159 1972 163
rect 1966 158 1972 159
rect 1823 138 1827 139
rect 1823 133 1827 134
rect 1879 138 1883 139
rect 1879 133 1883 134
rect 1911 138 1915 139
rect 1911 133 1915 134
rect 1943 138 1947 139
rect 1943 133 1947 134
rect 1824 114 1826 133
rect 1846 131 1852 132
rect 1846 127 1847 131
rect 1851 127 1852 131
rect 1846 126 1852 127
rect 1822 113 1828 114
rect 1758 108 1764 109
rect 1778 111 1784 112
rect 1726 106 1732 107
rect 1778 107 1779 111
rect 1783 107 1784 111
rect 1822 109 1823 113
rect 1827 109 1828 113
rect 1848 112 1850 126
rect 1880 114 1882 133
rect 1902 131 1908 132
rect 1902 127 1903 131
rect 1907 127 1908 131
rect 1902 126 1908 127
rect 1878 113 1884 114
rect 1822 108 1828 109
rect 1846 111 1852 112
rect 1778 106 1784 107
rect 1846 107 1847 111
rect 1851 107 1852 111
rect 1878 109 1879 113
rect 1883 109 1884 113
rect 1904 112 1906 126
rect 1944 114 1946 133
rect 1942 113 1948 114
rect 1878 108 1884 109
rect 1902 111 1908 112
rect 1846 106 1852 107
rect 1902 107 1903 111
rect 1907 107 1908 111
rect 1942 109 1943 113
rect 1947 109 1948 113
rect 1968 112 1970 158
rect 2008 139 2010 178
rect 2120 139 2122 178
rect 2007 138 2011 139
rect 2007 133 2011 134
rect 2071 138 2075 139
rect 2071 133 2075 134
rect 2119 138 2123 139
rect 2119 133 2123 134
rect 2008 114 2010 133
rect 2072 114 2074 133
rect 2128 132 2130 178
rect 2232 139 2234 178
rect 2328 164 2330 234
rect 2358 220 2364 221
rect 2358 216 2359 220
rect 2363 216 2364 220
rect 2358 215 2364 216
rect 2438 220 2444 221
rect 2438 216 2439 220
rect 2443 216 2444 220
rect 2438 215 2444 216
rect 2360 211 2362 215
rect 2440 211 2442 215
rect 2335 210 2339 211
rect 2335 205 2339 206
rect 2359 210 2363 211
rect 2359 205 2363 206
rect 2439 210 2443 211
rect 2439 205 2443 206
rect 2334 204 2340 205
rect 2334 200 2335 204
rect 2339 200 2340 204
rect 2334 199 2340 200
rect 2438 204 2444 205
rect 2438 200 2439 204
rect 2443 200 2444 204
rect 2438 199 2444 200
rect 2350 183 2356 184
rect 2350 179 2351 183
rect 2355 179 2356 183
rect 2350 178 2356 179
rect 2454 183 2460 184
rect 2454 179 2455 183
rect 2459 179 2460 183
rect 2454 178 2460 179
rect 2462 183 2468 184
rect 2462 179 2463 183
rect 2467 179 2468 183
rect 2462 178 2468 179
rect 2326 163 2332 164
rect 2326 159 2327 163
rect 2331 159 2332 163
rect 2326 158 2332 159
rect 2352 139 2354 178
rect 2456 139 2458 178
rect 2143 138 2147 139
rect 2143 133 2147 134
rect 2223 138 2227 139
rect 2223 133 2227 134
rect 2231 138 2235 139
rect 2231 133 2235 134
rect 2303 138 2307 139
rect 2303 133 2307 134
rect 2351 138 2355 139
rect 2351 133 2355 134
rect 2391 138 2395 139
rect 2391 133 2395 134
rect 2455 138 2459 139
rect 2455 133 2459 134
rect 2126 131 2132 132
rect 2126 127 2127 131
rect 2131 127 2132 131
rect 2126 126 2132 127
rect 2144 114 2146 133
rect 2166 131 2172 132
rect 2166 127 2167 131
rect 2171 127 2172 131
rect 2166 126 2172 127
rect 2006 113 2012 114
rect 1942 108 1948 109
rect 1966 111 1972 112
rect 1902 106 1908 107
rect 1966 107 1967 111
rect 1971 107 1972 111
rect 2006 109 2007 113
rect 2011 109 2012 113
rect 2006 108 2012 109
rect 2070 113 2076 114
rect 2070 109 2071 113
rect 2075 109 2076 113
rect 2070 108 2076 109
rect 2142 113 2148 114
rect 2142 109 2143 113
rect 2147 109 2148 113
rect 2168 112 2170 126
rect 2224 114 2226 133
rect 2246 131 2252 132
rect 2246 127 2247 131
rect 2251 127 2252 131
rect 2246 126 2252 127
rect 2222 113 2228 114
rect 2142 108 2148 109
rect 2166 111 2172 112
rect 1966 106 1972 107
rect 2166 107 2167 111
rect 2171 107 2172 111
rect 2222 109 2223 113
rect 2227 109 2228 113
rect 2248 112 2250 126
rect 2304 114 2306 133
rect 2392 114 2394 133
rect 2456 114 2458 133
rect 2464 132 2466 178
rect 2472 164 2474 234
rect 2502 223 2508 224
rect 2502 219 2503 223
rect 2507 219 2508 223
rect 2502 218 2508 219
rect 2504 211 2506 218
rect 2503 210 2507 211
rect 2503 205 2507 206
rect 2504 202 2506 205
rect 2502 201 2508 202
rect 2502 197 2503 201
rect 2507 197 2508 201
rect 2502 196 2508 197
rect 2502 184 2508 185
rect 2502 180 2503 184
rect 2507 180 2508 184
rect 2502 179 2508 180
rect 2470 163 2476 164
rect 2470 159 2471 163
rect 2475 159 2476 163
rect 2470 158 2476 159
rect 2504 139 2506 179
rect 2503 138 2507 139
rect 2503 133 2507 134
rect 2462 131 2468 132
rect 2462 127 2463 131
rect 2467 127 2468 131
rect 2462 126 2468 127
rect 2302 113 2308 114
rect 2222 108 2228 109
rect 2246 111 2252 112
rect 2166 106 2172 107
rect 2246 107 2247 111
rect 2251 107 2252 111
rect 2302 109 2303 113
rect 2307 109 2308 113
rect 2302 108 2308 109
rect 2390 113 2396 114
rect 2390 109 2391 113
rect 2395 109 2396 113
rect 2390 108 2396 109
rect 2454 113 2460 114
rect 2504 113 2506 133
rect 2454 109 2455 113
rect 2459 109 2460 113
rect 2454 108 2460 109
rect 2502 112 2508 113
rect 2502 108 2503 112
rect 2507 108 2508 112
rect 2502 107 2508 108
rect 2246 106 2252 107
rect 1286 102 1292 103
rect 1134 99 1140 100
rect 1288 99 1290 102
rect 111 98 115 99
rect 111 93 115 94
rect 135 98 139 99
rect 135 93 139 94
rect 191 98 195 99
rect 191 93 195 94
rect 247 98 251 99
rect 247 93 251 94
rect 303 98 307 99
rect 303 93 307 94
rect 359 98 363 99
rect 359 93 363 94
rect 415 98 419 99
rect 415 93 419 94
rect 471 98 475 99
rect 471 93 475 94
rect 527 98 531 99
rect 527 93 531 94
rect 583 98 587 99
rect 583 93 587 94
rect 639 98 643 99
rect 639 93 643 94
rect 695 98 699 99
rect 695 93 699 94
rect 751 98 755 99
rect 751 93 755 94
rect 815 98 819 99
rect 815 93 819 94
rect 879 98 883 99
rect 879 93 883 94
rect 943 98 947 99
rect 943 93 947 94
rect 1007 98 1011 99
rect 1007 93 1011 94
rect 1071 98 1075 99
rect 1071 93 1075 94
rect 1135 98 1139 99
rect 1135 93 1139 94
rect 1287 98 1291 99
rect 1287 93 1291 94
rect 1326 95 1332 96
rect 1326 91 1327 95
rect 1331 91 1332 95
rect 2502 95 2508 96
rect 1326 90 1332 91
rect 1350 92 1356 93
rect 1328 87 1330 90
rect 1350 88 1351 92
rect 1355 88 1356 92
rect 1350 87 1356 88
rect 1406 92 1412 93
rect 1406 88 1407 92
rect 1411 88 1412 92
rect 1406 87 1412 88
rect 1462 92 1468 93
rect 1462 88 1463 92
rect 1467 88 1468 92
rect 1462 87 1468 88
rect 1518 92 1524 93
rect 1518 88 1519 92
rect 1523 88 1524 92
rect 1518 87 1524 88
rect 1574 92 1580 93
rect 1574 88 1575 92
rect 1579 88 1580 92
rect 1574 87 1580 88
rect 1630 92 1636 93
rect 1630 88 1631 92
rect 1635 88 1636 92
rect 1630 87 1636 88
rect 1686 92 1692 93
rect 1686 88 1687 92
rect 1691 88 1692 92
rect 1686 87 1692 88
rect 1742 92 1748 93
rect 1742 88 1743 92
rect 1747 88 1748 92
rect 1742 87 1748 88
rect 1806 92 1812 93
rect 1806 88 1807 92
rect 1811 88 1812 92
rect 1806 87 1812 88
rect 1862 92 1868 93
rect 1862 88 1863 92
rect 1867 88 1868 92
rect 1862 87 1868 88
rect 1926 92 1932 93
rect 1926 88 1927 92
rect 1931 88 1932 92
rect 1926 87 1932 88
rect 1990 92 1996 93
rect 1990 88 1991 92
rect 1995 88 1996 92
rect 1990 87 1996 88
rect 2054 92 2060 93
rect 2054 88 2055 92
rect 2059 88 2060 92
rect 2054 87 2060 88
rect 2126 92 2132 93
rect 2126 88 2127 92
rect 2131 88 2132 92
rect 2126 87 2132 88
rect 2206 92 2212 93
rect 2206 88 2207 92
rect 2211 88 2212 92
rect 2206 87 2212 88
rect 2286 92 2292 93
rect 2286 88 2287 92
rect 2291 88 2292 92
rect 2286 87 2292 88
rect 2374 92 2380 93
rect 2374 88 2375 92
rect 2379 88 2380 92
rect 2374 87 2380 88
rect 2438 92 2444 93
rect 2438 88 2439 92
rect 2443 88 2444 92
rect 2502 91 2503 95
rect 2507 91 2508 95
rect 2502 90 2508 91
rect 2438 87 2444 88
rect 2504 87 2506 90
rect 1327 86 1331 87
rect 1327 81 1331 82
rect 1351 86 1355 87
rect 1351 81 1355 82
rect 1407 86 1411 87
rect 1407 81 1411 82
rect 1463 86 1467 87
rect 1463 81 1467 82
rect 1519 86 1523 87
rect 1519 81 1523 82
rect 1575 86 1579 87
rect 1575 81 1579 82
rect 1631 86 1635 87
rect 1631 81 1635 82
rect 1687 86 1691 87
rect 1687 81 1691 82
rect 1743 86 1747 87
rect 1743 81 1747 82
rect 1807 86 1811 87
rect 1807 81 1811 82
rect 1863 86 1867 87
rect 1863 81 1867 82
rect 1927 86 1931 87
rect 1927 81 1931 82
rect 1991 86 1995 87
rect 1991 81 1995 82
rect 2055 86 2059 87
rect 2055 81 2059 82
rect 2127 86 2131 87
rect 2127 81 2131 82
rect 2207 86 2211 87
rect 2207 81 2211 82
rect 2287 86 2291 87
rect 2287 81 2291 82
rect 2375 86 2379 87
rect 2375 81 2379 82
rect 2439 86 2443 87
rect 2439 81 2443 82
rect 2503 86 2507 87
rect 2503 81 2507 82
<< m4c >>
rect 111 2578 115 2582
rect 135 2578 139 2582
rect 191 2578 195 2582
rect 247 2578 251 2582
rect 303 2578 307 2582
rect 359 2578 363 2582
rect 1287 2578 1291 2582
rect 1327 2558 1331 2562
rect 1495 2558 1499 2562
rect 1551 2558 1555 2562
rect 1607 2558 1611 2562
rect 1663 2558 1667 2562
rect 1719 2558 1723 2562
rect 1775 2558 1779 2562
rect 1831 2558 1835 2562
rect 1887 2558 1891 2562
rect 1943 2558 1947 2562
rect 1999 2558 2003 2562
rect 2055 2558 2059 2562
rect 2111 2558 2115 2562
rect 2167 2558 2171 2562
rect 2503 2558 2507 2562
rect 111 2526 115 2530
rect 151 2526 155 2530
rect 207 2526 211 2530
rect 223 2526 227 2530
rect 263 2526 267 2530
rect 279 2526 283 2530
rect 319 2526 323 2530
rect 343 2526 347 2530
rect 375 2526 379 2530
rect 415 2526 419 2530
rect 487 2526 491 2530
rect 551 2526 555 2530
rect 615 2526 619 2530
rect 679 2526 683 2530
rect 743 2526 747 2530
rect 807 2526 811 2530
rect 871 2526 875 2530
rect 935 2526 939 2530
rect 999 2526 1003 2530
rect 1063 2526 1067 2530
rect 1287 2526 1291 2530
rect 111 2466 115 2470
rect 167 2466 171 2470
rect 207 2466 211 2470
rect 223 2466 227 2470
rect 263 2466 267 2470
rect 279 2466 283 2470
rect 327 2466 331 2470
rect 335 2466 339 2470
rect 391 2466 395 2470
rect 399 2466 403 2470
rect 447 2466 451 2470
rect 471 2466 475 2470
rect 503 2466 507 2470
rect 535 2466 539 2470
rect 559 2466 563 2470
rect 1327 2506 1331 2510
rect 1911 2520 1915 2524
rect 1511 2506 1515 2510
rect 599 2466 603 2470
rect 615 2466 619 2470
rect 663 2466 667 2470
rect 671 2466 675 2470
rect 727 2466 731 2470
rect 783 2466 787 2470
rect 791 2466 795 2470
rect 839 2466 843 2470
rect 855 2466 859 2470
rect 895 2466 899 2470
rect 919 2466 923 2470
rect 951 2466 955 2470
rect 983 2466 987 2470
rect 1007 2466 1011 2470
rect 1047 2466 1051 2470
rect 1063 2466 1067 2470
rect 167 2448 171 2452
rect 495 2448 499 2452
rect 567 2448 571 2452
rect 875 2448 879 2452
rect 111 2402 115 2406
rect 183 2402 187 2406
rect 239 2402 243 2406
rect 295 2402 299 2406
rect 351 2402 355 2406
rect 407 2402 411 2406
rect 463 2402 467 2406
rect 519 2402 523 2406
rect 575 2402 579 2406
rect 631 2402 635 2406
rect 687 2402 691 2406
rect 743 2402 747 2406
rect 799 2402 803 2406
rect 855 2402 859 2406
rect 911 2402 915 2406
rect 1543 2506 1547 2510
rect 1567 2506 1571 2510
rect 1607 2506 1611 2510
rect 1623 2506 1627 2510
rect 1679 2506 1683 2510
rect 1735 2506 1739 2510
rect 1751 2506 1755 2510
rect 1791 2506 1795 2510
rect 1823 2506 1827 2510
rect 1847 2506 1851 2510
rect 1895 2506 1899 2510
rect 1903 2506 1907 2510
rect 1527 2488 1531 2492
rect 1287 2466 1291 2470
rect 1327 2450 1331 2454
rect 1527 2450 1531 2454
rect 1543 2450 1547 2454
rect 1843 2488 1847 2492
rect 2191 2520 2195 2524
rect 1959 2506 1963 2510
rect 1967 2506 1971 2510
rect 2015 2506 2019 2510
rect 2039 2506 2043 2510
rect 2071 2506 2075 2510
rect 2111 2506 2115 2510
rect 2127 2506 2131 2510
rect 2183 2506 2187 2510
rect 2503 2506 2507 2510
rect 1591 2450 1595 2454
rect 1607 2450 1611 2454
rect 1663 2450 1667 2454
rect 1671 2450 1675 2454
rect 1735 2450 1739 2454
rect 1743 2450 1747 2454
rect 1807 2450 1811 2454
rect 1815 2450 1819 2454
rect 1879 2450 1883 2454
rect 1951 2450 1955 2454
rect 2023 2450 2027 2454
rect 2095 2450 2099 2454
rect 2167 2450 2171 2454
rect 967 2402 971 2406
rect 1023 2402 1027 2406
rect 1079 2402 1083 2406
rect 1287 2402 1291 2406
rect 1327 2394 1331 2398
rect 1559 2394 1563 2398
rect 1567 2394 1571 2398
rect 1623 2394 1627 2398
rect 1679 2394 1683 2398
rect 1687 2394 1691 2398
rect 1735 2394 1739 2398
rect 1759 2394 1763 2398
rect 1791 2394 1795 2398
rect 111 2342 115 2346
rect 319 2342 323 2346
rect 391 2342 395 2346
rect 463 2342 467 2346
rect 503 2342 507 2346
rect 535 2342 539 2346
rect 111 2282 115 2286
rect 175 2282 179 2286
rect 271 2282 275 2286
rect 335 2282 339 2286
rect 375 2282 379 2286
rect 407 2282 411 2286
rect 559 2342 563 2346
rect 607 2342 611 2346
rect 615 2342 619 2346
rect 671 2342 675 2346
rect 679 2342 683 2346
rect 743 2342 747 2346
rect 807 2342 811 2346
rect 863 2342 867 2346
rect 927 2342 931 2346
rect 991 2342 995 2346
rect 1055 2342 1059 2346
rect 1111 2342 1115 2346
rect 1167 2342 1171 2346
rect 1223 2342 1227 2346
rect 1287 2342 1291 2346
rect 1327 2334 1331 2338
rect 1471 2334 1475 2338
rect 1535 2334 1539 2338
rect 1551 2334 1555 2338
rect 1607 2334 1611 2338
rect 1663 2334 1667 2338
rect 1687 2334 1691 2338
rect 1719 2334 1723 2338
rect 1759 2334 1763 2338
rect 1775 2334 1779 2338
rect 479 2282 483 2286
rect 551 2282 555 2286
rect 591 2282 595 2286
rect 623 2282 627 2286
rect 695 2282 699 2286
rect 703 2282 707 2286
rect 759 2282 763 2286
rect 807 2282 811 2286
rect 823 2282 827 2286
rect 879 2282 883 2286
rect 911 2282 915 2286
rect 943 2282 947 2286
rect 1007 2282 1011 2286
rect 1015 2282 1019 2286
rect 1071 2282 1075 2286
rect 1127 2282 1131 2286
rect 1183 2282 1187 2286
rect 1239 2282 1243 2286
rect 111 2230 115 2234
rect 143 2230 147 2234
rect 159 2230 163 2234
rect 231 2230 235 2234
rect 255 2230 259 2234
rect 319 2230 323 2234
rect 359 2230 363 2234
rect 415 2230 419 2234
rect 463 2230 467 2234
rect 519 2230 523 2234
rect 575 2230 579 2234
rect 623 2230 627 2234
rect 687 2230 691 2234
rect 727 2230 731 2234
rect 791 2230 795 2234
rect 831 2230 835 2234
rect 895 2230 899 2234
rect 111 2178 115 2182
rect 159 2178 163 2182
rect 247 2178 251 2182
rect 255 2178 259 2182
rect 335 2178 339 2182
rect 351 2178 355 2182
rect 431 2178 435 2182
rect 455 2178 459 2182
rect 535 2178 539 2182
rect 559 2178 563 2182
rect 639 2178 643 2182
rect 935 2230 939 2234
rect 999 2230 1003 2234
rect 1039 2230 1043 2234
rect 1831 2394 1835 2398
rect 1855 2394 1859 2398
rect 1895 2394 1899 2398
rect 1919 2394 1923 2398
rect 1967 2394 1971 2398
rect 2503 2450 2507 2454
rect 1983 2394 1987 2398
rect 2039 2394 2043 2398
rect 2047 2394 2051 2398
rect 2111 2394 2115 2398
rect 2183 2394 2187 2398
rect 2503 2394 2507 2398
rect 1831 2334 1835 2338
rect 1839 2334 1843 2338
rect 1287 2282 1291 2286
rect 1327 2282 1331 2286
rect 1383 2282 1387 2286
rect 1479 2282 1483 2286
rect 1903 2334 1907 2338
rect 1967 2334 1971 2338
rect 1983 2334 1987 2338
rect 2031 2334 2035 2338
rect 2063 2334 2067 2338
rect 2095 2334 2099 2338
rect 2143 2334 2147 2338
rect 2503 2334 2507 2338
rect 1487 2282 1491 2286
rect 1111 2230 1115 2234
rect 1143 2230 1147 2234
rect 1223 2230 1227 2234
rect 1287 2230 1291 2234
rect 1327 2230 1331 2234
rect 1367 2230 1371 2234
rect 1551 2282 1555 2286
rect 1583 2282 1587 2286
rect 1623 2282 1627 2286
rect 1687 2282 1691 2286
rect 1703 2282 1707 2286
rect 1775 2282 1779 2286
rect 1791 2282 1795 2286
rect 1847 2282 1851 2286
rect 1903 2282 1907 2286
rect 1919 2282 1923 2286
rect 1999 2282 2003 2286
rect 2015 2282 2019 2286
rect 2079 2282 2083 2286
rect 2127 2282 2131 2286
rect 2159 2282 2163 2286
rect 2239 2282 2243 2286
rect 2503 2282 2507 2286
rect 1463 2230 1467 2234
rect 1487 2230 1491 2234
rect 1567 2230 1571 2234
rect 1607 2230 1611 2234
rect 1671 2230 1675 2234
rect 1719 2230 1723 2234
rect 1775 2230 1779 2234
rect 1815 2230 1819 2234
rect 1887 2230 1891 2234
rect 1903 2230 1907 2234
rect 1983 2230 1987 2234
rect 1999 2230 2003 2234
rect 2055 2230 2059 2234
rect 2111 2230 2115 2234
rect 2127 2230 2131 2234
rect 2191 2230 2195 2234
rect 2223 2230 2227 2234
rect 2255 2230 2259 2234
rect 2319 2230 2323 2234
rect 2383 2230 2387 2234
rect 2439 2230 2443 2234
rect 2503 2230 2507 2234
rect 1719 2216 1723 2220
rect 2247 2216 2251 2220
rect 663 2178 667 2182
rect 743 2178 747 2182
rect 767 2178 771 2182
rect 847 2178 851 2182
rect 863 2178 867 2182
rect 951 2178 955 2182
rect 959 2178 963 2182
rect 1055 2178 1059 2182
rect 1159 2178 1163 2182
rect 1239 2178 1243 2182
rect 1287 2178 1291 2182
rect 111 2126 115 2130
rect 239 2126 243 2130
rect 303 2126 307 2130
rect 335 2126 339 2130
rect 359 2126 363 2130
rect 423 2126 427 2130
rect 439 2126 443 2130
rect 487 2126 491 2130
rect 543 2126 547 2130
rect 559 2126 563 2130
rect 631 2126 635 2130
rect 647 2126 651 2130
rect 711 2126 715 2130
rect 751 2126 755 2130
rect 799 2126 803 2130
rect 847 2126 851 2130
rect 887 2126 891 2130
rect 943 2126 947 2130
rect 975 2126 979 2130
rect 111 2070 115 2074
rect 319 2070 323 2074
rect 375 2070 379 2074
rect 399 2070 403 2074
rect 439 2070 443 2074
rect 455 2070 459 2074
rect 503 2070 507 2074
rect 511 2070 515 2074
rect 575 2070 579 2074
rect 639 2070 643 2074
rect 647 2070 651 2074
rect 711 2070 715 2074
rect 727 2070 731 2074
rect 791 2070 795 2074
rect 815 2070 819 2074
rect 1039 2126 1043 2130
rect 1063 2126 1067 2130
rect 1143 2126 1147 2130
rect 1151 2126 1155 2130
rect 1223 2126 1227 2130
rect 1327 2158 1331 2162
rect 1383 2158 1387 2162
rect 1407 2158 1411 2162
rect 1503 2158 1507 2162
rect 1623 2158 1627 2162
rect 1735 2158 1739 2162
rect 1815 2158 1819 2162
rect 1831 2158 1835 2162
rect 1919 2158 1923 2162
rect 1991 2158 1995 2162
rect 1999 2158 2003 2162
rect 2071 2158 2075 2162
rect 2143 2158 2147 2162
rect 2159 2158 2163 2162
rect 2207 2158 2211 2162
rect 2271 2158 2275 2162
rect 2319 2158 2323 2162
rect 2335 2158 2339 2162
rect 2399 2158 2403 2162
rect 2455 2158 2459 2162
rect 1287 2126 1291 2130
rect 1327 2106 1331 2110
rect 1383 2106 1387 2110
rect 1391 2106 1395 2110
rect 1551 2106 1555 2110
rect 1607 2106 1611 2110
rect 1711 2106 1715 2110
rect 863 2070 867 2074
rect 903 2070 907 2074
rect 943 2070 947 2074
rect 991 2070 995 2074
rect 1023 2070 1027 2074
rect 1079 2070 1083 2074
rect 1103 2070 1107 2074
rect 111 2014 115 2018
rect 231 2014 235 2018
rect 287 2014 291 2018
rect 359 2014 363 2018
rect 383 2014 387 2018
rect 231 1976 235 1980
rect 111 1958 115 1962
rect 151 1958 155 1962
rect 215 1958 219 1962
rect 247 1958 251 1962
rect 303 1958 307 1962
rect 319 1958 323 1962
rect 375 1958 379 1962
rect 167 1936 171 1940
rect 439 2014 443 2018
rect 495 2014 499 2018
rect 535 2014 539 2018
rect 559 2014 563 2018
rect 623 2014 627 2018
rect 631 2014 635 2018
rect 695 2014 699 2018
rect 655 1976 659 1980
rect 735 2014 739 2018
rect 775 2014 779 2018
rect 847 2014 851 2018
rect 927 2014 931 2018
rect 959 2014 963 2018
rect 2503 2158 2507 2162
rect 1799 2106 1803 2110
rect 1855 2106 1859 2110
rect 1975 2106 1979 2110
rect 1991 2106 1995 2110
rect 1167 2070 1171 2074
rect 1183 2070 1187 2074
rect 1239 2070 1243 2074
rect 1287 2070 1291 2074
rect 1327 2050 1331 2054
rect 1399 2050 1403 2054
rect 1447 2050 1451 2054
rect 1551 2050 1555 2054
rect 1567 2050 1571 2054
rect 1655 2050 1659 2054
rect 1727 2050 1731 2054
rect 1751 2050 1755 2054
rect 1839 2050 1843 2054
rect 1871 2050 1875 2054
rect 1007 2014 1011 2018
rect 1079 2014 1083 2018
rect 1087 2014 1091 2018
rect 1167 2014 1171 2018
rect 1199 2014 1203 2018
rect 1223 2014 1227 2018
rect 1287 2014 1291 2018
rect 1327 1994 1331 1998
rect 1431 1994 1435 1998
rect 1455 1994 1459 1998
rect 1511 1994 1515 1998
rect 1535 1994 1539 1998
rect 439 1958 443 1962
rect 455 1958 459 1962
rect 551 1958 555 1962
rect 583 1958 587 1962
rect 647 1958 651 1962
rect 743 1958 747 1962
rect 751 1958 755 1962
rect 863 1958 867 1962
rect 603 1936 607 1940
rect 919 1958 923 1962
rect 975 1958 979 1962
rect 1095 1958 1099 1962
rect 111 1898 115 1902
rect 135 1898 139 1902
rect 191 1898 195 1902
rect 199 1898 203 1902
rect 271 1898 275 1902
rect 303 1898 307 1902
rect 111 1846 115 1850
rect 151 1846 155 1850
rect 359 1898 363 1902
rect 423 1898 427 1902
rect 455 1898 459 1902
rect 543 1898 547 1902
rect 567 1898 571 1902
rect 631 1898 635 1902
rect 719 1898 723 1902
rect 727 1898 731 1902
rect 207 1846 211 1850
rect 287 1846 291 1850
rect 295 1846 299 1850
rect 375 1846 379 1850
rect 391 1846 395 1850
rect 471 1846 475 1850
rect 495 1846 499 1850
rect 559 1846 563 1850
rect 799 1898 803 1902
rect 871 1898 875 1902
rect 903 1898 907 1902
rect 943 1898 947 1902
rect 1015 1898 1019 1902
rect 2119 2106 2123 2110
rect 2143 2106 2147 2110
rect 2239 2106 2243 2110
rect 2303 2106 2307 2110
rect 2367 2106 2371 2110
rect 2439 2106 2443 2110
rect 2503 2106 2507 2110
rect 1927 2050 1931 2054
rect 2007 2050 2011 2054
rect 2023 2050 2027 2054
rect 2119 2050 2123 2054
rect 2135 2050 2139 2054
rect 2255 2050 2259 2054
rect 2383 2050 2387 2054
rect 2503 2050 2507 2054
rect 1575 1994 1579 1998
rect 1639 1994 1643 1998
rect 1703 1994 1707 1998
rect 1735 1994 1739 1998
rect 1767 1994 1771 1998
rect 1215 1958 1219 1962
rect 1287 1958 1291 1962
rect 1327 1938 1331 1942
rect 1471 1938 1475 1942
rect 1527 1938 1531 1942
rect 1567 1938 1571 1942
rect 1591 1938 1595 1942
rect 1631 1938 1635 1942
rect 1655 1938 1659 1942
rect 1703 1938 1707 1942
rect 1823 1994 1827 1998
rect 1831 1994 1835 1998
rect 1895 1994 1899 1998
rect 1911 1994 1915 1998
rect 1959 1994 1963 1998
rect 2007 1994 2011 1998
rect 2031 1994 2035 1998
rect 2103 1994 2107 1998
rect 2503 1994 2507 1998
rect 1719 1938 1723 1942
rect 1775 1938 1779 1942
rect 1783 1938 1787 1942
rect 1847 1938 1851 1942
rect 1911 1938 1915 1942
rect 1919 1938 1923 1942
rect 1975 1938 1979 1942
rect 1999 1938 2003 1942
rect 2047 1938 2051 1942
rect 2087 1938 2091 1942
rect 2183 1938 2187 1942
rect 2279 1938 2283 1942
rect 2375 1938 2379 1942
rect 2455 1938 2459 1942
rect 2503 1938 2507 1942
rect 1079 1898 1083 1902
rect 1087 1898 1091 1902
rect 1159 1898 1163 1902
rect 1287 1898 1291 1902
rect 1327 1882 1331 1886
rect 1551 1882 1555 1886
rect 1607 1882 1611 1886
rect 1615 1882 1619 1886
rect 1663 1882 1667 1886
rect 1687 1882 1691 1886
rect 1727 1882 1731 1886
rect 1759 1882 1763 1886
rect 591 1846 595 1850
rect 647 1846 651 1850
rect 687 1846 691 1850
rect 735 1846 739 1850
rect 775 1846 779 1850
rect 815 1846 819 1850
rect 855 1846 859 1850
rect 887 1846 891 1850
rect 927 1846 931 1850
rect 111 1782 115 1786
rect 135 1782 139 1786
rect 191 1782 195 1786
rect 199 1782 203 1786
rect 279 1782 283 1786
rect 295 1782 299 1786
rect 375 1782 379 1786
rect 399 1782 403 1786
rect 479 1782 483 1786
rect 503 1782 507 1786
rect 575 1782 579 1786
rect 607 1782 611 1786
rect 135 1768 139 1772
rect 511 1768 515 1772
rect 111 1726 115 1730
rect 151 1726 155 1730
rect 167 1726 171 1730
rect 215 1726 219 1730
rect 239 1726 243 1730
rect 311 1726 315 1730
rect 319 1726 323 1730
rect 407 1726 411 1730
rect 415 1726 419 1730
rect 503 1726 507 1730
rect 519 1726 523 1730
rect 671 1782 675 1786
rect 703 1782 707 1786
rect 759 1782 763 1786
rect 799 1782 803 1786
rect 839 1782 843 1786
rect 887 1782 891 1786
rect 911 1782 915 1786
rect 959 1846 963 1850
rect 1799 1882 1803 1886
rect 1831 1882 1835 1886
rect 1871 1882 1875 1886
rect 1903 1882 1907 1886
rect 1943 1882 1947 1886
rect 1983 1882 1987 1886
rect 2007 1882 2011 1886
rect 2071 1882 2075 1886
rect 2135 1882 2139 1886
rect 2167 1882 2171 1886
rect 2199 1882 2203 1886
rect 2263 1882 2267 1886
rect 999 1846 1003 1850
rect 1031 1846 1035 1850
rect 1079 1846 1083 1850
rect 1103 1846 1107 1850
rect 1159 1846 1163 1850
rect 1175 1846 1179 1850
rect 1287 1846 1291 1850
rect 1327 1826 1331 1830
rect 1623 1826 1627 1830
rect 1631 1826 1635 1830
rect 1679 1826 1683 1830
rect 1719 1826 1723 1830
rect 1743 1826 1747 1830
rect 1815 1826 1819 1830
rect 1887 1826 1891 1830
rect 1927 1826 1931 1830
rect 1959 1826 1963 1830
rect 975 1782 979 1786
rect 983 1782 987 1786
rect 1063 1782 1067 1786
rect 1143 1782 1147 1786
rect 1151 1782 1155 1786
rect 607 1726 611 1730
rect 623 1726 627 1730
rect 711 1726 715 1730
rect 719 1726 723 1730
rect 815 1726 819 1730
rect 823 1726 827 1730
rect 903 1726 907 1730
rect 935 1726 939 1730
rect 111 1670 115 1674
rect 151 1670 155 1674
rect 223 1670 227 1674
rect 255 1670 259 1674
rect 303 1670 307 1674
rect 319 1670 323 1674
rect 391 1670 395 1674
rect 399 1670 403 1674
rect 487 1670 491 1674
rect 575 1670 579 1674
rect 591 1670 595 1674
rect 111 1614 115 1618
rect 271 1614 275 1618
rect 303 1614 307 1618
rect 335 1614 339 1618
rect 359 1614 363 1618
rect 415 1614 419 1618
rect 431 1614 435 1618
rect 503 1614 507 1618
rect 511 1614 515 1618
rect 591 1614 595 1618
rect 599 1614 603 1618
rect 111 1562 115 1566
rect 247 1562 251 1566
rect 671 1670 675 1674
rect 695 1670 699 1674
rect 767 1670 771 1674
rect 807 1670 811 1674
rect 863 1670 867 1674
rect 991 1726 995 1730
rect 1287 1782 1291 1786
rect 1327 1774 1331 1778
rect 1527 1774 1531 1778
rect 1607 1774 1611 1778
rect 1615 1774 1619 1778
rect 2327 1882 2331 1886
rect 2359 1882 2363 1886
rect 2383 1882 2387 1886
rect 2439 1882 2443 1886
rect 2023 1826 2027 1830
rect 2055 1826 2059 1830
rect 2087 1826 2091 1830
rect 2151 1826 2155 1830
rect 2191 1826 2195 1830
rect 2215 1826 2219 1830
rect 2279 1826 2283 1830
rect 2335 1826 2339 1830
rect 2343 1826 2347 1830
rect 2399 1826 2403 1830
rect 2455 1826 2459 1830
rect 1695 1774 1699 1778
rect 1703 1774 1707 1778
rect 1791 1774 1795 1778
rect 1799 1774 1803 1778
rect 1879 1774 1883 1778
rect 1911 1774 1915 1778
rect 1967 1774 1971 1778
rect 2039 1774 2043 1778
rect 2055 1774 2059 1778
rect 2135 1774 2139 1778
rect 2175 1774 2179 1778
rect 1655 1752 1659 1756
rect 1915 1752 1919 1756
rect 1047 1726 1051 1730
rect 1079 1726 1083 1730
rect 1159 1726 1163 1730
rect 1167 1726 1171 1730
rect 1287 1726 1291 1730
rect 1327 1718 1331 1722
rect 1399 1718 1403 1722
rect 1463 1718 1467 1722
rect 1543 1718 1547 1722
rect 919 1670 923 1674
rect 959 1670 963 1674
rect 1031 1670 1035 1674
rect 1063 1670 1067 1674
rect 1143 1670 1147 1674
rect 1167 1670 1171 1674
rect 687 1614 691 1618
rect 695 1614 699 1618
rect 287 1562 291 1566
rect 319 1562 323 1566
rect 343 1562 347 1566
rect 399 1562 403 1566
rect 415 1562 419 1566
rect 111 1502 115 1506
rect 263 1502 267 1506
rect 279 1502 283 1506
rect 335 1502 339 1506
rect 343 1502 347 1506
rect 487 1562 491 1566
rect 495 1562 499 1566
rect 583 1562 587 1566
rect 671 1562 675 1566
rect 679 1562 683 1566
rect 783 1614 787 1618
rect 791 1614 795 1618
rect 879 1614 883 1618
rect 895 1614 899 1618
rect 759 1562 763 1566
rect 775 1562 779 1566
rect 975 1614 979 1618
rect 1007 1614 1011 1618
rect 1079 1614 1083 1618
rect 1287 1670 1291 1674
rect 1327 1662 1331 1666
rect 1351 1662 1355 1666
rect 1383 1662 1387 1666
rect 1407 1662 1411 1666
rect 1623 1718 1627 1722
rect 1631 1718 1635 1722
rect 1711 1718 1715 1722
rect 1727 1718 1731 1722
rect 1807 1718 1811 1722
rect 1823 1718 1827 1722
rect 1895 1718 1899 1722
rect 1919 1718 1923 1722
rect 1983 1718 1987 1722
rect 2015 1718 2019 1722
rect 2071 1718 2075 1722
rect 1595 1696 1599 1700
rect 1843 1696 1847 1700
rect 2215 1774 2219 1778
rect 2295 1774 2299 1778
rect 2319 1774 2323 1778
rect 2503 1882 2507 1886
rect 2503 1826 2507 1830
rect 2375 1774 2379 1778
rect 2439 1774 2443 1778
rect 2111 1718 2115 1722
rect 2151 1718 2155 1722
rect 2199 1718 2203 1722
rect 2231 1718 2235 1722
rect 2287 1718 2291 1722
rect 2311 1718 2315 1722
rect 2383 1718 2387 1722
rect 2391 1718 2395 1722
rect 2455 1718 2459 1722
rect 2503 1774 2507 1778
rect 2503 1718 2507 1722
rect 1447 1662 1451 1666
rect 1495 1662 1499 1666
rect 1527 1662 1531 1666
rect 1583 1662 1587 1666
rect 1615 1662 1619 1666
rect 1679 1662 1683 1666
rect 1711 1662 1715 1666
rect 1783 1662 1787 1666
rect 1807 1662 1811 1666
rect 1895 1662 1899 1666
rect 1903 1662 1907 1666
rect 1999 1662 2003 1666
rect 2023 1662 2027 1666
rect 1415 1640 1419 1644
rect 1703 1640 1707 1644
rect 1119 1614 1123 1618
rect 1183 1614 1187 1618
rect 1287 1614 1291 1618
rect 847 1562 851 1566
rect 879 1562 883 1566
rect 927 1562 931 1566
rect 991 1562 995 1566
rect 1007 1562 1011 1566
rect 415 1502 419 1506
rect 495 1502 499 1506
rect 503 1502 507 1506
rect 575 1502 579 1506
rect 599 1502 603 1506
rect 655 1502 659 1506
rect 111 1446 115 1450
rect 191 1446 195 1450
rect 255 1446 259 1450
rect 263 1446 267 1450
rect 327 1446 331 1450
rect 399 1446 403 1450
rect 407 1446 411 1450
rect 479 1446 483 1450
rect 503 1446 507 1450
rect 559 1446 563 1450
rect 607 1446 611 1450
rect 687 1502 691 1506
rect 735 1502 739 1506
rect 775 1502 779 1506
rect 815 1502 819 1506
rect 863 1502 867 1506
rect 1087 1562 1091 1566
rect 1103 1562 1107 1566
rect 1167 1562 1171 1566
rect 1223 1562 1227 1566
rect 1327 1610 1331 1614
rect 1367 1610 1371 1614
rect 1423 1610 1427 1614
rect 1479 1610 1483 1614
rect 1511 1610 1515 1614
rect 1559 1610 1563 1614
rect 1599 1610 1603 1614
rect 1639 1610 1643 1614
rect 1695 1610 1699 1614
rect 1719 1610 1723 1614
rect 1791 1610 1795 1614
rect 1799 1610 1803 1614
rect 1871 1610 1875 1614
rect 1911 1610 1915 1614
rect 2095 1662 2099 1666
rect 2159 1662 2163 1666
rect 2183 1662 2187 1666
rect 2271 1662 2275 1666
rect 2303 1662 2307 1666
rect 2367 1662 2371 1666
rect 2439 1662 2443 1666
rect 2503 1662 2507 1666
rect 1951 1610 1955 1614
rect 2031 1610 2035 1614
rect 2039 1610 2043 1614
rect 2175 1610 2179 1614
rect 2319 1610 2323 1614
rect 2455 1610 2459 1614
rect 2503 1610 2507 1614
rect 1287 1562 1291 1566
rect 1327 1558 1331 1562
rect 1351 1558 1355 1562
rect 1407 1558 1411 1562
rect 1463 1558 1467 1562
rect 1471 1558 1475 1562
rect 1543 1558 1547 1562
rect 1607 1558 1611 1562
rect 1623 1558 1627 1562
rect 1703 1558 1707 1562
rect 1735 1558 1739 1562
rect 1775 1558 1779 1562
rect 1855 1558 1859 1562
rect 1871 1558 1875 1562
rect 1935 1558 1939 1562
rect 2007 1558 2011 1562
rect 2015 1558 2019 1562
rect 2503 1558 2507 1562
rect 895 1502 899 1506
rect 943 1502 947 1506
rect 975 1502 979 1506
rect 1023 1502 1027 1506
rect 1055 1502 1059 1506
rect 1103 1502 1107 1506
rect 1143 1502 1147 1506
rect 1183 1502 1187 1506
rect 1239 1502 1243 1506
rect 1287 1502 1291 1506
rect 1327 1506 1331 1510
rect 1367 1506 1371 1510
rect 639 1446 643 1450
rect 711 1446 715 1450
rect 719 1446 723 1450
rect 799 1446 803 1450
rect 815 1446 819 1450
rect 1423 1506 1427 1510
rect 1479 1506 1483 1510
rect 1487 1506 1491 1510
rect 1551 1506 1555 1510
rect 1623 1506 1627 1510
rect 1631 1506 1635 1510
rect 1711 1506 1715 1510
rect 1751 1506 1755 1510
rect 879 1446 883 1450
rect 919 1446 923 1450
rect 959 1446 963 1450
rect 1023 1446 1027 1450
rect 1039 1446 1043 1450
rect 1127 1446 1131 1450
rect 111 1390 115 1394
rect 151 1390 155 1394
rect 207 1390 211 1394
rect 223 1390 227 1394
rect 271 1390 275 1394
rect 295 1390 299 1394
rect 343 1390 347 1394
rect 359 1390 363 1394
rect 423 1390 427 1394
rect 431 1390 435 1394
rect 503 1390 507 1394
rect 519 1390 523 1394
rect 583 1390 587 1394
rect 623 1390 627 1394
rect 663 1390 667 1394
rect 111 1322 115 1326
rect 135 1322 139 1326
rect 207 1322 211 1326
rect 239 1322 243 1326
rect 111 1262 115 1266
rect 151 1262 155 1266
rect 279 1322 283 1326
rect 343 1322 347 1326
rect 367 1322 371 1326
rect 415 1322 419 1326
rect 479 1322 483 1326
rect 487 1322 491 1326
rect 567 1322 571 1326
rect 583 1322 587 1326
rect 647 1322 651 1326
rect 727 1390 731 1394
rect 751 1390 755 1394
rect 831 1390 835 1394
rect 839 1390 843 1394
rect 1223 1446 1227 1450
rect 1287 1446 1291 1450
rect 1327 1446 1331 1450
rect 1351 1446 1355 1450
rect 1359 1446 1363 1450
rect 1407 1446 1411 1450
rect 1447 1446 1451 1450
rect 1463 1446 1467 1450
rect 1535 1446 1539 1450
rect 1791 1506 1795 1510
rect 1871 1506 1875 1510
rect 1887 1506 1891 1510
rect 1951 1506 1955 1510
rect 2023 1506 2027 1510
rect 2031 1506 2035 1510
rect 2119 1506 2123 1510
rect 2503 1506 2507 1510
rect 1615 1446 1619 1450
rect 1631 1446 1635 1450
rect 1695 1446 1699 1450
rect 1727 1446 1731 1450
rect 1775 1446 1779 1450
rect 1815 1446 1819 1450
rect 927 1390 931 1394
rect 935 1390 939 1394
rect 1015 1390 1019 1394
rect 1039 1390 1043 1394
rect 1103 1390 1107 1394
rect 1143 1390 1147 1394
rect 1199 1390 1203 1394
rect 1239 1390 1243 1394
rect 1855 1446 1859 1450
rect 1903 1446 1907 1450
rect 1935 1446 1939 1450
rect 1991 1446 1995 1450
rect 2015 1446 2019 1450
rect 2071 1446 2075 1450
rect 2103 1446 2107 1450
rect 2159 1446 2163 1450
rect 2247 1446 2251 1450
rect 2503 1446 2507 1450
rect 1287 1390 1291 1394
rect 1327 1394 1331 1398
rect 1375 1394 1379 1398
rect 1463 1394 1467 1398
rect 1551 1394 1555 1398
rect 1567 1394 1571 1398
rect 1647 1394 1651 1398
rect 1735 1394 1739 1398
rect 1743 1394 1747 1398
rect 1831 1394 1835 1398
rect 1919 1394 1923 1398
rect 2007 1394 2011 1398
rect 2087 1394 2091 1398
rect 2095 1394 2099 1398
rect 2175 1394 2179 1398
rect 2247 1394 2251 1398
rect 2263 1394 2267 1398
rect 2319 1394 2323 1398
rect 2399 1394 2403 1398
rect 2455 1394 2459 1398
rect 2503 1394 2507 1398
rect 687 1322 691 1326
rect 735 1322 739 1326
rect 783 1322 787 1326
rect 823 1322 827 1326
rect 879 1322 883 1326
rect 911 1322 915 1326
rect 215 1262 219 1266
rect 255 1262 259 1266
rect 303 1262 307 1266
rect 383 1262 387 1266
rect 391 1262 395 1266
rect 471 1262 475 1266
rect 495 1262 499 1266
rect 551 1262 555 1266
rect 111 1206 115 1210
rect 135 1206 139 1210
rect 191 1206 195 1210
rect 199 1206 203 1210
rect 271 1206 275 1210
rect 287 1206 291 1210
rect 351 1206 355 1210
rect 375 1206 379 1210
rect 111 1150 115 1154
rect 151 1150 155 1154
rect 183 1150 187 1154
rect 207 1150 211 1154
rect 279 1150 283 1154
rect 287 1150 291 1154
rect 367 1150 371 1154
rect 375 1150 379 1154
rect 431 1206 435 1210
rect 455 1206 459 1210
rect 599 1262 603 1266
rect 623 1262 627 1266
rect 695 1262 699 1266
rect 703 1262 707 1266
rect 1327 1342 1331 1346
rect 1551 1342 1555 1346
rect 1583 1342 1587 1346
rect 1631 1342 1635 1346
rect 1647 1342 1651 1346
rect 1719 1342 1723 1346
rect 1727 1342 1731 1346
rect 1807 1342 1811 1346
rect 1815 1342 1819 1346
rect 1895 1342 1899 1346
rect 1903 1342 1907 1346
rect 975 1322 979 1326
rect 999 1322 1003 1326
rect 1087 1322 1091 1326
rect 1183 1322 1187 1326
rect 1287 1322 1291 1326
rect 1983 1342 1987 1346
rect 1991 1342 1995 1346
rect 2063 1342 2067 1346
rect 2079 1342 2083 1346
rect 2143 1342 2147 1346
rect 2159 1342 2163 1346
rect 2223 1342 2227 1346
rect 2231 1342 2235 1346
rect 2303 1342 2307 1346
rect 1327 1290 1331 1294
rect 1567 1290 1571 1294
rect 767 1262 771 1266
rect 799 1262 803 1266
rect 839 1262 843 1266
rect 895 1262 899 1266
rect 919 1262 923 1266
rect 991 1262 995 1266
rect 1287 1262 1291 1266
rect 1599 1290 1603 1294
rect 1631 1290 1635 1294
rect 1663 1290 1667 1294
rect 1711 1290 1715 1294
rect 1743 1290 1747 1294
rect 1327 1234 1331 1238
rect 511 1206 515 1210
rect 535 1206 539 1210
rect 583 1206 587 1210
rect 607 1206 611 1210
rect 447 1150 451 1154
rect 471 1150 475 1154
rect 1519 1234 1523 1238
rect 1551 1234 1555 1238
rect 1575 1234 1579 1238
rect 1799 1290 1803 1294
rect 1823 1290 1827 1294
rect 1895 1290 1899 1294
rect 1911 1290 1915 1294
rect 1991 1290 1995 1294
rect 1999 1290 2003 1294
rect 2079 1290 2083 1294
rect 2095 1290 2099 1294
rect 2159 1290 2163 1294
rect 2207 1290 2211 1294
rect 2239 1290 2243 1294
rect 1615 1234 1619 1238
rect 1631 1234 1635 1238
rect 1687 1234 1691 1238
rect 1695 1234 1699 1238
rect 647 1206 651 1210
rect 679 1206 683 1210
rect 719 1206 723 1210
rect 751 1206 755 1210
rect 791 1206 795 1210
rect 823 1206 827 1210
rect 863 1206 867 1210
rect 903 1206 907 1210
rect 1287 1206 1291 1210
rect 1743 1234 1747 1238
rect 1783 1234 1787 1238
rect 1799 1234 1803 1238
rect 1855 1234 1859 1238
rect 1879 1234 1883 1238
rect 1911 1234 1915 1238
rect 1967 1234 1971 1238
rect 1975 1234 1979 1238
rect 2031 1234 2035 1238
rect 2383 1342 2387 1346
rect 2439 1342 2443 1346
rect 2503 1342 2507 1346
rect 2319 1290 2323 1294
rect 2079 1234 2083 1238
rect 2103 1234 2107 1238
rect 2183 1234 2187 1238
rect 2191 1234 2195 1238
rect 2271 1234 2275 1238
rect 2303 1234 2307 1238
rect 2367 1234 2371 1238
rect 2399 1290 2403 1294
rect 2455 1290 2459 1294
rect 2439 1234 2443 1238
rect 1327 1178 1331 1182
rect 1535 1178 1539 1182
rect 1567 1178 1571 1182
rect 1591 1178 1595 1182
rect 1631 1178 1635 1182
rect 1647 1178 1651 1182
rect 1703 1178 1707 1182
rect 1759 1178 1763 1182
rect 1791 1178 1795 1182
rect 1815 1178 1819 1182
rect 527 1150 531 1154
rect 567 1150 571 1154
rect 599 1150 603 1154
rect 655 1150 659 1154
rect 663 1150 667 1154
rect 735 1150 739 1154
rect 807 1150 811 1154
rect 879 1150 883 1154
rect 959 1150 963 1154
rect 1039 1150 1043 1154
rect 1287 1150 1291 1154
rect 111 1090 115 1094
rect 167 1090 171 1094
rect 207 1090 211 1094
rect 263 1090 267 1094
rect 279 1090 283 1094
rect 359 1090 363 1094
rect 447 1090 451 1094
rect 455 1090 459 1094
rect 543 1090 547 1094
rect 551 1090 555 1094
rect 1327 1126 1331 1130
rect 1383 1126 1387 1130
rect 1447 1126 1451 1130
rect 1519 1126 1523 1130
rect 1551 1126 1555 1130
rect 1591 1126 1595 1130
rect 1615 1126 1619 1130
rect 1671 1126 1675 1130
rect 1687 1126 1691 1130
rect 1751 1126 1755 1130
rect 1775 1126 1779 1130
rect 639 1090 643 1094
rect 719 1090 723 1094
rect 727 1090 731 1094
rect 791 1090 795 1094
rect 815 1090 819 1094
rect 863 1090 867 1094
rect 895 1090 899 1094
rect 943 1090 947 1094
rect 975 1090 979 1094
rect 1023 1090 1027 1094
rect 1055 1090 1059 1094
rect 111 1030 115 1034
rect 223 1030 227 1034
rect 295 1030 299 1034
rect 375 1030 379 1034
rect 383 1030 387 1034
rect 463 1030 467 1034
rect 479 1030 483 1034
rect 559 1030 563 1034
rect 575 1030 579 1034
rect 1871 1178 1875 1182
rect 1903 1178 1907 1182
rect 1927 1178 1931 1182
rect 1983 1178 1987 1182
rect 2031 1178 2035 1182
rect 2047 1178 2051 1182
rect 2119 1178 2123 1182
rect 2175 1178 2179 1182
rect 2199 1178 2203 1182
rect 2287 1178 2291 1182
rect 2327 1178 2331 1182
rect 2383 1178 2387 1182
rect 2455 1178 2459 1182
rect 2503 1290 2507 1294
rect 2503 1234 2507 1238
rect 2503 1178 2507 1182
rect 1831 1126 1835 1130
rect 1887 1126 1891 1130
rect 1911 1126 1915 1130
rect 1143 1090 1147 1094
rect 1287 1090 1291 1094
rect 1983 1126 1987 1130
rect 2015 1126 2019 1130
rect 2055 1126 2059 1130
rect 2135 1126 2139 1130
rect 2159 1126 2163 1130
rect 2215 1126 2219 1130
rect 2311 1126 2315 1130
rect 2439 1126 2443 1130
rect 1327 1066 1331 1070
rect 1367 1066 1371 1070
rect 1399 1066 1403 1070
rect 1455 1066 1459 1070
rect 1463 1066 1467 1070
rect 1535 1066 1539 1070
rect 1575 1066 1579 1070
rect 1607 1066 1611 1070
rect 1687 1066 1691 1070
rect 1695 1066 1699 1070
rect 1767 1066 1771 1070
rect 1815 1066 1819 1070
rect 655 1030 659 1034
rect 671 1030 675 1034
rect 743 1030 747 1034
rect 767 1030 771 1034
rect 831 1030 835 1034
rect 855 1030 859 1034
rect 911 1030 915 1034
rect 943 1030 947 1034
rect 991 1030 995 1034
rect 1023 1030 1027 1034
rect 1071 1030 1075 1034
rect 1103 1030 1107 1034
rect 1159 1030 1163 1034
rect 1183 1030 1187 1034
rect 1239 1030 1243 1034
rect 1287 1030 1291 1034
rect 111 978 115 982
rect 271 978 275 982
rect 279 978 283 982
rect 359 978 363 982
rect 367 978 371 982
rect 455 978 459 982
rect 463 978 467 982
rect 551 978 555 982
rect 559 978 563 982
rect 655 978 659 982
rect 751 978 755 982
rect 839 978 843 982
rect 927 978 931 982
rect 1007 978 1011 982
rect 1087 978 1091 982
rect 1167 978 1171 982
rect 111 918 115 922
rect 271 918 275 922
rect 287 918 291 922
rect 343 918 347 922
rect 375 918 379 922
rect 423 918 427 922
rect 111 862 115 866
rect 247 862 251 866
rect 255 862 259 866
rect 1327 1010 1331 1014
rect 1351 1010 1355 1014
rect 1439 1010 1443 1014
rect 1511 1010 1515 1014
rect 1559 1010 1563 1014
rect 1679 1010 1683 1014
rect 1223 978 1227 982
rect 1847 1066 1851 1070
rect 1927 1066 1931 1070
rect 1999 1066 2003 1070
rect 2039 1066 2043 1070
rect 2071 1066 2075 1070
rect 2151 1066 2155 1070
rect 2231 1066 2235 1070
rect 2255 1066 2259 1070
rect 2367 1066 2371 1070
rect 2455 1066 2459 1070
rect 1799 1010 1803 1014
rect 1823 1010 1827 1014
rect 1911 1010 1915 1014
rect 1951 1010 1955 1014
rect 2023 1010 2027 1014
rect 2071 1010 2075 1014
rect 2135 1010 2139 1014
rect 2175 1010 2179 1014
rect 2239 1010 2243 1014
rect 2271 1010 2275 1014
rect 2351 1010 2355 1014
rect 2367 1010 2371 1014
rect 1287 978 1291 982
rect 471 918 475 922
rect 519 918 523 922
rect 567 918 571 922
rect 615 918 619 922
rect 671 918 675 922
rect 711 918 715 922
rect 767 918 771 922
rect 807 918 811 922
rect 855 918 859 922
rect 903 918 907 922
rect 943 918 947 922
rect 991 918 995 922
rect 1023 918 1027 922
rect 1087 918 1091 922
rect 1103 918 1107 922
rect 1183 918 1187 922
rect 311 862 315 866
rect 327 862 331 866
rect 375 862 379 866
rect 407 862 411 866
rect 439 862 443 866
rect 503 862 507 866
rect 567 862 571 866
rect 599 862 603 866
rect 631 862 635 866
rect 695 862 699 866
rect 111 806 115 810
rect 215 806 219 810
rect 263 806 267 810
rect 303 806 307 810
rect 111 754 115 758
rect 135 754 139 758
rect 327 806 331 810
rect 391 806 395 810
rect 455 806 459 810
rect 479 806 483 810
rect 519 806 523 810
rect 559 806 563 810
rect 583 806 587 810
rect 631 806 635 810
rect 647 806 651 810
rect 759 862 763 866
rect 791 862 795 866
rect 831 862 835 866
rect 887 862 891 866
rect 903 862 907 866
rect 1327 946 1331 950
rect 1367 946 1371 950
rect 1823 968 1827 972
rect 2439 1010 2443 1014
rect 2375 968 2379 972
rect 1423 946 1427 950
rect 1503 946 1507 950
rect 1527 946 1531 950
rect 1607 946 1611 950
rect 1695 946 1699 950
rect 1719 946 1723 950
rect 1831 946 1835 950
rect 1839 946 1843 950
rect 1935 946 1939 950
rect 1967 946 1971 950
rect 2031 946 2035 950
rect 2087 946 2091 950
rect 2127 946 2131 950
rect 2191 946 2195 950
rect 2215 946 2219 950
rect 2287 946 2291 950
rect 2295 946 2299 950
rect 2375 946 2379 950
rect 2383 946 2387 950
rect 1239 918 1243 922
rect 1287 918 1291 922
rect 1327 890 1331 894
rect 1351 890 1355 894
rect 1407 890 1411 894
rect 1431 890 1435 894
rect 975 862 979 866
rect 1071 862 1075 866
rect 1167 862 1171 866
rect 1287 862 1291 866
rect 1487 890 1491 894
rect 1551 890 1555 894
rect 1591 890 1595 894
rect 1623 890 1627 894
rect 1703 890 1707 894
rect 1791 890 1795 894
rect 1815 890 1819 894
rect 1895 890 1899 894
rect 1919 890 1923 894
rect 2015 890 2019 894
rect 2111 890 2115 894
rect 2143 890 2147 894
rect 1327 834 1331 838
rect 1447 834 1451 838
rect 1503 834 1507 838
rect 1567 834 1571 838
rect 1591 834 1595 838
rect 1639 834 1643 838
rect 1647 834 1651 838
rect 1703 834 1707 838
rect 1719 834 1723 838
rect 1767 834 1771 838
rect 1807 834 1811 838
rect 1847 834 1851 838
rect 1911 834 1915 838
rect 703 806 707 810
rect 711 806 715 810
rect 767 806 771 810
rect 775 806 779 810
rect 831 806 835 810
rect 847 806 851 810
rect 895 806 899 810
rect 919 806 923 810
rect 967 806 971 810
rect 1039 806 1043 810
rect 1287 806 1291 810
rect 2199 890 2203 894
rect 2279 890 2283 894
rect 2359 890 2363 894
rect 2423 890 2427 894
rect 2439 890 2443 894
rect 2455 946 2459 950
rect 2503 1126 2507 1130
rect 2503 1066 2507 1070
rect 2503 1010 2507 1014
rect 2503 946 2507 950
rect 1927 834 1931 838
rect 2015 834 2019 838
rect 2031 834 2035 838
rect 2103 834 2107 838
rect 2159 834 2163 838
rect 2191 834 2195 838
rect 2287 834 2291 838
rect 2295 834 2299 838
rect 2383 834 2387 838
rect 199 754 203 758
rect 255 754 259 758
rect 287 754 291 758
rect 375 754 379 758
rect 391 754 395 758
rect 463 754 467 758
rect 519 754 523 758
rect 543 754 547 758
rect 615 754 619 758
rect 647 754 651 758
rect 687 754 691 758
rect 751 754 755 758
rect 775 754 779 758
rect 111 702 115 706
rect 151 702 155 706
rect 207 702 211 706
rect 271 702 275 706
rect 295 702 299 706
rect 391 702 395 706
rect 407 702 411 706
rect 111 646 115 650
rect 135 646 139 650
rect 151 646 155 650
rect 191 646 195 650
rect 263 646 267 650
rect 279 646 283 650
rect 503 702 507 706
rect 535 702 539 706
rect 623 702 627 706
rect 663 702 667 706
rect 815 754 819 758
rect 879 754 883 758
rect 903 754 907 758
rect 951 754 955 758
rect 1023 754 1027 758
rect 1039 754 1043 758
rect 1327 778 1331 782
rect 1567 778 1571 782
rect 1575 778 1579 782
rect 1623 778 1627 782
rect 1631 778 1635 782
rect 1687 778 1691 782
rect 1751 778 1755 782
rect 1759 778 1763 782
rect 1831 778 1835 782
rect 1287 754 1291 758
rect 1327 726 1331 730
rect 1367 726 1371 730
rect 1431 726 1435 730
rect 1527 726 1531 730
rect 1583 726 1587 730
rect 743 702 747 706
rect 791 702 795 706
rect 871 702 875 706
rect 919 702 923 706
rect 999 702 1003 706
rect 1055 702 1059 706
rect 1127 702 1131 706
rect 1239 702 1243 706
rect 1287 702 1291 706
rect 1631 726 1635 730
rect 1639 726 1643 730
rect 367 646 371 650
rect 375 646 379 650
rect 463 646 467 650
rect 487 646 491 650
rect 559 646 563 650
rect 607 646 611 650
rect 111 594 115 598
rect 151 594 155 598
rect 167 594 171 598
rect 239 594 243 598
rect 279 594 283 598
rect 335 594 339 598
rect 383 594 387 598
rect 111 534 115 538
rect 135 534 139 538
rect 143 534 147 538
rect 223 534 227 538
rect 239 534 243 538
rect 655 646 659 650
rect 727 646 731 650
rect 751 646 755 650
rect 847 646 851 650
rect 855 646 859 650
rect 943 646 947 650
rect 1703 726 1707 730
rect 1911 778 1915 782
rect 1919 778 1923 782
rect 1999 778 2003 782
rect 2015 778 2019 782
rect 2087 778 2091 782
rect 2119 778 2123 782
rect 2175 778 2179 782
rect 2231 778 2235 782
rect 2271 778 2275 782
rect 2343 778 2347 782
rect 2367 778 2371 782
rect 2439 834 2443 838
rect 2455 834 2459 838
rect 2503 890 2507 894
rect 2503 834 2507 838
rect 2439 778 2443 782
rect 1735 726 1739 730
rect 1775 726 1779 730
rect 1839 726 1843 730
rect 1847 726 1851 730
rect 1935 726 1939 730
rect 1943 726 1947 730
rect 2031 726 2035 730
rect 2047 726 2051 730
rect 2135 726 2139 730
rect 1327 662 1331 666
rect 983 646 987 650
rect 1039 646 1043 650
rect 1111 646 1115 650
rect 1143 646 1147 650
rect 1223 646 1227 650
rect 1287 646 1291 650
rect 431 594 435 598
rect 479 594 483 598
rect 535 594 539 598
rect 575 594 579 598
rect 631 594 635 598
rect 671 594 675 598
rect 727 594 731 598
rect 767 594 771 598
rect 823 594 827 598
rect 319 534 323 538
rect 335 534 339 538
rect 415 534 419 538
rect 431 534 435 538
rect 519 534 523 538
rect 527 534 531 538
rect 615 534 619 538
rect 623 534 627 538
rect 111 478 115 482
rect 151 478 155 482
rect 159 478 163 482
rect 207 478 211 482
rect 255 478 259 482
rect 287 478 291 482
rect 351 478 355 482
rect 375 478 379 482
rect 447 478 451 482
rect 111 426 115 430
rect 135 426 139 430
rect 191 426 195 430
rect 271 426 275 430
rect 279 426 283 430
rect 711 534 715 538
rect 863 594 867 598
rect 911 594 915 598
rect 959 594 963 598
rect 999 594 1003 598
rect 1055 594 1059 598
rect 1087 594 1091 598
rect 1159 594 1163 598
rect 1351 662 1355 666
rect 1415 662 1419 666
rect 1511 662 1515 666
rect 1607 662 1611 666
rect 1615 662 1619 666
rect 1711 662 1715 666
rect 1719 662 1723 666
rect 1823 662 1827 666
rect 2151 726 2155 730
rect 2247 726 2251 730
rect 2255 726 2259 730
rect 2359 726 2363 730
rect 2367 726 2371 730
rect 2455 726 2459 730
rect 2503 778 2507 782
rect 2503 726 2507 730
rect 1927 662 1931 666
rect 1935 662 1939 666
rect 2031 662 2035 666
rect 2055 662 2059 666
rect 2135 662 2139 666
rect 2183 662 2187 666
rect 2239 662 2243 666
rect 2319 662 2323 666
rect 2351 662 2355 666
rect 2439 662 2443 666
rect 1327 610 1331 614
rect 1367 610 1371 614
rect 1383 610 1387 614
rect 1431 610 1435 614
rect 1463 610 1467 614
rect 1527 610 1531 614
rect 1551 610 1555 614
rect 1623 610 1627 614
rect 1647 610 1651 614
rect 1727 610 1731 614
rect 1743 610 1747 614
rect 1183 594 1187 598
rect 1239 594 1243 598
rect 1287 594 1291 598
rect 791 534 795 538
rect 807 534 811 538
rect 871 534 875 538
rect 895 534 899 538
rect 463 478 467 482
rect 543 478 547 482
rect 559 478 563 482
rect 639 478 643 482
rect 655 478 659 482
rect 727 478 731 482
rect 751 478 755 482
rect 807 478 811 482
rect 359 426 363 430
rect 383 426 387 430
rect 111 370 115 374
rect 151 370 155 374
rect 447 426 451 430
rect 495 426 499 430
rect 543 426 547 430
rect 607 426 611 430
rect 639 426 643 430
rect 719 426 723 430
rect 735 426 739 430
rect 1327 558 1331 562
rect 1367 558 1371 562
rect 1375 558 1379 562
rect 951 534 955 538
rect 983 534 987 538
rect 1031 534 1035 538
rect 1071 534 1075 538
rect 1167 534 1171 538
rect 1287 534 1291 538
rect 1447 558 1451 562
rect 1455 558 1459 562
rect 1535 558 1539 562
rect 1551 558 1555 562
rect 1839 610 1843 614
rect 1847 610 1851 614
rect 1951 610 1955 614
rect 1959 610 1963 614
rect 1631 558 1635 562
rect 1647 558 1651 562
rect 1727 558 1731 562
rect 1751 558 1755 562
rect 1831 558 1835 562
rect 1855 558 1859 562
rect 2071 610 2075 614
rect 2079 610 2083 614
rect 2199 610 2203 614
rect 2207 610 2211 614
rect 2335 610 2339 614
rect 2343 610 2347 614
rect 2455 610 2459 614
rect 2503 662 2507 666
rect 2503 610 2507 614
rect 1943 558 1947 562
rect 1959 558 1963 562
rect 2055 558 2059 562
rect 2063 558 2067 562
rect 2151 558 2155 562
rect 2191 558 2195 562
rect 1327 502 1331 506
rect 1367 502 1371 506
rect 1391 502 1395 506
rect 1455 502 1459 506
rect 1471 502 1475 506
rect 847 478 851 482
rect 887 478 891 482
rect 951 478 955 482
rect 967 478 971 482
rect 1047 478 1051 482
rect 1055 478 1059 482
rect 1159 478 1163 482
rect 1239 478 1243 482
rect 1287 478 1291 482
rect 1567 502 1571 506
rect 1575 502 1579 506
rect 1663 502 1667 506
rect 1695 502 1699 506
rect 1767 502 1771 506
rect 1807 502 1811 506
rect 831 426 835 430
rect 935 426 939 430
rect 1039 426 1043 430
rect 1143 426 1147 430
rect 207 370 211 374
rect 231 370 235 374
rect 295 370 299 374
rect 335 370 339 374
rect 399 370 403 374
rect 439 370 443 374
rect 511 370 515 374
rect 543 370 547 374
rect 623 370 627 374
rect 647 370 651 374
rect 735 370 739 374
rect 751 370 755 374
rect 111 314 115 318
rect 135 314 139 318
rect 215 314 219 318
rect 319 314 323 318
rect 423 314 427 318
rect 527 314 531 318
rect 535 314 539 318
rect 111 262 115 266
rect 151 262 155 266
rect 223 262 227 266
rect 231 262 235 266
rect 319 262 323 266
rect 335 262 339 266
rect 111 206 115 210
rect 135 206 139 210
rect 183 206 187 210
rect 207 206 211 210
rect 279 206 283 210
rect 303 206 307 210
rect 631 314 635 318
rect 639 314 643 318
rect 847 370 851 374
rect 935 370 939 374
rect 951 370 955 374
rect 1015 370 1019 374
rect 1055 370 1059 374
rect 1327 438 1331 442
rect 1351 438 1355 442
rect 1439 438 1443 442
rect 1559 438 1563 442
rect 1583 438 1587 442
rect 1223 426 1227 430
rect 1287 426 1291 430
rect 1871 502 1875 506
rect 1919 502 1923 506
rect 2255 558 2259 562
rect 2327 558 2331 562
rect 2359 558 2363 562
rect 2439 558 2443 562
rect 1975 502 1979 506
rect 2023 502 2027 506
rect 2071 502 2075 506
rect 2119 502 2123 506
rect 2167 502 2171 506
rect 2207 502 2211 506
rect 2271 502 2275 506
rect 1639 438 1643 442
rect 1679 438 1683 442
rect 1695 438 1699 442
rect 1759 438 1763 442
rect 1791 438 1795 442
rect 1831 438 1835 442
rect 1903 438 1907 442
rect 1911 438 1915 442
rect 1327 382 1331 386
rect 1599 382 1603 386
rect 1655 382 1659 386
rect 1679 382 1683 386
rect 1711 382 1715 386
rect 1735 382 1739 386
rect 1775 382 1779 386
rect 1799 382 1803 386
rect 1847 382 1851 386
rect 1871 382 1875 386
rect 1095 370 1099 374
rect 1159 370 1163 374
rect 1175 370 1179 374
rect 1239 370 1243 374
rect 1287 370 1291 374
rect 735 314 739 318
rect 743 314 747 318
rect 831 314 835 318
rect 847 314 851 318
rect 919 314 923 318
rect 943 314 947 318
rect 999 314 1003 318
rect 1039 314 1043 318
rect 1079 314 1083 318
rect 1143 314 1147 318
rect 1159 314 1163 318
rect 1223 314 1227 318
rect 423 262 427 266
rect 439 262 443 266
rect 535 262 539 266
rect 551 262 555 266
rect 647 262 651 266
rect 655 262 659 266
rect 759 262 763 266
rect 863 262 867 266
rect 871 262 875 266
rect 383 206 387 210
rect 407 206 411 210
rect 487 206 491 210
rect 519 206 523 210
rect 591 206 595 210
rect 631 206 635 210
rect 111 146 115 150
rect 151 146 155 150
rect 199 146 203 150
rect 207 146 211 150
rect 263 146 267 150
rect 295 146 299 150
rect 319 146 323 150
rect 375 146 379 150
rect 399 146 403 150
rect 431 146 435 150
rect 695 206 699 210
rect 959 262 963 266
rect 983 262 987 266
rect 1055 262 1059 266
rect 1103 262 1107 266
rect 1159 262 1163 266
rect 1327 322 1331 326
rect 1351 322 1355 326
rect 1455 322 1459 326
rect 1583 322 1587 326
rect 1287 314 1291 318
rect 1663 322 1667 326
rect 1711 322 1715 326
rect 1719 322 1723 326
rect 1783 322 1787 326
rect 1839 322 1843 326
rect 1855 322 1859 326
rect 1927 382 1931 386
rect 1943 382 1947 386
rect 2295 502 2299 506
rect 2375 502 2379 506
rect 2383 502 2387 506
rect 2503 558 2507 562
rect 2455 502 2459 506
rect 1991 438 1995 442
rect 2007 438 2011 442
rect 2079 438 2083 442
rect 2103 438 2107 442
rect 2007 382 2011 386
rect 2023 382 2027 386
rect 2095 382 2099 386
rect 2175 438 2179 442
rect 2191 438 2195 442
rect 2271 438 2275 442
rect 2279 438 2283 442
rect 2367 438 2371 442
rect 2111 382 2115 386
rect 2191 382 2195 386
rect 2199 382 2203 386
rect 2287 382 2291 386
rect 2375 382 2379 386
rect 2383 382 2387 386
rect 2439 438 2443 442
rect 2455 382 2459 386
rect 1927 322 1931 326
rect 1951 322 1955 326
rect 2007 322 2011 326
rect 2063 322 2067 326
rect 2095 322 2099 326
rect 2167 322 2171 326
rect 2183 322 2187 326
rect 1223 262 1227 266
rect 1239 262 1243 266
rect 1287 262 1291 266
rect 1327 262 1331 266
rect 1367 262 1371 266
rect 1447 262 1451 266
rect 1471 262 1475 266
rect 1551 262 1555 266
rect 1599 262 1603 266
rect 1655 262 1659 266
rect 1727 262 1731 266
rect 1759 262 1763 266
rect 743 206 747 210
rect 799 206 803 210
rect 855 206 859 210
rect 895 206 899 210
rect 967 206 971 210
rect 999 206 1003 210
rect 1087 206 1091 210
rect 1103 206 1107 210
rect 1207 206 1211 210
rect 1287 206 1291 210
rect 1327 206 1331 210
rect 1351 206 1355 210
rect 1407 206 1411 210
rect 1431 206 1435 210
rect 487 146 491 150
rect 503 146 507 150
rect 543 146 547 150
rect 599 146 603 150
rect 607 146 611 150
rect 655 146 659 150
rect 711 146 715 150
rect 767 146 771 150
rect 815 146 819 150
rect 831 146 835 150
rect 895 146 899 150
rect 911 146 915 150
rect 959 146 963 150
rect 1015 146 1019 150
rect 1023 146 1027 150
rect 1087 146 1091 150
rect 1119 146 1123 150
rect 1151 146 1155 150
rect 1287 146 1291 150
rect 1327 134 1331 138
rect 1367 134 1371 138
rect 1471 206 1475 210
rect 1535 206 1539 210
rect 1551 206 1555 210
rect 1855 262 1859 266
rect 1863 262 1867 266
rect 1967 262 1971 266
rect 1639 206 1643 210
rect 1719 206 1723 210
rect 1743 206 1747 210
rect 1807 206 1811 210
rect 2071 262 2075 266
rect 2079 262 2083 266
rect 2263 322 2267 326
rect 2271 322 2275 326
rect 2359 322 2363 326
rect 2175 262 2179 266
rect 2183 262 2187 266
rect 2271 262 2275 266
rect 2279 262 2283 266
rect 2439 322 2443 326
rect 2503 502 2507 506
rect 2503 438 2507 442
rect 2503 382 2507 386
rect 2503 322 2507 326
rect 2375 262 2379 266
rect 2455 262 2459 266
rect 2503 262 2507 266
rect 1847 206 1851 210
rect 1895 206 1899 210
rect 1951 206 1955 210
rect 1991 206 1995 210
rect 2055 206 2059 210
rect 2103 206 2107 210
rect 2159 206 2163 210
rect 2215 206 2219 210
rect 2255 206 2259 210
rect 1423 134 1427 138
rect 1479 134 1483 138
rect 1487 134 1491 138
rect 1535 134 1539 138
rect 1567 134 1571 138
rect 1591 134 1595 138
rect 1647 134 1651 138
rect 1655 134 1659 138
rect 1703 134 1707 138
rect 1735 134 1739 138
rect 1759 134 1763 138
rect 1823 134 1827 138
rect 1879 134 1883 138
rect 1911 134 1915 138
rect 1943 134 1947 138
rect 2007 134 2011 138
rect 2071 134 2075 138
rect 2119 134 2123 138
rect 2335 206 2339 210
rect 2359 206 2363 210
rect 2439 206 2443 210
rect 2143 134 2147 138
rect 2223 134 2227 138
rect 2231 134 2235 138
rect 2303 134 2307 138
rect 2351 134 2355 138
rect 2391 134 2395 138
rect 2455 134 2459 138
rect 2503 206 2507 210
rect 2503 134 2507 138
rect 111 94 115 98
rect 135 94 139 98
rect 191 94 195 98
rect 247 94 251 98
rect 303 94 307 98
rect 359 94 363 98
rect 415 94 419 98
rect 471 94 475 98
rect 527 94 531 98
rect 583 94 587 98
rect 639 94 643 98
rect 695 94 699 98
rect 751 94 755 98
rect 815 94 819 98
rect 879 94 883 98
rect 943 94 947 98
rect 1007 94 1011 98
rect 1071 94 1075 98
rect 1135 94 1139 98
rect 1287 94 1291 98
rect 1327 82 1331 86
rect 1351 82 1355 86
rect 1407 82 1411 86
rect 1463 82 1467 86
rect 1519 82 1523 86
rect 1575 82 1579 86
rect 1631 82 1635 86
rect 1687 82 1691 86
rect 1743 82 1747 86
rect 1807 82 1811 86
rect 1863 82 1867 86
rect 1927 82 1931 86
rect 1991 82 1995 86
rect 2055 82 2059 86
rect 2127 82 2131 86
rect 2207 82 2211 86
rect 2287 82 2291 86
rect 2375 82 2379 86
rect 2439 82 2443 86
rect 2503 82 2507 86
<< m4 >>
rect 84 2577 85 2583
rect 91 2582 1299 2583
rect 91 2578 111 2582
rect 115 2578 135 2582
rect 139 2578 191 2582
rect 195 2578 247 2582
rect 251 2578 303 2582
rect 307 2578 359 2582
rect 363 2578 1287 2582
rect 1291 2578 1299 2582
rect 91 2577 1299 2578
rect 1305 2577 1306 2583
rect 1298 2557 1299 2563
rect 1305 2562 2527 2563
rect 1305 2558 1327 2562
rect 1331 2558 1495 2562
rect 1499 2558 1551 2562
rect 1555 2558 1607 2562
rect 1611 2558 1663 2562
rect 1667 2558 1719 2562
rect 1723 2558 1775 2562
rect 1779 2558 1831 2562
rect 1835 2558 1887 2562
rect 1891 2558 1943 2562
rect 1947 2558 1999 2562
rect 2003 2558 2055 2562
rect 2059 2558 2111 2562
rect 2115 2558 2167 2562
rect 2171 2558 2503 2562
rect 2507 2558 2527 2562
rect 1305 2557 2527 2558
rect 2533 2557 2534 2563
rect 96 2525 97 2531
rect 103 2530 1311 2531
rect 103 2526 111 2530
rect 115 2526 151 2530
rect 155 2526 207 2530
rect 211 2526 223 2530
rect 227 2526 263 2530
rect 267 2526 279 2530
rect 283 2526 319 2530
rect 323 2526 343 2530
rect 347 2526 375 2530
rect 379 2526 415 2530
rect 419 2526 487 2530
rect 491 2526 551 2530
rect 555 2526 615 2530
rect 619 2526 679 2530
rect 683 2526 743 2530
rect 747 2526 807 2530
rect 811 2526 871 2530
rect 875 2526 935 2530
rect 939 2526 999 2530
rect 1003 2526 1063 2530
rect 1067 2526 1287 2530
rect 1291 2526 1311 2530
rect 103 2525 1311 2526
rect 1317 2525 1318 2531
rect 1910 2524 1916 2525
rect 2190 2524 2196 2525
rect 1910 2520 1911 2524
rect 1915 2520 2191 2524
rect 2195 2520 2196 2524
rect 1910 2519 1916 2520
rect 2190 2519 2196 2520
rect 1310 2505 1311 2511
rect 1317 2510 2539 2511
rect 1317 2506 1327 2510
rect 1331 2506 1511 2510
rect 1515 2506 1543 2510
rect 1547 2506 1567 2510
rect 1571 2506 1607 2510
rect 1611 2506 1623 2510
rect 1627 2506 1679 2510
rect 1683 2506 1735 2510
rect 1739 2506 1751 2510
rect 1755 2506 1791 2510
rect 1795 2506 1823 2510
rect 1827 2506 1847 2510
rect 1851 2506 1895 2510
rect 1899 2506 1903 2510
rect 1907 2506 1959 2510
rect 1963 2506 1967 2510
rect 1971 2506 2015 2510
rect 2019 2506 2039 2510
rect 2043 2506 2071 2510
rect 2075 2506 2111 2510
rect 2115 2506 2127 2510
rect 2131 2506 2183 2510
rect 2187 2506 2503 2510
rect 2507 2506 2539 2510
rect 1317 2505 2539 2506
rect 2545 2505 2546 2511
rect 1526 2492 1532 2493
rect 1842 2492 1848 2493
rect 1526 2488 1527 2492
rect 1531 2488 1843 2492
rect 1847 2488 1848 2492
rect 1526 2487 1532 2488
rect 1842 2487 1848 2488
rect 84 2465 85 2471
rect 91 2470 1299 2471
rect 91 2466 111 2470
rect 115 2466 167 2470
rect 171 2466 207 2470
rect 211 2466 223 2470
rect 227 2466 263 2470
rect 267 2466 279 2470
rect 283 2466 327 2470
rect 331 2466 335 2470
rect 339 2466 391 2470
rect 395 2466 399 2470
rect 403 2466 447 2470
rect 451 2466 471 2470
rect 475 2466 503 2470
rect 507 2466 535 2470
rect 539 2466 559 2470
rect 563 2466 599 2470
rect 603 2466 615 2470
rect 619 2466 663 2470
rect 667 2466 671 2470
rect 675 2466 727 2470
rect 731 2466 783 2470
rect 787 2466 791 2470
rect 795 2466 839 2470
rect 843 2466 855 2470
rect 859 2466 895 2470
rect 899 2466 919 2470
rect 923 2466 951 2470
rect 955 2466 983 2470
rect 987 2466 1007 2470
rect 1011 2466 1047 2470
rect 1051 2466 1063 2470
rect 1067 2466 1287 2470
rect 1291 2466 1299 2470
rect 91 2465 1299 2466
rect 1305 2465 1306 2471
rect 166 2452 172 2453
rect 494 2452 500 2453
rect 166 2448 167 2452
rect 171 2448 495 2452
rect 499 2448 500 2452
rect 166 2447 172 2448
rect 494 2447 500 2448
rect 566 2452 572 2453
rect 874 2452 880 2453
rect 566 2448 567 2452
rect 571 2448 875 2452
rect 879 2448 880 2452
rect 1298 2449 1299 2455
rect 1305 2454 2527 2455
rect 1305 2450 1327 2454
rect 1331 2450 1527 2454
rect 1531 2450 1543 2454
rect 1547 2450 1591 2454
rect 1595 2450 1607 2454
rect 1611 2450 1663 2454
rect 1667 2450 1671 2454
rect 1675 2450 1735 2454
rect 1739 2450 1743 2454
rect 1747 2450 1807 2454
rect 1811 2450 1815 2454
rect 1819 2450 1879 2454
rect 1883 2450 1951 2454
rect 1955 2450 2023 2454
rect 2027 2450 2095 2454
rect 2099 2450 2167 2454
rect 2171 2450 2503 2454
rect 2507 2450 2527 2454
rect 1305 2449 2527 2450
rect 2533 2449 2534 2455
rect 566 2447 572 2448
rect 874 2447 880 2448
rect 96 2401 97 2407
rect 103 2406 1311 2407
rect 103 2402 111 2406
rect 115 2402 183 2406
rect 187 2402 239 2406
rect 243 2402 295 2406
rect 299 2402 351 2406
rect 355 2402 407 2406
rect 411 2402 463 2406
rect 467 2402 519 2406
rect 523 2402 575 2406
rect 579 2402 631 2406
rect 635 2402 687 2406
rect 691 2402 743 2406
rect 747 2402 799 2406
rect 803 2402 855 2406
rect 859 2402 911 2406
rect 915 2402 967 2406
rect 971 2402 1023 2406
rect 1027 2402 1079 2406
rect 1083 2402 1287 2406
rect 1291 2402 1311 2406
rect 103 2401 1311 2402
rect 1317 2401 1318 2407
rect 1310 2399 1318 2401
rect 1310 2393 1311 2399
rect 1317 2398 2539 2399
rect 1317 2394 1327 2398
rect 1331 2394 1559 2398
rect 1563 2394 1567 2398
rect 1571 2394 1623 2398
rect 1627 2394 1679 2398
rect 1683 2394 1687 2398
rect 1691 2394 1735 2398
rect 1739 2394 1759 2398
rect 1763 2394 1791 2398
rect 1795 2394 1831 2398
rect 1835 2394 1855 2398
rect 1859 2394 1895 2398
rect 1899 2394 1919 2398
rect 1923 2394 1967 2398
rect 1971 2394 1983 2398
rect 1987 2394 2039 2398
rect 2043 2394 2047 2398
rect 2051 2394 2111 2398
rect 2115 2394 2183 2398
rect 2187 2394 2503 2398
rect 2507 2394 2539 2398
rect 1317 2393 2539 2394
rect 2545 2393 2546 2399
rect 84 2341 85 2347
rect 91 2346 1299 2347
rect 91 2342 111 2346
rect 115 2342 319 2346
rect 323 2342 391 2346
rect 395 2342 463 2346
rect 467 2342 503 2346
rect 507 2342 535 2346
rect 539 2342 559 2346
rect 563 2342 607 2346
rect 611 2342 615 2346
rect 619 2342 671 2346
rect 675 2342 679 2346
rect 683 2342 743 2346
rect 747 2342 807 2346
rect 811 2342 863 2346
rect 867 2342 927 2346
rect 931 2342 991 2346
rect 995 2342 1055 2346
rect 1059 2342 1111 2346
rect 1115 2342 1167 2346
rect 1171 2342 1223 2346
rect 1227 2342 1287 2346
rect 1291 2342 1299 2346
rect 91 2341 1299 2342
rect 1305 2341 1306 2347
rect 1298 2339 1306 2341
rect 1298 2333 1299 2339
rect 1305 2338 2527 2339
rect 1305 2334 1327 2338
rect 1331 2334 1471 2338
rect 1475 2334 1535 2338
rect 1539 2334 1551 2338
rect 1555 2334 1607 2338
rect 1611 2334 1663 2338
rect 1667 2334 1687 2338
rect 1691 2334 1719 2338
rect 1723 2334 1759 2338
rect 1763 2334 1775 2338
rect 1779 2334 1831 2338
rect 1835 2334 1839 2338
rect 1843 2334 1903 2338
rect 1907 2334 1967 2338
rect 1971 2334 1983 2338
rect 1987 2334 2031 2338
rect 2035 2334 2063 2338
rect 2067 2334 2095 2338
rect 2099 2334 2143 2338
rect 2147 2334 2503 2338
rect 2507 2334 2527 2338
rect 1305 2333 2527 2334
rect 2533 2333 2534 2339
rect 96 2281 97 2287
rect 103 2286 1311 2287
rect 103 2282 111 2286
rect 115 2282 175 2286
rect 179 2282 271 2286
rect 275 2282 335 2286
rect 339 2282 375 2286
rect 379 2282 407 2286
rect 411 2282 479 2286
rect 483 2282 551 2286
rect 555 2282 591 2286
rect 595 2282 623 2286
rect 627 2282 695 2286
rect 699 2282 703 2286
rect 707 2282 759 2286
rect 763 2282 807 2286
rect 811 2282 823 2286
rect 827 2282 879 2286
rect 883 2282 911 2286
rect 915 2282 943 2286
rect 947 2282 1007 2286
rect 1011 2282 1015 2286
rect 1019 2282 1071 2286
rect 1075 2282 1127 2286
rect 1131 2282 1183 2286
rect 1187 2282 1239 2286
rect 1243 2282 1287 2286
rect 1291 2282 1311 2286
rect 103 2281 1311 2282
rect 1317 2286 2546 2287
rect 1317 2282 1327 2286
rect 1331 2282 1383 2286
rect 1387 2282 1479 2286
rect 1483 2282 1487 2286
rect 1491 2282 1551 2286
rect 1555 2282 1583 2286
rect 1587 2282 1623 2286
rect 1627 2282 1687 2286
rect 1691 2282 1703 2286
rect 1707 2282 1775 2286
rect 1779 2282 1791 2286
rect 1795 2282 1847 2286
rect 1851 2282 1903 2286
rect 1907 2282 1919 2286
rect 1923 2282 1999 2286
rect 2003 2282 2015 2286
rect 2019 2282 2079 2286
rect 2083 2282 2127 2286
rect 2131 2282 2159 2286
rect 2163 2282 2239 2286
rect 2243 2282 2503 2286
rect 2507 2282 2546 2286
rect 1317 2281 2546 2282
rect 84 2229 85 2235
rect 91 2234 1299 2235
rect 91 2230 111 2234
rect 115 2230 143 2234
rect 147 2230 159 2234
rect 163 2230 231 2234
rect 235 2230 255 2234
rect 259 2230 319 2234
rect 323 2230 359 2234
rect 363 2230 415 2234
rect 419 2230 463 2234
rect 467 2230 519 2234
rect 523 2230 575 2234
rect 579 2230 623 2234
rect 627 2230 687 2234
rect 691 2230 727 2234
rect 731 2230 791 2234
rect 795 2230 831 2234
rect 835 2230 895 2234
rect 899 2230 935 2234
rect 939 2230 999 2234
rect 1003 2230 1039 2234
rect 1043 2230 1111 2234
rect 1115 2230 1143 2234
rect 1147 2230 1223 2234
rect 1227 2230 1287 2234
rect 1291 2230 1299 2234
rect 91 2229 1299 2230
rect 1305 2234 2534 2235
rect 1305 2230 1327 2234
rect 1331 2230 1367 2234
rect 1371 2230 1463 2234
rect 1467 2230 1487 2234
rect 1491 2230 1567 2234
rect 1571 2230 1607 2234
rect 1611 2230 1671 2234
rect 1675 2230 1719 2234
rect 1723 2230 1775 2234
rect 1779 2230 1815 2234
rect 1819 2230 1887 2234
rect 1891 2230 1903 2234
rect 1907 2230 1983 2234
rect 1987 2230 1999 2234
rect 2003 2230 2055 2234
rect 2059 2230 2111 2234
rect 2115 2230 2127 2234
rect 2131 2230 2191 2234
rect 2195 2230 2223 2234
rect 2227 2230 2255 2234
rect 2259 2230 2319 2234
rect 2323 2230 2383 2234
rect 2387 2230 2439 2234
rect 2443 2230 2503 2234
rect 2507 2230 2534 2234
rect 1305 2229 2534 2230
rect 1718 2220 1724 2221
rect 2246 2220 2252 2221
rect 1718 2216 1719 2220
rect 1723 2216 2247 2220
rect 2251 2216 2252 2220
rect 1718 2215 1724 2216
rect 2246 2215 2252 2216
rect 96 2177 97 2183
rect 103 2182 1311 2183
rect 103 2178 111 2182
rect 115 2178 159 2182
rect 163 2178 247 2182
rect 251 2178 255 2182
rect 259 2178 335 2182
rect 339 2178 351 2182
rect 355 2178 431 2182
rect 435 2178 455 2182
rect 459 2178 535 2182
rect 539 2178 559 2182
rect 563 2178 639 2182
rect 643 2178 663 2182
rect 667 2178 743 2182
rect 747 2178 767 2182
rect 771 2178 847 2182
rect 851 2178 863 2182
rect 867 2178 951 2182
rect 955 2178 959 2182
rect 963 2178 1055 2182
rect 1059 2178 1159 2182
rect 1163 2178 1239 2182
rect 1243 2178 1287 2182
rect 1291 2178 1311 2182
rect 103 2177 1311 2178
rect 1317 2177 1318 2183
rect 1310 2157 1311 2163
rect 1317 2162 2539 2163
rect 1317 2158 1327 2162
rect 1331 2158 1383 2162
rect 1387 2158 1407 2162
rect 1411 2158 1503 2162
rect 1507 2158 1623 2162
rect 1627 2158 1735 2162
rect 1739 2158 1815 2162
rect 1819 2158 1831 2162
rect 1835 2158 1919 2162
rect 1923 2158 1991 2162
rect 1995 2158 1999 2162
rect 2003 2158 2071 2162
rect 2075 2158 2143 2162
rect 2147 2158 2159 2162
rect 2163 2158 2207 2162
rect 2211 2158 2271 2162
rect 2275 2158 2319 2162
rect 2323 2158 2335 2162
rect 2339 2158 2399 2162
rect 2403 2158 2455 2162
rect 2459 2158 2503 2162
rect 2507 2158 2539 2162
rect 1317 2157 2539 2158
rect 2545 2157 2546 2163
rect 84 2125 85 2131
rect 91 2130 1299 2131
rect 91 2126 111 2130
rect 115 2126 239 2130
rect 243 2126 303 2130
rect 307 2126 335 2130
rect 339 2126 359 2130
rect 363 2126 423 2130
rect 427 2126 439 2130
rect 443 2126 487 2130
rect 491 2126 543 2130
rect 547 2126 559 2130
rect 563 2126 631 2130
rect 635 2126 647 2130
rect 651 2126 711 2130
rect 715 2126 751 2130
rect 755 2126 799 2130
rect 803 2126 847 2130
rect 851 2126 887 2130
rect 891 2126 943 2130
rect 947 2126 975 2130
rect 979 2126 1039 2130
rect 1043 2126 1063 2130
rect 1067 2126 1143 2130
rect 1147 2126 1151 2130
rect 1155 2126 1223 2130
rect 1227 2126 1287 2130
rect 1291 2126 1299 2130
rect 91 2125 1299 2126
rect 1305 2125 1306 2131
rect 1298 2105 1299 2111
rect 1305 2110 2527 2111
rect 1305 2106 1327 2110
rect 1331 2106 1383 2110
rect 1387 2106 1391 2110
rect 1395 2106 1551 2110
rect 1555 2106 1607 2110
rect 1611 2106 1711 2110
rect 1715 2106 1799 2110
rect 1803 2106 1855 2110
rect 1859 2106 1975 2110
rect 1979 2106 1991 2110
rect 1995 2106 2119 2110
rect 2123 2106 2143 2110
rect 2147 2106 2239 2110
rect 2243 2106 2303 2110
rect 2307 2106 2367 2110
rect 2371 2106 2439 2110
rect 2443 2106 2503 2110
rect 2507 2106 2527 2110
rect 1305 2105 2527 2106
rect 2533 2105 2534 2111
rect 96 2069 97 2075
rect 103 2074 1311 2075
rect 103 2070 111 2074
rect 115 2070 319 2074
rect 323 2070 375 2074
rect 379 2070 399 2074
rect 403 2070 439 2074
rect 443 2070 455 2074
rect 459 2070 503 2074
rect 507 2070 511 2074
rect 515 2070 575 2074
rect 579 2070 639 2074
rect 643 2070 647 2074
rect 651 2070 711 2074
rect 715 2070 727 2074
rect 731 2070 791 2074
rect 795 2070 815 2074
rect 819 2070 863 2074
rect 867 2070 903 2074
rect 907 2070 943 2074
rect 947 2070 991 2074
rect 995 2070 1023 2074
rect 1027 2070 1079 2074
rect 1083 2070 1103 2074
rect 1107 2070 1167 2074
rect 1171 2070 1183 2074
rect 1187 2070 1239 2074
rect 1243 2070 1287 2074
rect 1291 2070 1311 2074
rect 103 2069 1311 2070
rect 1317 2069 1318 2075
rect 1310 2049 1311 2055
rect 1317 2054 2539 2055
rect 1317 2050 1327 2054
rect 1331 2050 1399 2054
rect 1403 2050 1447 2054
rect 1451 2050 1551 2054
rect 1555 2050 1567 2054
rect 1571 2050 1655 2054
rect 1659 2050 1727 2054
rect 1731 2050 1751 2054
rect 1755 2050 1839 2054
rect 1843 2050 1871 2054
rect 1875 2050 1927 2054
rect 1931 2050 2007 2054
rect 2011 2050 2023 2054
rect 2027 2050 2119 2054
rect 2123 2050 2135 2054
rect 2139 2050 2255 2054
rect 2259 2050 2383 2054
rect 2387 2050 2503 2054
rect 2507 2050 2539 2054
rect 1317 2049 2539 2050
rect 2545 2049 2546 2055
rect 84 2013 85 2019
rect 91 2018 1299 2019
rect 91 2014 111 2018
rect 115 2014 231 2018
rect 235 2014 287 2018
rect 291 2014 359 2018
rect 363 2014 383 2018
rect 387 2014 439 2018
rect 443 2014 495 2018
rect 499 2014 535 2018
rect 539 2014 559 2018
rect 563 2014 623 2018
rect 627 2014 631 2018
rect 635 2014 695 2018
rect 699 2014 735 2018
rect 739 2014 775 2018
rect 779 2014 847 2018
rect 851 2014 927 2018
rect 931 2014 959 2018
rect 963 2014 1007 2018
rect 1011 2014 1079 2018
rect 1083 2014 1087 2018
rect 1091 2014 1167 2018
rect 1171 2014 1199 2018
rect 1203 2014 1223 2018
rect 1227 2014 1287 2018
rect 1291 2014 1299 2018
rect 91 2013 1299 2014
rect 1305 2013 1306 2019
rect 1298 1993 1299 1999
rect 1305 1998 2527 1999
rect 1305 1994 1327 1998
rect 1331 1994 1431 1998
rect 1435 1994 1455 1998
rect 1459 1994 1511 1998
rect 1515 1994 1535 1998
rect 1539 1994 1575 1998
rect 1579 1994 1639 1998
rect 1643 1994 1703 1998
rect 1707 1994 1735 1998
rect 1739 1994 1767 1998
rect 1771 1994 1823 1998
rect 1827 1994 1831 1998
rect 1835 1994 1895 1998
rect 1899 1994 1911 1998
rect 1915 1994 1959 1998
rect 1963 1994 2007 1998
rect 2011 1994 2031 1998
rect 2035 1994 2103 1998
rect 2107 1994 2503 1998
rect 2507 1994 2527 1998
rect 1305 1993 2527 1994
rect 2533 1993 2534 1999
rect 230 1980 236 1981
rect 654 1980 660 1981
rect 230 1976 231 1980
rect 235 1976 655 1980
rect 659 1976 660 1980
rect 230 1975 236 1976
rect 654 1975 660 1976
rect 96 1957 97 1963
rect 103 1962 1311 1963
rect 103 1958 111 1962
rect 115 1958 151 1962
rect 155 1958 215 1962
rect 219 1958 247 1962
rect 251 1958 303 1962
rect 307 1958 319 1962
rect 323 1958 375 1962
rect 379 1958 439 1962
rect 443 1958 455 1962
rect 459 1958 551 1962
rect 555 1958 583 1962
rect 587 1958 647 1962
rect 651 1958 743 1962
rect 747 1958 751 1962
rect 755 1958 863 1962
rect 867 1958 919 1962
rect 923 1958 975 1962
rect 979 1958 1095 1962
rect 1099 1958 1215 1962
rect 1219 1958 1287 1962
rect 1291 1958 1311 1962
rect 103 1957 1311 1958
rect 1317 1957 1318 1963
rect 166 1940 172 1941
rect 602 1940 608 1941
rect 166 1936 167 1940
rect 171 1936 603 1940
rect 607 1936 608 1940
rect 1310 1937 1311 1943
rect 1317 1942 2539 1943
rect 1317 1938 1327 1942
rect 1331 1938 1471 1942
rect 1475 1938 1527 1942
rect 1531 1938 1567 1942
rect 1571 1938 1591 1942
rect 1595 1938 1631 1942
rect 1635 1938 1655 1942
rect 1659 1938 1703 1942
rect 1707 1938 1719 1942
rect 1723 1938 1775 1942
rect 1779 1938 1783 1942
rect 1787 1938 1847 1942
rect 1851 1938 1911 1942
rect 1915 1938 1919 1942
rect 1923 1938 1975 1942
rect 1979 1938 1999 1942
rect 2003 1938 2047 1942
rect 2051 1938 2087 1942
rect 2091 1938 2183 1942
rect 2187 1938 2279 1942
rect 2283 1938 2375 1942
rect 2379 1938 2455 1942
rect 2459 1938 2503 1942
rect 2507 1938 2539 1942
rect 1317 1937 2539 1938
rect 2545 1937 2546 1943
rect 166 1935 172 1936
rect 602 1935 608 1936
rect 84 1897 85 1903
rect 91 1902 1299 1903
rect 91 1898 111 1902
rect 115 1898 135 1902
rect 139 1898 191 1902
rect 195 1898 199 1902
rect 203 1898 271 1902
rect 275 1898 303 1902
rect 307 1898 359 1902
rect 363 1898 423 1902
rect 427 1898 455 1902
rect 459 1898 543 1902
rect 547 1898 567 1902
rect 571 1898 631 1902
rect 635 1898 719 1902
rect 723 1898 727 1902
rect 731 1898 799 1902
rect 803 1898 871 1902
rect 875 1898 903 1902
rect 907 1898 943 1902
rect 947 1898 1015 1902
rect 1019 1898 1079 1902
rect 1083 1898 1087 1902
rect 1091 1898 1159 1902
rect 1163 1898 1287 1902
rect 1291 1898 1299 1902
rect 91 1897 1299 1898
rect 1305 1897 1306 1903
rect 1298 1881 1299 1887
rect 1305 1886 2527 1887
rect 1305 1882 1327 1886
rect 1331 1882 1551 1886
rect 1555 1882 1607 1886
rect 1611 1882 1615 1886
rect 1619 1882 1663 1886
rect 1667 1882 1687 1886
rect 1691 1882 1727 1886
rect 1731 1882 1759 1886
rect 1763 1882 1799 1886
rect 1803 1882 1831 1886
rect 1835 1882 1871 1886
rect 1875 1882 1903 1886
rect 1907 1882 1943 1886
rect 1947 1882 1983 1886
rect 1987 1882 2007 1886
rect 2011 1882 2071 1886
rect 2075 1882 2135 1886
rect 2139 1882 2167 1886
rect 2171 1882 2199 1886
rect 2203 1882 2263 1886
rect 2267 1882 2327 1886
rect 2331 1882 2359 1886
rect 2363 1882 2383 1886
rect 2387 1882 2439 1886
rect 2443 1882 2503 1886
rect 2507 1882 2527 1886
rect 1305 1881 2527 1882
rect 2533 1881 2534 1887
rect 96 1845 97 1851
rect 103 1850 1311 1851
rect 103 1846 111 1850
rect 115 1846 151 1850
rect 155 1846 207 1850
rect 211 1846 287 1850
rect 291 1846 295 1850
rect 299 1846 375 1850
rect 379 1846 391 1850
rect 395 1846 471 1850
rect 475 1846 495 1850
rect 499 1846 559 1850
rect 563 1846 591 1850
rect 595 1846 647 1850
rect 651 1846 687 1850
rect 691 1846 735 1850
rect 739 1846 775 1850
rect 779 1846 815 1850
rect 819 1846 855 1850
rect 859 1846 887 1850
rect 891 1846 927 1850
rect 931 1846 959 1850
rect 963 1846 999 1850
rect 1003 1846 1031 1850
rect 1035 1846 1079 1850
rect 1083 1846 1103 1850
rect 1107 1846 1159 1850
rect 1163 1846 1175 1850
rect 1179 1846 1287 1850
rect 1291 1846 1311 1850
rect 103 1845 1311 1846
rect 1317 1845 1318 1851
rect 1310 1825 1311 1831
rect 1317 1830 2539 1831
rect 1317 1826 1327 1830
rect 1331 1826 1623 1830
rect 1627 1826 1631 1830
rect 1635 1826 1679 1830
rect 1683 1826 1719 1830
rect 1723 1826 1743 1830
rect 1747 1826 1815 1830
rect 1819 1826 1887 1830
rect 1891 1826 1927 1830
rect 1931 1826 1959 1830
rect 1963 1826 2023 1830
rect 2027 1826 2055 1830
rect 2059 1826 2087 1830
rect 2091 1826 2151 1830
rect 2155 1826 2191 1830
rect 2195 1826 2215 1830
rect 2219 1826 2279 1830
rect 2283 1826 2335 1830
rect 2339 1826 2343 1830
rect 2347 1826 2399 1830
rect 2403 1826 2455 1830
rect 2459 1826 2503 1830
rect 2507 1826 2539 1830
rect 1317 1825 2539 1826
rect 2545 1825 2546 1831
rect 84 1781 85 1787
rect 91 1786 1299 1787
rect 91 1782 111 1786
rect 115 1782 135 1786
rect 139 1782 191 1786
rect 195 1782 199 1786
rect 203 1782 279 1786
rect 283 1782 295 1786
rect 299 1782 375 1786
rect 379 1782 399 1786
rect 403 1782 479 1786
rect 483 1782 503 1786
rect 507 1782 575 1786
rect 579 1782 607 1786
rect 611 1782 671 1786
rect 675 1782 703 1786
rect 707 1782 759 1786
rect 763 1782 799 1786
rect 803 1782 839 1786
rect 843 1782 887 1786
rect 891 1782 911 1786
rect 915 1782 975 1786
rect 979 1782 983 1786
rect 987 1782 1063 1786
rect 1067 1782 1143 1786
rect 1147 1782 1151 1786
rect 1155 1782 1287 1786
rect 1291 1782 1299 1786
rect 91 1781 1299 1782
rect 1305 1781 1306 1787
rect 1298 1779 1306 1781
rect 1298 1773 1299 1779
rect 1305 1778 2527 1779
rect 1305 1774 1327 1778
rect 1331 1774 1527 1778
rect 1531 1774 1607 1778
rect 1611 1774 1615 1778
rect 1619 1774 1695 1778
rect 1699 1774 1703 1778
rect 1707 1774 1791 1778
rect 1795 1774 1799 1778
rect 1803 1774 1879 1778
rect 1883 1774 1911 1778
rect 1915 1774 1967 1778
rect 1971 1774 2039 1778
rect 2043 1774 2055 1778
rect 2059 1774 2135 1778
rect 2139 1774 2175 1778
rect 2179 1774 2215 1778
rect 2219 1774 2295 1778
rect 2299 1774 2319 1778
rect 2323 1774 2375 1778
rect 2379 1774 2439 1778
rect 2443 1774 2503 1778
rect 2507 1774 2527 1778
rect 1305 1773 2527 1774
rect 2533 1773 2534 1779
rect 134 1772 140 1773
rect 510 1772 516 1773
rect 134 1768 135 1772
rect 139 1768 511 1772
rect 515 1768 516 1772
rect 134 1767 140 1768
rect 510 1767 516 1768
rect 1654 1756 1660 1757
rect 1914 1756 1920 1757
rect 1654 1752 1655 1756
rect 1659 1752 1915 1756
rect 1919 1752 1920 1756
rect 1654 1751 1660 1752
rect 1914 1751 1920 1752
rect 96 1725 97 1731
rect 103 1730 1311 1731
rect 103 1726 111 1730
rect 115 1726 151 1730
rect 155 1726 167 1730
rect 171 1726 215 1730
rect 219 1726 239 1730
rect 243 1726 311 1730
rect 315 1726 319 1730
rect 323 1726 407 1730
rect 411 1726 415 1730
rect 419 1726 503 1730
rect 507 1726 519 1730
rect 523 1726 607 1730
rect 611 1726 623 1730
rect 627 1726 711 1730
rect 715 1726 719 1730
rect 723 1726 815 1730
rect 819 1726 823 1730
rect 827 1726 903 1730
rect 907 1726 935 1730
rect 939 1726 991 1730
rect 995 1726 1047 1730
rect 1051 1726 1079 1730
rect 1083 1726 1159 1730
rect 1163 1726 1167 1730
rect 1171 1726 1287 1730
rect 1291 1726 1311 1730
rect 103 1725 1311 1726
rect 1317 1725 1318 1731
rect 1310 1723 1318 1725
rect 1310 1717 1311 1723
rect 1317 1722 2539 1723
rect 1317 1718 1327 1722
rect 1331 1718 1399 1722
rect 1403 1718 1463 1722
rect 1467 1718 1543 1722
rect 1547 1718 1623 1722
rect 1627 1718 1631 1722
rect 1635 1718 1711 1722
rect 1715 1718 1727 1722
rect 1731 1718 1807 1722
rect 1811 1718 1823 1722
rect 1827 1718 1895 1722
rect 1899 1718 1919 1722
rect 1923 1718 1983 1722
rect 1987 1718 2015 1722
rect 2019 1718 2071 1722
rect 2075 1718 2111 1722
rect 2115 1718 2151 1722
rect 2155 1718 2199 1722
rect 2203 1718 2231 1722
rect 2235 1718 2287 1722
rect 2291 1718 2311 1722
rect 2315 1718 2383 1722
rect 2387 1718 2391 1722
rect 2395 1718 2455 1722
rect 2459 1718 2503 1722
rect 2507 1718 2539 1722
rect 1317 1717 2539 1718
rect 2545 1717 2546 1723
rect 1594 1700 1600 1701
rect 1842 1700 1848 1701
rect 1594 1696 1595 1700
rect 1599 1696 1843 1700
rect 1847 1696 1848 1700
rect 1594 1695 1600 1696
rect 1842 1695 1848 1696
rect 84 1669 85 1675
rect 91 1674 1299 1675
rect 91 1670 111 1674
rect 115 1670 151 1674
rect 155 1670 223 1674
rect 227 1670 255 1674
rect 259 1670 303 1674
rect 307 1670 319 1674
rect 323 1670 391 1674
rect 395 1670 399 1674
rect 403 1670 487 1674
rect 491 1670 575 1674
rect 579 1670 591 1674
rect 595 1670 671 1674
rect 675 1670 695 1674
rect 699 1670 767 1674
rect 771 1670 807 1674
rect 811 1670 863 1674
rect 867 1670 919 1674
rect 923 1670 959 1674
rect 963 1670 1031 1674
rect 1035 1670 1063 1674
rect 1067 1670 1143 1674
rect 1147 1670 1167 1674
rect 1171 1670 1287 1674
rect 1291 1670 1299 1674
rect 91 1669 1299 1670
rect 1305 1669 1306 1675
rect 1298 1667 1306 1669
rect 1298 1661 1299 1667
rect 1305 1666 2527 1667
rect 1305 1662 1327 1666
rect 1331 1662 1351 1666
rect 1355 1662 1383 1666
rect 1387 1662 1407 1666
rect 1411 1662 1447 1666
rect 1451 1662 1495 1666
rect 1499 1662 1527 1666
rect 1531 1662 1583 1666
rect 1587 1662 1615 1666
rect 1619 1662 1679 1666
rect 1683 1662 1711 1666
rect 1715 1662 1783 1666
rect 1787 1662 1807 1666
rect 1811 1662 1895 1666
rect 1899 1662 1903 1666
rect 1907 1662 1999 1666
rect 2003 1662 2023 1666
rect 2027 1662 2095 1666
rect 2099 1662 2159 1666
rect 2163 1662 2183 1666
rect 2187 1662 2271 1666
rect 2275 1662 2303 1666
rect 2307 1662 2367 1666
rect 2371 1662 2439 1666
rect 2443 1662 2503 1666
rect 2507 1662 2527 1666
rect 1305 1661 2527 1662
rect 2533 1661 2534 1667
rect 1414 1644 1420 1645
rect 1702 1644 1708 1645
rect 1414 1640 1415 1644
rect 1419 1640 1703 1644
rect 1707 1640 1708 1644
rect 1414 1639 1420 1640
rect 1702 1639 1708 1640
rect 96 1613 97 1619
rect 103 1618 1311 1619
rect 103 1614 111 1618
rect 115 1614 271 1618
rect 275 1614 303 1618
rect 307 1614 335 1618
rect 339 1614 359 1618
rect 363 1614 415 1618
rect 419 1614 431 1618
rect 435 1614 503 1618
rect 507 1614 511 1618
rect 515 1614 591 1618
rect 595 1614 599 1618
rect 603 1614 687 1618
rect 691 1614 695 1618
rect 699 1614 783 1618
rect 787 1614 791 1618
rect 795 1614 879 1618
rect 883 1614 895 1618
rect 899 1614 975 1618
rect 979 1614 1007 1618
rect 1011 1614 1079 1618
rect 1083 1614 1119 1618
rect 1123 1614 1183 1618
rect 1187 1614 1287 1618
rect 1291 1614 1311 1618
rect 103 1613 1311 1614
rect 1317 1615 1318 1619
rect 1317 1614 2546 1615
rect 1317 1613 1327 1614
rect 1310 1610 1327 1613
rect 1331 1610 1367 1614
rect 1371 1610 1423 1614
rect 1427 1610 1479 1614
rect 1483 1610 1511 1614
rect 1515 1610 1559 1614
rect 1563 1610 1599 1614
rect 1603 1610 1639 1614
rect 1643 1610 1695 1614
rect 1699 1610 1719 1614
rect 1723 1610 1791 1614
rect 1795 1610 1799 1614
rect 1803 1610 1871 1614
rect 1875 1610 1911 1614
rect 1915 1610 1951 1614
rect 1955 1610 2031 1614
rect 2035 1610 2039 1614
rect 2043 1610 2175 1614
rect 2179 1610 2319 1614
rect 2323 1610 2455 1614
rect 2459 1610 2503 1614
rect 2507 1610 2546 1614
rect 1310 1609 2546 1610
rect 84 1561 85 1567
rect 91 1566 1299 1567
rect 91 1562 111 1566
rect 115 1562 247 1566
rect 251 1562 287 1566
rect 291 1562 319 1566
rect 323 1562 343 1566
rect 347 1562 399 1566
rect 403 1562 415 1566
rect 419 1562 487 1566
rect 491 1562 495 1566
rect 499 1562 583 1566
rect 587 1562 671 1566
rect 675 1562 679 1566
rect 683 1562 759 1566
rect 763 1562 775 1566
rect 779 1562 847 1566
rect 851 1562 879 1566
rect 883 1562 927 1566
rect 931 1562 991 1566
rect 995 1562 1007 1566
rect 1011 1562 1087 1566
rect 1091 1562 1103 1566
rect 1107 1562 1167 1566
rect 1171 1562 1223 1566
rect 1227 1562 1287 1566
rect 1291 1562 1299 1566
rect 91 1561 1299 1562
rect 1305 1563 1306 1567
rect 1305 1562 2534 1563
rect 1305 1561 1327 1562
rect 1298 1558 1327 1561
rect 1331 1558 1351 1562
rect 1355 1558 1407 1562
rect 1411 1558 1463 1562
rect 1467 1558 1471 1562
rect 1475 1558 1543 1562
rect 1547 1558 1607 1562
rect 1611 1558 1623 1562
rect 1627 1558 1703 1562
rect 1707 1558 1735 1562
rect 1739 1558 1775 1562
rect 1779 1558 1855 1562
rect 1859 1558 1871 1562
rect 1875 1558 1935 1562
rect 1939 1558 2007 1562
rect 2011 1558 2015 1562
rect 2019 1558 2503 1562
rect 2507 1558 2534 1562
rect 1298 1557 2534 1558
rect 1310 1510 2546 1511
rect 1310 1507 1327 1510
rect 96 1501 97 1507
rect 103 1506 1311 1507
rect 103 1502 111 1506
rect 115 1502 263 1506
rect 267 1502 279 1506
rect 283 1502 335 1506
rect 339 1502 343 1506
rect 347 1502 415 1506
rect 419 1502 495 1506
rect 499 1502 503 1506
rect 507 1502 575 1506
rect 579 1502 599 1506
rect 603 1502 655 1506
rect 659 1502 687 1506
rect 691 1502 735 1506
rect 739 1502 775 1506
rect 779 1502 815 1506
rect 819 1502 863 1506
rect 867 1502 895 1506
rect 899 1502 943 1506
rect 947 1502 975 1506
rect 979 1502 1023 1506
rect 1027 1502 1055 1506
rect 1059 1502 1103 1506
rect 1107 1502 1143 1506
rect 1147 1502 1183 1506
rect 1187 1502 1239 1506
rect 1243 1502 1287 1506
rect 1291 1502 1311 1506
rect 103 1501 1311 1502
rect 1317 1506 1327 1507
rect 1331 1506 1367 1510
rect 1371 1506 1423 1510
rect 1427 1506 1479 1510
rect 1483 1506 1487 1510
rect 1491 1506 1551 1510
rect 1555 1506 1623 1510
rect 1627 1506 1631 1510
rect 1635 1506 1711 1510
rect 1715 1506 1751 1510
rect 1755 1506 1791 1510
rect 1795 1506 1871 1510
rect 1875 1506 1887 1510
rect 1891 1506 1951 1510
rect 1955 1506 2023 1510
rect 2027 1506 2031 1510
rect 2035 1506 2119 1510
rect 2123 1506 2503 1510
rect 2507 1506 2546 1510
rect 1317 1505 2546 1506
rect 1317 1501 1318 1505
rect 84 1445 85 1451
rect 91 1450 1299 1451
rect 91 1446 111 1450
rect 115 1446 191 1450
rect 195 1446 255 1450
rect 259 1446 263 1450
rect 267 1446 327 1450
rect 331 1446 399 1450
rect 403 1446 407 1450
rect 411 1446 479 1450
rect 483 1446 503 1450
rect 507 1446 559 1450
rect 563 1446 607 1450
rect 611 1446 639 1450
rect 643 1446 711 1450
rect 715 1446 719 1450
rect 723 1446 799 1450
rect 803 1446 815 1450
rect 819 1446 879 1450
rect 883 1446 919 1450
rect 923 1446 959 1450
rect 963 1446 1023 1450
rect 1027 1446 1039 1450
rect 1043 1446 1127 1450
rect 1131 1446 1223 1450
rect 1227 1446 1287 1450
rect 1291 1446 1299 1450
rect 91 1445 1299 1446
rect 1305 1450 2534 1451
rect 1305 1446 1327 1450
rect 1331 1446 1351 1450
rect 1355 1446 1359 1450
rect 1363 1446 1407 1450
rect 1411 1446 1447 1450
rect 1451 1446 1463 1450
rect 1467 1446 1535 1450
rect 1539 1446 1615 1450
rect 1619 1446 1631 1450
rect 1635 1446 1695 1450
rect 1699 1446 1727 1450
rect 1731 1446 1775 1450
rect 1779 1446 1815 1450
rect 1819 1446 1855 1450
rect 1859 1446 1903 1450
rect 1907 1446 1935 1450
rect 1939 1446 1991 1450
rect 1995 1446 2015 1450
rect 2019 1446 2071 1450
rect 2075 1446 2103 1450
rect 2107 1446 2159 1450
rect 2163 1446 2247 1450
rect 2251 1446 2503 1450
rect 2507 1446 2534 1450
rect 1305 1445 2534 1446
rect 1310 1398 2546 1399
rect 1310 1395 1327 1398
rect 96 1389 97 1395
rect 103 1394 1311 1395
rect 103 1390 111 1394
rect 115 1390 151 1394
rect 155 1390 207 1394
rect 211 1390 223 1394
rect 227 1390 271 1394
rect 275 1390 295 1394
rect 299 1390 343 1394
rect 347 1390 359 1394
rect 363 1390 423 1394
rect 427 1390 431 1394
rect 435 1390 503 1394
rect 507 1390 519 1394
rect 523 1390 583 1394
rect 587 1390 623 1394
rect 627 1390 663 1394
rect 667 1390 727 1394
rect 731 1390 751 1394
rect 755 1390 831 1394
rect 835 1390 839 1394
rect 843 1390 927 1394
rect 931 1390 935 1394
rect 939 1390 1015 1394
rect 1019 1390 1039 1394
rect 1043 1390 1103 1394
rect 1107 1390 1143 1394
rect 1147 1390 1199 1394
rect 1203 1390 1239 1394
rect 1243 1390 1287 1394
rect 1291 1390 1311 1394
rect 103 1389 1311 1390
rect 1317 1394 1327 1395
rect 1331 1394 1375 1398
rect 1379 1394 1463 1398
rect 1467 1394 1551 1398
rect 1555 1394 1567 1398
rect 1571 1394 1647 1398
rect 1651 1394 1735 1398
rect 1739 1394 1743 1398
rect 1747 1394 1831 1398
rect 1835 1394 1919 1398
rect 1923 1394 2007 1398
rect 2011 1394 2087 1398
rect 2091 1394 2095 1398
rect 2099 1394 2175 1398
rect 2179 1394 2247 1398
rect 2251 1394 2263 1398
rect 2267 1394 2319 1398
rect 2323 1394 2399 1398
rect 2403 1394 2455 1398
rect 2459 1394 2503 1398
rect 2507 1394 2546 1398
rect 1317 1393 2546 1394
rect 1317 1389 1318 1393
rect 1298 1341 1299 1347
rect 1305 1346 2527 1347
rect 1305 1342 1327 1346
rect 1331 1342 1551 1346
rect 1555 1342 1583 1346
rect 1587 1342 1631 1346
rect 1635 1342 1647 1346
rect 1651 1342 1719 1346
rect 1723 1342 1727 1346
rect 1731 1342 1807 1346
rect 1811 1342 1815 1346
rect 1819 1342 1895 1346
rect 1899 1342 1903 1346
rect 1907 1342 1983 1346
rect 1987 1342 1991 1346
rect 1995 1342 2063 1346
rect 2067 1342 2079 1346
rect 2083 1342 2143 1346
rect 2147 1342 2159 1346
rect 2163 1342 2223 1346
rect 2227 1342 2231 1346
rect 2235 1342 2303 1346
rect 2307 1342 2383 1346
rect 2387 1342 2439 1346
rect 2443 1342 2503 1346
rect 2507 1342 2527 1346
rect 1305 1341 2527 1342
rect 2533 1341 2534 1347
rect 84 1321 85 1327
rect 91 1326 1299 1327
rect 91 1322 111 1326
rect 115 1322 135 1326
rect 139 1322 207 1326
rect 211 1322 239 1326
rect 243 1322 279 1326
rect 283 1322 343 1326
rect 347 1322 367 1326
rect 371 1322 415 1326
rect 419 1322 479 1326
rect 483 1322 487 1326
rect 491 1322 567 1326
rect 571 1322 583 1326
rect 587 1322 647 1326
rect 651 1322 687 1326
rect 691 1322 735 1326
rect 739 1322 783 1326
rect 787 1322 823 1326
rect 827 1322 879 1326
rect 883 1322 911 1326
rect 915 1322 975 1326
rect 979 1322 999 1326
rect 1003 1322 1087 1326
rect 1091 1322 1183 1326
rect 1187 1322 1287 1326
rect 1291 1322 1299 1326
rect 91 1321 1299 1322
rect 1305 1321 1306 1327
rect 1310 1289 1311 1295
rect 1317 1294 2539 1295
rect 1317 1290 1327 1294
rect 1331 1290 1567 1294
rect 1571 1290 1599 1294
rect 1603 1290 1631 1294
rect 1635 1290 1663 1294
rect 1667 1290 1711 1294
rect 1715 1290 1743 1294
rect 1747 1290 1799 1294
rect 1803 1290 1823 1294
rect 1827 1290 1895 1294
rect 1899 1290 1911 1294
rect 1915 1290 1991 1294
rect 1995 1290 1999 1294
rect 2003 1290 2079 1294
rect 2083 1290 2095 1294
rect 2099 1290 2159 1294
rect 2163 1290 2207 1294
rect 2211 1290 2239 1294
rect 2243 1290 2319 1294
rect 2323 1290 2399 1294
rect 2403 1290 2455 1294
rect 2459 1290 2503 1294
rect 2507 1290 2539 1294
rect 1317 1289 2539 1290
rect 2545 1289 2546 1295
rect 96 1261 97 1267
rect 103 1266 1311 1267
rect 103 1262 111 1266
rect 115 1262 151 1266
rect 155 1262 215 1266
rect 219 1262 255 1266
rect 259 1262 303 1266
rect 307 1262 383 1266
rect 387 1262 391 1266
rect 395 1262 471 1266
rect 475 1262 495 1266
rect 499 1262 551 1266
rect 555 1262 599 1266
rect 603 1262 623 1266
rect 627 1262 695 1266
rect 699 1262 703 1266
rect 707 1262 767 1266
rect 771 1262 799 1266
rect 803 1262 839 1266
rect 843 1262 895 1266
rect 899 1262 919 1266
rect 923 1262 991 1266
rect 995 1262 1287 1266
rect 1291 1262 1311 1266
rect 103 1261 1311 1262
rect 1317 1261 1318 1267
rect 1298 1233 1299 1239
rect 1305 1238 2527 1239
rect 1305 1234 1327 1238
rect 1331 1234 1519 1238
rect 1523 1234 1551 1238
rect 1555 1234 1575 1238
rect 1579 1234 1615 1238
rect 1619 1234 1631 1238
rect 1635 1234 1687 1238
rect 1691 1234 1695 1238
rect 1699 1234 1743 1238
rect 1747 1234 1783 1238
rect 1787 1234 1799 1238
rect 1803 1234 1855 1238
rect 1859 1234 1879 1238
rect 1883 1234 1911 1238
rect 1915 1234 1967 1238
rect 1971 1234 1975 1238
rect 1979 1234 2031 1238
rect 2035 1234 2079 1238
rect 2083 1234 2103 1238
rect 2107 1234 2183 1238
rect 2187 1234 2191 1238
rect 2195 1234 2271 1238
rect 2275 1234 2303 1238
rect 2307 1234 2367 1238
rect 2371 1234 2439 1238
rect 2443 1234 2503 1238
rect 2507 1234 2527 1238
rect 1305 1233 2527 1234
rect 2533 1233 2534 1239
rect 84 1205 85 1211
rect 91 1210 1299 1211
rect 91 1206 111 1210
rect 115 1206 135 1210
rect 139 1206 191 1210
rect 195 1206 199 1210
rect 203 1206 271 1210
rect 275 1206 287 1210
rect 291 1206 351 1210
rect 355 1206 375 1210
rect 379 1206 431 1210
rect 435 1206 455 1210
rect 459 1206 511 1210
rect 515 1206 535 1210
rect 539 1206 583 1210
rect 587 1206 607 1210
rect 611 1206 647 1210
rect 651 1206 679 1210
rect 683 1206 719 1210
rect 723 1206 751 1210
rect 755 1206 791 1210
rect 795 1206 823 1210
rect 827 1206 863 1210
rect 867 1206 903 1210
rect 907 1206 1287 1210
rect 1291 1206 1299 1210
rect 91 1205 1299 1206
rect 1305 1205 1306 1211
rect 1310 1177 1311 1183
rect 1317 1182 2539 1183
rect 1317 1178 1327 1182
rect 1331 1178 1535 1182
rect 1539 1178 1567 1182
rect 1571 1178 1591 1182
rect 1595 1178 1631 1182
rect 1635 1178 1647 1182
rect 1651 1178 1703 1182
rect 1707 1178 1759 1182
rect 1763 1178 1791 1182
rect 1795 1178 1815 1182
rect 1819 1178 1871 1182
rect 1875 1178 1903 1182
rect 1907 1178 1927 1182
rect 1931 1178 1983 1182
rect 1987 1178 2031 1182
rect 2035 1178 2047 1182
rect 2051 1178 2119 1182
rect 2123 1178 2175 1182
rect 2179 1178 2199 1182
rect 2203 1178 2287 1182
rect 2291 1178 2327 1182
rect 2331 1178 2383 1182
rect 2387 1178 2455 1182
rect 2459 1178 2503 1182
rect 2507 1178 2539 1182
rect 1317 1177 2539 1178
rect 2545 1177 2546 1183
rect 96 1149 97 1155
rect 103 1154 1311 1155
rect 103 1150 111 1154
rect 115 1150 151 1154
rect 155 1150 183 1154
rect 187 1150 207 1154
rect 211 1150 279 1154
rect 283 1150 287 1154
rect 291 1150 367 1154
rect 371 1150 375 1154
rect 379 1150 447 1154
rect 451 1150 471 1154
rect 475 1150 527 1154
rect 531 1150 567 1154
rect 571 1150 599 1154
rect 603 1150 655 1154
rect 659 1150 663 1154
rect 667 1150 735 1154
rect 739 1150 807 1154
rect 811 1150 879 1154
rect 883 1150 959 1154
rect 963 1150 1039 1154
rect 1043 1150 1287 1154
rect 1291 1150 1311 1154
rect 103 1149 1311 1150
rect 1317 1149 1318 1155
rect 1298 1125 1299 1131
rect 1305 1130 2527 1131
rect 1305 1126 1327 1130
rect 1331 1126 1383 1130
rect 1387 1126 1447 1130
rect 1451 1126 1519 1130
rect 1523 1126 1551 1130
rect 1555 1126 1591 1130
rect 1595 1126 1615 1130
rect 1619 1126 1671 1130
rect 1675 1126 1687 1130
rect 1691 1126 1751 1130
rect 1755 1126 1775 1130
rect 1779 1126 1831 1130
rect 1835 1126 1887 1130
rect 1891 1126 1911 1130
rect 1915 1126 1983 1130
rect 1987 1126 2015 1130
rect 2019 1126 2055 1130
rect 2059 1126 2135 1130
rect 2139 1126 2159 1130
rect 2163 1126 2215 1130
rect 2219 1126 2311 1130
rect 2315 1126 2439 1130
rect 2443 1126 2503 1130
rect 2507 1126 2527 1130
rect 1305 1125 2527 1126
rect 2533 1125 2534 1131
rect 84 1089 85 1095
rect 91 1094 1299 1095
rect 91 1090 111 1094
rect 115 1090 167 1094
rect 171 1090 207 1094
rect 211 1090 263 1094
rect 267 1090 279 1094
rect 283 1090 359 1094
rect 363 1090 447 1094
rect 451 1090 455 1094
rect 459 1090 543 1094
rect 547 1090 551 1094
rect 555 1090 639 1094
rect 643 1090 719 1094
rect 723 1090 727 1094
rect 731 1090 791 1094
rect 795 1090 815 1094
rect 819 1090 863 1094
rect 867 1090 895 1094
rect 899 1090 943 1094
rect 947 1090 975 1094
rect 979 1090 1023 1094
rect 1027 1090 1055 1094
rect 1059 1090 1143 1094
rect 1147 1090 1287 1094
rect 1291 1090 1299 1094
rect 91 1089 1299 1090
rect 1305 1089 1306 1095
rect 1310 1065 1311 1071
rect 1317 1070 2539 1071
rect 1317 1066 1327 1070
rect 1331 1066 1367 1070
rect 1371 1066 1399 1070
rect 1403 1066 1455 1070
rect 1459 1066 1463 1070
rect 1467 1066 1535 1070
rect 1539 1066 1575 1070
rect 1579 1066 1607 1070
rect 1611 1066 1687 1070
rect 1691 1066 1695 1070
rect 1699 1066 1767 1070
rect 1771 1066 1815 1070
rect 1819 1066 1847 1070
rect 1851 1066 1927 1070
rect 1931 1066 1999 1070
rect 2003 1066 2039 1070
rect 2043 1066 2071 1070
rect 2075 1066 2151 1070
rect 2155 1066 2231 1070
rect 2235 1066 2255 1070
rect 2259 1066 2367 1070
rect 2371 1066 2455 1070
rect 2459 1066 2503 1070
rect 2507 1066 2539 1070
rect 1317 1065 2539 1066
rect 2545 1065 2546 1071
rect 96 1029 97 1035
rect 103 1034 1311 1035
rect 103 1030 111 1034
rect 115 1030 223 1034
rect 227 1030 295 1034
rect 299 1030 375 1034
rect 379 1030 383 1034
rect 387 1030 463 1034
rect 467 1030 479 1034
rect 483 1030 559 1034
rect 563 1030 575 1034
rect 579 1030 655 1034
rect 659 1030 671 1034
rect 675 1030 743 1034
rect 747 1030 767 1034
rect 771 1030 831 1034
rect 835 1030 855 1034
rect 859 1030 911 1034
rect 915 1030 943 1034
rect 947 1030 991 1034
rect 995 1030 1023 1034
rect 1027 1030 1071 1034
rect 1075 1030 1103 1034
rect 1107 1030 1159 1034
rect 1163 1030 1183 1034
rect 1187 1030 1239 1034
rect 1243 1030 1287 1034
rect 1291 1030 1311 1034
rect 103 1029 1311 1030
rect 1317 1029 1318 1035
rect 1298 1009 1299 1015
rect 1305 1014 2527 1015
rect 1305 1010 1327 1014
rect 1331 1010 1351 1014
rect 1355 1010 1439 1014
rect 1443 1010 1511 1014
rect 1515 1010 1559 1014
rect 1563 1010 1679 1014
rect 1683 1010 1799 1014
rect 1803 1010 1823 1014
rect 1827 1010 1911 1014
rect 1915 1010 1951 1014
rect 1955 1010 2023 1014
rect 2027 1010 2071 1014
rect 2075 1010 2135 1014
rect 2139 1010 2175 1014
rect 2179 1010 2239 1014
rect 2243 1010 2271 1014
rect 2275 1010 2351 1014
rect 2355 1010 2367 1014
rect 2371 1010 2439 1014
rect 2443 1010 2503 1014
rect 2507 1010 2527 1014
rect 1305 1009 2527 1010
rect 2533 1009 2534 1015
rect 84 977 85 983
rect 91 982 1299 983
rect 91 978 111 982
rect 115 978 271 982
rect 275 978 279 982
rect 283 978 359 982
rect 363 978 367 982
rect 371 978 455 982
rect 459 978 463 982
rect 467 978 551 982
rect 555 978 559 982
rect 563 978 655 982
rect 659 978 751 982
rect 755 978 839 982
rect 843 978 927 982
rect 931 978 1007 982
rect 1011 978 1087 982
rect 1091 978 1167 982
rect 1171 978 1223 982
rect 1227 978 1287 982
rect 1291 978 1299 982
rect 91 977 1299 978
rect 1305 977 1306 983
rect 1822 972 1828 973
rect 2374 972 2380 973
rect 1822 968 1823 972
rect 1827 968 2375 972
rect 2379 968 2380 972
rect 1822 967 1828 968
rect 2374 967 2380 968
rect 1310 945 1311 951
rect 1317 950 2539 951
rect 1317 946 1327 950
rect 1331 946 1367 950
rect 1371 946 1423 950
rect 1427 946 1503 950
rect 1507 946 1527 950
rect 1531 946 1607 950
rect 1611 946 1695 950
rect 1699 946 1719 950
rect 1723 946 1831 950
rect 1835 946 1839 950
rect 1843 946 1935 950
rect 1939 946 1967 950
rect 1971 946 2031 950
rect 2035 946 2087 950
rect 2091 946 2127 950
rect 2131 946 2191 950
rect 2195 946 2215 950
rect 2219 946 2287 950
rect 2291 946 2295 950
rect 2299 946 2375 950
rect 2379 946 2383 950
rect 2387 946 2455 950
rect 2459 946 2503 950
rect 2507 946 2539 950
rect 1317 945 2539 946
rect 2545 945 2546 951
rect 96 917 97 923
rect 103 922 1311 923
rect 103 918 111 922
rect 115 918 271 922
rect 275 918 287 922
rect 291 918 343 922
rect 347 918 375 922
rect 379 918 423 922
rect 427 918 471 922
rect 475 918 519 922
rect 523 918 567 922
rect 571 918 615 922
rect 619 918 671 922
rect 675 918 711 922
rect 715 918 767 922
rect 771 918 807 922
rect 811 918 855 922
rect 859 918 903 922
rect 907 918 943 922
rect 947 918 991 922
rect 995 918 1023 922
rect 1027 918 1087 922
rect 1091 918 1103 922
rect 1107 918 1183 922
rect 1187 918 1239 922
rect 1243 918 1287 922
rect 1291 918 1311 922
rect 103 917 1311 918
rect 1317 917 1318 923
rect 1298 889 1299 895
rect 1305 894 2527 895
rect 1305 890 1327 894
rect 1331 890 1351 894
rect 1355 890 1407 894
rect 1411 890 1431 894
rect 1435 890 1487 894
rect 1491 890 1551 894
rect 1555 890 1591 894
rect 1595 890 1623 894
rect 1627 890 1703 894
rect 1707 890 1791 894
rect 1795 890 1815 894
rect 1819 890 1895 894
rect 1899 890 1919 894
rect 1923 890 2015 894
rect 2019 890 2111 894
rect 2115 890 2143 894
rect 2147 890 2199 894
rect 2203 890 2279 894
rect 2283 890 2359 894
rect 2363 890 2423 894
rect 2427 890 2439 894
rect 2443 890 2503 894
rect 2507 890 2527 894
rect 1305 889 2527 890
rect 2533 889 2534 895
rect 84 861 85 867
rect 91 866 1299 867
rect 91 862 111 866
rect 115 862 247 866
rect 251 862 255 866
rect 259 862 311 866
rect 315 862 327 866
rect 331 862 375 866
rect 379 862 407 866
rect 411 862 439 866
rect 443 862 503 866
rect 507 862 567 866
rect 571 862 599 866
rect 603 862 631 866
rect 635 862 695 866
rect 699 862 759 866
rect 763 862 791 866
rect 795 862 831 866
rect 835 862 887 866
rect 891 862 903 866
rect 907 862 975 866
rect 979 862 1071 866
rect 1075 862 1167 866
rect 1171 862 1287 866
rect 1291 862 1299 866
rect 91 861 1299 862
rect 1305 861 1306 867
rect 1310 833 1311 839
rect 1317 838 2539 839
rect 1317 834 1327 838
rect 1331 834 1447 838
rect 1451 834 1503 838
rect 1507 834 1567 838
rect 1571 834 1591 838
rect 1595 834 1639 838
rect 1643 834 1647 838
rect 1651 834 1703 838
rect 1707 834 1719 838
rect 1723 834 1767 838
rect 1771 834 1807 838
rect 1811 834 1847 838
rect 1851 834 1911 838
rect 1915 834 1927 838
rect 1931 834 2015 838
rect 2019 834 2031 838
rect 2035 834 2103 838
rect 2107 834 2159 838
rect 2163 834 2191 838
rect 2195 834 2287 838
rect 2291 834 2295 838
rect 2299 834 2383 838
rect 2387 834 2439 838
rect 2443 834 2455 838
rect 2459 834 2503 838
rect 2507 834 2539 838
rect 1317 833 2539 834
rect 2545 833 2546 839
rect 96 805 97 811
rect 103 810 1311 811
rect 103 806 111 810
rect 115 806 215 810
rect 219 806 263 810
rect 267 806 303 810
rect 307 806 327 810
rect 331 806 391 810
rect 395 806 455 810
rect 459 806 479 810
rect 483 806 519 810
rect 523 806 559 810
rect 563 806 583 810
rect 587 806 631 810
rect 635 806 647 810
rect 651 806 703 810
rect 707 806 711 810
rect 715 806 767 810
rect 771 806 775 810
rect 779 806 831 810
rect 835 806 847 810
rect 851 806 895 810
rect 899 806 919 810
rect 923 806 967 810
rect 971 806 1039 810
rect 1043 806 1287 810
rect 1291 806 1311 810
rect 103 805 1311 806
rect 1317 805 1318 811
rect 1298 777 1299 783
rect 1305 782 2527 783
rect 1305 778 1327 782
rect 1331 778 1567 782
rect 1571 778 1575 782
rect 1579 778 1623 782
rect 1627 778 1631 782
rect 1635 778 1687 782
rect 1691 778 1751 782
rect 1755 778 1759 782
rect 1763 778 1831 782
rect 1835 778 1911 782
rect 1915 778 1919 782
rect 1923 778 1999 782
rect 2003 778 2015 782
rect 2019 778 2087 782
rect 2091 778 2119 782
rect 2123 778 2175 782
rect 2179 778 2231 782
rect 2235 778 2271 782
rect 2275 778 2343 782
rect 2347 778 2367 782
rect 2371 778 2439 782
rect 2443 778 2503 782
rect 2507 778 2527 782
rect 1305 777 2527 778
rect 2533 777 2534 783
rect 84 753 85 759
rect 91 758 1299 759
rect 91 754 111 758
rect 115 754 135 758
rect 139 754 199 758
rect 203 754 255 758
rect 259 754 287 758
rect 291 754 375 758
rect 379 754 391 758
rect 395 754 463 758
rect 467 754 519 758
rect 523 754 543 758
rect 547 754 615 758
rect 619 754 647 758
rect 651 754 687 758
rect 691 754 751 758
rect 755 754 775 758
rect 779 754 815 758
rect 819 754 879 758
rect 883 754 903 758
rect 907 754 951 758
rect 955 754 1023 758
rect 1027 754 1039 758
rect 1043 754 1287 758
rect 1291 754 1299 758
rect 91 753 1299 754
rect 1305 753 1306 759
rect 1310 725 1311 731
rect 1317 730 2539 731
rect 1317 726 1327 730
rect 1331 726 1367 730
rect 1371 726 1431 730
rect 1435 726 1527 730
rect 1531 726 1583 730
rect 1587 726 1631 730
rect 1635 726 1639 730
rect 1643 726 1703 730
rect 1707 726 1735 730
rect 1739 726 1775 730
rect 1779 726 1839 730
rect 1843 726 1847 730
rect 1851 726 1935 730
rect 1939 726 1943 730
rect 1947 726 2031 730
rect 2035 726 2047 730
rect 2051 726 2135 730
rect 2139 726 2151 730
rect 2155 726 2247 730
rect 2251 726 2255 730
rect 2259 726 2359 730
rect 2363 726 2367 730
rect 2371 726 2455 730
rect 2459 726 2503 730
rect 2507 726 2539 730
rect 1317 725 2539 726
rect 2545 725 2546 731
rect 96 701 97 707
rect 103 706 1311 707
rect 103 702 111 706
rect 115 702 151 706
rect 155 702 207 706
rect 211 702 271 706
rect 275 702 295 706
rect 299 702 391 706
rect 395 702 407 706
rect 411 702 503 706
rect 507 702 535 706
rect 539 702 623 706
rect 627 702 663 706
rect 667 702 743 706
rect 747 702 791 706
rect 795 702 871 706
rect 875 702 919 706
rect 923 702 999 706
rect 1003 702 1055 706
rect 1059 702 1127 706
rect 1131 702 1239 706
rect 1243 702 1287 706
rect 1291 702 1311 706
rect 103 701 1311 702
rect 1317 701 1318 707
rect 1298 661 1299 667
rect 1305 666 2527 667
rect 1305 662 1327 666
rect 1331 662 1351 666
rect 1355 662 1415 666
rect 1419 662 1511 666
rect 1515 662 1607 666
rect 1611 662 1615 666
rect 1619 662 1711 666
rect 1715 662 1719 666
rect 1723 662 1823 666
rect 1827 662 1927 666
rect 1931 662 1935 666
rect 1939 662 2031 666
rect 2035 662 2055 666
rect 2059 662 2135 666
rect 2139 662 2183 666
rect 2187 662 2239 666
rect 2243 662 2319 666
rect 2323 662 2351 666
rect 2355 662 2439 666
rect 2443 662 2503 666
rect 2507 662 2527 666
rect 1305 661 2527 662
rect 2533 661 2534 667
rect 84 645 85 651
rect 91 650 1299 651
rect 91 646 111 650
rect 115 646 135 650
rect 139 646 151 650
rect 155 646 191 650
rect 195 646 263 650
rect 267 646 279 650
rect 283 646 367 650
rect 371 646 375 650
rect 379 646 463 650
rect 467 646 487 650
rect 491 646 559 650
rect 563 646 607 650
rect 611 646 655 650
rect 659 646 727 650
rect 731 646 751 650
rect 755 646 847 650
rect 851 646 855 650
rect 859 646 943 650
rect 947 646 983 650
rect 987 646 1039 650
rect 1043 646 1111 650
rect 1115 646 1143 650
rect 1147 646 1223 650
rect 1227 646 1287 650
rect 1291 646 1299 650
rect 91 645 1299 646
rect 1305 645 1306 651
rect 1310 609 1311 615
rect 1317 614 2539 615
rect 1317 610 1327 614
rect 1331 610 1367 614
rect 1371 610 1383 614
rect 1387 610 1431 614
rect 1435 610 1463 614
rect 1467 610 1527 614
rect 1531 610 1551 614
rect 1555 610 1623 614
rect 1627 610 1647 614
rect 1651 610 1727 614
rect 1731 610 1743 614
rect 1747 610 1839 614
rect 1843 610 1847 614
rect 1851 610 1951 614
rect 1955 610 1959 614
rect 1963 610 2071 614
rect 2075 610 2079 614
rect 2083 610 2199 614
rect 2203 610 2207 614
rect 2211 610 2335 614
rect 2339 610 2343 614
rect 2347 610 2455 614
rect 2459 610 2503 614
rect 2507 610 2539 614
rect 1317 609 2539 610
rect 2545 609 2546 615
rect 96 593 97 599
rect 103 598 1311 599
rect 103 594 111 598
rect 115 594 151 598
rect 155 594 167 598
rect 171 594 239 598
rect 243 594 279 598
rect 283 594 335 598
rect 339 594 383 598
rect 387 594 431 598
rect 435 594 479 598
rect 483 594 535 598
rect 539 594 575 598
rect 579 594 631 598
rect 635 594 671 598
rect 675 594 727 598
rect 731 594 767 598
rect 771 594 823 598
rect 827 594 863 598
rect 867 594 911 598
rect 915 594 959 598
rect 963 594 999 598
rect 1003 594 1055 598
rect 1059 594 1087 598
rect 1091 594 1159 598
rect 1163 594 1183 598
rect 1187 594 1239 598
rect 1243 594 1287 598
rect 1291 594 1311 598
rect 103 593 1311 594
rect 1317 593 1318 599
rect 1298 557 1299 563
rect 1305 562 2527 563
rect 1305 558 1327 562
rect 1331 558 1367 562
rect 1371 558 1375 562
rect 1379 558 1447 562
rect 1451 558 1455 562
rect 1459 558 1535 562
rect 1539 558 1551 562
rect 1555 558 1631 562
rect 1635 558 1647 562
rect 1651 558 1727 562
rect 1731 558 1751 562
rect 1755 558 1831 562
rect 1835 558 1855 562
rect 1859 558 1943 562
rect 1947 558 1959 562
rect 1963 558 2055 562
rect 2059 558 2063 562
rect 2067 558 2151 562
rect 2155 558 2191 562
rect 2195 558 2255 562
rect 2259 558 2327 562
rect 2331 558 2359 562
rect 2363 558 2439 562
rect 2443 558 2503 562
rect 2507 558 2527 562
rect 1305 557 2527 558
rect 2533 557 2534 563
rect 84 533 85 539
rect 91 538 1299 539
rect 91 534 111 538
rect 115 534 135 538
rect 139 534 143 538
rect 147 534 223 538
rect 227 534 239 538
rect 243 534 319 538
rect 323 534 335 538
rect 339 534 415 538
rect 419 534 431 538
rect 435 534 519 538
rect 523 534 527 538
rect 531 534 615 538
rect 619 534 623 538
rect 627 534 711 538
rect 715 534 791 538
rect 795 534 807 538
rect 811 534 871 538
rect 875 534 895 538
rect 899 534 951 538
rect 955 534 983 538
rect 987 534 1031 538
rect 1035 534 1071 538
rect 1075 534 1167 538
rect 1171 534 1287 538
rect 1291 534 1299 538
rect 91 533 1299 534
rect 1305 533 1306 539
rect 1310 501 1311 507
rect 1317 506 2539 507
rect 1317 502 1327 506
rect 1331 502 1367 506
rect 1371 502 1391 506
rect 1395 502 1455 506
rect 1459 502 1471 506
rect 1475 502 1567 506
rect 1571 502 1575 506
rect 1579 502 1663 506
rect 1667 502 1695 506
rect 1699 502 1767 506
rect 1771 502 1807 506
rect 1811 502 1871 506
rect 1875 502 1919 506
rect 1923 502 1975 506
rect 1979 502 2023 506
rect 2027 502 2071 506
rect 2075 502 2119 506
rect 2123 502 2167 506
rect 2171 502 2207 506
rect 2211 502 2271 506
rect 2275 502 2295 506
rect 2299 502 2375 506
rect 2379 502 2383 506
rect 2387 502 2455 506
rect 2459 502 2503 506
rect 2507 502 2539 506
rect 1317 501 2539 502
rect 2545 501 2546 507
rect 96 477 97 483
rect 103 482 1311 483
rect 103 478 111 482
rect 115 478 151 482
rect 155 478 159 482
rect 163 478 207 482
rect 211 478 255 482
rect 259 478 287 482
rect 291 478 351 482
rect 355 478 375 482
rect 379 478 447 482
rect 451 478 463 482
rect 467 478 543 482
rect 547 478 559 482
rect 563 478 639 482
rect 643 478 655 482
rect 659 478 727 482
rect 731 478 751 482
rect 755 478 807 482
rect 811 478 847 482
rect 851 478 887 482
rect 891 478 951 482
rect 955 478 967 482
rect 971 478 1047 482
rect 1051 478 1055 482
rect 1059 478 1159 482
rect 1163 478 1239 482
rect 1243 478 1287 482
rect 1291 478 1311 482
rect 103 477 1311 478
rect 1317 477 1318 483
rect 1298 437 1299 443
rect 1305 442 2527 443
rect 1305 438 1327 442
rect 1331 438 1351 442
rect 1355 438 1439 442
rect 1443 438 1559 442
rect 1563 438 1583 442
rect 1587 438 1639 442
rect 1643 438 1679 442
rect 1683 438 1695 442
rect 1699 438 1759 442
rect 1763 438 1791 442
rect 1795 438 1831 442
rect 1835 438 1903 442
rect 1907 438 1911 442
rect 1915 438 1991 442
rect 1995 438 2007 442
rect 2011 438 2079 442
rect 2083 438 2103 442
rect 2107 438 2175 442
rect 2179 438 2191 442
rect 2195 438 2271 442
rect 2275 438 2279 442
rect 2283 438 2367 442
rect 2371 438 2439 442
rect 2443 438 2503 442
rect 2507 438 2527 442
rect 1305 437 2527 438
rect 2533 437 2534 443
rect 84 425 85 431
rect 91 430 1299 431
rect 91 426 111 430
rect 115 426 135 430
rect 139 426 191 430
rect 195 426 271 430
rect 275 426 279 430
rect 283 426 359 430
rect 363 426 383 430
rect 387 426 447 430
rect 451 426 495 430
rect 499 426 543 430
rect 547 426 607 430
rect 611 426 639 430
rect 643 426 719 430
rect 723 426 735 430
rect 739 426 831 430
rect 835 426 935 430
rect 939 426 1039 430
rect 1043 426 1143 430
rect 1147 426 1223 430
rect 1227 426 1287 430
rect 1291 426 1299 430
rect 91 425 1299 426
rect 1305 425 1306 431
rect 1310 381 1311 387
rect 1317 386 2539 387
rect 1317 382 1327 386
rect 1331 382 1599 386
rect 1603 382 1655 386
rect 1659 382 1679 386
rect 1683 382 1711 386
rect 1715 382 1735 386
rect 1739 382 1775 386
rect 1779 382 1799 386
rect 1803 382 1847 386
rect 1851 382 1871 386
rect 1875 382 1927 386
rect 1931 382 1943 386
rect 1947 382 2007 386
rect 2011 382 2023 386
rect 2027 382 2095 386
rect 2099 382 2111 386
rect 2115 382 2191 386
rect 2195 382 2199 386
rect 2203 382 2287 386
rect 2291 382 2375 386
rect 2379 382 2383 386
rect 2387 382 2455 386
rect 2459 382 2503 386
rect 2507 382 2539 386
rect 1317 381 2539 382
rect 2545 381 2546 387
rect 96 369 97 375
rect 103 374 1311 375
rect 103 370 111 374
rect 115 370 151 374
rect 155 370 207 374
rect 211 370 231 374
rect 235 370 295 374
rect 299 370 335 374
rect 339 370 399 374
rect 403 370 439 374
rect 443 370 511 374
rect 515 370 543 374
rect 547 370 623 374
rect 627 370 647 374
rect 651 370 735 374
rect 739 370 751 374
rect 755 370 847 374
rect 851 370 935 374
rect 939 370 951 374
rect 955 370 1015 374
rect 1019 370 1055 374
rect 1059 370 1095 374
rect 1099 370 1159 374
rect 1163 370 1175 374
rect 1179 370 1239 374
rect 1243 370 1287 374
rect 1291 370 1311 374
rect 103 369 1311 370
rect 1317 369 1318 375
rect 1298 321 1299 327
rect 1305 326 2527 327
rect 1305 322 1327 326
rect 1331 322 1351 326
rect 1355 322 1455 326
rect 1459 322 1583 326
rect 1587 322 1663 326
rect 1667 322 1711 326
rect 1715 322 1719 326
rect 1723 322 1783 326
rect 1787 322 1839 326
rect 1843 322 1855 326
rect 1859 322 1927 326
rect 1931 322 1951 326
rect 1955 322 2007 326
rect 2011 322 2063 326
rect 2067 322 2095 326
rect 2099 322 2167 326
rect 2171 322 2183 326
rect 2187 322 2263 326
rect 2267 322 2271 326
rect 2275 322 2359 326
rect 2363 322 2439 326
rect 2443 322 2503 326
rect 2507 322 2527 326
rect 1305 321 2527 322
rect 2533 321 2534 327
rect 1298 319 1306 321
rect 84 313 85 319
rect 91 318 1299 319
rect 91 314 111 318
rect 115 314 135 318
rect 139 314 215 318
rect 219 314 319 318
rect 323 314 423 318
rect 427 314 527 318
rect 531 314 535 318
rect 539 314 631 318
rect 635 314 639 318
rect 643 314 735 318
rect 739 314 743 318
rect 747 314 831 318
rect 835 314 847 318
rect 851 314 919 318
rect 923 314 943 318
rect 947 314 999 318
rect 1003 314 1039 318
rect 1043 314 1079 318
rect 1083 314 1143 318
rect 1147 314 1159 318
rect 1163 314 1223 318
rect 1227 314 1287 318
rect 1291 314 1299 318
rect 91 313 1299 314
rect 1305 313 1306 319
rect 96 261 97 267
rect 103 266 1311 267
rect 103 262 111 266
rect 115 262 151 266
rect 155 262 223 266
rect 227 262 231 266
rect 235 262 319 266
rect 323 262 335 266
rect 339 262 423 266
rect 427 262 439 266
rect 443 262 535 266
rect 539 262 551 266
rect 555 262 647 266
rect 651 262 655 266
rect 659 262 759 266
rect 763 262 863 266
rect 867 262 871 266
rect 875 262 959 266
rect 963 262 983 266
rect 987 262 1055 266
rect 1059 262 1103 266
rect 1107 262 1159 266
rect 1163 262 1223 266
rect 1227 262 1239 266
rect 1243 262 1287 266
rect 1291 262 1311 266
rect 103 261 1311 262
rect 1317 266 2546 267
rect 1317 262 1327 266
rect 1331 262 1367 266
rect 1371 262 1447 266
rect 1451 262 1471 266
rect 1475 262 1551 266
rect 1555 262 1599 266
rect 1603 262 1655 266
rect 1659 262 1727 266
rect 1731 262 1759 266
rect 1763 262 1855 266
rect 1859 262 1863 266
rect 1867 262 1967 266
rect 1971 262 2071 266
rect 2075 262 2079 266
rect 2083 262 2175 266
rect 2179 262 2183 266
rect 2187 262 2271 266
rect 2275 262 2279 266
rect 2283 262 2375 266
rect 2379 262 2455 266
rect 2459 262 2503 266
rect 2507 262 2546 266
rect 1317 261 2546 262
rect 84 205 85 211
rect 91 210 1299 211
rect 91 206 111 210
rect 115 206 135 210
rect 139 206 183 210
rect 187 206 207 210
rect 211 206 279 210
rect 283 206 303 210
rect 307 206 383 210
rect 387 206 407 210
rect 411 206 487 210
rect 491 206 519 210
rect 523 206 591 210
rect 595 206 631 210
rect 635 206 695 210
rect 699 206 743 210
rect 747 206 799 210
rect 803 206 855 210
rect 859 206 895 210
rect 899 206 967 210
rect 971 206 999 210
rect 1003 206 1087 210
rect 1091 206 1103 210
rect 1107 206 1207 210
rect 1211 206 1287 210
rect 1291 206 1299 210
rect 91 205 1299 206
rect 1305 210 2534 211
rect 1305 206 1327 210
rect 1331 206 1351 210
rect 1355 206 1407 210
rect 1411 206 1431 210
rect 1435 206 1471 210
rect 1475 206 1535 210
rect 1539 206 1551 210
rect 1555 206 1639 210
rect 1643 206 1719 210
rect 1723 206 1743 210
rect 1747 206 1807 210
rect 1811 206 1847 210
rect 1851 206 1895 210
rect 1899 206 1951 210
rect 1955 206 1991 210
rect 1995 206 2055 210
rect 2059 206 2103 210
rect 2107 206 2159 210
rect 2163 206 2215 210
rect 2219 206 2255 210
rect 2259 206 2335 210
rect 2339 206 2359 210
rect 2363 206 2439 210
rect 2443 206 2503 210
rect 2507 206 2534 210
rect 1305 205 2534 206
rect 96 145 97 151
rect 103 150 1311 151
rect 103 146 111 150
rect 115 146 151 150
rect 155 146 199 150
rect 203 146 207 150
rect 211 146 263 150
rect 267 146 295 150
rect 299 146 319 150
rect 323 146 375 150
rect 379 146 399 150
rect 403 146 431 150
rect 435 146 487 150
rect 491 146 503 150
rect 507 146 543 150
rect 547 146 599 150
rect 603 146 607 150
rect 611 146 655 150
rect 659 146 711 150
rect 715 146 767 150
rect 771 146 815 150
rect 819 146 831 150
rect 835 146 895 150
rect 899 146 911 150
rect 915 146 959 150
rect 963 146 1015 150
rect 1019 146 1023 150
rect 1027 146 1087 150
rect 1091 146 1119 150
rect 1123 146 1151 150
rect 1155 146 1287 150
rect 1291 146 1311 150
rect 103 145 1311 146
rect 1317 145 1318 151
rect 1310 133 1311 139
rect 1317 138 2539 139
rect 1317 134 1327 138
rect 1331 134 1367 138
rect 1371 134 1423 138
rect 1427 134 1479 138
rect 1483 134 1487 138
rect 1491 134 1535 138
rect 1539 134 1567 138
rect 1571 134 1591 138
rect 1595 134 1647 138
rect 1651 134 1655 138
rect 1659 134 1703 138
rect 1707 134 1735 138
rect 1739 134 1759 138
rect 1763 134 1823 138
rect 1827 134 1879 138
rect 1883 134 1911 138
rect 1915 134 1943 138
rect 1947 134 2007 138
rect 2011 134 2071 138
rect 2075 134 2119 138
rect 2123 134 2143 138
rect 2147 134 2223 138
rect 2227 134 2231 138
rect 2235 134 2303 138
rect 2307 134 2351 138
rect 2355 134 2391 138
rect 2395 134 2455 138
rect 2459 134 2503 138
rect 2507 134 2539 138
rect 1317 133 2539 134
rect 2545 133 2546 139
rect 84 93 85 99
rect 91 98 1299 99
rect 91 94 111 98
rect 115 94 135 98
rect 139 94 191 98
rect 195 94 247 98
rect 251 94 303 98
rect 307 94 359 98
rect 363 94 415 98
rect 419 94 471 98
rect 475 94 527 98
rect 531 94 583 98
rect 587 94 639 98
rect 643 94 695 98
rect 699 94 751 98
rect 755 94 815 98
rect 819 94 879 98
rect 883 94 943 98
rect 947 94 1007 98
rect 1011 94 1071 98
rect 1075 94 1135 98
rect 1139 94 1287 98
rect 1291 94 1299 98
rect 91 93 1299 94
rect 1305 93 1306 99
rect 1298 81 1299 87
rect 1305 86 2527 87
rect 1305 82 1327 86
rect 1331 82 1351 86
rect 1355 82 1407 86
rect 1411 82 1463 86
rect 1467 82 1519 86
rect 1523 82 1575 86
rect 1579 82 1631 86
rect 1635 82 1687 86
rect 1691 82 1743 86
rect 1747 82 1807 86
rect 1811 82 1863 86
rect 1867 82 1927 86
rect 1931 82 1991 86
rect 1995 82 2055 86
rect 2059 82 2127 86
rect 2131 82 2207 86
rect 2211 82 2287 86
rect 2291 82 2375 86
rect 2379 82 2439 86
rect 2443 82 2503 86
rect 2507 82 2527 86
rect 1305 81 2527 82
rect 2533 81 2534 87
<< m5c >>
rect 85 2577 91 2583
rect 1299 2577 1305 2583
rect 1299 2557 1305 2563
rect 2527 2557 2533 2563
rect 97 2525 103 2531
rect 1311 2525 1317 2531
rect 1311 2505 1317 2511
rect 2539 2505 2545 2511
rect 85 2465 91 2471
rect 1299 2465 1305 2471
rect 1299 2449 1305 2455
rect 2527 2449 2533 2455
rect 97 2401 103 2407
rect 1311 2401 1317 2407
rect 1311 2393 1317 2399
rect 2539 2393 2545 2399
rect 85 2341 91 2347
rect 1299 2341 1305 2347
rect 1299 2333 1305 2339
rect 2527 2333 2533 2339
rect 97 2281 103 2287
rect 1311 2281 1317 2287
rect 85 2229 91 2235
rect 1299 2229 1305 2235
rect 97 2177 103 2183
rect 1311 2177 1317 2183
rect 1311 2157 1317 2163
rect 2539 2157 2545 2163
rect 85 2125 91 2131
rect 1299 2125 1305 2131
rect 1299 2105 1305 2111
rect 2527 2105 2533 2111
rect 97 2069 103 2075
rect 1311 2069 1317 2075
rect 1311 2049 1317 2055
rect 2539 2049 2545 2055
rect 85 2013 91 2019
rect 1299 2013 1305 2019
rect 1299 1993 1305 1999
rect 2527 1993 2533 1999
rect 97 1957 103 1963
rect 1311 1957 1317 1963
rect 1311 1937 1317 1943
rect 2539 1937 2545 1943
rect 85 1897 91 1903
rect 1299 1897 1305 1903
rect 1299 1881 1305 1887
rect 2527 1881 2533 1887
rect 97 1845 103 1851
rect 1311 1845 1317 1851
rect 1311 1825 1317 1831
rect 2539 1825 2545 1831
rect 85 1781 91 1787
rect 1299 1781 1305 1787
rect 1299 1773 1305 1779
rect 2527 1773 2533 1779
rect 97 1725 103 1731
rect 1311 1725 1317 1731
rect 1311 1717 1317 1723
rect 2539 1717 2545 1723
rect 85 1669 91 1675
rect 1299 1669 1305 1675
rect 1299 1661 1305 1667
rect 2527 1661 2533 1667
rect 97 1613 103 1619
rect 1311 1613 1317 1619
rect 85 1561 91 1567
rect 1299 1561 1305 1567
rect 97 1501 103 1507
rect 1311 1501 1317 1507
rect 85 1445 91 1451
rect 1299 1445 1305 1451
rect 97 1389 103 1395
rect 1311 1389 1317 1395
rect 1299 1341 1305 1347
rect 2527 1341 2533 1347
rect 85 1321 91 1327
rect 1299 1321 1305 1327
rect 1311 1289 1317 1295
rect 2539 1289 2545 1295
rect 97 1261 103 1267
rect 1311 1261 1317 1267
rect 1299 1233 1305 1239
rect 2527 1233 2533 1239
rect 85 1205 91 1211
rect 1299 1205 1305 1211
rect 1311 1177 1317 1183
rect 2539 1177 2545 1183
rect 97 1149 103 1155
rect 1311 1149 1317 1155
rect 1299 1125 1305 1131
rect 2527 1125 2533 1131
rect 85 1089 91 1095
rect 1299 1089 1305 1095
rect 1311 1065 1317 1071
rect 2539 1065 2545 1071
rect 97 1029 103 1035
rect 1311 1029 1317 1035
rect 1299 1009 1305 1015
rect 2527 1009 2533 1015
rect 85 977 91 983
rect 1299 977 1305 983
rect 1311 945 1317 951
rect 2539 945 2545 951
rect 97 917 103 923
rect 1311 917 1317 923
rect 1299 889 1305 895
rect 2527 889 2533 895
rect 85 861 91 867
rect 1299 861 1305 867
rect 1311 833 1317 839
rect 2539 833 2545 839
rect 97 805 103 811
rect 1311 805 1317 811
rect 1299 777 1305 783
rect 2527 777 2533 783
rect 85 753 91 759
rect 1299 753 1305 759
rect 1311 725 1317 731
rect 2539 725 2545 731
rect 97 701 103 707
rect 1311 701 1317 707
rect 1299 661 1305 667
rect 2527 661 2533 667
rect 85 645 91 651
rect 1299 645 1305 651
rect 1311 609 1317 615
rect 2539 609 2545 615
rect 97 593 103 599
rect 1311 593 1317 599
rect 1299 557 1305 563
rect 2527 557 2533 563
rect 85 533 91 539
rect 1299 533 1305 539
rect 1311 501 1317 507
rect 2539 501 2545 507
rect 97 477 103 483
rect 1311 477 1317 483
rect 1299 437 1305 443
rect 2527 437 2533 443
rect 85 425 91 431
rect 1299 425 1305 431
rect 1311 381 1317 387
rect 2539 381 2545 387
rect 97 369 103 375
rect 1311 369 1317 375
rect 1299 321 1305 327
rect 2527 321 2533 327
rect 85 313 91 319
rect 1299 313 1305 319
rect 97 261 103 267
rect 1311 261 1317 267
rect 85 205 91 211
rect 1299 205 1305 211
rect 97 145 103 151
rect 1311 145 1317 151
rect 1311 133 1317 139
rect 2539 133 2545 139
rect 85 93 91 99
rect 1299 93 1305 99
rect 1299 81 1305 87
rect 2527 81 2533 87
<< m5 >>
rect 84 2583 92 2592
rect 84 2577 85 2583
rect 91 2577 92 2583
rect 84 2471 92 2577
rect 84 2465 85 2471
rect 91 2465 92 2471
rect 84 2347 92 2465
rect 84 2341 85 2347
rect 91 2341 92 2347
rect 84 2235 92 2341
rect 84 2229 85 2235
rect 91 2229 92 2235
rect 84 2131 92 2229
rect 84 2125 85 2131
rect 91 2125 92 2131
rect 84 2019 92 2125
rect 84 2013 85 2019
rect 91 2013 92 2019
rect 84 1903 92 2013
rect 84 1897 85 1903
rect 91 1897 92 1903
rect 84 1787 92 1897
rect 84 1781 85 1787
rect 91 1781 92 1787
rect 84 1675 92 1781
rect 84 1669 85 1675
rect 91 1669 92 1675
rect 84 1567 92 1669
rect 84 1561 85 1567
rect 91 1561 92 1567
rect 84 1451 92 1561
rect 84 1445 85 1451
rect 91 1445 92 1451
rect 84 1327 92 1445
rect 84 1321 85 1327
rect 91 1321 92 1327
rect 84 1211 92 1321
rect 84 1205 85 1211
rect 91 1205 92 1211
rect 84 1095 92 1205
rect 84 1089 85 1095
rect 91 1089 92 1095
rect 84 983 92 1089
rect 84 977 85 983
rect 91 977 92 983
rect 84 867 92 977
rect 84 861 85 867
rect 91 861 92 867
rect 84 759 92 861
rect 84 753 85 759
rect 91 753 92 759
rect 84 651 92 753
rect 84 645 85 651
rect 91 645 92 651
rect 84 539 92 645
rect 84 533 85 539
rect 91 533 92 539
rect 84 431 92 533
rect 84 425 85 431
rect 91 425 92 431
rect 84 319 92 425
rect 84 313 85 319
rect 91 313 92 319
rect 84 211 92 313
rect 84 205 85 211
rect 91 205 92 211
rect 84 99 92 205
rect 84 93 85 99
rect 91 93 92 99
rect 84 72 92 93
rect 96 2531 104 2592
rect 96 2525 97 2531
rect 103 2525 104 2531
rect 96 2407 104 2525
rect 96 2401 97 2407
rect 103 2401 104 2407
rect 96 2287 104 2401
rect 96 2281 97 2287
rect 103 2281 104 2287
rect 96 2183 104 2281
rect 96 2177 97 2183
rect 103 2177 104 2183
rect 96 2075 104 2177
rect 96 2069 97 2075
rect 103 2069 104 2075
rect 96 1963 104 2069
rect 96 1957 97 1963
rect 103 1957 104 1963
rect 96 1851 104 1957
rect 96 1845 97 1851
rect 103 1845 104 1851
rect 96 1731 104 1845
rect 96 1725 97 1731
rect 103 1725 104 1731
rect 96 1619 104 1725
rect 96 1613 97 1619
rect 103 1613 104 1619
rect 96 1507 104 1613
rect 96 1501 97 1507
rect 103 1501 104 1507
rect 96 1395 104 1501
rect 96 1389 97 1395
rect 103 1389 104 1395
rect 96 1267 104 1389
rect 96 1261 97 1267
rect 103 1261 104 1267
rect 96 1155 104 1261
rect 96 1149 97 1155
rect 103 1149 104 1155
rect 96 1035 104 1149
rect 96 1029 97 1035
rect 103 1029 104 1035
rect 96 923 104 1029
rect 96 917 97 923
rect 103 917 104 923
rect 96 811 104 917
rect 96 805 97 811
rect 103 805 104 811
rect 96 707 104 805
rect 96 701 97 707
rect 103 701 104 707
rect 96 599 104 701
rect 96 593 97 599
rect 103 593 104 599
rect 96 483 104 593
rect 96 477 97 483
rect 103 477 104 483
rect 96 375 104 477
rect 96 369 97 375
rect 103 369 104 375
rect 96 267 104 369
rect 96 261 97 267
rect 103 261 104 267
rect 96 151 104 261
rect 96 145 97 151
rect 103 145 104 151
rect 96 72 104 145
rect 1298 2583 1306 2592
rect 1298 2577 1299 2583
rect 1305 2577 1306 2583
rect 1298 2563 1306 2577
rect 1298 2557 1299 2563
rect 1305 2557 1306 2563
rect 1298 2471 1306 2557
rect 1298 2465 1299 2471
rect 1305 2465 1306 2471
rect 1298 2455 1306 2465
rect 1298 2449 1299 2455
rect 1305 2449 1306 2455
rect 1298 2347 1306 2449
rect 1298 2341 1299 2347
rect 1305 2341 1306 2347
rect 1298 2339 1306 2341
rect 1298 2333 1299 2339
rect 1305 2333 1306 2339
rect 1298 2235 1306 2333
rect 1298 2229 1299 2235
rect 1305 2229 1306 2235
rect 1298 2131 1306 2229
rect 1298 2125 1299 2131
rect 1305 2125 1306 2131
rect 1298 2111 1306 2125
rect 1298 2105 1299 2111
rect 1305 2105 1306 2111
rect 1298 2019 1306 2105
rect 1298 2013 1299 2019
rect 1305 2013 1306 2019
rect 1298 1999 1306 2013
rect 1298 1993 1299 1999
rect 1305 1993 1306 1999
rect 1298 1903 1306 1993
rect 1298 1897 1299 1903
rect 1305 1897 1306 1903
rect 1298 1887 1306 1897
rect 1298 1881 1299 1887
rect 1305 1881 1306 1887
rect 1298 1787 1306 1881
rect 1298 1781 1299 1787
rect 1305 1781 1306 1787
rect 1298 1779 1306 1781
rect 1298 1773 1299 1779
rect 1305 1773 1306 1779
rect 1298 1675 1306 1773
rect 1298 1669 1299 1675
rect 1305 1669 1306 1675
rect 1298 1667 1306 1669
rect 1298 1661 1299 1667
rect 1305 1661 1306 1667
rect 1298 1567 1306 1661
rect 1298 1561 1299 1567
rect 1305 1561 1306 1567
rect 1298 1451 1306 1561
rect 1298 1445 1299 1451
rect 1305 1445 1306 1451
rect 1298 1347 1306 1445
rect 1298 1341 1299 1347
rect 1305 1341 1306 1347
rect 1298 1327 1306 1341
rect 1298 1321 1299 1327
rect 1305 1321 1306 1327
rect 1298 1239 1306 1321
rect 1298 1233 1299 1239
rect 1305 1233 1306 1239
rect 1298 1211 1306 1233
rect 1298 1205 1299 1211
rect 1305 1205 1306 1211
rect 1298 1131 1306 1205
rect 1298 1125 1299 1131
rect 1305 1125 1306 1131
rect 1298 1095 1306 1125
rect 1298 1089 1299 1095
rect 1305 1089 1306 1095
rect 1298 1015 1306 1089
rect 1298 1009 1299 1015
rect 1305 1009 1306 1015
rect 1298 983 1306 1009
rect 1298 977 1299 983
rect 1305 977 1306 983
rect 1298 895 1306 977
rect 1298 889 1299 895
rect 1305 889 1306 895
rect 1298 867 1306 889
rect 1298 861 1299 867
rect 1305 861 1306 867
rect 1298 783 1306 861
rect 1298 777 1299 783
rect 1305 777 1306 783
rect 1298 759 1306 777
rect 1298 753 1299 759
rect 1305 753 1306 759
rect 1298 667 1306 753
rect 1298 661 1299 667
rect 1305 661 1306 667
rect 1298 651 1306 661
rect 1298 645 1299 651
rect 1305 645 1306 651
rect 1298 563 1306 645
rect 1298 557 1299 563
rect 1305 557 1306 563
rect 1298 539 1306 557
rect 1298 533 1299 539
rect 1305 533 1306 539
rect 1298 443 1306 533
rect 1298 437 1299 443
rect 1305 437 1306 443
rect 1298 431 1306 437
rect 1298 425 1299 431
rect 1305 425 1306 431
rect 1298 327 1306 425
rect 1298 321 1299 327
rect 1305 321 1306 327
rect 1298 319 1306 321
rect 1298 313 1299 319
rect 1305 313 1306 319
rect 1298 211 1306 313
rect 1298 205 1299 211
rect 1305 205 1306 211
rect 1298 99 1306 205
rect 1298 93 1299 99
rect 1305 93 1306 99
rect 1298 87 1306 93
rect 1298 81 1299 87
rect 1305 81 1306 87
rect 1298 72 1306 81
rect 1310 2531 1318 2592
rect 1310 2525 1311 2531
rect 1317 2525 1318 2531
rect 1310 2511 1318 2525
rect 1310 2505 1311 2511
rect 1317 2505 1318 2511
rect 1310 2407 1318 2505
rect 1310 2401 1311 2407
rect 1317 2401 1318 2407
rect 1310 2399 1318 2401
rect 1310 2393 1311 2399
rect 1317 2393 1318 2399
rect 1310 2287 1318 2393
rect 1310 2281 1311 2287
rect 1317 2281 1318 2287
rect 1310 2183 1318 2281
rect 1310 2177 1311 2183
rect 1317 2177 1318 2183
rect 1310 2163 1318 2177
rect 1310 2157 1311 2163
rect 1317 2157 1318 2163
rect 1310 2075 1318 2157
rect 1310 2069 1311 2075
rect 1317 2069 1318 2075
rect 1310 2055 1318 2069
rect 1310 2049 1311 2055
rect 1317 2049 1318 2055
rect 1310 1963 1318 2049
rect 1310 1957 1311 1963
rect 1317 1957 1318 1963
rect 1310 1943 1318 1957
rect 1310 1937 1311 1943
rect 1317 1937 1318 1943
rect 1310 1851 1318 1937
rect 1310 1845 1311 1851
rect 1317 1845 1318 1851
rect 1310 1831 1318 1845
rect 1310 1825 1311 1831
rect 1317 1825 1318 1831
rect 1310 1731 1318 1825
rect 1310 1725 1311 1731
rect 1317 1725 1318 1731
rect 1310 1723 1318 1725
rect 1310 1717 1311 1723
rect 1317 1717 1318 1723
rect 1310 1619 1318 1717
rect 1310 1613 1311 1619
rect 1317 1613 1318 1619
rect 1310 1507 1318 1613
rect 1310 1501 1311 1507
rect 1317 1501 1318 1507
rect 1310 1395 1318 1501
rect 1310 1389 1311 1395
rect 1317 1389 1318 1395
rect 1310 1295 1318 1389
rect 1310 1289 1311 1295
rect 1317 1289 1318 1295
rect 1310 1267 1318 1289
rect 1310 1261 1311 1267
rect 1317 1261 1318 1267
rect 1310 1183 1318 1261
rect 1310 1177 1311 1183
rect 1317 1177 1318 1183
rect 1310 1155 1318 1177
rect 1310 1149 1311 1155
rect 1317 1149 1318 1155
rect 1310 1071 1318 1149
rect 1310 1065 1311 1071
rect 1317 1065 1318 1071
rect 1310 1035 1318 1065
rect 1310 1029 1311 1035
rect 1317 1029 1318 1035
rect 1310 951 1318 1029
rect 1310 945 1311 951
rect 1317 945 1318 951
rect 1310 923 1318 945
rect 1310 917 1311 923
rect 1317 917 1318 923
rect 1310 839 1318 917
rect 1310 833 1311 839
rect 1317 833 1318 839
rect 1310 811 1318 833
rect 1310 805 1311 811
rect 1317 805 1318 811
rect 1310 731 1318 805
rect 1310 725 1311 731
rect 1317 725 1318 731
rect 1310 707 1318 725
rect 1310 701 1311 707
rect 1317 701 1318 707
rect 1310 615 1318 701
rect 1310 609 1311 615
rect 1317 609 1318 615
rect 1310 599 1318 609
rect 1310 593 1311 599
rect 1317 593 1318 599
rect 1310 507 1318 593
rect 1310 501 1311 507
rect 1317 501 1318 507
rect 1310 483 1318 501
rect 1310 477 1311 483
rect 1317 477 1318 483
rect 1310 387 1318 477
rect 1310 381 1311 387
rect 1317 381 1318 387
rect 1310 375 1318 381
rect 1310 369 1311 375
rect 1317 369 1318 375
rect 1310 267 1318 369
rect 1310 261 1311 267
rect 1317 261 1318 267
rect 1310 151 1318 261
rect 1310 145 1311 151
rect 1317 145 1318 151
rect 1310 139 1318 145
rect 1310 133 1311 139
rect 1317 133 1318 139
rect 1310 72 1318 133
rect 2526 2563 2534 2592
rect 2526 2557 2527 2563
rect 2533 2557 2534 2563
rect 2526 2455 2534 2557
rect 2526 2449 2527 2455
rect 2533 2449 2534 2455
rect 2526 2339 2534 2449
rect 2526 2333 2527 2339
rect 2533 2333 2534 2339
rect 2526 2111 2534 2333
rect 2526 2105 2527 2111
rect 2533 2105 2534 2111
rect 2526 1999 2534 2105
rect 2526 1993 2527 1999
rect 2533 1993 2534 1999
rect 2526 1887 2534 1993
rect 2526 1881 2527 1887
rect 2533 1881 2534 1887
rect 2526 1779 2534 1881
rect 2526 1773 2527 1779
rect 2533 1773 2534 1779
rect 2526 1667 2534 1773
rect 2526 1661 2527 1667
rect 2533 1661 2534 1667
rect 2526 1347 2534 1661
rect 2526 1341 2527 1347
rect 2533 1341 2534 1347
rect 2526 1239 2534 1341
rect 2526 1233 2527 1239
rect 2533 1233 2534 1239
rect 2526 1131 2534 1233
rect 2526 1125 2527 1131
rect 2533 1125 2534 1131
rect 2526 1015 2534 1125
rect 2526 1009 2527 1015
rect 2533 1009 2534 1015
rect 2526 895 2534 1009
rect 2526 889 2527 895
rect 2533 889 2534 895
rect 2526 783 2534 889
rect 2526 777 2527 783
rect 2533 777 2534 783
rect 2526 667 2534 777
rect 2526 661 2527 667
rect 2533 661 2534 667
rect 2526 563 2534 661
rect 2526 557 2527 563
rect 2533 557 2534 563
rect 2526 443 2534 557
rect 2526 437 2527 443
rect 2533 437 2534 443
rect 2526 327 2534 437
rect 2526 321 2527 327
rect 2533 321 2534 327
rect 2526 87 2534 321
rect 2526 81 2527 87
rect 2533 81 2534 87
rect 2526 72 2534 81
rect 2538 2511 2546 2592
rect 2538 2505 2539 2511
rect 2545 2505 2546 2511
rect 2538 2399 2546 2505
rect 2538 2393 2539 2399
rect 2545 2393 2546 2399
rect 2538 2163 2546 2393
rect 2538 2157 2539 2163
rect 2545 2157 2546 2163
rect 2538 2055 2546 2157
rect 2538 2049 2539 2055
rect 2545 2049 2546 2055
rect 2538 1943 2546 2049
rect 2538 1937 2539 1943
rect 2545 1937 2546 1943
rect 2538 1831 2546 1937
rect 2538 1825 2539 1831
rect 2545 1825 2546 1831
rect 2538 1723 2546 1825
rect 2538 1717 2539 1723
rect 2545 1717 2546 1723
rect 2538 1295 2546 1717
rect 2538 1289 2539 1295
rect 2545 1289 2546 1295
rect 2538 1183 2546 1289
rect 2538 1177 2539 1183
rect 2545 1177 2546 1183
rect 2538 1071 2546 1177
rect 2538 1065 2539 1071
rect 2545 1065 2546 1071
rect 2538 951 2546 1065
rect 2538 945 2539 951
rect 2545 945 2546 951
rect 2538 839 2546 945
rect 2538 833 2539 839
rect 2545 833 2546 839
rect 2538 731 2546 833
rect 2538 725 2539 731
rect 2545 725 2546 731
rect 2538 615 2546 725
rect 2538 609 2539 615
rect 2545 609 2546 615
rect 2538 507 2546 609
rect 2538 501 2539 507
rect 2545 501 2546 507
rect 2538 387 2546 501
rect 2538 381 2539 387
rect 2545 381 2546 387
rect 2538 139 2546 381
rect 2538 133 2539 139
rect 2545 133 2546 139
rect 2538 72 2546 133
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__175
timestamp 1731220673
transform 1 0 2496 0 -1 2556
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220673
transform 1 0 1320 0 -1 2556
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220673
transform 1 0 2496 0 1 2460
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220673
transform 1 0 1320 0 1 2460
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220673
transform 1 0 2496 0 -1 2448
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220673
transform 1 0 1320 0 -1 2448
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220673
transform 1 0 2496 0 1 2348
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220673
transform 1 0 1320 0 1 2348
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220673
transform 1 0 2496 0 -1 2332
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220673
transform 1 0 1320 0 -1 2332
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220673
transform 1 0 2496 0 1 2236
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220673
transform 1 0 1320 0 1 2236
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220673
transform 1 0 2496 0 -1 2228
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220673
transform 1 0 1320 0 -1 2228
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220673
transform 1 0 2496 0 1 2112
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220673
transform 1 0 1320 0 1 2112
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220673
transform 1 0 2496 0 -1 2104
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220673
transform 1 0 1320 0 -1 2104
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220673
transform 1 0 2496 0 1 2004
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220673
transform 1 0 1320 0 1 2004
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220673
transform 1 0 2496 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220673
transform 1 0 1320 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220673
transform 1 0 2496 0 1 1892
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220673
transform 1 0 1320 0 1 1892
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220673
transform 1 0 2496 0 -1 1880
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220673
transform 1 0 1320 0 -1 1880
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220673
transform 1 0 2496 0 1 1780
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220673
transform 1 0 1320 0 1 1780
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220673
transform 1 0 2496 0 -1 1772
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220673
transform 1 0 1320 0 -1 1772
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220673
transform 1 0 2496 0 1 1672
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220673
transform 1 0 1320 0 1 1672
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220673
transform 1 0 2496 0 -1 1660
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220673
transform 1 0 1320 0 -1 1660
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220673
transform 1 0 2496 0 1 1564
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220673
transform 1 0 1320 0 1 1564
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220673
transform 1 0 2496 0 -1 1556
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220673
transform 1 0 1320 0 -1 1556
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220673
transform 1 0 2496 0 1 1460
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220673
transform 1 0 1320 0 1 1460
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220673
transform 1 0 2496 0 -1 1444
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220673
transform 1 0 1320 0 -1 1444
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220673
transform 1 0 2496 0 1 1348
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220673
transform 1 0 1320 0 1 1348
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220673
transform 1 0 2496 0 -1 1340
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220673
transform 1 0 1320 0 -1 1340
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220673
transform 1 0 2496 0 1 1244
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220673
transform 1 0 1320 0 1 1244
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220673
transform 1 0 2496 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220673
transform 1 0 1320 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220673
transform 1 0 2496 0 1 1132
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220673
transform 1 0 1320 0 1 1132
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220673
transform 1 0 2496 0 -1 1124
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220673
transform 1 0 1320 0 -1 1124
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220673
transform 1 0 2496 0 1 1020
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220673
transform 1 0 1320 0 1 1020
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220673
transform 1 0 2496 0 -1 1008
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220673
transform 1 0 1320 0 -1 1008
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220673
transform 1 0 2496 0 1 900
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220673
transform 1 0 1320 0 1 900
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220673
transform 1 0 2496 0 -1 888
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220673
transform 1 0 1320 0 -1 888
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220673
transform 1 0 2496 0 1 788
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220673
transform 1 0 1320 0 1 788
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220673
transform 1 0 2496 0 -1 776
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220673
transform 1 0 1320 0 -1 776
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220673
transform 1 0 2496 0 1 680
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220673
transform 1 0 1320 0 1 680
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220673
transform 1 0 2496 0 -1 660
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220673
transform 1 0 1320 0 -1 660
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220673
transform 1 0 2496 0 1 564
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220673
transform 1 0 1320 0 1 564
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220673
transform 1 0 2496 0 -1 556
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220673
transform 1 0 1320 0 -1 556
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220673
transform 1 0 2496 0 1 456
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220673
transform 1 0 1320 0 1 456
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220673
transform 1 0 2496 0 -1 436
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220673
transform 1 0 1320 0 -1 436
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220673
transform 1 0 2496 0 1 336
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220673
transform 1 0 1320 0 1 336
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220673
transform 1 0 2496 0 -1 320
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220673
transform 1 0 1320 0 -1 320
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220673
transform 1 0 2496 0 1 216
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220673
transform 1 0 1320 0 1 216
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220673
transform 1 0 2496 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220673
transform 1 0 1320 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220673
transform 1 0 2496 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220673
transform 1 0 1320 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220673
transform 1 0 1280 0 -1 2576
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220673
transform 1 0 104 0 -1 2576
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220673
transform 1 0 1280 0 1 2480
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220673
transform 1 0 104 0 1 2480
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220673
transform 1 0 1280 0 -1 2464
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220673
transform 1 0 104 0 -1 2464
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220673
transform 1 0 1280 0 1 2356
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220673
transform 1 0 104 0 1 2356
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220673
transform 1 0 1280 0 -1 2340
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220673
transform 1 0 104 0 -1 2340
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220673
transform 1 0 1280 0 1 2236
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220673
transform 1 0 104 0 1 2236
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220673
transform 1 0 1280 0 -1 2228
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220673
transform 1 0 104 0 -1 2228
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220673
transform 1 0 1280 0 1 2132
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220673
transform 1 0 104 0 1 2132
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220673
transform 1 0 1280 0 -1 2124
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220673
transform 1 0 104 0 -1 2124
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220673
transform 1 0 1280 0 1 2024
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220673
transform 1 0 104 0 1 2024
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220673
transform 1 0 1280 0 -1 2012
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220673
transform 1 0 104 0 -1 2012
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220673
transform 1 0 1280 0 1 1912
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220673
transform 1 0 104 0 1 1912
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220673
transform 1 0 1280 0 -1 1896
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220673
transform 1 0 104 0 -1 1896
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220673
transform 1 0 1280 0 1 1800
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220673
transform 1 0 104 0 1 1800
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220673
transform 1 0 1280 0 -1 1780
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220673
transform 1 0 104 0 -1 1780
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220673
transform 1 0 1280 0 1 1680
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220673
transform 1 0 104 0 1 1680
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220673
transform 1 0 1280 0 -1 1668
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220673
transform 1 0 104 0 -1 1668
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220673
transform 1 0 1280 0 1 1568
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220673
transform 1 0 104 0 1 1568
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220673
transform 1 0 1280 0 -1 1560
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220673
transform 1 0 104 0 -1 1560
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220673
transform 1 0 1280 0 1 1456
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220673
transform 1 0 104 0 1 1456
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220673
transform 1 0 1280 0 -1 1444
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220673
transform 1 0 104 0 -1 1444
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220673
transform 1 0 1280 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220673
transform 1 0 104 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220673
transform 1 0 1280 0 -1 1320
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220673
transform 1 0 104 0 -1 1320
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220673
transform 1 0 1280 0 1 1216
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220673
transform 1 0 104 0 1 1216
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220673
transform 1 0 1280 0 -1 1204
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220673
transform 1 0 104 0 -1 1204
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220673
transform 1 0 1280 0 1 1104
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220673
transform 1 0 104 0 1 1104
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220673
transform 1 0 1280 0 -1 1088
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220673
transform 1 0 104 0 -1 1088
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220673
transform 1 0 1280 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220673
transform 1 0 104 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220673
transform 1 0 1280 0 -1 976
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220673
transform 1 0 104 0 -1 976
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220673
transform 1 0 1280 0 1 872
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220673
transform 1 0 104 0 1 872
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220673
transform 1 0 1280 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220673
transform 1 0 104 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220673
transform 1 0 1280 0 1 760
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220673
transform 1 0 104 0 1 760
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220673
transform 1 0 1280 0 -1 752
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220673
transform 1 0 104 0 -1 752
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220673
transform 1 0 1280 0 1 656
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220673
transform 1 0 104 0 1 656
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220673
transform 1 0 1280 0 -1 644
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220673
transform 1 0 104 0 -1 644
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220673
transform 1 0 1280 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220673
transform 1 0 104 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220673
transform 1 0 1280 0 -1 532
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220673
transform 1 0 104 0 -1 532
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220673
transform 1 0 1280 0 1 432
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220673
transform 1 0 104 0 1 432
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220673
transform 1 0 1280 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220673
transform 1 0 104 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220673
transform 1 0 1280 0 1 324
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220673
transform 1 0 104 0 1 324
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220673
transform 1 0 1280 0 -1 312
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220673
transform 1 0 104 0 -1 312
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220673
transform 1 0 1280 0 1 216
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220673
transform 1 0 104 0 1 216
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220673
transform 1 0 1280 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220673
transform 1 0 104 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220673
transform 1 0 1280 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220673
transform 1 0 104 0 1 100
box 7 3 12 24
use _0_0std_0_0cells_0_0OR2X1  tst_5999_6
timestamp 1731220673
transform 1 0 2368 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5998_6
timestamp 1731220673
transform 1 0 2432 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5997_6
timestamp 1731220673
transform 1 0 2432 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5996_6
timestamp 1731220673
transform 1 0 2432 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5995_6
timestamp 1731220673
transform 1 0 2352 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5994_6
timestamp 1731220673
transform 1 0 2256 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5993_6
timestamp 1731220673
transform 1 0 2352 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5992_6
timestamp 1731220673
transform 1 0 2352 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5991_6
timestamp 1731220673
transform 1 0 2360 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5990_6
timestamp 1731220673
transform 1 0 2360 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5989_6
timestamp 1731220673
transform 1 0 2272 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5988_6
timestamp 1731220673
transform 1 0 2248 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5987_6
timestamp 1731220673
transform 1 0 2144 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5986_6
timestamp 1731220673
transform 1 0 2048 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5985_6
timestamp 1731220673
transform 1 0 2184 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5984_6
timestamp 1731220673
transform 1 0 2320 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5983_6
timestamp 1731220673
transform 1 0 2312 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5982_6
timestamp 1731220673
transform 1 0 2176 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5981_6
timestamp 1731220673
transform 1 0 2048 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5980_6
timestamp 1731220673
transform 1 0 2024 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5979_6
timestamp 1731220673
transform 1 0 1920 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5978_6
timestamp 1731220673
transform 1 0 1816 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5977_6
timestamp 1731220673
transform 1 0 1816 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5976_6
timestamp 1731220673
transform 1 0 1928 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5975_6
timestamp 1731220673
transform 1 0 2056 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5974_6
timestamp 1731220673
transform 1 0 1936 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5973_6
timestamp 1731220673
transform 1 0 1824 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5972_6
timestamp 1731220673
transform 1 0 1848 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5971_6
timestamp 1731220673
transform 1 0 1952 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5970_6
timestamp 1731220673
transform 1 0 1896 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5969_6
timestamp 1731220673
transform 1 0 1920 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5968_6
timestamp 1731220673
transform 1 0 1832 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5967_6
timestamp 1731220673
transform 1 0 1944 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5966_6
timestamp 1731220673
transform 1 0 1944 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5965_6
timestamp 1731220673
transform 1 0 1840 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5964_6
timestamp 1731220673
transform 1 0 1800 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5963_6
timestamp 1731220673
transform 1 0 1888 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5962_6
timestamp 1731220673
transform 1 0 1984 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5961_6
timestamp 1731220673
transform 1 0 1920 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5960_6
timestamp 1731220673
transform 1 0 1856 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5959_6
timestamp 1731220673
transform 1 0 1800 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5958_6
timestamp 1731220673
transform 1 0 1984 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5957_6
timestamp 1731220673
transform 1 0 2048 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5956_6
timestamp 1731220673
transform 1 0 2280 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5955_6
timestamp 1731220673
transform 1 0 2200 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5954_6
timestamp 1731220673
transform 1 0 2120 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5953_6
timestamp 1731220673
transform 1 0 2096 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5952_6
timestamp 1731220673
transform 1 0 2208 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5951_6
timestamp 1731220673
transform 1 0 2328 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5950_6
timestamp 1731220673
transform 1 0 2248 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5949_6
timestamp 1731220673
transform 1 0 2152 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5948_6
timestamp 1731220673
transform 1 0 2048 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5947_6
timestamp 1731220673
transform 1 0 2056 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5946_6
timestamp 1731220673
transform 1 0 2160 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5945_6
timestamp 1731220673
transform 1 0 2176 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5944_6
timestamp 1731220673
transform 1 0 2264 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5943_6
timestamp 1731220673
transform 1 0 2264 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5942_6
timestamp 1731220673
transform 1 0 2168 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5941_6
timestamp 1731220673
transform 1 0 2096 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5940_6
timestamp 1731220673
transform 1 0 2000 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5939_6
timestamp 1731220673
transform 1 0 2184 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5938_6
timestamp 1731220673
transform 1 0 2352 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5937_6
timestamp 1731220673
transform 1 0 2432 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5936_6
timestamp 1731220673
transform 1 0 2432 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5935_6
timestamp 1731220673
transform 1 0 2432 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5934_6
timestamp 1731220673
transform 1 0 2432 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5933_6
timestamp 1731220673
transform 1 0 2432 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5932_6
timestamp 1731220673
transform 1 0 2432 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5931_6
timestamp 1731220673
transform 1 0 2432 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5930_6
timestamp 1731220673
transform 1 0 2432 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5929_6
timestamp 1731220673
transform 1 0 2432 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5928_6
timestamp 1731220673
transform 1 0 2432 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5927_6
timestamp 1731220673
transform 1 0 2432 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5926_6
timestamp 1731220673
transform 1 0 2432 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5925_6
timestamp 1731220673
transform 1 0 2432 0 1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5924_6
timestamp 1731220673
transform 1 0 2432 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5923_6
timestamp 1731220673
transform 1 0 2432 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5922_6
timestamp 1731220673
transform 1 0 2432 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5921_6
timestamp 1731220673
transform 1 0 2376 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5920_6
timestamp 1731220673
transform 1 0 2376 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5919_6
timestamp 1731220673
transform 1 0 2360 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5918_6
timestamp 1731220673
transform 1 0 2432 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5917_6
timestamp 1731220673
transform 1 0 2416 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5916_6
timestamp 1731220673
transform 1 0 2360 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5915_6
timestamp 1731220673
transform 1 0 2264 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5914_6
timestamp 1731220673
transform 1 0 2168 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5913_6
timestamp 1731220673
transform 1 0 2336 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5912_6
timestamp 1731220673
transform 1 0 2344 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5911_6
timestamp 1731220673
transform 1 0 2232 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5910_6
timestamp 1731220673
transform 1 0 2128 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5909_6
timestamp 1731220673
transform 1 0 2224 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5908_6
timestamp 1731220673
transform 1 0 2112 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5907_6
timestamp 1731220673
transform 1 0 2008 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5906_6
timestamp 1731220673
transform 1 0 1912 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5905_6
timestamp 1731220673
transform 1 0 2080 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5904_6
timestamp 1731220673
transform 1 0 1992 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5903_6
timestamp 1731220673
transform 1 0 1904 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5902_6
timestamp 1731220673
transform 1 0 1888 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5901_6
timestamp 1731220673
transform 1 0 1784 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5900_6
timestamp 1731220673
transform 1 0 2008 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5899_6
timestamp 1731220673
transform 1 0 2272 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5898_6
timestamp 1731220673
transform 1 0 2136 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5897_6
timestamp 1731220673
transform 1 0 2104 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5896_6
timestamp 1731220673
transform 1 0 2008 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5895_6
timestamp 1731220673
transform 1 0 1912 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5894_6
timestamp 1731220673
transform 1 0 2192 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5893_6
timestamp 1731220673
transform 1 0 2272 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5892_6
timestamp 1731220673
transform 1 0 2352 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5891_6
timestamp 1731220673
transform 1 0 2360 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5890_6
timestamp 1731220673
transform 1 0 2264 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5889_6
timestamp 1731220673
transform 1 0 2168 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5888_6
timestamp 1731220673
transform 1 0 2064 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5887_6
timestamp 1731220673
transform 1 0 1944 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5886_6
timestamp 1731220673
transform 1 0 1816 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5885_6
timestamp 1731220673
transform 1 0 2344 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5884_6
timestamp 1731220673
transform 1 0 2232 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5883_6
timestamp 1731220673
transform 1 0 2128 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5882_6
timestamp 1731220673
transform 1 0 2016 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5881_6
timestamp 1731220673
transform 1 0 1904 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5880_6
timestamp 1731220673
transform 1 0 2208 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5879_6
timestamp 1731220673
transform 1 0 2128 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5878_6
timestamp 1731220673
transform 1 0 2048 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5877_6
timestamp 1731220673
transform 1 0 1976 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5876_6
timestamp 1731220673
transform 1 0 1904 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5875_6
timestamp 1731220673
transform 1 0 1824 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5874_6
timestamp 1731220673
transform 1 0 1880 0 1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5873_6
timestamp 1731220673
transform 1 0 2008 0 1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5872_6
timestamp 1731220673
transform 1 0 2152 0 1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5871_6
timestamp 1731220673
transform 1 0 2304 0 1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5870_6
timestamp 1731220673
transform 1 0 2264 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5869_6
timestamp 1731220673
transform 1 0 2176 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5868_6
timestamp 1731220673
transform 1 0 2096 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5867_6
timestamp 1731220673
transform 1 0 2072 0 1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5866_6
timestamp 1731220673
transform 1 0 2184 0 1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5865_6
timestamp 1731220673
transform 1 0 2296 0 1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5864_6
timestamp 1731220673
transform 1 0 2216 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5863_6
timestamp 1731220673
transform 1 0 2136 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5862_6
timestamp 1731220673
transform 1 0 2056 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5861_6
timestamp 1731220673
transform 1 0 2296 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5860_6
timestamp 1731220673
transform 1 0 2296 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5859_6
timestamp 1731220673
transform 1 0 2224 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5858_6
timestamp 1731220673
transform 1 0 2152 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5857_6
timestamp 1731220673
transform 1 0 2072 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5856_6
timestamp 1731220673
transform 1 0 1984 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5855_6
timestamp 1731220673
transform 1 0 2240 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5854_6
timestamp 1731220673
transform 1 0 2152 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5853_6
timestamp 1731220673
transform 1 0 2064 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5852_6
timestamp 1731220673
transform 1 0 1984 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5851_6
timestamp 1731220673
transform 1 0 1896 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5850_6
timestamp 1731220673
transform 1 0 1808 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5849_6
timestamp 1731220673
transform 1 0 2096 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5848_6
timestamp 1731220673
transform 1 0 2008 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5847_6
timestamp 1731220673
transform 1 0 1928 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5846_6
timestamp 1731220673
transform 1 0 1848 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5845_6
timestamp 1731220673
transform 1 0 1768 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5844_6
timestamp 1731220673
transform 1 0 2000 0 -1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5843_6
timestamp 1731220673
transform 1 0 1864 0 -1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5842_6
timestamp 1731220673
transform 1 0 1728 0 -1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5841_6
timestamp 1731220673
transform 1 0 1600 0 -1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5840_6
timestamp 1731220673
transform 1 0 1464 0 -1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5839_6
timestamp 1731220673
transform 1 0 1696 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5838_6
timestamp 1731220673
transform 1 0 1768 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5837_6
timestamp 1731220673
transform 1 0 1848 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5836_6
timestamp 1731220673
transform 1 0 2008 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5835_6
timestamp 1731220673
transform 1 0 1928 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5834_6
timestamp 1731220673
transform 1 0 1888 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5833_6
timestamp 1731220673
transform 1 0 1776 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5832_6
timestamp 1731220673
transform 1 0 2296 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5831_6
timestamp 1731220673
transform 1 0 2152 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5830_6
timestamp 1731220673
transform 1 0 2016 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5829_6
timestamp 1731220673
transform 1 0 1992 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5828_6
timestamp 1731220673
transform 1 0 1896 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5827_6
timestamp 1731220673
transform 1 0 2176 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5826_6
timestamp 1731220673
transform 1 0 2088 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5825_6
timestamp 1731220673
transform 1 0 2048 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5824_6
timestamp 1731220673
transform 1 0 1960 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5823_6
timestamp 1731220673
transform 1 0 2128 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5822_6
timestamp 1731220673
transform 1 0 2208 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5821_6
timestamp 1731220673
transform 1 0 2168 0 1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5820_6
timestamp 1731220673
transform 1 0 2312 0 1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5819_6
timestamp 1731220673
transform 1 0 2288 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5818_6
timestamp 1731220673
transform 1 0 2368 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5817_6
timestamp 1731220673
transform 1 0 2360 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5816_6
timestamp 1731220673
transform 1 0 2264 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5815_6
timestamp 1731220673
transform 1 0 2432 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5814_6
timestamp 1731220673
transform 1 0 2432 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5813_6
timestamp 1731220673
transform 1 0 2432 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5812_6
timestamp 1731220673
transform 1 0 2432 0 1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5811_6
timestamp 1731220673
transform 1 0 2432 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5810_6
timestamp 1731220673
transform 1 0 2432 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5809_6
timestamp 1731220673
transform 1 0 2352 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5808_6
timestamp 1731220673
transform 1 0 2376 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5807_6
timestamp 1731220673
transform 1 0 2320 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5806_6
timestamp 1731220673
transform 1 0 2256 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5805_6
timestamp 1731220673
transform 1 0 2192 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5804_6
timestamp 1731220673
transform 1 0 2128 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5803_6
timestamp 1731220673
transform 1 0 2064 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5802_6
timestamp 1731220673
transform 1 0 2000 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5801_6
timestamp 1731220673
transform 1 0 2256 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5800_6
timestamp 1731220673
transform 1 0 2160 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5799_6
timestamp 1731220673
transform 1 0 2064 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5798_6
timestamp 1731220673
transform 1 0 1976 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5797_6
timestamp 1731220673
transform 1 0 1896 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5796_6
timestamp 1731220673
transform 1 0 2024 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5795_6
timestamp 1731220673
transform 1 0 1952 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5794_6
timestamp 1731220673
transform 1 0 1888 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5793_6
timestamp 1731220673
transform 1 0 1824 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5792_6
timestamp 1731220673
transform 1 0 1760 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5791_6
timestamp 1731220673
transform 1 0 1728 0 1 2000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5790_6
timestamp 1731220673
transform 1 0 1816 0 1 2000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5789_6
timestamp 1731220673
transform 1 0 2096 0 1 2000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5788_6
timestamp 1731220673
transform 1 0 2000 0 1 2000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5787_6
timestamp 1731220673
transform 1 0 1904 0 1 2000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5786_6
timestamp 1731220673
transform 1 0 1848 0 -1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5785_6
timestamp 1731220673
transform 1 0 1984 0 -1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5784_6
timestamp 1731220673
transform 1 0 2360 0 -1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5783_6
timestamp 1731220673
transform 1 0 2232 0 -1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5782_6
timestamp 1731220673
transform 1 0 2112 0 -1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5781_6
timestamp 1731220673
transform 1 0 1968 0 1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5780_6
timestamp 1731220673
transform 1 0 1792 0 1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5779_6
timestamp 1731220673
transform 1 0 2136 0 1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5778_6
timestamp 1731220673
transform 1 0 2296 0 1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5777_6
timestamp 1731220673
transform 1 0 2432 0 1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5776_6
timestamp 1731220673
transform 1 0 2432 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5775_6
timestamp 1731220673
transform 1 0 2376 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5774_6
timestamp 1731220673
transform 1 0 2312 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5773_6
timestamp 1731220673
transform 1 0 2248 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5772_6
timestamp 1731220673
transform 1 0 2184 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5771_6
timestamp 1731220673
transform 1 0 2120 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5770_6
timestamp 1731220673
transform 1 0 2048 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5769_6
timestamp 1731220673
transform 1 0 1976 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5768_6
timestamp 1731220673
transform 1 0 1896 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5767_6
timestamp 1731220673
transform 1 0 1808 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5766_6
timestamp 1731220673
transform 1 0 1712 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5765_6
timestamp 1731220673
transform 1 0 2216 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5764_6
timestamp 1731220673
transform 1 0 2104 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5763_6
timestamp 1731220673
transform 1 0 1992 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5762_6
timestamp 1731220673
transform 1 0 1880 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5761_6
timestamp 1731220673
transform 1 0 2136 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5760_6
timestamp 1731220673
transform 1 0 2056 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5759_6
timestamp 1731220673
transform 1 0 1976 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5758_6
timestamp 1731220673
transform 1 0 1896 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5757_6
timestamp 1731220673
transform 1 0 1824 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5756_6
timestamp 1731220673
transform 1 0 1832 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5755_6
timestamp 1731220673
transform 1 0 1896 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5754_6
timestamp 1731220673
transform 1 0 2088 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5753_6
timestamp 1731220673
transform 1 0 2024 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5752_6
timestamp 1731220673
transform 1 0 1960 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5751_6
timestamp 1731220673
transform 1 0 1944 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5750_6
timestamp 1731220673
transform 1 0 1872 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5749_6
timestamp 1731220673
transform 1 0 2016 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5748_6
timestamp 1731220673
transform 1 0 2088 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5747_6
timestamp 1731220673
transform 1 0 2160 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5746_6
timestamp 1731220673
transform 1 0 2160 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5745_6
timestamp 1731220673
transform 1 0 2088 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5744_6
timestamp 1731220673
transform 1 0 2016 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5743_6
timestamp 1731220673
transform 1 0 1944 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5742_6
timestamp 1731220673
transform 1 0 1872 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5741_6
timestamp 1731220673
transform 1 0 2160 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5740_6
timestamp 1731220673
transform 1 0 2104 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5739_6
timestamp 1731220673
transform 1 0 2048 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5738_6
timestamp 1731220673
transform 1 0 1992 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5737_6
timestamp 1731220673
transform 1 0 1936 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5736_6
timestamp 1731220673
transform 1 0 1880 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5735_6
timestamp 1731220673
transform 1 0 1824 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5734_6
timestamp 1731220673
transform 1 0 1768 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5733_6
timestamp 1731220673
transform 1 0 1712 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5732_6
timestamp 1731220673
transform 1 0 1656 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5731_6
timestamp 1731220673
transform 1 0 1600 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5730_6
timestamp 1731220673
transform 1 0 1544 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5729_6
timestamp 1731220673
transform 1 0 1488 0 -1 2560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5728_6
timestamp 1731220673
transform 1 0 1800 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5727_6
timestamp 1731220673
transform 1 0 1728 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5726_6
timestamp 1731220673
transform 1 0 1656 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5725_6
timestamp 1731220673
transform 1 0 1584 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5724_6
timestamp 1731220673
transform 1 0 1520 0 1 2456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5723_6
timestamp 1731220673
transform 1 0 1536 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5722_6
timestamp 1731220673
transform 1 0 1600 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5721_6
timestamp 1731220673
transform 1 0 1664 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5720_6
timestamp 1731220673
transform 1 0 1736 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5719_6
timestamp 1731220673
transform 1 0 1808 0 -1 2452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5718_6
timestamp 1731220673
transform 1 0 1768 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5717_6
timestamp 1731220673
transform 1 0 1712 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5716_6
timestamp 1731220673
transform 1 0 1656 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5715_6
timestamp 1731220673
transform 1 0 1600 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5714_6
timestamp 1731220673
transform 1 0 1544 0 1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5713_6
timestamp 1731220673
transform 1 0 1752 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5712_6
timestamp 1731220673
transform 1 0 1680 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5711_6
timestamp 1731220673
transform 1 0 1600 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5710_6
timestamp 1731220673
transform 1 0 1528 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5709_6
timestamp 1731220673
transform 1 0 1464 0 -1 2336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5708_6
timestamp 1731220673
transform 1 0 1768 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5707_6
timestamp 1731220673
transform 1 0 1664 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5706_6
timestamp 1731220673
transform 1 0 1560 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5705_6
timestamp 1731220673
transform 1 0 1456 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5704_6
timestamp 1731220673
transform 1 0 1360 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5703_6
timestamp 1731220673
transform 1 0 1360 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5702_6
timestamp 1731220673
transform 1 0 1600 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5701_6
timestamp 1731220673
transform 1 0 1480 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5700_6
timestamp 1731220673
transform 1 0 1384 0 1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5699_6
timestamp 1731220673
transform 1 0 1600 0 1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5698_6
timestamp 1731220673
transform 1 0 1704 0 -1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5697_6
timestamp 1731220673
transform 1 0 1544 0 -1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5696_6
timestamp 1731220673
transform 1 0 1376 0 -1 2108
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5695_6
timestamp 1731220673
transform 1 0 1424 0 1 2000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5694_6
timestamp 1731220673
transform 1 0 1632 0 1 2000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5693_6
timestamp 1731220673
transform 1 0 1528 0 1 2000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5692_6
timestamp 1731220673
transform 1 0 1504 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5691_6
timestamp 1731220673
transform 1 0 1448 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5690_6
timestamp 1731220673
transform 1 0 1568 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5689_6
timestamp 1731220673
transform 1 0 1632 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5688_6
timestamp 1731220673
transform 1 0 1696 0 -1 1996
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5687_6
timestamp 1731220673
transform 1 0 1680 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5686_6
timestamp 1731220673
transform 1 0 1608 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5685_6
timestamp 1731220673
transform 1 0 1544 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5684_6
timestamp 1731220673
transform 1 0 1824 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5683_6
timestamp 1731220673
transform 1 0 1752 0 1 1888
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5682_6
timestamp 1731220673
transform 1 0 1720 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5681_6
timestamp 1731220673
transform 1 0 1656 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5680_6
timestamp 1731220673
transform 1 0 1600 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5679_6
timestamp 1731220673
transform 1 0 1792 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5678_6
timestamp 1731220673
transform 1 0 1864 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5677_6
timestamp 1731220673
transform 1 0 1936 0 -1 1884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5676_6
timestamp 1731220673
transform 1 0 2032 0 1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5675_6
timestamp 1731220673
transform 1 0 1904 0 1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5674_6
timestamp 1731220673
transform 1 0 1792 0 1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5673_6
timestamp 1731220673
transform 1 0 1696 0 1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5672_6
timestamp 1731220673
transform 1 0 1608 0 1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5671_6
timestamp 1731220673
transform 1 0 1872 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5670_6
timestamp 1731220673
transform 1 0 1784 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5669_6
timestamp 1731220673
transform 1 0 1688 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5668_6
timestamp 1731220673
transform 1 0 1600 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5667_6
timestamp 1731220673
transform 1 0 1520 0 -1 1776
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5666_6
timestamp 1731220673
transform 1 0 1800 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5665_6
timestamp 1731220673
transform 1 0 1704 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5664_6
timestamp 1731220673
transform 1 0 1608 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5663_6
timestamp 1731220673
transform 1 0 1520 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5662_6
timestamp 1731220673
transform 1 0 1440 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5661_6
timestamp 1731220673
transform 1 0 1376 0 1 1668
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5660_6
timestamp 1731220673
transform 1 0 1672 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5659_6
timestamp 1731220673
transform 1 0 1576 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5658_6
timestamp 1731220673
transform 1 0 1488 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5657_6
timestamp 1731220673
transform 1 0 1400 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5656_6
timestamp 1731220673
transform 1 0 1344 0 -1 1664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5655_6
timestamp 1731220673
transform 1 0 1616 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5654_6
timestamp 1731220673
transform 1 0 1536 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5653_6
timestamp 1731220673
transform 1 0 1456 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5652_6
timestamp 1731220673
transform 1 0 1400 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5651_6
timestamp 1731220673
transform 1 0 1344 0 1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5650_6
timestamp 1731220673
transform 1 0 1216 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5649_6
timestamp 1731220673
transform 1 0 1160 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5648_6
timestamp 1731220673
transform 1 0 1080 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5647_6
timestamp 1731220673
transform 1 0 1344 0 -1 1560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5646_6
timestamp 1731220673
transform 1 0 1344 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5645_6
timestamp 1731220673
transform 1 0 1400 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5644_6
timestamp 1731220673
transform 1 0 1456 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5643_6
timestamp 1731220673
transform 1 0 1688 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5642_6
timestamp 1731220673
transform 1 0 1608 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5641_6
timestamp 1731220673
transform 1 0 1528 0 1 1456
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5640_6
timestamp 1731220673
transform 1 0 1528 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5639_6
timestamp 1731220673
transform 1 0 1440 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5638_6
timestamp 1731220673
transform 1 0 1352 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5637_6
timestamp 1731220673
transform 1 0 1624 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5636_6
timestamp 1731220673
transform 1 0 1720 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5635_6
timestamp 1731220673
transform 1 0 1712 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5634_6
timestamp 1731220673
transform 1 0 1624 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5633_6
timestamp 1731220673
transform 1 0 1544 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5632_6
timestamp 1731220673
transform 1 0 1808 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5631_6
timestamp 1731220673
transform 1 0 1896 0 1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5630_6
timestamp 1731220673
transform 1 0 1888 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5629_6
timestamp 1731220673
transform 1 0 1800 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5628_6
timestamp 1731220673
transform 1 0 1976 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5627_6
timestamp 1731220673
transform 1 0 1968 0 1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5626_6
timestamp 1731220673
transform 1 0 2024 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5625_6
timestamp 1731220673
transform 1 0 1960 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5624_6
timestamp 1731220673
transform 1 0 1904 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5623_6
timestamp 1731220673
transform 1 0 1848 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5622_6
timestamp 1731220673
transform 1 0 1792 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5621_6
timestamp 1731220673
transform 1 0 1736 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5620_6
timestamp 1731220673
transform 1 0 1680 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5619_6
timestamp 1731220673
transform 1 0 1624 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5618_6
timestamp 1731220673
transform 1 0 1688 0 1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5617_6
timestamp 1731220673
transform 1 0 1872 0 1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5616_6
timestamp 1731220673
transform 1 0 1776 0 1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5615_6
timestamp 1731220673
transform 1 0 1720 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5614_6
timestamp 1731220673
transform 1 0 1640 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5613_6
timestamp 1731220673
transform 1 0 1576 0 -1 1344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5612_6
timestamp 1731220673
transform 1 0 1544 0 1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5611_6
timestamp 1731220673
transform 1 0 1608 0 1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5610_6
timestamp 1731220673
transform 1 0 1568 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5609_6
timestamp 1731220673
transform 1 0 1512 0 -1 1236
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5608_6
timestamp 1731220673
transform 1 0 1768 0 1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5607_6
timestamp 1731220673
transform 1 0 1680 0 1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5606_6
timestamp 1731220673
transform 1 0 1608 0 1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5605_6
timestamp 1731220673
transform 1 0 1544 0 1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5604_6
timestamp 1731220673
transform 1 0 1744 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5603_6
timestamp 1731220673
transform 1 0 1664 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5602_6
timestamp 1731220673
transform 1 0 1584 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5601_6
timestamp 1731220673
transform 1 0 1512 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5600_6
timestamp 1731220673
transform 1 0 1440 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5599_6
timestamp 1731220673
transform 1 0 1376 0 -1 1128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5598_6
timestamp 1731220673
transform 1 0 1792 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5597_6
timestamp 1731220673
transform 1 0 1672 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5596_6
timestamp 1731220673
transform 1 0 1552 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5595_6
timestamp 1731220673
transform 1 0 1432 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5594_6
timestamp 1731220673
transform 1 0 1344 0 1 1016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5593_6
timestamp 1731220673
transform 1 0 1672 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5592_6
timestamp 1731220673
transform 1 0 1504 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5591_6
timestamp 1731220673
transform 1 0 1216 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5590_6
timestamp 1731220673
transform 1 0 1160 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5589_6
timestamp 1731220673
transform 1 0 1080 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5588_6
timestamp 1731220673
transform 1 0 1000 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5587_6
timestamp 1731220673
transform 1 0 920 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5586_6
timestamp 1731220673
transform 1 0 832 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5585_6
timestamp 1731220673
transform 1 0 744 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5584_6
timestamp 1731220673
transform 1 0 1080 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5583_6
timestamp 1731220673
transform 1 0 1160 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5582_6
timestamp 1731220673
transform 1 0 1160 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5581_6
timestamp 1731220673
transform 1 0 1064 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5580_6
timestamp 1731220673
transform 1 0 968 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5579_6
timestamp 1731220673
transform 1 0 880 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5578_6
timestamp 1731220673
transform 1 0 784 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5577_6
timestamp 1731220673
transform 1 0 896 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5576_6
timestamp 1731220673
transform 1 0 824 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5575_6
timestamp 1731220673
transform 1 0 752 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5574_6
timestamp 1731220673
transform 1 0 688 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5573_6
timestamp 1731220673
transform 1 0 624 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5572_6
timestamp 1731220673
transform 1 0 680 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5571_6
timestamp 1731220673
transform 1 0 608 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5570_6
timestamp 1731220673
transform 1 0 536 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5569_6
timestamp 1731220673
transform 1 0 456 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5568_6
timestamp 1731220673
transform 1 0 368 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5567_6
timestamp 1731220673
transform 1 0 560 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5566_6
timestamp 1731220673
transform 1 0 496 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5565_6
timestamp 1731220673
transform 1 0 432 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5564_6
timestamp 1731220673
transform 1 0 368 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5563_6
timestamp 1731220673
transform 1 0 688 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5562_6
timestamp 1731220673
transform 1 0 592 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5561_6
timestamp 1731220673
transform 1 0 496 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5560_6
timestamp 1731220673
transform 1 0 400 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5559_6
timestamp 1731220673
transform 1 0 448 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5558_6
timestamp 1731220673
transform 1 0 352 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5557_6
timestamp 1731220673
transform 1 0 264 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5556_6
timestamp 1731220673
transform 1 0 272 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5555_6
timestamp 1731220673
transform 1 0 360 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5554_6
timestamp 1731220673
transform 1 0 456 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5553_6
timestamp 1731220673
transform 1 0 440 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5552_6
timestamp 1731220673
transform 1 0 352 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5551_6
timestamp 1731220673
transform 1 0 272 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5550_6
timestamp 1731220673
transform 1 0 200 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5549_6
timestamp 1731220673
transform 1 0 160 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5548_6
timestamp 1731220673
transform 1 0 256 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5547_6
timestamp 1731220673
transform 1 0 352 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5546_6
timestamp 1731220673
transform 1 0 344 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5545_6
timestamp 1731220673
transform 1 0 264 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5544_6
timestamp 1731220673
transform 1 0 184 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5543_6
timestamp 1731220673
transform 1 0 128 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5542_6
timestamp 1731220673
transform 1 0 368 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5541_6
timestamp 1731220673
transform 1 0 280 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5540_6
timestamp 1731220673
transform 1 0 192 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5539_6
timestamp 1731220673
transform 1 0 128 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5538_6
timestamp 1731220673
transform 1 0 128 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5537_6
timestamp 1731220673
transform 1 0 360 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5536_6
timestamp 1731220673
transform 1 0 232 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5535_6
timestamp 1731220673
transform 1 0 200 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5534_6
timestamp 1731220673
transform 1 0 128 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5533_6
timestamp 1731220673
transform 1 0 184 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5532_6
timestamp 1731220673
transform 1 0 248 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5531_6
timestamp 1731220673
transform 1 0 256 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5530_6
timestamp 1731220673
transform 1 0 240 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5529_6
timestamp 1731220673
transform 1 0 488 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5528_6
timestamp 1731220673
transform 1 0 576 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5527_6
timestamp 1731220673
transform 1 0 568 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5526_6
timestamp 1731220673
transform 1 0 584 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5525_6
timestamp 1731220673
transform 1 0 496 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5524_6
timestamp 1731220673
transform 1 0 600 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5523_6
timestamp 1731220673
transform 1 0 568 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5522_6
timestamp 1731220673
transform 1 0 536 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5521_6
timestamp 1731220673
transform 1 0 624 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5520_6
timestamp 1731220673
transform 1 0 720 0 1 1908
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5519_6
timestamp 1731220673
transform 1 0 896 0 1 1908
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5518_6
timestamp 1731220673
transform 1 0 840 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5517_6
timestamp 1731220673
transform 1 0 728 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5516_6
timestamp 1731220673
transform 1 0 688 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5515_6
timestamp 1731220673
transform 1 0 768 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5514_6
timestamp 1731220673
transform 1 0 920 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5513_6
timestamp 1731220673
transform 1 0 840 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5512_6
timestamp 1731220673
transform 1 0 792 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5511_6
timestamp 1731220673
transform 1 0 704 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5510_6
timestamp 1731220673
transform 1 0 880 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5509_6
timestamp 1731220673
transform 1 0 968 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5508_6
timestamp 1731220673
transform 1 0 936 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5507_6
timestamp 1731220673
transform 1 0 840 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5506_6
timestamp 1731220673
transform 1 0 744 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5505_6
timestamp 1731220673
transform 1 0 640 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5504_6
timestamp 1731220673
transform 1 0 616 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5503_6
timestamp 1731220673
transform 1 0 720 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5502_6
timestamp 1731220673
transform 1 0 824 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5501_6
timestamp 1731220673
transform 1 0 928 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5500_6
timestamp 1731220673
transform 1 0 888 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5499_6
timestamp 1731220673
transform 1 0 784 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5498_6
timestamp 1731220673
transform 1 0 680 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5497_6
timestamp 1731220673
transform 1 0 672 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5496_6
timestamp 1731220673
transform 1 0 600 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5495_6
timestamp 1731220673
transform 1 0 736 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5494_6
timestamp 1731220673
transform 1 0 800 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5493_6
timestamp 1731220673
transform 1 0 856 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5492_6
timestamp 1731220673
transform 1 0 920 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5491_6
timestamp 1731220673
transform 1 0 984 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5490_6
timestamp 1731220673
transform 1 0 1048 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5489_6
timestamp 1731220673
transform 1 0 1104 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5488_6
timestamp 1731220673
transform 1 0 1160 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5487_6
timestamp 1731220673
transform 1 0 1216 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5486_6
timestamp 1731220673
transform 1 0 1216 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5485_6
timestamp 1731220673
transform 1 0 1104 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5484_6
timestamp 1731220673
transform 1 0 992 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5483_6
timestamp 1731220673
transform 1 0 1032 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5482_6
timestamp 1731220673
transform 1 0 1216 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5481_6
timestamp 1731220673
transform 1 0 1136 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5480_6
timestamp 1731220673
transform 1 0 1032 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5479_6
timestamp 1731220673
transform 1 0 1136 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5478_6
timestamp 1731220673
transform 1 0 1216 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5477_6
timestamp 1731220673
transform 1 0 1216 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5476_6
timestamp 1731220673
transform 1 0 1144 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5475_6
timestamp 1731220673
transform 1 0 1056 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5474_6
timestamp 1731220673
transform 1 0 1216 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5473_6
timestamp 1731220673
transform 1 0 1160 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5472_6
timestamp 1731220673
transform 1 0 1080 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5471_6
timestamp 1731220673
transform 1 0 1000 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5470_6
timestamp 1731220673
transform 1 0 952 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5469_6
timestamp 1731220673
transform 1 0 1192 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5468_6
timestamp 1731220673
transform 1 0 1072 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5467_6
timestamp 1731220673
transform 1 0 1072 0 1 1908
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5466_6
timestamp 1731220673
transform 1 0 1008 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5465_6
timestamp 1731220673
transform 1 0 904 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5464_6
timestamp 1731220673
transform 1 0 880 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5463_6
timestamp 1731220673
transform 1 0 912 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5462_6
timestamp 1731220673
transform 1 0 856 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5461_6
timestamp 1731220673
transform 1 0 872 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5460_6
timestamp 1731220673
transform 1 0 752 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5459_6
timestamp 1731220673
transform 1 0 712 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5458_6
timestamp 1731220673
transform 1 0 792 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5457_6
timestamp 1731220673
transform 1 0 808 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5456_6
timestamp 1731220673
transform 1 0 816 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5455_6
timestamp 1731220673
transform 1 0 728 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5454_6
timestamp 1731220673
transform 1 0 576 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5453_6
timestamp 1731220673
transform 1 0 472 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5452_6
timestamp 1731220673
transform 1 0 528 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5451_6
timestamp 1731220673
transform 1 0 448 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5450_6
timestamp 1731220673
transform 1 0 424 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5449_6
timestamp 1731220673
transform 1 0 504 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5448_6
timestamp 1731220673
transform 1 0 448 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5447_6
timestamp 1731220673
transform 1 0 544 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5446_6
timestamp 1731220673
transform 1 0 536 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5445_6
timestamp 1731220673
transform 1 0 632 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5444_6
timestamp 1731220673
transform 1 0 552 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5443_6
timestamp 1731220673
transform 1 0 648 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5442_6
timestamp 1731220673
transform 1 0 648 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5441_6
timestamp 1731220673
transform 1 0 544 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5440_6
timestamp 1731220673
transform 1 0 320 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5439_6
timestamp 1731220673
transform 1 0 248 0 1 868
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5438_6
timestamp 1731220673
transform 1 0 240 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5437_6
timestamp 1731220673
transform 1 0 304 0 -1 864
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5436_6
timestamp 1731220673
transform 1 0 280 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5435_6
timestamp 1731220673
transform 1 0 192 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5434_6
timestamp 1731220673
transform 1 0 128 0 -1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5433_6
timestamp 1731220673
transform 1 0 248 0 -1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5432_6
timestamp 1731220673
transform 1 0 384 0 -1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5431_6
timestamp 1731220673
transform 1 0 480 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5430_6
timestamp 1731220673
transform 1 0 368 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5429_6
timestamp 1731220673
transform 1 0 272 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5428_6
timestamp 1731220673
transform 1 0 184 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5427_6
timestamp 1731220673
transform 1 0 128 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5426_6
timestamp 1731220673
transform 1 0 256 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5425_6
timestamp 1731220673
transform 1 0 144 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5424_6
timestamp 1731220673
transform 1 0 128 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5423_6
timestamp 1731220673
transform 1 0 216 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5422_6
timestamp 1731220673
transform 1 0 312 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5421_6
timestamp 1731220673
transform 1 0 232 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5420_6
timestamp 1731220673
transform 1 0 136 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5419_6
timestamp 1731220673
transform 1 0 128 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5418_6
timestamp 1731220673
transform 1 0 184 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5417_6
timestamp 1731220673
transform 1 0 272 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5416_6
timestamp 1731220673
transform 1 0 184 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5415_6
timestamp 1731220673
transform 1 0 128 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5414_6
timestamp 1731220673
transform 1 0 128 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5413_6
timestamp 1731220673
transform 1 0 208 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5412_6
timestamp 1731220673
transform 1 0 208 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5411_6
timestamp 1731220673
transform 1 0 128 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5410_6
timestamp 1731220673
transform 1 0 128 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5409_6
timestamp 1731220673
transform 1 0 200 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5408_6
timestamp 1731220673
transform 1 0 296 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5407_6
timestamp 1731220673
transform 1 0 272 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5406_6
timestamp 1731220673
transform 1 0 176 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5405_6
timestamp 1731220673
transform 1 0 184 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5404_6
timestamp 1731220673
transform 1 0 128 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5403_6
timestamp 1731220673
transform 1 0 240 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5402_6
timestamp 1731220673
transform 1 0 296 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5401_6
timestamp 1731220673
transform 1 0 352 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5400_6
timestamp 1731220673
transform 1 0 408 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5399_6
timestamp 1731220673
transform 1 0 576 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5398_6
timestamp 1731220673
transform 1 0 520 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5397_6
timestamp 1731220673
transform 1 0 464 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5396_6
timestamp 1731220673
transform 1 0 376 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5395_6
timestamp 1731220673
transform 1 0 480 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5394_6
timestamp 1731220673
transform 1 0 584 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5393_6
timestamp 1731220673
transform 1 0 624 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5392_6
timestamp 1731220673
transform 1 0 512 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5391_6
timestamp 1731220673
transform 1 0 400 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5390_6
timestamp 1731220673
transform 1 0 312 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5389_6
timestamp 1731220673
transform 1 0 416 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5388_6
timestamp 1731220673
transform 1 0 528 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5387_6
timestamp 1731220673
transform 1 0 520 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5386_6
timestamp 1731220673
transform 1 0 416 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5385_6
timestamp 1731220673
transform 1 0 312 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5384_6
timestamp 1731220673
transform 1 0 600 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5383_6
timestamp 1731220673
transform 1 0 488 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5382_6
timestamp 1731220673
transform 1 0 376 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5381_6
timestamp 1731220673
transform 1 0 352 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5380_6
timestamp 1731220673
transform 1 0 264 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5379_6
timestamp 1731220673
transform 1 0 536 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5378_6
timestamp 1731220673
transform 1 0 440 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5377_6
timestamp 1731220673
transform 1 0 424 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5376_6
timestamp 1731220673
transform 1 0 328 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5375_6
timestamp 1731220673
transform 1 0 520 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5374_6
timestamp 1731220673
transform 1 0 608 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5373_6
timestamp 1731220673
transform 1 0 512 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5372_6
timestamp 1731220673
transform 1 0 408 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5371_6
timestamp 1731220673
transform 1 0 360 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5370_6
timestamp 1731220673
transform 1 0 456 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5369_6
timestamp 1731220673
transform 1 0 552 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5368_6
timestamp 1731220673
transform 1 0 648 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5367_6
timestamp 1731220673
transform 1 0 600 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5366_6
timestamp 1731220673
transform 1 0 720 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5365_6
timestamp 1731220673
transform 1 0 640 0 -1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5364_6
timestamp 1731220673
transform 1 0 512 0 -1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5363_6
timestamp 1731220673
transform 1 0 768 0 -1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5362_6
timestamp 1731220673
transform 1 0 744 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5361_6
timestamp 1731220673
transform 1 0 808 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5360_6
timestamp 1731220673
transform 1 0 872 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5359_6
timestamp 1731220673
transform 1 0 944 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5358_6
timestamp 1731220673
transform 1 0 1016 0 1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5357_6
timestamp 1731220673
transform 1 0 1032 0 -1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5356_6
timestamp 1731220673
transform 1 0 896 0 -1 756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5355_6
timestamp 1731220673
transform 1 0 848 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5354_6
timestamp 1731220673
transform 1 0 976 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5353_6
timestamp 1731220673
transform 1 0 936 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5352_6
timestamp 1731220673
transform 1 0 840 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5351_6
timestamp 1731220673
transform 1 0 744 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5350_6
timestamp 1731220673
transform 1 0 800 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5349_6
timestamp 1731220673
transform 1 0 704 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5348_6
timestamp 1731220673
transform 1 0 704 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5347_6
timestamp 1731220673
transform 1 0 616 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5346_6
timestamp 1731220673
transform 1 0 632 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5345_6
timestamp 1731220673
transform 1 0 728 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5344_6
timestamp 1731220673
transform 1 0 712 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5343_6
timestamp 1731220673
transform 1 0 728 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5342_6
timestamp 1731220673
transform 1 0 624 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5341_6
timestamp 1731220673
transform 1 0 632 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5340_6
timestamp 1731220673
transform 1 0 736 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5339_6
timestamp 1731220673
transform 1 0 840 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5338_6
timestamp 1731220673
transform 1 0 848 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5337_6
timestamp 1731220673
transform 1 0 736 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5336_6
timestamp 1731220673
transform 1 0 688 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5335_6
timestamp 1731220673
transform 1 0 792 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5334_6
timestamp 1731220673
transform 1 0 744 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5333_6
timestamp 1731220673
transform 1 0 688 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5332_6
timestamp 1731220673
transform 1 0 632 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5331_6
timestamp 1731220673
transform 1 0 808 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5330_6
timestamp 1731220673
transform 1 0 872 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5329_6
timestamp 1731220673
transform 1 0 936 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5328_6
timestamp 1731220673
transform 1 0 1000 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5327_6
timestamp 1731220673
transform 1 0 1064 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5326_6
timestamp 1731220673
transform 1 0 1128 0 1 96
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5325_6
timestamp 1731220673
transform 1 0 1096 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5324_6
timestamp 1731220673
transform 1 0 992 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5323_6
timestamp 1731220673
transform 1 0 888 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5322_6
timestamp 1731220673
transform 1 0 960 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5321_6
timestamp 1731220673
transform 1 0 1080 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5320_6
timestamp 1731220673
transform 1 0 1200 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5319_6
timestamp 1731220673
transform 1 0 1136 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5318_6
timestamp 1731220673
transform 1 0 1032 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5317_6
timestamp 1731220673
transform 1 0 936 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5316_6
timestamp 1731220673
transform 1 0 912 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5315_6
timestamp 1731220673
transform 1 0 824 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5314_6
timestamp 1731220673
transform 1 0 992 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5313_6
timestamp 1731220673
transform 1 0 928 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5312_6
timestamp 1731220673
transform 1 0 824 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5311_6
timestamp 1731220673
transform 1 0 1032 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5310_6
timestamp 1731220673
transform 1 0 928 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5309_6
timestamp 1731220673
transform 1 0 824 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5308_6
timestamp 1731220673
transform 1 0 784 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5307_6
timestamp 1731220673
transform 1 0 864 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5306_6
timestamp 1731220673
transform 1 0 1024 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5305_6
timestamp 1731220673
transform 1 0 944 0 -1 536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5304_6
timestamp 1731220673
transform 1 0 888 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5303_6
timestamp 1731220673
transform 1 0 976 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5302_6
timestamp 1731220673
transform 1 0 1064 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5301_6
timestamp 1731220673
transform 1 0 1160 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5300_6
timestamp 1731220673
transform 1 0 1136 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5299_6
timestamp 1731220673
transform 1 0 1032 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5298_6
timestamp 1731220673
transform 1 0 1216 0 -1 648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5297_6
timestamp 1731220673
transform 1 0 1600 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5296_6
timestamp 1731220673
transform 1 0 1704 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5295_6
timestamp 1731220673
transform 1 0 1720 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5294_6
timestamp 1731220673
transform 1 0 1624 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5293_6
timestamp 1731220673
transform 1 0 1528 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5292_6
timestamp 1731220673
transform 1 0 1544 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5291_6
timestamp 1731220673
transform 1 0 1640 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5290_6
timestamp 1731220673
transform 1 0 1744 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5289_6
timestamp 1731220673
transform 1 0 1784 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5288_6
timestamp 1731220673
transform 1 0 1672 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5287_6
timestamp 1731220673
transform 1 0 1552 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5286_6
timestamp 1731220673
transform 1 0 1576 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5285_6
timestamp 1731220673
transform 1 0 1632 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5284_6
timestamp 1731220673
transform 1 0 1688 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5283_6
timestamp 1731220673
transform 1 0 1752 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5282_6
timestamp 1731220673
transform 1 0 1824 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5281_6
timestamp 1731220673
transform 1 0 2000 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5280_6
timestamp 1731220673
transform 1 0 2088 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5279_6
timestamp 1731220673
transform 1 0 2072 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5278_6
timestamp 1731220673
transform 1 0 1984 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5277_6
timestamp 1731220673
transform 1 0 1904 0 -1 440
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5276_6
timestamp 1731220673
transform 1 0 1848 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5275_6
timestamp 1731220673
transform 1 0 1776 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5274_6
timestamp 1731220673
transform 1 0 1712 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5273_6
timestamp 1731220673
transform 1 0 1656 0 1 332
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5272_6
timestamp 1731220673
transform 1 0 1576 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5271_6
timestamp 1731220673
transform 1 0 1448 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5270_6
timestamp 1731220673
transform 1 0 1704 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5269_6
timestamp 1731220673
transform 1 0 1736 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5268_6
timestamp 1731220673
transform 1 0 1632 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5267_6
timestamp 1731220673
transform 1 0 1528 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5266_6
timestamp 1731220673
transform 1 0 1544 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5265_6
timestamp 1731220673
transform 1 0 1632 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5264_6
timestamp 1731220673
transform 1 0 1712 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5263_6
timestamp 1731220673
transform 1 0 1736 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5262_6
timestamp 1731220673
transform 1 0 1680 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5261_6
timestamp 1731220673
transform 1 0 1624 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5260_6
timestamp 1731220673
transform 1 0 1568 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5259_6
timestamp 1731220673
transform 1 0 1512 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5258_6
timestamp 1731220673
transform 1 0 1456 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5257_6
timestamp 1731220673
transform 1 0 1400 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5256_6
timestamp 1731220673
transform 1 0 1344 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5255_6
timestamp 1731220673
transform 1 0 1344 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5254_6
timestamp 1731220673
transform 1 0 1400 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5253_6
timestamp 1731220673
transform 1 0 1464 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5252_6
timestamp 1731220673
transform 1 0 1424 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5251_6
timestamp 1731220673
transform 1 0 1344 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5250_6
timestamp 1731220673
transform 1 0 1344 0 -1 324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5249_6
timestamp 1731220673
transform 1 0 1216 0 -1 316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5248_6
timestamp 1731220673
transform 1 0 1216 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5247_6
timestamp 1731220673
transform 1 0 1152 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5246_6
timestamp 1731220673
transform 1 0 1072 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5245_6
timestamp 1731220673
transform 1 0 1032 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5244_6
timestamp 1731220673
transform 1 0 1216 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5243_6
timestamp 1731220673
transform 1 0 1136 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5242_6
timestamp 1731220673
transform 1 0 1136 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5241_6
timestamp 1731220673
transform 1 0 1216 0 1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5240_6
timestamp 1731220673
transform 1 0 1344 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5239_6
timestamp 1731220673
transform 1 0 1432 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5238_6
timestamp 1731220673
transform 1 0 1448 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5237_6
timestamp 1731220673
transform 1 0 1368 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5236_6
timestamp 1731220673
transform 1 0 1360 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5235_6
timestamp 1731220673
transform 1 0 1440 0 1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5234_6
timestamp 1731220673
transform 1 0 1504 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5233_6
timestamp 1731220673
transform 1 0 1408 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5232_6
timestamp 1731220673
transform 1 0 1344 0 -1 664
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5231_6
timestamp 1731220673
transform 1 0 1216 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5230_6
timestamp 1731220673
transform 1 0 1104 0 1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5229_6
timestamp 1731220673
transform 1 0 1344 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5228_6
timestamp 1731220673
transform 1 0 1408 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5227_6
timestamp 1731220673
transform 1 0 1504 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5226_6
timestamp 1731220673
transform 1 0 1608 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5225_6
timestamp 1731220673
transform 1 0 1712 0 1 676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5224_6
timestamp 1731220673
transform 1 0 1680 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5223_6
timestamp 1731220673
transform 1 0 1616 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5222_6
timestamp 1731220673
transform 1 0 1560 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5221_6
timestamp 1731220673
transform 1 0 1752 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5220_6
timestamp 1731220673
transform 1 0 1824 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5219_6
timestamp 1731220673
transform 1 0 1824 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5218_6
timestamp 1731220673
transform 1 0 1744 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5217_6
timestamp 1731220673
transform 1 0 1680 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5216_6
timestamp 1731220673
transform 1 0 1624 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5215_6
timestamp 1731220673
transform 1 0 1568 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5214_6
timestamp 1731220673
transform 1 0 1696 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5213_6
timestamp 1731220673
transform 1 0 1616 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5212_6
timestamp 1731220673
transform 1 0 1544 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5211_6
timestamp 1731220673
transform 1 0 1480 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5210_6
timestamp 1731220673
transform 1 0 1424 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5209_6
timestamp 1731220673
transform 1 0 1808 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5208_6
timestamp 1731220673
transform 1 0 1696 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5207_6
timestamp 1731220673
transform 1 0 1584 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5206_6
timestamp 1731220673
transform 1 0 1480 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5205_6
timestamp 1731220673
transform 1 0 1400 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5204_6
timestamp 1731220673
transform 1 0 1344 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5203_6
timestamp 1731220673
transform 1 0 1344 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5202_6
timestamp 1731220673
transform 1 0 1216 0 -1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5201_6
timestamp 1731220673
transform 1 0 1000 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5200_6
timestamp 1731220673
transform 1 0 920 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5199_6
timestamp 1731220673
transform 1 0 832 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5198_6
timestamp 1731220673
transform 1 0 744 0 1 980
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5197_6
timestamp 1731220673
transform 1 0 1136 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5196_6
timestamp 1731220673
transform 1 0 1048 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5195_6
timestamp 1731220673
transform 1 0 968 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5194_6
timestamp 1731220673
transform 1 0 888 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5193_6
timestamp 1731220673
transform 1 0 808 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5192_6
timestamp 1731220673
transform 1 0 720 0 -1 1092
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5191_6
timestamp 1731220673
transform 1 0 1016 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5190_6
timestamp 1731220673
transform 1 0 936 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5189_6
timestamp 1731220673
transform 1 0 856 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5188_6
timestamp 1731220673
transform 1 0 784 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5187_6
timestamp 1731220673
transform 1 0 712 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5186_6
timestamp 1731220673
transform 1 0 632 0 1 1100
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5185_6
timestamp 1731220673
transform 1 0 856 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5184_6
timestamp 1731220673
transform 1 0 784 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5183_6
timestamp 1731220673
transform 1 0 712 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5182_6
timestamp 1731220673
transform 1 0 640 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5181_6
timestamp 1731220673
transform 1 0 576 0 -1 1208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5180_6
timestamp 1731220673
transform 1 0 600 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5179_6
timestamp 1731220673
transform 1 0 672 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5178_6
timestamp 1731220673
transform 1 0 896 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5177_6
timestamp 1731220673
transform 1 0 816 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5176_6
timestamp 1731220673
transform 1 0 744 0 1 1212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5175_6
timestamp 1731220673
transform 1 0 680 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5174_6
timestamp 1731220673
transform 1 0 776 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5173_6
timestamp 1731220673
transform 1 0 872 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5172_6
timestamp 1731220673
transform 1 0 968 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5171_6
timestamp 1731220673
transform 1 0 904 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5170_6
timestamp 1731220673
transform 1 0 992 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5169_6
timestamp 1731220673
transform 1 0 1080 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5168_6
timestamp 1731220673
transform 1 0 1176 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5167_6
timestamp 1731220673
transform 1 0 1216 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5166_6
timestamp 1731220673
transform 1 0 1120 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5165_6
timestamp 1731220673
transform 1 0 1016 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5164_6
timestamp 1731220673
transform 1 0 912 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5163_6
timestamp 1731220673
transform 1 0 1120 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5162_6
timestamp 1731220673
transform 1 0 1032 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5161_6
timestamp 1731220673
transform 1 0 952 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5160_6
timestamp 1731220673
transform 1 0 872 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5159_6
timestamp 1731220673
transform 1 0 840 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5158_6
timestamp 1731220673
transform 1 0 920 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5157_6
timestamp 1731220673
transform 1 0 1000 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5156_6
timestamp 1731220673
transform 1 0 984 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5155_6
timestamp 1731220673
transform 1 0 1096 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5154_6
timestamp 1731220673
transform 1 0 1056 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5153_6
timestamp 1731220673
transform 1 0 952 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5152_6
timestamp 1731220673
transform 1 0 1160 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5151_6
timestamp 1731220673
transform 1 0 1136 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5150_6
timestamp 1731220673
transform 1 0 1024 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5149_6
timestamp 1731220673
transform 1 0 968 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5148_6
timestamp 1731220673
transform 1 0 1056 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5147_6
timestamp 1731220673
transform 1 0 1144 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5146_6
timestamp 1731220673
transform 1 0 1136 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5145_6
timestamp 1731220673
transform 1 0 1056 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5144_6
timestamp 1731220673
transform 1 0 976 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5143_6
timestamp 1731220673
transform 1 0 1152 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5142_6
timestamp 1731220673
transform 1 0 1080 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5141_6
timestamp 1731220673
transform 1 0 936 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5140_6
timestamp 1731220673
transform 1 0 864 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5139_6
timestamp 1731220673
transform 1 0 792 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5138_6
timestamp 1731220673
transform 1 0 712 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5137_6
timestamp 1731220673
transform 1 0 664 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5136_6
timestamp 1731220673
transform 1 0 752 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5135_6
timestamp 1731220673
transform 1 0 832 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5134_6
timestamp 1731220673
transform 1 0 792 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5133_6
timestamp 1731220673
transform 1 0 696 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5132_6
timestamp 1731220673
transform 1 0 688 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5131_6
timestamp 1731220673
transform 1 0 800 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5130_6
timestamp 1731220673
transform 1 0 760 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5129_6
timestamp 1731220673
transform 1 0 664 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5128_6
timestamp 1731220673
transform 1 0 768 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5127_6
timestamp 1731220673
transform 1 0 672 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5126_6
timestamp 1731220673
transform 1 0 664 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5125_6
timestamp 1731220673
transform 1 0 632 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5124_6
timestamp 1731220673
transform 1 0 552 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5123_6
timestamp 1731220673
transform 1 0 600 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5122_6
timestamp 1731220673
transform 1 0 704 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5121_6
timestamp 1731220673
transform 1 0 640 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5120_6
timestamp 1731220673
transform 1 0 560 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5119_6
timestamp 1731220673
transform 1 0 480 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5118_6
timestamp 1731220673
transform 1 0 408 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5117_6
timestamp 1731220673
transform 1 0 336 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5116_6
timestamp 1731220673
transform 1 0 272 0 1 1340
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5115_6
timestamp 1731220673
transform 1 0 320 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5114_6
timestamp 1731220673
transform 1 0 400 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5113_6
timestamp 1731220673
transform 1 0 496 0 -1 1448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5112_6
timestamp 1731220673
transform 1 0 472 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5111_6
timestamp 1731220673
transform 1 0 392 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5110_6
timestamp 1731220673
transform 1 0 320 0 1 1452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5109_6
timestamp 1731220673
transform 1 0 312 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5108_6
timestamp 1731220673
transform 1 0 392 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5107_6
timestamp 1731220673
transform 1 0 576 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5106_6
timestamp 1731220673
transform 1 0 480 0 -1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5105_6
timestamp 1731220673
transform 1 0 408 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5104_6
timestamp 1731220673
transform 1 0 336 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5103_6
timestamp 1731220673
transform 1 0 280 0 1 1564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5102_6
timestamp 1731220673
transform 1 0 480 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5101_6
timestamp 1731220673
transform 1 0 392 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5100_6
timestamp 1731220673
transform 1 0 312 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_599_6
timestamp 1731220673
transform 1 0 248 0 -1 1672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_598_6
timestamp 1731220673
transform 1 0 480 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_597_6
timestamp 1731220673
transform 1 0 384 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_596_6
timestamp 1731220673
transform 1 0 296 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_595_6
timestamp 1731220673
transform 1 0 216 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_594_6
timestamp 1731220673
transform 1 0 144 0 1 1676
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_593_6
timestamp 1731220673
transform 1 0 392 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_592_6
timestamp 1731220673
transform 1 0 288 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_591_6
timestamp 1731220673
transform 1 0 192 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_590_6
timestamp 1731220673
transform 1 0 128 0 -1 1784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_589_6
timestamp 1731220673
transform 1 0 472 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_588_6
timestamp 1731220673
transform 1 0 368 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_587_6
timestamp 1731220673
transform 1 0 272 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_586_6
timestamp 1731220673
transform 1 0 184 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_585_6
timestamp 1731220673
transform 1 0 128 0 1 1796
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_584_6
timestamp 1731220673
transform 1 0 128 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_583_6
timestamp 1731220673
transform 1 0 184 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_582_6
timestamp 1731220673
transform 1 0 264 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_581_6
timestamp 1731220673
transform 1 0 448 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_580_6
timestamp 1731220673
transform 1 0 352 0 -1 1900
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_579_6
timestamp 1731220673
transform 1 0 296 0 1 1908
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_578_6
timestamp 1731220673
transform 1 0 192 0 1 1908
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_577_6
timestamp 1731220673
transform 1 0 128 0 1 1908
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_576_6
timestamp 1731220673
transform 1 0 560 0 1 1908
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_575_6
timestamp 1731220673
transform 1 0 416 0 1 1908
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_574_6
timestamp 1731220673
transform 1 0 352 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_573_6
timestamp 1731220673
transform 1 0 280 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_572_6
timestamp 1731220673
transform 1 0 224 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_571_6
timestamp 1731220673
transform 1 0 624 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_570_6
timestamp 1731220673
transform 1 0 528 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_569_6
timestamp 1731220673
transform 1 0 432 0 -1 2016
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_568_6
timestamp 1731220673
transform 1 0 376 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_567_6
timestamp 1731220673
transform 1 0 432 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_566_6
timestamp 1731220673
transform 1 0 488 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_565_6
timestamp 1731220673
transform 1 0 552 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_564_6
timestamp 1731220673
transform 1 0 616 0 1 2020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_563_6
timestamp 1731220673
transform 1 0 624 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_562_6
timestamp 1731220673
transform 1 0 552 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_561_6
timestamp 1731220673
transform 1 0 480 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_560_6
timestamp 1731220673
transform 1 0 416 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_559_6
timestamp 1731220673
transform 1 0 352 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_558_6
timestamp 1731220673
transform 1 0 296 0 -1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_557_6
timestamp 1731220673
transform 1 0 536 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_556_6
timestamp 1731220673
transform 1 0 432 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_555_6
timestamp 1731220673
transform 1 0 328 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_554_6
timestamp 1731220673
transform 1 0 232 0 1 2128
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_553_6
timestamp 1731220673
transform 1 0 512 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_552_6
timestamp 1731220673
transform 1 0 408 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_551_6
timestamp 1731220673
transform 1 0 312 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_550_6
timestamp 1731220673
transform 1 0 224 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_549_6
timestamp 1731220673
transform 1 0 136 0 -1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_548_6
timestamp 1731220673
transform 1 0 152 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_547_6
timestamp 1731220673
transform 1 0 248 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_546_6
timestamp 1731220673
transform 1 0 352 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_545_6
timestamp 1731220673
transform 1 0 568 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_544_6
timestamp 1731220673
transform 1 0 456 0 1 2232
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_543_6
timestamp 1731220673
transform 1 0 384 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_542_6
timestamp 1731220673
transform 1 0 312 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_541_6
timestamp 1731220673
transform 1 0 456 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_540_6
timestamp 1731220673
transform 1 0 528 0 -1 2344
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_539_6
timestamp 1731220673
transform 1 0 496 0 1 2352
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_538_6
timestamp 1731220673
transform 1 0 552 0 1 2352
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_537_6
timestamp 1731220673
transform 1 0 608 0 1 2352
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_536_6
timestamp 1731220673
transform 1 0 664 0 1 2352
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_535_6
timestamp 1731220673
transform 1 0 888 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_534_6
timestamp 1731220673
transform 1 0 944 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_533_6
timestamp 1731220673
transform 1 0 1000 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_532_6
timestamp 1731220673
transform 1 0 1056 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_531_6
timestamp 1731220673
transform 1 0 1040 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_530_6
timestamp 1731220673
transform 1 0 976 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_529_6
timestamp 1731220673
transform 1 0 912 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_528_6
timestamp 1731220673
transform 1 0 848 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_527_6
timestamp 1731220673
transform 1 0 784 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_526_6
timestamp 1731220673
transform 1 0 720 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_525_6
timestamp 1731220673
transform 1 0 656 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_524_6
timestamp 1731220673
transform 1 0 592 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_523_6
timestamp 1731220673
transform 1 0 528 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_522_6
timestamp 1731220673
transform 1 0 832 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_521_6
timestamp 1731220673
transform 1 0 776 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_520_6
timestamp 1731220673
transform 1 0 720 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_519_6
timestamp 1731220673
transform 1 0 664 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_518_6
timestamp 1731220673
transform 1 0 608 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_517_6
timestamp 1731220673
transform 1 0 552 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_516_6
timestamp 1731220673
transform 1 0 496 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_515_6
timestamp 1731220673
transform 1 0 440 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_514_6
timestamp 1731220673
transform 1 0 384 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_513_6
timestamp 1731220673
transform 1 0 328 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_512_6
timestamp 1731220673
transform 1 0 272 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_511_6
timestamp 1731220673
transform 1 0 216 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_510_6
timestamp 1731220673
transform 1 0 160 0 -1 2468
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_59_6
timestamp 1731220673
transform 1 0 464 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_58_6
timestamp 1731220673
transform 1 0 392 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_57_6
timestamp 1731220673
transform 1 0 320 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_56_6
timestamp 1731220673
transform 1 0 256 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_55_6
timestamp 1731220673
transform 1 0 200 0 1 2476
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_54_6
timestamp 1731220673
transform 1 0 352 0 -1 2580
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_53_6
timestamp 1731220673
transform 1 0 296 0 -1 2580
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_52_6
timestamp 1731220673
transform 1 0 240 0 -1 2580
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_51_6
timestamp 1731220673
transform 1 0 184 0 -1 2580
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_50_6
timestamp 1731220673
transform 1 0 128 0 -1 2580
box 4 4 48 48
<< end >>
