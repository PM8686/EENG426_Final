magic
tech sky130l
timestamp 1731220380
<< m2 >>
rect 550 2630 556 2631
rect 550 2626 551 2630
rect 555 2626 556 2630
rect 550 2625 556 2626
rect 606 2630 612 2631
rect 606 2626 607 2630
rect 611 2626 612 2630
rect 606 2625 612 2626
rect 662 2630 668 2631
rect 662 2626 663 2630
rect 667 2626 668 2630
rect 662 2625 668 2626
rect 718 2630 724 2631
rect 718 2626 719 2630
rect 723 2626 724 2630
rect 718 2625 724 2626
rect 774 2630 780 2631
rect 774 2626 775 2630
rect 779 2626 780 2630
rect 774 2625 780 2626
rect 1550 2626 1556 2627
rect 1550 2622 1551 2626
rect 1555 2622 1556 2626
rect 110 2621 116 2622
rect 110 2617 111 2621
rect 115 2617 116 2621
rect 110 2616 116 2617
rect 1326 2621 1332 2622
rect 1550 2621 1556 2622
rect 1606 2626 1612 2627
rect 1606 2622 1607 2626
rect 1611 2622 1612 2626
rect 1606 2621 1612 2622
rect 1662 2626 1668 2627
rect 1662 2622 1663 2626
rect 1667 2622 1668 2626
rect 1662 2621 1668 2622
rect 1718 2626 1724 2627
rect 1718 2622 1719 2626
rect 1723 2622 1724 2626
rect 1718 2621 1724 2622
rect 1774 2626 1780 2627
rect 1774 2622 1775 2626
rect 1779 2622 1780 2626
rect 1774 2621 1780 2622
rect 1830 2626 1836 2627
rect 1830 2622 1831 2626
rect 1835 2622 1836 2626
rect 1830 2621 1836 2622
rect 1886 2626 1892 2627
rect 1886 2622 1887 2626
rect 1891 2622 1892 2626
rect 1886 2621 1892 2622
rect 1942 2626 1948 2627
rect 1942 2622 1943 2626
rect 1947 2622 1948 2626
rect 1942 2621 1948 2622
rect 1998 2626 2004 2627
rect 1998 2622 1999 2626
rect 2003 2622 2004 2626
rect 1998 2621 2004 2622
rect 2054 2626 2060 2627
rect 2054 2622 2055 2626
rect 2059 2622 2060 2626
rect 2054 2621 2060 2622
rect 2110 2626 2116 2627
rect 2110 2622 2111 2626
rect 2115 2622 2116 2626
rect 2110 2621 2116 2622
rect 2166 2626 2172 2627
rect 2166 2622 2167 2626
rect 2171 2622 2172 2626
rect 2166 2621 2172 2622
rect 1326 2617 1327 2621
rect 1331 2617 1332 2621
rect 1326 2616 1332 2617
rect 1366 2617 1372 2618
rect 1366 2613 1367 2617
rect 1371 2613 1372 2617
rect 1366 2612 1372 2613
rect 2582 2617 2588 2618
rect 2582 2613 2583 2617
rect 2587 2613 2588 2617
rect 2582 2612 2588 2613
rect 110 2604 116 2605
rect 1326 2604 1332 2605
rect 110 2600 111 2604
rect 115 2600 116 2604
rect 110 2599 116 2600
rect 534 2603 540 2604
rect 534 2599 535 2603
rect 539 2599 540 2603
rect 534 2598 540 2599
rect 590 2603 596 2604
rect 590 2599 591 2603
rect 595 2599 596 2603
rect 590 2598 596 2599
rect 646 2603 652 2604
rect 646 2599 647 2603
rect 651 2599 652 2603
rect 646 2598 652 2599
rect 702 2603 708 2604
rect 702 2599 703 2603
rect 707 2599 708 2603
rect 702 2598 708 2599
rect 758 2603 764 2604
rect 758 2599 759 2603
rect 763 2599 764 2603
rect 1326 2600 1327 2604
rect 1331 2600 1332 2604
rect 1326 2599 1332 2600
rect 1366 2600 1372 2601
rect 2582 2600 2588 2601
rect 758 2598 764 2599
rect 1366 2596 1367 2600
rect 1371 2596 1372 2600
rect 1366 2595 1372 2596
rect 1534 2599 1540 2600
rect 1534 2595 1535 2599
rect 1539 2595 1540 2599
rect 1534 2594 1540 2595
rect 1590 2599 1596 2600
rect 1590 2595 1591 2599
rect 1595 2595 1596 2599
rect 1590 2594 1596 2595
rect 1646 2599 1652 2600
rect 1646 2595 1647 2599
rect 1651 2595 1652 2599
rect 1646 2594 1652 2595
rect 1702 2599 1708 2600
rect 1702 2595 1703 2599
rect 1707 2595 1708 2599
rect 1702 2594 1708 2595
rect 1758 2599 1764 2600
rect 1758 2595 1759 2599
rect 1763 2595 1764 2599
rect 1758 2594 1764 2595
rect 1814 2599 1820 2600
rect 1814 2595 1815 2599
rect 1819 2595 1820 2599
rect 1814 2594 1820 2595
rect 1870 2599 1876 2600
rect 1870 2595 1871 2599
rect 1875 2595 1876 2599
rect 1870 2594 1876 2595
rect 1926 2599 1932 2600
rect 1926 2595 1927 2599
rect 1931 2595 1932 2599
rect 1926 2594 1932 2595
rect 1982 2599 1988 2600
rect 1982 2595 1983 2599
rect 1987 2595 1988 2599
rect 1982 2594 1988 2595
rect 2038 2599 2044 2600
rect 2038 2595 2039 2599
rect 2043 2595 2044 2599
rect 2038 2594 2044 2595
rect 2094 2599 2100 2600
rect 2094 2595 2095 2599
rect 2099 2595 2100 2599
rect 2094 2594 2100 2595
rect 2150 2599 2156 2600
rect 2150 2595 2151 2599
rect 2155 2595 2156 2599
rect 2582 2596 2583 2600
rect 2587 2596 2588 2600
rect 2582 2595 2588 2596
rect 2150 2594 2156 2595
rect 214 2569 220 2570
rect 110 2568 116 2569
rect 110 2564 111 2568
rect 115 2564 116 2568
rect 214 2565 215 2569
rect 219 2565 220 2569
rect 214 2564 220 2565
rect 270 2569 276 2570
rect 270 2565 271 2569
rect 275 2565 276 2569
rect 270 2564 276 2565
rect 326 2569 332 2570
rect 326 2565 327 2569
rect 331 2565 332 2569
rect 326 2564 332 2565
rect 382 2569 388 2570
rect 382 2565 383 2569
rect 387 2565 388 2569
rect 382 2564 388 2565
rect 438 2569 444 2570
rect 438 2565 439 2569
rect 443 2565 444 2569
rect 438 2564 444 2565
rect 494 2569 500 2570
rect 494 2565 495 2569
rect 499 2565 500 2569
rect 494 2564 500 2565
rect 550 2569 556 2570
rect 550 2565 551 2569
rect 555 2565 556 2569
rect 550 2564 556 2565
rect 606 2569 612 2570
rect 606 2565 607 2569
rect 611 2565 612 2569
rect 606 2564 612 2565
rect 662 2569 668 2570
rect 662 2565 663 2569
rect 667 2565 668 2569
rect 662 2564 668 2565
rect 718 2569 724 2570
rect 718 2565 719 2569
rect 723 2565 724 2569
rect 718 2564 724 2565
rect 774 2569 780 2570
rect 774 2565 775 2569
rect 779 2565 780 2569
rect 774 2564 780 2565
rect 830 2569 836 2570
rect 830 2565 831 2569
rect 835 2565 836 2569
rect 830 2564 836 2565
rect 886 2569 892 2570
rect 886 2565 887 2569
rect 891 2565 892 2569
rect 886 2564 892 2565
rect 942 2569 948 2570
rect 942 2565 943 2569
rect 947 2565 948 2569
rect 942 2564 948 2565
rect 998 2569 1004 2570
rect 998 2565 999 2569
rect 1003 2565 1004 2569
rect 998 2564 1004 2565
rect 1054 2569 1060 2570
rect 1054 2565 1055 2569
rect 1059 2565 1060 2569
rect 1054 2564 1060 2565
rect 1110 2569 1116 2570
rect 1110 2565 1111 2569
rect 1115 2565 1116 2569
rect 1110 2564 1116 2565
rect 1326 2568 1332 2569
rect 1326 2564 1327 2568
rect 1331 2564 1332 2568
rect 1438 2565 1444 2566
rect 110 2563 116 2564
rect 1326 2563 1332 2564
rect 1366 2564 1372 2565
rect 1366 2560 1367 2564
rect 1371 2560 1372 2564
rect 1438 2561 1439 2565
rect 1443 2561 1444 2565
rect 1438 2560 1444 2561
rect 1542 2565 1548 2566
rect 1542 2561 1543 2565
rect 1547 2561 1548 2565
rect 1542 2560 1548 2561
rect 1654 2565 1660 2566
rect 1654 2561 1655 2565
rect 1659 2561 1660 2565
rect 1654 2560 1660 2561
rect 1766 2565 1772 2566
rect 1766 2561 1767 2565
rect 1771 2561 1772 2565
rect 1766 2560 1772 2561
rect 1878 2565 1884 2566
rect 1878 2561 1879 2565
rect 1883 2561 1884 2565
rect 1878 2560 1884 2561
rect 1990 2565 1996 2566
rect 1990 2561 1991 2565
rect 1995 2561 1996 2565
rect 1990 2560 1996 2561
rect 2110 2565 2116 2566
rect 2110 2561 2111 2565
rect 2115 2561 2116 2565
rect 2110 2560 2116 2561
rect 2230 2565 2236 2566
rect 2230 2561 2231 2565
rect 2235 2561 2236 2565
rect 2230 2560 2236 2561
rect 2350 2565 2356 2566
rect 2350 2561 2351 2565
rect 2355 2561 2356 2565
rect 2350 2560 2356 2561
rect 2582 2564 2588 2565
rect 2582 2560 2583 2564
rect 2587 2560 2588 2564
rect 1366 2559 1372 2560
rect 2582 2559 2588 2560
rect 110 2551 116 2552
rect 110 2547 111 2551
rect 115 2547 116 2551
rect 110 2546 116 2547
rect 1326 2551 1332 2552
rect 1326 2547 1327 2551
rect 1331 2547 1332 2551
rect 1326 2546 1332 2547
rect 1366 2547 1372 2548
rect 1366 2543 1367 2547
rect 1371 2543 1372 2547
rect 230 2542 236 2543
rect 230 2538 231 2542
rect 235 2538 236 2542
rect 230 2537 236 2538
rect 286 2542 292 2543
rect 286 2538 287 2542
rect 291 2538 292 2542
rect 286 2537 292 2538
rect 342 2542 348 2543
rect 342 2538 343 2542
rect 347 2538 348 2542
rect 342 2537 348 2538
rect 398 2542 404 2543
rect 398 2538 399 2542
rect 403 2538 404 2542
rect 398 2537 404 2538
rect 454 2542 460 2543
rect 454 2538 455 2542
rect 459 2538 460 2542
rect 454 2537 460 2538
rect 510 2542 516 2543
rect 510 2538 511 2542
rect 515 2538 516 2542
rect 510 2537 516 2538
rect 566 2542 572 2543
rect 566 2538 567 2542
rect 571 2538 572 2542
rect 566 2537 572 2538
rect 622 2542 628 2543
rect 622 2538 623 2542
rect 627 2538 628 2542
rect 622 2537 628 2538
rect 678 2542 684 2543
rect 678 2538 679 2542
rect 683 2538 684 2542
rect 678 2537 684 2538
rect 734 2542 740 2543
rect 734 2538 735 2542
rect 739 2538 740 2542
rect 734 2537 740 2538
rect 790 2542 796 2543
rect 790 2538 791 2542
rect 795 2538 796 2542
rect 790 2537 796 2538
rect 846 2542 852 2543
rect 846 2538 847 2542
rect 851 2538 852 2542
rect 846 2537 852 2538
rect 902 2542 908 2543
rect 902 2538 903 2542
rect 907 2538 908 2542
rect 902 2537 908 2538
rect 958 2542 964 2543
rect 958 2538 959 2542
rect 963 2538 964 2542
rect 958 2537 964 2538
rect 1014 2542 1020 2543
rect 1014 2538 1015 2542
rect 1019 2538 1020 2542
rect 1014 2537 1020 2538
rect 1070 2542 1076 2543
rect 1070 2538 1071 2542
rect 1075 2538 1076 2542
rect 1070 2537 1076 2538
rect 1126 2542 1132 2543
rect 1366 2542 1372 2543
rect 2582 2547 2588 2548
rect 2582 2543 2583 2547
rect 2587 2543 2588 2547
rect 2582 2542 2588 2543
rect 1126 2538 1127 2542
rect 1131 2538 1132 2542
rect 1126 2537 1132 2538
rect 1454 2538 1460 2539
rect 1454 2534 1455 2538
rect 1459 2534 1460 2538
rect 1454 2533 1460 2534
rect 1558 2538 1564 2539
rect 1558 2534 1559 2538
rect 1563 2534 1564 2538
rect 1558 2533 1564 2534
rect 1670 2538 1676 2539
rect 1670 2534 1671 2538
rect 1675 2534 1676 2538
rect 1670 2533 1676 2534
rect 1782 2538 1788 2539
rect 1782 2534 1783 2538
rect 1787 2534 1788 2538
rect 1782 2533 1788 2534
rect 1894 2538 1900 2539
rect 1894 2534 1895 2538
rect 1899 2534 1900 2538
rect 1894 2533 1900 2534
rect 2006 2538 2012 2539
rect 2006 2534 2007 2538
rect 2011 2534 2012 2538
rect 2006 2533 2012 2534
rect 2126 2538 2132 2539
rect 2126 2534 2127 2538
rect 2131 2534 2132 2538
rect 2126 2533 2132 2534
rect 2246 2538 2252 2539
rect 2246 2534 2247 2538
rect 2251 2534 2252 2538
rect 2246 2533 2252 2534
rect 2366 2538 2372 2539
rect 2366 2534 2367 2538
rect 2371 2534 2372 2538
rect 2366 2533 2372 2534
rect 366 2514 372 2515
rect 366 2510 367 2514
rect 371 2510 372 2514
rect 366 2509 372 2510
rect 422 2514 428 2515
rect 422 2510 423 2514
rect 427 2510 428 2514
rect 422 2509 428 2510
rect 486 2514 492 2515
rect 486 2510 487 2514
rect 491 2510 492 2514
rect 486 2509 492 2510
rect 550 2514 556 2515
rect 550 2510 551 2514
rect 555 2510 556 2514
rect 550 2509 556 2510
rect 614 2514 620 2515
rect 614 2510 615 2514
rect 619 2510 620 2514
rect 614 2509 620 2510
rect 678 2514 684 2515
rect 678 2510 679 2514
rect 683 2510 684 2514
rect 678 2509 684 2510
rect 742 2514 748 2515
rect 742 2510 743 2514
rect 747 2510 748 2514
rect 742 2509 748 2510
rect 806 2514 812 2515
rect 806 2510 807 2514
rect 811 2510 812 2514
rect 806 2509 812 2510
rect 870 2514 876 2515
rect 870 2510 871 2514
rect 875 2510 876 2514
rect 870 2509 876 2510
rect 942 2514 948 2515
rect 942 2510 943 2514
rect 947 2510 948 2514
rect 942 2509 948 2510
rect 1014 2514 1020 2515
rect 1014 2510 1015 2514
rect 1019 2510 1020 2514
rect 1014 2509 1020 2510
rect 1550 2506 1556 2507
rect 110 2505 116 2506
rect 110 2501 111 2505
rect 115 2501 116 2505
rect 110 2500 116 2501
rect 1326 2505 1332 2506
rect 1326 2501 1327 2505
rect 1331 2501 1332 2505
rect 1550 2502 1551 2506
rect 1555 2502 1556 2506
rect 1550 2501 1556 2502
rect 1630 2506 1636 2507
rect 1630 2502 1631 2506
rect 1635 2502 1636 2506
rect 1630 2501 1636 2502
rect 1718 2506 1724 2507
rect 1718 2502 1719 2506
rect 1723 2502 1724 2506
rect 1718 2501 1724 2502
rect 1806 2506 1812 2507
rect 1806 2502 1807 2506
rect 1811 2502 1812 2506
rect 1806 2501 1812 2502
rect 1902 2506 1908 2507
rect 1902 2502 1903 2506
rect 1907 2502 1908 2506
rect 1902 2501 1908 2502
rect 1998 2506 2004 2507
rect 1998 2502 1999 2506
rect 2003 2502 2004 2506
rect 1998 2501 2004 2502
rect 2094 2506 2100 2507
rect 2094 2502 2095 2506
rect 2099 2502 2100 2506
rect 2094 2501 2100 2502
rect 2190 2506 2196 2507
rect 2190 2502 2191 2506
rect 2195 2502 2196 2506
rect 2190 2501 2196 2502
rect 2294 2506 2300 2507
rect 2294 2502 2295 2506
rect 2299 2502 2300 2506
rect 2294 2501 2300 2502
rect 2398 2506 2404 2507
rect 2398 2502 2399 2506
rect 2403 2502 2404 2506
rect 2398 2501 2404 2502
rect 1326 2500 1332 2501
rect 1366 2497 1372 2498
rect 1366 2493 1367 2497
rect 1371 2493 1372 2497
rect 1366 2492 1372 2493
rect 2582 2497 2588 2498
rect 2582 2493 2583 2497
rect 2587 2493 2588 2497
rect 2582 2492 2588 2493
rect 110 2488 116 2489
rect 1326 2488 1332 2489
rect 110 2484 111 2488
rect 115 2484 116 2488
rect 110 2483 116 2484
rect 350 2487 356 2488
rect 350 2483 351 2487
rect 355 2483 356 2487
rect 350 2482 356 2483
rect 406 2487 412 2488
rect 406 2483 407 2487
rect 411 2483 412 2487
rect 406 2482 412 2483
rect 470 2487 476 2488
rect 470 2483 471 2487
rect 475 2483 476 2487
rect 470 2482 476 2483
rect 534 2487 540 2488
rect 534 2483 535 2487
rect 539 2483 540 2487
rect 534 2482 540 2483
rect 598 2487 604 2488
rect 598 2483 599 2487
rect 603 2483 604 2487
rect 598 2482 604 2483
rect 662 2487 668 2488
rect 662 2483 663 2487
rect 667 2483 668 2487
rect 662 2482 668 2483
rect 726 2487 732 2488
rect 726 2483 727 2487
rect 731 2483 732 2487
rect 726 2482 732 2483
rect 790 2487 796 2488
rect 790 2483 791 2487
rect 795 2483 796 2487
rect 790 2482 796 2483
rect 854 2487 860 2488
rect 854 2483 855 2487
rect 859 2483 860 2487
rect 854 2482 860 2483
rect 926 2487 932 2488
rect 926 2483 927 2487
rect 931 2483 932 2487
rect 926 2482 932 2483
rect 998 2487 1004 2488
rect 998 2483 999 2487
rect 1003 2483 1004 2487
rect 1326 2484 1327 2488
rect 1331 2484 1332 2488
rect 1326 2483 1332 2484
rect 998 2482 1004 2483
rect 1366 2480 1372 2481
rect 2582 2480 2588 2481
rect 1366 2476 1367 2480
rect 1371 2476 1372 2480
rect 1366 2475 1372 2476
rect 1534 2479 1540 2480
rect 1534 2475 1535 2479
rect 1539 2475 1540 2479
rect 1534 2474 1540 2475
rect 1614 2479 1620 2480
rect 1614 2475 1615 2479
rect 1619 2475 1620 2479
rect 1614 2474 1620 2475
rect 1702 2479 1708 2480
rect 1702 2475 1703 2479
rect 1707 2475 1708 2479
rect 1702 2474 1708 2475
rect 1790 2479 1796 2480
rect 1790 2475 1791 2479
rect 1795 2475 1796 2479
rect 1790 2474 1796 2475
rect 1886 2479 1892 2480
rect 1886 2475 1887 2479
rect 1891 2475 1892 2479
rect 1886 2474 1892 2475
rect 1982 2479 1988 2480
rect 1982 2475 1983 2479
rect 1987 2475 1988 2479
rect 1982 2474 1988 2475
rect 2078 2479 2084 2480
rect 2078 2475 2079 2479
rect 2083 2475 2084 2479
rect 2078 2474 2084 2475
rect 2174 2479 2180 2480
rect 2174 2475 2175 2479
rect 2179 2475 2180 2479
rect 2174 2474 2180 2475
rect 2278 2479 2284 2480
rect 2278 2475 2279 2479
rect 2283 2475 2284 2479
rect 2278 2474 2284 2475
rect 2382 2479 2388 2480
rect 2382 2475 2383 2479
rect 2387 2475 2388 2479
rect 2582 2476 2583 2480
rect 2587 2476 2588 2480
rect 2582 2475 2588 2476
rect 2382 2474 2388 2475
rect 270 2449 276 2450
rect 110 2448 116 2449
rect 110 2444 111 2448
rect 115 2444 116 2448
rect 270 2445 271 2449
rect 275 2445 276 2449
rect 270 2444 276 2445
rect 334 2449 340 2450
rect 334 2445 335 2449
rect 339 2445 340 2449
rect 334 2444 340 2445
rect 398 2449 404 2450
rect 398 2445 399 2449
rect 403 2445 404 2449
rect 398 2444 404 2445
rect 470 2449 476 2450
rect 470 2445 471 2449
rect 475 2445 476 2449
rect 470 2444 476 2445
rect 550 2449 556 2450
rect 550 2445 551 2449
rect 555 2445 556 2449
rect 550 2444 556 2445
rect 630 2449 636 2450
rect 630 2445 631 2449
rect 635 2445 636 2449
rect 630 2444 636 2445
rect 710 2449 716 2450
rect 710 2445 711 2449
rect 715 2445 716 2449
rect 710 2444 716 2445
rect 782 2449 788 2450
rect 782 2445 783 2449
rect 787 2445 788 2449
rect 782 2444 788 2445
rect 862 2449 868 2450
rect 862 2445 863 2449
rect 867 2445 868 2449
rect 862 2444 868 2445
rect 942 2449 948 2450
rect 942 2445 943 2449
rect 947 2445 948 2449
rect 942 2444 948 2445
rect 1022 2449 1028 2450
rect 1022 2445 1023 2449
rect 1027 2445 1028 2449
rect 1022 2444 1028 2445
rect 1326 2448 1332 2449
rect 1326 2444 1327 2448
rect 1331 2444 1332 2448
rect 1646 2445 1652 2446
rect 110 2443 116 2444
rect 1326 2443 1332 2444
rect 1366 2444 1372 2445
rect 1366 2440 1367 2444
rect 1371 2440 1372 2444
rect 1646 2441 1647 2445
rect 1651 2441 1652 2445
rect 1646 2440 1652 2441
rect 1702 2445 1708 2446
rect 1702 2441 1703 2445
rect 1707 2441 1708 2445
rect 1702 2440 1708 2441
rect 1766 2445 1772 2446
rect 1766 2441 1767 2445
rect 1771 2441 1772 2445
rect 1766 2440 1772 2441
rect 1838 2445 1844 2446
rect 1838 2441 1839 2445
rect 1843 2441 1844 2445
rect 1838 2440 1844 2441
rect 1910 2445 1916 2446
rect 1910 2441 1911 2445
rect 1915 2441 1916 2445
rect 1910 2440 1916 2441
rect 1990 2445 1996 2446
rect 1990 2441 1991 2445
rect 1995 2441 1996 2445
rect 1990 2440 1996 2441
rect 2078 2445 2084 2446
rect 2078 2441 2079 2445
rect 2083 2441 2084 2445
rect 2078 2440 2084 2441
rect 2166 2445 2172 2446
rect 2166 2441 2167 2445
rect 2171 2441 2172 2445
rect 2166 2440 2172 2441
rect 2262 2445 2268 2446
rect 2262 2441 2263 2445
rect 2267 2441 2268 2445
rect 2262 2440 2268 2441
rect 2358 2445 2364 2446
rect 2358 2441 2359 2445
rect 2363 2441 2364 2445
rect 2358 2440 2364 2441
rect 2454 2445 2460 2446
rect 2454 2441 2455 2445
rect 2459 2441 2460 2445
rect 2454 2440 2460 2441
rect 2526 2445 2532 2446
rect 2526 2441 2527 2445
rect 2531 2441 2532 2445
rect 2526 2440 2532 2441
rect 2582 2444 2588 2445
rect 2582 2440 2583 2444
rect 2587 2440 2588 2444
rect 1366 2439 1372 2440
rect 2582 2439 2588 2440
rect 110 2431 116 2432
rect 110 2427 111 2431
rect 115 2427 116 2431
rect 110 2426 116 2427
rect 1326 2431 1332 2432
rect 1326 2427 1327 2431
rect 1331 2427 1332 2431
rect 1326 2426 1332 2427
rect 1366 2427 1372 2428
rect 1366 2423 1367 2427
rect 1371 2423 1372 2427
rect 286 2422 292 2423
rect 286 2418 287 2422
rect 291 2418 292 2422
rect 286 2417 292 2418
rect 350 2422 356 2423
rect 350 2418 351 2422
rect 355 2418 356 2422
rect 350 2417 356 2418
rect 414 2422 420 2423
rect 414 2418 415 2422
rect 419 2418 420 2422
rect 414 2417 420 2418
rect 486 2422 492 2423
rect 486 2418 487 2422
rect 491 2418 492 2422
rect 486 2417 492 2418
rect 566 2422 572 2423
rect 566 2418 567 2422
rect 571 2418 572 2422
rect 566 2417 572 2418
rect 646 2422 652 2423
rect 646 2418 647 2422
rect 651 2418 652 2422
rect 646 2417 652 2418
rect 726 2422 732 2423
rect 726 2418 727 2422
rect 731 2418 732 2422
rect 726 2417 732 2418
rect 798 2422 804 2423
rect 798 2418 799 2422
rect 803 2418 804 2422
rect 798 2417 804 2418
rect 878 2422 884 2423
rect 878 2418 879 2422
rect 883 2418 884 2422
rect 878 2417 884 2418
rect 958 2422 964 2423
rect 958 2418 959 2422
rect 963 2418 964 2422
rect 958 2417 964 2418
rect 1038 2422 1044 2423
rect 1366 2422 1372 2423
rect 2582 2427 2588 2428
rect 2582 2423 2583 2427
rect 2587 2423 2588 2427
rect 2582 2422 2588 2423
rect 1038 2418 1039 2422
rect 1043 2418 1044 2422
rect 1038 2417 1044 2418
rect 1662 2418 1668 2419
rect 1662 2414 1663 2418
rect 1667 2414 1668 2418
rect 1662 2413 1668 2414
rect 1718 2418 1724 2419
rect 1718 2414 1719 2418
rect 1723 2414 1724 2418
rect 1718 2413 1724 2414
rect 1782 2418 1788 2419
rect 1782 2414 1783 2418
rect 1787 2414 1788 2418
rect 1782 2413 1788 2414
rect 1854 2418 1860 2419
rect 1854 2414 1855 2418
rect 1859 2414 1860 2418
rect 1854 2413 1860 2414
rect 1926 2418 1932 2419
rect 1926 2414 1927 2418
rect 1931 2414 1932 2418
rect 1926 2413 1932 2414
rect 2006 2418 2012 2419
rect 2006 2414 2007 2418
rect 2011 2414 2012 2418
rect 2006 2413 2012 2414
rect 2094 2418 2100 2419
rect 2094 2414 2095 2418
rect 2099 2414 2100 2418
rect 2094 2413 2100 2414
rect 2182 2418 2188 2419
rect 2182 2414 2183 2418
rect 2187 2414 2188 2418
rect 2182 2413 2188 2414
rect 2278 2418 2284 2419
rect 2278 2414 2279 2418
rect 2283 2414 2284 2418
rect 2278 2413 2284 2414
rect 2374 2418 2380 2419
rect 2374 2414 2375 2418
rect 2379 2414 2380 2418
rect 2374 2413 2380 2414
rect 2470 2418 2476 2419
rect 2470 2414 2471 2418
rect 2475 2414 2476 2418
rect 2470 2413 2476 2414
rect 2542 2418 2548 2419
rect 2542 2414 2543 2418
rect 2547 2414 2548 2418
rect 2542 2413 2548 2414
rect 246 2394 252 2395
rect 246 2390 247 2394
rect 251 2390 252 2394
rect 246 2389 252 2390
rect 334 2394 340 2395
rect 334 2390 335 2394
rect 339 2390 340 2394
rect 334 2389 340 2390
rect 430 2394 436 2395
rect 430 2390 431 2394
rect 435 2390 436 2394
rect 430 2389 436 2390
rect 526 2394 532 2395
rect 526 2390 527 2394
rect 531 2390 532 2394
rect 526 2389 532 2390
rect 630 2394 636 2395
rect 630 2390 631 2394
rect 635 2390 636 2394
rect 630 2389 636 2390
rect 726 2394 732 2395
rect 726 2390 727 2394
rect 731 2390 732 2394
rect 726 2389 732 2390
rect 822 2394 828 2395
rect 822 2390 823 2394
rect 827 2390 828 2394
rect 822 2389 828 2390
rect 918 2394 924 2395
rect 918 2390 919 2394
rect 923 2390 924 2394
rect 918 2389 924 2390
rect 1014 2394 1020 2395
rect 1014 2390 1015 2394
rect 1019 2390 1020 2394
rect 1014 2389 1020 2390
rect 1110 2394 1116 2395
rect 1110 2390 1111 2394
rect 1115 2390 1116 2394
rect 1110 2389 1116 2390
rect 1454 2390 1460 2391
rect 1454 2386 1455 2390
rect 1459 2386 1460 2390
rect 110 2385 116 2386
rect 110 2381 111 2385
rect 115 2381 116 2385
rect 110 2380 116 2381
rect 1326 2385 1332 2386
rect 1454 2385 1460 2386
rect 1558 2390 1564 2391
rect 1558 2386 1559 2390
rect 1563 2386 1564 2390
rect 1558 2385 1564 2386
rect 1662 2390 1668 2391
rect 1662 2386 1663 2390
rect 1667 2386 1668 2390
rect 1662 2385 1668 2386
rect 1758 2390 1764 2391
rect 1758 2386 1759 2390
rect 1763 2386 1764 2390
rect 1758 2385 1764 2386
rect 1854 2390 1860 2391
rect 1854 2386 1855 2390
rect 1859 2386 1860 2390
rect 1854 2385 1860 2386
rect 1942 2390 1948 2391
rect 1942 2386 1943 2390
rect 1947 2386 1948 2390
rect 1942 2385 1948 2386
rect 2038 2390 2044 2391
rect 2038 2386 2039 2390
rect 2043 2386 2044 2390
rect 2038 2385 2044 2386
rect 2134 2390 2140 2391
rect 2134 2386 2135 2390
rect 2139 2386 2140 2390
rect 2134 2385 2140 2386
rect 2230 2390 2236 2391
rect 2230 2386 2231 2390
rect 2235 2386 2236 2390
rect 2230 2385 2236 2386
rect 2334 2390 2340 2391
rect 2334 2386 2335 2390
rect 2339 2386 2340 2390
rect 2334 2385 2340 2386
rect 2446 2390 2452 2391
rect 2446 2386 2447 2390
rect 2451 2386 2452 2390
rect 2446 2385 2452 2386
rect 2542 2390 2548 2391
rect 2542 2386 2543 2390
rect 2547 2386 2548 2390
rect 2542 2385 2548 2386
rect 1326 2381 1327 2385
rect 1331 2381 1332 2385
rect 1326 2380 1332 2381
rect 1366 2381 1372 2382
rect 1366 2377 1367 2381
rect 1371 2377 1372 2381
rect 1366 2376 1372 2377
rect 2582 2381 2588 2382
rect 2582 2377 2583 2381
rect 2587 2377 2588 2381
rect 2582 2376 2588 2377
rect 110 2368 116 2369
rect 1326 2368 1332 2369
rect 110 2364 111 2368
rect 115 2364 116 2368
rect 110 2363 116 2364
rect 230 2367 236 2368
rect 230 2363 231 2367
rect 235 2363 236 2367
rect 230 2362 236 2363
rect 318 2367 324 2368
rect 318 2363 319 2367
rect 323 2363 324 2367
rect 318 2362 324 2363
rect 414 2367 420 2368
rect 414 2363 415 2367
rect 419 2363 420 2367
rect 414 2362 420 2363
rect 510 2367 516 2368
rect 510 2363 511 2367
rect 515 2363 516 2367
rect 510 2362 516 2363
rect 614 2367 620 2368
rect 614 2363 615 2367
rect 619 2363 620 2367
rect 614 2362 620 2363
rect 710 2367 716 2368
rect 710 2363 711 2367
rect 715 2363 716 2367
rect 710 2362 716 2363
rect 806 2367 812 2368
rect 806 2363 807 2367
rect 811 2363 812 2367
rect 806 2362 812 2363
rect 902 2367 908 2368
rect 902 2363 903 2367
rect 907 2363 908 2367
rect 902 2362 908 2363
rect 998 2367 1004 2368
rect 998 2363 999 2367
rect 1003 2363 1004 2367
rect 998 2362 1004 2363
rect 1094 2367 1100 2368
rect 1094 2363 1095 2367
rect 1099 2363 1100 2367
rect 1326 2364 1327 2368
rect 1331 2364 1332 2368
rect 1326 2363 1332 2364
rect 1366 2364 1372 2365
rect 2582 2364 2588 2365
rect 1094 2362 1100 2363
rect 1366 2360 1367 2364
rect 1371 2360 1372 2364
rect 1366 2359 1372 2360
rect 1438 2363 1444 2364
rect 1438 2359 1439 2363
rect 1443 2359 1444 2363
rect 1438 2358 1444 2359
rect 1542 2363 1548 2364
rect 1542 2359 1543 2363
rect 1547 2359 1548 2363
rect 1542 2358 1548 2359
rect 1646 2363 1652 2364
rect 1646 2359 1647 2363
rect 1651 2359 1652 2363
rect 1646 2358 1652 2359
rect 1742 2363 1748 2364
rect 1742 2359 1743 2363
rect 1747 2359 1748 2363
rect 1742 2358 1748 2359
rect 1838 2363 1844 2364
rect 1838 2359 1839 2363
rect 1843 2359 1844 2363
rect 1838 2358 1844 2359
rect 1926 2363 1932 2364
rect 1926 2359 1927 2363
rect 1931 2359 1932 2363
rect 1926 2358 1932 2359
rect 2022 2363 2028 2364
rect 2022 2359 2023 2363
rect 2027 2359 2028 2363
rect 2022 2358 2028 2359
rect 2118 2363 2124 2364
rect 2118 2359 2119 2363
rect 2123 2359 2124 2363
rect 2118 2358 2124 2359
rect 2214 2363 2220 2364
rect 2214 2359 2215 2363
rect 2219 2359 2220 2363
rect 2214 2358 2220 2359
rect 2318 2363 2324 2364
rect 2318 2359 2319 2363
rect 2323 2359 2324 2363
rect 2318 2358 2324 2359
rect 2430 2363 2436 2364
rect 2430 2359 2431 2363
rect 2435 2359 2436 2363
rect 2430 2358 2436 2359
rect 2526 2363 2532 2364
rect 2526 2359 2527 2363
rect 2531 2359 2532 2363
rect 2582 2360 2583 2364
rect 2587 2360 2588 2364
rect 2582 2359 2588 2360
rect 2526 2358 2532 2359
rect 158 2333 164 2334
rect 110 2332 116 2333
rect 110 2328 111 2332
rect 115 2328 116 2332
rect 158 2329 159 2333
rect 163 2329 164 2333
rect 158 2328 164 2329
rect 262 2333 268 2334
rect 262 2329 263 2333
rect 267 2329 268 2333
rect 262 2328 268 2329
rect 374 2333 380 2334
rect 374 2329 375 2333
rect 379 2329 380 2333
rect 374 2328 380 2329
rect 486 2333 492 2334
rect 486 2329 487 2333
rect 491 2329 492 2333
rect 486 2328 492 2329
rect 598 2333 604 2334
rect 598 2329 599 2333
rect 603 2329 604 2333
rect 598 2328 604 2329
rect 710 2333 716 2334
rect 710 2329 711 2333
rect 715 2329 716 2333
rect 710 2328 716 2329
rect 814 2333 820 2334
rect 814 2329 815 2333
rect 819 2329 820 2333
rect 814 2328 820 2329
rect 910 2333 916 2334
rect 910 2329 911 2333
rect 915 2329 916 2333
rect 910 2328 916 2329
rect 1006 2333 1012 2334
rect 1006 2329 1007 2333
rect 1011 2329 1012 2333
rect 1006 2328 1012 2329
rect 1102 2333 1108 2334
rect 1102 2329 1103 2333
rect 1107 2329 1108 2333
rect 1102 2328 1108 2329
rect 1198 2333 1204 2334
rect 1198 2329 1199 2333
rect 1203 2329 1204 2333
rect 1198 2328 1204 2329
rect 1326 2332 1332 2333
rect 1326 2328 1327 2332
rect 1331 2328 1332 2332
rect 1398 2329 1404 2330
rect 110 2327 116 2328
rect 1326 2327 1332 2328
rect 1366 2328 1372 2329
rect 1366 2324 1367 2328
rect 1371 2324 1372 2328
rect 1398 2325 1399 2329
rect 1403 2325 1404 2329
rect 1398 2324 1404 2325
rect 1454 2329 1460 2330
rect 1454 2325 1455 2329
rect 1459 2325 1460 2329
rect 1454 2324 1460 2325
rect 1510 2329 1516 2330
rect 1510 2325 1511 2329
rect 1515 2325 1516 2329
rect 1510 2324 1516 2325
rect 1566 2329 1572 2330
rect 1566 2325 1567 2329
rect 1571 2325 1572 2329
rect 1566 2324 1572 2325
rect 1638 2329 1644 2330
rect 1638 2325 1639 2329
rect 1643 2325 1644 2329
rect 1638 2324 1644 2325
rect 1726 2329 1732 2330
rect 1726 2325 1727 2329
rect 1731 2325 1732 2329
rect 1726 2324 1732 2325
rect 1822 2329 1828 2330
rect 1822 2325 1823 2329
rect 1827 2325 1828 2329
rect 1822 2324 1828 2325
rect 1942 2329 1948 2330
rect 1942 2325 1943 2329
rect 1947 2325 1948 2329
rect 1942 2324 1948 2325
rect 2078 2329 2084 2330
rect 2078 2325 2079 2329
rect 2083 2325 2084 2329
rect 2078 2324 2084 2325
rect 2222 2329 2228 2330
rect 2222 2325 2223 2329
rect 2227 2325 2228 2329
rect 2222 2324 2228 2325
rect 2382 2329 2388 2330
rect 2382 2325 2383 2329
rect 2387 2325 2388 2329
rect 2382 2324 2388 2325
rect 2526 2329 2532 2330
rect 2526 2325 2527 2329
rect 2531 2325 2532 2329
rect 2526 2324 2532 2325
rect 2582 2328 2588 2329
rect 2582 2324 2583 2328
rect 2587 2324 2588 2328
rect 1366 2323 1372 2324
rect 2582 2323 2588 2324
rect 110 2315 116 2316
rect 110 2311 111 2315
rect 115 2311 116 2315
rect 110 2310 116 2311
rect 1326 2315 1332 2316
rect 1326 2311 1327 2315
rect 1331 2311 1332 2315
rect 1326 2310 1332 2311
rect 1366 2311 1372 2312
rect 1366 2307 1367 2311
rect 1371 2307 1372 2311
rect 174 2306 180 2307
rect 174 2302 175 2306
rect 179 2302 180 2306
rect 174 2301 180 2302
rect 278 2306 284 2307
rect 278 2302 279 2306
rect 283 2302 284 2306
rect 278 2301 284 2302
rect 390 2306 396 2307
rect 390 2302 391 2306
rect 395 2302 396 2306
rect 390 2301 396 2302
rect 502 2306 508 2307
rect 502 2302 503 2306
rect 507 2302 508 2306
rect 502 2301 508 2302
rect 614 2306 620 2307
rect 614 2302 615 2306
rect 619 2302 620 2306
rect 614 2301 620 2302
rect 726 2306 732 2307
rect 726 2302 727 2306
rect 731 2302 732 2306
rect 726 2301 732 2302
rect 830 2306 836 2307
rect 830 2302 831 2306
rect 835 2302 836 2306
rect 830 2301 836 2302
rect 926 2306 932 2307
rect 926 2302 927 2306
rect 931 2302 932 2306
rect 926 2301 932 2302
rect 1022 2306 1028 2307
rect 1022 2302 1023 2306
rect 1027 2302 1028 2306
rect 1022 2301 1028 2302
rect 1118 2306 1124 2307
rect 1118 2302 1119 2306
rect 1123 2302 1124 2306
rect 1118 2301 1124 2302
rect 1214 2306 1220 2307
rect 1366 2306 1372 2307
rect 2582 2311 2588 2312
rect 2582 2307 2583 2311
rect 2587 2307 2588 2311
rect 2582 2306 2588 2307
rect 1214 2302 1215 2306
rect 1219 2302 1220 2306
rect 1214 2301 1220 2302
rect 1414 2302 1420 2303
rect 1414 2298 1415 2302
rect 1419 2298 1420 2302
rect 1414 2297 1420 2298
rect 1470 2302 1476 2303
rect 1470 2298 1471 2302
rect 1475 2298 1476 2302
rect 1470 2297 1476 2298
rect 1526 2302 1532 2303
rect 1526 2298 1527 2302
rect 1531 2298 1532 2302
rect 1526 2297 1532 2298
rect 1582 2302 1588 2303
rect 1582 2298 1583 2302
rect 1587 2298 1588 2302
rect 1582 2297 1588 2298
rect 1654 2302 1660 2303
rect 1654 2298 1655 2302
rect 1659 2298 1660 2302
rect 1654 2297 1660 2298
rect 1742 2302 1748 2303
rect 1742 2298 1743 2302
rect 1747 2298 1748 2302
rect 1742 2297 1748 2298
rect 1838 2302 1844 2303
rect 1838 2298 1839 2302
rect 1843 2298 1844 2302
rect 1838 2297 1844 2298
rect 1958 2302 1964 2303
rect 1958 2298 1959 2302
rect 1963 2298 1964 2302
rect 1958 2297 1964 2298
rect 2094 2302 2100 2303
rect 2094 2298 2095 2302
rect 2099 2298 2100 2302
rect 2094 2297 2100 2298
rect 2238 2302 2244 2303
rect 2238 2298 2239 2302
rect 2243 2298 2244 2302
rect 2238 2297 2244 2298
rect 2398 2302 2404 2303
rect 2398 2298 2399 2302
rect 2403 2298 2404 2302
rect 2398 2297 2404 2298
rect 2542 2302 2548 2303
rect 2542 2298 2543 2302
rect 2547 2298 2548 2302
rect 2542 2297 2548 2298
rect 158 2278 164 2279
rect 158 2274 159 2278
rect 163 2274 164 2278
rect 158 2273 164 2274
rect 246 2278 252 2279
rect 246 2274 247 2278
rect 251 2274 252 2278
rect 246 2273 252 2274
rect 374 2278 380 2279
rect 374 2274 375 2278
rect 379 2274 380 2278
rect 374 2273 380 2274
rect 510 2278 516 2279
rect 510 2274 511 2278
rect 515 2274 516 2278
rect 510 2273 516 2274
rect 638 2278 644 2279
rect 638 2274 639 2278
rect 643 2274 644 2278
rect 638 2273 644 2274
rect 766 2278 772 2279
rect 766 2274 767 2278
rect 771 2274 772 2278
rect 766 2273 772 2274
rect 886 2278 892 2279
rect 886 2274 887 2278
rect 891 2274 892 2278
rect 886 2273 892 2274
rect 998 2278 1004 2279
rect 998 2274 999 2278
rect 1003 2274 1004 2278
rect 998 2273 1004 2274
rect 1102 2278 1108 2279
rect 1102 2274 1103 2278
rect 1107 2274 1108 2278
rect 1102 2273 1108 2274
rect 1206 2278 1212 2279
rect 1206 2274 1207 2278
rect 1211 2274 1212 2278
rect 1206 2273 1212 2274
rect 1286 2278 1292 2279
rect 1286 2274 1287 2278
rect 1291 2274 1292 2278
rect 1286 2273 1292 2274
rect 1414 2270 1420 2271
rect 110 2269 116 2270
rect 110 2265 111 2269
rect 115 2265 116 2269
rect 110 2264 116 2265
rect 1326 2269 1332 2270
rect 1326 2265 1327 2269
rect 1331 2265 1332 2269
rect 1414 2266 1415 2270
rect 1419 2266 1420 2270
rect 1414 2265 1420 2266
rect 1494 2270 1500 2271
rect 1494 2266 1495 2270
rect 1499 2266 1500 2270
rect 1494 2265 1500 2266
rect 1614 2270 1620 2271
rect 1614 2266 1615 2270
rect 1619 2266 1620 2270
rect 1614 2265 1620 2266
rect 1734 2270 1740 2271
rect 1734 2266 1735 2270
rect 1739 2266 1740 2270
rect 1734 2265 1740 2266
rect 1854 2270 1860 2271
rect 1854 2266 1855 2270
rect 1859 2266 1860 2270
rect 1854 2265 1860 2266
rect 1966 2270 1972 2271
rect 1966 2266 1967 2270
rect 1971 2266 1972 2270
rect 1966 2265 1972 2266
rect 2070 2270 2076 2271
rect 2070 2266 2071 2270
rect 2075 2266 2076 2270
rect 2070 2265 2076 2266
rect 2166 2270 2172 2271
rect 2166 2266 2167 2270
rect 2171 2266 2172 2270
rect 2166 2265 2172 2266
rect 2254 2270 2260 2271
rect 2254 2266 2255 2270
rect 2259 2266 2260 2270
rect 2254 2265 2260 2266
rect 2334 2270 2340 2271
rect 2334 2266 2335 2270
rect 2339 2266 2340 2270
rect 2334 2265 2340 2266
rect 2406 2270 2412 2271
rect 2406 2266 2407 2270
rect 2411 2266 2412 2270
rect 2406 2265 2412 2266
rect 2486 2270 2492 2271
rect 2486 2266 2487 2270
rect 2491 2266 2492 2270
rect 2486 2265 2492 2266
rect 2542 2270 2548 2271
rect 2542 2266 2543 2270
rect 2547 2266 2548 2270
rect 2542 2265 2548 2266
rect 1326 2264 1332 2265
rect 1366 2261 1372 2262
rect 1366 2257 1367 2261
rect 1371 2257 1372 2261
rect 1366 2256 1372 2257
rect 2582 2261 2588 2262
rect 2582 2257 2583 2261
rect 2587 2257 2588 2261
rect 2582 2256 2588 2257
rect 110 2252 116 2253
rect 1326 2252 1332 2253
rect 110 2248 111 2252
rect 115 2248 116 2252
rect 110 2247 116 2248
rect 142 2251 148 2252
rect 142 2247 143 2251
rect 147 2247 148 2251
rect 142 2246 148 2247
rect 230 2251 236 2252
rect 230 2247 231 2251
rect 235 2247 236 2251
rect 230 2246 236 2247
rect 358 2251 364 2252
rect 358 2247 359 2251
rect 363 2247 364 2251
rect 358 2246 364 2247
rect 494 2251 500 2252
rect 494 2247 495 2251
rect 499 2247 500 2251
rect 494 2246 500 2247
rect 622 2251 628 2252
rect 622 2247 623 2251
rect 627 2247 628 2251
rect 622 2246 628 2247
rect 750 2251 756 2252
rect 750 2247 751 2251
rect 755 2247 756 2251
rect 750 2246 756 2247
rect 870 2251 876 2252
rect 870 2247 871 2251
rect 875 2247 876 2251
rect 870 2246 876 2247
rect 982 2251 988 2252
rect 982 2247 983 2251
rect 987 2247 988 2251
rect 982 2246 988 2247
rect 1086 2251 1092 2252
rect 1086 2247 1087 2251
rect 1091 2247 1092 2251
rect 1086 2246 1092 2247
rect 1190 2251 1196 2252
rect 1190 2247 1191 2251
rect 1195 2247 1196 2251
rect 1190 2246 1196 2247
rect 1270 2251 1276 2252
rect 1270 2247 1271 2251
rect 1275 2247 1276 2251
rect 1326 2248 1327 2252
rect 1331 2248 1332 2252
rect 1326 2247 1332 2248
rect 1270 2246 1276 2247
rect 1366 2244 1372 2245
rect 2582 2244 2588 2245
rect 1366 2240 1367 2244
rect 1371 2240 1372 2244
rect 1366 2239 1372 2240
rect 1398 2243 1404 2244
rect 1398 2239 1399 2243
rect 1403 2239 1404 2243
rect 1398 2238 1404 2239
rect 1478 2243 1484 2244
rect 1478 2239 1479 2243
rect 1483 2239 1484 2243
rect 1478 2238 1484 2239
rect 1598 2243 1604 2244
rect 1598 2239 1599 2243
rect 1603 2239 1604 2243
rect 1598 2238 1604 2239
rect 1718 2243 1724 2244
rect 1718 2239 1719 2243
rect 1723 2239 1724 2243
rect 1718 2238 1724 2239
rect 1838 2243 1844 2244
rect 1838 2239 1839 2243
rect 1843 2239 1844 2243
rect 1838 2238 1844 2239
rect 1950 2243 1956 2244
rect 1950 2239 1951 2243
rect 1955 2239 1956 2243
rect 1950 2238 1956 2239
rect 2054 2243 2060 2244
rect 2054 2239 2055 2243
rect 2059 2239 2060 2243
rect 2054 2238 2060 2239
rect 2150 2243 2156 2244
rect 2150 2239 2151 2243
rect 2155 2239 2156 2243
rect 2150 2238 2156 2239
rect 2238 2243 2244 2244
rect 2238 2239 2239 2243
rect 2243 2239 2244 2243
rect 2238 2238 2244 2239
rect 2318 2243 2324 2244
rect 2318 2239 2319 2243
rect 2323 2239 2324 2243
rect 2318 2238 2324 2239
rect 2390 2243 2396 2244
rect 2390 2239 2391 2243
rect 2395 2239 2396 2243
rect 2390 2238 2396 2239
rect 2470 2243 2476 2244
rect 2470 2239 2471 2243
rect 2475 2239 2476 2243
rect 2470 2238 2476 2239
rect 2526 2243 2532 2244
rect 2526 2239 2527 2243
rect 2531 2239 2532 2243
rect 2582 2240 2583 2244
rect 2587 2240 2588 2244
rect 2582 2239 2588 2240
rect 2526 2238 2532 2239
rect 142 2209 148 2210
rect 110 2208 116 2209
rect 110 2204 111 2208
rect 115 2204 116 2208
rect 142 2205 143 2209
rect 147 2205 148 2209
rect 142 2204 148 2205
rect 230 2209 236 2210
rect 230 2205 231 2209
rect 235 2205 236 2209
rect 230 2204 236 2205
rect 358 2209 364 2210
rect 358 2205 359 2209
rect 363 2205 364 2209
rect 358 2204 364 2205
rect 494 2209 500 2210
rect 494 2205 495 2209
rect 499 2205 500 2209
rect 494 2204 500 2205
rect 622 2209 628 2210
rect 622 2205 623 2209
rect 627 2205 628 2209
rect 622 2204 628 2205
rect 750 2209 756 2210
rect 750 2205 751 2209
rect 755 2205 756 2209
rect 750 2204 756 2205
rect 870 2209 876 2210
rect 870 2205 871 2209
rect 875 2205 876 2209
rect 870 2204 876 2205
rect 982 2209 988 2210
rect 982 2205 983 2209
rect 987 2205 988 2209
rect 982 2204 988 2205
rect 1086 2209 1092 2210
rect 1086 2205 1087 2209
rect 1091 2205 1092 2209
rect 1086 2204 1092 2205
rect 1190 2209 1196 2210
rect 1190 2205 1191 2209
rect 1195 2205 1196 2209
rect 1190 2204 1196 2205
rect 1270 2209 1276 2210
rect 1270 2205 1271 2209
rect 1275 2205 1276 2209
rect 1270 2204 1276 2205
rect 1326 2208 1332 2209
rect 1326 2204 1327 2208
rect 1331 2204 1332 2208
rect 110 2203 116 2204
rect 1326 2203 1332 2204
rect 1454 2197 1460 2198
rect 1366 2196 1372 2197
rect 1366 2192 1367 2196
rect 1371 2192 1372 2196
rect 1454 2193 1455 2197
rect 1459 2193 1460 2197
rect 1454 2192 1460 2193
rect 1534 2197 1540 2198
rect 1534 2193 1535 2197
rect 1539 2193 1540 2197
rect 1534 2192 1540 2193
rect 1630 2197 1636 2198
rect 1630 2193 1631 2197
rect 1635 2193 1636 2197
rect 1630 2192 1636 2193
rect 1742 2197 1748 2198
rect 1742 2193 1743 2197
rect 1747 2193 1748 2197
rect 1742 2192 1748 2193
rect 1862 2197 1868 2198
rect 1862 2193 1863 2197
rect 1867 2193 1868 2197
rect 1862 2192 1868 2193
rect 1982 2197 1988 2198
rect 1982 2193 1983 2197
rect 1987 2193 1988 2197
rect 1982 2192 1988 2193
rect 2094 2197 2100 2198
rect 2094 2193 2095 2197
rect 2099 2193 2100 2197
rect 2094 2192 2100 2193
rect 2206 2197 2212 2198
rect 2206 2193 2207 2197
rect 2211 2193 2212 2197
rect 2206 2192 2212 2193
rect 2310 2197 2316 2198
rect 2310 2193 2311 2197
rect 2315 2193 2316 2197
rect 2310 2192 2316 2193
rect 2422 2197 2428 2198
rect 2422 2193 2423 2197
rect 2427 2193 2428 2197
rect 2422 2192 2428 2193
rect 2526 2197 2532 2198
rect 2526 2193 2527 2197
rect 2531 2193 2532 2197
rect 2526 2192 2532 2193
rect 2582 2196 2588 2197
rect 2582 2192 2583 2196
rect 2587 2192 2588 2196
rect 110 2191 116 2192
rect 110 2187 111 2191
rect 115 2187 116 2191
rect 110 2186 116 2187
rect 1326 2191 1332 2192
rect 1366 2191 1372 2192
rect 2582 2191 2588 2192
rect 1326 2187 1327 2191
rect 1331 2187 1332 2191
rect 1326 2186 1332 2187
rect 158 2182 164 2183
rect 158 2178 159 2182
rect 163 2178 164 2182
rect 158 2177 164 2178
rect 246 2182 252 2183
rect 246 2178 247 2182
rect 251 2178 252 2182
rect 246 2177 252 2178
rect 374 2182 380 2183
rect 374 2178 375 2182
rect 379 2178 380 2182
rect 374 2177 380 2178
rect 510 2182 516 2183
rect 510 2178 511 2182
rect 515 2178 516 2182
rect 510 2177 516 2178
rect 638 2182 644 2183
rect 638 2178 639 2182
rect 643 2178 644 2182
rect 638 2177 644 2178
rect 766 2182 772 2183
rect 766 2178 767 2182
rect 771 2178 772 2182
rect 766 2177 772 2178
rect 886 2182 892 2183
rect 886 2178 887 2182
rect 891 2178 892 2182
rect 886 2177 892 2178
rect 998 2182 1004 2183
rect 998 2178 999 2182
rect 1003 2178 1004 2182
rect 998 2177 1004 2178
rect 1102 2182 1108 2183
rect 1102 2178 1103 2182
rect 1107 2178 1108 2182
rect 1102 2177 1108 2178
rect 1206 2182 1212 2183
rect 1206 2178 1207 2182
rect 1211 2178 1212 2182
rect 1206 2177 1212 2178
rect 1286 2182 1292 2183
rect 1286 2178 1287 2182
rect 1291 2178 1292 2182
rect 1286 2177 1292 2178
rect 1366 2179 1372 2180
rect 1366 2175 1367 2179
rect 1371 2175 1372 2179
rect 1366 2174 1372 2175
rect 2582 2179 2588 2180
rect 2582 2175 2583 2179
rect 2587 2175 2588 2179
rect 2582 2174 2588 2175
rect 1470 2170 1476 2171
rect 1470 2166 1471 2170
rect 1475 2166 1476 2170
rect 1470 2165 1476 2166
rect 1550 2170 1556 2171
rect 1550 2166 1551 2170
rect 1555 2166 1556 2170
rect 1550 2165 1556 2166
rect 1646 2170 1652 2171
rect 1646 2166 1647 2170
rect 1651 2166 1652 2170
rect 1646 2165 1652 2166
rect 1758 2170 1764 2171
rect 1758 2166 1759 2170
rect 1763 2166 1764 2170
rect 1758 2165 1764 2166
rect 1878 2170 1884 2171
rect 1878 2166 1879 2170
rect 1883 2166 1884 2170
rect 1878 2165 1884 2166
rect 1998 2170 2004 2171
rect 1998 2166 1999 2170
rect 2003 2166 2004 2170
rect 1998 2165 2004 2166
rect 2110 2170 2116 2171
rect 2110 2166 2111 2170
rect 2115 2166 2116 2170
rect 2110 2165 2116 2166
rect 2222 2170 2228 2171
rect 2222 2166 2223 2170
rect 2227 2166 2228 2170
rect 2222 2165 2228 2166
rect 2326 2170 2332 2171
rect 2326 2166 2327 2170
rect 2331 2166 2332 2170
rect 2326 2165 2332 2166
rect 2438 2170 2444 2171
rect 2438 2166 2439 2170
rect 2443 2166 2444 2170
rect 2438 2165 2444 2166
rect 2542 2170 2548 2171
rect 2542 2166 2543 2170
rect 2547 2166 2548 2170
rect 2542 2165 2548 2166
rect 158 2154 164 2155
rect 158 2150 159 2154
rect 163 2150 164 2154
rect 158 2149 164 2150
rect 214 2154 220 2155
rect 214 2150 215 2154
rect 219 2150 220 2154
rect 214 2149 220 2150
rect 310 2154 316 2155
rect 310 2150 311 2154
rect 315 2150 316 2154
rect 310 2149 316 2150
rect 422 2154 428 2155
rect 422 2150 423 2154
rect 427 2150 428 2154
rect 422 2149 428 2150
rect 542 2154 548 2155
rect 542 2150 543 2154
rect 547 2150 548 2154
rect 542 2149 548 2150
rect 662 2154 668 2155
rect 662 2150 663 2154
rect 667 2150 668 2154
rect 662 2149 668 2150
rect 774 2154 780 2155
rect 774 2150 775 2154
rect 779 2150 780 2154
rect 774 2149 780 2150
rect 878 2154 884 2155
rect 878 2150 879 2154
rect 883 2150 884 2154
rect 878 2149 884 2150
rect 974 2154 980 2155
rect 974 2150 975 2154
rect 979 2150 980 2154
rect 974 2149 980 2150
rect 1070 2154 1076 2155
rect 1070 2150 1071 2154
rect 1075 2150 1076 2154
rect 1070 2149 1076 2150
rect 1166 2154 1172 2155
rect 1166 2150 1167 2154
rect 1171 2150 1172 2154
rect 1166 2149 1172 2150
rect 1270 2154 1276 2155
rect 1270 2150 1271 2154
rect 1275 2150 1276 2154
rect 1270 2149 1276 2150
rect 1534 2146 1540 2147
rect 110 2145 116 2146
rect 110 2141 111 2145
rect 115 2141 116 2145
rect 110 2140 116 2141
rect 1326 2145 1332 2146
rect 1326 2141 1327 2145
rect 1331 2141 1332 2145
rect 1534 2142 1535 2146
rect 1539 2142 1540 2146
rect 1534 2141 1540 2142
rect 1630 2146 1636 2147
rect 1630 2142 1631 2146
rect 1635 2142 1636 2146
rect 1630 2141 1636 2142
rect 1734 2146 1740 2147
rect 1734 2142 1735 2146
rect 1739 2142 1740 2146
rect 1734 2141 1740 2142
rect 1838 2146 1844 2147
rect 1838 2142 1839 2146
rect 1843 2142 1844 2146
rect 1838 2141 1844 2142
rect 1950 2146 1956 2147
rect 1950 2142 1951 2146
rect 1955 2142 1956 2146
rect 1950 2141 1956 2142
rect 2054 2146 2060 2147
rect 2054 2142 2055 2146
rect 2059 2142 2060 2146
rect 2054 2141 2060 2142
rect 2158 2146 2164 2147
rect 2158 2142 2159 2146
rect 2163 2142 2164 2146
rect 2158 2141 2164 2142
rect 2262 2146 2268 2147
rect 2262 2142 2263 2146
rect 2267 2142 2268 2146
rect 2262 2141 2268 2142
rect 2358 2146 2364 2147
rect 2358 2142 2359 2146
rect 2363 2142 2364 2146
rect 2358 2141 2364 2142
rect 2462 2146 2468 2147
rect 2462 2142 2463 2146
rect 2467 2142 2468 2146
rect 2462 2141 2468 2142
rect 2542 2146 2548 2147
rect 2542 2142 2543 2146
rect 2547 2142 2548 2146
rect 2542 2141 2548 2142
rect 1326 2140 1332 2141
rect 1366 2137 1372 2138
rect 1366 2133 1367 2137
rect 1371 2133 1372 2137
rect 1366 2132 1372 2133
rect 2582 2137 2588 2138
rect 2582 2133 2583 2137
rect 2587 2133 2588 2137
rect 2582 2132 2588 2133
rect 110 2128 116 2129
rect 1326 2128 1332 2129
rect 110 2124 111 2128
rect 115 2124 116 2128
rect 110 2123 116 2124
rect 142 2127 148 2128
rect 142 2123 143 2127
rect 147 2123 148 2127
rect 142 2122 148 2123
rect 198 2127 204 2128
rect 198 2123 199 2127
rect 203 2123 204 2127
rect 198 2122 204 2123
rect 294 2127 300 2128
rect 294 2123 295 2127
rect 299 2123 300 2127
rect 294 2122 300 2123
rect 406 2127 412 2128
rect 406 2123 407 2127
rect 411 2123 412 2127
rect 406 2122 412 2123
rect 526 2127 532 2128
rect 526 2123 527 2127
rect 531 2123 532 2127
rect 526 2122 532 2123
rect 646 2127 652 2128
rect 646 2123 647 2127
rect 651 2123 652 2127
rect 646 2122 652 2123
rect 758 2127 764 2128
rect 758 2123 759 2127
rect 763 2123 764 2127
rect 758 2122 764 2123
rect 862 2127 868 2128
rect 862 2123 863 2127
rect 867 2123 868 2127
rect 862 2122 868 2123
rect 958 2127 964 2128
rect 958 2123 959 2127
rect 963 2123 964 2127
rect 958 2122 964 2123
rect 1054 2127 1060 2128
rect 1054 2123 1055 2127
rect 1059 2123 1060 2127
rect 1054 2122 1060 2123
rect 1150 2127 1156 2128
rect 1150 2123 1151 2127
rect 1155 2123 1156 2127
rect 1150 2122 1156 2123
rect 1254 2127 1260 2128
rect 1254 2123 1255 2127
rect 1259 2123 1260 2127
rect 1326 2124 1327 2128
rect 1331 2124 1332 2128
rect 1326 2123 1332 2124
rect 1254 2122 1260 2123
rect 1366 2120 1372 2121
rect 2582 2120 2588 2121
rect 1366 2116 1367 2120
rect 1371 2116 1372 2120
rect 1366 2115 1372 2116
rect 1518 2119 1524 2120
rect 1518 2115 1519 2119
rect 1523 2115 1524 2119
rect 1518 2114 1524 2115
rect 1614 2119 1620 2120
rect 1614 2115 1615 2119
rect 1619 2115 1620 2119
rect 1614 2114 1620 2115
rect 1718 2119 1724 2120
rect 1718 2115 1719 2119
rect 1723 2115 1724 2119
rect 1718 2114 1724 2115
rect 1822 2119 1828 2120
rect 1822 2115 1823 2119
rect 1827 2115 1828 2119
rect 1822 2114 1828 2115
rect 1934 2119 1940 2120
rect 1934 2115 1935 2119
rect 1939 2115 1940 2119
rect 1934 2114 1940 2115
rect 2038 2119 2044 2120
rect 2038 2115 2039 2119
rect 2043 2115 2044 2119
rect 2038 2114 2044 2115
rect 2142 2119 2148 2120
rect 2142 2115 2143 2119
rect 2147 2115 2148 2119
rect 2142 2114 2148 2115
rect 2246 2119 2252 2120
rect 2246 2115 2247 2119
rect 2251 2115 2252 2119
rect 2246 2114 2252 2115
rect 2342 2119 2348 2120
rect 2342 2115 2343 2119
rect 2347 2115 2348 2119
rect 2342 2114 2348 2115
rect 2446 2119 2452 2120
rect 2446 2115 2447 2119
rect 2451 2115 2452 2119
rect 2446 2114 2452 2115
rect 2526 2119 2532 2120
rect 2526 2115 2527 2119
rect 2531 2115 2532 2119
rect 2582 2116 2583 2120
rect 2587 2116 2588 2120
rect 2582 2115 2588 2116
rect 2526 2114 2532 2115
rect 262 2085 268 2086
rect 110 2084 116 2085
rect 110 2080 111 2084
rect 115 2080 116 2084
rect 262 2081 263 2085
rect 267 2081 268 2085
rect 262 2080 268 2081
rect 326 2085 332 2086
rect 326 2081 327 2085
rect 331 2081 332 2085
rect 326 2080 332 2081
rect 398 2085 404 2086
rect 398 2081 399 2085
rect 403 2081 404 2085
rect 398 2080 404 2081
rect 478 2085 484 2086
rect 478 2081 479 2085
rect 483 2081 484 2085
rect 478 2080 484 2081
rect 566 2085 572 2086
rect 566 2081 567 2085
rect 571 2081 572 2085
rect 566 2080 572 2081
rect 654 2085 660 2086
rect 654 2081 655 2085
rect 659 2081 660 2085
rect 654 2080 660 2081
rect 734 2085 740 2086
rect 734 2081 735 2085
rect 739 2081 740 2085
rect 734 2080 740 2081
rect 814 2085 820 2086
rect 814 2081 815 2085
rect 819 2081 820 2085
rect 814 2080 820 2081
rect 886 2085 892 2086
rect 886 2081 887 2085
rect 891 2081 892 2085
rect 886 2080 892 2081
rect 966 2085 972 2086
rect 966 2081 967 2085
rect 971 2081 972 2085
rect 966 2080 972 2081
rect 1046 2085 1052 2086
rect 1046 2081 1047 2085
rect 1051 2081 1052 2085
rect 1046 2080 1052 2081
rect 1126 2085 1132 2086
rect 1430 2085 1436 2086
rect 1126 2081 1127 2085
rect 1131 2081 1132 2085
rect 1126 2080 1132 2081
rect 1326 2084 1332 2085
rect 1326 2080 1327 2084
rect 1331 2080 1332 2084
rect 110 2079 116 2080
rect 1326 2079 1332 2080
rect 1366 2084 1372 2085
rect 1366 2080 1367 2084
rect 1371 2080 1372 2084
rect 1430 2081 1431 2085
rect 1435 2081 1436 2085
rect 1430 2080 1436 2081
rect 1534 2085 1540 2086
rect 1534 2081 1535 2085
rect 1539 2081 1540 2085
rect 1534 2080 1540 2081
rect 1646 2085 1652 2086
rect 1646 2081 1647 2085
rect 1651 2081 1652 2085
rect 1646 2080 1652 2081
rect 1758 2085 1764 2086
rect 1758 2081 1759 2085
rect 1763 2081 1764 2085
rect 1758 2080 1764 2081
rect 1862 2085 1868 2086
rect 1862 2081 1863 2085
rect 1867 2081 1868 2085
rect 1862 2080 1868 2081
rect 1966 2085 1972 2086
rect 1966 2081 1967 2085
rect 1971 2081 1972 2085
rect 1966 2080 1972 2081
rect 2070 2085 2076 2086
rect 2070 2081 2071 2085
rect 2075 2081 2076 2085
rect 2070 2080 2076 2081
rect 2174 2085 2180 2086
rect 2174 2081 2175 2085
rect 2179 2081 2180 2085
rect 2174 2080 2180 2081
rect 2270 2085 2276 2086
rect 2270 2081 2271 2085
rect 2275 2081 2276 2085
rect 2270 2080 2276 2081
rect 2358 2085 2364 2086
rect 2358 2081 2359 2085
rect 2363 2081 2364 2085
rect 2358 2080 2364 2081
rect 2454 2085 2460 2086
rect 2454 2081 2455 2085
rect 2459 2081 2460 2085
rect 2454 2080 2460 2081
rect 2526 2085 2532 2086
rect 2526 2081 2527 2085
rect 2531 2081 2532 2085
rect 2526 2080 2532 2081
rect 2582 2084 2588 2085
rect 2582 2080 2583 2084
rect 2587 2080 2588 2084
rect 1366 2079 1372 2080
rect 2582 2079 2588 2080
rect 110 2067 116 2068
rect 110 2063 111 2067
rect 115 2063 116 2067
rect 110 2062 116 2063
rect 1326 2067 1332 2068
rect 1326 2063 1327 2067
rect 1331 2063 1332 2067
rect 1326 2062 1332 2063
rect 1366 2067 1372 2068
rect 1366 2063 1367 2067
rect 1371 2063 1372 2067
rect 1366 2062 1372 2063
rect 2582 2067 2588 2068
rect 2582 2063 2583 2067
rect 2587 2063 2588 2067
rect 2582 2062 2588 2063
rect 278 2058 284 2059
rect 278 2054 279 2058
rect 283 2054 284 2058
rect 278 2053 284 2054
rect 342 2058 348 2059
rect 342 2054 343 2058
rect 347 2054 348 2058
rect 342 2053 348 2054
rect 414 2058 420 2059
rect 414 2054 415 2058
rect 419 2054 420 2058
rect 414 2053 420 2054
rect 494 2058 500 2059
rect 494 2054 495 2058
rect 499 2054 500 2058
rect 494 2053 500 2054
rect 582 2058 588 2059
rect 582 2054 583 2058
rect 587 2054 588 2058
rect 582 2053 588 2054
rect 670 2058 676 2059
rect 670 2054 671 2058
rect 675 2054 676 2058
rect 670 2053 676 2054
rect 750 2058 756 2059
rect 750 2054 751 2058
rect 755 2054 756 2058
rect 750 2053 756 2054
rect 830 2058 836 2059
rect 830 2054 831 2058
rect 835 2054 836 2058
rect 830 2053 836 2054
rect 902 2058 908 2059
rect 902 2054 903 2058
rect 907 2054 908 2058
rect 902 2053 908 2054
rect 982 2058 988 2059
rect 982 2054 983 2058
rect 987 2054 988 2058
rect 982 2053 988 2054
rect 1062 2058 1068 2059
rect 1062 2054 1063 2058
rect 1067 2054 1068 2058
rect 1062 2053 1068 2054
rect 1142 2058 1148 2059
rect 1142 2054 1143 2058
rect 1147 2054 1148 2058
rect 1142 2053 1148 2054
rect 1446 2058 1452 2059
rect 1446 2054 1447 2058
rect 1451 2054 1452 2058
rect 1446 2053 1452 2054
rect 1550 2058 1556 2059
rect 1550 2054 1551 2058
rect 1555 2054 1556 2058
rect 1550 2053 1556 2054
rect 1662 2058 1668 2059
rect 1662 2054 1663 2058
rect 1667 2054 1668 2058
rect 1662 2053 1668 2054
rect 1774 2058 1780 2059
rect 1774 2054 1775 2058
rect 1779 2054 1780 2058
rect 1774 2053 1780 2054
rect 1878 2058 1884 2059
rect 1878 2054 1879 2058
rect 1883 2054 1884 2058
rect 1878 2053 1884 2054
rect 1982 2058 1988 2059
rect 1982 2054 1983 2058
rect 1987 2054 1988 2058
rect 1982 2053 1988 2054
rect 2086 2058 2092 2059
rect 2086 2054 2087 2058
rect 2091 2054 2092 2058
rect 2086 2053 2092 2054
rect 2190 2058 2196 2059
rect 2190 2054 2191 2058
rect 2195 2054 2196 2058
rect 2190 2053 2196 2054
rect 2286 2058 2292 2059
rect 2286 2054 2287 2058
rect 2291 2054 2292 2058
rect 2286 2053 2292 2054
rect 2374 2058 2380 2059
rect 2374 2054 2375 2058
rect 2379 2054 2380 2058
rect 2374 2053 2380 2054
rect 2470 2058 2476 2059
rect 2470 2054 2471 2058
rect 2475 2054 2476 2058
rect 2470 2053 2476 2054
rect 2542 2058 2548 2059
rect 2542 2054 2543 2058
rect 2547 2054 2548 2058
rect 2542 2053 2548 2054
rect 1414 2034 1420 2035
rect 1414 2030 1415 2034
rect 1419 2030 1420 2034
rect 1414 2029 1420 2030
rect 1502 2034 1508 2035
rect 1502 2030 1503 2034
rect 1507 2030 1508 2034
rect 1502 2029 1508 2030
rect 1606 2034 1612 2035
rect 1606 2030 1607 2034
rect 1611 2030 1612 2034
rect 1606 2029 1612 2030
rect 1710 2034 1716 2035
rect 1710 2030 1711 2034
rect 1715 2030 1716 2034
rect 1710 2029 1716 2030
rect 1806 2034 1812 2035
rect 1806 2030 1807 2034
rect 1811 2030 1812 2034
rect 1806 2029 1812 2030
rect 1902 2034 1908 2035
rect 1902 2030 1903 2034
rect 1907 2030 1908 2034
rect 1902 2029 1908 2030
rect 2006 2034 2012 2035
rect 2006 2030 2007 2034
rect 2011 2030 2012 2034
rect 2006 2029 2012 2030
rect 2110 2034 2116 2035
rect 2110 2030 2111 2034
rect 2115 2030 2116 2034
rect 2110 2029 2116 2030
rect 2214 2034 2220 2035
rect 2214 2030 2215 2034
rect 2219 2030 2220 2034
rect 2214 2029 2220 2030
rect 2326 2034 2332 2035
rect 2326 2030 2327 2034
rect 2331 2030 2332 2034
rect 2326 2029 2332 2030
rect 2446 2034 2452 2035
rect 2446 2030 2447 2034
rect 2451 2030 2452 2034
rect 2446 2029 2452 2030
rect 2542 2034 2548 2035
rect 2542 2030 2543 2034
rect 2547 2030 2548 2034
rect 2542 2029 2548 2030
rect 414 2026 420 2027
rect 414 2022 415 2026
rect 419 2022 420 2026
rect 414 2021 420 2022
rect 470 2026 476 2027
rect 470 2022 471 2026
rect 475 2022 476 2026
rect 470 2021 476 2022
rect 526 2026 532 2027
rect 526 2022 527 2026
rect 531 2022 532 2026
rect 526 2021 532 2022
rect 582 2026 588 2027
rect 582 2022 583 2026
rect 587 2022 588 2026
rect 582 2021 588 2022
rect 638 2026 644 2027
rect 638 2022 639 2026
rect 643 2022 644 2026
rect 638 2021 644 2022
rect 694 2026 700 2027
rect 694 2022 695 2026
rect 699 2022 700 2026
rect 694 2021 700 2022
rect 750 2026 756 2027
rect 750 2022 751 2026
rect 755 2022 756 2026
rect 750 2021 756 2022
rect 806 2026 812 2027
rect 806 2022 807 2026
rect 811 2022 812 2026
rect 806 2021 812 2022
rect 862 2026 868 2027
rect 862 2022 863 2026
rect 867 2022 868 2026
rect 862 2021 868 2022
rect 918 2026 924 2027
rect 918 2022 919 2026
rect 923 2022 924 2026
rect 918 2021 924 2022
rect 974 2026 980 2027
rect 974 2022 975 2026
rect 979 2022 980 2026
rect 974 2021 980 2022
rect 1030 2026 1036 2027
rect 1030 2022 1031 2026
rect 1035 2022 1036 2026
rect 1030 2021 1036 2022
rect 1366 2025 1372 2026
rect 1366 2021 1367 2025
rect 1371 2021 1372 2025
rect 1366 2020 1372 2021
rect 2582 2025 2588 2026
rect 2582 2021 2583 2025
rect 2587 2021 2588 2025
rect 2582 2020 2588 2021
rect 110 2017 116 2018
rect 110 2013 111 2017
rect 115 2013 116 2017
rect 110 2012 116 2013
rect 1326 2017 1332 2018
rect 1326 2013 1327 2017
rect 1331 2013 1332 2017
rect 1326 2012 1332 2013
rect 1366 2008 1372 2009
rect 2582 2008 2588 2009
rect 1366 2004 1367 2008
rect 1371 2004 1372 2008
rect 1366 2003 1372 2004
rect 1398 2007 1404 2008
rect 1398 2003 1399 2007
rect 1403 2003 1404 2007
rect 1398 2002 1404 2003
rect 1486 2007 1492 2008
rect 1486 2003 1487 2007
rect 1491 2003 1492 2007
rect 1486 2002 1492 2003
rect 1590 2007 1596 2008
rect 1590 2003 1591 2007
rect 1595 2003 1596 2007
rect 1590 2002 1596 2003
rect 1694 2007 1700 2008
rect 1694 2003 1695 2007
rect 1699 2003 1700 2007
rect 1694 2002 1700 2003
rect 1790 2007 1796 2008
rect 1790 2003 1791 2007
rect 1795 2003 1796 2007
rect 1790 2002 1796 2003
rect 1886 2007 1892 2008
rect 1886 2003 1887 2007
rect 1891 2003 1892 2007
rect 1886 2002 1892 2003
rect 1990 2007 1996 2008
rect 1990 2003 1991 2007
rect 1995 2003 1996 2007
rect 1990 2002 1996 2003
rect 2094 2007 2100 2008
rect 2094 2003 2095 2007
rect 2099 2003 2100 2007
rect 2094 2002 2100 2003
rect 2198 2007 2204 2008
rect 2198 2003 2199 2007
rect 2203 2003 2204 2007
rect 2198 2002 2204 2003
rect 2310 2007 2316 2008
rect 2310 2003 2311 2007
rect 2315 2003 2316 2007
rect 2310 2002 2316 2003
rect 2430 2007 2436 2008
rect 2430 2003 2431 2007
rect 2435 2003 2436 2007
rect 2430 2002 2436 2003
rect 2526 2007 2532 2008
rect 2526 2003 2527 2007
rect 2531 2003 2532 2007
rect 2582 2004 2583 2008
rect 2587 2004 2588 2008
rect 2582 2003 2588 2004
rect 2526 2002 2532 2003
rect 110 2000 116 2001
rect 1326 2000 1332 2001
rect 110 1996 111 2000
rect 115 1996 116 2000
rect 110 1995 116 1996
rect 398 1999 404 2000
rect 398 1995 399 1999
rect 403 1995 404 1999
rect 398 1994 404 1995
rect 454 1999 460 2000
rect 454 1995 455 1999
rect 459 1995 460 1999
rect 454 1994 460 1995
rect 510 1999 516 2000
rect 510 1995 511 1999
rect 515 1995 516 1999
rect 510 1994 516 1995
rect 566 1999 572 2000
rect 566 1995 567 1999
rect 571 1995 572 1999
rect 566 1994 572 1995
rect 622 1999 628 2000
rect 622 1995 623 1999
rect 627 1995 628 1999
rect 622 1994 628 1995
rect 678 1999 684 2000
rect 678 1995 679 1999
rect 683 1995 684 1999
rect 678 1994 684 1995
rect 734 1999 740 2000
rect 734 1995 735 1999
rect 739 1995 740 1999
rect 734 1994 740 1995
rect 790 1999 796 2000
rect 790 1995 791 1999
rect 795 1995 796 1999
rect 790 1994 796 1995
rect 846 1999 852 2000
rect 846 1995 847 1999
rect 851 1995 852 1999
rect 846 1994 852 1995
rect 902 1999 908 2000
rect 902 1995 903 1999
rect 907 1995 908 1999
rect 902 1994 908 1995
rect 958 1999 964 2000
rect 958 1995 959 1999
rect 963 1995 964 1999
rect 958 1994 964 1995
rect 1014 1999 1020 2000
rect 1014 1995 1015 1999
rect 1019 1995 1020 1999
rect 1326 1996 1327 2000
rect 1331 1996 1332 2000
rect 1326 1995 1332 1996
rect 1014 1994 1020 1995
rect 1398 1973 1404 1974
rect 1366 1972 1372 1973
rect 1366 1968 1367 1972
rect 1371 1968 1372 1972
rect 1398 1969 1399 1973
rect 1403 1969 1404 1973
rect 1398 1968 1404 1969
rect 1478 1973 1484 1974
rect 1478 1969 1479 1973
rect 1483 1969 1484 1973
rect 1478 1968 1484 1969
rect 1582 1973 1588 1974
rect 1582 1969 1583 1973
rect 1587 1969 1588 1973
rect 1582 1968 1588 1969
rect 1678 1973 1684 1974
rect 1678 1969 1679 1973
rect 1683 1969 1684 1973
rect 1678 1968 1684 1969
rect 1766 1973 1772 1974
rect 1766 1969 1767 1973
rect 1771 1969 1772 1973
rect 1766 1968 1772 1969
rect 1846 1973 1852 1974
rect 1846 1969 1847 1973
rect 1851 1969 1852 1973
rect 1846 1968 1852 1969
rect 1926 1973 1932 1974
rect 1926 1969 1927 1973
rect 1931 1969 1932 1973
rect 1926 1968 1932 1969
rect 2006 1973 2012 1974
rect 2006 1969 2007 1973
rect 2011 1969 2012 1973
rect 2006 1968 2012 1969
rect 2086 1973 2092 1974
rect 2086 1969 2087 1973
rect 2091 1969 2092 1973
rect 2086 1968 2092 1969
rect 2582 1972 2588 1973
rect 2582 1968 2583 1972
rect 2587 1968 2588 1972
rect 1366 1967 1372 1968
rect 2582 1967 2588 1968
rect 334 1961 340 1962
rect 110 1960 116 1961
rect 110 1956 111 1960
rect 115 1956 116 1960
rect 334 1957 335 1961
rect 339 1957 340 1961
rect 334 1956 340 1957
rect 390 1961 396 1962
rect 390 1957 391 1961
rect 395 1957 396 1961
rect 390 1956 396 1957
rect 446 1961 452 1962
rect 446 1957 447 1961
rect 451 1957 452 1961
rect 446 1956 452 1957
rect 502 1961 508 1962
rect 502 1957 503 1961
rect 507 1957 508 1961
rect 502 1956 508 1957
rect 566 1961 572 1962
rect 566 1957 567 1961
rect 571 1957 572 1961
rect 566 1956 572 1957
rect 646 1961 652 1962
rect 646 1957 647 1961
rect 651 1957 652 1961
rect 646 1956 652 1957
rect 742 1961 748 1962
rect 742 1957 743 1961
rect 747 1957 748 1961
rect 742 1956 748 1957
rect 862 1961 868 1962
rect 862 1957 863 1961
rect 867 1957 868 1961
rect 862 1956 868 1957
rect 998 1961 1004 1962
rect 998 1957 999 1961
rect 1003 1957 1004 1961
rect 998 1956 1004 1957
rect 1142 1961 1148 1962
rect 1142 1957 1143 1961
rect 1147 1957 1148 1961
rect 1142 1956 1148 1957
rect 1270 1961 1276 1962
rect 1270 1957 1271 1961
rect 1275 1957 1276 1961
rect 1270 1956 1276 1957
rect 1326 1960 1332 1961
rect 1326 1956 1327 1960
rect 1331 1956 1332 1960
rect 110 1955 116 1956
rect 1326 1955 1332 1956
rect 1366 1955 1372 1956
rect 1366 1951 1367 1955
rect 1371 1951 1372 1955
rect 1366 1950 1372 1951
rect 2582 1955 2588 1956
rect 2582 1951 2583 1955
rect 2587 1951 2588 1955
rect 2582 1950 2588 1951
rect 1414 1946 1420 1947
rect 110 1943 116 1944
rect 110 1939 111 1943
rect 115 1939 116 1943
rect 110 1938 116 1939
rect 1326 1943 1332 1944
rect 1326 1939 1327 1943
rect 1331 1939 1332 1943
rect 1414 1942 1415 1946
rect 1419 1942 1420 1946
rect 1414 1941 1420 1942
rect 1494 1946 1500 1947
rect 1494 1942 1495 1946
rect 1499 1942 1500 1946
rect 1494 1941 1500 1942
rect 1598 1946 1604 1947
rect 1598 1942 1599 1946
rect 1603 1942 1604 1946
rect 1598 1941 1604 1942
rect 1694 1946 1700 1947
rect 1694 1942 1695 1946
rect 1699 1942 1700 1946
rect 1694 1941 1700 1942
rect 1782 1946 1788 1947
rect 1782 1942 1783 1946
rect 1787 1942 1788 1946
rect 1782 1941 1788 1942
rect 1862 1946 1868 1947
rect 1862 1942 1863 1946
rect 1867 1942 1868 1946
rect 1862 1941 1868 1942
rect 1942 1946 1948 1947
rect 1942 1942 1943 1946
rect 1947 1942 1948 1946
rect 1942 1941 1948 1942
rect 2022 1946 2028 1947
rect 2022 1942 2023 1946
rect 2027 1942 2028 1946
rect 2022 1941 2028 1942
rect 2102 1946 2108 1947
rect 2102 1942 2103 1946
rect 2107 1942 2108 1946
rect 2102 1941 2108 1942
rect 1326 1938 1332 1939
rect 350 1934 356 1935
rect 350 1930 351 1934
rect 355 1930 356 1934
rect 350 1929 356 1930
rect 406 1934 412 1935
rect 406 1930 407 1934
rect 411 1930 412 1934
rect 406 1929 412 1930
rect 462 1934 468 1935
rect 462 1930 463 1934
rect 467 1930 468 1934
rect 462 1929 468 1930
rect 518 1934 524 1935
rect 518 1930 519 1934
rect 523 1930 524 1934
rect 518 1929 524 1930
rect 582 1934 588 1935
rect 582 1930 583 1934
rect 587 1930 588 1934
rect 582 1929 588 1930
rect 662 1934 668 1935
rect 662 1930 663 1934
rect 667 1930 668 1934
rect 662 1929 668 1930
rect 758 1934 764 1935
rect 758 1930 759 1934
rect 763 1930 764 1934
rect 758 1929 764 1930
rect 878 1934 884 1935
rect 878 1930 879 1934
rect 883 1930 884 1934
rect 878 1929 884 1930
rect 1014 1934 1020 1935
rect 1014 1930 1015 1934
rect 1019 1930 1020 1934
rect 1014 1929 1020 1930
rect 1158 1934 1164 1935
rect 1158 1930 1159 1934
rect 1163 1930 1164 1934
rect 1158 1929 1164 1930
rect 1286 1934 1292 1935
rect 1286 1930 1287 1934
rect 1291 1930 1292 1934
rect 1286 1929 1292 1930
rect 1718 1918 1724 1919
rect 1718 1914 1719 1918
rect 1723 1914 1724 1918
rect 1718 1913 1724 1914
rect 1774 1918 1780 1919
rect 1774 1914 1775 1918
rect 1779 1914 1780 1918
rect 1774 1913 1780 1914
rect 1830 1918 1836 1919
rect 1830 1914 1831 1918
rect 1835 1914 1836 1918
rect 1830 1913 1836 1914
rect 1886 1918 1892 1919
rect 1886 1914 1887 1918
rect 1891 1914 1892 1918
rect 1886 1913 1892 1914
rect 1942 1918 1948 1919
rect 1942 1914 1943 1918
rect 1947 1914 1948 1918
rect 1942 1913 1948 1914
rect 1998 1918 2004 1919
rect 1998 1914 1999 1918
rect 2003 1914 2004 1918
rect 1998 1913 2004 1914
rect 2054 1918 2060 1919
rect 2054 1914 2055 1918
rect 2059 1914 2060 1918
rect 2054 1913 2060 1914
rect 2118 1918 2124 1919
rect 2118 1914 2119 1918
rect 2123 1914 2124 1918
rect 2118 1913 2124 1914
rect 158 1910 164 1911
rect 158 1906 159 1910
rect 163 1906 164 1910
rect 158 1905 164 1906
rect 230 1910 236 1911
rect 230 1906 231 1910
rect 235 1906 236 1910
rect 230 1905 236 1906
rect 326 1910 332 1911
rect 326 1906 327 1910
rect 331 1906 332 1910
rect 326 1905 332 1906
rect 430 1910 436 1911
rect 430 1906 431 1910
rect 435 1906 436 1910
rect 430 1905 436 1906
rect 542 1910 548 1911
rect 542 1906 543 1910
rect 547 1906 548 1910
rect 542 1905 548 1906
rect 654 1910 660 1911
rect 654 1906 655 1910
rect 659 1906 660 1910
rect 654 1905 660 1906
rect 766 1910 772 1911
rect 766 1906 767 1910
rect 771 1906 772 1910
rect 766 1905 772 1906
rect 878 1910 884 1911
rect 878 1906 879 1910
rect 883 1906 884 1910
rect 878 1905 884 1906
rect 982 1910 988 1911
rect 982 1906 983 1910
rect 987 1906 988 1910
rect 982 1905 988 1906
rect 1086 1910 1092 1911
rect 1086 1906 1087 1910
rect 1091 1906 1092 1910
rect 1086 1905 1092 1906
rect 1198 1910 1204 1911
rect 1198 1906 1199 1910
rect 1203 1906 1204 1910
rect 1198 1905 1204 1906
rect 1286 1910 1292 1911
rect 1286 1906 1287 1910
rect 1291 1906 1292 1910
rect 1286 1905 1292 1906
rect 1366 1909 1372 1910
rect 1366 1905 1367 1909
rect 1371 1905 1372 1909
rect 1366 1904 1372 1905
rect 2582 1909 2588 1910
rect 2582 1905 2583 1909
rect 2587 1905 2588 1909
rect 2582 1904 2588 1905
rect 110 1901 116 1902
rect 110 1897 111 1901
rect 115 1897 116 1901
rect 110 1896 116 1897
rect 1326 1901 1332 1902
rect 1326 1897 1327 1901
rect 1331 1897 1332 1901
rect 1326 1896 1332 1897
rect 1366 1892 1372 1893
rect 2582 1892 2588 1893
rect 1366 1888 1367 1892
rect 1371 1888 1372 1892
rect 1366 1887 1372 1888
rect 1702 1891 1708 1892
rect 1702 1887 1703 1891
rect 1707 1887 1708 1891
rect 1702 1886 1708 1887
rect 1758 1891 1764 1892
rect 1758 1887 1759 1891
rect 1763 1887 1764 1891
rect 1758 1886 1764 1887
rect 1814 1891 1820 1892
rect 1814 1887 1815 1891
rect 1819 1887 1820 1891
rect 1814 1886 1820 1887
rect 1870 1891 1876 1892
rect 1870 1887 1871 1891
rect 1875 1887 1876 1891
rect 1870 1886 1876 1887
rect 1926 1891 1932 1892
rect 1926 1887 1927 1891
rect 1931 1887 1932 1891
rect 1926 1886 1932 1887
rect 1982 1891 1988 1892
rect 1982 1887 1983 1891
rect 1987 1887 1988 1891
rect 1982 1886 1988 1887
rect 2038 1891 2044 1892
rect 2038 1887 2039 1891
rect 2043 1887 2044 1891
rect 2038 1886 2044 1887
rect 2102 1891 2108 1892
rect 2102 1887 2103 1891
rect 2107 1887 2108 1891
rect 2582 1888 2583 1892
rect 2587 1888 2588 1892
rect 2582 1887 2588 1888
rect 2102 1886 2108 1887
rect 110 1884 116 1885
rect 1326 1884 1332 1885
rect 110 1880 111 1884
rect 115 1880 116 1884
rect 110 1879 116 1880
rect 142 1883 148 1884
rect 142 1879 143 1883
rect 147 1879 148 1883
rect 142 1878 148 1879
rect 214 1883 220 1884
rect 214 1879 215 1883
rect 219 1879 220 1883
rect 214 1878 220 1879
rect 310 1883 316 1884
rect 310 1879 311 1883
rect 315 1879 316 1883
rect 310 1878 316 1879
rect 414 1883 420 1884
rect 414 1879 415 1883
rect 419 1879 420 1883
rect 414 1878 420 1879
rect 526 1883 532 1884
rect 526 1879 527 1883
rect 531 1879 532 1883
rect 526 1878 532 1879
rect 638 1883 644 1884
rect 638 1879 639 1883
rect 643 1879 644 1883
rect 638 1878 644 1879
rect 750 1883 756 1884
rect 750 1879 751 1883
rect 755 1879 756 1883
rect 750 1878 756 1879
rect 862 1883 868 1884
rect 862 1879 863 1883
rect 867 1879 868 1883
rect 862 1878 868 1879
rect 966 1883 972 1884
rect 966 1879 967 1883
rect 971 1879 972 1883
rect 966 1878 972 1879
rect 1070 1883 1076 1884
rect 1070 1879 1071 1883
rect 1075 1879 1076 1883
rect 1070 1878 1076 1879
rect 1182 1883 1188 1884
rect 1182 1879 1183 1883
rect 1187 1879 1188 1883
rect 1182 1878 1188 1879
rect 1270 1883 1276 1884
rect 1270 1879 1271 1883
rect 1275 1879 1276 1883
rect 1326 1880 1327 1884
rect 1331 1880 1332 1884
rect 1326 1879 1332 1880
rect 1270 1878 1276 1879
rect 1398 1853 1404 1854
rect 1366 1852 1372 1853
rect 1366 1848 1367 1852
rect 1371 1848 1372 1852
rect 1398 1849 1399 1853
rect 1403 1849 1404 1853
rect 1398 1848 1404 1849
rect 1462 1853 1468 1854
rect 1462 1849 1463 1853
rect 1467 1849 1468 1853
rect 1462 1848 1468 1849
rect 1558 1853 1564 1854
rect 1558 1849 1559 1853
rect 1563 1849 1564 1853
rect 1558 1848 1564 1849
rect 1654 1853 1660 1854
rect 1654 1849 1655 1853
rect 1659 1849 1660 1853
rect 1654 1848 1660 1849
rect 1742 1853 1748 1854
rect 1742 1849 1743 1853
rect 1747 1849 1748 1853
rect 1742 1848 1748 1849
rect 1830 1853 1836 1854
rect 1830 1849 1831 1853
rect 1835 1849 1836 1853
rect 1830 1848 1836 1849
rect 1918 1853 1924 1854
rect 1918 1849 1919 1853
rect 1923 1849 1924 1853
rect 1918 1848 1924 1849
rect 2006 1853 2012 1854
rect 2006 1849 2007 1853
rect 2011 1849 2012 1853
rect 2006 1848 2012 1849
rect 2094 1853 2100 1854
rect 2094 1849 2095 1853
rect 2099 1849 2100 1853
rect 2094 1848 2100 1849
rect 2182 1853 2188 1854
rect 2182 1849 2183 1853
rect 2187 1849 2188 1853
rect 2182 1848 2188 1849
rect 2582 1852 2588 1853
rect 2582 1848 2583 1852
rect 2587 1848 2588 1852
rect 1366 1847 1372 1848
rect 2582 1847 2588 1848
rect 142 1841 148 1842
rect 110 1840 116 1841
rect 110 1836 111 1840
rect 115 1836 116 1840
rect 142 1837 143 1841
rect 147 1837 148 1841
rect 142 1836 148 1837
rect 198 1841 204 1842
rect 198 1837 199 1841
rect 203 1837 204 1841
rect 198 1836 204 1837
rect 262 1841 268 1842
rect 262 1837 263 1841
rect 267 1837 268 1841
rect 262 1836 268 1837
rect 350 1841 356 1842
rect 350 1837 351 1841
rect 355 1837 356 1841
rect 350 1836 356 1837
rect 438 1841 444 1842
rect 438 1837 439 1841
rect 443 1837 444 1841
rect 438 1836 444 1837
rect 534 1841 540 1842
rect 534 1837 535 1841
rect 539 1837 540 1841
rect 534 1836 540 1837
rect 622 1841 628 1842
rect 622 1837 623 1841
rect 627 1837 628 1841
rect 622 1836 628 1837
rect 710 1841 716 1842
rect 710 1837 711 1841
rect 715 1837 716 1841
rect 710 1836 716 1837
rect 790 1841 796 1842
rect 790 1837 791 1841
rect 795 1837 796 1841
rect 790 1836 796 1837
rect 870 1841 876 1842
rect 870 1837 871 1841
rect 875 1837 876 1841
rect 870 1836 876 1837
rect 950 1841 956 1842
rect 950 1837 951 1841
rect 955 1837 956 1841
rect 950 1836 956 1837
rect 1038 1841 1044 1842
rect 1038 1837 1039 1841
rect 1043 1837 1044 1841
rect 1038 1836 1044 1837
rect 1326 1840 1332 1841
rect 1326 1836 1327 1840
rect 1331 1836 1332 1840
rect 110 1835 116 1836
rect 1326 1835 1332 1836
rect 1366 1835 1372 1836
rect 1366 1831 1367 1835
rect 1371 1831 1372 1835
rect 1366 1830 1372 1831
rect 2582 1835 2588 1836
rect 2582 1831 2583 1835
rect 2587 1831 2588 1835
rect 2582 1830 2588 1831
rect 1414 1826 1420 1827
rect 110 1823 116 1824
rect 110 1819 111 1823
rect 115 1819 116 1823
rect 110 1818 116 1819
rect 1326 1823 1332 1824
rect 1326 1819 1327 1823
rect 1331 1819 1332 1823
rect 1414 1822 1415 1826
rect 1419 1822 1420 1826
rect 1414 1821 1420 1822
rect 1478 1826 1484 1827
rect 1478 1822 1479 1826
rect 1483 1822 1484 1826
rect 1478 1821 1484 1822
rect 1574 1826 1580 1827
rect 1574 1822 1575 1826
rect 1579 1822 1580 1826
rect 1574 1821 1580 1822
rect 1670 1826 1676 1827
rect 1670 1822 1671 1826
rect 1675 1822 1676 1826
rect 1670 1821 1676 1822
rect 1758 1826 1764 1827
rect 1758 1822 1759 1826
rect 1763 1822 1764 1826
rect 1758 1821 1764 1822
rect 1846 1826 1852 1827
rect 1846 1822 1847 1826
rect 1851 1822 1852 1826
rect 1846 1821 1852 1822
rect 1934 1826 1940 1827
rect 1934 1822 1935 1826
rect 1939 1822 1940 1826
rect 1934 1821 1940 1822
rect 2022 1826 2028 1827
rect 2022 1822 2023 1826
rect 2027 1822 2028 1826
rect 2022 1821 2028 1822
rect 2110 1826 2116 1827
rect 2110 1822 2111 1826
rect 2115 1822 2116 1826
rect 2110 1821 2116 1822
rect 2198 1826 2204 1827
rect 2198 1822 2199 1826
rect 2203 1822 2204 1826
rect 2198 1821 2204 1822
rect 1326 1818 1332 1819
rect 158 1814 164 1815
rect 158 1810 159 1814
rect 163 1810 164 1814
rect 158 1809 164 1810
rect 214 1814 220 1815
rect 214 1810 215 1814
rect 219 1810 220 1814
rect 214 1809 220 1810
rect 278 1814 284 1815
rect 278 1810 279 1814
rect 283 1810 284 1814
rect 278 1809 284 1810
rect 366 1814 372 1815
rect 366 1810 367 1814
rect 371 1810 372 1814
rect 366 1809 372 1810
rect 454 1814 460 1815
rect 454 1810 455 1814
rect 459 1810 460 1814
rect 454 1809 460 1810
rect 550 1814 556 1815
rect 550 1810 551 1814
rect 555 1810 556 1814
rect 550 1809 556 1810
rect 638 1814 644 1815
rect 638 1810 639 1814
rect 643 1810 644 1814
rect 638 1809 644 1810
rect 726 1814 732 1815
rect 726 1810 727 1814
rect 731 1810 732 1814
rect 726 1809 732 1810
rect 806 1814 812 1815
rect 806 1810 807 1814
rect 811 1810 812 1814
rect 806 1809 812 1810
rect 886 1814 892 1815
rect 886 1810 887 1814
rect 891 1810 892 1814
rect 886 1809 892 1810
rect 966 1814 972 1815
rect 966 1810 967 1814
rect 971 1810 972 1814
rect 966 1809 972 1810
rect 1054 1814 1060 1815
rect 1054 1810 1055 1814
rect 1059 1810 1060 1814
rect 1054 1809 1060 1810
rect 1414 1802 1420 1803
rect 1414 1798 1415 1802
rect 1419 1798 1420 1802
rect 1414 1797 1420 1798
rect 1510 1802 1516 1803
rect 1510 1798 1511 1802
rect 1515 1798 1516 1802
rect 1510 1797 1516 1798
rect 1622 1802 1628 1803
rect 1622 1798 1623 1802
rect 1627 1798 1628 1802
rect 1622 1797 1628 1798
rect 1734 1802 1740 1803
rect 1734 1798 1735 1802
rect 1739 1798 1740 1802
rect 1734 1797 1740 1798
rect 1838 1802 1844 1803
rect 1838 1798 1839 1802
rect 1843 1798 1844 1802
rect 1838 1797 1844 1798
rect 1950 1802 1956 1803
rect 1950 1798 1951 1802
rect 1955 1798 1956 1802
rect 1950 1797 1956 1798
rect 2062 1802 2068 1803
rect 2062 1798 2063 1802
rect 2067 1798 2068 1802
rect 2062 1797 2068 1798
rect 2182 1802 2188 1803
rect 2182 1798 2183 1802
rect 2187 1798 2188 1802
rect 2182 1797 2188 1798
rect 2302 1802 2308 1803
rect 2302 1798 2303 1802
rect 2307 1798 2308 1802
rect 2302 1797 2308 1798
rect 2430 1802 2436 1803
rect 2430 1798 2431 1802
rect 2435 1798 2436 1802
rect 2430 1797 2436 1798
rect 2542 1802 2548 1803
rect 2542 1798 2543 1802
rect 2547 1798 2548 1802
rect 2542 1797 2548 1798
rect 1366 1793 1372 1794
rect 1366 1789 1367 1793
rect 1371 1789 1372 1793
rect 1366 1788 1372 1789
rect 2582 1793 2588 1794
rect 2582 1789 2583 1793
rect 2587 1789 2588 1793
rect 2582 1788 2588 1789
rect 230 1786 236 1787
rect 230 1782 231 1786
rect 235 1782 236 1786
rect 230 1781 236 1782
rect 294 1786 300 1787
rect 294 1782 295 1786
rect 299 1782 300 1786
rect 294 1781 300 1782
rect 366 1786 372 1787
rect 366 1782 367 1786
rect 371 1782 372 1786
rect 366 1781 372 1782
rect 446 1786 452 1787
rect 446 1782 447 1786
rect 451 1782 452 1786
rect 446 1781 452 1782
rect 534 1786 540 1787
rect 534 1782 535 1786
rect 539 1782 540 1786
rect 534 1781 540 1782
rect 622 1786 628 1787
rect 622 1782 623 1786
rect 627 1782 628 1786
rect 622 1781 628 1782
rect 710 1786 716 1787
rect 710 1782 711 1786
rect 715 1782 716 1786
rect 710 1781 716 1782
rect 790 1786 796 1787
rect 790 1782 791 1786
rect 795 1782 796 1786
rect 790 1781 796 1782
rect 870 1786 876 1787
rect 870 1782 871 1786
rect 875 1782 876 1786
rect 870 1781 876 1782
rect 950 1786 956 1787
rect 950 1782 951 1786
rect 955 1782 956 1786
rect 950 1781 956 1782
rect 1030 1786 1036 1787
rect 1030 1782 1031 1786
rect 1035 1782 1036 1786
rect 1030 1781 1036 1782
rect 1118 1786 1124 1787
rect 1118 1782 1119 1786
rect 1123 1782 1124 1786
rect 1118 1781 1124 1782
rect 110 1777 116 1778
rect 110 1773 111 1777
rect 115 1773 116 1777
rect 110 1772 116 1773
rect 1326 1777 1332 1778
rect 1326 1773 1327 1777
rect 1331 1773 1332 1777
rect 1326 1772 1332 1773
rect 1366 1776 1372 1777
rect 2582 1776 2588 1777
rect 1366 1772 1367 1776
rect 1371 1772 1372 1776
rect 1366 1771 1372 1772
rect 1398 1775 1404 1776
rect 1398 1771 1399 1775
rect 1403 1771 1404 1775
rect 1398 1770 1404 1771
rect 1494 1775 1500 1776
rect 1494 1771 1495 1775
rect 1499 1771 1500 1775
rect 1494 1770 1500 1771
rect 1606 1775 1612 1776
rect 1606 1771 1607 1775
rect 1611 1771 1612 1775
rect 1606 1770 1612 1771
rect 1718 1775 1724 1776
rect 1718 1771 1719 1775
rect 1723 1771 1724 1775
rect 1718 1770 1724 1771
rect 1822 1775 1828 1776
rect 1822 1771 1823 1775
rect 1827 1771 1828 1775
rect 1822 1770 1828 1771
rect 1934 1775 1940 1776
rect 1934 1771 1935 1775
rect 1939 1771 1940 1775
rect 1934 1770 1940 1771
rect 2046 1775 2052 1776
rect 2046 1771 2047 1775
rect 2051 1771 2052 1775
rect 2046 1770 2052 1771
rect 2166 1775 2172 1776
rect 2166 1771 2167 1775
rect 2171 1771 2172 1775
rect 2166 1770 2172 1771
rect 2286 1775 2292 1776
rect 2286 1771 2287 1775
rect 2291 1771 2292 1775
rect 2286 1770 2292 1771
rect 2414 1775 2420 1776
rect 2414 1771 2415 1775
rect 2419 1771 2420 1775
rect 2414 1770 2420 1771
rect 2526 1775 2532 1776
rect 2526 1771 2527 1775
rect 2531 1771 2532 1775
rect 2582 1772 2583 1776
rect 2587 1772 2588 1776
rect 2582 1771 2588 1772
rect 2526 1770 2532 1771
rect 110 1760 116 1761
rect 1326 1760 1332 1761
rect 110 1756 111 1760
rect 115 1756 116 1760
rect 110 1755 116 1756
rect 214 1759 220 1760
rect 214 1755 215 1759
rect 219 1755 220 1759
rect 214 1754 220 1755
rect 278 1759 284 1760
rect 278 1755 279 1759
rect 283 1755 284 1759
rect 278 1754 284 1755
rect 350 1759 356 1760
rect 350 1755 351 1759
rect 355 1755 356 1759
rect 350 1754 356 1755
rect 430 1759 436 1760
rect 430 1755 431 1759
rect 435 1755 436 1759
rect 430 1754 436 1755
rect 518 1759 524 1760
rect 518 1755 519 1759
rect 523 1755 524 1759
rect 518 1754 524 1755
rect 606 1759 612 1760
rect 606 1755 607 1759
rect 611 1755 612 1759
rect 606 1754 612 1755
rect 694 1759 700 1760
rect 694 1755 695 1759
rect 699 1755 700 1759
rect 694 1754 700 1755
rect 774 1759 780 1760
rect 774 1755 775 1759
rect 779 1755 780 1759
rect 774 1754 780 1755
rect 854 1759 860 1760
rect 854 1755 855 1759
rect 859 1755 860 1759
rect 854 1754 860 1755
rect 934 1759 940 1760
rect 934 1755 935 1759
rect 939 1755 940 1759
rect 934 1754 940 1755
rect 1014 1759 1020 1760
rect 1014 1755 1015 1759
rect 1019 1755 1020 1759
rect 1014 1754 1020 1755
rect 1102 1759 1108 1760
rect 1102 1755 1103 1759
rect 1107 1755 1108 1759
rect 1326 1756 1327 1760
rect 1331 1756 1332 1760
rect 1326 1755 1332 1756
rect 1102 1754 1108 1755
rect 1438 1741 1444 1742
rect 1366 1740 1372 1741
rect 1366 1736 1367 1740
rect 1371 1736 1372 1740
rect 1438 1737 1439 1741
rect 1443 1737 1444 1741
rect 1438 1736 1444 1737
rect 1518 1741 1524 1742
rect 1518 1737 1519 1741
rect 1523 1737 1524 1741
rect 1518 1736 1524 1737
rect 1614 1741 1620 1742
rect 1614 1737 1615 1741
rect 1619 1737 1620 1741
rect 1614 1736 1620 1737
rect 1718 1741 1724 1742
rect 1718 1737 1719 1741
rect 1723 1737 1724 1741
rect 1718 1736 1724 1737
rect 1822 1741 1828 1742
rect 1822 1737 1823 1741
rect 1827 1737 1828 1741
rect 1822 1736 1828 1737
rect 1926 1741 1932 1742
rect 1926 1737 1927 1741
rect 1931 1737 1932 1741
rect 1926 1736 1932 1737
rect 2022 1741 2028 1742
rect 2022 1737 2023 1741
rect 2027 1737 2028 1741
rect 2022 1736 2028 1737
rect 2118 1741 2124 1742
rect 2118 1737 2119 1741
rect 2123 1737 2124 1741
rect 2118 1736 2124 1737
rect 2206 1741 2212 1742
rect 2206 1737 2207 1741
rect 2211 1737 2212 1741
rect 2206 1736 2212 1737
rect 2286 1741 2292 1742
rect 2286 1737 2287 1741
rect 2291 1737 2292 1741
rect 2286 1736 2292 1737
rect 2374 1741 2380 1742
rect 2374 1737 2375 1741
rect 2379 1737 2380 1741
rect 2374 1736 2380 1737
rect 2462 1741 2468 1742
rect 2462 1737 2463 1741
rect 2467 1737 2468 1741
rect 2462 1736 2468 1737
rect 2526 1741 2532 1742
rect 2526 1737 2527 1741
rect 2531 1737 2532 1741
rect 2526 1736 2532 1737
rect 2582 1740 2588 1741
rect 2582 1736 2583 1740
rect 2587 1736 2588 1740
rect 1366 1735 1372 1736
rect 2582 1735 2588 1736
rect 1366 1723 1372 1724
rect 350 1721 356 1722
rect 110 1720 116 1721
rect 110 1716 111 1720
rect 115 1716 116 1720
rect 350 1717 351 1721
rect 355 1717 356 1721
rect 350 1716 356 1717
rect 406 1721 412 1722
rect 406 1717 407 1721
rect 411 1717 412 1721
rect 406 1716 412 1717
rect 470 1721 476 1722
rect 470 1717 471 1721
rect 475 1717 476 1721
rect 470 1716 476 1717
rect 550 1721 556 1722
rect 550 1717 551 1721
rect 555 1717 556 1721
rect 550 1716 556 1717
rect 638 1721 644 1722
rect 638 1717 639 1721
rect 643 1717 644 1721
rect 638 1716 644 1717
rect 726 1721 732 1722
rect 726 1717 727 1721
rect 731 1717 732 1721
rect 726 1716 732 1717
rect 822 1721 828 1722
rect 822 1717 823 1721
rect 827 1717 828 1721
rect 822 1716 828 1717
rect 918 1721 924 1722
rect 918 1717 919 1721
rect 923 1717 924 1721
rect 918 1716 924 1717
rect 1014 1721 1020 1722
rect 1014 1717 1015 1721
rect 1019 1717 1020 1721
rect 1014 1716 1020 1717
rect 1110 1721 1116 1722
rect 1110 1717 1111 1721
rect 1115 1717 1116 1721
rect 1110 1716 1116 1717
rect 1206 1721 1212 1722
rect 1206 1717 1207 1721
rect 1211 1717 1212 1721
rect 1206 1716 1212 1717
rect 1326 1720 1332 1721
rect 1326 1716 1327 1720
rect 1331 1716 1332 1720
rect 1366 1719 1367 1723
rect 1371 1719 1372 1723
rect 1366 1718 1372 1719
rect 2582 1723 2588 1724
rect 2582 1719 2583 1723
rect 2587 1719 2588 1723
rect 2582 1718 2588 1719
rect 110 1715 116 1716
rect 1326 1715 1332 1716
rect 1454 1714 1460 1715
rect 1454 1710 1455 1714
rect 1459 1710 1460 1714
rect 1454 1709 1460 1710
rect 1534 1714 1540 1715
rect 1534 1710 1535 1714
rect 1539 1710 1540 1714
rect 1534 1709 1540 1710
rect 1630 1714 1636 1715
rect 1630 1710 1631 1714
rect 1635 1710 1636 1714
rect 1630 1709 1636 1710
rect 1734 1714 1740 1715
rect 1734 1710 1735 1714
rect 1739 1710 1740 1714
rect 1734 1709 1740 1710
rect 1838 1714 1844 1715
rect 1838 1710 1839 1714
rect 1843 1710 1844 1714
rect 1838 1709 1844 1710
rect 1942 1714 1948 1715
rect 1942 1710 1943 1714
rect 1947 1710 1948 1714
rect 1942 1709 1948 1710
rect 2038 1714 2044 1715
rect 2038 1710 2039 1714
rect 2043 1710 2044 1714
rect 2038 1709 2044 1710
rect 2134 1714 2140 1715
rect 2134 1710 2135 1714
rect 2139 1710 2140 1714
rect 2134 1709 2140 1710
rect 2222 1714 2228 1715
rect 2222 1710 2223 1714
rect 2227 1710 2228 1714
rect 2222 1709 2228 1710
rect 2302 1714 2308 1715
rect 2302 1710 2303 1714
rect 2307 1710 2308 1714
rect 2302 1709 2308 1710
rect 2390 1714 2396 1715
rect 2390 1710 2391 1714
rect 2395 1710 2396 1714
rect 2390 1709 2396 1710
rect 2478 1714 2484 1715
rect 2478 1710 2479 1714
rect 2483 1710 2484 1714
rect 2478 1709 2484 1710
rect 2542 1714 2548 1715
rect 2542 1710 2543 1714
rect 2547 1710 2548 1714
rect 2542 1709 2548 1710
rect 110 1703 116 1704
rect 110 1699 111 1703
rect 115 1699 116 1703
rect 110 1698 116 1699
rect 1326 1703 1332 1704
rect 1326 1699 1327 1703
rect 1331 1699 1332 1703
rect 1326 1698 1332 1699
rect 366 1694 372 1695
rect 366 1690 367 1694
rect 371 1690 372 1694
rect 366 1689 372 1690
rect 422 1694 428 1695
rect 422 1690 423 1694
rect 427 1690 428 1694
rect 422 1689 428 1690
rect 486 1694 492 1695
rect 486 1690 487 1694
rect 491 1690 492 1694
rect 486 1689 492 1690
rect 566 1694 572 1695
rect 566 1690 567 1694
rect 571 1690 572 1694
rect 566 1689 572 1690
rect 654 1694 660 1695
rect 654 1690 655 1694
rect 659 1690 660 1694
rect 654 1689 660 1690
rect 742 1694 748 1695
rect 742 1690 743 1694
rect 747 1690 748 1694
rect 742 1689 748 1690
rect 838 1694 844 1695
rect 838 1690 839 1694
rect 843 1690 844 1694
rect 838 1689 844 1690
rect 934 1694 940 1695
rect 934 1690 935 1694
rect 939 1690 940 1694
rect 934 1689 940 1690
rect 1030 1694 1036 1695
rect 1030 1690 1031 1694
rect 1035 1690 1036 1694
rect 1030 1689 1036 1690
rect 1126 1694 1132 1695
rect 1126 1690 1127 1694
rect 1131 1690 1132 1694
rect 1126 1689 1132 1690
rect 1222 1694 1228 1695
rect 1222 1690 1223 1694
rect 1227 1690 1228 1694
rect 1222 1689 1228 1690
rect 1558 1678 1564 1679
rect 1558 1674 1559 1678
rect 1563 1674 1564 1678
rect 1558 1673 1564 1674
rect 1630 1678 1636 1679
rect 1630 1674 1631 1678
rect 1635 1674 1636 1678
rect 1630 1673 1636 1674
rect 1710 1678 1716 1679
rect 1710 1674 1711 1678
rect 1715 1674 1716 1678
rect 1710 1673 1716 1674
rect 1798 1678 1804 1679
rect 1798 1674 1799 1678
rect 1803 1674 1804 1678
rect 1798 1673 1804 1674
rect 1886 1678 1892 1679
rect 1886 1674 1887 1678
rect 1891 1674 1892 1678
rect 1886 1673 1892 1674
rect 1974 1678 1980 1679
rect 1974 1674 1975 1678
rect 1979 1674 1980 1678
rect 1974 1673 1980 1674
rect 2062 1678 2068 1679
rect 2062 1674 2063 1678
rect 2067 1674 2068 1678
rect 2062 1673 2068 1674
rect 2142 1678 2148 1679
rect 2142 1674 2143 1678
rect 2147 1674 2148 1678
rect 2142 1673 2148 1674
rect 2214 1678 2220 1679
rect 2214 1674 2215 1678
rect 2219 1674 2220 1678
rect 2214 1673 2220 1674
rect 2286 1678 2292 1679
rect 2286 1674 2287 1678
rect 2291 1674 2292 1678
rect 2286 1673 2292 1674
rect 2350 1678 2356 1679
rect 2350 1674 2351 1678
rect 2355 1674 2356 1678
rect 2350 1673 2356 1674
rect 2422 1678 2428 1679
rect 2422 1674 2423 1678
rect 2427 1674 2428 1678
rect 2422 1673 2428 1674
rect 2486 1678 2492 1679
rect 2486 1674 2487 1678
rect 2491 1674 2492 1678
rect 2486 1673 2492 1674
rect 2542 1678 2548 1679
rect 2542 1674 2543 1678
rect 2547 1674 2548 1678
rect 2542 1673 2548 1674
rect 1366 1669 1372 1670
rect 398 1666 404 1667
rect 398 1662 399 1666
rect 403 1662 404 1666
rect 398 1661 404 1662
rect 454 1666 460 1667
rect 454 1662 455 1666
rect 459 1662 460 1666
rect 454 1661 460 1662
rect 510 1666 516 1667
rect 510 1662 511 1666
rect 515 1662 516 1666
rect 510 1661 516 1662
rect 574 1666 580 1667
rect 574 1662 575 1666
rect 579 1662 580 1666
rect 574 1661 580 1662
rect 646 1666 652 1667
rect 646 1662 647 1666
rect 651 1662 652 1666
rect 646 1661 652 1662
rect 726 1666 732 1667
rect 726 1662 727 1666
rect 731 1662 732 1666
rect 726 1661 732 1662
rect 806 1666 812 1667
rect 806 1662 807 1666
rect 811 1662 812 1666
rect 806 1661 812 1662
rect 886 1666 892 1667
rect 886 1662 887 1666
rect 891 1662 892 1666
rect 886 1661 892 1662
rect 966 1666 972 1667
rect 966 1662 967 1666
rect 971 1662 972 1666
rect 966 1661 972 1662
rect 1046 1666 1052 1667
rect 1046 1662 1047 1666
rect 1051 1662 1052 1666
rect 1046 1661 1052 1662
rect 1134 1666 1140 1667
rect 1134 1662 1135 1666
rect 1139 1662 1140 1666
rect 1134 1661 1140 1662
rect 1222 1666 1228 1667
rect 1222 1662 1223 1666
rect 1227 1662 1228 1666
rect 1222 1661 1228 1662
rect 1286 1666 1292 1667
rect 1286 1662 1287 1666
rect 1291 1662 1292 1666
rect 1366 1665 1367 1669
rect 1371 1665 1372 1669
rect 1366 1664 1372 1665
rect 2582 1669 2588 1670
rect 2582 1665 2583 1669
rect 2587 1665 2588 1669
rect 2582 1664 2588 1665
rect 1286 1661 1292 1662
rect 110 1657 116 1658
rect 110 1653 111 1657
rect 115 1653 116 1657
rect 110 1652 116 1653
rect 1326 1657 1332 1658
rect 1326 1653 1327 1657
rect 1331 1653 1332 1657
rect 1326 1652 1332 1653
rect 1366 1652 1372 1653
rect 2582 1652 2588 1653
rect 1366 1648 1367 1652
rect 1371 1648 1372 1652
rect 1366 1647 1372 1648
rect 1542 1651 1548 1652
rect 1542 1647 1543 1651
rect 1547 1647 1548 1651
rect 1542 1646 1548 1647
rect 1614 1651 1620 1652
rect 1614 1647 1615 1651
rect 1619 1647 1620 1651
rect 1614 1646 1620 1647
rect 1694 1651 1700 1652
rect 1694 1647 1695 1651
rect 1699 1647 1700 1651
rect 1694 1646 1700 1647
rect 1782 1651 1788 1652
rect 1782 1647 1783 1651
rect 1787 1647 1788 1651
rect 1782 1646 1788 1647
rect 1870 1651 1876 1652
rect 1870 1647 1871 1651
rect 1875 1647 1876 1651
rect 1870 1646 1876 1647
rect 1958 1651 1964 1652
rect 1958 1647 1959 1651
rect 1963 1647 1964 1651
rect 1958 1646 1964 1647
rect 2046 1651 2052 1652
rect 2046 1647 2047 1651
rect 2051 1647 2052 1651
rect 2046 1646 2052 1647
rect 2126 1651 2132 1652
rect 2126 1647 2127 1651
rect 2131 1647 2132 1651
rect 2126 1646 2132 1647
rect 2198 1651 2204 1652
rect 2198 1647 2199 1651
rect 2203 1647 2204 1651
rect 2198 1646 2204 1647
rect 2270 1651 2276 1652
rect 2270 1647 2271 1651
rect 2275 1647 2276 1651
rect 2270 1646 2276 1647
rect 2334 1651 2340 1652
rect 2334 1647 2335 1651
rect 2339 1647 2340 1651
rect 2334 1646 2340 1647
rect 2406 1651 2412 1652
rect 2406 1647 2407 1651
rect 2411 1647 2412 1651
rect 2406 1646 2412 1647
rect 2470 1651 2476 1652
rect 2470 1647 2471 1651
rect 2475 1647 2476 1651
rect 2470 1646 2476 1647
rect 2526 1651 2532 1652
rect 2526 1647 2527 1651
rect 2531 1647 2532 1651
rect 2582 1648 2583 1652
rect 2587 1648 2588 1652
rect 2582 1647 2588 1648
rect 2526 1646 2532 1647
rect 110 1640 116 1641
rect 1326 1640 1332 1641
rect 110 1636 111 1640
rect 115 1636 116 1640
rect 110 1635 116 1636
rect 382 1639 388 1640
rect 382 1635 383 1639
rect 387 1635 388 1639
rect 382 1634 388 1635
rect 438 1639 444 1640
rect 438 1635 439 1639
rect 443 1635 444 1639
rect 438 1634 444 1635
rect 494 1639 500 1640
rect 494 1635 495 1639
rect 499 1635 500 1639
rect 494 1634 500 1635
rect 558 1639 564 1640
rect 558 1635 559 1639
rect 563 1635 564 1639
rect 558 1634 564 1635
rect 630 1639 636 1640
rect 630 1635 631 1639
rect 635 1635 636 1639
rect 630 1634 636 1635
rect 710 1639 716 1640
rect 710 1635 711 1639
rect 715 1635 716 1639
rect 710 1634 716 1635
rect 790 1639 796 1640
rect 790 1635 791 1639
rect 795 1635 796 1639
rect 790 1634 796 1635
rect 870 1639 876 1640
rect 870 1635 871 1639
rect 875 1635 876 1639
rect 870 1634 876 1635
rect 950 1639 956 1640
rect 950 1635 951 1639
rect 955 1635 956 1639
rect 950 1634 956 1635
rect 1030 1639 1036 1640
rect 1030 1635 1031 1639
rect 1035 1635 1036 1639
rect 1030 1634 1036 1635
rect 1118 1639 1124 1640
rect 1118 1635 1119 1639
rect 1123 1635 1124 1639
rect 1118 1634 1124 1635
rect 1206 1639 1212 1640
rect 1206 1635 1207 1639
rect 1211 1635 1212 1639
rect 1206 1634 1212 1635
rect 1270 1639 1276 1640
rect 1270 1635 1271 1639
rect 1275 1635 1276 1639
rect 1326 1636 1327 1640
rect 1331 1636 1332 1640
rect 1326 1635 1332 1636
rect 1270 1634 1276 1635
rect 1574 1605 1580 1606
rect 1366 1604 1372 1605
rect 1366 1600 1367 1604
rect 1371 1600 1372 1604
rect 1574 1601 1575 1605
rect 1579 1601 1580 1605
rect 1574 1600 1580 1601
rect 1630 1605 1636 1606
rect 1630 1601 1631 1605
rect 1635 1601 1636 1605
rect 1630 1600 1636 1601
rect 1686 1605 1692 1606
rect 1686 1601 1687 1605
rect 1691 1601 1692 1605
rect 1686 1600 1692 1601
rect 1750 1605 1756 1606
rect 1750 1601 1751 1605
rect 1755 1601 1756 1605
rect 1750 1600 1756 1601
rect 1830 1605 1836 1606
rect 1830 1601 1831 1605
rect 1835 1601 1836 1605
rect 1830 1600 1836 1601
rect 1918 1605 1924 1606
rect 1918 1601 1919 1605
rect 1923 1601 1924 1605
rect 1918 1600 1924 1601
rect 2006 1605 2012 1606
rect 2006 1601 2007 1605
rect 2011 1601 2012 1605
rect 2006 1600 2012 1601
rect 2102 1605 2108 1606
rect 2102 1601 2103 1605
rect 2107 1601 2108 1605
rect 2102 1600 2108 1601
rect 2206 1605 2212 1606
rect 2206 1601 2207 1605
rect 2211 1601 2212 1605
rect 2206 1600 2212 1601
rect 2318 1605 2324 1606
rect 2318 1601 2319 1605
rect 2323 1601 2324 1605
rect 2318 1600 2324 1601
rect 2430 1605 2436 1606
rect 2430 1601 2431 1605
rect 2435 1601 2436 1605
rect 2430 1600 2436 1601
rect 2526 1605 2532 1606
rect 2526 1601 2527 1605
rect 2531 1601 2532 1605
rect 2526 1600 2532 1601
rect 2582 1604 2588 1605
rect 2582 1600 2583 1604
rect 2587 1600 2588 1604
rect 1366 1599 1372 1600
rect 2582 1599 2588 1600
rect 286 1589 292 1590
rect 110 1588 116 1589
rect 110 1584 111 1588
rect 115 1584 116 1588
rect 286 1585 287 1589
rect 291 1585 292 1589
rect 286 1584 292 1585
rect 366 1589 372 1590
rect 366 1585 367 1589
rect 371 1585 372 1589
rect 366 1584 372 1585
rect 454 1589 460 1590
rect 454 1585 455 1589
rect 459 1585 460 1589
rect 454 1584 460 1585
rect 550 1589 556 1590
rect 550 1585 551 1589
rect 555 1585 556 1589
rect 550 1584 556 1585
rect 646 1589 652 1590
rect 646 1585 647 1589
rect 651 1585 652 1589
rect 646 1584 652 1585
rect 734 1589 740 1590
rect 734 1585 735 1589
rect 739 1585 740 1589
rect 734 1584 740 1585
rect 822 1589 828 1590
rect 822 1585 823 1589
rect 827 1585 828 1589
rect 822 1584 828 1585
rect 902 1589 908 1590
rect 902 1585 903 1589
rect 907 1585 908 1589
rect 902 1584 908 1585
rect 982 1589 988 1590
rect 982 1585 983 1589
rect 987 1585 988 1589
rect 982 1584 988 1585
rect 1062 1589 1068 1590
rect 1062 1585 1063 1589
rect 1067 1585 1068 1589
rect 1062 1584 1068 1585
rect 1150 1589 1156 1590
rect 1150 1585 1151 1589
rect 1155 1585 1156 1589
rect 1150 1584 1156 1585
rect 1326 1588 1332 1589
rect 1326 1584 1327 1588
rect 1331 1584 1332 1588
rect 110 1583 116 1584
rect 1326 1583 1332 1584
rect 1366 1587 1372 1588
rect 1366 1583 1367 1587
rect 1371 1583 1372 1587
rect 1366 1582 1372 1583
rect 2582 1587 2588 1588
rect 2582 1583 2583 1587
rect 2587 1583 2588 1587
rect 2582 1582 2588 1583
rect 1590 1578 1596 1579
rect 1590 1574 1591 1578
rect 1595 1574 1596 1578
rect 1590 1573 1596 1574
rect 1646 1578 1652 1579
rect 1646 1574 1647 1578
rect 1651 1574 1652 1578
rect 1646 1573 1652 1574
rect 1702 1578 1708 1579
rect 1702 1574 1703 1578
rect 1707 1574 1708 1578
rect 1702 1573 1708 1574
rect 1766 1578 1772 1579
rect 1766 1574 1767 1578
rect 1771 1574 1772 1578
rect 1766 1573 1772 1574
rect 1846 1578 1852 1579
rect 1846 1574 1847 1578
rect 1851 1574 1852 1578
rect 1846 1573 1852 1574
rect 1934 1578 1940 1579
rect 1934 1574 1935 1578
rect 1939 1574 1940 1578
rect 1934 1573 1940 1574
rect 2022 1578 2028 1579
rect 2022 1574 2023 1578
rect 2027 1574 2028 1578
rect 2022 1573 2028 1574
rect 2118 1578 2124 1579
rect 2118 1574 2119 1578
rect 2123 1574 2124 1578
rect 2118 1573 2124 1574
rect 2222 1578 2228 1579
rect 2222 1574 2223 1578
rect 2227 1574 2228 1578
rect 2222 1573 2228 1574
rect 2334 1578 2340 1579
rect 2334 1574 2335 1578
rect 2339 1574 2340 1578
rect 2334 1573 2340 1574
rect 2446 1578 2452 1579
rect 2446 1574 2447 1578
rect 2451 1574 2452 1578
rect 2446 1573 2452 1574
rect 2542 1578 2548 1579
rect 2542 1574 2543 1578
rect 2547 1574 2548 1578
rect 2542 1573 2548 1574
rect 110 1571 116 1572
rect 110 1567 111 1571
rect 115 1567 116 1571
rect 110 1566 116 1567
rect 1326 1571 1332 1572
rect 1326 1567 1327 1571
rect 1331 1567 1332 1571
rect 1326 1566 1332 1567
rect 302 1562 308 1563
rect 302 1558 303 1562
rect 307 1558 308 1562
rect 302 1557 308 1558
rect 382 1562 388 1563
rect 382 1558 383 1562
rect 387 1558 388 1562
rect 382 1557 388 1558
rect 470 1562 476 1563
rect 470 1558 471 1562
rect 475 1558 476 1562
rect 470 1557 476 1558
rect 566 1562 572 1563
rect 566 1558 567 1562
rect 571 1558 572 1562
rect 566 1557 572 1558
rect 662 1562 668 1563
rect 662 1558 663 1562
rect 667 1558 668 1562
rect 662 1557 668 1558
rect 750 1562 756 1563
rect 750 1558 751 1562
rect 755 1558 756 1562
rect 750 1557 756 1558
rect 838 1562 844 1563
rect 838 1558 839 1562
rect 843 1558 844 1562
rect 838 1557 844 1558
rect 918 1562 924 1563
rect 918 1558 919 1562
rect 923 1558 924 1562
rect 918 1557 924 1558
rect 998 1562 1004 1563
rect 998 1558 999 1562
rect 1003 1558 1004 1562
rect 998 1557 1004 1558
rect 1078 1562 1084 1563
rect 1078 1558 1079 1562
rect 1083 1558 1084 1562
rect 1078 1557 1084 1558
rect 1166 1562 1172 1563
rect 1166 1558 1167 1562
rect 1171 1558 1172 1562
rect 1166 1557 1172 1558
rect 1678 1550 1684 1551
rect 1678 1546 1679 1550
rect 1683 1546 1684 1550
rect 1678 1545 1684 1546
rect 1734 1550 1740 1551
rect 1734 1546 1735 1550
rect 1739 1546 1740 1550
rect 1734 1545 1740 1546
rect 1790 1550 1796 1551
rect 1790 1546 1791 1550
rect 1795 1546 1796 1550
rect 1790 1545 1796 1546
rect 1854 1550 1860 1551
rect 1854 1546 1855 1550
rect 1859 1546 1860 1550
rect 1854 1545 1860 1546
rect 1926 1550 1932 1551
rect 1926 1546 1927 1550
rect 1931 1546 1932 1550
rect 1926 1545 1932 1546
rect 2006 1550 2012 1551
rect 2006 1546 2007 1550
rect 2011 1546 2012 1550
rect 2006 1545 2012 1546
rect 2086 1550 2092 1551
rect 2086 1546 2087 1550
rect 2091 1546 2092 1550
rect 2086 1545 2092 1546
rect 2166 1550 2172 1551
rect 2166 1546 2167 1550
rect 2171 1546 2172 1550
rect 2166 1545 2172 1546
rect 2246 1550 2252 1551
rect 2246 1546 2247 1550
rect 2251 1546 2252 1550
rect 2246 1545 2252 1546
rect 2326 1550 2332 1551
rect 2326 1546 2327 1550
rect 2331 1546 2332 1550
rect 2326 1545 2332 1546
rect 2406 1550 2412 1551
rect 2406 1546 2407 1550
rect 2411 1546 2412 1550
rect 2406 1545 2412 1546
rect 2486 1550 2492 1551
rect 2486 1546 2487 1550
rect 2491 1546 2492 1550
rect 2486 1545 2492 1546
rect 2542 1550 2548 1551
rect 2542 1546 2543 1550
rect 2547 1546 2548 1550
rect 2542 1545 2548 1546
rect 1366 1541 1372 1542
rect 278 1538 284 1539
rect 278 1534 279 1538
rect 283 1534 284 1538
rect 278 1533 284 1534
rect 334 1538 340 1539
rect 334 1534 335 1538
rect 339 1534 340 1538
rect 334 1533 340 1534
rect 398 1538 404 1539
rect 398 1534 399 1538
rect 403 1534 404 1538
rect 398 1533 404 1534
rect 470 1538 476 1539
rect 470 1534 471 1538
rect 475 1534 476 1538
rect 470 1533 476 1534
rect 542 1538 548 1539
rect 542 1534 543 1538
rect 547 1534 548 1538
rect 542 1533 548 1534
rect 614 1538 620 1539
rect 614 1534 615 1538
rect 619 1534 620 1538
rect 614 1533 620 1534
rect 686 1538 692 1539
rect 686 1534 687 1538
rect 691 1534 692 1538
rect 686 1533 692 1534
rect 758 1538 764 1539
rect 758 1534 759 1538
rect 763 1534 764 1538
rect 758 1533 764 1534
rect 830 1538 836 1539
rect 830 1534 831 1538
rect 835 1534 836 1538
rect 830 1533 836 1534
rect 902 1538 908 1539
rect 902 1534 903 1538
rect 907 1534 908 1538
rect 902 1533 908 1534
rect 974 1538 980 1539
rect 974 1534 975 1538
rect 979 1534 980 1538
rect 974 1533 980 1534
rect 1054 1538 1060 1539
rect 1054 1534 1055 1538
rect 1059 1534 1060 1538
rect 1366 1537 1367 1541
rect 1371 1537 1372 1541
rect 1366 1536 1372 1537
rect 2582 1541 2588 1542
rect 2582 1537 2583 1541
rect 2587 1537 2588 1541
rect 2582 1536 2588 1537
rect 1054 1533 1060 1534
rect 110 1529 116 1530
rect 110 1525 111 1529
rect 115 1525 116 1529
rect 110 1524 116 1525
rect 1326 1529 1332 1530
rect 1326 1525 1327 1529
rect 1331 1525 1332 1529
rect 1326 1524 1332 1525
rect 1366 1524 1372 1525
rect 2582 1524 2588 1525
rect 1366 1520 1367 1524
rect 1371 1520 1372 1524
rect 1366 1519 1372 1520
rect 1662 1523 1668 1524
rect 1662 1519 1663 1523
rect 1667 1519 1668 1523
rect 1662 1518 1668 1519
rect 1718 1523 1724 1524
rect 1718 1519 1719 1523
rect 1723 1519 1724 1523
rect 1718 1518 1724 1519
rect 1774 1523 1780 1524
rect 1774 1519 1775 1523
rect 1779 1519 1780 1523
rect 1774 1518 1780 1519
rect 1838 1523 1844 1524
rect 1838 1519 1839 1523
rect 1843 1519 1844 1523
rect 1838 1518 1844 1519
rect 1910 1523 1916 1524
rect 1910 1519 1911 1523
rect 1915 1519 1916 1523
rect 1910 1518 1916 1519
rect 1990 1523 1996 1524
rect 1990 1519 1991 1523
rect 1995 1519 1996 1523
rect 1990 1518 1996 1519
rect 2070 1523 2076 1524
rect 2070 1519 2071 1523
rect 2075 1519 2076 1523
rect 2070 1518 2076 1519
rect 2150 1523 2156 1524
rect 2150 1519 2151 1523
rect 2155 1519 2156 1523
rect 2150 1518 2156 1519
rect 2230 1523 2236 1524
rect 2230 1519 2231 1523
rect 2235 1519 2236 1523
rect 2230 1518 2236 1519
rect 2310 1523 2316 1524
rect 2310 1519 2311 1523
rect 2315 1519 2316 1523
rect 2310 1518 2316 1519
rect 2390 1523 2396 1524
rect 2390 1519 2391 1523
rect 2395 1519 2396 1523
rect 2390 1518 2396 1519
rect 2470 1523 2476 1524
rect 2470 1519 2471 1523
rect 2475 1519 2476 1523
rect 2470 1518 2476 1519
rect 2526 1523 2532 1524
rect 2526 1519 2527 1523
rect 2531 1519 2532 1523
rect 2582 1520 2583 1524
rect 2587 1520 2588 1524
rect 2582 1519 2588 1520
rect 2526 1518 2532 1519
rect 110 1512 116 1513
rect 1326 1512 1332 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 110 1507 116 1508
rect 262 1511 268 1512
rect 262 1507 263 1511
rect 267 1507 268 1511
rect 262 1506 268 1507
rect 318 1511 324 1512
rect 318 1507 319 1511
rect 323 1507 324 1511
rect 318 1506 324 1507
rect 382 1511 388 1512
rect 382 1507 383 1511
rect 387 1507 388 1511
rect 382 1506 388 1507
rect 454 1511 460 1512
rect 454 1507 455 1511
rect 459 1507 460 1511
rect 454 1506 460 1507
rect 526 1511 532 1512
rect 526 1507 527 1511
rect 531 1507 532 1511
rect 526 1506 532 1507
rect 598 1511 604 1512
rect 598 1507 599 1511
rect 603 1507 604 1511
rect 598 1506 604 1507
rect 670 1511 676 1512
rect 670 1507 671 1511
rect 675 1507 676 1511
rect 670 1506 676 1507
rect 742 1511 748 1512
rect 742 1507 743 1511
rect 747 1507 748 1511
rect 742 1506 748 1507
rect 814 1511 820 1512
rect 814 1507 815 1511
rect 819 1507 820 1511
rect 814 1506 820 1507
rect 886 1511 892 1512
rect 886 1507 887 1511
rect 891 1507 892 1511
rect 886 1506 892 1507
rect 958 1511 964 1512
rect 958 1507 959 1511
rect 963 1507 964 1511
rect 958 1506 964 1507
rect 1038 1511 1044 1512
rect 1038 1507 1039 1511
rect 1043 1507 1044 1511
rect 1326 1508 1327 1512
rect 1331 1508 1332 1512
rect 1326 1507 1332 1508
rect 1038 1506 1044 1507
rect 1518 1481 1524 1482
rect 1366 1480 1372 1481
rect 1366 1476 1367 1480
rect 1371 1476 1372 1480
rect 1518 1477 1519 1481
rect 1523 1477 1524 1481
rect 1518 1476 1524 1477
rect 1574 1481 1580 1482
rect 1574 1477 1575 1481
rect 1579 1477 1580 1481
rect 1574 1476 1580 1477
rect 1646 1481 1652 1482
rect 1646 1477 1647 1481
rect 1651 1477 1652 1481
rect 1646 1476 1652 1477
rect 1726 1481 1732 1482
rect 1726 1477 1727 1481
rect 1731 1477 1732 1481
rect 1726 1476 1732 1477
rect 1806 1481 1812 1482
rect 1806 1477 1807 1481
rect 1811 1477 1812 1481
rect 1806 1476 1812 1477
rect 1894 1481 1900 1482
rect 1894 1477 1895 1481
rect 1899 1477 1900 1481
rect 1894 1476 1900 1477
rect 1982 1481 1988 1482
rect 1982 1477 1983 1481
rect 1987 1477 1988 1481
rect 1982 1476 1988 1477
rect 2070 1481 2076 1482
rect 2070 1477 2071 1481
rect 2075 1477 2076 1481
rect 2070 1476 2076 1477
rect 2150 1481 2156 1482
rect 2150 1477 2151 1481
rect 2155 1477 2156 1481
rect 2150 1476 2156 1477
rect 2230 1481 2236 1482
rect 2230 1477 2231 1481
rect 2235 1477 2236 1481
rect 2230 1476 2236 1477
rect 2310 1481 2316 1482
rect 2310 1477 2311 1481
rect 2315 1477 2316 1481
rect 2310 1476 2316 1477
rect 2390 1481 2396 1482
rect 2390 1477 2391 1481
rect 2395 1477 2396 1481
rect 2390 1476 2396 1477
rect 2470 1481 2476 1482
rect 2470 1477 2471 1481
rect 2475 1477 2476 1481
rect 2470 1476 2476 1477
rect 2526 1481 2532 1482
rect 2526 1477 2527 1481
rect 2531 1477 2532 1481
rect 2526 1476 2532 1477
rect 2582 1480 2588 1481
rect 2582 1476 2583 1480
rect 2587 1476 2588 1480
rect 1366 1475 1372 1476
rect 2582 1475 2588 1476
rect 198 1473 204 1474
rect 110 1472 116 1473
rect 110 1468 111 1472
rect 115 1468 116 1472
rect 198 1469 199 1473
rect 203 1469 204 1473
rect 198 1468 204 1469
rect 286 1473 292 1474
rect 286 1469 287 1473
rect 291 1469 292 1473
rect 286 1468 292 1469
rect 382 1473 388 1474
rect 382 1469 383 1473
rect 387 1469 388 1473
rect 382 1468 388 1469
rect 486 1473 492 1474
rect 486 1469 487 1473
rect 491 1469 492 1473
rect 486 1468 492 1469
rect 582 1473 588 1474
rect 582 1469 583 1473
rect 587 1469 588 1473
rect 582 1468 588 1469
rect 678 1473 684 1474
rect 678 1469 679 1473
rect 683 1469 684 1473
rect 678 1468 684 1469
rect 774 1473 780 1474
rect 774 1469 775 1473
rect 779 1469 780 1473
rect 774 1468 780 1469
rect 862 1473 868 1474
rect 862 1469 863 1473
rect 867 1469 868 1473
rect 862 1468 868 1469
rect 950 1473 956 1474
rect 950 1469 951 1473
rect 955 1469 956 1473
rect 950 1468 956 1469
rect 1038 1473 1044 1474
rect 1038 1469 1039 1473
rect 1043 1469 1044 1473
rect 1038 1468 1044 1469
rect 1134 1473 1140 1474
rect 1134 1469 1135 1473
rect 1139 1469 1140 1473
rect 1134 1468 1140 1469
rect 1326 1472 1332 1473
rect 1326 1468 1327 1472
rect 1331 1468 1332 1472
rect 110 1467 116 1468
rect 1326 1467 1332 1468
rect 1366 1463 1372 1464
rect 1366 1459 1367 1463
rect 1371 1459 1372 1463
rect 1366 1458 1372 1459
rect 2582 1463 2588 1464
rect 2582 1459 2583 1463
rect 2587 1459 2588 1463
rect 2582 1458 2588 1459
rect 110 1455 116 1456
rect 110 1451 111 1455
rect 115 1451 116 1455
rect 110 1450 116 1451
rect 1326 1455 1332 1456
rect 1326 1451 1327 1455
rect 1331 1451 1332 1455
rect 1326 1450 1332 1451
rect 1534 1454 1540 1455
rect 1534 1450 1535 1454
rect 1539 1450 1540 1454
rect 1534 1449 1540 1450
rect 1590 1454 1596 1455
rect 1590 1450 1591 1454
rect 1595 1450 1596 1454
rect 1590 1449 1596 1450
rect 1662 1454 1668 1455
rect 1662 1450 1663 1454
rect 1667 1450 1668 1454
rect 1662 1449 1668 1450
rect 1742 1454 1748 1455
rect 1742 1450 1743 1454
rect 1747 1450 1748 1454
rect 1742 1449 1748 1450
rect 1822 1454 1828 1455
rect 1822 1450 1823 1454
rect 1827 1450 1828 1454
rect 1822 1449 1828 1450
rect 1910 1454 1916 1455
rect 1910 1450 1911 1454
rect 1915 1450 1916 1454
rect 1910 1449 1916 1450
rect 1998 1454 2004 1455
rect 1998 1450 1999 1454
rect 2003 1450 2004 1454
rect 1998 1449 2004 1450
rect 2086 1454 2092 1455
rect 2086 1450 2087 1454
rect 2091 1450 2092 1454
rect 2086 1449 2092 1450
rect 2166 1454 2172 1455
rect 2166 1450 2167 1454
rect 2171 1450 2172 1454
rect 2166 1449 2172 1450
rect 2246 1454 2252 1455
rect 2246 1450 2247 1454
rect 2251 1450 2252 1454
rect 2246 1449 2252 1450
rect 2326 1454 2332 1455
rect 2326 1450 2327 1454
rect 2331 1450 2332 1454
rect 2326 1449 2332 1450
rect 2406 1454 2412 1455
rect 2406 1450 2407 1454
rect 2411 1450 2412 1454
rect 2406 1449 2412 1450
rect 2486 1454 2492 1455
rect 2486 1450 2487 1454
rect 2491 1450 2492 1454
rect 2486 1449 2492 1450
rect 2542 1454 2548 1455
rect 2542 1450 2543 1454
rect 2547 1450 2548 1454
rect 2542 1449 2548 1450
rect 214 1446 220 1447
rect 214 1442 215 1446
rect 219 1442 220 1446
rect 214 1441 220 1442
rect 302 1446 308 1447
rect 302 1442 303 1446
rect 307 1442 308 1446
rect 302 1441 308 1442
rect 398 1446 404 1447
rect 398 1442 399 1446
rect 403 1442 404 1446
rect 398 1441 404 1442
rect 502 1446 508 1447
rect 502 1442 503 1446
rect 507 1442 508 1446
rect 502 1441 508 1442
rect 598 1446 604 1447
rect 598 1442 599 1446
rect 603 1442 604 1446
rect 598 1441 604 1442
rect 694 1446 700 1447
rect 694 1442 695 1446
rect 699 1442 700 1446
rect 694 1441 700 1442
rect 790 1446 796 1447
rect 790 1442 791 1446
rect 795 1442 796 1446
rect 790 1441 796 1442
rect 878 1446 884 1447
rect 878 1442 879 1446
rect 883 1442 884 1446
rect 878 1441 884 1442
rect 966 1446 972 1447
rect 966 1442 967 1446
rect 971 1442 972 1446
rect 966 1441 972 1442
rect 1054 1446 1060 1447
rect 1054 1442 1055 1446
rect 1059 1442 1060 1446
rect 1054 1441 1060 1442
rect 1150 1446 1156 1447
rect 1150 1442 1151 1446
rect 1155 1442 1156 1446
rect 1150 1441 1156 1442
rect 1414 1422 1420 1423
rect 158 1418 164 1419
rect 158 1414 159 1418
rect 163 1414 164 1418
rect 158 1413 164 1414
rect 246 1418 252 1419
rect 246 1414 247 1418
rect 251 1414 252 1418
rect 246 1413 252 1414
rect 342 1418 348 1419
rect 342 1414 343 1418
rect 347 1414 348 1418
rect 342 1413 348 1414
rect 446 1418 452 1419
rect 446 1414 447 1418
rect 451 1414 452 1418
rect 446 1413 452 1414
rect 550 1418 556 1419
rect 550 1414 551 1418
rect 555 1414 556 1418
rect 550 1413 556 1414
rect 662 1418 668 1419
rect 662 1414 663 1418
rect 667 1414 668 1418
rect 662 1413 668 1414
rect 766 1418 772 1419
rect 766 1414 767 1418
rect 771 1414 772 1418
rect 766 1413 772 1414
rect 878 1418 884 1419
rect 878 1414 879 1418
rect 883 1414 884 1418
rect 878 1413 884 1414
rect 990 1418 996 1419
rect 990 1414 991 1418
rect 995 1414 996 1418
rect 990 1413 996 1414
rect 1102 1418 1108 1419
rect 1102 1414 1103 1418
rect 1107 1414 1108 1418
rect 1102 1413 1108 1414
rect 1214 1418 1220 1419
rect 1214 1414 1215 1418
rect 1219 1414 1220 1418
rect 1414 1418 1415 1422
rect 1419 1418 1420 1422
rect 1414 1417 1420 1418
rect 1470 1422 1476 1423
rect 1470 1418 1471 1422
rect 1475 1418 1476 1422
rect 1470 1417 1476 1418
rect 1534 1422 1540 1423
rect 1534 1418 1535 1422
rect 1539 1418 1540 1422
rect 1534 1417 1540 1418
rect 1622 1422 1628 1423
rect 1622 1418 1623 1422
rect 1627 1418 1628 1422
rect 1622 1417 1628 1418
rect 1718 1422 1724 1423
rect 1718 1418 1719 1422
rect 1723 1418 1724 1422
rect 1718 1417 1724 1418
rect 1822 1422 1828 1423
rect 1822 1418 1823 1422
rect 1827 1418 1828 1422
rect 1822 1417 1828 1418
rect 1926 1422 1932 1423
rect 1926 1418 1927 1422
rect 1931 1418 1932 1422
rect 1926 1417 1932 1418
rect 2022 1422 2028 1423
rect 2022 1418 2023 1422
rect 2027 1418 2028 1422
rect 2022 1417 2028 1418
rect 2118 1422 2124 1423
rect 2118 1418 2119 1422
rect 2123 1418 2124 1422
rect 2118 1417 2124 1418
rect 2214 1422 2220 1423
rect 2214 1418 2215 1422
rect 2219 1418 2220 1422
rect 2214 1417 2220 1418
rect 2302 1422 2308 1423
rect 2302 1418 2303 1422
rect 2307 1418 2308 1422
rect 2302 1417 2308 1418
rect 2390 1422 2396 1423
rect 2390 1418 2391 1422
rect 2395 1418 2396 1422
rect 2390 1417 2396 1418
rect 2478 1422 2484 1423
rect 2478 1418 2479 1422
rect 2483 1418 2484 1422
rect 2478 1417 2484 1418
rect 2542 1422 2548 1423
rect 2542 1418 2543 1422
rect 2547 1418 2548 1422
rect 2542 1417 2548 1418
rect 1214 1413 1220 1414
rect 1366 1413 1372 1414
rect 110 1409 116 1410
rect 110 1405 111 1409
rect 115 1405 116 1409
rect 110 1404 116 1405
rect 1326 1409 1332 1410
rect 1326 1405 1327 1409
rect 1331 1405 1332 1409
rect 1366 1409 1367 1413
rect 1371 1409 1372 1413
rect 1366 1408 1372 1409
rect 2582 1413 2588 1414
rect 2582 1409 2583 1413
rect 2587 1409 2588 1413
rect 2582 1408 2588 1409
rect 1326 1404 1332 1405
rect 1366 1396 1372 1397
rect 2582 1396 2588 1397
rect 110 1392 116 1393
rect 1326 1392 1332 1393
rect 110 1388 111 1392
rect 115 1388 116 1392
rect 110 1387 116 1388
rect 142 1391 148 1392
rect 142 1387 143 1391
rect 147 1387 148 1391
rect 142 1386 148 1387
rect 230 1391 236 1392
rect 230 1387 231 1391
rect 235 1387 236 1391
rect 230 1386 236 1387
rect 326 1391 332 1392
rect 326 1387 327 1391
rect 331 1387 332 1391
rect 326 1386 332 1387
rect 430 1391 436 1392
rect 430 1387 431 1391
rect 435 1387 436 1391
rect 430 1386 436 1387
rect 534 1391 540 1392
rect 534 1387 535 1391
rect 539 1387 540 1391
rect 534 1386 540 1387
rect 646 1391 652 1392
rect 646 1387 647 1391
rect 651 1387 652 1391
rect 646 1386 652 1387
rect 750 1391 756 1392
rect 750 1387 751 1391
rect 755 1387 756 1391
rect 750 1386 756 1387
rect 862 1391 868 1392
rect 862 1387 863 1391
rect 867 1387 868 1391
rect 862 1386 868 1387
rect 974 1391 980 1392
rect 974 1387 975 1391
rect 979 1387 980 1391
rect 974 1386 980 1387
rect 1086 1391 1092 1392
rect 1086 1387 1087 1391
rect 1091 1387 1092 1391
rect 1086 1386 1092 1387
rect 1198 1391 1204 1392
rect 1198 1387 1199 1391
rect 1203 1387 1204 1391
rect 1326 1388 1327 1392
rect 1331 1388 1332 1392
rect 1366 1392 1367 1396
rect 1371 1392 1372 1396
rect 1366 1391 1372 1392
rect 1398 1395 1404 1396
rect 1398 1391 1399 1395
rect 1403 1391 1404 1395
rect 1398 1390 1404 1391
rect 1454 1395 1460 1396
rect 1454 1391 1455 1395
rect 1459 1391 1460 1395
rect 1454 1390 1460 1391
rect 1518 1395 1524 1396
rect 1518 1391 1519 1395
rect 1523 1391 1524 1395
rect 1518 1390 1524 1391
rect 1606 1395 1612 1396
rect 1606 1391 1607 1395
rect 1611 1391 1612 1395
rect 1606 1390 1612 1391
rect 1702 1395 1708 1396
rect 1702 1391 1703 1395
rect 1707 1391 1708 1395
rect 1702 1390 1708 1391
rect 1806 1395 1812 1396
rect 1806 1391 1807 1395
rect 1811 1391 1812 1395
rect 1806 1390 1812 1391
rect 1910 1395 1916 1396
rect 1910 1391 1911 1395
rect 1915 1391 1916 1395
rect 1910 1390 1916 1391
rect 2006 1395 2012 1396
rect 2006 1391 2007 1395
rect 2011 1391 2012 1395
rect 2006 1390 2012 1391
rect 2102 1395 2108 1396
rect 2102 1391 2103 1395
rect 2107 1391 2108 1395
rect 2102 1390 2108 1391
rect 2198 1395 2204 1396
rect 2198 1391 2199 1395
rect 2203 1391 2204 1395
rect 2198 1390 2204 1391
rect 2286 1395 2292 1396
rect 2286 1391 2287 1395
rect 2291 1391 2292 1395
rect 2286 1390 2292 1391
rect 2374 1395 2380 1396
rect 2374 1391 2375 1395
rect 2379 1391 2380 1395
rect 2374 1390 2380 1391
rect 2462 1395 2468 1396
rect 2462 1391 2463 1395
rect 2467 1391 2468 1395
rect 2462 1390 2468 1391
rect 2526 1395 2532 1396
rect 2526 1391 2527 1395
rect 2531 1391 2532 1395
rect 2582 1392 2583 1396
rect 2587 1392 2588 1396
rect 2582 1391 2588 1392
rect 2526 1390 2532 1391
rect 1326 1387 1332 1388
rect 1198 1386 1204 1387
rect 142 1357 148 1358
rect 110 1356 116 1357
rect 110 1352 111 1356
rect 115 1352 116 1356
rect 142 1353 143 1357
rect 147 1353 148 1357
rect 142 1352 148 1353
rect 206 1357 212 1358
rect 206 1353 207 1357
rect 211 1353 212 1357
rect 206 1352 212 1353
rect 294 1357 300 1358
rect 294 1353 295 1357
rect 299 1353 300 1357
rect 294 1352 300 1353
rect 398 1357 404 1358
rect 398 1353 399 1357
rect 403 1353 404 1357
rect 398 1352 404 1353
rect 510 1357 516 1358
rect 510 1353 511 1357
rect 515 1353 516 1357
rect 510 1352 516 1353
rect 622 1357 628 1358
rect 622 1353 623 1357
rect 627 1353 628 1357
rect 622 1352 628 1353
rect 734 1357 740 1358
rect 734 1353 735 1357
rect 739 1353 740 1357
rect 734 1352 740 1353
rect 846 1357 852 1358
rect 846 1353 847 1357
rect 851 1353 852 1357
rect 846 1352 852 1353
rect 958 1357 964 1358
rect 958 1353 959 1357
rect 963 1353 964 1357
rect 958 1352 964 1353
rect 1070 1357 1076 1358
rect 1070 1353 1071 1357
rect 1075 1353 1076 1357
rect 1070 1352 1076 1353
rect 1182 1357 1188 1358
rect 1182 1353 1183 1357
rect 1187 1353 1188 1357
rect 1182 1352 1188 1353
rect 1270 1357 1276 1358
rect 1270 1353 1271 1357
rect 1275 1353 1276 1357
rect 1270 1352 1276 1353
rect 1326 1356 1332 1357
rect 1326 1352 1327 1356
rect 1331 1352 1332 1356
rect 1398 1353 1404 1354
rect 110 1351 116 1352
rect 1326 1351 1332 1352
rect 1366 1352 1372 1353
rect 1366 1348 1367 1352
rect 1371 1348 1372 1352
rect 1398 1349 1399 1353
rect 1403 1349 1404 1353
rect 1398 1348 1404 1349
rect 1454 1353 1460 1354
rect 1454 1349 1455 1353
rect 1459 1349 1460 1353
rect 1454 1348 1460 1349
rect 1542 1353 1548 1354
rect 1542 1349 1543 1353
rect 1547 1349 1548 1353
rect 1542 1348 1548 1349
rect 1630 1353 1636 1354
rect 1630 1349 1631 1353
rect 1635 1349 1636 1353
rect 1630 1348 1636 1349
rect 1718 1353 1724 1354
rect 1718 1349 1719 1353
rect 1723 1349 1724 1353
rect 1718 1348 1724 1349
rect 1806 1353 1812 1354
rect 1806 1349 1807 1353
rect 1811 1349 1812 1353
rect 1806 1348 1812 1349
rect 1886 1353 1892 1354
rect 1886 1349 1887 1353
rect 1891 1349 1892 1353
rect 1886 1348 1892 1349
rect 1966 1353 1972 1354
rect 1966 1349 1967 1353
rect 1971 1349 1972 1353
rect 1966 1348 1972 1349
rect 2046 1353 2052 1354
rect 2046 1349 2047 1353
rect 2051 1349 2052 1353
rect 2046 1348 2052 1349
rect 2126 1353 2132 1354
rect 2126 1349 2127 1353
rect 2131 1349 2132 1353
rect 2126 1348 2132 1349
rect 2206 1353 2212 1354
rect 2206 1349 2207 1353
rect 2211 1349 2212 1353
rect 2206 1348 2212 1349
rect 2582 1352 2588 1353
rect 2582 1348 2583 1352
rect 2587 1348 2588 1352
rect 1366 1347 1372 1348
rect 2582 1347 2588 1348
rect 110 1339 116 1340
rect 110 1335 111 1339
rect 115 1335 116 1339
rect 110 1334 116 1335
rect 1326 1339 1332 1340
rect 1326 1335 1327 1339
rect 1331 1335 1332 1339
rect 1326 1334 1332 1335
rect 1366 1335 1372 1336
rect 1366 1331 1367 1335
rect 1371 1331 1372 1335
rect 158 1330 164 1331
rect 158 1326 159 1330
rect 163 1326 164 1330
rect 158 1325 164 1326
rect 222 1330 228 1331
rect 222 1326 223 1330
rect 227 1326 228 1330
rect 222 1325 228 1326
rect 310 1330 316 1331
rect 310 1326 311 1330
rect 315 1326 316 1330
rect 310 1325 316 1326
rect 414 1330 420 1331
rect 414 1326 415 1330
rect 419 1326 420 1330
rect 414 1325 420 1326
rect 526 1330 532 1331
rect 526 1326 527 1330
rect 531 1326 532 1330
rect 526 1325 532 1326
rect 638 1330 644 1331
rect 638 1326 639 1330
rect 643 1326 644 1330
rect 638 1325 644 1326
rect 750 1330 756 1331
rect 750 1326 751 1330
rect 755 1326 756 1330
rect 750 1325 756 1326
rect 862 1330 868 1331
rect 862 1326 863 1330
rect 867 1326 868 1330
rect 862 1325 868 1326
rect 974 1330 980 1331
rect 974 1326 975 1330
rect 979 1326 980 1330
rect 974 1325 980 1326
rect 1086 1330 1092 1331
rect 1086 1326 1087 1330
rect 1091 1326 1092 1330
rect 1086 1325 1092 1326
rect 1198 1330 1204 1331
rect 1198 1326 1199 1330
rect 1203 1326 1204 1330
rect 1198 1325 1204 1326
rect 1286 1330 1292 1331
rect 1366 1330 1372 1331
rect 2582 1335 2588 1336
rect 2582 1331 2583 1335
rect 2587 1331 2588 1335
rect 2582 1330 2588 1331
rect 1286 1326 1287 1330
rect 1291 1326 1292 1330
rect 1286 1325 1292 1326
rect 1414 1326 1420 1327
rect 1414 1322 1415 1326
rect 1419 1322 1420 1326
rect 1414 1321 1420 1322
rect 1470 1326 1476 1327
rect 1470 1322 1471 1326
rect 1475 1322 1476 1326
rect 1470 1321 1476 1322
rect 1558 1326 1564 1327
rect 1558 1322 1559 1326
rect 1563 1322 1564 1326
rect 1558 1321 1564 1322
rect 1646 1326 1652 1327
rect 1646 1322 1647 1326
rect 1651 1322 1652 1326
rect 1646 1321 1652 1322
rect 1734 1326 1740 1327
rect 1734 1322 1735 1326
rect 1739 1322 1740 1326
rect 1734 1321 1740 1322
rect 1822 1326 1828 1327
rect 1822 1322 1823 1326
rect 1827 1322 1828 1326
rect 1822 1321 1828 1322
rect 1902 1326 1908 1327
rect 1902 1322 1903 1326
rect 1907 1322 1908 1326
rect 1902 1321 1908 1322
rect 1982 1326 1988 1327
rect 1982 1322 1983 1326
rect 1987 1322 1988 1326
rect 1982 1321 1988 1322
rect 2062 1326 2068 1327
rect 2062 1322 2063 1326
rect 2067 1322 2068 1326
rect 2062 1321 2068 1322
rect 2142 1326 2148 1327
rect 2142 1322 2143 1326
rect 2147 1322 2148 1326
rect 2142 1321 2148 1322
rect 2222 1326 2228 1327
rect 2222 1322 2223 1326
rect 2227 1322 2228 1326
rect 2222 1321 2228 1322
rect 158 1306 164 1307
rect 158 1302 159 1306
rect 163 1302 164 1306
rect 158 1301 164 1302
rect 230 1306 236 1307
rect 230 1302 231 1306
rect 235 1302 236 1306
rect 230 1301 236 1302
rect 326 1306 332 1307
rect 326 1302 327 1306
rect 331 1302 332 1306
rect 326 1301 332 1302
rect 430 1306 436 1307
rect 430 1302 431 1306
rect 435 1302 436 1306
rect 430 1301 436 1302
rect 534 1306 540 1307
rect 534 1302 535 1306
rect 539 1302 540 1306
rect 534 1301 540 1302
rect 630 1306 636 1307
rect 630 1302 631 1306
rect 635 1302 636 1306
rect 630 1301 636 1302
rect 726 1306 732 1307
rect 726 1302 727 1306
rect 731 1302 732 1306
rect 726 1301 732 1302
rect 822 1306 828 1307
rect 822 1302 823 1306
rect 827 1302 828 1306
rect 822 1301 828 1302
rect 910 1306 916 1307
rect 910 1302 911 1306
rect 915 1302 916 1306
rect 910 1301 916 1302
rect 990 1306 996 1307
rect 990 1302 991 1306
rect 995 1302 996 1306
rect 990 1301 996 1302
rect 1070 1306 1076 1307
rect 1070 1302 1071 1306
rect 1075 1302 1076 1306
rect 1070 1301 1076 1302
rect 1150 1306 1156 1307
rect 1150 1302 1151 1306
rect 1155 1302 1156 1306
rect 1150 1301 1156 1302
rect 1230 1306 1236 1307
rect 1230 1302 1231 1306
rect 1235 1302 1236 1306
rect 1230 1301 1236 1302
rect 1286 1306 1292 1307
rect 1286 1302 1287 1306
rect 1291 1302 1292 1306
rect 1286 1301 1292 1302
rect 1670 1298 1676 1299
rect 110 1297 116 1298
rect 110 1293 111 1297
rect 115 1293 116 1297
rect 110 1292 116 1293
rect 1326 1297 1332 1298
rect 1326 1293 1327 1297
rect 1331 1293 1332 1297
rect 1670 1294 1671 1298
rect 1675 1294 1676 1298
rect 1670 1293 1676 1294
rect 1766 1298 1772 1299
rect 1766 1294 1767 1298
rect 1771 1294 1772 1298
rect 1766 1293 1772 1294
rect 1862 1298 1868 1299
rect 1862 1294 1863 1298
rect 1867 1294 1868 1298
rect 1862 1293 1868 1294
rect 1958 1298 1964 1299
rect 1958 1294 1959 1298
rect 1963 1294 1964 1298
rect 1958 1293 1964 1294
rect 2046 1298 2052 1299
rect 2046 1294 2047 1298
rect 2051 1294 2052 1298
rect 2046 1293 2052 1294
rect 2134 1298 2140 1299
rect 2134 1294 2135 1298
rect 2139 1294 2140 1298
rect 2134 1293 2140 1294
rect 2230 1298 2236 1299
rect 2230 1294 2231 1298
rect 2235 1294 2236 1298
rect 2230 1293 2236 1294
rect 1326 1292 1332 1293
rect 1366 1289 1372 1290
rect 1366 1285 1367 1289
rect 1371 1285 1372 1289
rect 1366 1284 1372 1285
rect 2582 1289 2588 1290
rect 2582 1285 2583 1289
rect 2587 1285 2588 1289
rect 2582 1284 2588 1285
rect 110 1280 116 1281
rect 1326 1280 1332 1281
rect 110 1276 111 1280
rect 115 1276 116 1280
rect 110 1275 116 1276
rect 142 1279 148 1280
rect 142 1275 143 1279
rect 147 1275 148 1279
rect 142 1274 148 1275
rect 214 1279 220 1280
rect 214 1275 215 1279
rect 219 1275 220 1279
rect 214 1274 220 1275
rect 310 1279 316 1280
rect 310 1275 311 1279
rect 315 1275 316 1279
rect 310 1274 316 1275
rect 414 1279 420 1280
rect 414 1275 415 1279
rect 419 1275 420 1279
rect 414 1274 420 1275
rect 518 1279 524 1280
rect 518 1275 519 1279
rect 523 1275 524 1279
rect 518 1274 524 1275
rect 614 1279 620 1280
rect 614 1275 615 1279
rect 619 1275 620 1279
rect 614 1274 620 1275
rect 710 1279 716 1280
rect 710 1275 711 1279
rect 715 1275 716 1279
rect 710 1274 716 1275
rect 806 1279 812 1280
rect 806 1275 807 1279
rect 811 1275 812 1279
rect 806 1274 812 1275
rect 894 1279 900 1280
rect 894 1275 895 1279
rect 899 1275 900 1279
rect 894 1274 900 1275
rect 974 1279 980 1280
rect 974 1275 975 1279
rect 979 1275 980 1279
rect 974 1274 980 1275
rect 1054 1279 1060 1280
rect 1054 1275 1055 1279
rect 1059 1275 1060 1279
rect 1054 1274 1060 1275
rect 1134 1279 1140 1280
rect 1134 1275 1135 1279
rect 1139 1275 1140 1279
rect 1134 1274 1140 1275
rect 1214 1279 1220 1280
rect 1214 1275 1215 1279
rect 1219 1275 1220 1279
rect 1214 1274 1220 1275
rect 1270 1279 1276 1280
rect 1270 1275 1271 1279
rect 1275 1275 1276 1279
rect 1326 1276 1327 1280
rect 1331 1276 1332 1280
rect 1326 1275 1332 1276
rect 1270 1274 1276 1275
rect 1366 1272 1372 1273
rect 2582 1272 2588 1273
rect 1366 1268 1367 1272
rect 1371 1268 1372 1272
rect 1366 1267 1372 1268
rect 1654 1271 1660 1272
rect 1654 1267 1655 1271
rect 1659 1267 1660 1271
rect 1654 1266 1660 1267
rect 1750 1271 1756 1272
rect 1750 1267 1751 1271
rect 1755 1267 1756 1271
rect 1750 1266 1756 1267
rect 1846 1271 1852 1272
rect 1846 1267 1847 1271
rect 1851 1267 1852 1271
rect 1846 1266 1852 1267
rect 1942 1271 1948 1272
rect 1942 1267 1943 1271
rect 1947 1267 1948 1271
rect 1942 1266 1948 1267
rect 2030 1271 2036 1272
rect 2030 1267 2031 1271
rect 2035 1267 2036 1271
rect 2030 1266 2036 1267
rect 2118 1271 2124 1272
rect 2118 1267 2119 1271
rect 2123 1267 2124 1271
rect 2118 1266 2124 1267
rect 2214 1271 2220 1272
rect 2214 1267 2215 1271
rect 2219 1267 2220 1271
rect 2582 1268 2583 1272
rect 2587 1268 2588 1272
rect 2582 1267 2588 1268
rect 2214 1266 2220 1267
rect 1494 1237 1500 1238
rect 1366 1236 1372 1237
rect 142 1233 148 1234
rect 110 1232 116 1233
rect 110 1228 111 1232
rect 115 1228 116 1232
rect 142 1229 143 1233
rect 147 1229 148 1233
rect 142 1228 148 1229
rect 198 1233 204 1234
rect 198 1229 199 1233
rect 203 1229 204 1233
rect 198 1228 204 1229
rect 278 1233 284 1234
rect 278 1229 279 1233
rect 283 1229 284 1233
rect 278 1228 284 1229
rect 358 1233 364 1234
rect 358 1229 359 1233
rect 363 1229 364 1233
rect 358 1228 364 1229
rect 438 1233 444 1234
rect 438 1229 439 1233
rect 443 1229 444 1233
rect 438 1228 444 1229
rect 518 1233 524 1234
rect 518 1229 519 1233
rect 523 1229 524 1233
rect 518 1228 524 1229
rect 598 1233 604 1234
rect 598 1229 599 1233
rect 603 1229 604 1233
rect 598 1228 604 1229
rect 670 1233 676 1234
rect 670 1229 671 1233
rect 675 1229 676 1233
rect 670 1228 676 1229
rect 742 1233 748 1234
rect 742 1229 743 1233
rect 747 1229 748 1233
rect 742 1228 748 1229
rect 814 1233 820 1234
rect 814 1229 815 1233
rect 819 1229 820 1233
rect 814 1228 820 1229
rect 894 1233 900 1234
rect 894 1229 895 1233
rect 899 1229 900 1233
rect 894 1228 900 1229
rect 1326 1232 1332 1233
rect 1326 1228 1327 1232
rect 1331 1228 1332 1232
rect 1366 1232 1367 1236
rect 1371 1232 1372 1236
rect 1494 1233 1495 1237
rect 1499 1233 1500 1237
rect 1494 1232 1500 1233
rect 1558 1237 1564 1238
rect 1558 1233 1559 1237
rect 1563 1233 1564 1237
rect 1558 1232 1564 1233
rect 1622 1237 1628 1238
rect 1622 1233 1623 1237
rect 1627 1233 1628 1237
rect 1622 1232 1628 1233
rect 1686 1237 1692 1238
rect 1686 1233 1687 1237
rect 1691 1233 1692 1237
rect 1686 1232 1692 1233
rect 1758 1237 1764 1238
rect 1758 1233 1759 1237
rect 1763 1233 1764 1237
rect 1758 1232 1764 1233
rect 1822 1237 1828 1238
rect 1822 1233 1823 1237
rect 1827 1233 1828 1237
rect 1822 1232 1828 1233
rect 1886 1237 1892 1238
rect 1886 1233 1887 1237
rect 1891 1233 1892 1237
rect 1886 1232 1892 1233
rect 1950 1237 1956 1238
rect 1950 1233 1951 1237
rect 1955 1233 1956 1237
rect 1950 1232 1956 1233
rect 2014 1237 2020 1238
rect 2014 1233 2015 1237
rect 2019 1233 2020 1237
rect 2014 1232 2020 1233
rect 2078 1237 2084 1238
rect 2078 1233 2079 1237
rect 2083 1233 2084 1237
rect 2078 1232 2084 1233
rect 2150 1237 2156 1238
rect 2150 1233 2151 1237
rect 2155 1233 2156 1237
rect 2150 1232 2156 1233
rect 2222 1237 2228 1238
rect 2222 1233 2223 1237
rect 2227 1233 2228 1237
rect 2222 1232 2228 1233
rect 2294 1237 2300 1238
rect 2294 1233 2295 1237
rect 2299 1233 2300 1237
rect 2294 1232 2300 1233
rect 2582 1236 2588 1237
rect 2582 1232 2583 1236
rect 2587 1232 2588 1236
rect 1366 1231 1372 1232
rect 2582 1231 2588 1232
rect 110 1227 116 1228
rect 1326 1227 1332 1228
rect 1366 1219 1372 1220
rect 110 1215 116 1216
rect 110 1211 111 1215
rect 115 1211 116 1215
rect 110 1210 116 1211
rect 1326 1215 1332 1216
rect 1326 1211 1327 1215
rect 1331 1211 1332 1215
rect 1366 1215 1367 1219
rect 1371 1215 1372 1219
rect 1366 1214 1372 1215
rect 2582 1219 2588 1220
rect 2582 1215 2583 1219
rect 2587 1215 2588 1219
rect 2582 1214 2588 1215
rect 1326 1210 1332 1211
rect 1510 1210 1516 1211
rect 158 1206 164 1207
rect 158 1202 159 1206
rect 163 1202 164 1206
rect 158 1201 164 1202
rect 214 1206 220 1207
rect 214 1202 215 1206
rect 219 1202 220 1206
rect 214 1201 220 1202
rect 294 1206 300 1207
rect 294 1202 295 1206
rect 299 1202 300 1206
rect 294 1201 300 1202
rect 374 1206 380 1207
rect 374 1202 375 1206
rect 379 1202 380 1206
rect 374 1201 380 1202
rect 454 1206 460 1207
rect 454 1202 455 1206
rect 459 1202 460 1206
rect 454 1201 460 1202
rect 534 1206 540 1207
rect 534 1202 535 1206
rect 539 1202 540 1206
rect 534 1201 540 1202
rect 614 1206 620 1207
rect 614 1202 615 1206
rect 619 1202 620 1206
rect 614 1201 620 1202
rect 686 1206 692 1207
rect 686 1202 687 1206
rect 691 1202 692 1206
rect 686 1201 692 1202
rect 758 1206 764 1207
rect 758 1202 759 1206
rect 763 1202 764 1206
rect 758 1201 764 1202
rect 830 1206 836 1207
rect 830 1202 831 1206
rect 835 1202 836 1206
rect 830 1201 836 1202
rect 910 1206 916 1207
rect 910 1202 911 1206
rect 915 1202 916 1206
rect 1510 1206 1511 1210
rect 1515 1206 1516 1210
rect 1510 1205 1516 1206
rect 1574 1210 1580 1211
rect 1574 1206 1575 1210
rect 1579 1206 1580 1210
rect 1574 1205 1580 1206
rect 1638 1210 1644 1211
rect 1638 1206 1639 1210
rect 1643 1206 1644 1210
rect 1638 1205 1644 1206
rect 1702 1210 1708 1211
rect 1702 1206 1703 1210
rect 1707 1206 1708 1210
rect 1702 1205 1708 1206
rect 1774 1210 1780 1211
rect 1774 1206 1775 1210
rect 1779 1206 1780 1210
rect 1774 1205 1780 1206
rect 1838 1210 1844 1211
rect 1838 1206 1839 1210
rect 1843 1206 1844 1210
rect 1838 1205 1844 1206
rect 1902 1210 1908 1211
rect 1902 1206 1903 1210
rect 1907 1206 1908 1210
rect 1902 1205 1908 1206
rect 1966 1210 1972 1211
rect 1966 1206 1967 1210
rect 1971 1206 1972 1210
rect 1966 1205 1972 1206
rect 2030 1210 2036 1211
rect 2030 1206 2031 1210
rect 2035 1206 2036 1210
rect 2030 1205 2036 1206
rect 2094 1210 2100 1211
rect 2094 1206 2095 1210
rect 2099 1206 2100 1210
rect 2094 1205 2100 1206
rect 2166 1210 2172 1211
rect 2166 1206 2167 1210
rect 2171 1206 2172 1210
rect 2166 1205 2172 1206
rect 2238 1210 2244 1211
rect 2238 1206 2239 1210
rect 2243 1206 2244 1210
rect 2238 1205 2244 1206
rect 2310 1210 2316 1211
rect 2310 1206 2311 1210
rect 2315 1206 2316 1210
rect 2310 1205 2316 1206
rect 910 1201 916 1202
rect 158 1178 164 1179
rect 158 1174 159 1178
rect 163 1174 164 1178
rect 158 1173 164 1174
rect 238 1178 244 1179
rect 238 1174 239 1178
rect 243 1174 244 1178
rect 238 1173 244 1174
rect 326 1178 332 1179
rect 326 1174 327 1178
rect 331 1174 332 1178
rect 326 1173 332 1174
rect 422 1178 428 1179
rect 422 1174 423 1178
rect 427 1174 428 1178
rect 422 1173 428 1174
rect 510 1178 516 1179
rect 510 1174 511 1178
rect 515 1174 516 1178
rect 510 1173 516 1174
rect 598 1178 604 1179
rect 598 1174 599 1178
rect 603 1174 604 1178
rect 598 1173 604 1174
rect 686 1178 692 1179
rect 686 1174 687 1178
rect 691 1174 692 1178
rect 686 1173 692 1174
rect 766 1178 772 1179
rect 766 1174 767 1178
rect 771 1174 772 1178
rect 766 1173 772 1174
rect 838 1178 844 1179
rect 838 1174 839 1178
rect 843 1174 844 1178
rect 838 1173 844 1174
rect 910 1178 916 1179
rect 910 1174 911 1178
rect 915 1174 916 1178
rect 910 1173 916 1174
rect 982 1178 988 1179
rect 982 1174 983 1178
rect 987 1174 988 1178
rect 982 1173 988 1174
rect 1062 1178 1068 1179
rect 1062 1174 1063 1178
rect 1067 1174 1068 1178
rect 1062 1173 1068 1174
rect 1414 1178 1420 1179
rect 1414 1174 1415 1178
rect 1419 1174 1420 1178
rect 1414 1173 1420 1174
rect 1502 1178 1508 1179
rect 1502 1174 1503 1178
rect 1507 1174 1508 1178
rect 1502 1173 1508 1174
rect 1598 1178 1604 1179
rect 1598 1174 1599 1178
rect 1603 1174 1604 1178
rect 1598 1173 1604 1174
rect 1702 1178 1708 1179
rect 1702 1174 1703 1178
rect 1707 1174 1708 1178
rect 1702 1173 1708 1174
rect 1806 1178 1812 1179
rect 1806 1174 1807 1178
rect 1811 1174 1812 1178
rect 1806 1173 1812 1174
rect 1910 1178 1916 1179
rect 1910 1174 1911 1178
rect 1915 1174 1916 1178
rect 1910 1173 1916 1174
rect 2014 1178 2020 1179
rect 2014 1174 2015 1178
rect 2019 1174 2020 1178
rect 2014 1173 2020 1174
rect 2110 1178 2116 1179
rect 2110 1174 2111 1178
rect 2115 1174 2116 1178
rect 2110 1173 2116 1174
rect 2206 1178 2212 1179
rect 2206 1174 2207 1178
rect 2211 1174 2212 1178
rect 2206 1173 2212 1174
rect 2302 1178 2308 1179
rect 2302 1174 2303 1178
rect 2307 1174 2308 1178
rect 2302 1173 2308 1174
rect 2398 1178 2404 1179
rect 2398 1174 2399 1178
rect 2403 1174 2404 1178
rect 2398 1173 2404 1174
rect 110 1169 116 1170
rect 110 1165 111 1169
rect 115 1165 116 1169
rect 110 1164 116 1165
rect 1326 1169 1332 1170
rect 1326 1165 1327 1169
rect 1331 1165 1332 1169
rect 1326 1164 1332 1165
rect 1366 1169 1372 1170
rect 1366 1165 1367 1169
rect 1371 1165 1372 1169
rect 1366 1164 1372 1165
rect 2582 1169 2588 1170
rect 2582 1165 2583 1169
rect 2587 1165 2588 1169
rect 2582 1164 2588 1165
rect 110 1152 116 1153
rect 1326 1152 1332 1153
rect 110 1148 111 1152
rect 115 1148 116 1152
rect 110 1147 116 1148
rect 142 1151 148 1152
rect 142 1147 143 1151
rect 147 1147 148 1151
rect 142 1146 148 1147
rect 222 1151 228 1152
rect 222 1147 223 1151
rect 227 1147 228 1151
rect 222 1146 228 1147
rect 310 1151 316 1152
rect 310 1147 311 1151
rect 315 1147 316 1151
rect 310 1146 316 1147
rect 406 1151 412 1152
rect 406 1147 407 1151
rect 411 1147 412 1151
rect 406 1146 412 1147
rect 494 1151 500 1152
rect 494 1147 495 1151
rect 499 1147 500 1151
rect 494 1146 500 1147
rect 582 1151 588 1152
rect 582 1147 583 1151
rect 587 1147 588 1151
rect 582 1146 588 1147
rect 670 1151 676 1152
rect 670 1147 671 1151
rect 675 1147 676 1151
rect 670 1146 676 1147
rect 750 1151 756 1152
rect 750 1147 751 1151
rect 755 1147 756 1151
rect 750 1146 756 1147
rect 822 1151 828 1152
rect 822 1147 823 1151
rect 827 1147 828 1151
rect 822 1146 828 1147
rect 894 1151 900 1152
rect 894 1147 895 1151
rect 899 1147 900 1151
rect 894 1146 900 1147
rect 966 1151 972 1152
rect 966 1147 967 1151
rect 971 1147 972 1151
rect 966 1146 972 1147
rect 1046 1151 1052 1152
rect 1046 1147 1047 1151
rect 1051 1147 1052 1151
rect 1326 1148 1327 1152
rect 1331 1148 1332 1152
rect 1326 1147 1332 1148
rect 1366 1152 1372 1153
rect 2582 1152 2588 1153
rect 1366 1148 1367 1152
rect 1371 1148 1372 1152
rect 1366 1147 1372 1148
rect 1398 1151 1404 1152
rect 1398 1147 1399 1151
rect 1403 1147 1404 1151
rect 1046 1146 1052 1147
rect 1398 1146 1404 1147
rect 1486 1151 1492 1152
rect 1486 1147 1487 1151
rect 1491 1147 1492 1151
rect 1486 1146 1492 1147
rect 1582 1151 1588 1152
rect 1582 1147 1583 1151
rect 1587 1147 1588 1151
rect 1582 1146 1588 1147
rect 1686 1151 1692 1152
rect 1686 1147 1687 1151
rect 1691 1147 1692 1151
rect 1686 1146 1692 1147
rect 1790 1151 1796 1152
rect 1790 1147 1791 1151
rect 1795 1147 1796 1151
rect 1790 1146 1796 1147
rect 1894 1151 1900 1152
rect 1894 1147 1895 1151
rect 1899 1147 1900 1151
rect 1894 1146 1900 1147
rect 1998 1151 2004 1152
rect 1998 1147 1999 1151
rect 2003 1147 2004 1151
rect 1998 1146 2004 1147
rect 2094 1151 2100 1152
rect 2094 1147 2095 1151
rect 2099 1147 2100 1151
rect 2094 1146 2100 1147
rect 2190 1151 2196 1152
rect 2190 1147 2191 1151
rect 2195 1147 2196 1151
rect 2190 1146 2196 1147
rect 2286 1151 2292 1152
rect 2286 1147 2287 1151
rect 2291 1147 2292 1151
rect 2286 1146 2292 1147
rect 2382 1151 2388 1152
rect 2382 1147 2383 1151
rect 2387 1147 2388 1151
rect 2582 1148 2583 1152
rect 2587 1148 2588 1152
rect 2582 1147 2588 1148
rect 2382 1146 2388 1147
rect 1398 1113 1404 1114
rect 1366 1112 1372 1113
rect 222 1109 228 1110
rect 110 1108 116 1109
rect 110 1104 111 1108
rect 115 1104 116 1108
rect 222 1105 223 1109
rect 227 1105 228 1109
rect 222 1104 228 1105
rect 318 1109 324 1110
rect 318 1105 319 1109
rect 323 1105 324 1109
rect 318 1104 324 1105
rect 422 1109 428 1110
rect 422 1105 423 1109
rect 427 1105 428 1109
rect 422 1104 428 1105
rect 526 1109 532 1110
rect 526 1105 527 1109
rect 531 1105 532 1109
rect 526 1104 532 1105
rect 630 1109 636 1110
rect 630 1105 631 1109
rect 635 1105 636 1109
rect 630 1104 636 1105
rect 726 1109 732 1110
rect 726 1105 727 1109
rect 731 1105 732 1109
rect 726 1104 732 1105
rect 822 1109 828 1110
rect 822 1105 823 1109
rect 827 1105 828 1109
rect 822 1104 828 1105
rect 910 1109 916 1110
rect 910 1105 911 1109
rect 915 1105 916 1109
rect 910 1104 916 1105
rect 990 1109 996 1110
rect 990 1105 991 1109
rect 995 1105 996 1109
rect 990 1104 996 1105
rect 1078 1109 1084 1110
rect 1078 1105 1079 1109
rect 1083 1105 1084 1109
rect 1078 1104 1084 1105
rect 1166 1109 1172 1110
rect 1166 1105 1167 1109
rect 1171 1105 1172 1109
rect 1166 1104 1172 1105
rect 1326 1108 1332 1109
rect 1326 1104 1327 1108
rect 1331 1104 1332 1108
rect 1366 1108 1367 1112
rect 1371 1108 1372 1112
rect 1398 1109 1399 1113
rect 1403 1109 1404 1113
rect 1398 1108 1404 1109
rect 1478 1113 1484 1114
rect 1478 1109 1479 1113
rect 1483 1109 1484 1113
rect 1478 1108 1484 1109
rect 1582 1113 1588 1114
rect 1582 1109 1583 1113
rect 1587 1109 1588 1113
rect 1582 1108 1588 1109
rect 1686 1113 1692 1114
rect 1686 1109 1687 1113
rect 1691 1109 1692 1113
rect 1686 1108 1692 1109
rect 1790 1113 1796 1114
rect 1790 1109 1791 1113
rect 1795 1109 1796 1113
rect 1790 1108 1796 1109
rect 1886 1113 1892 1114
rect 1886 1109 1887 1113
rect 1891 1109 1892 1113
rect 1886 1108 1892 1109
rect 1974 1113 1980 1114
rect 1974 1109 1975 1113
rect 1979 1109 1980 1113
rect 1974 1108 1980 1109
rect 2062 1113 2068 1114
rect 2062 1109 2063 1113
rect 2067 1109 2068 1113
rect 2062 1108 2068 1109
rect 2142 1113 2148 1114
rect 2142 1109 2143 1113
rect 2147 1109 2148 1113
rect 2142 1108 2148 1109
rect 2214 1113 2220 1114
rect 2214 1109 2215 1113
rect 2219 1109 2220 1113
rect 2214 1108 2220 1109
rect 2278 1113 2284 1114
rect 2278 1109 2279 1113
rect 2283 1109 2284 1113
rect 2278 1108 2284 1109
rect 2342 1113 2348 1114
rect 2342 1109 2343 1113
rect 2347 1109 2348 1113
rect 2342 1108 2348 1109
rect 2406 1113 2412 1114
rect 2406 1109 2407 1113
rect 2411 1109 2412 1113
rect 2406 1108 2412 1109
rect 2470 1113 2476 1114
rect 2470 1109 2471 1113
rect 2475 1109 2476 1113
rect 2470 1108 2476 1109
rect 2526 1113 2532 1114
rect 2526 1109 2527 1113
rect 2531 1109 2532 1113
rect 2526 1108 2532 1109
rect 2582 1112 2588 1113
rect 2582 1108 2583 1112
rect 2587 1108 2588 1112
rect 1366 1107 1372 1108
rect 2582 1107 2588 1108
rect 110 1103 116 1104
rect 1326 1103 1332 1104
rect 1366 1095 1372 1096
rect 110 1091 116 1092
rect 110 1087 111 1091
rect 115 1087 116 1091
rect 110 1086 116 1087
rect 1326 1091 1332 1092
rect 1326 1087 1327 1091
rect 1331 1087 1332 1091
rect 1366 1091 1367 1095
rect 1371 1091 1372 1095
rect 1366 1090 1372 1091
rect 2582 1095 2588 1096
rect 2582 1091 2583 1095
rect 2587 1091 2588 1095
rect 2582 1090 2588 1091
rect 1326 1086 1332 1087
rect 1414 1086 1420 1087
rect 238 1082 244 1083
rect 238 1078 239 1082
rect 243 1078 244 1082
rect 238 1077 244 1078
rect 334 1082 340 1083
rect 334 1078 335 1082
rect 339 1078 340 1082
rect 334 1077 340 1078
rect 438 1082 444 1083
rect 438 1078 439 1082
rect 443 1078 444 1082
rect 438 1077 444 1078
rect 542 1082 548 1083
rect 542 1078 543 1082
rect 547 1078 548 1082
rect 542 1077 548 1078
rect 646 1082 652 1083
rect 646 1078 647 1082
rect 651 1078 652 1082
rect 646 1077 652 1078
rect 742 1082 748 1083
rect 742 1078 743 1082
rect 747 1078 748 1082
rect 742 1077 748 1078
rect 838 1082 844 1083
rect 838 1078 839 1082
rect 843 1078 844 1082
rect 838 1077 844 1078
rect 926 1082 932 1083
rect 926 1078 927 1082
rect 931 1078 932 1082
rect 926 1077 932 1078
rect 1006 1082 1012 1083
rect 1006 1078 1007 1082
rect 1011 1078 1012 1082
rect 1006 1077 1012 1078
rect 1094 1082 1100 1083
rect 1094 1078 1095 1082
rect 1099 1078 1100 1082
rect 1094 1077 1100 1078
rect 1182 1082 1188 1083
rect 1182 1078 1183 1082
rect 1187 1078 1188 1082
rect 1414 1082 1415 1086
rect 1419 1082 1420 1086
rect 1414 1081 1420 1082
rect 1494 1086 1500 1087
rect 1494 1082 1495 1086
rect 1499 1082 1500 1086
rect 1494 1081 1500 1082
rect 1598 1086 1604 1087
rect 1598 1082 1599 1086
rect 1603 1082 1604 1086
rect 1598 1081 1604 1082
rect 1702 1086 1708 1087
rect 1702 1082 1703 1086
rect 1707 1082 1708 1086
rect 1702 1081 1708 1082
rect 1806 1086 1812 1087
rect 1806 1082 1807 1086
rect 1811 1082 1812 1086
rect 1806 1081 1812 1082
rect 1902 1086 1908 1087
rect 1902 1082 1903 1086
rect 1907 1082 1908 1086
rect 1902 1081 1908 1082
rect 1990 1086 1996 1087
rect 1990 1082 1991 1086
rect 1995 1082 1996 1086
rect 1990 1081 1996 1082
rect 2078 1086 2084 1087
rect 2078 1082 2079 1086
rect 2083 1082 2084 1086
rect 2078 1081 2084 1082
rect 2158 1086 2164 1087
rect 2158 1082 2159 1086
rect 2163 1082 2164 1086
rect 2158 1081 2164 1082
rect 2230 1086 2236 1087
rect 2230 1082 2231 1086
rect 2235 1082 2236 1086
rect 2230 1081 2236 1082
rect 2294 1086 2300 1087
rect 2294 1082 2295 1086
rect 2299 1082 2300 1086
rect 2294 1081 2300 1082
rect 2358 1086 2364 1087
rect 2358 1082 2359 1086
rect 2363 1082 2364 1086
rect 2358 1081 2364 1082
rect 2422 1086 2428 1087
rect 2422 1082 2423 1086
rect 2427 1082 2428 1086
rect 2422 1081 2428 1082
rect 2486 1086 2492 1087
rect 2486 1082 2487 1086
rect 2491 1082 2492 1086
rect 2486 1081 2492 1082
rect 2542 1086 2548 1087
rect 2542 1082 2543 1086
rect 2547 1082 2548 1086
rect 2542 1081 2548 1082
rect 1182 1077 1188 1078
rect 1414 1058 1420 1059
rect 310 1054 316 1055
rect 310 1050 311 1054
rect 315 1050 316 1054
rect 310 1049 316 1050
rect 366 1054 372 1055
rect 366 1050 367 1054
rect 371 1050 372 1054
rect 366 1049 372 1050
rect 438 1054 444 1055
rect 438 1050 439 1054
rect 443 1050 444 1054
rect 438 1049 444 1050
rect 518 1054 524 1055
rect 518 1050 519 1054
rect 523 1050 524 1054
rect 518 1049 524 1050
rect 606 1054 612 1055
rect 606 1050 607 1054
rect 611 1050 612 1054
rect 606 1049 612 1050
rect 702 1054 708 1055
rect 702 1050 703 1054
rect 707 1050 708 1054
rect 702 1049 708 1050
rect 798 1054 804 1055
rect 798 1050 799 1054
rect 803 1050 804 1054
rect 798 1049 804 1050
rect 886 1054 892 1055
rect 886 1050 887 1054
rect 891 1050 892 1054
rect 886 1049 892 1050
rect 974 1054 980 1055
rect 974 1050 975 1054
rect 979 1050 980 1054
rect 974 1049 980 1050
rect 1054 1054 1060 1055
rect 1054 1050 1055 1054
rect 1059 1050 1060 1054
rect 1054 1049 1060 1050
rect 1134 1054 1140 1055
rect 1134 1050 1135 1054
rect 1139 1050 1140 1054
rect 1134 1049 1140 1050
rect 1222 1054 1228 1055
rect 1222 1050 1223 1054
rect 1227 1050 1228 1054
rect 1222 1049 1228 1050
rect 1286 1054 1292 1055
rect 1286 1050 1287 1054
rect 1291 1050 1292 1054
rect 1414 1054 1415 1058
rect 1419 1054 1420 1058
rect 1414 1053 1420 1054
rect 1470 1058 1476 1059
rect 1470 1054 1471 1058
rect 1475 1054 1476 1058
rect 1470 1053 1476 1054
rect 1534 1058 1540 1059
rect 1534 1054 1535 1058
rect 1539 1054 1540 1058
rect 1534 1053 1540 1054
rect 1622 1058 1628 1059
rect 1622 1054 1623 1058
rect 1627 1054 1628 1058
rect 1622 1053 1628 1054
rect 1726 1058 1732 1059
rect 1726 1054 1727 1058
rect 1731 1054 1732 1058
rect 1726 1053 1732 1054
rect 1838 1058 1844 1059
rect 1838 1054 1839 1058
rect 1843 1054 1844 1058
rect 1838 1053 1844 1054
rect 1950 1058 1956 1059
rect 1950 1054 1951 1058
rect 1955 1054 1956 1058
rect 1950 1053 1956 1054
rect 2062 1058 2068 1059
rect 2062 1054 2063 1058
rect 2067 1054 2068 1058
rect 2062 1053 2068 1054
rect 2166 1058 2172 1059
rect 2166 1054 2167 1058
rect 2171 1054 2172 1058
rect 2166 1053 2172 1054
rect 2270 1058 2276 1059
rect 2270 1054 2271 1058
rect 2275 1054 2276 1058
rect 2270 1053 2276 1054
rect 2366 1058 2372 1059
rect 2366 1054 2367 1058
rect 2371 1054 2372 1058
rect 2366 1053 2372 1054
rect 2462 1058 2468 1059
rect 2462 1054 2463 1058
rect 2467 1054 2468 1058
rect 2462 1053 2468 1054
rect 2542 1058 2548 1059
rect 2542 1054 2543 1058
rect 2547 1054 2548 1058
rect 2542 1053 2548 1054
rect 1286 1049 1292 1050
rect 1366 1049 1372 1050
rect 110 1045 116 1046
rect 110 1041 111 1045
rect 115 1041 116 1045
rect 110 1040 116 1041
rect 1326 1045 1332 1046
rect 1326 1041 1327 1045
rect 1331 1041 1332 1045
rect 1366 1045 1367 1049
rect 1371 1045 1372 1049
rect 1366 1044 1372 1045
rect 2582 1049 2588 1050
rect 2582 1045 2583 1049
rect 2587 1045 2588 1049
rect 2582 1044 2588 1045
rect 1326 1040 1332 1041
rect 1366 1032 1372 1033
rect 2582 1032 2588 1033
rect 110 1028 116 1029
rect 1326 1028 1332 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 110 1023 116 1024
rect 294 1027 300 1028
rect 294 1023 295 1027
rect 299 1023 300 1027
rect 294 1022 300 1023
rect 350 1027 356 1028
rect 350 1023 351 1027
rect 355 1023 356 1027
rect 350 1022 356 1023
rect 422 1027 428 1028
rect 422 1023 423 1027
rect 427 1023 428 1027
rect 422 1022 428 1023
rect 502 1027 508 1028
rect 502 1023 503 1027
rect 507 1023 508 1027
rect 502 1022 508 1023
rect 590 1027 596 1028
rect 590 1023 591 1027
rect 595 1023 596 1027
rect 590 1022 596 1023
rect 686 1027 692 1028
rect 686 1023 687 1027
rect 691 1023 692 1027
rect 686 1022 692 1023
rect 782 1027 788 1028
rect 782 1023 783 1027
rect 787 1023 788 1027
rect 782 1022 788 1023
rect 870 1027 876 1028
rect 870 1023 871 1027
rect 875 1023 876 1027
rect 870 1022 876 1023
rect 958 1027 964 1028
rect 958 1023 959 1027
rect 963 1023 964 1027
rect 958 1022 964 1023
rect 1038 1027 1044 1028
rect 1038 1023 1039 1027
rect 1043 1023 1044 1027
rect 1038 1022 1044 1023
rect 1118 1027 1124 1028
rect 1118 1023 1119 1027
rect 1123 1023 1124 1027
rect 1118 1022 1124 1023
rect 1206 1027 1212 1028
rect 1206 1023 1207 1027
rect 1211 1023 1212 1027
rect 1206 1022 1212 1023
rect 1270 1027 1276 1028
rect 1270 1023 1271 1027
rect 1275 1023 1276 1027
rect 1326 1024 1327 1028
rect 1331 1024 1332 1028
rect 1366 1028 1367 1032
rect 1371 1028 1372 1032
rect 1366 1027 1372 1028
rect 1398 1031 1404 1032
rect 1398 1027 1399 1031
rect 1403 1027 1404 1031
rect 1398 1026 1404 1027
rect 1454 1031 1460 1032
rect 1454 1027 1455 1031
rect 1459 1027 1460 1031
rect 1454 1026 1460 1027
rect 1518 1031 1524 1032
rect 1518 1027 1519 1031
rect 1523 1027 1524 1031
rect 1518 1026 1524 1027
rect 1606 1031 1612 1032
rect 1606 1027 1607 1031
rect 1611 1027 1612 1031
rect 1606 1026 1612 1027
rect 1710 1031 1716 1032
rect 1710 1027 1711 1031
rect 1715 1027 1716 1031
rect 1710 1026 1716 1027
rect 1822 1031 1828 1032
rect 1822 1027 1823 1031
rect 1827 1027 1828 1031
rect 1822 1026 1828 1027
rect 1934 1031 1940 1032
rect 1934 1027 1935 1031
rect 1939 1027 1940 1031
rect 1934 1026 1940 1027
rect 2046 1031 2052 1032
rect 2046 1027 2047 1031
rect 2051 1027 2052 1031
rect 2046 1026 2052 1027
rect 2150 1031 2156 1032
rect 2150 1027 2151 1031
rect 2155 1027 2156 1031
rect 2150 1026 2156 1027
rect 2254 1031 2260 1032
rect 2254 1027 2255 1031
rect 2259 1027 2260 1031
rect 2254 1026 2260 1027
rect 2350 1031 2356 1032
rect 2350 1027 2351 1031
rect 2355 1027 2356 1031
rect 2350 1026 2356 1027
rect 2446 1031 2452 1032
rect 2446 1027 2447 1031
rect 2451 1027 2452 1031
rect 2446 1026 2452 1027
rect 2526 1031 2532 1032
rect 2526 1027 2527 1031
rect 2531 1027 2532 1031
rect 2582 1028 2583 1032
rect 2587 1028 2588 1032
rect 2582 1027 2588 1028
rect 2526 1026 2532 1027
rect 1326 1023 1332 1024
rect 1270 1022 1276 1023
rect 414 989 420 990
rect 110 988 116 989
rect 110 984 111 988
rect 115 984 116 988
rect 414 985 415 989
rect 419 985 420 989
rect 414 984 420 985
rect 470 989 476 990
rect 470 985 471 989
rect 475 985 476 989
rect 470 984 476 985
rect 526 989 532 990
rect 526 985 527 989
rect 531 985 532 989
rect 526 984 532 985
rect 590 989 596 990
rect 590 985 591 989
rect 595 985 596 989
rect 590 984 596 985
rect 654 989 660 990
rect 654 985 655 989
rect 659 985 660 989
rect 654 984 660 985
rect 718 989 724 990
rect 718 985 719 989
rect 723 985 724 989
rect 718 984 724 985
rect 782 989 788 990
rect 782 985 783 989
rect 787 985 788 989
rect 782 984 788 985
rect 846 989 852 990
rect 846 985 847 989
rect 851 985 852 989
rect 846 984 852 985
rect 910 989 916 990
rect 910 985 911 989
rect 915 985 916 989
rect 910 984 916 985
rect 974 989 980 990
rect 974 985 975 989
rect 979 985 980 989
rect 974 984 980 985
rect 1038 989 1044 990
rect 1038 985 1039 989
rect 1043 985 1044 989
rect 1038 984 1044 985
rect 1102 989 1108 990
rect 1102 985 1103 989
rect 1107 985 1108 989
rect 1102 984 1108 985
rect 1158 989 1164 990
rect 1158 985 1159 989
rect 1163 985 1164 989
rect 1158 984 1164 985
rect 1214 989 1220 990
rect 1214 985 1215 989
rect 1219 985 1220 989
rect 1214 984 1220 985
rect 1270 989 1276 990
rect 1270 985 1271 989
rect 1275 985 1276 989
rect 1270 984 1276 985
rect 1326 988 1332 989
rect 1326 984 1327 988
rect 1331 984 1332 988
rect 110 983 116 984
rect 1326 983 1332 984
rect 1398 981 1404 982
rect 1366 980 1372 981
rect 1366 976 1367 980
rect 1371 976 1372 980
rect 1398 977 1399 981
rect 1403 977 1404 981
rect 1398 976 1404 977
rect 1454 981 1460 982
rect 1454 977 1455 981
rect 1459 977 1460 981
rect 1454 976 1460 977
rect 1510 981 1516 982
rect 1510 977 1511 981
rect 1515 977 1516 981
rect 1510 976 1516 977
rect 1566 981 1572 982
rect 1566 977 1567 981
rect 1571 977 1572 981
rect 1566 976 1572 977
rect 1638 981 1644 982
rect 1638 977 1639 981
rect 1643 977 1644 981
rect 1638 976 1644 977
rect 1718 981 1724 982
rect 1718 977 1719 981
rect 1723 977 1724 981
rect 1718 976 1724 977
rect 1806 981 1812 982
rect 1806 977 1807 981
rect 1811 977 1812 981
rect 1806 976 1812 977
rect 1902 981 1908 982
rect 1902 977 1903 981
rect 1907 977 1908 981
rect 1902 976 1908 977
rect 2014 981 2020 982
rect 2014 977 2015 981
rect 2019 977 2020 981
rect 2014 976 2020 977
rect 2142 981 2148 982
rect 2142 977 2143 981
rect 2147 977 2148 981
rect 2142 976 2148 977
rect 2270 981 2276 982
rect 2270 977 2271 981
rect 2275 977 2276 981
rect 2270 976 2276 977
rect 2406 981 2412 982
rect 2406 977 2407 981
rect 2411 977 2412 981
rect 2406 976 2412 977
rect 2526 981 2532 982
rect 2526 977 2527 981
rect 2531 977 2532 981
rect 2526 976 2532 977
rect 2582 980 2588 981
rect 2582 976 2583 980
rect 2587 976 2588 980
rect 1366 975 1372 976
rect 2582 975 2588 976
rect 110 971 116 972
rect 110 967 111 971
rect 115 967 116 971
rect 110 966 116 967
rect 1326 971 1332 972
rect 1326 967 1327 971
rect 1331 967 1332 971
rect 1326 966 1332 967
rect 1366 963 1372 964
rect 430 962 436 963
rect 430 958 431 962
rect 435 958 436 962
rect 430 957 436 958
rect 486 962 492 963
rect 486 958 487 962
rect 491 958 492 962
rect 486 957 492 958
rect 542 962 548 963
rect 542 958 543 962
rect 547 958 548 962
rect 542 957 548 958
rect 606 962 612 963
rect 606 958 607 962
rect 611 958 612 962
rect 606 957 612 958
rect 670 962 676 963
rect 670 958 671 962
rect 675 958 676 962
rect 670 957 676 958
rect 734 962 740 963
rect 734 958 735 962
rect 739 958 740 962
rect 734 957 740 958
rect 798 962 804 963
rect 798 958 799 962
rect 803 958 804 962
rect 798 957 804 958
rect 862 962 868 963
rect 862 958 863 962
rect 867 958 868 962
rect 862 957 868 958
rect 926 962 932 963
rect 926 958 927 962
rect 931 958 932 962
rect 926 957 932 958
rect 990 962 996 963
rect 990 958 991 962
rect 995 958 996 962
rect 990 957 996 958
rect 1054 962 1060 963
rect 1054 958 1055 962
rect 1059 958 1060 962
rect 1054 957 1060 958
rect 1118 962 1124 963
rect 1118 958 1119 962
rect 1123 958 1124 962
rect 1118 957 1124 958
rect 1174 962 1180 963
rect 1174 958 1175 962
rect 1179 958 1180 962
rect 1174 957 1180 958
rect 1230 962 1236 963
rect 1230 958 1231 962
rect 1235 958 1236 962
rect 1230 957 1236 958
rect 1286 962 1292 963
rect 1286 958 1287 962
rect 1291 958 1292 962
rect 1366 959 1367 963
rect 1371 959 1372 963
rect 1366 958 1372 959
rect 2582 963 2588 964
rect 2582 959 2583 963
rect 2587 959 2588 963
rect 2582 958 2588 959
rect 1286 957 1292 958
rect 1414 954 1420 955
rect 1414 950 1415 954
rect 1419 950 1420 954
rect 1414 949 1420 950
rect 1470 954 1476 955
rect 1470 950 1471 954
rect 1475 950 1476 954
rect 1470 949 1476 950
rect 1526 954 1532 955
rect 1526 950 1527 954
rect 1531 950 1532 954
rect 1526 949 1532 950
rect 1582 954 1588 955
rect 1582 950 1583 954
rect 1587 950 1588 954
rect 1582 949 1588 950
rect 1654 954 1660 955
rect 1654 950 1655 954
rect 1659 950 1660 954
rect 1654 949 1660 950
rect 1734 954 1740 955
rect 1734 950 1735 954
rect 1739 950 1740 954
rect 1734 949 1740 950
rect 1822 954 1828 955
rect 1822 950 1823 954
rect 1827 950 1828 954
rect 1822 949 1828 950
rect 1918 954 1924 955
rect 1918 950 1919 954
rect 1923 950 1924 954
rect 1918 949 1924 950
rect 2030 954 2036 955
rect 2030 950 2031 954
rect 2035 950 2036 954
rect 2030 949 2036 950
rect 2158 954 2164 955
rect 2158 950 2159 954
rect 2163 950 2164 954
rect 2158 949 2164 950
rect 2286 954 2292 955
rect 2286 950 2287 954
rect 2291 950 2292 954
rect 2286 949 2292 950
rect 2422 954 2428 955
rect 2422 950 2423 954
rect 2427 950 2428 954
rect 2422 949 2428 950
rect 2542 954 2548 955
rect 2542 950 2543 954
rect 2547 950 2548 954
rect 2542 949 2548 950
rect 422 934 428 935
rect 422 930 423 934
rect 427 930 428 934
rect 422 929 428 930
rect 478 934 484 935
rect 478 930 479 934
rect 483 930 484 934
rect 478 929 484 930
rect 534 934 540 935
rect 534 930 535 934
rect 539 930 540 934
rect 534 929 540 930
rect 590 934 596 935
rect 590 930 591 934
rect 595 930 596 934
rect 590 929 596 930
rect 646 934 652 935
rect 646 930 647 934
rect 651 930 652 934
rect 646 929 652 930
rect 702 934 708 935
rect 702 930 703 934
rect 707 930 708 934
rect 702 929 708 930
rect 758 934 764 935
rect 758 930 759 934
rect 763 930 764 934
rect 758 929 764 930
rect 814 934 820 935
rect 814 930 815 934
rect 819 930 820 934
rect 814 929 820 930
rect 110 925 116 926
rect 110 921 111 925
rect 115 921 116 925
rect 110 920 116 921
rect 1326 925 1332 926
rect 1326 921 1327 925
rect 1331 921 1332 925
rect 1326 920 1332 921
rect 1414 922 1420 923
rect 1414 918 1415 922
rect 1419 918 1420 922
rect 1414 917 1420 918
rect 1470 922 1476 923
rect 1470 918 1471 922
rect 1475 918 1476 922
rect 1470 917 1476 918
rect 1526 922 1532 923
rect 1526 918 1527 922
rect 1531 918 1532 922
rect 1526 917 1532 918
rect 1614 922 1620 923
rect 1614 918 1615 922
rect 1619 918 1620 922
rect 1614 917 1620 918
rect 1710 922 1716 923
rect 1710 918 1711 922
rect 1715 918 1716 922
rect 1710 917 1716 918
rect 1822 922 1828 923
rect 1822 918 1823 922
rect 1827 918 1828 922
rect 1822 917 1828 918
rect 1942 922 1948 923
rect 1942 918 1943 922
rect 1947 918 1948 922
rect 1942 917 1948 918
rect 2062 922 2068 923
rect 2062 918 2063 922
rect 2067 918 2068 922
rect 2062 917 2068 918
rect 2182 922 2188 923
rect 2182 918 2183 922
rect 2187 918 2188 922
rect 2182 917 2188 918
rect 2310 922 2316 923
rect 2310 918 2311 922
rect 2315 918 2316 922
rect 2310 917 2316 918
rect 2438 922 2444 923
rect 2438 918 2439 922
rect 2443 918 2444 922
rect 2438 917 2444 918
rect 2542 922 2548 923
rect 2542 918 2543 922
rect 2547 918 2548 922
rect 2542 917 2548 918
rect 1366 913 1372 914
rect 1366 909 1367 913
rect 1371 909 1372 913
rect 110 908 116 909
rect 1326 908 1332 909
rect 1366 908 1372 909
rect 2582 913 2588 914
rect 2582 909 2583 913
rect 2587 909 2588 913
rect 2582 908 2588 909
rect 110 904 111 908
rect 115 904 116 908
rect 110 903 116 904
rect 406 907 412 908
rect 406 903 407 907
rect 411 903 412 907
rect 406 902 412 903
rect 462 907 468 908
rect 462 903 463 907
rect 467 903 468 907
rect 462 902 468 903
rect 518 907 524 908
rect 518 903 519 907
rect 523 903 524 907
rect 518 902 524 903
rect 574 907 580 908
rect 574 903 575 907
rect 579 903 580 907
rect 574 902 580 903
rect 630 907 636 908
rect 630 903 631 907
rect 635 903 636 907
rect 630 902 636 903
rect 686 907 692 908
rect 686 903 687 907
rect 691 903 692 907
rect 686 902 692 903
rect 742 907 748 908
rect 742 903 743 907
rect 747 903 748 907
rect 742 902 748 903
rect 798 907 804 908
rect 798 903 799 907
rect 803 903 804 907
rect 1326 904 1327 908
rect 1331 904 1332 908
rect 1326 903 1332 904
rect 798 902 804 903
rect 1366 896 1372 897
rect 2582 896 2588 897
rect 1366 892 1367 896
rect 1371 892 1372 896
rect 1366 891 1372 892
rect 1398 895 1404 896
rect 1398 891 1399 895
rect 1403 891 1404 895
rect 1398 890 1404 891
rect 1454 895 1460 896
rect 1454 891 1455 895
rect 1459 891 1460 895
rect 1454 890 1460 891
rect 1510 895 1516 896
rect 1510 891 1511 895
rect 1515 891 1516 895
rect 1510 890 1516 891
rect 1598 895 1604 896
rect 1598 891 1599 895
rect 1603 891 1604 895
rect 1598 890 1604 891
rect 1694 895 1700 896
rect 1694 891 1695 895
rect 1699 891 1700 895
rect 1694 890 1700 891
rect 1806 895 1812 896
rect 1806 891 1807 895
rect 1811 891 1812 895
rect 1806 890 1812 891
rect 1926 895 1932 896
rect 1926 891 1927 895
rect 1931 891 1932 895
rect 1926 890 1932 891
rect 2046 895 2052 896
rect 2046 891 2047 895
rect 2051 891 2052 895
rect 2046 890 2052 891
rect 2166 895 2172 896
rect 2166 891 2167 895
rect 2171 891 2172 895
rect 2166 890 2172 891
rect 2294 895 2300 896
rect 2294 891 2295 895
rect 2299 891 2300 895
rect 2294 890 2300 891
rect 2422 895 2428 896
rect 2422 891 2423 895
rect 2427 891 2428 895
rect 2422 890 2428 891
rect 2526 895 2532 896
rect 2526 891 2527 895
rect 2531 891 2532 895
rect 2582 892 2583 896
rect 2587 892 2588 896
rect 2582 891 2588 892
rect 2526 890 2532 891
rect 278 873 284 874
rect 110 872 116 873
rect 110 868 111 872
rect 115 868 116 872
rect 278 869 279 873
rect 283 869 284 873
rect 278 868 284 869
rect 334 873 340 874
rect 334 869 335 873
rect 339 869 340 873
rect 334 868 340 869
rect 390 873 396 874
rect 390 869 391 873
rect 395 869 396 873
rect 390 868 396 869
rect 454 873 460 874
rect 454 869 455 873
rect 459 869 460 873
rect 454 868 460 869
rect 518 873 524 874
rect 518 869 519 873
rect 523 869 524 873
rect 518 868 524 869
rect 582 873 588 874
rect 582 869 583 873
rect 587 869 588 873
rect 582 868 588 869
rect 646 873 652 874
rect 646 869 647 873
rect 651 869 652 873
rect 646 868 652 869
rect 710 873 716 874
rect 710 869 711 873
rect 715 869 716 873
rect 710 868 716 869
rect 774 873 780 874
rect 774 869 775 873
rect 779 869 780 873
rect 774 868 780 869
rect 846 873 852 874
rect 846 869 847 873
rect 851 869 852 873
rect 846 868 852 869
rect 918 873 924 874
rect 918 869 919 873
rect 923 869 924 873
rect 918 868 924 869
rect 1326 872 1332 873
rect 1326 868 1327 872
rect 1331 868 1332 872
rect 110 867 116 868
rect 1326 867 1332 868
rect 1470 861 1476 862
rect 1366 860 1372 861
rect 1366 856 1367 860
rect 1371 856 1372 860
rect 1470 857 1471 861
rect 1475 857 1476 861
rect 1470 856 1476 857
rect 1550 861 1556 862
rect 1550 857 1551 861
rect 1555 857 1556 861
rect 1550 856 1556 857
rect 1638 861 1644 862
rect 1638 857 1639 861
rect 1643 857 1644 861
rect 1638 856 1644 857
rect 1726 861 1732 862
rect 1726 857 1727 861
rect 1731 857 1732 861
rect 1726 856 1732 857
rect 1814 861 1820 862
rect 1814 857 1815 861
rect 1819 857 1820 861
rect 1814 856 1820 857
rect 1902 861 1908 862
rect 1902 857 1903 861
rect 1907 857 1908 861
rect 1902 856 1908 857
rect 1990 861 1996 862
rect 1990 857 1991 861
rect 1995 857 1996 861
rect 1990 856 1996 857
rect 2070 861 2076 862
rect 2070 857 2071 861
rect 2075 857 2076 861
rect 2070 856 2076 857
rect 2142 861 2148 862
rect 2142 857 2143 861
rect 2147 857 2148 861
rect 2142 856 2148 857
rect 2214 861 2220 862
rect 2214 857 2215 861
rect 2219 857 2220 861
rect 2214 856 2220 857
rect 2278 861 2284 862
rect 2278 857 2279 861
rect 2283 857 2284 861
rect 2278 856 2284 857
rect 2342 861 2348 862
rect 2342 857 2343 861
rect 2347 857 2348 861
rect 2342 856 2348 857
rect 2406 861 2412 862
rect 2406 857 2407 861
rect 2411 857 2412 861
rect 2406 856 2412 857
rect 2470 861 2476 862
rect 2470 857 2471 861
rect 2475 857 2476 861
rect 2470 856 2476 857
rect 2526 861 2532 862
rect 2526 857 2527 861
rect 2531 857 2532 861
rect 2526 856 2532 857
rect 2582 860 2588 861
rect 2582 856 2583 860
rect 2587 856 2588 860
rect 110 855 116 856
rect 110 851 111 855
rect 115 851 116 855
rect 110 850 116 851
rect 1326 855 1332 856
rect 1366 855 1372 856
rect 2582 855 2588 856
rect 1326 851 1327 855
rect 1331 851 1332 855
rect 1326 850 1332 851
rect 294 846 300 847
rect 294 842 295 846
rect 299 842 300 846
rect 294 841 300 842
rect 350 846 356 847
rect 350 842 351 846
rect 355 842 356 846
rect 350 841 356 842
rect 406 846 412 847
rect 406 842 407 846
rect 411 842 412 846
rect 406 841 412 842
rect 470 846 476 847
rect 470 842 471 846
rect 475 842 476 846
rect 470 841 476 842
rect 534 846 540 847
rect 534 842 535 846
rect 539 842 540 846
rect 534 841 540 842
rect 598 846 604 847
rect 598 842 599 846
rect 603 842 604 846
rect 598 841 604 842
rect 662 846 668 847
rect 662 842 663 846
rect 667 842 668 846
rect 662 841 668 842
rect 726 846 732 847
rect 726 842 727 846
rect 731 842 732 846
rect 726 841 732 842
rect 790 846 796 847
rect 790 842 791 846
rect 795 842 796 846
rect 790 841 796 842
rect 862 846 868 847
rect 862 842 863 846
rect 867 842 868 846
rect 862 841 868 842
rect 934 846 940 847
rect 934 842 935 846
rect 939 842 940 846
rect 934 841 940 842
rect 1366 843 1372 844
rect 1366 839 1367 843
rect 1371 839 1372 843
rect 1366 838 1372 839
rect 2582 843 2588 844
rect 2582 839 2583 843
rect 2587 839 2588 843
rect 2582 838 2588 839
rect 1486 834 1492 835
rect 1486 830 1487 834
rect 1491 830 1492 834
rect 1486 829 1492 830
rect 1566 834 1572 835
rect 1566 830 1567 834
rect 1571 830 1572 834
rect 1566 829 1572 830
rect 1654 834 1660 835
rect 1654 830 1655 834
rect 1659 830 1660 834
rect 1654 829 1660 830
rect 1742 834 1748 835
rect 1742 830 1743 834
rect 1747 830 1748 834
rect 1742 829 1748 830
rect 1830 834 1836 835
rect 1830 830 1831 834
rect 1835 830 1836 834
rect 1830 829 1836 830
rect 1918 834 1924 835
rect 1918 830 1919 834
rect 1923 830 1924 834
rect 1918 829 1924 830
rect 2006 834 2012 835
rect 2006 830 2007 834
rect 2011 830 2012 834
rect 2006 829 2012 830
rect 2086 834 2092 835
rect 2086 830 2087 834
rect 2091 830 2092 834
rect 2086 829 2092 830
rect 2158 834 2164 835
rect 2158 830 2159 834
rect 2163 830 2164 834
rect 2158 829 2164 830
rect 2230 834 2236 835
rect 2230 830 2231 834
rect 2235 830 2236 834
rect 2230 829 2236 830
rect 2294 834 2300 835
rect 2294 830 2295 834
rect 2299 830 2300 834
rect 2294 829 2300 830
rect 2358 834 2364 835
rect 2358 830 2359 834
rect 2363 830 2364 834
rect 2358 829 2364 830
rect 2422 834 2428 835
rect 2422 830 2423 834
rect 2427 830 2428 834
rect 2422 829 2428 830
rect 2486 834 2492 835
rect 2486 830 2487 834
rect 2491 830 2492 834
rect 2486 829 2492 830
rect 2542 834 2548 835
rect 2542 830 2543 834
rect 2547 830 2548 834
rect 2542 829 2548 830
rect 166 814 172 815
rect 166 810 167 814
rect 171 810 172 814
rect 166 809 172 810
rect 230 814 236 815
rect 230 810 231 814
rect 235 810 236 814
rect 230 809 236 810
rect 310 814 316 815
rect 310 810 311 814
rect 315 810 316 814
rect 310 809 316 810
rect 398 814 404 815
rect 398 810 399 814
rect 403 810 404 814
rect 398 809 404 810
rect 486 814 492 815
rect 486 810 487 814
rect 491 810 492 814
rect 486 809 492 810
rect 582 814 588 815
rect 582 810 583 814
rect 587 810 588 814
rect 582 809 588 810
rect 670 814 676 815
rect 670 810 671 814
rect 675 810 676 814
rect 670 809 676 810
rect 758 814 764 815
rect 758 810 759 814
rect 763 810 764 814
rect 758 809 764 810
rect 838 814 844 815
rect 838 810 839 814
rect 843 810 844 814
rect 838 809 844 810
rect 918 814 924 815
rect 918 810 919 814
rect 923 810 924 814
rect 918 809 924 810
rect 1006 814 1012 815
rect 1006 810 1007 814
rect 1011 810 1012 814
rect 1006 809 1012 810
rect 1094 814 1100 815
rect 1094 810 1095 814
rect 1099 810 1100 814
rect 1094 809 1100 810
rect 110 805 116 806
rect 110 801 111 805
rect 115 801 116 805
rect 110 800 116 801
rect 1326 805 1332 806
rect 1326 801 1327 805
rect 1331 801 1332 805
rect 1326 800 1332 801
rect 1630 802 1636 803
rect 1630 798 1631 802
rect 1635 798 1636 802
rect 1630 797 1636 798
rect 1686 802 1692 803
rect 1686 798 1687 802
rect 1691 798 1692 802
rect 1686 797 1692 798
rect 1750 802 1756 803
rect 1750 798 1751 802
rect 1755 798 1756 802
rect 1750 797 1756 798
rect 1822 802 1828 803
rect 1822 798 1823 802
rect 1827 798 1828 802
rect 1822 797 1828 798
rect 1902 802 1908 803
rect 1902 798 1903 802
rect 1907 798 1908 802
rect 1902 797 1908 798
rect 1990 802 1996 803
rect 1990 798 1991 802
rect 1995 798 1996 802
rect 1990 797 1996 798
rect 2070 802 2076 803
rect 2070 798 2071 802
rect 2075 798 2076 802
rect 2070 797 2076 798
rect 2158 802 2164 803
rect 2158 798 2159 802
rect 2163 798 2164 802
rect 2158 797 2164 798
rect 2246 802 2252 803
rect 2246 798 2247 802
rect 2251 798 2252 802
rect 2246 797 2252 798
rect 2334 802 2340 803
rect 2334 798 2335 802
rect 2339 798 2340 802
rect 2334 797 2340 798
rect 2422 802 2428 803
rect 2422 798 2423 802
rect 2427 798 2428 802
rect 2422 797 2428 798
rect 1366 793 1372 794
rect 1366 789 1367 793
rect 1371 789 1372 793
rect 110 788 116 789
rect 1326 788 1332 789
rect 1366 788 1372 789
rect 2582 793 2588 794
rect 2582 789 2583 793
rect 2587 789 2588 793
rect 2582 788 2588 789
rect 110 784 111 788
rect 115 784 116 788
rect 110 783 116 784
rect 150 787 156 788
rect 150 783 151 787
rect 155 783 156 787
rect 150 782 156 783
rect 214 787 220 788
rect 214 783 215 787
rect 219 783 220 787
rect 214 782 220 783
rect 294 787 300 788
rect 294 783 295 787
rect 299 783 300 787
rect 294 782 300 783
rect 382 787 388 788
rect 382 783 383 787
rect 387 783 388 787
rect 382 782 388 783
rect 470 787 476 788
rect 470 783 471 787
rect 475 783 476 787
rect 470 782 476 783
rect 566 787 572 788
rect 566 783 567 787
rect 571 783 572 787
rect 566 782 572 783
rect 654 787 660 788
rect 654 783 655 787
rect 659 783 660 787
rect 654 782 660 783
rect 742 787 748 788
rect 742 783 743 787
rect 747 783 748 787
rect 742 782 748 783
rect 822 787 828 788
rect 822 783 823 787
rect 827 783 828 787
rect 822 782 828 783
rect 902 787 908 788
rect 902 783 903 787
rect 907 783 908 787
rect 902 782 908 783
rect 990 787 996 788
rect 990 783 991 787
rect 995 783 996 787
rect 990 782 996 783
rect 1078 787 1084 788
rect 1078 783 1079 787
rect 1083 783 1084 787
rect 1326 784 1327 788
rect 1331 784 1332 788
rect 1326 783 1332 784
rect 1078 782 1084 783
rect 1366 776 1372 777
rect 2582 776 2588 777
rect 1366 772 1367 776
rect 1371 772 1372 776
rect 1366 771 1372 772
rect 1614 775 1620 776
rect 1614 771 1615 775
rect 1619 771 1620 775
rect 1614 770 1620 771
rect 1670 775 1676 776
rect 1670 771 1671 775
rect 1675 771 1676 775
rect 1670 770 1676 771
rect 1734 775 1740 776
rect 1734 771 1735 775
rect 1739 771 1740 775
rect 1734 770 1740 771
rect 1806 775 1812 776
rect 1806 771 1807 775
rect 1811 771 1812 775
rect 1806 770 1812 771
rect 1886 775 1892 776
rect 1886 771 1887 775
rect 1891 771 1892 775
rect 1886 770 1892 771
rect 1974 775 1980 776
rect 1974 771 1975 775
rect 1979 771 1980 775
rect 1974 770 1980 771
rect 2054 775 2060 776
rect 2054 771 2055 775
rect 2059 771 2060 775
rect 2054 770 2060 771
rect 2142 775 2148 776
rect 2142 771 2143 775
rect 2147 771 2148 775
rect 2142 770 2148 771
rect 2230 775 2236 776
rect 2230 771 2231 775
rect 2235 771 2236 775
rect 2230 770 2236 771
rect 2318 775 2324 776
rect 2318 771 2319 775
rect 2323 771 2324 775
rect 2318 770 2324 771
rect 2406 775 2412 776
rect 2406 771 2407 775
rect 2411 771 2412 775
rect 2582 772 2583 776
rect 2587 772 2588 776
rect 2582 771 2588 772
rect 2406 770 2412 771
rect 142 745 148 746
rect 110 744 116 745
rect 110 740 111 744
rect 115 740 116 744
rect 142 741 143 745
rect 147 741 148 745
rect 142 740 148 741
rect 198 745 204 746
rect 198 741 199 745
rect 203 741 204 745
rect 198 740 204 741
rect 278 745 284 746
rect 278 741 279 745
rect 283 741 284 745
rect 278 740 284 741
rect 382 745 388 746
rect 382 741 383 745
rect 387 741 388 745
rect 382 740 388 741
rect 486 745 492 746
rect 486 741 487 745
rect 491 741 492 745
rect 486 740 492 741
rect 598 745 604 746
rect 598 741 599 745
rect 603 741 604 745
rect 598 740 604 741
rect 702 745 708 746
rect 702 741 703 745
rect 707 741 708 745
rect 702 740 708 741
rect 806 745 812 746
rect 806 741 807 745
rect 811 741 812 745
rect 806 740 812 741
rect 902 745 908 746
rect 902 741 903 745
rect 907 741 908 745
rect 902 740 908 741
rect 990 745 996 746
rect 990 741 991 745
rect 995 741 996 745
rect 990 740 996 741
rect 1078 745 1084 746
rect 1078 741 1079 745
rect 1083 741 1084 745
rect 1078 740 1084 741
rect 1174 745 1180 746
rect 1174 741 1175 745
rect 1179 741 1180 745
rect 1174 740 1180 741
rect 1326 744 1332 745
rect 1326 740 1327 744
rect 1331 740 1332 744
rect 110 739 116 740
rect 1326 739 1332 740
rect 1566 737 1572 738
rect 1366 736 1372 737
rect 1366 732 1367 736
rect 1371 732 1372 736
rect 1566 733 1567 737
rect 1571 733 1572 737
rect 1566 732 1572 733
rect 1622 737 1628 738
rect 1622 733 1623 737
rect 1627 733 1628 737
rect 1622 732 1628 733
rect 1686 737 1692 738
rect 1686 733 1687 737
rect 1691 733 1692 737
rect 1686 732 1692 733
rect 1758 737 1764 738
rect 1758 733 1759 737
rect 1763 733 1764 737
rect 1758 732 1764 733
rect 1838 737 1844 738
rect 1838 733 1839 737
rect 1843 733 1844 737
rect 1838 732 1844 733
rect 1918 737 1924 738
rect 1918 733 1919 737
rect 1923 733 1924 737
rect 1918 732 1924 733
rect 1998 737 2004 738
rect 1998 733 1999 737
rect 2003 733 2004 737
rect 1998 732 2004 733
rect 2078 737 2084 738
rect 2078 733 2079 737
rect 2083 733 2084 737
rect 2078 732 2084 733
rect 2158 737 2164 738
rect 2158 733 2159 737
rect 2163 733 2164 737
rect 2158 732 2164 733
rect 2246 737 2252 738
rect 2246 733 2247 737
rect 2251 733 2252 737
rect 2246 732 2252 733
rect 2334 737 2340 738
rect 2334 733 2335 737
rect 2339 733 2340 737
rect 2334 732 2340 733
rect 2582 736 2588 737
rect 2582 732 2583 736
rect 2587 732 2588 736
rect 1366 731 1372 732
rect 2582 731 2588 732
rect 110 727 116 728
rect 110 723 111 727
rect 115 723 116 727
rect 110 722 116 723
rect 1326 727 1332 728
rect 1326 723 1327 727
rect 1331 723 1332 727
rect 1326 722 1332 723
rect 1366 719 1372 720
rect 158 718 164 719
rect 158 714 159 718
rect 163 714 164 718
rect 158 713 164 714
rect 214 718 220 719
rect 214 714 215 718
rect 219 714 220 718
rect 214 713 220 714
rect 294 718 300 719
rect 294 714 295 718
rect 299 714 300 718
rect 294 713 300 714
rect 398 718 404 719
rect 398 714 399 718
rect 403 714 404 718
rect 398 713 404 714
rect 502 718 508 719
rect 502 714 503 718
rect 507 714 508 718
rect 502 713 508 714
rect 614 718 620 719
rect 614 714 615 718
rect 619 714 620 718
rect 614 713 620 714
rect 718 718 724 719
rect 718 714 719 718
rect 723 714 724 718
rect 718 713 724 714
rect 822 718 828 719
rect 822 714 823 718
rect 827 714 828 718
rect 822 713 828 714
rect 918 718 924 719
rect 918 714 919 718
rect 923 714 924 718
rect 918 713 924 714
rect 1006 718 1012 719
rect 1006 714 1007 718
rect 1011 714 1012 718
rect 1006 713 1012 714
rect 1094 718 1100 719
rect 1094 714 1095 718
rect 1099 714 1100 718
rect 1094 713 1100 714
rect 1190 718 1196 719
rect 1190 714 1191 718
rect 1195 714 1196 718
rect 1366 715 1367 719
rect 1371 715 1372 719
rect 1366 714 1372 715
rect 2582 719 2588 720
rect 2582 715 2583 719
rect 2587 715 2588 719
rect 2582 714 2588 715
rect 1190 713 1196 714
rect 1582 710 1588 711
rect 1582 706 1583 710
rect 1587 706 1588 710
rect 1582 705 1588 706
rect 1638 710 1644 711
rect 1638 706 1639 710
rect 1643 706 1644 710
rect 1638 705 1644 706
rect 1702 710 1708 711
rect 1702 706 1703 710
rect 1707 706 1708 710
rect 1702 705 1708 706
rect 1774 710 1780 711
rect 1774 706 1775 710
rect 1779 706 1780 710
rect 1774 705 1780 706
rect 1854 710 1860 711
rect 1854 706 1855 710
rect 1859 706 1860 710
rect 1854 705 1860 706
rect 1934 710 1940 711
rect 1934 706 1935 710
rect 1939 706 1940 710
rect 1934 705 1940 706
rect 2014 710 2020 711
rect 2014 706 2015 710
rect 2019 706 2020 710
rect 2014 705 2020 706
rect 2094 710 2100 711
rect 2094 706 2095 710
rect 2099 706 2100 710
rect 2094 705 2100 706
rect 2174 710 2180 711
rect 2174 706 2175 710
rect 2179 706 2180 710
rect 2174 705 2180 706
rect 2262 710 2268 711
rect 2262 706 2263 710
rect 2267 706 2268 710
rect 2262 705 2268 706
rect 2350 710 2356 711
rect 2350 706 2351 710
rect 2355 706 2356 710
rect 2350 705 2356 706
rect 158 690 164 691
rect 158 686 159 690
rect 163 686 164 690
rect 158 685 164 686
rect 214 690 220 691
rect 214 686 215 690
rect 219 686 220 690
rect 214 685 220 686
rect 278 690 284 691
rect 278 686 279 690
rect 283 686 284 690
rect 278 685 284 686
rect 358 690 364 691
rect 358 686 359 690
rect 363 686 364 690
rect 358 685 364 686
rect 446 690 452 691
rect 446 686 447 690
rect 451 686 452 690
rect 446 685 452 686
rect 534 690 540 691
rect 534 686 535 690
rect 539 686 540 690
rect 534 685 540 686
rect 622 690 628 691
rect 622 686 623 690
rect 627 686 628 690
rect 622 685 628 686
rect 710 690 716 691
rect 710 686 711 690
rect 715 686 716 690
rect 710 685 716 686
rect 790 690 796 691
rect 790 686 791 690
rect 795 686 796 690
rect 790 685 796 686
rect 870 690 876 691
rect 870 686 871 690
rect 875 686 876 690
rect 870 685 876 686
rect 950 690 956 691
rect 950 686 951 690
rect 955 686 956 690
rect 950 685 956 686
rect 1038 690 1044 691
rect 1038 686 1039 690
rect 1043 686 1044 690
rect 1038 685 1044 686
rect 1414 682 1420 683
rect 110 681 116 682
rect 110 677 111 681
rect 115 677 116 681
rect 110 676 116 677
rect 1326 681 1332 682
rect 1326 677 1327 681
rect 1331 677 1332 681
rect 1414 678 1415 682
rect 1419 678 1420 682
rect 1414 677 1420 678
rect 1510 682 1516 683
rect 1510 678 1511 682
rect 1515 678 1516 682
rect 1510 677 1516 678
rect 1614 682 1620 683
rect 1614 678 1615 682
rect 1619 678 1620 682
rect 1614 677 1620 678
rect 1718 682 1724 683
rect 1718 678 1719 682
rect 1723 678 1724 682
rect 1718 677 1724 678
rect 1822 682 1828 683
rect 1822 678 1823 682
rect 1827 678 1828 682
rect 1822 677 1828 678
rect 1926 682 1932 683
rect 1926 678 1927 682
rect 1931 678 1932 682
rect 1926 677 1932 678
rect 2022 682 2028 683
rect 2022 678 2023 682
rect 2027 678 2028 682
rect 2022 677 2028 678
rect 2118 682 2124 683
rect 2118 678 2119 682
rect 2123 678 2124 682
rect 2118 677 2124 678
rect 2206 682 2212 683
rect 2206 678 2207 682
rect 2211 678 2212 682
rect 2206 677 2212 678
rect 2294 682 2300 683
rect 2294 678 2295 682
rect 2299 678 2300 682
rect 2294 677 2300 678
rect 2390 682 2396 683
rect 2390 678 2391 682
rect 2395 678 2396 682
rect 2390 677 2396 678
rect 1326 676 1332 677
rect 1366 673 1372 674
rect 1366 669 1367 673
rect 1371 669 1372 673
rect 1366 668 1372 669
rect 2582 673 2588 674
rect 2582 669 2583 673
rect 2587 669 2588 673
rect 2582 668 2588 669
rect 110 664 116 665
rect 1326 664 1332 665
rect 110 660 111 664
rect 115 660 116 664
rect 110 659 116 660
rect 142 663 148 664
rect 142 659 143 663
rect 147 659 148 663
rect 142 658 148 659
rect 198 663 204 664
rect 198 659 199 663
rect 203 659 204 663
rect 198 658 204 659
rect 262 663 268 664
rect 262 659 263 663
rect 267 659 268 663
rect 262 658 268 659
rect 342 663 348 664
rect 342 659 343 663
rect 347 659 348 663
rect 342 658 348 659
rect 430 663 436 664
rect 430 659 431 663
rect 435 659 436 663
rect 430 658 436 659
rect 518 663 524 664
rect 518 659 519 663
rect 523 659 524 663
rect 518 658 524 659
rect 606 663 612 664
rect 606 659 607 663
rect 611 659 612 663
rect 606 658 612 659
rect 694 663 700 664
rect 694 659 695 663
rect 699 659 700 663
rect 694 658 700 659
rect 774 663 780 664
rect 774 659 775 663
rect 779 659 780 663
rect 774 658 780 659
rect 854 663 860 664
rect 854 659 855 663
rect 859 659 860 663
rect 854 658 860 659
rect 934 663 940 664
rect 934 659 935 663
rect 939 659 940 663
rect 934 658 940 659
rect 1022 663 1028 664
rect 1022 659 1023 663
rect 1027 659 1028 663
rect 1326 660 1327 664
rect 1331 660 1332 664
rect 1326 659 1332 660
rect 1022 658 1028 659
rect 1366 656 1372 657
rect 2582 656 2588 657
rect 1366 652 1367 656
rect 1371 652 1372 656
rect 1366 651 1372 652
rect 1398 655 1404 656
rect 1398 651 1399 655
rect 1403 651 1404 655
rect 1398 650 1404 651
rect 1494 655 1500 656
rect 1494 651 1495 655
rect 1499 651 1500 655
rect 1494 650 1500 651
rect 1598 655 1604 656
rect 1598 651 1599 655
rect 1603 651 1604 655
rect 1598 650 1604 651
rect 1702 655 1708 656
rect 1702 651 1703 655
rect 1707 651 1708 655
rect 1702 650 1708 651
rect 1806 655 1812 656
rect 1806 651 1807 655
rect 1811 651 1812 655
rect 1806 650 1812 651
rect 1910 655 1916 656
rect 1910 651 1911 655
rect 1915 651 1916 655
rect 1910 650 1916 651
rect 2006 655 2012 656
rect 2006 651 2007 655
rect 2011 651 2012 655
rect 2006 650 2012 651
rect 2102 655 2108 656
rect 2102 651 2103 655
rect 2107 651 2108 655
rect 2102 650 2108 651
rect 2190 655 2196 656
rect 2190 651 2191 655
rect 2195 651 2196 655
rect 2190 650 2196 651
rect 2278 655 2284 656
rect 2278 651 2279 655
rect 2283 651 2284 655
rect 2278 650 2284 651
rect 2374 655 2380 656
rect 2374 651 2375 655
rect 2379 651 2380 655
rect 2582 652 2583 656
rect 2587 652 2588 656
rect 2582 651 2588 652
rect 2374 650 2380 651
rect 142 621 148 622
rect 110 620 116 621
rect 110 616 111 620
rect 115 616 116 620
rect 142 617 143 621
rect 147 617 148 621
rect 142 616 148 617
rect 198 621 204 622
rect 198 617 199 621
rect 203 617 204 621
rect 198 616 204 617
rect 254 621 260 622
rect 254 617 255 621
rect 259 617 260 621
rect 254 616 260 617
rect 310 621 316 622
rect 310 617 311 621
rect 315 617 316 621
rect 310 616 316 617
rect 390 621 396 622
rect 390 617 391 621
rect 395 617 396 621
rect 390 616 396 617
rect 478 621 484 622
rect 478 617 479 621
rect 483 617 484 621
rect 478 616 484 617
rect 574 621 580 622
rect 574 617 575 621
rect 579 617 580 621
rect 574 616 580 617
rect 678 621 684 622
rect 678 617 679 621
rect 683 617 684 621
rect 678 616 684 617
rect 782 621 788 622
rect 782 617 783 621
rect 787 617 788 621
rect 782 616 788 617
rect 886 621 892 622
rect 886 617 887 621
rect 891 617 892 621
rect 886 616 892 617
rect 990 621 996 622
rect 990 617 991 621
rect 995 617 996 621
rect 990 616 996 617
rect 1086 621 1092 622
rect 1086 617 1087 621
rect 1091 617 1092 621
rect 1086 616 1092 617
rect 1190 621 1196 622
rect 1190 617 1191 621
rect 1195 617 1196 621
rect 1190 616 1196 617
rect 1270 621 1276 622
rect 1398 621 1404 622
rect 1270 617 1271 621
rect 1275 617 1276 621
rect 1270 616 1276 617
rect 1326 620 1332 621
rect 1326 616 1327 620
rect 1331 616 1332 620
rect 110 615 116 616
rect 1326 615 1332 616
rect 1366 620 1372 621
rect 1366 616 1367 620
rect 1371 616 1372 620
rect 1398 617 1399 621
rect 1403 617 1404 621
rect 1398 616 1404 617
rect 1510 621 1516 622
rect 1510 617 1511 621
rect 1515 617 1516 621
rect 1510 616 1516 617
rect 1646 621 1652 622
rect 1646 617 1647 621
rect 1651 617 1652 621
rect 1646 616 1652 617
rect 1782 621 1788 622
rect 1782 617 1783 621
rect 1787 617 1788 621
rect 1782 616 1788 617
rect 1910 621 1916 622
rect 1910 617 1911 621
rect 1915 617 1916 621
rect 1910 616 1916 617
rect 2038 621 2044 622
rect 2038 617 2039 621
rect 2043 617 2044 621
rect 2038 616 2044 617
rect 2158 621 2164 622
rect 2158 617 2159 621
rect 2163 617 2164 621
rect 2158 616 2164 617
rect 2278 621 2284 622
rect 2278 617 2279 621
rect 2283 617 2284 621
rect 2278 616 2284 617
rect 2406 621 2412 622
rect 2406 617 2407 621
rect 2411 617 2412 621
rect 2406 616 2412 617
rect 2582 620 2588 621
rect 2582 616 2583 620
rect 2587 616 2588 620
rect 1366 615 1372 616
rect 2582 615 2588 616
rect 110 603 116 604
rect 110 599 111 603
rect 115 599 116 603
rect 110 598 116 599
rect 1326 603 1332 604
rect 1326 599 1327 603
rect 1331 599 1332 603
rect 1326 598 1332 599
rect 1366 603 1372 604
rect 1366 599 1367 603
rect 1371 599 1372 603
rect 1366 598 1372 599
rect 2582 603 2588 604
rect 2582 599 2583 603
rect 2587 599 2588 603
rect 2582 598 2588 599
rect 158 594 164 595
rect 158 590 159 594
rect 163 590 164 594
rect 158 589 164 590
rect 214 594 220 595
rect 214 590 215 594
rect 219 590 220 594
rect 214 589 220 590
rect 270 594 276 595
rect 270 590 271 594
rect 275 590 276 594
rect 270 589 276 590
rect 326 594 332 595
rect 326 590 327 594
rect 331 590 332 594
rect 326 589 332 590
rect 406 594 412 595
rect 406 590 407 594
rect 411 590 412 594
rect 406 589 412 590
rect 494 594 500 595
rect 494 590 495 594
rect 499 590 500 594
rect 494 589 500 590
rect 590 594 596 595
rect 590 590 591 594
rect 595 590 596 594
rect 590 589 596 590
rect 694 594 700 595
rect 694 590 695 594
rect 699 590 700 594
rect 694 589 700 590
rect 798 594 804 595
rect 798 590 799 594
rect 803 590 804 594
rect 798 589 804 590
rect 902 594 908 595
rect 902 590 903 594
rect 907 590 908 594
rect 902 589 908 590
rect 1006 594 1012 595
rect 1006 590 1007 594
rect 1011 590 1012 594
rect 1006 589 1012 590
rect 1102 594 1108 595
rect 1102 590 1103 594
rect 1107 590 1108 594
rect 1102 589 1108 590
rect 1206 594 1212 595
rect 1206 590 1207 594
rect 1211 590 1212 594
rect 1206 589 1212 590
rect 1286 594 1292 595
rect 1286 590 1287 594
rect 1291 590 1292 594
rect 1286 589 1292 590
rect 1414 594 1420 595
rect 1414 590 1415 594
rect 1419 590 1420 594
rect 1414 589 1420 590
rect 1526 594 1532 595
rect 1526 590 1527 594
rect 1531 590 1532 594
rect 1526 589 1532 590
rect 1662 594 1668 595
rect 1662 590 1663 594
rect 1667 590 1668 594
rect 1662 589 1668 590
rect 1798 594 1804 595
rect 1798 590 1799 594
rect 1803 590 1804 594
rect 1798 589 1804 590
rect 1926 594 1932 595
rect 1926 590 1927 594
rect 1931 590 1932 594
rect 1926 589 1932 590
rect 2054 594 2060 595
rect 2054 590 2055 594
rect 2059 590 2060 594
rect 2054 589 2060 590
rect 2174 594 2180 595
rect 2174 590 2175 594
rect 2179 590 2180 594
rect 2174 589 2180 590
rect 2294 594 2300 595
rect 2294 590 2295 594
rect 2299 590 2300 594
rect 2294 589 2300 590
rect 2422 594 2428 595
rect 2422 590 2423 594
rect 2427 590 2428 594
rect 2422 589 2428 590
rect 198 566 204 567
rect 198 562 199 566
rect 203 562 204 566
rect 198 561 204 562
rect 262 566 268 567
rect 262 562 263 566
rect 267 562 268 566
rect 262 561 268 562
rect 334 566 340 567
rect 334 562 335 566
rect 339 562 340 566
rect 334 561 340 562
rect 414 566 420 567
rect 414 562 415 566
rect 419 562 420 566
rect 414 561 420 562
rect 510 566 516 567
rect 510 562 511 566
rect 515 562 516 566
rect 510 561 516 562
rect 614 566 620 567
rect 614 562 615 566
rect 619 562 620 566
rect 614 561 620 562
rect 718 566 724 567
rect 718 562 719 566
rect 723 562 724 566
rect 718 561 724 562
rect 830 566 836 567
rect 830 562 831 566
rect 835 562 836 566
rect 830 561 836 562
rect 942 566 948 567
rect 942 562 943 566
rect 947 562 948 566
rect 942 561 948 562
rect 1062 566 1068 567
rect 1062 562 1063 566
rect 1067 562 1068 566
rect 1062 561 1068 562
rect 1182 566 1188 567
rect 1182 562 1183 566
rect 1187 562 1188 566
rect 1182 561 1188 562
rect 1286 566 1292 567
rect 1286 562 1287 566
rect 1291 562 1292 566
rect 1286 561 1292 562
rect 1414 562 1420 563
rect 1414 558 1415 562
rect 1419 558 1420 562
rect 110 557 116 558
rect 110 553 111 557
rect 115 553 116 557
rect 110 552 116 553
rect 1326 557 1332 558
rect 1414 557 1420 558
rect 1470 562 1476 563
rect 1470 558 1471 562
rect 1475 558 1476 562
rect 1470 557 1476 558
rect 1550 562 1556 563
rect 1550 558 1551 562
rect 1555 558 1556 562
rect 1550 557 1556 558
rect 1646 562 1652 563
rect 1646 558 1647 562
rect 1651 558 1652 562
rect 1646 557 1652 558
rect 1750 562 1756 563
rect 1750 558 1751 562
rect 1755 558 1756 562
rect 1750 557 1756 558
rect 1854 562 1860 563
rect 1854 558 1855 562
rect 1859 558 1860 562
rect 1854 557 1860 558
rect 1958 562 1964 563
rect 1958 558 1959 562
rect 1963 558 1964 562
rect 1958 557 1964 558
rect 2054 562 2060 563
rect 2054 558 2055 562
rect 2059 558 2060 562
rect 2054 557 2060 558
rect 2150 562 2156 563
rect 2150 558 2151 562
rect 2155 558 2156 562
rect 2150 557 2156 558
rect 2238 562 2244 563
rect 2238 558 2239 562
rect 2243 558 2244 562
rect 2238 557 2244 558
rect 2318 562 2324 563
rect 2318 558 2319 562
rect 2323 558 2324 562
rect 2318 557 2324 558
rect 2398 562 2404 563
rect 2398 558 2399 562
rect 2403 558 2404 562
rect 2398 557 2404 558
rect 2478 562 2484 563
rect 2478 558 2479 562
rect 2483 558 2484 562
rect 2478 557 2484 558
rect 2542 562 2548 563
rect 2542 558 2543 562
rect 2547 558 2548 562
rect 2542 557 2548 558
rect 1326 553 1327 557
rect 1331 553 1332 557
rect 1326 552 1332 553
rect 1366 553 1372 554
rect 1366 549 1367 553
rect 1371 549 1372 553
rect 1366 548 1372 549
rect 2582 553 2588 554
rect 2582 549 2583 553
rect 2587 549 2588 553
rect 2582 548 2588 549
rect 110 540 116 541
rect 1326 540 1332 541
rect 110 536 111 540
rect 115 536 116 540
rect 110 535 116 536
rect 182 539 188 540
rect 182 535 183 539
rect 187 535 188 539
rect 182 534 188 535
rect 246 539 252 540
rect 246 535 247 539
rect 251 535 252 539
rect 246 534 252 535
rect 318 539 324 540
rect 318 535 319 539
rect 323 535 324 539
rect 318 534 324 535
rect 398 539 404 540
rect 398 535 399 539
rect 403 535 404 539
rect 398 534 404 535
rect 494 539 500 540
rect 494 535 495 539
rect 499 535 500 539
rect 494 534 500 535
rect 598 539 604 540
rect 598 535 599 539
rect 603 535 604 539
rect 598 534 604 535
rect 702 539 708 540
rect 702 535 703 539
rect 707 535 708 539
rect 702 534 708 535
rect 814 539 820 540
rect 814 535 815 539
rect 819 535 820 539
rect 814 534 820 535
rect 926 539 932 540
rect 926 535 927 539
rect 931 535 932 539
rect 926 534 932 535
rect 1046 539 1052 540
rect 1046 535 1047 539
rect 1051 535 1052 539
rect 1046 534 1052 535
rect 1166 539 1172 540
rect 1166 535 1167 539
rect 1171 535 1172 539
rect 1166 534 1172 535
rect 1270 539 1276 540
rect 1270 535 1271 539
rect 1275 535 1276 539
rect 1326 536 1327 540
rect 1331 536 1332 540
rect 1326 535 1332 536
rect 1366 536 1372 537
rect 2582 536 2588 537
rect 1270 534 1276 535
rect 1366 532 1367 536
rect 1371 532 1372 536
rect 1366 531 1372 532
rect 1398 535 1404 536
rect 1398 531 1399 535
rect 1403 531 1404 535
rect 1398 530 1404 531
rect 1454 535 1460 536
rect 1454 531 1455 535
rect 1459 531 1460 535
rect 1454 530 1460 531
rect 1534 535 1540 536
rect 1534 531 1535 535
rect 1539 531 1540 535
rect 1534 530 1540 531
rect 1630 535 1636 536
rect 1630 531 1631 535
rect 1635 531 1636 535
rect 1630 530 1636 531
rect 1734 535 1740 536
rect 1734 531 1735 535
rect 1739 531 1740 535
rect 1734 530 1740 531
rect 1838 535 1844 536
rect 1838 531 1839 535
rect 1843 531 1844 535
rect 1838 530 1844 531
rect 1942 535 1948 536
rect 1942 531 1943 535
rect 1947 531 1948 535
rect 1942 530 1948 531
rect 2038 535 2044 536
rect 2038 531 2039 535
rect 2043 531 2044 535
rect 2038 530 2044 531
rect 2134 535 2140 536
rect 2134 531 2135 535
rect 2139 531 2140 535
rect 2134 530 2140 531
rect 2222 535 2228 536
rect 2222 531 2223 535
rect 2227 531 2228 535
rect 2222 530 2228 531
rect 2302 535 2308 536
rect 2302 531 2303 535
rect 2307 531 2308 535
rect 2302 530 2308 531
rect 2382 535 2388 536
rect 2382 531 2383 535
rect 2387 531 2388 535
rect 2382 530 2388 531
rect 2462 535 2468 536
rect 2462 531 2463 535
rect 2467 531 2468 535
rect 2462 530 2468 531
rect 2526 535 2532 536
rect 2526 531 2527 535
rect 2531 531 2532 535
rect 2582 532 2583 536
rect 2587 532 2588 536
rect 2582 531 2588 532
rect 2526 530 2532 531
rect 1534 501 1540 502
rect 1366 500 1372 501
rect 302 497 308 498
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 302 493 303 497
rect 307 493 308 497
rect 302 492 308 493
rect 358 497 364 498
rect 358 493 359 497
rect 363 493 364 497
rect 358 492 364 493
rect 422 497 428 498
rect 422 493 423 497
rect 427 493 428 497
rect 422 492 428 493
rect 494 497 500 498
rect 494 493 495 497
rect 499 493 500 497
rect 494 492 500 493
rect 574 497 580 498
rect 574 493 575 497
rect 579 493 580 497
rect 574 492 580 493
rect 646 497 652 498
rect 646 493 647 497
rect 651 493 652 497
rect 646 492 652 493
rect 718 497 724 498
rect 718 493 719 497
rect 723 493 724 497
rect 718 492 724 493
rect 790 497 796 498
rect 790 493 791 497
rect 795 493 796 497
rect 790 492 796 493
rect 862 497 868 498
rect 862 493 863 497
rect 867 493 868 497
rect 862 492 868 493
rect 934 497 940 498
rect 934 493 935 497
rect 939 493 940 497
rect 934 492 940 493
rect 1006 497 1012 498
rect 1006 493 1007 497
rect 1011 493 1012 497
rect 1006 492 1012 493
rect 1086 497 1092 498
rect 1086 493 1087 497
rect 1091 493 1092 497
rect 1086 492 1092 493
rect 1326 496 1332 497
rect 1326 492 1327 496
rect 1331 492 1332 496
rect 1366 496 1367 500
rect 1371 496 1372 500
rect 1534 497 1535 501
rect 1539 497 1540 501
rect 1534 496 1540 497
rect 1598 501 1604 502
rect 1598 497 1599 501
rect 1603 497 1604 501
rect 1598 496 1604 497
rect 1670 501 1676 502
rect 1670 497 1671 501
rect 1675 497 1676 501
rect 1670 496 1676 497
rect 1750 501 1756 502
rect 1750 497 1751 501
rect 1755 497 1756 501
rect 1750 496 1756 497
rect 1838 501 1844 502
rect 1838 497 1839 501
rect 1843 497 1844 501
rect 1838 496 1844 497
rect 1926 501 1932 502
rect 1926 497 1927 501
rect 1931 497 1932 501
rect 1926 496 1932 497
rect 2014 501 2020 502
rect 2014 497 2015 501
rect 2019 497 2020 501
rect 2014 496 2020 497
rect 2094 501 2100 502
rect 2094 497 2095 501
rect 2099 497 2100 501
rect 2094 496 2100 497
rect 2174 501 2180 502
rect 2174 497 2175 501
rect 2179 497 2180 501
rect 2174 496 2180 497
rect 2254 501 2260 502
rect 2254 497 2255 501
rect 2259 497 2260 501
rect 2254 496 2260 497
rect 2326 501 2332 502
rect 2326 497 2327 501
rect 2331 497 2332 501
rect 2326 496 2332 497
rect 2398 501 2404 502
rect 2398 497 2399 501
rect 2403 497 2404 501
rect 2398 496 2404 497
rect 2470 501 2476 502
rect 2470 497 2471 501
rect 2475 497 2476 501
rect 2470 496 2476 497
rect 2526 501 2532 502
rect 2526 497 2527 501
rect 2531 497 2532 501
rect 2526 496 2532 497
rect 2582 500 2588 501
rect 2582 496 2583 500
rect 2587 496 2588 500
rect 1366 495 1372 496
rect 2582 495 2588 496
rect 110 491 116 492
rect 1326 491 1332 492
rect 1366 483 1372 484
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 110 474 116 475
rect 1326 479 1332 480
rect 1326 475 1327 479
rect 1331 475 1332 479
rect 1366 479 1367 483
rect 1371 479 1372 483
rect 1366 478 1372 479
rect 2582 483 2588 484
rect 2582 479 2583 483
rect 2587 479 2588 483
rect 2582 478 2588 479
rect 1326 474 1332 475
rect 1550 474 1556 475
rect 318 470 324 471
rect 318 466 319 470
rect 323 466 324 470
rect 318 465 324 466
rect 374 470 380 471
rect 374 466 375 470
rect 379 466 380 470
rect 374 465 380 466
rect 438 470 444 471
rect 438 466 439 470
rect 443 466 444 470
rect 438 465 444 466
rect 510 470 516 471
rect 510 466 511 470
rect 515 466 516 470
rect 510 465 516 466
rect 590 470 596 471
rect 590 466 591 470
rect 595 466 596 470
rect 590 465 596 466
rect 662 470 668 471
rect 662 466 663 470
rect 667 466 668 470
rect 662 465 668 466
rect 734 470 740 471
rect 734 466 735 470
rect 739 466 740 470
rect 734 465 740 466
rect 806 470 812 471
rect 806 466 807 470
rect 811 466 812 470
rect 806 465 812 466
rect 878 470 884 471
rect 878 466 879 470
rect 883 466 884 470
rect 878 465 884 466
rect 950 470 956 471
rect 950 466 951 470
rect 955 466 956 470
rect 950 465 956 466
rect 1022 470 1028 471
rect 1022 466 1023 470
rect 1027 466 1028 470
rect 1022 465 1028 466
rect 1102 470 1108 471
rect 1102 466 1103 470
rect 1107 466 1108 470
rect 1550 470 1551 474
rect 1555 470 1556 474
rect 1550 469 1556 470
rect 1614 474 1620 475
rect 1614 470 1615 474
rect 1619 470 1620 474
rect 1614 469 1620 470
rect 1686 474 1692 475
rect 1686 470 1687 474
rect 1691 470 1692 474
rect 1686 469 1692 470
rect 1766 474 1772 475
rect 1766 470 1767 474
rect 1771 470 1772 474
rect 1766 469 1772 470
rect 1854 474 1860 475
rect 1854 470 1855 474
rect 1859 470 1860 474
rect 1854 469 1860 470
rect 1942 474 1948 475
rect 1942 470 1943 474
rect 1947 470 1948 474
rect 1942 469 1948 470
rect 2030 474 2036 475
rect 2030 470 2031 474
rect 2035 470 2036 474
rect 2030 469 2036 470
rect 2110 474 2116 475
rect 2110 470 2111 474
rect 2115 470 2116 474
rect 2110 469 2116 470
rect 2190 474 2196 475
rect 2190 470 2191 474
rect 2195 470 2196 474
rect 2190 469 2196 470
rect 2270 474 2276 475
rect 2270 470 2271 474
rect 2275 470 2276 474
rect 2270 469 2276 470
rect 2342 474 2348 475
rect 2342 470 2343 474
rect 2347 470 2348 474
rect 2342 469 2348 470
rect 2414 474 2420 475
rect 2414 470 2415 474
rect 2419 470 2420 474
rect 2414 469 2420 470
rect 2486 474 2492 475
rect 2486 470 2487 474
rect 2491 470 2492 474
rect 2486 469 2492 470
rect 2542 474 2548 475
rect 2542 470 2543 474
rect 2547 470 2548 474
rect 2542 469 2548 470
rect 1102 465 1108 466
rect 454 442 460 443
rect 454 438 455 442
rect 459 438 460 442
rect 454 437 460 438
rect 510 442 516 443
rect 510 438 511 442
rect 515 438 516 442
rect 510 437 516 438
rect 574 442 580 443
rect 574 438 575 442
rect 579 438 580 442
rect 574 437 580 438
rect 646 442 652 443
rect 646 438 647 442
rect 651 438 652 442
rect 646 437 652 438
rect 726 442 732 443
rect 726 438 727 442
rect 731 438 732 442
rect 726 437 732 438
rect 798 442 804 443
rect 798 438 799 442
rect 803 438 804 442
rect 798 437 804 438
rect 870 442 876 443
rect 870 438 871 442
rect 875 438 876 442
rect 870 437 876 438
rect 942 442 948 443
rect 942 438 943 442
rect 947 438 948 442
rect 942 437 948 438
rect 1014 442 1020 443
rect 1014 438 1015 442
rect 1019 438 1020 442
rect 1014 437 1020 438
rect 1086 442 1092 443
rect 1086 438 1087 442
rect 1091 438 1092 442
rect 1086 437 1092 438
rect 1158 442 1164 443
rect 1158 438 1159 442
rect 1163 438 1164 442
rect 1158 437 1164 438
rect 1238 442 1244 443
rect 1238 438 1239 442
rect 1243 438 1244 442
rect 1238 437 1244 438
rect 1646 442 1652 443
rect 1646 438 1647 442
rect 1651 438 1652 442
rect 1646 437 1652 438
rect 1702 442 1708 443
rect 1702 438 1703 442
rect 1707 438 1708 442
rect 1702 437 1708 438
rect 1758 442 1764 443
rect 1758 438 1759 442
rect 1763 438 1764 442
rect 1758 437 1764 438
rect 1814 442 1820 443
rect 1814 438 1815 442
rect 1819 438 1820 442
rect 1814 437 1820 438
rect 1870 442 1876 443
rect 1870 438 1871 442
rect 1875 438 1876 442
rect 1870 437 1876 438
rect 1926 442 1932 443
rect 1926 438 1927 442
rect 1931 438 1932 442
rect 1926 437 1932 438
rect 1998 442 2004 443
rect 1998 438 1999 442
rect 2003 438 2004 442
rect 1998 437 2004 438
rect 2086 442 2092 443
rect 2086 438 2087 442
rect 2091 438 2092 442
rect 2086 437 2092 438
rect 2190 442 2196 443
rect 2190 438 2191 442
rect 2195 438 2196 442
rect 2190 437 2196 438
rect 2310 442 2316 443
rect 2310 438 2311 442
rect 2315 438 2316 442
rect 2310 437 2316 438
rect 2438 442 2444 443
rect 2438 438 2439 442
rect 2443 438 2444 442
rect 2438 437 2444 438
rect 2542 442 2548 443
rect 2542 438 2543 442
rect 2547 438 2548 442
rect 2542 437 2548 438
rect 110 433 116 434
rect 110 429 111 433
rect 115 429 116 433
rect 110 428 116 429
rect 1326 433 1332 434
rect 1326 429 1327 433
rect 1331 429 1332 433
rect 1326 428 1332 429
rect 1366 433 1372 434
rect 1366 429 1367 433
rect 1371 429 1372 433
rect 1366 428 1372 429
rect 2582 433 2588 434
rect 2582 429 2583 433
rect 2587 429 2588 433
rect 2582 428 2588 429
rect 110 416 116 417
rect 1326 416 1332 417
rect 110 412 111 416
rect 115 412 116 416
rect 110 411 116 412
rect 438 415 444 416
rect 438 411 439 415
rect 443 411 444 415
rect 438 410 444 411
rect 494 415 500 416
rect 494 411 495 415
rect 499 411 500 415
rect 494 410 500 411
rect 558 415 564 416
rect 558 411 559 415
rect 563 411 564 415
rect 558 410 564 411
rect 630 415 636 416
rect 630 411 631 415
rect 635 411 636 415
rect 630 410 636 411
rect 710 415 716 416
rect 710 411 711 415
rect 715 411 716 415
rect 710 410 716 411
rect 782 415 788 416
rect 782 411 783 415
rect 787 411 788 415
rect 782 410 788 411
rect 854 415 860 416
rect 854 411 855 415
rect 859 411 860 415
rect 854 410 860 411
rect 926 415 932 416
rect 926 411 927 415
rect 931 411 932 415
rect 926 410 932 411
rect 998 415 1004 416
rect 998 411 999 415
rect 1003 411 1004 415
rect 998 410 1004 411
rect 1070 415 1076 416
rect 1070 411 1071 415
rect 1075 411 1076 415
rect 1070 410 1076 411
rect 1142 415 1148 416
rect 1142 411 1143 415
rect 1147 411 1148 415
rect 1142 410 1148 411
rect 1222 415 1228 416
rect 1222 411 1223 415
rect 1227 411 1228 415
rect 1326 412 1327 416
rect 1331 412 1332 416
rect 1326 411 1332 412
rect 1366 416 1372 417
rect 2582 416 2588 417
rect 1366 412 1367 416
rect 1371 412 1372 416
rect 1366 411 1372 412
rect 1630 415 1636 416
rect 1630 411 1631 415
rect 1635 411 1636 415
rect 1222 410 1228 411
rect 1630 410 1636 411
rect 1686 415 1692 416
rect 1686 411 1687 415
rect 1691 411 1692 415
rect 1686 410 1692 411
rect 1742 415 1748 416
rect 1742 411 1743 415
rect 1747 411 1748 415
rect 1742 410 1748 411
rect 1798 415 1804 416
rect 1798 411 1799 415
rect 1803 411 1804 415
rect 1798 410 1804 411
rect 1854 415 1860 416
rect 1854 411 1855 415
rect 1859 411 1860 415
rect 1854 410 1860 411
rect 1910 415 1916 416
rect 1910 411 1911 415
rect 1915 411 1916 415
rect 1910 410 1916 411
rect 1982 415 1988 416
rect 1982 411 1983 415
rect 1987 411 1988 415
rect 1982 410 1988 411
rect 2070 415 2076 416
rect 2070 411 2071 415
rect 2075 411 2076 415
rect 2070 410 2076 411
rect 2174 415 2180 416
rect 2174 411 2175 415
rect 2179 411 2180 415
rect 2174 410 2180 411
rect 2294 415 2300 416
rect 2294 411 2295 415
rect 2299 411 2300 415
rect 2294 410 2300 411
rect 2422 415 2428 416
rect 2422 411 2423 415
rect 2427 411 2428 415
rect 2422 410 2428 411
rect 2526 415 2532 416
rect 2526 411 2527 415
rect 2531 411 2532 415
rect 2582 412 2583 416
rect 2587 412 2588 416
rect 2582 411 2588 412
rect 2526 410 2532 411
rect 1654 381 1660 382
rect 1366 380 1372 381
rect 414 377 420 378
rect 110 376 116 377
rect 110 372 111 376
rect 115 372 116 376
rect 414 373 415 377
rect 419 373 420 377
rect 414 372 420 373
rect 470 377 476 378
rect 470 373 471 377
rect 475 373 476 377
rect 470 372 476 373
rect 534 377 540 378
rect 534 373 535 377
rect 539 373 540 377
rect 534 372 540 373
rect 606 377 612 378
rect 606 373 607 377
rect 611 373 612 377
rect 606 372 612 373
rect 686 377 692 378
rect 686 373 687 377
rect 691 373 692 377
rect 686 372 692 373
rect 766 377 772 378
rect 766 373 767 377
rect 771 373 772 377
rect 766 372 772 373
rect 846 377 852 378
rect 846 373 847 377
rect 851 373 852 377
rect 846 372 852 373
rect 926 377 932 378
rect 926 373 927 377
rect 931 373 932 377
rect 926 372 932 373
rect 1006 377 1012 378
rect 1006 373 1007 377
rect 1011 373 1012 377
rect 1006 372 1012 373
rect 1086 377 1092 378
rect 1086 373 1087 377
rect 1091 373 1092 377
rect 1086 372 1092 373
rect 1174 377 1180 378
rect 1174 373 1175 377
rect 1179 373 1180 377
rect 1174 372 1180 373
rect 1262 377 1268 378
rect 1262 373 1263 377
rect 1267 373 1268 377
rect 1262 372 1268 373
rect 1326 376 1332 377
rect 1326 372 1327 376
rect 1331 372 1332 376
rect 1366 376 1367 380
rect 1371 376 1372 380
rect 1654 377 1655 381
rect 1659 377 1660 381
rect 1654 376 1660 377
rect 1710 381 1716 382
rect 1710 377 1711 381
rect 1715 377 1716 381
rect 1710 376 1716 377
rect 1766 381 1772 382
rect 1766 377 1767 381
rect 1771 377 1772 381
rect 1766 376 1772 377
rect 1822 381 1828 382
rect 1822 377 1823 381
rect 1827 377 1828 381
rect 1822 376 1828 377
rect 1878 381 1884 382
rect 1878 377 1879 381
rect 1883 377 1884 381
rect 1878 376 1884 377
rect 1950 381 1956 382
rect 1950 377 1951 381
rect 1955 377 1956 381
rect 1950 376 1956 377
rect 2038 381 2044 382
rect 2038 377 2039 381
rect 2043 377 2044 381
rect 2038 376 2044 377
rect 2150 381 2156 382
rect 2150 377 2151 381
rect 2155 377 2156 381
rect 2150 376 2156 377
rect 2278 381 2284 382
rect 2278 377 2279 381
rect 2283 377 2284 381
rect 2278 376 2284 377
rect 2414 381 2420 382
rect 2414 377 2415 381
rect 2419 377 2420 381
rect 2414 376 2420 377
rect 2526 381 2532 382
rect 2526 377 2527 381
rect 2531 377 2532 381
rect 2526 376 2532 377
rect 2582 380 2588 381
rect 2582 376 2583 380
rect 2587 376 2588 380
rect 1366 375 1372 376
rect 2582 375 2588 376
rect 110 371 116 372
rect 1326 371 1332 372
rect 1366 363 1372 364
rect 110 359 116 360
rect 110 355 111 359
rect 115 355 116 359
rect 110 354 116 355
rect 1326 359 1332 360
rect 1326 355 1327 359
rect 1331 355 1332 359
rect 1366 359 1367 363
rect 1371 359 1372 363
rect 1366 358 1372 359
rect 2582 363 2588 364
rect 2582 359 2583 363
rect 2587 359 2588 363
rect 2582 358 2588 359
rect 1326 354 1332 355
rect 1670 354 1676 355
rect 430 350 436 351
rect 430 346 431 350
rect 435 346 436 350
rect 430 345 436 346
rect 486 350 492 351
rect 486 346 487 350
rect 491 346 492 350
rect 486 345 492 346
rect 550 350 556 351
rect 550 346 551 350
rect 555 346 556 350
rect 550 345 556 346
rect 622 350 628 351
rect 622 346 623 350
rect 627 346 628 350
rect 622 345 628 346
rect 702 350 708 351
rect 702 346 703 350
rect 707 346 708 350
rect 702 345 708 346
rect 782 350 788 351
rect 782 346 783 350
rect 787 346 788 350
rect 782 345 788 346
rect 862 350 868 351
rect 862 346 863 350
rect 867 346 868 350
rect 862 345 868 346
rect 942 350 948 351
rect 942 346 943 350
rect 947 346 948 350
rect 942 345 948 346
rect 1022 350 1028 351
rect 1022 346 1023 350
rect 1027 346 1028 350
rect 1022 345 1028 346
rect 1102 350 1108 351
rect 1102 346 1103 350
rect 1107 346 1108 350
rect 1102 345 1108 346
rect 1190 350 1196 351
rect 1190 346 1191 350
rect 1195 346 1196 350
rect 1190 345 1196 346
rect 1278 350 1284 351
rect 1278 346 1279 350
rect 1283 346 1284 350
rect 1670 350 1671 354
rect 1675 350 1676 354
rect 1670 349 1676 350
rect 1726 354 1732 355
rect 1726 350 1727 354
rect 1731 350 1732 354
rect 1726 349 1732 350
rect 1782 354 1788 355
rect 1782 350 1783 354
rect 1787 350 1788 354
rect 1782 349 1788 350
rect 1838 354 1844 355
rect 1838 350 1839 354
rect 1843 350 1844 354
rect 1838 349 1844 350
rect 1894 354 1900 355
rect 1894 350 1895 354
rect 1899 350 1900 354
rect 1894 349 1900 350
rect 1966 354 1972 355
rect 1966 350 1967 354
rect 1971 350 1972 354
rect 1966 349 1972 350
rect 2054 354 2060 355
rect 2054 350 2055 354
rect 2059 350 2060 354
rect 2054 349 2060 350
rect 2166 354 2172 355
rect 2166 350 2167 354
rect 2171 350 2172 354
rect 2166 349 2172 350
rect 2294 354 2300 355
rect 2294 350 2295 354
rect 2299 350 2300 354
rect 2294 349 2300 350
rect 2430 354 2436 355
rect 2430 350 2431 354
rect 2435 350 2436 354
rect 2430 349 2436 350
rect 2542 354 2548 355
rect 2542 350 2543 354
rect 2547 350 2548 354
rect 2542 349 2548 350
rect 1278 345 1284 346
rect 462 322 468 323
rect 462 318 463 322
rect 467 318 468 322
rect 462 317 468 318
rect 518 322 524 323
rect 518 318 519 322
rect 523 318 524 322
rect 518 317 524 318
rect 574 322 580 323
rect 574 318 575 322
rect 579 318 580 322
rect 574 317 580 318
rect 630 322 636 323
rect 630 318 631 322
rect 635 318 636 322
rect 630 317 636 318
rect 694 322 700 323
rect 694 318 695 322
rect 699 318 700 322
rect 694 317 700 318
rect 766 322 772 323
rect 766 318 767 322
rect 771 318 772 322
rect 766 317 772 318
rect 846 322 852 323
rect 846 318 847 322
rect 851 318 852 322
rect 846 317 852 318
rect 926 322 932 323
rect 926 318 927 322
rect 931 318 932 322
rect 926 317 932 318
rect 1014 322 1020 323
rect 1014 318 1015 322
rect 1019 318 1020 322
rect 1014 317 1020 318
rect 1110 322 1116 323
rect 1110 318 1111 322
rect 1115 318 1116 322
rect 1110 317 1116 318
rect 1214 322 1220 323
rect 1214 318 1215 322
rect 1219 318 1220 322
rect 1214 317 1220 318
rect 1630 322 1636 323
rect 1630 318 1631 322
rect 1635 318 1636 322
rect 1630 317 1636 318
rect 1686 322 1692 323
rect 1686 318 1687 322
rect 1691 318 1692 322
rect 1686 317 1692 318
rect 1742 322 1748 323
rect 1742 318 1743 322
rect 1747 318 1748 322
rect 1742 317 1748 318
rect 1806 322 1812 323
rect 1806 318 1807 322
rect 1811 318 1812 322
rect 1806 317 1812 318
rect 1886 322 1892 323
rect 1886 318 1887 322
rect 1891 318 1892 322
rect 1886 317 1892 318
rect 1966 322 1972 323
rect 1966 318 1967 322
rect 1971 318 1972 322
rect 1966 317 1972 318
rect 2054 322 2060 323
rect 2054 318 2055 322
rect 2059 318 2060 322
rect 2054 317 2060 318
rect 2142 322 2148 323
rect 2142 318 2143 322
rect 2147 318 2148 322
rect 2142 317 2148 318
rect 2230 322 2236 323
rect 2230 318 2231 322
rect 2235 318 2236 322
rect 2230 317 2236 318
rect 2310 322 2316 323
rect 2310 318 2311 322
rect 2315 318 2316 322
rect 2310 317 2316 318
rect 2390 322 2396 323
rect 2390 318 2391 322
rect 2395 318 2396 322
rect 2390 317 2396 318
rect 2478 322 2484 323
rect 2478 318 2479 322
rect 2483 318 2484 322
rect 2478 317 2484 318
rect 2542 322 2548 323
rect 2542 318 2543 322
rect 2547 318 2548 322
rect 2542 317 2548 318
rect 110 313 116 314
rect 110 309 111 313
rect 115 309 116 313
rect 110 308 116 309
rect 1326 313 1332 314
rect 1326 309 1327 313
rect 1331 309 1332 313
rect 1326 308 1332 309
rect 1366 313 1372 314
rect 1366 309 1367 313
rect 1371 309 1372 313
rect 1366 308 1372 309
rect 2582 313 2588 314
rect 2582 309 2583 313
rect 2587 309 2588 313
rect 2582 308 2588 309
rect 110 296 116 297
rect 1326 296 1332 297
rect 110 292 111 296
rect 115 292 116 296
rect 110 291 116 292
rect 446 295 452 296
rect 446 291 447 295
rect 451 291 452 295
rect 446 290 452 291
rect 502 295 508 296
rect 502 291 503 295
rect 507 291 508 295
rect 502 290 508 291
rect 558 295 564 296
rect 558 291 559 295
rect 563 291 564 295
rect 558 290 564 291
rect 614 295 620 296
rect 614 291 615 295
rect 619 291 620 295
rect 614 290 620 291
rect 678 295 684 296
rect 678 291 679 295
rect 683 291 684 295
rect 678 290 684 291
rect 750 295 756 296
rect 750 291 751 295
rect 755 291 756 295
rect 750 290 756 291
rect 830 295 836 296
rect 830 291 831 295
rect 835 291 836 295
rect 830 290 836 291
rect 910 295 916 296
rect 910 291 911 295
rect 915 291 916 295
rect 910 290 916 291
rect 998 295 1004 296
rect 998 291 999 295
rect 1003 291 1004 295
rect 998 290 1004 291
rect 1094 295 1100 296
rect 1094 291 1095 295
rect 1099 291 1100 295
rect 1094 290 1100 291
rect 1198 295 1204 296
rect 1198 291 1199 295
rect 1203 291 1204 295
rect 1326 292 1327 296
rect 1331 292 1332 296
rect 1326 291 1332 292
rect 1366 296 1372 297
rect 2582 296 2588 297
rect 1366 292 1367 296
rect 1371 292 1372 296
rect 1366 291 1372 292
rect 1614 295 1620 296
rect 1614 291 1615 295
rect 1619 291 1620 295
rect 1198 290 1204 291
rect 1614 290 1620 291
rect 1670 295 1676 296
rect 1670 291 1671 295
rect 1675 291 1676 295
rect 1670 290 1676 291
rect 1726 295 1732 296
rect 1726 291 1727 295
rect 1731 291 1732 295
rect 1726 290 1732 291
rect 1790 295 1796 296
rect 1790 291 1791 295
rect 1795 291 1796 295
rect 1790 290 1796 291
rect 1870 295 1876 296
rect 1870 291 1871 295
rect 1875 291 1876 295
rect 1870 290 1876 291
rect 1950 295 1956 296
rect 1950 291 1951 295
rect 1955 291 1956 295
rect 1950 290 1956 291
rect 2038 295 2044 296
rect 2038 291 2039 295
rect 2043 291 2044 295
rect 2038 290 2044 291
rect 2126 295 2132 296
rect 2126 291 2127 295
rect 2131 291 2132 295
rect 2126 290 2132 291
rect 2214 295 2220 296
rect 2214 291 2215 295
rect 2219 291 2220 295
rect 2214 290 2220 291
rect 2294 295 2300 296
rect 2294 291 2295 295
rect 2299 291 2300 295
rect 2294 290 2300 291
rect 2374 295 2380 296
rect 2374 291 2375 295
rect 2379 291 2380 295
rect 2374 290 2380 291
rect 2462 295 2468 296
rect 2462 291 2463 295
rect 2467 291 2468 295
rect 2462 290 2468 291
rect 2526 295 2532 296
rect 2526 291 2527 295
rect 2531 291 2532 295
rect 2582 292 2583 296
rect 2587 292 2588 296
rect 2582 291 2588 292
rect 2526 290 2532 291
rect 1534 261 1540 262
rect 1366 260 1372 261
rect 286 257 292 258
rect 110 256 116 257
rect 110 252 111 256
rect 115 252 116 256
rect 286 253 287 257
rect 291 253 292 257
rect 286 252 292 253
rect 358 257 364 258
rect 358 253 359 257
rect 363 253 364 257
rect 358 252 364 253
rect 438 257 444 258
rect 438 253 439 257
rect 443 253 444 257
rect 438 252 444 253
rect 526 257 532 258
rect 526 253 527 257
rect 531 253 532 257
rect 526 252 532 253
rect 622 257 628 258
rect 622 253 623 257
rect 627 253 628 257
rect 622 252 628 253
rect 718 257 724 258
rect 718 253 719 257
rect 723 253 724 257
rect 718 252 724 253
rect 822 257 828 258
rect 822 253 823 257
rect 827 253 828 257
rect 822 252 828 253
rect 926 257 932 258
rect 926 253 927 257
rect 931 253 932 257
rect 926 252 932 253
rect 1030 257 1036 258
rect 1030 253 1031 257
rect 1035 253 1036 257
rect 1030 252 1036 253
rect 1142 257 1148 258
rect 1142 253 1143 257
rect 1147 253 1148 257
rect 1142 252 1148 253
rect 1254 257 1260 258
rect 1254 253 1255 257
rect 1259 253 1260 257
rect 1254 252 1260 253
rect 1326 256 1332 257
rect 1326 252 1327 256
rect 1331 252 1332 256
rect 1366 256 1367 260
rect 1371 256 1372 260
rect 1534 257 1535 261
rect 1539 257 1540 261
rect 1534 256 1540 257
rect 1606 261 1612 262
rect 1606 257 1607 261
rect 1611 257 1612 261
rect 1606 256 1612 257
rect 1686 261 1692 262
rect 1686 257 1687 261
rect 1691 257 1692 261
rect 1686 256 1692 257
rect 1774 261 1780 262
rect 1774 257 1775 261
rect 1779 257 1780 261
rect 1774 256 1780 257
rect 1862 261 1868 262
rect 1862 257 1863 261
rect 1867 257 1868 261
rect 1862 256 1868 257
rect 1950 261 1956 262
rect 1950 257 1951 261
rect 1955 257 1956 261
rect 1950 256 1956 257
rect 2038 261 2044 262
rect 2038 257 2039 261
rect 2043 257 2044 261
rect 2038 256 2044 257
rect 2118 261 2124 262
rect 2118 257 2119 261
rect 2123 257 2124 261
rect 2118 256 2124 257
rect 2198 261 2204 262
rect 2198 257 2199 261
rect 2203 257 2204 261
rect 2198 256 2204 257
rect 2270 261 2276 262
rect 2270 257 2271 261
rect 2275 257 2276 261
rect 2270 256 2276 257
rect 2334 261 2340 262
rect 2334 257 2335 261
rect 2339 257 2340 261
rect 2334 256 2340 257
rect 2406 261 2412 262
rect 2406 257 2407 261
rect 2411 257 2412 261
rect 2406 256 2412 257
rect 2470 261 2476 262
rect 2470 257 2471 261
rect 2475 257 2476 261
rect 2470 256 2476 257
rect 2526 261 2532 262
rect 2526 257 2527 261
rect 2531 257 2532 261
rect 2526 256 2532 257
rect 2582 260 2588 261
rect 2582 256 2583 260
rect 2587 256 2588 260
rect 1366 255 1372 256
rect 2582 255 2588 256
rect 110 251 116 252
rect 1326 251 1332 252
rect 1366 243 1372 244
rect 110 239 116 240
rect 110 235 111 239
rect 115 235 116 239
rect 110 234 116 235
rect 1326 239 1332 240
rect 1326 235 1327 239
rect 1331 235 1332 239
rect 1366 239 1367 243
rect 1371 239 1372 243
rect 1366 238 1372 239
rect 2582 243 2588 244
rect 2582 239 2583 243
rect 2587 239 2588 243
rect 2582 238 2588 239
rect 1326 234 1332 235
rect 1550 234 1556 235
rect 302 230 308 231
rect 302 226 303 230
rect 307 226 308 230
rect 302 225 308 226
rect 374 230 380 231
rect 374 226 375 230
rect 379 226 380 230
rect 374 225 380 226
rect 454 230 460 231
rect 454 226 455 230
rect 459 226 460 230
rect 454 225 460 226
rect 542 230 548 231
rect 542 226 543 230
rect 547 226 548 230
rect 542 225 548 226
rect 638 230 644 231
rect 638 226 639 230
rect 643 226 644 230
rect 638 225 644 226
rect 734 230 740 231
rect 734 226 735 230
rect 739 226 740 230
rect 734 225 740 226
rect 838 230 844 231
rect 838 226 839 230
rect 843 226 844 230
rect 838 225 844 226
rect 942 230 948 231
rect 942 226 943 230
rect 947 226 948 230
rect 942 225 948 226
rect 1046 230 1052 231
rect 1046 226 1047 230
rect 1051 226 1052 230
rect 1046 225 1052 226
rect 1158 230 1164 231
rect 1158 226 1159 230
rect 1163 226 1164 230
rect 1158 225 1164 226
rect 1270 230 1276 231
rect 1270 226 1271 230
rect 1275 226 1276 230
rect 1550 230 1551 234
rect 1555 230 1556 234
rect 1550 229 1556 230
rect 1622 234 1628 235
rect 1622 230 1623 234
rect 1627 230 1628 234
rect 1622 229 1628 230
rect 1702 234 1708 235
rect 1702 230 1703 234
rect 1707 230 1708 234
rect 1702 229 1708 230
rect 1790 234 1796 235
rect 1790 230 1791 234
rect 1795 230 1796 234
rect 1790 229 1796 230
rect 1878 234 1884 235
rect 1878 230 1879 234
rect 1883 230 1884 234
rect 1878 229 1884 230
rect 1966 234 1972 235
rect 1966 230 1967 234
rect 1971 230 1972 234
rect 1966 229 1972 230
rect 2054 234 2060 235
rect 2054 230 2055 234
rect 2059 230 2060 234
rect 2054 229 2060 230
rect 2134 234 2140 235
rect 2134 230 2135 234
rect 2139 230 2140 234
rect 2134 229 2140 230
rect 2214 234 2220 235
rect 2214 230 2215 234
rect 2219 230 2220 234
rect 2214 229 2220 230
rect 2286 234 2292 235
rect 2286 230 2287 234
rect 2291 230 2292 234
rect 2286 229 2292 230
rect 2350 234 2356 235
rect 2350 230 2351 234
rect 2355 230 2356 234
rect 2350 229 2356 230
rect 2422 234 2428 235
rect 2422 230 2423 234
rect 2427 230 2428 234
rect 2422 229 2428 230
rect 2486 234 2492 235
rect 2486 230 2487 234
rect 2491 230 2492 234
rect 2486 229 2492 230
rect 2542 234 2548 235
rect 2542 230 2543 234
rect 2547 230 2548 234
rect 2542 229 2548 230
rect 1270 225 1276 226
rect 1414 210 1420 211
rect 198 206 204 207
rect 198 202 199 206
rect 203 202 204 206
rect 198 201 204 202
rect 270 206 276 207
rect 270 202 271 206
rect 275 202 276 206
rect 270 201 276 202
rect 358 206 364 207
rect 358 202 359 206
rect 363 202 364 206
rect 358 201 364 202
rect 462 206 468 207
rect 462 202 463 206
rect 467 202 468 206
rect 462 201 468 202
rect 566 206 572 207
rect 566 202 567 206
rect 571 202 572 206
rect 566 201 572 202
rect 678 206 684 207
rect 678 202 679 206
rect 683 202 684 206
rect 678 201 684 202
rect 790 206 796 207
rect 790 202 791 206
rect 795 202 796 206
rect 790 201 796 202
rect 910 206 916 207
rect 910 202 911 206
rect 915 202 916 206
rect 910 201 916 202
rect 1030 206 1036 207
rect 1030 202 1031 206
rect 1035 202 1036 206
rect 1030 201 1036 202
rect 1150 206 1156 207
rect 1150 202 1151 206
rect 1155 202 1156 206
rect 1150 201 1156 202
rect 1270 206 1276 207
rect 1270 202 1271 206
rect 1275 202 1276 206
rect 1414 206 1415 210
rect 1419 206 1420 210
rect 1414 205 1420 206
rect 1478 210 1484 211
rect 1478 206 1479 210
rect 1483 206 1484 210
rect 1478 205 1484 206
rect 1558 210 1564 211
rect 1558 206 1559 210
rect 1563 206 1564 210
rect 1558 205 1564 206
rect 1654 210 1660 211
rect 1654 206 1655 210
rect 1659 206 1660 210
rect 1654 205 1660 206
rect 1750 210 1756 211
rect 1750 206 1751 210
rect 1755 206 1756 210
rect 1750 205 1756 206
rect 1854 210 1860 211
rect 1854 206 1855 210
rect 1859 206 1860 210
rect 1854 205 1860 206
rect 1958 210 1964 211
rect 1958 206 1959 210
rect 1963 206 1964 210
rect 1958 205 1964 206
rect 2062 210 2068 211
rect 2062 206 2063 210
rect 2067 206 2068 210
rect 2062 205 2068 206
rect 2166 210 2172 211
rect 2166 206 2167 210
rect 2171 206 2172 210
rect 2166 205 2172 206
rect 2262 210 2268 211
rect 2262 206 2263 210
rect 2267 206 2268 210
rect 2262 205 2268 206
rect 2358 210 2364 211
rect 2358 206 2359 210
rect 2363 206 2364 210
rect 2358 205 2364 206
rect 2462 210 2468 211
rect 2462 206 2463 210
rect 2467 206 2468 210
rect 2462 205 2468 206
rect 2542 210 2548 211
rect 2542 206 2543 210
rect 2547 206 2548 210
rect 2542 205 2548 206
rect 1270 201 1276 202
rect 1366 201 1372 202
rect 110 197 116 198
rect 110 193 111 197
rect 115 193 116 197
rect 110 192 116 193
rect 1326 197 1332 198
rect 1326 193 1327 197
rect 1331 193 1332 197
rect 1366 197 1367 201
rect 1371 197 1372 201
rect 1366 196 1372 197
rect 2582 201 2588 202
rect 2582 197 2583 201
rect 2587 197 2588 201
rect 2582 196 2588 197
rect 1326 192 1332 193
rect 1366 184 1372 185
rect 2582 184 2588 185
rect 110 180 116 181
rect 1326 180 1332 181
rect 110 176 111 180
rect 115 176 116 180
rect 110 175 116 176
rect 182 179 188 180
rect 182 175 183 179
rect 187 175 188 179
rect 182 174 188 175
rect 254 179 260 180
rect 254 175 255 179
rect 259 175 260 179
rect 254 174 260 175
rect 342 179 348 180
rect 342 175 343 179
rect 347 175 348 179
rect 342 174 348 175
rect 446 179 452 180
rect 446 175 447 179
rect 451 175 452 179
rect 446 174 452 175
rect 550 179 556 180
rect 550 175 551 179
rect 555 175 556 179
rect 550 174 556 175
rect 662 179 668 180
rect 662 175 663 179
rect 667 175 668 179
rect 662 174 668 175
rect 774 179 780 180
rect 774 175 775 179
rect 779 175 780 179
rect 774 174 780 175
rect 894 179 900 180
rect 894 175 895 179
rect 899 175 900 179
rect 894 174 900 175
rect 1014 179 1020 180
rect 1014 175 1015 179
rect 1019 175 1020 179
rect 1014 174 1020 175
rect 1134 179 1140 180
rect 1134 175 1135 179
rect 1139 175 1140 179
rect 1134 174 1140 175
rect 1254 179 1260 180
rect 1254 175 1255 179
rect 1259 175 1260 179
rect 1326 176 1327 180
rect 1331 176 1332 180
rect 1366 180 1367 184
rect 1371 180 1372 184
rect 1366 179 1372 180
rect 1398 183 1404 184
rect 1398 179 1399 183
rect 1403 179 1404 183
rect 1398 178 1404 179
rect 1462 183 1468 184
rect 1462 179 1463 183
rect 1467 179 1468 183
rect 1462 178 1468 179
rect 1542 183 1548 184
rect 1542 179 1543 183
rect 1547 179 1548 183
rect 1542 178 1548 179
rect 1638 183 1644 184
rect 1638 179 1639 183
rect 1643 179 1644 183
rect 1638 178 1644 179
rect 1734 183 1740 184
rect 1734 179 1735 183
rect 1739 179 1740 183
rect 1734 178 1740 179
rect 1838 183 1844 184
rect 1838 179 1839 183
rect 1843 179 1844 183
rect 1838 178 1844 179
rect 1942 183 1948 184
rect 1942 179 1943 183
rect 1947 179 1948 183
rect 1942 178 1948 179
rect 2046 183 2052 184
rect 2046 179 2047 183
rect 2051 179 2052 183
rect 2046 178 2052 179
rect 2150 183 2156 184
rect 2150 179 2151 183
rect 2155 179 2156 183
rect 2150 178 2156 179
rect 2246 183 2252 184
rect 2246 179 2247 183
rect 2251 179 2252 183
rect 2246 178 2252 179
rect 2342 183 2348 184
rect 2342 179 2343 183
rect 2347 179 2348 183
rect 2342 178 2348 179
rect 2446 183 2452 184
rect 2446 179 2447 183
rect 2451 179 2452 183
rect 2446 178 2452 179
rect 2526 183 2532 184
rect 2526 179 2527 183
rect 2531 179 2532 183
rect 2582 180 2583 184
rect 2587 180 2588 184
rect 2582 179 2588 180
rect 2526 178 2532 179
rect 1326 175 1332 176
rect 1254 174 1260 175
rect 1398 133 1404 134
rect 1366 132 1372 133
rect 1366 128 1367 132
rect 1371 128 1372 132
rect 1398 129 1399 133
rect 1403 129 1404 133
rect 1398 128 1404 129
rect 1454 133 1460 134
rect 1454 129 1455 133
rect 1459 129 1460 133
rect 1454 128 1460 129
rect 1510 133 1516 134
rect 1510 129 1511 133
rect 1515 129 1516 133
rect 1510 128 1516 129
rect 1566 133 1572 134
rect 1566 129 1567 133
rect 1571 129 1572 133
rect 1566 128 1572 129
rect 1630 133 1636 134
rect 1630 129 1631 133
rect 1635 129 1636 133
rect 1630 128 1636 129
rect 1710 133 1716 134
rect 1710 129 1711 133
rect 1715 129 1716 133
rect 1710 128 1716 129
rect 1790 133 1796 134
rect 1790 129 1791 133
rect 1795 129 1796 133
rect 1790 128 1796 129
rect 1870 133 1876 134
rect 1870 129 1871 133
rect 1875 129 1876 133
rect 1870 128 1876 129
rect 1942 133 1948 134
rect 1942 129 1943 133
rect 1947 129 1948 133
rect 1942 128 1948 129
rect 2014 133 2020 134
rect 2014 129 2015 133
rect 2019 129 2020 133
rect 2014 128 2020 129
rect 2078 133 2084 134
rect 2078 129 2079 133
rect 2083 129 2084 133
rect 2078 128 2084 129
rect 2142 133 2148 134
rect 2142 129 2143 133
rect 2147 129 2148 133
rect 2142 128 2148 129
rect 2206 133 2212 134
rect 2206 129 2207 133
rect 2211 129 2212 133
rect 2206 128 2212 129
rect 2270 133 2276 134
rect 2270 129 2271 133
rect 2275 129 2276 133
rect 2270 128 2276 129
rect 2342 133 2348 134
rect 2342 129 2343 133
rect 2347 129 2348 133
rect 2342 128 2348 129
rect 2414 133 2420 134
rect 2414 129 2415 133
rect 2419 129 2420 133
rect 2414 128 2420 129
rect 2582 132 2588 133
rect 2582 128 2583 132
rect 2587 128 2588 132
rect 1366 127 1372 128
rect 2582 127 2588 128
rect 142 121 148 122
rect 110 120 116 121
rect 110 116 111 120
rect 115 116 116 120
rect 142 117 143 121
rect 147 117 148 121
rect 142 116 148 117
rect 198 121 204 122
rect 198 117 199 121
rect 203 117 204 121
rect 198 116 204 117
rect 254 121 260 122
rect 254 117 255 121
rect 259 117 260 121
rect 254 116 260 117
rect 310 121 316 122
rect 310 117 311 121
rect 315 117 316 121
rect 310 116 316 117
rect 366 121 372 122
rect 366 117 367 121
rect 371 117 372 121
rect 366 116 372 117
rect 422 121 428 122
rect 422 117 423 121
rect 427 117 428 121
rect 422 116 428 117
rect 478 121 484 122
rect 478 117 479 121
rect 483 117 484 121
rect 478 116 484 117
rect 534 121 540 122
rect 534 117 535 121
rect 539 117 540 121
rect 534 116 540 117
rect 590 121 596 122
rect 590 117 591 121
rect 595 117 596 121
rect 590 116 596 117
rect 646 121 652 122
rect 646 117 647 121
rect 651 117 652 121
rect 646 116 652 117
rect 702 121 708 122
rect 702 117 703 121
rect 707 117 708 121
rect 702 116 708 117
rect 758 121 764 122
rect 758 117 759 121
rect 763 117 764 121
rect 758 116 764 117
rect 822 121 828 122
rect 822 117 823 121
rect 827 117 828 121
rect 822 116 828 117
rect 886 121 892 122
rect 886 117 887 121
rect 891 117 892 121
rect 886 116 892 117
rect 950 121 956 122
rect 950 117 951 121
rect 955 117 956 121
rect 950 116 956 117
rect 1014 121 1020 122
rect 1014 117 1015 121
rect 1019 117 1020 121
rect 1014 116 1020 117
rect 1078 121 1084 122
rect 1078 117 1079 121
rect 1083 117 1084 121
rect 1078 116 1084 117
rect 1150 121 1156 122
rect 1150 117 1151 121
rect 1155 117 1156 121
rect 1150 116 1156 117
rect 1214 121 1220 122
rect 1214 117 1215 121
rect 1219 117 1220 121
rect 1214 116 1220 117
rect 1270 121 1276 122
rect 1270 117 1271 121
rect 1275 117 1276 121
rect 1270 116 1276 117
rect 1326 120 1332 121
rect 1326 116 1327 120
rect 1331 116 1332 120
rect 110 115 116 116
rect 1326 115 1332 116
rect 1366 115 1372 116
rect 1366 111 1367 115
rect 1371 111 1372 115
rect 1366 110 1372 111
rect 2582 115 2588 116
rect 2582 111 2583 115
rect 2587 111 2588 115
rect 2582 110 2588 111
rect 1414 106 1420 107
rect 110 103 116 104
rect 110 99 111 103
rect 115 99 116 103
rect 110 98 116 99
rect 1326 103 1332 104
rect 1326 99 1327 103
rect 1331 99 1332 103
rect 1414 102 1415 106
rect 1419 102 1420 106
rect 1414 101 1420 102
rect 1470 106 1476 107
rect 1470 102 1471 106
rect 1475 102 1476 106
rect 1470 101 1476 102
rect 1526 106 1532 107
rect 1526 102 1527 106
rect 1531 102 1532 106
rect 1526 101 1532 102
rect 1582 106 1588 107
rect 1582 102 1583 106
rect 1587 102 1588 106
rect 1582 101 1588 102
rect 1646 106 1652 107
rect 1646 102 1647 106
rect 1651 102 1652 106
rect 1646 101 1652 102
rect 1726 106 1732 107
rect 1726 102 1727 106
rect 1731 102 1732 106
rect 1726 101 1732 102
rect 1806 106 1812 107
rect 1806 102 1807 106
rect 1811 102 1812 106
rect 1806 101 1812 102
rect 1886 106 1892 107
rect 1886 102 1887 106
rect 1891 102 1892 106
rect 1886 101 1892 102
rect 1958 106 1964 107
rect 1958 102 1959 106
rect 1963 102 1964 106
rect 1958 101 1964 102
rect 2030 106 2036 107
rect 2030 102 2031 106
rect 2035 102 2036 106
rect 2030 101 2036 102
rect 2094 106 2100 107
rect 2094 102 2095 106
rect 2099 102 2100 106
rect 2094 101 2100 102
rect 2158 106 2164 107
rect 2158 102 2159 106
rect 2163 102 2164 106
rect 2158 101 2164 102
rect 2222 106 2228 107
rect 2222 102 2223 106
rect 2227 102 2228 106
rect 2222 101 2228 102
rect 2286 106 2292 107
rect 2286 102 2287 106
rect 2291 102 2292 106
rect 2286 101 2292 102
rect 2358 106 2364 107
rect 2358 102 2359 106
rect 2363 102 2364 106
rect 2358 101 2364 102
rect 2430 106 2436 107
rect 2430 102 2431 106
rect 2435 102 2436 106
rect 2430 101 2436 102
rect 1326 98 1332 99
rect 158 94 164 95
rect 158 90 159 94
rect 163 90 164 94
rect 158 89 164 90
rect 214 94 220 95
rect 214 90 215 94
rect 219 90 220 94
rect 214 89 220 90
rect 270 94 276 95
rect 270 90 271 94
rect 275 90 276 94
rect 270 89 276 90
rect 326 94 332 95
rect 326 90 327 94
rect 331 90 332 94
rect 326 89 332 90
rect 382 94 388 95
rect 382 90 383 94
rect 387 90 388 94
rect 382 89 388 90
rect 438 94 444 95
rect 438 90 439 94
rect 443 90 444 94
rect 438 89 444 90
rect 494 94 500 95
rect 494 90 495 94
rect 499 90 500 94
rect 494 89 500 90
rect 550 94 556 95
rect 550 90 551 94
rect 555 90 556 94
rect 550 89 556 90
rect 606 94 612 95
rect 606 90 607 94
rect 611 90 612 94
rect 606 89 612 90
rect 662 94 668 95
rect 662 90 663 94
rect 667 90 668 94
rect 662 89 668 90
rect 718 94 724 95
rect 718 90 719 94
rect 723 90 724 94
rect 718 89 724 90
rect 774 94 780 95
rect 774 90 775 94
rect 779 90 780 94
rect 774 89 780 90
rect 838 94 844 95
rect 838 90 839 94
rect 843 90 844 94
rect 838 89 844 90
rect 902 94 908 95
rect 902 90 903 94
rect 907 90 908 94
rect 902 89 908 90
rect 966 94 972 95
rect 966 90 967 94
rect 971 90 972 94
rect 966 89 972 90
rect 1030 94 1036 95
rect 1030 90 1031 94
rect 1035 90 1036 94
rect 1030 89 1036 90
rect 1094 94 1100 95
rect 1094 90 1095 94
rect 1099 90 1100 94
rect 1094 89 1100 90
rect 1166 94 1172 95
rect 1166 90 1167 94
rect 1171 90 1172 94
rect 1166 89 1172 90
rect 1230 94 1236 95
rect 1230 90 1231 94
rect 1235 90 1236 94
rect 1230 89 1236 90
rect 1286 94 1292 95
rect 1286 90 1287 94
rect 1291 90 1292 94
rect 1286 89 1292 90
<< m3c >>
rect 551 2626 555 2630
rect 607 2626 611 2630
rect 663 2626 667 2630
rect 719 2626 723 2630
rect 775 2626 779 2630
rect 1551 2622 1555 2626
rect 111 2617 115 2621
rect 1607 2622 1611 2626
rect 1663 2622 1667 2626
rect 1719 2622 1723 2626
rect 1775 2622 1779 2626
rect 1831 2622 1835 2626
rect 1887 2622 1891 2626
rect 1943 2622 1947 2626
rect 1999 2622 2003 2626
rect 2055 2622 2059 2626
rect 2111 2622 2115 2626
rect 2167 2622 2171 2626
rect 1327 2617 1331 2621
rect 1367 2613 1371 2617
rect 2583 2613 2587 2617
rect 111 2600 115 2604
rect 535 2599 539 2603
rect 591 2599 595 2603
rect 647 2599 651 2603
rect 703 2599 707 2603
rect 759 2599 763 2603
rect 1327 2600 1331 2604
rect 1367 2596 1371 2600
rect 1535 2595 1539 2599
rect 1591 2595 1595 2599
rect 1647 2595 1651 2599
rect 1703 2595 1707 2599
rect 1759 2595 1763 2599
rect 1815 2595 1819 2599
rect 1871 2595 1875 2599
rect 1927 2595 1931 2599
rect 1983 2595 1987 2599
rect 2039 2595 2043 2599
rect 2095 2595 2099 2599
rect 2151 2595 2155 2599
rect 2583 2596 2587 2600
rect 111 2564 115 2568
rect 215 2565 219 2569
rect 271 2565 275 2569
rect 327 2565 331 2569
rect 383 2565 387 2569
rect 439 2565 443 2569
rect 495 2565 499 2569
rect 551 2565 555 2569
rect 607 2565 611 2569
rect 663 2565 667 2569
rect 719 2565 723 2569
rect 775 2565 779 2569
rect 831 2565 835 2569
rect 887 2565 891 2569
rect 943 2565 947 2569
rect 999 2565 1003 2569
rect 1055 2565 1059 2569
rect 1111 2565 1115 2569
rect 1327 2564 1331 2568
rect 1367 2560 1371 2564
rect 1439 2561 1443 2565
rect 1543 2561 1547 2565
rect 1655 2561 1659 2565
rect 1767 2561 1771 2565
rect 1879 2561 1883 2565
rect 1991 2561 1995 2565
rect 2111 2561 2115 2565
rect 2231 2561 2235 2565
rect 2351 2561 2355 2565
rect 2583 2560 2587 2564
rect 111 2547 115 2551
rect 1327 2547 1331 2551
rect 1367 2543 1371 2547
rect 231 2538 235 2542
rect 287 2538 291 2542
rect 343 2538 347 2542
rect 399 2538 403 2542
rect 455 2538 459 2542
rect 511 2538 515 2542
rect 567 2538 571 2542
rect 623 2538 627 2542
rect 679 2538 683 2542
rect 735 2538 739 2542
rect 791 2538 795 2542
rect 847 2538 851 2542
rect 903 2538 907 2542
rect 959 2538 963 2542
rect 1015 2538 1019 2542
rect 1071 2538 1075 2542
rect 2583 2543 2587 2547
rect 1127 2538 1131 2542
rect 1455 2534 1459 2538
rect 1559 2534 1563 2538
rect 1671 2534 1675 2538
rect 1783 2534 1787 2538
rect 1895 2534 1899 2538
rect 2007 2534 2011 2538
rect 2127 2534 2131 2538
rect 2247 2534 2251 2538
rect 2367 2534 2371 2538
rect 367 2510 371 2514
rect 423 2510 427 2514
rect 487 2510 491 2514
rect 551 2510 555 2514
rect 615 2510 619 2514
rect 679 2510 683 2514
rect 743 2510 747 2514
rect 807 2510 811 2514
rect 871 2510 875 2514
rect 943 2510 947 2514
rect 1015 2510 1019 2514
rect 111 2501 115 2505
rect 1327 2501 1331 2505
rect 1551 2502 1555 2506
rect 1631 2502 1635 2506
rect 1719 2502 1723 2506
rect 1807 2502 1811 2506
rect 1903 2502 1907 2506
rect 1999 2502 2003 2506
rect 2095 2502 2099 2506
rect 2191 2502 2195 2506
rect 2295 2502 2299 2506
rect 2399 2502 2403 2506
rect 1367 2493 1371 2497
rect 2583 2493 2587 2497
rect 111 2484 115 2488
rect 351 2483 355 2487
rect 407 2483 411 2487
rect 471 2483 475 2487
rect 535 2483 539 2487
rect 599 2483 603 2487
rect 663 2483 667 2487
rect 727 2483 731 2487
rect 791 2483 795 2487
rect 855 2483 859 2487
rect 927 2483 931 2487
rect 999 2483 1003 2487
rect 1327 2484 1331 2488
rect 1367 2476 1371 2480
rect 1535 2475 1539 2479
rect 1615 2475 1619 2479
rect 1703 2475 1707 2479
rect 1791 2475 1795 2479
rect 1887 2475 1891 2479
rect 1983 2475 1987 2479
rect 2079 2475 2083 2479
rect 2175 2475 2179 2479
rect 2279 2475 2283 2479
rect 2383 2475 2387 2479
rect 2583 2476 2587 2480
rect 111 2444 115 2448
rect 271 2445 275 2449
rect 335 2445 339 2449
rect 399 2445 403 2449
rect 471 2445 475 2449
rect 551 2445 555 2449
rect 631 2445 635 2449
rect 711 2445 715 2449
rect 783 2445 787 2449
rect 863 2445 867 2449
rect 943 2445 947 2449
rect 1023 2445 1027 2449
rect 1327 2444 1331 2448
rect 1367 2440 1371 2444
rect 1647 2441 1651 2445
rect 1703 2441 1707 2445
rect 1767 2441 1771 2445
rect 1839 2441 1843 2445
rect 1911 2441 1915 2445
rect 1991 2441 1995 2445
rect 2079 2441 2083 2445
rect 2167 2441 2171 2445
rect 2263 2441 2267 2445
rect 2359 2441 2363 2445
rect 2455 2441 2459 2445
rect 2527 2441 2531 2445
rect 2583 2440 2587 2444
rect 111 2427 115 2431
rect 1327 2427 1331 2431
rect 1367 2423 1371 2427
rect 287 2418 291 2422
rect 351 2418 355 2422
rect 415 2418 419 2422
rect 487 2418 491 2422
rect 567 2418 571 2422
rect 647 2418 651 2422
rect 727 2418 731 2422
rect 799 2418 803 2422
rect 879 2418 883 2422
rect 959 2418 963 2422
rect 2583 2423 2587 2427
rect 1039 2418 1043 2422
rect 1663 2414 1667 2418
rect 1719 2414 1723 2418
rect 1783 2414 1787 2418
rect 1855 2414 1859 2418
rect 1927 2414 1931 2418
rect 2007 2414 2011 2418
rect 2095 2414 2099 2418
rect 2183 2414 2187 2418
rect 2279 2414 2283 2418
rect 2375 2414 2379 2418
rect 2471 2414 2475 2418
rect 2543 2414 2547 2418
rect 247 2390 251 2394
rect 335 2390 339 2394
rect 431 2390 435 2394
rect 527 2390 531 2394
rect 631 2390 635 2394
rect 727 2390 731 2394
rect 823 2390 827 2394
rect 919 2390 923 2394
rect 1015 2390 1019 2394
rect 1111 2390 1115 2394
rect 1455 2386 1459 2390
rect 111 2381 115 2385
rect 1559 2386 1563 2390
rect 1663 2386 1667 2390
rect 1759 2386 1763 2390
rect 1855 2386 1859 2390
rect 1943 2386 1947 2390
rect 2039 2386 2043 2390
rect 2135 2386 2139 2390
rect 2231 2386 2235 2390
rect 2335 2386 2339 2390
rect 2447 2386 2451 2390
rect 2543 2386 2547 2390
rect 1327 2381 1331 2385
rect 1367 2377 1371 2381
rect 2583 2377 2587 2381
rect 111 2364 115 2368
rect 231 2363 235 2367
rect 319 2363 323 2367
rect 415 2363 419 2367
rect 511 2363 515 2367
rect 615 2363 619 2367
rect 711 2363 715 2367
rect 807 2363 811 2367
rect 903 2363 907 2367
rect 999 2363 1003 2367
rect 1095 2363 1099 2367
rect 1327 2364 1331 2368
rect 1367 2360 1371 2364
rect 1439 2359 1443 2363
rect 1543 2359 1547 2363
rect 1647 2359 1651 2363
rect 1743 2359 1747 2363
rect 1839 2359 1843 2363
rect 1927 2359 1931 2363
rect 2023 2359 2027 2363
rect 2119 2359 2123 2363
rect 2215 2359 2219 2363
rect 2319 2359 2323 2363
rect 2431 2359 2435 2363
rect 2527 2359 2531 2363
rect 2583 2360 2587 2364
rect 111 2328 115 2332
rect 159 2329 163 2333
rect 263 2329 267 2333
rect 375 2329 379 2333
rect 487 2329 491 2333
rect 599 2329 603 2333
rect 711 2329 715 2333
rect 815 2329 819 2333
rect 911 2329 915 2333
rect 1007 2329 1011 2333
rect 1103 2329 1107 2333
rect 1199 2329 1203 2333
rect 1327 2328 1331 2332
rect 1367 2324 1371 2328
rect 1399 2325 1403 2329
rect 1455 2325 1459 2329
rect 1511 2325 1515 2329
rect 1567 2325 1571 2329
rect 1639 2325 1643 2329
rect 1727 2325 1731 2329
rect 1823 2325 1827 2329
rect 1943 2325 1947 2329
rect 2079 2325 2083 2329
rect 2223 2325 2227 2329
rect 2383 2325 2387 2329
rect 2527 2325 2531 2329
rect 2583 2324 2587 2328
rect 111 2311 115 2315
rect 1327 2311 1331 2315
rect 1367 2307 1371 2311
rect 175 2302 179 2306
rect 279 2302 283 2306
rect 391 2302 395 2306
rect 503 2302 507 2306
rect 615 2302 619 2306
rect 727 2302 731 2306
rect 831 2302 835 2306
rect 927 2302 931 2306
rect 1023 2302 1027 2306
rect 1119 2302 1123 2306
rect 2583 2307 2587 2311
rect 1215 2302 1219 2306
rect 1415 2298 1419 2302
rect 1471 2298 1475 2302
rect 1527 2298 1531 2302
rect 1583 2298 1587 2302
rect 1655 2298 1659 2302
rect 1743 2298 1747 2302
rect 1839 2298 1843 2302
rect 1959 2298 1963 2302
rect 2095 2298 2099 2302
rect 2239 2298 2243 2302
rect 2399 2298 2403 2302
rect 2543 2298 2547 2302
rect 159 2274 163 2278
rect 247 2274 251 2278
rect 375 2274 379 2278
rect 511 2274 515 2278
rect 639 2274 643 2278
rect 767 2274 771 2278
rect 887 2274 891 2278
rect 999 2274 1003 2278
rect 1103 2274 1107 2278
rect 1207 2274 1211 2278
rect 1287 2274 1291 2278
rect 111 2265 115 2269
rect 1327 2265 1331 2269
rect 1415 2266 1419 2270
rect 1495 2266 1499 2270
rect 1615 2266 1619 2270
rect 1735 2266 1739 2270
rect 1855 2266 1859 2270
rect 1967 2266 1971 2270
rect 2071 2266 2075 2270
rect 2167 2266 2171 2270
rect 2255 2266 2259 2270
rect 2335 2266 2339 2270
rect 2407 2266 2411 2270
rect 2487 2266 2491 2270
rect 2543 2266 2547 2270
rect 1367 2257 1371 2261
rect 2583 2257 2587 2261
rect 111 2248 115 2252
rect 143 2247 147 2251
rect 231 2247 235 2251
rect 359 2247 363 2251
rect 495 2247 499 2251
rect 623 2247 627 2251
rect 751 2247 755 2251
rect 871 2247 875 2251
rect 983 2247 987 2251
rect 1087 2247 1091 2251
rect 1191 2247 1195 2251
rect 1271 2247 1275 2251
rect 1327 2248 1331 2252
rect 1367 2240 1371 2244
rect 1399 2239 1403 2243
rect 1479 2239 1483 2243
rect 1599 2239 1603 2243
rect 1719 2239 1723 2243
rect 1839 2239 1843 2243
rect 1951 2239 1955 2243
rect 2055 2239 2059 2243
rect 2151 2239 2155 2243
rect 2239 2239 2243 2243
rect 2319 2239 2323 2243
rect 2391 2239 2395 2243
rect 2471 2239 2475 2243
rect 2527 2239 2531 2243
rect 2583 2240 2587 2244
rect 111 2204 115 2208
rect 143 2205 147 2209
rect 231 2205 235 2209
rect 359 2205 363 2209
rect 495 2205 499 2209
rect 623 2205 627 2209
rect 751 2205 755 2209
rect 871 2205 875 2209
rect 983 2205 987 2209
rect 1087 2205 1091 2209
rect 1191 2205 1195 2209
rect 1271 2205 1275 2209
rect 1327 2204 1331 2208
rect 1367 2192 1371 2196
rect 1455 2193 1459 2197
rect 1535 2193 1539 2197
rect 1631 2193 1635 2197
rect 1743 2193 1747 2197
rect 1863 2193 1867 2197
rect 1983 2193 1987 2197
rect 2095 2193 2099 2197
rect 2207 2193 2211 2197
rect 2311 2193 2315 2197
rect 2423 2193 2427 2197
rect 2527 2193 2531 2197
rect 2583 2192 2587 2196
rect 111 2187 115 2191
rect 1327 2187 1331 2191
rect 159 2178 163 2182
rect 247 2178 251 2182
rect 375 2178 379 2182
rect 511 2178 515 2182
rect 639 2178 643 2182
rect 767 2178 771 2182
rect 887 2178 891 2182
rect 999 2178 1003 2182
rect 1103 2178 1107 2182
rect 1207 2178 1211 2182
rect 1287 2178 1291 2182
rect 1367 2175 1371 2179
rect 2583 2175 2587 2179
rect 1471 2166 1475 2170
rect 1551 2166 1555 2170
rect 1647 2166 1651 2170
rect 1759 2166 1763 2170
rect 1879 2166 1883 2170
rect 1999 2166 2003 2170
rect 2111 2166 2115 2170
rect 2223 2166 2227 2170
rect 2327 2166 2331 2170
rect 2439 2166 2443 2170
rect 2543 2166 2547 2170
rect 159 2150 163 2154
rect 215 2150 219 2154
rect 311 2150 315 2154
rect 423 2150 427 2154
rect 543 2150 547 2154
rect 663 2150 667 2154
rect 775 2150 779 2154
rect 879 2150 883 2154
rect 975 2150 979 2154
rect 1071 2150 1075 2154
rect 1167 2150 1171 2154
rect 1271 2150 1275 2154
rect 111 2141 115 2145
rect 1327 2141 1331 2145
rect 1535 2142 1539 2146
rect 1631 2142 1635 2146
rect 1735 2142 1739 2146
rect 1839 2142 1843 2146
rect 1951 2142 1955 2146
rect 2055 2142 2059 2146
rect 2159 2142 2163 2146
rect 2263 2142 2267 2146
rect 2359 2142 2363 2146
rect 2463 2142 2467 2146
rect 2543 2142 2547 2146
rect 1367 2133 1371 2137
rect 2583 2133 2587 2137
rect 111 2124 115 2128
rect 143 2123 147 2127
rect 199 2123 203 2127
rect 295 2123 299 2127
rect 407 2123 411 2127
rect 527 2123 531 2127
rect 647 2123 651 2127
rect 759 2123 763 2127
rect 863 2123 867 2127
rect 959 2123 963 2127
rect 1055 2123 1059 2127
rect 1151 2123 1155 2127
rect 1255 2123 1259 2127
rect 1327 2124 1331 2128
rect 1367 2116 1371 2120
rect 1519 2115 1523 2119
rect 1615 2115 1619 2119
rect 1719 2115 1723 2119
rect 1823 2115 1827 2119
rect 1935 2115 1939 2119
rect 2039 2115 2043 2119
rect 2143 2115 2147 2119
rect 2247 2115 2251 2119
rect 2343 2115 2347 2119
rect 2447 2115 2451 2119
rect 2527 2115 2531 2119
rect 2583 2116 2587 2120
rect 111 2080 115 2084
rect 263 2081 267 2085
rect 327 2081 331 2085
rect 399 2081 403 2085
rect 479 2081 483 2085
rect 567 2081 571 2085
rect 655 2081 659 2085
rect 735 2081 739 2085
rect 815 2081 819 2085
rect 887 2081 891 2085
rect 967 2081 971 2085
rect 1047 2081 1051 2085
rect 1127 2081 1131 2085
rect 1327 2080 1331 2084
rect 1367 2080 1371 2084
rect 1431 2081 1435 2085
rect 1535 2081 1539 2085
rect 1647 2081 1651 2085
rect 1759 2081 1763 2085
rect 1863 2081 1867 2085
rect 1967 2081 1971 2085
rect 2071 2081 2075 2085
rect 2175 2081 2179 2085
rect 2271 2081 2275 2085
rect 2359 2081 2363 2085
rect 2455 2081 2459 2085
rect 2527 2081 2531 2085
rect 2583 2080 2587 2084
rect 111 2063 115 2067
rect 1327 2063 1331 2067
rect 1367 2063 1371 2067
rect 2583 2063 2587 2067
rect 279 2054 283 2058
rect 343 2054 347 2058
rect 415 2054 419 2058
rect 495 2054 499 2058
rect 583 2054 587 2058
rect 671 2054 675 2058
rect 751 2054 755 2058
rect 831 2054 835 2058
rect 903 2054 907 2058
rect 983 2054 987 2058
rect 1063 2054 1067 2058
rect 1143 2054 1147 2058
rect 1447 2054 1451 2058
rect 1551 2054 1555 2058
rect 1663 2054 1667 2058
rect 1775 2054 1779 2058
rect 1879 2054 1883 2058
rect 1983 2054 1987 2058
rect 2087 2054 2091 2058
rect 2191 2054 2195 2058
rect 2287 2054 2291 2058
rect 2375 2054 2379 2058
rect 2471 2054 2475 2058
rect 2543 2054 2547 2058
rect 1415 2030 1419 2034
rect 1503 2030 1507 2034
rect 1607 2030 1611 2034
rect 1711 2030 1715 2034
rect 1807 2030 1811 2034
rect 1903 2030 1907 2034
rect 2007 2030 2011 2034
rect 2111 2030 2115 2034
rect 2215 2030 2219 2034
rect 2327 2030 2331 2034
rect 2447 2030 2451 2034
rect 2543 2030 2547 2034
rect 415 2022 419 2026
rect 471 2022 475 2026
rect 527 2022 531 2026
rect 583 2022 587 2026
rect 639 2022 643 2026
rect 695 2022 699 2026
rect 751 2022 755 2026
rect 807 2022 811 2026
rect 863 2022 867 2026
rect 919 2022 923 2026
rect 975 2022 979 2026
rect 1031 2022 1035 2026
rect 1367 2021 1371 2025
rect 2583 2021 2587 2025
rect 111 2013 115 2017
rect 1327 2013 1331 2017
rect 1367 2004 1371 2008
rect 1399 2003 1403 2007
rect 1487 2003 1491 2007
rect 1591 2003 1595 2007
rect 1695 2003 1699 2007
rect 1791 2003 1795 2007
rect 1887 2003 1891 2007
rect 1991 2003 1995 2007
rect 2095 2003 2099 2007
rect 2199 2003 2203 2007
rect 2311 2003 2315 2007
rect 2431 2003 2435 2007
rect 2527 2003 2531 2007
rect 2583 2004 2587 2008
rect 111 1996 115 2000
rect 399 1995 403 1999
rect 455 1995 459 1999
rect 511 1995 515 1999
rect 567 1995 571 1999
rect 623 1995 627 1999
rect 679 1995 683 1999
rect 735 1995 739 1999
rect 791 1995 795 1999
rect 847 1995 851 1999
rect 903 1995 907 1999
rect 959 1995 963 1999
rect 1015 1995 1019 1999
rect 1327 1996 1331 2000
rect 1367 1968 1371 1972
rect 1399 1969 1403 1973
rect 1479 1969 1483 1973
rect 1583 1969 1587 1973
rect 1679 1969 1683 1973
rect 1767 1969 1771 1973
rect 1847 1969 1851 1973
rect 1927 1969 1931 1973
rect 2007 1969 2011 1973
rect 2087 1969 2091 1973
rect 2583 1968 2587 1972
rect 111 1956 115 1960
rect 335 1957 339 1961
rect 391 1957 395 1961
rect 447 1957 451 1961
rect 503 1957 507 1961
rect 567 1957 571 1961
rect 647 1957 651 1961
rect 743 1957 747 1961
rect 863 1957 867 1961
rect 999 1957 1003 1961
rect 1143 1957 1147 1961
rect 1271 1957 1275 1961
rect 1327 1956 1331 1960
rect 1367 1951 1371 1955
rect 2583 1951 2587 1955
rect 111 1939 115 1943
rect 1327 1939 1331 1943
rect 1415 1942 1419 1946
rect 1495 1942 1499 1946
rect 1599 1942 1603 1946
rect 1695 1942 1699 1946
rect 1783 1942 1787 1946
rect 1863 1942 1867 1946
rect 1943 1942 1947 1946
rect 2023 1942 2027 1946
rect 2103 1942 2107 1946
rect 351 1930 355 1934
rect 407 1930 411 1934
rect 463 1930 467 1934
rect 519 1930 523 1934
rect 583 1930 587 1934
rect 663 1930 667 1934
rect 759 1930 763 1934
rect 879 1930 883 1934
rect 1015 1930 1019 1934
rect 1159 1930 1163 1934
rect 1287 1930 1291 1934
rect 1719 1914 1723 1918
rect 1775 1914 1779 1918
rect 1831 1914 1835 1918
rect 1887 1914 1891 1918
rect 1943 1914 1947 1918
rect 1999 1914 2003 1918
rect 2055 1914 2059 1918
rect 2119 1914 2123 1918
rect 159 1906 163 1910
rect 231 1906 235 1910
rect 327 1906 331 1910
rect 431 1906 435 1910
rect 543 1906 547 1910
rect 655 1906 659 1910
rect 767 1906 771 1910
rect 879 1906 883 1910
rect 983 1906 987 1910
rect 1087 1906 1091 1910
rect 1199 1906 1203 1910
rect 1287 1906 1291 1910
rect 1367 1905 1371 1909
rect 2583 1905 2587 1909
rect 111 1897 115 1901
rect 1327 1897 1331 1901
rect 1367 1888 1371 1892
rect 1703 1887 1707 1891
rect 1759 1887 1763 1891
rect 1815 1887 1819 1891
rect 1871 1887 1875 1891
rect 1927 1887 1931 1891
rect 1983 1887 1987 1891
rect 2039 1887 2043 1891
rect 2103 1887 2107 1891
rect 2583 1888 2587 1892
rect 111 1880 115 1884
rect 143 1879 147 1883
rect 215 1879 219 1883
rect 311 1879 315 1883
rect 415 1879 419 1883
rect 527 1879 531 1883
rect 639 1879 643 1883
rect 751 1879 755 1883
rect 863 1879 867 1883
rect 967 1879 971 1883
rect 1071 1879 1075 1883
rect 1183 1879 1187 1883
rect 1271 1879 1275 1883
rect 1327 1880 1331 1884
rect 1367 1848 1371 1852
rect 1399 1849 1403 1853
rect 1463 1849 1467 1853
rect 1559 1849 1563 1853
rect 1655 1849 1659 1853
rect 1743 1849 1747 1853
rect 1831 1849 1835 1853
rect 1919 1849 1923 1853
rect 2007 1849 2011 1853
rect 2095 1849 2099 1853
rect 2183 1849 2187 1853
rect 2583 1848 2587 1852
rect 111 1836 115 1840
rect 143 1837 147 1841
rect 199 1837 203 1841
rect 263 1837 267 1841
rect 351 1837 355 1841
rect 439 1837 443 1841
rect 535 1837 539 1841
rect 623 1837 627 1841
rect 711 1837 715 1841
rect 791 1837 795 1841
rect 871 1837 875 1841
rect 951 1837 955 1841
rect 1039 1837 1043 1841
rect 1327 1836 1331 1840
rect 1367 1831 1371 1835
rect 2583 1831 2587 1835
rect 111 1819 115 1823
rect 1327 1819 1331 1823
rect 1415 1822 1419 1826
rect 1479 1822 1483 1826
rect 1575 1822 1579 1826
rect 1671 1822 1675 1826
rect 1759 1822 1763 1826
rect 1847 1822 1851 1826
rect 1935 1822 1939 1826
rect 2023 1822 2027 1826
rect 2111 1822 2115 1826
rect 2199 1822 2203 1826
rect 159 1810 163 1814
rect 215 1810 219 1814
rect 279 1810 283 1814
rect 367 1810 371 1814
rect 455 1810 459 1814
rect 551 1810 555 1814
rect 639 1810 643 1814
rect 727 1810 731 1814
rect 807 1810 811 1814
rect 887 1810 891 1814
rect 967 1810 971 1814
rect 1055 1810 1059 1814
rect 1415 1798 1419 1802
rect 1511 1798 1515 1802
rect 1623 1798 1627 1802
rect 1735 1798 1739 1802
rect 1839 1798 1843 1802
rect 1951 1798 1955 1802
rect 2063 1798 2067 1802
rect 2183 1798 2187 1802
rect 2303 1798 2307 1802
rect 2431 1798 2435 1802
rect 2543 1798 2547 1802
rect 1367 1789 1371 1793
rect 2583 1789 2587 1793
rect 231 1782 235 1786
rect 295 1782 299 1786
rect 367 1782 371 1786
rect 447 1782 451 1786
rect 535 1782 539 1786
rect 623 1782 627 1786
rect 711 1782 715 1786
rect 791 1782 795 1786
rect 871 1782 875 1786
rect 951 1782 955 1786
rect 1031 1782 1035 1786
rect 1119 1782 1123 1786
rect 111 1773 115 1777
rect 1327 1773 1331 1777
rect 1367 1772 1371 1776
rect 1399 1771 1403 1775
rect 1495 1771 1499 1775
rect 1607 1771 1611 1775
rect 1719 1771 1723 1775
rect 1823 1771 1827 1775
rect 1935 1771 1939 1775
rect 2047 1771 2051 1775
rect 2167 1771 2171 1775
rect 2287 1771 2291 1775
rect 2415 1771 2419 1775
rect 2527 1771 2531 1775
rect 2583 1772 2587 1776
rect 111 1756 115 1760
rect 215 1755 219 1759
rect 279 1755 283 1759
rect 351 1755 355 1759
rect 431 1755 435 1759
rect 519 1755 523 1759
rect 607 1755 611 1759
rect 695 1755 699 1759
rect 775 1755 779 1759
rect 855 1755 859 1759
rect 935 1755 939 1759
rect 1015 1755 1019 1759
rect 1103 1755 1107 1759
rect 1327 1756 1331 1760
rect 1367 1736 1371 1740
rect 1439 1737 1443 1741
rect 1519 1737 1523 1741
rect 1615 1737 1619 1741
rect 1719 1737 1723 1741
rect 1823 1737 1827 1741
rect 1927 1737 1931 1741
rect 2023 1737 2027 1741
rect 2119 1737 2123 1741
rect 2207 1737 2211 1741
rect 2287 1737 2291 1741
rect 2375 1737 2379 1741
rect 2463 1737 2467 1741
rect 2527 1737 2531 1741
rect 2583 1736 2587 1740
rect 111 1716 115 1720
rect 351 1717 355 1721
rect 407 1717 411 1721
rect 471 1717 475 1721
rect 551 1717 555 1721
rect 639 1717 643 1721
rect 727 1717 731 1721
rect 823 1717 827 1721
rect 919 1717 923 1721
rect 1015 1717 1019 1721
rect 1111 1717 1115 1721
rect 1207 1717 1211 1721
rect 1327 1716 1331 1720
rect 1367 1719 1371 1723
rect 2583 1719 2587 1723
rect 1455 1710 1459 1714
rect 1535 1710 1539 1714
rect 1631 1710 1635 1714
rect 1735 1710 1739 1714
rect 1839 1710 1843 1714
rect 1943 1710 1947 1714
rect 2039 1710 2043 1714
rect 2135 1710 2139 1714
rect 2223 1710 2227 1714
rect 2303 1710 2307 1714
rect 2391 1710 2395 1714
rect 2479 1710 2483 1714
rect 2543 1710 2547 1714
rect 111 1699 115 1703
rect 1327 1699 1331 1703
rect 367 1690 371 1694
rect 423 1690 427 1694
rect 487 1690 491 1694
rect 567 1690 571 1694
rect 655 1690 659 1694
rect 743 1690 747 1694
rect 839 1690 843 1694
rect 935 1690 939 1694
rect 1031 1690 1035 1694
rect 1127 1690 1131 1694
rect 1223 1690 1227 1694
rect 1559 1674 1563 1678
rect 1631 1674 1635 1678
rect 1711 1674 1715 1678
rect 1799 1674 1803 1678
rect 1887 1674 1891 1678
rect 1975 1674 1979 1678
rect 2063 1674 2067 1678
rect 2143 1674 2147 1678
rect 2215 1674 2219 1678
rect 2287 1674 2291 1678
rect 2351 1674 2355 1678
rect 2423 1674 2427 1678
rect 2487 1674 2491 1678
rect 2543 1674 2547 1678
rect 399 1662 403 1666
rect 455 1662 459 1666
rect 511 1662 515 1666
rect 575 1662 579 1666
rect 647 1662 651 1666
rect 727 1662 731 1666
rect 807 1662 811 1666
rect 887 1662 891 1666
rect 967 1662 971 1666
rect 1047 1662 1051 1666
rect 1135 1662 1139 1666
rect 1223 1662 1227 1666
rect 1287 1662 1291 1666
rect 1367 1665 1371 1669
rect 2583 1665 2587 1669
rect 111 1653 115 1657
rect 1327 1653 1331 1657
rect 1367 1648 1371 1652
rect 1543 1647 1547 1651
rect 1615 1647 1619 1651
rect 1695 1647 1699 1651
rect 1783 1647 1787 1651
rect 1871 1647 1875 1651
rect 1959 1647 1963 1651
rect 2047 1647 2051 1651
rect 2127 1647 2131 1651
rect 2199 1647 2203 1651
rect 2271 1647 2275 1651
rect 2335 1647 2339 1651
rect 2407 1647 2411 1651
rect 2471 1647 2475 1651
rect 2527 1647 2531 1651
rect 2583 1648 2587 1652
rect 111 1636 115 1640
rect 383 1635 387 1639
rect 439 1635 443 1639
rect 495 1635 499 1639
rect 559 1635 563 1639
rect 631 1635 635 1639
rect 711 1635 715 1639
rect 791 1635 795 1639
rect 871 1635 875 1639
rect 951 1635 955 1639
rect 1031 1635 1035 1639
rect 1119 1635 1123 1639
rect 1207 1635 1211 1639
rect 1271 1635 1275 1639
rect 1327 1636 1331 1640
rect 1367 1600 1371 1604
rect 1575 1601 1579 1605
rect 1631 1601 1635 1605
rect 1687 1601 1691 1605
rect 1751 1601 1755 1605
rect 1831 1601 1835 1605
rect 1919 1601 1923 1605
rect 2007 1601 2011 1605
rect 2103 1601 2107 1605
rect 2207 1601 2211 1605
rect 2319 1601 2323 1605
rect 2431 1601 2435 1605
rect 2527 1601 2531 1605
rect 2583 1600 2587 1604
rect 111 1584 115 1588
rect 287 1585 291 1589
rect 367 1585 371 1589
rect 455 1585 459 1589
rect 551 1585 555 1589
rect 647 1585 651 1589
rect 735 1585 739 1589
rect 823 1585 827 1589
rect 903 1585 907 1589
rect 983 1585 987 1589
rect 1063 1585 1067 1589
rect 1151 1585 1155 1589
rect 1327 1584 1331 1588
rect 1367 1583 1371 1587
rect 2583 1583 2587 1587
rect 1591 1574 1595 1578
rect 1647 1574 1651 1578
rect 1703 1574 1707 1578
rect 1767 1574 1771 1578
rect 1847 1574 1851 1578
rect 1935 1574 1939 1578
rect 2023 1574 2027 1578
rect 2119 1574 2123 1578
rect 2223 1574 2227 1578
rect 2335 1574 2339 1578
rect 2447 1574 2451 1578
rect 2543 1574 2547 1578
rect 111 1567 115 1571
rect 1327 1567 1331 1571
rect 303 1558 307 1562
rect 383 1558 387 1562
rect 471 1558 475 1562
rect 567 1558 571 1562
rect 663 1558 667 1562
rect 751 1558 755 1562
rect 839 1558 843 1562
rect 919 1558 923 1562
rect 999 1558 1003 1562
rect 1079 1558 1083 1562
rect 1167 1558 1171 1562
rect 1679 1546 1683 1550
rect 1735 1546 1739 1550
rect 1791 1546 1795 1550
rect 1855 1546 1859 1550
rect 1927 1546 1931 1550
rect 2007 1546 2011 1550
rect 2087 1546 2091 1550
rect 2167 1546 2171 1550
rect 2247 1546 2251 1550
rect 2327 1546 2331 1550
rect 2407 1546 2411 1550
rect 2487 1546 2491 1550
rect 2543 1546 2547 1550
rect 279 1534 283 1538
rect 335 1534 339 1538
rect 399 1534 403 1538
rect 471 1534 475 1538
rect 543 1534 547 1538
rect 615 1534 619 1538
rect 687 1534 691 1538
rect 759 1534 763 1538
rect 831 1534 835 1538
rect 903 1534 907 1538
rect 975 1534 979 1538
rect 1055 1534 1059 1538
rect 1367 1537 1371 1541
rect 2583 1537 2587 1541
rect 111 1525 115 1529
rect 1327 1525 1331 1529
rect 1367 1520 1371 1524
rect 1663 1519 1667 1523
rect 1719 1519 1723 1523
rect 1775 1519 1779 1523
rect 1839 1519 1843 1523
rect 1911 1519 1915 1523
rect 1991 1519 1995 1523
rect 2071 1519 2075 1523
rect 2151 1519 2155 1523
rect 2231 1519 2235 1523
rect 2311 1519 2315 1523
rect 2391 1519 2395 1523
rect 2471 1519 2475 1523
rect 2527 1519 2531 1523
rect 2583 1520 2587 1524
rect 111 1508 115 1512
rect 263 1507 267 1511
rect 319 1507 323 1511
rect 383 1507 387 1511
rect 455 1507 459 1511
rect 527 1507 531 1511
rect 599 1507 603 1511
rect 671 1507 675 1511
rect 743 1507 747 1511
rect 815 1507 819 1511
rect 887 1507 891 1511
rect 959 1507 963 1511
rect 1039 1507 1043 1511
rect 1327 1508 1331 1512
rect 1367 1476 1371 1480
rect 1519 1477 1523 1481
rect 1575 1477 1579 1481
rect 1647 1477 1651 1481
rect 1727 1477 1731 1481
rect 1807 1477 1811 1481
rect 1895 1477 1899 1481
rect 1983 1477 1987 1481
rect 2071 1477 2075 1481
rect 2151 1477 2155 1481
rect 2231 1477 2235 1481
rect 2311 1477 2315 1481
rect 2391 1477 2395 1481
rect 2471 1477 2475 1481
rect 2527 1477 2531 1481
rect 2583 1476 2587 1480
rect 111 1468 115 1472
rect 199 1469 203 1473
rect 287 1469 291 1473
rect 383 1469 387 1473
rect 487 1469 491 1473
rect 583 1469 587 1473
rect 679 1469 683 1473
rect 775 1469 779 1473
rect 863 1469 867 1473
rect 951 1469 955 1473
rect 1039 1469 1043 1473
rect 1135 1469 1139 1473
rect 1327 1468 1331 1472
rect 1367 1459 1371 1463
rect 2583 1459 2587 1463
rect 111 1451 115 1455
rect 1327 1451 1331 1455
rect 1535 1450 1539 1454
rect 1591 1450 1595 1454
rect 1663 1450 1667 1454
rect 1743 1450 1747 1454
rect 1823 1450 1827 1454
rect 1911 1450 1915 1454
rect 1999 1450 2003 1454
rect 2087 1450 2091 1454
rect 2167 1450 2171 1454
rect 2247 1450 2251 1454
rect 2327 1450 2331 1454
rect 2407 1450 2411 1454
rect 2487 1450 2491 1454
rect 2543 1450 2547 1454
rect 215 1442 219 1446
rect 303 1442 307 1446
rect 399 1442 403 1446
rect 503 1442 507 1446
rect 599 1442 603 1446
rect 695 1442 699 1446
rect 791 1442 795 1446
rect 879 1442 883 1446
rect 967 1442 971 1446
rect 1055 1442 1059 1446
rect 1151 1442 1155 1446
rect 159 1414 163 1418
rect 247 1414 251 1418
rect 343 1414 347 1418
rect 447 1414 451 1418
rect 551 1414 555 1418
rect 663 1414 667 1418
rect 767 1414 771 1418
rect 879 1414 883 1418
rect 991 1414 995 1418
rect 1103 1414 1107 1418
rect 1215 1414 1219 1418
rect 1415 1418 1419 1422
rect 1471 1418 1475 1422
rect 1535 1418 1539 1422
rect 1623 1418 1627 1422
rect 1719 1418 1723 1422
rect 1823 1418 1827 1422
rect 1927 1418 1931 1422
rect 2023 1418 2027 1422
rect 2119 1418 2123 1422
rect 2215 1418 2219 1422
rect 2303 1418 2307 1422
rect 2391 1418 2395 1422
rect 2479 1418 2483 1422
rect 2543 1418 2547 1422
rect 111 1405 115 1409
rect 1327 1405 1331 1409
rect 1367 1409 1371 1413
rect 2583 1409 2587 1413
rect 111 1388 115 1392
rect 143 1387 147 1391
rect 231 1387 235 1391
rect 327 1387 331 1391
rect 431 1387 435 1391
rect 535 1387 539 1391
rect 647 1387 651 1391
rect 751 1387 755 1391
rect 863 1387 867 1391
rect 975 1387 979 1391
rect 1087 1387 1091 1391
rect 1199 1387 1203 1391
rect 1327 1388 1331 1392
rect 1367 1392 1371 1396
rect 1399 1391 1403 1395
rect 1455 1391 1459 1395
rect 1519 1391 1523 1395
rect 1607 1391 1611 1395
rect 1703 1391 1707 1395
rect 1807 1391 1811 1395
rect 1911 1391 1915 1395
rect 2007 1391 2011 1395
rect 2103 1391 2107 1395
rect 2199 1391 2203 1395
rect 2287 1391 2291 1395
rect 2375 1391 2379 1395
rect 2463 1391 2467 1395
rect 2527 1391 2531 1395
rect 2583 1392 2587 1396
rect 111 1352 115 1356
rect 143 1353 147 1357
rect 207 1353 211 1357
rect 295 1353 299 1357
rect 399 1353 403 1357
rect 511 1353 515 1357
rect 623 1353 627 1357
rect 735 1353 739 1357
rect 847 1353 851 1357
rect 959 1353 963 1357
rect 1071 1353 1075 1357
rect 1183 1353 1187 1357
rect 1271 1353 1275 1357
rect 1327 1352 1331 1356
rect 1367 1348 1371 1352
rect 1399 1349 1403 1353
rect 1455 1349 1459 1353
rect 1543 1349 1547 1353
rect 1631 1349 1635 1353
rect 1719 1349 1723 1353
rect 1807 1349 1811 1353
rect 1887 1349 1891 1353
rect 1967 1349 1971 1353
rect 2047 1349 2051 1353
rect 2127 1349 2131 1353
rect 2207 1349 2211 1353
rect 2583 1348 2587 1352
rect 111 1335 115 1339
rect 1327 1335 1331 1339
rect 1367 1331 1371 1335
rect 159 1326 163 1330
rect 223 1326 227 1330
rect 311 1326 315 1330
rect 415 1326 419 1330
rect 527 1326 531 1330
rect 639 1326 643 1330
rect 751 1326 755 1330
rect 863 1326 867 1330
rect 975 1326 979 1330
rect 1087 1326 1091 1330
rect 1199 1326 1203 1330
rect 2583 1331 2587 1335
rect 1287 1326 1291 1330
rect 1415 1322 1419 1326
rect 1471 1322 1475 1326
rect 1559 1322 1563 1326
rect 1647 1322 1651 1326
rect 1735 1322 1739 1326
rect 1823 1322 1827 1326
rect 1903 1322 1907 1326
rect 1983 1322 1987 1326
rect 2063 1322 2067 1326
rect 2143 1322 2147 1326
rect 2223 1322 2227 1326
rect 159 1302 163 1306
rect 231 1302 235 1306
rect 327 1302 331 1306
rect 431 1302 435 1306
rect 535 1302 539 1306
rect 631 1302 635 1306
rect 727 1302 731 1306
rect 823 1302 827 1306
rect 911 1302 915 1306
rect 991 1302 995 1306
rect 1071 1302 1075 1306
rect 1151 1302 1155 1306
rect 1231 1302 1235 1306
rect 1287 1302 1291 1306
rect 111 1293 115 1297
rect 1327 1293 1331 1297
rect 1671 1294 1675 1298
rect 1767 1294 1771 1298
rect 1863 1294 1867 1298
rect 1959 1294 1963 1298
rect 2047 1294 2051 1298
rect 2135 1294 2139 1298
rect 2231 1294 2235 1298
rect 1367 1285 1371 1289
rect 2583 1285 2587 1289
rect 111 1276 115 1280
rect 143 1275 147 1279
rect 215 1275 219 1279
rect 311 1275 315 1279
rect 415 1275 419 1279
rect 519 1275 523 1279
rect 615 1275 619 1279
rect 711 1275 715 1279
rect 807 1275 811 1279
rect 895 1275 899 1279
rect 975 1275 979 1279
rect 1055 1275 1059 1279
rect 1135 1275 1139 1279
rect 1215 1275 1219 1279
rect 1271 1275 1275 1279
rect 1327 1276 1331 1280
rect 1367 1268 1371 1272
rect 1655 1267 1659 1271
rect 1751 1267 1755 1271
rect 1847 1267 1851 1271
rect 1943 1267 1947 1271
rect 2031 1267 2035 1271
rect 2119 1267 2123 1271
rect 2215 1267 2219 1271
rect 2583 1268 2587 1272
rect 111 1228 115 1232
rect 143 1229 147 1233
rect 199 1229 203 1233
rect 279 1229 283 1233
rect 359 1229 363 1233
rect 439 1229 443 1233
rect 519 1229 523 1233
rect 599 1229 603 1233
rect 671 1229 675 1233
rect 743 1229 747 1233
rect 815 1229 819 1233
rect 895 1229 899 1233
rect 1327 1228 1331 1232
rect 1367 1232 1371 1236
rect 1495 1233 1499 1237
rect 1559 1233 1563 1237
rect 1623 1233 1627 1237
rect 1687 1233 1691 1237
rect 1759 1233 1763 1237
rect 1823 1233 1827 1237
rect 1887 1233 1891 1237
rect 1951 1233 1955 1237
rect 2015 1233 2019 1237
rect 2079 1233 2083 1237
rect 2151 1233 2155 1237
rect 2223 1233 2227 1237
rect 2295 1233 2299 1237
rect 2583 1232 2587 1236
rect 111 1211 115 1215
rect 1327 1211 1331 1215
rect 1367 1215 1371 1219
rect 2583 1215 2587 1219
rect 159 1202 163 1206
rect 215 1202 219 1206
rect 295 1202 299 1206
rect 375 1202 379 1206
rect 455 1202 459 1206
rect 535 1202 539 1206
rect 615 1202 619 1206
rect 687 1202 691 1206
rect 759 1202 763 1206
rect 831 1202 835 1206
rect 911 1202 915 1206
rect 1511 1206 1515 1210
rect 1575 1206 1579 1210
rect 1639 1206 1643 1210
rect 1703 1206 1707 1210
rect 1775 1206 1779 1210
rect 1839 1206 1843 1210
rect 1903 1206 1907 1210
rect 1967 1206 1971 1210
rect 2031 1206 2035 1210
rect 2095 1206 2099 1210
rect 2167 1206 2171 1210
rect 2239 1206 2243 1210
rect 2311 1206 2315 1210
rect 159 1174 163 1178
rect 239 1174 243 1178
rect 327 1174 331 1178
rect 423 1174 427 1178
rect 511 1174 515 1178
rect 599 1174 603 1178
rect 687 1174 691 1178
rect 767 1174 771 1178
rect 839 1174 843 1178
rect 911 1174 915 1178
rect 983 1174 987 1178
rect 1063 1174 1067 1178
rect 1415 1174 1419 1178
rect 1503 1174 1507 1178
rect 1599 1174 1603 1178
rect 1703 1174 1707 1178
rect 1807 1174 1811 1178
rect 1911 1174 1915 1178
rect 2015 1174 2019 1178
rect 2111 1174 2115 1178
rect 2207 1174 2211 1178
rect 2303 1174 2307 1178
rect 2399 1174 2403 1178
rect 111 1165 115 1169
rect 1327 1165 1331 1169
rect 1367 1165 1371 1169
rect 2583 1165 2587 1169
rect 111 1148 115 1152
rect 143 1147 147 1151
rect 223 1147 227 1151
rect 311 1147 315 1151
rect 407 1147 411 1151
rect 495 1147 499 1151
rect 583 1147 587 1151
rect 671 1147 675 1151
rect 751 1147 755 1151
rect 823 1147 827 1151
rect 895 1147 899 1151
rect 967 1147 971 1151
rect 1047 1147 1051 1151
rect 1327 1148 1331 1152
rect 1367 1148 1371 1152
rect 1399 1147 1403 1151
rect 1487 1147 1491 1151
rect 1583 1147 1587 1151
rect 1687 1147 1691 1151
rect 1791 1147 1795 1151
rect 1895 1147 1899 1151
rect 1999 1147 2003 1151
rect 2095 1147 2099 1151
rect 2191 1147 2195 1151
rect 2287 1147 2291 1151
rect 2383 1147 2387 1151
rect 2583 1148 2587 1152
rect 111 1104 115 1108
rect 223 1105 227 1109
rect 319 1105 323 1109
rect 423 1105 427 1109
rect 527 1105 531 1109
rect 631 1105 635 1109
rect 727 1105 731 1109
rect 823 1105 827 1109
rect 911 1105 915 1109
rect 991 1105 995 1109
rect 1079 1105 1083 1109
rect 1167 1105 1171 1109
rect 1327 1104 1331 1108
rect 1367 1108 1371 1112
rect 1399 1109 1403 1113
rect 1479 1109 1483 1113
rect 1583 1109 1587 1113
rect 1687 1109 1691 1113
rect 1791 1109 1795 1113
rect 1887 1109 1891 1113
rect 1975 1109 1979 1113
rect 2063 1109 2067 1113
rect 2143 1109 2147 1113
rect 2215 1109 2219 1113
rect 2279 1109 2283 1113
rect 2343 1109 2347 1113
rect 2407 1109 2411 1113
rect 2471 1109 2475 1113
rect 2527 1109 2531 1113
rect 2583 1108 2587 1112
rect 111 1087 115 1091
rect 1327 1087 1331 1091
rect 1367 1091 1371 1095
rect 2583 1091 2587 1095
rect 239 1078 243 1082
rect 335 1078 339 1082
rect 439 1078 443 1082
rect 543 1078 547 1082
rect 647 1078 651 1082
rect 743 1078 747 1082
rect 839 1078 843 1082
rect 927 1078 931 1082
rect 1007 1078 1011 1082
rect 1095 1078 1099 1082
rect 1183 1078 1187 1082
rect 1415 1082 1419 1086
rect 1495 1082 1499 1086
rect 1599 1082 1603 1086
rect 1703 1082 1707 1086
rect 1807 1082 1811 1086
rect 1903 1082 1907 1086
rect 1991 1082 1995 1086
rect 2079 1082 2083 1086
rect 2159 1082 2163 1086
rect 2231 1082 2235 1086
rect 2295 1082 2299 1086
rect 2359 1082 2363 1086
rect 2423 1082 2427 1086
rect 2487 1082 2491 1086
rect 2543 1082 2547 1086
rect 311 1050 315 1054
rect 367 1050 371 1054
rect 439 1050 443 1054
rect 519 1050 523 1054
rect 607 1050 611 1054
rect 703 1050 707 1054
rect 799 1050 803 1054
rect 887 1050 891 1054
rect 975 1050 979 1054
rect 1055 1050 1059 1054
rect 1135 1050 1139 1054
rect 1223 1050 1227 1054
rect 1287 1050 1291 1054
rect 1415 1054 1419 1058
rect 1471 1054 1475 1058
rect 1535 1054 1539 1058
rect 1623 1054 1627 1058
rect 1727 1054 1731 1058
rect 1839 1054 1843 1058
rect 1951 1054 1955 1058
rect 2063 1054 2067 1058
rect 2167 1054 2171 1058
rect 2271 1054 2275 1058
rect 2367 1054 2371 1058
rect 2463 1054 2467 1058
rect 2543 1054 2547 1058
rect 111 1041 115 1045
rect 1327 1041 1331 1045
rect 1367 1045 1371 1049
rect 2583 1045 2587 1049
rect 111 1024 115 1028
rect 295 1023 299 1027
rect 351 1023 355 1027
rect 423 1023 427 1027
rect 503 1023 507 1027
rect 591 1023 595 1027
rect 687 1023 691 1027
rect 783 1023 787 1027
rect 871 1023 875 1027
rect 959 1023 963 1027
rect 1039 1023 1043 1027
rect 1119 1023 1123 1027
rect 1207 1023 1211 1027
rect 1271 1023 1275 1027
rect 1327 1024 1331 1028
rect 1367 1028 1371 1032
rect 1399 1027 1403 1031
rect 1455 1027 1459 1031
rect 1519 1027 1523 1031
rect 1607 1027 1611 1031
rect 1711 1027 1715 1031
rect 1823 1027 1827 1031
rect 1935 1027 1939 1031
rect 2047 1027 2051 1031
rect 2151 1027 2155 1031
rect 2255 1027 2259 1031
rect 2351 1027 2355 1031
rect 2447 1027 2451 1031
rect 2527 1027 2531 1031
rect 2583 1028 2587 1032
rect 111 984 115 988
rect 415 985 419 989
rect 471 985 475 989
rect 527 985 531 989
rect 591 985 595 989
rect 655 985 659 989
rect 719 985 723 989
rect 783 985 787 989
rect 847 985 851 989
rect 911 985 915 989
rect 975 985 979 989
rect 1039 985 1043 989
rect 1103 985 1107 989
rect 1159 985 1163 989
rect 1215 985 1219 989
rect 1271 985 1275 989
rect 1327 984 1331 988
rect 1367 976 1371 980
rect 1399 977 1403 981
rect 1455 977 1459 981
rect 1511 977 1515 981
rect 1567 977 1571 981
rect 1639 977 1643 981
rect 1719 977 1723 981
rect 1807 977 1811 981
rect 1903 977 1907 981
rect 2015 977 2019 981
rect 2143 977 2147 981
rect 2271 977 2275 981
rect 2407 977 2411 981
rect 2527 977 2531 981
rect 2583 976 2587 980
rect 111 967 115 971
rect 1327 967 1331 971
rect 431 958 435 962
rect 487 958 491 962
rect 543 958 547 962
rect 607 958 611 962
rect 671 958 675 962
rect 735 958 739 962
rect 799 958 803 962
rect 863 958 867 962
rect 927 958 931 962
rect 991 958 995 962
rect 1055 958 1059 962
rect 1119 958 1123 962
rect 1175 958 1179 962
rect 1231 958 1235 962
rect 1287 958 1291 962
rect 1367 959 1371 963
rect 2583 959 2587 963
rect 1415 950 1419 954
rect 1471 950 1475 954
rect 1527 950 1531 954
rect 1583 950 1587 954
rect 1655 950 1659 954
rect 1735 950 1739 954
rect 1823 950 1827 954
rect 1919 950 1923 954
rect 2031 950 2035 954
rect 2159 950 2163 954
rect 2287 950 2291 954
rect 2423 950 2427 954
rect 2543 950 2547 954
rect 423 930 427 934
rect 479 930 483 934
rect 535 930 539 934
rect 591 930 595 934
rect 647 930 651 934
rect 703 930 707 934
rect 759 930 763 934
rect 815 930 819 934
rect 111 921 115 925
rect 1327 921 1331 925
rect 1415 918 1419 922
rect 1471 918 1475 922
rect 1527 918 1531 922
rect 1615 918 1619 922
rect 1711 918 1715 922
rect 1823 918 1827 922
rect 1943 918 1947 922
rect 2063 918 2067 922
rect 2183 918 2187 922
rect 2311 918 2315 922
rect 2439 918 2443 922
rect 2543 918 2547 922
rect 1367 909 1371 913
rect 2583 909 2587 913
rect 111 904 115 908
rect 407 903 411 907
rect 463 903 467 907
rect 519 903 523 907
rect 575 903 579 907
rect 631 903 635 907
rect 687 903 691 907
rect 743 903 747 907
rect 799 903 803 907
rect 1327 904 1331 908
rect 1367 892 1371 896
rect 1399 891 1403 895
rect 1455 891 1459 895
rect 1511 891 1515 895
rect 1599 891 1603 895
rect 1695 891 1699 895
rect 1807 891 1811 895
rect 1927 891 1931 895
rect 2047 891 2051 895
rect 2167 891 2171 895
rect 2295 891 2299 895
rect 2423 891 2427 895
rect 2527 891 2531 895
rect 2583 892 2587 896
rect 111 868 115 872
rect 279 869 283 873
rect 335 869 339 873
rect 391 869 395 873
rect 455 869 459 873
rect 519 869 523 873
rect 583 869 587 873
rect 647 869 651 873
rect 711 869 715 873
rect 775 869 779 873
rect 847 869 851 873
rect 919 869 923 873
rect 1327 868 1331 872
rect 1367 856 1371 860
rect 1471 857 1475 861
rect 1551 857 1555 861
rect 1639 857 1643 861
rect 1727 857 1731 861
rect 1815 857 1819 861
rect 1903 857 1907 861
rect 1991 857 1995 861
rect 2071 857 2075 861
rect 2143 857 2147 861
rect 2215 857 2219 861
rect 2279 857 2283 861
rect 2343 857 2347 861
rect 2407 857 2411 861
rect 2471 857 2475 861
rect 2527 857 2531 861
rect 2583 856 2587 860
rect 111 851 115 855
rect 1327 851 1331 855
rect 295 842 299 846
rect 351 842 355 846
rect 407 842 411 846
rect 471 842 475 846
rect 535 842 539 846
rect 599 842 603 846
rect 663 842 667 846
rect 727 842 731 846
rect 791 842 795 846
rect 863 842 867 846
rect 935 842 939 846
rect 1367 839 1371 843
rect 2583 839 2587 843
rect 1487 830 1491 834
rect 1567 830 1571 834
rect 1655 830 1659 834
rect 1743 830 1747 834
rect 1831 830 1835 834
rect 1919 830 1923 834
rect 2007 830 2011 834
rect 2087 830 2091 834
rect 2159 830 2163 834
rect 2231 830 2235 834
rect 2295 830 2299 834
rect 2359 830 2363 834
rect 2423 830 2427 834
rect 2487 830 2491 834
rect 2543 830 2547 834
rect 167 810 171 814
rect 231 810 235 814
rect 311 810 315 814
rect 399 810 403 814
rect 487 810 491 814
rect 583 810 587 814
rect 671 810 675 814
rect 759 810 763 814
rect 839 810 843 814
rect 919 810 923 814
rect 1007 810 1011 814
rect 1095 810 1099 814
rect 111 801 115 805
rect 1327 801 1331 805
rect 1631 798 1635 802
rect 1687 798 1691 802
rect 1751 798 1755 802
rect 1823 798 1827 802
rect 1903 798 1907 802
rect 1991 798 1995 802
rect 2071 798 2075 802
rect 2159 798 2163 802
rect 2247 798 2251 802
rect 2335 798 2339 802
rect 2423 798 2427 802
rect 1367 789 1371 793
rect 2583 789 2587 793
rect 111 784 115 788
rect 151 783 155 787
rect 215 783 219 787
rect 295 783 299 787
rect 383 783 387 787
rect 471 783 475 787
rect 567 783 571 787
rect 655 783 659 787
rect 743 783 747 787
rect 823 783 827 787
rect 903 783 907 787
rect 991 783 995 787
rect 1079 783 1083 787
rect 1327 784 1331 788
rect 1367 772 1371 776
rect 1615 771 1619 775
rect 1671 771 1675 775
rect 1735 771 1739 775
rect 1807 771 1811 775
rect 1887 771 1891 775
rect 1975 771 1979 775
rect 2055 771 2059 775
rect 2143 771 2147 775
rect 2231 771 2235 775
rect 2319 771 2323 775
rect 2407 771 2411 775
rect 2583 772 2587 776
rect 111 740 115 744
rect 143 741 147 745
rect 199 741 203 745
rect 279 741 283 745
rect 383 741 387 745
rect 487 741 491 745
rect 599 741 603 745
rect 703 741 707 745
rect 807 741 811 745
rect 903 741 907 745
rect 991 741 995 745
rect 1079 741 1083 745
rect 1175 741 1179 745
rect 1327 740 1331 744
rect 1367 732 1371 736
rect 1567 733 1571 737
rect 1623 733 1627 737
rect 1687 733 1691 737
rect 1759 733 1763 737
rect 1839 733 1843 737
rect 1919 733 1923 737
rect 1999 733 2003 737
rect 2079 733 2083 737
rect 2159 733 2163 737
rect 2247 733 2251 737
rect 2335 733 2339 737
rect 2583 732 2587 736
rect 111 723 115 727
rect 1327 723 1331 727
rect 159 714 163 718
rect 215 714 219 718
rect 295 714 299 718
rect 399 714 403 718
rect 503 714 507 718
rect 615 714 619 718
rect 719 714 723 718
rect 823 714 827 718
rect 919 714 923 718
rect 1007 714 1011 718
rect 1095 714 1099 718
rect 1191 714 1195 718
rect 1367 715 1371 719
rect 2583 715 2587 719
rect 1583 706 1587 710
rect 1639 706 1643 710
rect 1703 706 1707 710
rect 1775 706 1779 710
rect 1855 706 1859 710
rect 1935 706 1939 710
rect 2015 706 2019 710
rect 2095 706 2099 710
rect 2175 706 2179 710
rect 2263 706 2267 710
rect 2351 706 2355 710
rect 159 686 163 690
rect 215 686 219 690
rect 279 686 283 690
rect 359 686 363 690
rect 447 686 451 690
rect 535 686 539 690
rect 623 686 627 690
rect 711 686 715 690
rect 791 686 795 690
rect 871 686 875 690
rect 951 686 955 690
rect 1039 686 1043 690
rect 111 677 115 681
rect 1327 677 1331 681
rect 1415 678 1419 682
rect 1511 678 1515 682
rect 1615 678 1619 682
rect 1719 678 1723 682
rect 1823 678 1827 682
rect 1927 678 1931 682
rect 2023 678 2027 682
rect 2119 678 2123 682
rect 2207 678 2211 682
rect 2295 678 2299 682
rect 2391 678 2395 682
rect 1367 669 1371 673
rect 2583 669 2587 673
rect 111 660 115 664
rect 143 659 147 663
rect 199 659 203 663
rect 263 659 267 663
rect 343 659 347 663
rect 431 659 435 663
rect 519 659 523 663
rect 607 659 611 663
rect 695 659 699 663
rect 775 659 779 663
rect 855 659 859 663
rect 935 659 939 663
rect 1023 659 1027 663
rect 1327 660 1331 664
rect 1367 652 1371 656
rect 1399 651 1403 655
rect 1495 651 1499 655
rect 1599 651 1603 655
rect 1703 651 1707 655
rect 1807 651 1811 655
rect 1911 651 1915 655
rect 2007 651 2011 655
rect 2103 651 2107 655
rect 2191 651 2195 655
rect 2279 651 2283 655
rect 2375 651 2379 655
rect 2583 652 2587 656
rect 111 616 115 620
rect 143 617 147 621
rect 199 617 203 621
rect 255 617 259 621
rect 311 617 315 621
rect 391 617 395 621
rect 479 617 483 621
rect 575 617 579 621
rect 679 617 683 621
rect 783 617 787 621
rect 887 617 891 621
rect 991 617 995 621
rect 1087 617 1091 621
rect 1191 617 1195 621
rect 1271 617 1275 621
rect 1327 616 1331 620
rect 1367 616 1371 620
rect 1399 617 1403 621
rect 1511 617 1515 621
rect 1647 617 1651 621
rect 1783 617 1787 621
rect 1911 617 1915 621
rect 2039 617 2043 621
rect 2159 617 2163 621
rect 2279 617 2283 621
rect 2407 617 2411 621
rect 2583 616 2587 620
rect 111 599 115 603
rect 1327 599 1331 603
rect 1367 599 1371 603
rect 2583 599 2587 603
rect 159 590 163 594
rect 215 590 219 594
rect 271 590 275 594
rect 327 590 331 594
rect 407 590 411 594
rect 495 590 499 594
rect 591 590 595 594
rect 695 590 699 594
rect 799 590 803 594
rect 903 590 907 594
rect 1007 590 1011 594
rect 1103 590 1107 594
rect 1207 590 1211 594
rect 1287 590 1291 594
rect 1415 590 1419 594
rect 1527 590 1531 594
rect 1663 590 1667 594
rect 1799 590 1803 594
rect 1927 590 1931 594
rect 2055 590 2059 594
rect 2175 590 2179 594
rect 2295 590 2299 594
rect 2423 590 2427 594
rect 199 562 203 566
rect 263 562 267 566
rect 335 562 339 566
rect 415 562 419 566
rect 511 562 515 566
rect 615 562 619 566
rect 719 562 723 566
rect 831 562 835 566
rect 943 562 947 566
rect 1063 562 1067 566
rect 1183 562 1187 566
rect 1287 562 1291 566
rect 1415 558 1419 562
rect 111 553 115 557
rect 1471 558 1475 562
rect 1551 558 1555 562
rect 1647 558 1651 562
rect 1751 558 1755 562
rect 1855 558 1859 562
rect 1959 558 1963 562
rect 2055 558 2059 562
rect 2151 558 2155 562
rect 2239 558 2243 562
rect 2319 558 2323 562
rect 2399 558 2403 562
rect 2479 558 2483 562
rect 2543 558 2547 562
rect 1327 553 1331 557
rect 1367 549 1371 553
rect 2583 549 2587 553
rect 111 536 115 540
rect 183 535 187 539
rect 247 535 251 539
rect 319 535 323 539
rect 399 535 403 539
rect 495 535 499 539
rect 599 535 603 539
rect 703 535 707 539
rect 815 535 819 539
rect 927 535 931 539
rect 1047 535 1051 539
rect 1167 535 1171 539
rect 1271 535 1275 539
rect 1327 536 1331 540
rect 1367 532 1371 536
rect 1399 531 1403 535
rect 1455 531 1459 535
rect 1535 531 1539 535
rect 1631 531 1635 535
rect 1735 531 1739 535
rect 1839 531 1843 535
rect 1943 531 1947 535
rect 2039 531 2043 535
rect 2135 531 2139 535
rect 2223 531 2227 535
rect 2303 531 2307 535
rect 2383 531 2387 535
rect 2463 531 2467 535
rect 2527 531 2531 535
rect 2583 532 2587 536
rect 111 492 115 496
rect 303 493 307 497
rect 359 493 363 497
rect 423 493 427 497
rect 495 493 499 497
rect 575 493 579 497
rect 647 493 651 497
rect 719 493 723 497
rect 791 493 795 497
rect 863 493 867 497
rect 935 493 939 497
rect 1007 493 1011 497
rect 1087 493 1091 497
rect 1327 492 1331 496
rect 1367 496 1371 500
rect 1535 497 1539 501
rect 1599 497 1603 501
rect 1671 497 1675 501
rect 1751 497 1755 501
rect 1839 497 1843 501
rect 1927 497 1931 501
rect 2015 497 2019 501
rect 2095 497 2099 501
rect 2175 497 2179 501
rect 2255 497 2259 501
rect 2327 497 2331 501
rect 2399 497 2403 501
rect 2471 497 2475 501
rect 2527 497 2531 501
rect 2583 496 2587 500
rect 111 475 115 479
rect 1327 475 1331 479
rect 1367 479 1371 483
rect 2583 479 2587 483
rect 319 466 323 470
rect 375 466 379 470
rect 439 466 443 470
rect 511 466 515 470
rect 591 466 595 470
rect 663 466 667 470
rect 735 466 739 470
rect 807 466 811 470
rect 879 466 883 470
rect 951 466 955 470
rect 1023 466 1027 470
rect 1103 466 1107 470
rect 1551 470 1555 474
rect 1615 470 1619 474
rect 1687 470 1691 474
rect 1767 470 1771 474
rect 1855 470 1859 474
rect 1943 470 1947 474
rect 2031 470 2035 474
rect 2111 470 2115 474
rect 2191 470 2195 474
rect 2271 470 2275 474
rect 2343 470 2347 474
rect 2415 470 2419 474
rect 2487 470 2491 474
rect 2543 470 2547 474
rect 455 438 459 442
rect 511 438 515 442
rect 575 438 579 442
rect 647 438 651 442
rect 727 438 731 442
rect 799 438 803 442
rect 871 438 875 442
rect 943 438 947 442
rect 1015 438 1019 442
rect 1087 438 1091 442
rect 1159 438 1163 442
rect 1239 438 1243 442
rect 1647 438 1651 442
rect 1703 438 1707 442
rect 1759 438 1763 442
rect 1815 438 1819 442
rect 1871 438 1875 442
rect 1927 438 1931 442
rect 1999 438 2003 442
rect 2087 438 2091 442
rect 2191 438 2195 442
rect 2311 438 2315 442
rect 2439 438 2443 442
rect 2543 438 2547 442
rect 111 429 115 433
rect 1327 429 1331 433
rect 1367 429 1371 433
rect 2583 429 2587 433
rect 111 412 115 416
rect 439 411 443 415
rect 495 411 499 415
rect 559 411 563 415
rect 631 411 635 415
rect 711 411 715 415
rect 783 411 787 415
rect 855 411 859 415
rect 927 411 931 415
rect 999 411 1003 415
rect 1071 411 1075 415
rect 1143 411 1147 415
rect 1223 411 1227 415
rect 1327 412 1331 416
rect 1367 412 1371 416
rect 1631 411 1635 415
rect 1687 411 1691 415
rect 1743 411 1747 415
rect 1799 411 1803 415
rect 1855 411 1859 415
rect 1911 411 1915 415
rect 1983 411 1987 415
rect 2071 411 2075 415
rect 2175 411 2179 415
rect 2295 411 2299 415
rect 2423 411 2427 415
rect 2527 411 2531 415
rect 2583 412 2587 416
rect 111 372 115 376
rect 415 373 419 377
rect 471 373 475 377
rect 535 373 539 377
rect 607 373 611 377
rect 687 373 691 377
rect 767 373 771 377
rect 847 373 851 377
rect 927 373 931 377
rect 1007 373 1011 377
rect 1087 373 1091 377
rect 1175 373 1179 377
rect 1263 373 1267 377
rect 1327 372 1331 376
rect 1367 376 1371 380
rect 1655 377 1659 381
rect 1711 377 1715 381
rect 1767 377 1771 381
rect 1823 377 1827 381
rect 1879 377 1883 381
rect 1951 377 1955 381
rect 2039 377 2043 381
rect 2151 377 2155 381
rect 2279 377 2283 381
rect 2415 377 2419 381
rect 2527 377 2531 381
rect 2583 376 2587 380
rect 111 355 115 359
rect 1327 355 1331 359
rect 1367 359 1371 363
rect 2583 359 2587 363
rect 431 346 435 350
rect 487 346 491 350
rect 551 346 555 350
rect 623 346 627 350
rect 703 346 707 350
rect 783 346 787 350
rect 863 346 867 350
rect 943 346 947 350
rect 1023 346 1027 350
rect 1103 346 1107 350
rect 1191 346 1195 350
rect 1279 346 1283 350
rect 1671 350 1675 354
rect 1727 350 1731 354
rect 1783 350 1787 354
rect 1839 350 1843 354
rect 1895 350 1899 354
rect 1967 350 1971 354
rect 2055 350 2059 354
rect 2167 350 2171 354
rect 2295 350 2299 354
rect 2431 350 2435 354
rect 2543 350 2547 354
rect 463 318 467 322
rect 519 318 523 322
rect 575 318 579 322
rect 631 318 635 322
rect 695 318 699 322
rect 767 318 771 322
rect 847 318 851 322
rect 927 318 931 322
rect 1015 318 1019 322
rect 1111 318 1115 322
rect 1215 318 1219 322
rect 1631 318 1635 322
rect 1687 318 1691 322
rect 1743 318 1747 322
rect 1807 318 1811 322
rect 1887 318 1891 322
rect 1967 318 1971 322
rect 2055 318 2059 322
rect 2143 318 2147 322
rect 2231 318 2235 322
rect 2311 318 2315 322
rect 2391 318 2395 322
rect 2479 318 2483 322
rect 2543 318 2547 322
rect 111 309 115 313
rect 1327 309 1331 313
rect 1367 309 1371 313
rect 2583 309 2587 313
rect 111 292 115 296
rect 447 291 451 295
rect 503 291 507 295
rect 559 291 563 295
rect 615 291 619 295
rect 679 291 683 295
rect 751 291 755 295
rect 831 291 835 295
rect 911 291 915 295
rect 999 291 1003 295
rect 1095 291 1099 295
rect 1199 291 1203 295
rect 1327 292 1331 296
rect 1367 292 1371 296
rect 1615 291 1619 295
rect 1671 291 1675 295
rect 1727 291 1731 295
rect 1791 291 1795 295
rect 1871 291 1875 295
rect 1951 291 1955 295
rect 2039 291 2043 295
rect 2127 291 2131 295
rect 2215 291 2219 295
rect 2295 291 2299 295
rect 2375 291 2379 295
rect 2463 291 2467 295
rect 2527 291 2531 295
rect 2583 292 2587 296
rect 111 252 115 256
rect 287 253 291 257
rect 359 253 363 257
rect 439 253 443 257
rect 527 253 531 257
rect 623 253 627 257
rect 719 253 723 257
rect 823 253 827 257
rect 927 253 931 257
rect 1031 253 1035 257
rect 1143 253 1147 257
rect 1255 253 1259 257
rect 1327 252 1331 256
rect 1367 256 1371 260
rect 1535 257 1539 261
rect 1607 257 1611 261
rect 1687 257 1691 261
rect 1775 257 1779 261
rect 1863 257 1867 261
rect 1951 257 1955 261
rect 2039 257 2043 261
rect 2119 257 2123 261
rect 2199 257 2203 261
rect 2271 257 2275 261
rect 2335 257 2339 261
rect 2407 257 2411 261
rect 2471 257 2475 261
rect 2527 257 2531 261
rect 2583 256 2587 260
rect 111 235 115 239
rect 1327 235 1331 239
rect 1367 239 1371 243
rect 2583 239 2587 243
rect 303 226 307 230
rect 375 226 379 230
rect 455 226 459 230
rect 543 226 547 230
rect 639 226 643 230
rect 735 226 739 230
rect 839 226 843 230
rect 943 226 947 230
rect 1047 226 1051 230
rect 1159 226 1163 230
rect 1271 226 1275 230
rect 1551 230 1555 234
rect 1623 230 1627 234
rect 1703 230 1707 234
rect 1791 230 1795 234
rect 1879 230 1883 234
rect 1967 230 1971 234
rect 2055 230 2059 234
rect 2135 230 2139 234
rect 2215 230 2219 234
rect 2287 230 2291 234
rect 2351 230 2355 234
rect 2423 230 2427 234
rect 2487 230 2491 234
rect 2543 230 2547 234
rect 199 202 203 206
rect 271 202 275 206
rect 359 202 363 206
rect 463 202 467 206
rect 567 202 571 206
rect 679 202 683 206
rect 791 202 795 206
rect 911 202 915 206
rect 1031 202 1035 206
rect 1151 202 1155 206
rect 1271 202 1275 206
rect 1415 206 1419 210
rect 1479 206 1483 210
rect 1559 206 1563 210
rect 1655 206 1659 210
rect 1751 206 1755 210
rect 1855 206 1859 210
rect 1959 206 1963 210
rect 2063 206 2067 210
rect 2167 206 2171 210
rect 2263 206 2267 210
rect 2359 206 2363 210
rect 2463 206 2467 210
rect 2543 206 2547 210
rect 111 193 115 197
rect 1327 193 1331 197
rect 1367 197 1371 201
rect 2583 197 2587 201
rect 111 176 115 180
rect 183 175 187 179
rect 255 175 259 179
rect 343 175 347 179
rect 447 175 451 179
rect 551 175 555 179
rect 663 175 667 179
rect 775 175 779 179
rect 895 175 899 179
rect 1015 175 1019 179
rect 1135 175 1139 179
rect 1255 175 1259 179
rect 1327 176 1331 180
rect 1367 180 1371 184
rect 1399 179 1403 183
rect 1463 179 1467 183
rect 1543 179 1547 183
rect 1639 179 1643 183
rect 1735 179 1739 183
rect 1839 179 1843 183
rect 1943 179 1947 183
rect 2047 179 2051 183
rect 2151 179 2155 183
rect 2247 179 2251 183
rect 2343 179 2347 183
rect 2447 179 2451 183
rect 2527 179 2531 183
rect 2583 180 2587 184
rect 1367 128 1371 132
rect 1399 129 1403 133
rect 1455 129 1459 133
rect 1511 129 1515 133
rect 1567 129 1571 133
rect 1631 129 1635 133
rect 1711 129 1715 133
rect 1791 129 1795 133
rect 1871 129 1875 133
rect 1943 129 1947 133
rect 2015 129 2019 133
rect 2079 129 2083 133
rect 2143 129 2147 133
rect 2207 129 2211 133
rect 2271 129 2275 133
rect 2343 129 2347 133
rect 2415 129 2419 133
rect 2583 128 2587 132
rect 111 116 115 120
rect 143 117 147 121
rect 199 117 203 121
rect 255 117 259 121
rect 311 117 315 121
rect 367 117 371 121
rect 423 117 427 121
rect 479 117 483 121
rect 535 117 539 121
rect 591 117 595 121
rect 647 117 651 121
rect 703 117 707 121
rect 759 117 763 121
rect 823 117 827 121
rect 887 117 891 121
rect 951 117 955 121
rect 1015 117 1019 121
rect 1079 117 1083 121
rect 1151 117 1155 121
rect 1215 117 1219 121
rect 1271 117 1275 121
rect 1327 116 1331 120
rect 1367 111 1371 115
rect 2583 111 2587 115
rect 111 99 115 103
rect 1327 99 1331 103
rect 1415 102 1419 106
rect 1471 102 1475 106
rect 1527 102 1531 106
rect 1583 102 1587 106
rect 1647 102 1651 106
rect 1727 102 1731 106
rect 1807 102 1811 106
rect 1887 102 1891 106
rect 1959 102 1963 106
rect 2031 102 2035 106
rect 2095 102 2099 106
rect 2159 102 2163 106
rect 2223 102 2227 106
rect 2287 102 2291 106
rect 2359 102 2363 106
rect 2431 102 2435 106
rect 159 90 163 94
rect 215 90 219 94
rect 271 90 275 94
rect 327 90 331 94
rect 383 90 387 94
rect 439 90 443 94
rect 495 90 499 94
rect 551 90 555 94
rect 607 90 611 94
rect 663 90 667 94
rect 719 90 723 94
rect 775 90 779 94
rect 839 90 843 94
rect 903 90 907 94
rect 967 90 971 94
rect 1031 90 1035 94
rect 1095 90 1099 94
rect 1167 90 1171 94
rect 1231 90 1235 94
rect 1287 90 1291 94
<< m3 >>
rect 111 2642 115 2643
rect 111 2637 115 2638
rect 551 2642 555 2643
rect 551 2637 555 2638
rect 607 2642 611 2643
rect 607 2637 611 2638
rect 663 2642 667 2643
rect 663 2637 667 2638
rect 719 2642 723 2643
rect 719 2637 723 2638
rect 775 2642 779 2643
rect 775 2637 779 2638
rect 1327 2642 1331 2643
rect 1327 2637 1331 2638
rect 1367 2638 1371 2639
rect 112 2622 114 2637
rect 552 2631 554 2637
rect 608 2631 610 2637
rect 664 2631 666 2637
rect 720 2631 722 2637
rect 776 2631 778 2637
rect 550 2630 556 2631
rect 550 2626 551 2630
rect 555 2626 556 2630
rect 550 2625 556 2626
rect 606 2630 612 2631
rect 606 2626 607 2630
rect 611 2626 612 2630
rect 606 2625 612 2626
rect 662 2630 668 2631
rect 662 2626 663 2630
rect 667 2626 668 2630
rect 662 2625 668 2626
rect 718 2630 724 2631
rect 718 2626 719 2630
rect 723 2626 724 2630
rect 718 2625 724 2626
rect 774 2630 780 2631
rect 774 2626 775 2630
rect 779 2626 780 2630
rect 774 2625 780 2626
rect 1328 2622 1330 2637
rect 1367 2633 1371 2634
rect 1551 2638 1555 2639
rect 1551 2633 1555 2634
rect 1607 2638 1611 2639
rect 1607 2633 1611 2634
rect 1663 2638 1667 2639
rect 1663 2633 1667 2634
rect 1719 2638 1723 2639
rect 1719 2633 1723 2634
rect 1775 2638 1779 2639
rect 1775 2633 1779 2634
rect 1831 2638 1835 2639
rect 1831 2633 1835 2634
rect 1887 2638 1891 2639
rect 1887 2633 1891 2634
rect 1943 2638 1947 2639
rect 1943 2633 1947 2634
rect 1999 2638 2003 2639
rect 1999 2633 2003 2634
rect 2055 2638 2059 2639
rect 2055 2633 2059 2634
rect 2111 2638 2115 2639
rect 2111 2633 2115 2634
rect 2167 2638 2171 2639
rect 2167 2633 2171 2634
rect 2583 2638 2587 2639
rect 2583 2633 2587 2634
rect 110 2621 116 2622
rect 110 2617 111 2621
rect 115 2617 116 2621
rect 110 2616 116 2617
rect 1326 2621 1332 2622
rect 1326 2617 1327 2621
rect 1331 2617 1332 2621
rect 1368 2618 1370 2633
rect 1552 2627 1554 2633
rect 1608 2627 1610 2633
rect 1664 2627 1666 2633
rect 1720 2627 1722 2633
rect 1776 2627 1778 2633
rect 1832 2627 1834 2633
rect 1888 2627 1890 2633
rect 1944 2627 1946 2633
rect 2000 2627 2002 2633
rect 2056 2627 2058 2633
rect 2112 2627 2114 2633
rect 2168 2627 2170 2633
rect 1550 2626 1556 2627
rect 1550 2622 1551 2626
rect 1555 2622 1556 2626
rect 1550 2621 1556 2622
rect 1606 2626 1612 2627
rect 1606 2622 1607 2626
rect 1611 2622 1612 2626
rect 1606 2621 1612 2622
rect 1662 2626 1668 2627
rect 1662 2622 1663 2626
rect 1667 2622 1668 2626
rect 1662 2621 1668 2622
rect 1718 2626 1724 2627
rect 1718 2622 1719 2626
rect 1723 2622 1724 2626
rect 1718 2621 1724 2622
rect 1774 2626 1780 2627
rect 1774 2622 1775 2626
rect 1779 2622 1780 2626
rect 1774 2621 1780 2622
rect 1830 2626 1836 2627
rect 1830 2622 1831 2626
rect 1835 2622 1836 2626
rect 1830 2621 1836 2622
rect 1886 2626 1892 2627
rect 1886 2622 1887 2626
rect 1891 2622 1892 2626
rect 1886 2621 1892 2622
rect 1942 2626 1948 2627
rect 1942 2622 1943 2626
rect 1947 2622 1948 2626
rect 1942 2621 1948 2622
rect 1998 2626 2004 2627
rect 1998 2622 1999 2626
rect 2003 2622 2004 2626
rect 1998 2621 2004 2622
rect 2054 2626 2060 2627
rect 2054 2622 2055 2626
rect 2059 2622 2060 2626
rect 2054 2621 2060 2622
rect 2110 2626 2116 2627
rect 2110 2622 2111 2626
rect 2115 2622 2116 2626
rect 2110 2621 2116 2622
rect 2166 2626 2172 2627
rect 2166 2622 2167 2626
rect 2171 2622 2172 2626
rect 2166 2621 2172 2622
rect 2584 2618 2586 2633
rect 1326 2616 1332 2617
rect 1366 2617 1372 2618
rect 1366 2613 1367 2617
rect 1371 2613 1372 2617
rect 1366 2612 1372 2613
rect 2582 2617 2588 2618
rect 2582 2613 2583 2617
rect 2587 2613 2588 2617
rect 2582 2612 2588 2613
rect 110 2604 116 2605
rect 1326 2604 1332 2605
rect 110 2600 111 2604
rect 115 2600 116 2604
rect 110 2599 116 2600
rect 534 2603 540 2604
rect 534 2599 535 2603
rect 539 2599 540 2603
rect 112 2587 114 2599
rect 534 2598 540 2599
rect 590 2603 596 2604
rect 590 2599 591 2603
rect 595 2599 596 2603
rect 590 2598 596 2599
rect 646 2603 652 2604
rect 646 2599 647 2603
rect 651 2599 652 2603
rect 646 2598 652 2599
rect 702 2603 708 2604
rect 702 2599 703 2603
rect 707 2599 708 2603
rect 702 2598 708 2599
rect 758 2603 764 2604
rect 758 2599 759 2603
rect 763 2599 764 2603
rect 1326 2600 1327 2604
rect 1331 2600 1332 2604
rect 1326 2599 1332 2600
rect 1366 2600 1372 2601
rect 2582 2600 2588 2601
rect 758 2598 764 2599
rect 536 2587 538 2598
rect 592 2587 594 2598
rect 648 2587 650 2598
rect 704 2587 706 2598
rect 760 2587 762 2598
rect 1328 2587 1330 2599
rect 1366 2596 1367 2600
rect 1371 2596 1372 2600
rect 1366 2595 1372 2596
rect 1534 2599 1540 2600
rect 1534 2595 1535 2599
rect 1539 2595 1540 2599
rect 111 2586 115 2587
rect 111 2581 115 2582
rect 215 2586 219 2587
rect 215 2581 219 2582
rect 271 2586 275 2587
rect 271 2581 275 2582
rect 327 2586 331 2587
rect 327 2581 331 2582
rect 383 2586 387 2587
rect 383 2581 387 2582
rect 439 2586 443 2587
rect 439 2581 443 2582
rect 495 2586 499 2587
rect 495 2581 499 2582
rect 535 2586 539 2587
rect 535 2581 539 2582
rect 551 2586 555 2587
rect 551 2581 555 2582
rect 591 2586 595 2587
rect 591 2581 595 2582
rect 607 2586 611 2587
rect 607 2581 611 2582
rect 647 2586 651 2587
rect 647 2581 651 2582
rect 663 2586 667 2587
rect 663 2581 667 2582
rect 703 2586 707 2587
rect 703 2581 707 2582
rect 719 2586 723 2587
rect 719 2581 723 2582
rect 759 2586 763 2587
rect 759 2581 763 2582
rect 775 2586 779 2587
rect 775 2581 779 2582
rect 831 2586 835 2587
rect 831 2581 835 2582
rect 887 2586 891 2587
rect 887 2581 891 2582
rect 943 2586 947 2587
rect 943 2581 947 2582
rect 999 2586 1003 2587
rect 999 2581 1003 2582
rect 1055 2586 1059 2587
rect 1055 2581 1059 2582
rect 1111 2586 1115 2587
rect 1111 2581 1115 2582
rect 1327 2586 1331 2587
rect 1368 2583 1370 2595
rect 1534 2594 1540 2595
rect 1590 2599 1596 2600
rect 1590 2595 1591 2599
rect 1595 2595 1596 2599
rect 1590 2594 1596 2595
rect 1646 2599 1652 2600
rect 1646 2595 1647 2599
rect 1651 2595 1652 2599
rect 1646 2594 1652 2595
rect 1702 2599 1708 2600
rect 1702 2595 1703 2599
rect 1707 2595 1708 2599
rect 1702 2594 1708 2595
rect 1758 2599 1764 2600
rect 1758 2595 1759 2599
rect 1763 2595 1764 2599
rect 1758 2594 1764 2595
rect 1814 2599 1820 2600
rect 1814 2595 1815 2599
rect 1819 2595 1820 2599
rect 1814 2594 1820 2595
rect 1870 2599 1876 2600
rect 1870 2595 1871 2599
rect 1875 2595 1876 2599
rect 1870 2594 1876 2595
rect 1926 2599 1932 2600
rect 1926 2595 1927 2599
rect 1931 2595 1932 2599
rect 1926 2594 1932 2595
rect 1982 2599 1988 2600
rect 1982 2595 1983 2599
rect 1987 2595 1988 2599
rect 1982 2594 1988 2595
rect 2038 2599 2044 2600
rect 2038 2595 2039 2599
rect 2043 2595 2044 2599
rect 2038 2594 2044 2595
rect 2094 2599 2100 2600
rect 2094 2595 2095 2599
rect 2099 2595 2100 2599
rect 2094 2594 2100 2595
rect 2150 2599 2156 2600
rect 2150 2595 2151 2599
rect 2155 2595 2156 2599
rect 2582 2596 2583 2600
rect 2587 2596 2588 2600
rect 2582 2595 2588 2596
rect 2150 2594 2156 2595
rect 1536 2583 1538 2594
rect 1592 2583 1594 2594
rect 1648 2583 1650 2594
rect 1704 2583 1706 2594
rect 1760 2583 1762 2594
rect 1816 2583 1818 2594
rect 1872 2583 1874 2594
rect 1928 2583 1930 2594
rect 1984 2583 1986 2594
rect 2040 2583 2042 2594
rect 2096 2583 2098 2594
rect 2152 2583 2154 2594
rect 2584 2583 2586 2595
rect 1327 2581 1331 2582
rect 1367 2582 1371 2583
rect 112 2569 114 2581
rect 216 2570 218 2581
rect 272 2570 274 2581
rect 328 2570 330 2581
rect 384 2570 386 2581
rect 440 2570 442 2581
rect 496 2570 498 2581
rect 552 2570 554 2581
rect 608 2570 610 2581
rect 664 2570 666 2581
rect 720 2570 722 2581
rect 776 2570 778 2581
rect 832 2570 834 2581
rect 888 2570 890 2581
rect 944 2570 946 2581
rect 1000 2570 1002 2581
rect 1056 2570 1058 2581
rect 1112 2570 1114 2581
rect 214 2569 220 2570
rect 110 2568 116 2569
rect 110 2564 111 2568
rect 115 2564 116 2568
rect 214 2565 215 2569
rect 219 2565 220 2569
rect 214 2564 220 2565
rect 270 2569 276 2570
rect 270 2565 271 2569
rect 275 2565 276 2569
rect 270 2564 276 2565
rect 326 2569 332 2570
rect 326 2565 327 2569
rect 331 2565 332 2569
rect 326 2564 332 2565
rect 382 2569 388 2570
rect 382 2565 383 2569
rect 387 2565 388 2569
rect 382 2564 388 2565
rect 438 2569 444 2570
rect 438 2565 439 2569
rect 443 2565 444 2569
rect 438 2564 444 2565
rect 494 2569 500 2570
rect 494 2565 495 2569
rect 499 2565 500 2569
rect 494 2564 500 2565
rect 550 2569 556 2570
rect 550 2565 551 2569
rect 555 2565 556 2569
rect 550 2564 556 2565
rect 606 2569 612 2570
rect 606 2565 607 2569
rect 611 2565 612 2569
rect 606 2564 612 2565
rect 662 2569 668 2570
rect 662 2565 663 2569
rect 667 2565 668 2569
rect 662 2564 668 2565
rect 718 2569 724 2570
rect 718 2565 719 2569
rect 723 2565 724 2569
rect 718 2564 724 2565
rect 774 2569 780 2570
rect 774 2565 775 2569
rect 779 2565 780 2569
rect 774 2564 780 2565
rect 830 2569 836 2570
rect 830 2565 831 2569
rect 835 2565 836 2569
rect 830 2564 836 2565
rect 886 2569 892 2570
rect 886 2565 887 2569
rect 891 2565 892 2569
rect 886 2564 892 2565
rect 942 2569 948 2570
rect 942 2565 943 2569
rect 947 2565 948 2569
rect 942 2564 948 2565
rect 998 2569 1004 2570
rect 998 2565 999 2569
rect 1003 2565 1004 2569
rect 998 2564 1004 2565
rect 1054 2569 1060 2570
rect 1054 2565 1055 2569
rect 1059 2565 1060 2569
rect 1054 2564 1060 2565
rect 1110 2569 1116 2570
rect 1328 2569 1330 2581
rect 1367 2577 1371 2578
rect 1439 2582 1443 2583
rect 1439 2577 1443 2578
rect 1535 2582 1539 2583
rect 1535 2577 1539 2578
rect 1543 2582 1547 2583
rect 1543 2577 1547 2578
rect 1591 2582 1595 2583
rect 1591 2577 1595 2578
rect 1647 2582 1651 2583
rect 1647 2577 1651 2578
rect 1655 2582 1659 2583
rect 1655 2577 1659 2578
rect 1703 2582 1707 2583
rect 1703 2577 1707 2578
rect 1759 2582 1763 2583
rect 1759 2577 1763 2578
rect 1767 2582 1771 2583
rect 1767 2577 1771 2578
rect 1815 2582 1819 2583
rect 1815 2577 1819 2578
rect 1871 2582 1875 2583
rect 1871 2577 1875 2578
rect 1879 2582 1883 2583
rect 1879 2577 1883 2578
rect 1927 2582 1931 2583
rect 1927 2577 1931 2578
rect 1983 2582 1987 2583
rect 1983 2577 1987 2578
rect 1991 2582 1995 2583
rect 1991 2577 1995 2578
rect 2039 2582 2043 2583
rect 2039 2577 2043 2578
rect 2095 2582 2099 2583
rect 2095 2577 2099 2578
rect 2111 2582 2115 2583
rect 2111 2577 2115 2578
rect 2151 2582 2155 2583
rect 2151 2577 2155 2578
rect 2231 2582 2235 2583
rect 2231 2577 2235 2578
rect 2351 2582 2355 2583
rect 2351 2577 2355 2578
rect 2583 2582 2587 2583
rect 2583 2577 2587 2578
rect 1110 2565 1111 2569
rect 1115 2565 1116 2569
rect 1110 2564 1116 2565
rect 1326 2568 1332 2569
rect 1326 2564 1327 2568
rect 1331 2564 1332 2568
rect 1368 2565 1370 2577
rect 1440 2566 1442 2577
rect 1544 2566 1546 2577
rect 1656 2566 1658 2577
rect 1768 2566 1770 2577
rect 1880 2566 1882 2577
rect 1992 2566 1994 2577
rect 2112 2566 2114 2577
rect 2232 2566 2234 2577
rect 2352 2566 2354 2577
rect 1438 2565 1444 2566
rect 110 2563 116 2564
rect 1326 2563 1332 2564
rect 1366 2564 1372 2565
rect 1366 2560 1367 2564
rect 1371 2560 1372 2564
rect 1438 2561 1439 2565
rect 1443 2561 1444 2565
rect 1438 2560 1444 2561
rect 1542 2565 1548 2566
rect 1542 2561 1543 2565
rect 1547 2561 1548 2565
rect 1542 2560 1548 2561
rect 1654 2565 1660 2566
rect 1654 2561 1655 2565
rect 1659 2561 1660 2565
rect 1654 2560 1660 2561
rect 1766 2565 1772 2566
rect 1766 2561 1767 2565
rect 1771 2561 1772 2565
rect 1766 2560 1772 2561
rect 1878 2565 1884 2566
rect 1878 2561 1879 2565
rect 1883 2561 1884 2565
rect 1878 2560 1884 2561
rect 1990 2565 1996 2566
rect 1990 2561 1991 2565
rect 1995 2561 1996 2565
rect 1990 2560 1996 2561
rect 2110 2565 2116 2566
rect 2110 2561 2111 2565
rect 2115 2561 2116 2565
rect 2110 2560 2116 2561
rect 2230 2565 2236 2566
rect 2230 2561 2231 2565
rect 2235 2561 2236 2565
rect 2230 2560 2236 2561
rect 2350 2565 2356 2566
rect 2584 2565 2586 2577
rect 2350 2561 2351 2565
rect 2355 2561 2356 2565
rect 2350 2560 2356 2561
rect 2582 2564 2588 2565
rect 2582 2560 2583 2564
rect 2587 2560 2588 2564
rect 1366 2559 1372 2560
rect 2582 2559 2588 2560
rect 110 2551 116 2552
rect 110 2547 111 2551
rect 115 2547 116 2551
rect 110 2546 116 2547
rect 1326 2551 1332 2552
rect 1326 2547 1327 2551
rect 1331 2547 1332 2551
rect 1326 2546 1332 2547
rect 1366 2547 1372 2548
rect 112 2527 114 2546
rect 230 2542 236 2543
rect 230 2538 231 2542
rect 235 2538 236 2542
rect 230 2537 236 2538
rect 286 2542 292 2543
rect 286 2538 287 2542
rect 291 2538 292 2542
rect 286 2537 292 2538
rect 342 2542 348 2543
rect 342 2538 343 2542
rect 347 2538 348 2542
rect 342 2537 348 2538
rect 398 2542 404 2543
rect 398 2538 399 2542
rect 403 2538 404 2542
rect 398 2537 404 2538
rect 454 2542 460 2543
rect 454 2538 455 2542
rect 459 2538 460 2542
rect 454 2537 460 2538
rect 510 2542 516 2543
rect 510 2538 511 2542
rect 515 2538 516 2542
rect 510 2537 516 2538
rect 566 2542 572 2543
rect 566 2538 567 2542
rect 571 2538 572 2542
rect 566 2537 572 2538
rect 622 2542 628 2543
rect 622 2538 623 2542
rect 627 2538 628 2542
rect 622 2537 628 2538
rect 678 2542 684 2543
rect 678 2538 679 2542
rect 683 2538 684 2542
rect 678 2537 684 2538
rect 734 2542 740 2543
rect 734 2538 735 2542
rect 739 2538 740 2542
rect 734 2537 740 2538
rect 790 2542 796 2543
rect 790 2538 791 2542
rect 795 2538 796 2542
rect 790 2537 796 2538
rect 846 2542 852 2543
rect 846 2538 847 2542
rect 851 2538 852 2542
rect 846 2537 852 2538
rect 902 2542 908 2543
rect 902 2538 903 2542
rect 907 2538 908 2542
rect 902 2537 908 2538
rect 958 2542 964 2543
rect 958 2538 959 2542
rect 963 2538 964 2542
rect 958 2537 964 2538
rect 1014 2542 1020 2543
rect 1014 2538 1015 2542
rect 1019 2538 1020 2542
rect 1014 2537 1020 2538
rect 1070 2542 1076 2543
rect 1070 2538 1071 2542
rect 1075 2538 1076 2542
rect 1070 2537 1076 2538
rect 1126 2542 1132 2543
rect 1126 2538 1127 2542
rect 1131 2538 1132 2542
rect 1126 2537 1132 2538
rect 232 2527 234 2537
rect 288 2527 290 2537
rect 344 2527 346 2537
rect 400 2527 402 2537
rect 456 2527 458 2537
rect 512 2527 514 2537
rect 568 2527 570 2537
rect 624 2527 626 2537
rect 680 2527 682 2537
rect 736 2527 738 2537
rect 792 2527 794 2537
rect 848 2527 850 2537
rect 904 2527 906 2537
rect 960 2527 962 2537
rect 1016 2527 1018 2537
rect 1072 2527 1074 2537
rect 1128 2527 1130 2537
rect 1328 2527 1330 2546
rect 1366 2543 1367 2547
rect 1371 2543 1372 2547
rect 1366 2542 1372 2543
rect 2582 2547 2588 2548
rect 2582 2543 2583 2547
rect 2587 2543 2588 2547
rect 2582 2542 2588 2543
rect 111 2526 115 2527
rect 111 2521 115 2522
rect 231 2526 235 2527
rect 231 2521 235 2522
rect 287 2526 291 2527
rect 287 2521 291 2522
rect 343 2526 347 2527
rect 343 2521 347 2522
rect 367 2526 371 2527
rect 367 2521 371 2522
rect 399 2526 403 2527
rect 399 2521 403 2522
rect 423 2526 427 2527
rect 423 2521 427 2522
rect 455 2526 459 2527
rect 455 2521 459 2522
rect 487 2526 491 2527
rect 487 2521 491 2522
rect 511 2526 515 2527
rect 511 2521 515 2522
rect 551 2526 555 2527
rect 551 2521 555 2522
rect 567 2526 571 2527
rect 567 2521 571 2522
rect 615 2526 619 2527
rect 615 2521 619 2522
rect 623 2526 627 2527
rect 623 2521 627 2522
rect 679 2526 683 2527
rect 679 2521 683 2522
rect 735 2526 739 2527
rect 735 2521 739 2522
rect 743 2526 747 2527
rect 743 2521 747 2522
rect 791 2526 795 2527
rect 791 2521 795 2522
rect 807 2526 811 2527
rect 807 2521 811 2522
rect 847 2526 851 2527
rect 847 2521 851 2522
rect 871 2526 875 2527
rect 871 2521 875 2522
rect 903 2526 907 2527
rect 903 2521 907 2522
rect 943 2526 947 2527
rect 943 2521 947 2522
rect 959 2526 963 2527
rect 959 2521 963 2522
rect 1015 2526 1019 2527
rect 1015 2521 1019 2522
rect 1071 2526 1075 2527
rect 1071 2521 1075 2522
rect 1127 2526 1131 2527
rect 1127 2521 1131 2522
rect 1327 2526 1331 2527
rect 1327 2521 1331 2522
rect 112 2506 114 2521
rect 368 2515 370 2521
rect 424 2515 426 2521
rect 488 2515 490 2521
rect 552 2515 554 2521
rect 616 2515 618 2521
rect 680 2515 682 2521
rect 744 2515 746 2521
rect 808 2515 810 2521
rect 872 2515 874 2521
rect 944 2515 946 2521
rect 1016 2515 1018 2521
rect 366 2514 372 2515
rect 366 2510 367 2514
rect 371 2510 372 2514
rect 366 2509 372 2510
rect 422 2514 428 2515
rect 422 2510 423 2514
rect 427 2510 428 2514
rect 422 2509 428 2510
rect 486 2514 492 2515
rect 486 2510 487 2514
rect 491 2510 492 2514
rect 486 2509 492 2510
rect 550 2514 556 2515
rect 550 2510 551 2514
rect 555 2510 556 2514
rect 550 2509 556 2510
rect 614 2514 620 2515
rect 614 2510 615 2514
rect 619 2510 620 2514
rect 614 2509 620 2510
rect 678 2514 684 2515
rect 678 2510 679 2514
rect 683 2510 684 2514
rect 678 2509 684 2510
rect 742 2514 748 2515
rect 742 2510 743 2514
rect 747 2510 748 2514
rect 742 2509 748 2510
rect 806 2514 812 2515
rect 806 2510 807 2514
rect 811 2510 812 2514
rect 806 2509 812 2510
rect 870 2514 876 2515
rect 870 2510 871 2514
rect 875 2510 876 2514
rect 870 2509 876 2510
rect 942 2514 948 2515
rect 942 2510 943 2514
rect 947 2510 948 2514
rect 942 2509 948 2510
rect 1014 2514 1020 2515
rect 1014 2510 1015 2514
rect 1019 2510 1020 2514
rect 1014 2509 1020 2510
rect 1328 2506 1330 2521
rect 1368 2519 1370 2542
rect 1454 2538 1460 2539
rect 1454 2534 1455 2538
rect 1459 2534 1460 2538
rect 1454 2533 1460 2534
rect 1558 2538 1564 2539
rect 1558 2534 1559 2538
rect 1563 2534 1564 2538
rect 1558 2533 1564 2534
rect 1670 2538 1676 2539
rect 1670 2534 1671 2538
rect 1675 2534 1676 2538
rect 1670 2533 1676 2534
rect 1782 2538 1788 2539
rect 1782 2534 1783 2538
rect 1787 2534 1788 2538
rect 1782 2533 1788 2534
rect 1894 2538 1900 2539
rect 1894 2534 1895 2538
rect 1899 2534 1900 2538
rect 1894 2533 1900 2534
rect 2006 2538 2012 2539
rect 2006 2534 2007 2538
rect 2011 2534 2012 2538
rect 2006 2533 2012 2534
rect 2126 2538 2132 2539
rect 2126 2534 2127 2538
rect 2131 2534 2132 2538
rect 2126 2533 2132 2534
rect 2246 2538 2252 2539
rect 2246 2534 2247 2538
rect 2251 2534 2252 2538
rect 2246 2533 2252 2534
rect 2366 2538 2372 2539
rect 2366 2534 2367 2538
rect 2371 2534 2372 2538
rect 2366 2533 2372 2534
rect 1456 2519 1458 2533
rect 1560 2519 1562 2533
rect 1672 2519 1674 2533
rect 1784 2519 1786 2533
rect 1896 2519 1898 2533
rect 2008 2519 2010 2533
rect 2128 2519 2130 2533
rect 2248 2519 2250 2533
rect 2368 2519 2370 2533
rect 2584 2519 2586 2542
rect 1367 2518 1371 2519
rect 1367 2513 1371 2514
rect 1455 2518 1459 2519
rect 1455 2513 1459 2514
rect 1551 2518 1555 2519
rect 1551 2513 1555 2514
rect 1559 2518 1563 2519
rect 1559 2513 1563 2514
rect 1631 2518 1635 2519
rect 1631 2513 1635 2514
rect 1671 2518 1675 2519
rect 1671 2513 1675 2514
rect 1719 2518 1723 2519
rect 1719 2513 1723 2514
rect 1783 2518 1787 2519
rect 1783 2513 1787 2514
rect 1807 2518 1811 2519
rect 1807 2513 1811 2514
rect 1895 2518 1899 2519
rect 1895 2513 1899 2514
rect 1903 2518 1907 2519
rect 1903 2513 1907 2514
rect 1999 2518 2003 2519
rect 1999 2513 2003 2514
rect 2007 2518 2011 2519
rect 2007 2513 2011 2514
rect 2095 2518 2099 2519
rect 2095 2513 2099 2514
rect 2127 2518 2131 2519
rect 2127 2513 2131 2514
rect 2191 2518 2195 2519
rect 2191 2513 2195 2514
rect 2247 2518 2251 2519
rect 2247 2513 2251 2514
rect 2295 2518 2299 2519
rect 2295 2513 2299 2514
rect 2367 2518 2371 2519
rect 2367 2513 2371 2514
rect 2399 2518 2403 2519
rect 2399 2513 2403 2514
rect 2583 2518 2587 2519
rect 2583 2513 2587 2514
rect 110 2505 116 2506
rect 110 2501 111 2505
rect 115 2501 116 2505
rect 110 2500 116 2501
rect 1326 2505 1332 2506
rect 1326 2501 1327 2505
rect 1331 2501 1332 2505
rect 1326 2500 1332 2501
rect 1368 2498 1370 2513
rect 1552 2507 1554 2513
rect 1632 2507 1634 2513
rect 1720 2507 1722 2513
rect 1808 2507 1810 2513
rect 1904 2507 1906 2513
rect 2000 2507 2002 2513
rect 2096 2507 2098 2513
rect 2192 2507 2194 2513
rect 2296 2507 2298 2513
rect 2400 2507 2402 2513
rect 1550 2506 1556 2507
rect 1550 2502 1551 2506
rect 1555 2502 1556 2506
rect 1550 2501 1556 2502
rect 1630 2506 1636 2507
rect 1630 2502 1631 2506
rect 1635 2502 1636 2506
rect 1630 2501 1636 2502
rect 1718 2506 1724 2507
rect 1718 2502 1719 2506
rect 1723 2502 1724 2506
rect 1718 2501 1724 2502
rect 1806 2506 1812 2507
rect 1806 2502 1807 2506
rect 1811 2502 1812 2506
rect 1806 2501 1812 2502
rect 1902 2506 1908 2507
rect 1902 2502 1903 2506
rect 1907 2502 1908 2506
rect 1902 2501 1908 2502
rect 1998 2506 2004 2507
rect 1998 2502 1999 2506
rect 2003 2502 2004 2506
rect 1998 2501 2004 2502
rect 2094 2506 2100 2507
rect 2094 2502 2095 2506
rect 2099 2502 2100 2506
rect 2094 2501 2100 2502
rect 2190 2506 2196 2507
rect 2190 2502 2191 2506
rect 2195 2502 2196 2506
rect 2190 2501 2196 2502
rect 2294 2506 2300 2507
rect 2294 2502 2295 2506
rect 2299 2502 2300 2506
rect 2294 2501 2300 2502
rect 2398 2506 2404 2507
rect 2398 2502 2399 2506
rect 2403 2502 2404 2506
rect 2398 2501 2404 2502
rect 2584 2498 2586 2513
rect 1366 2497 1372 2498
rect 1366 2493 1367 2497
rect 1371 2493 1372 2497
rect 1366 2492 1372 2493
rect 2582 2497 2588 2498
rect 2582 2493 2583 2497
rect 2587 2493 2588 2497
rect 2582 2492 2588 2493
rect 110 2488 116 2489
rect 1326 2488 1332 2489
rect 110 2484 111 2488
rect 115 2484 116 2488
rect 110 2483 116 2484
rect 350 2487 356 2488
rect 350 2483 351 2487
rect 355 2483 356 2487
rect 112 2467 114 2483
rect 350 2482 356 2483
rect 406 2487 412 2488
rect 406 2483 407 2487
rect 411 2483 412 2487
rect 406 2482 412 2483
rect 470 2487 476 2488
rect 470 2483 471 2487
rect 475 2483 476 2487
rect 470 2482 476 2483
rect 534 2487 540 2488
rect 534 2483 535 2487
rect 539 2483 540 2487
rect 534 2482 540 2483
rect 598 2487 604 2488
rect 598 2483 599 2487
rect 603 2483 604 2487
rect 598 2482 604 2483
rect 662 2487 668 2488
rect 662 2483 663 2487
rect 667 2483 668 2487
rect 662 2482 668 2483
rect 726 2487 732 2488
rect 726 2483 727 2487
rect 731 2483 732 2487
rect 726 2482 732 2483
rect 790 2487 796 2488
rect 790 2483 791 2487
rect 795 2483 796 2487
rect 790 2482 796 2483
rect 854 2487 860 2488
rect 854 2483 855 2487
rect 859 2483 860 2487
rect 854 2482 860 2483
rect 926 2487 932 2488
rect 926 2483 927 2487
rect 931 2483 932 2487
rect 926 2482 932 2483
rect 998 2487 1004 2488
rect 998 2483 999 2487
rect 1003 2483 1004 2487
rect 1326 2484 1327 2488
rect 1331 2484 1332 2488
rect 1326 2483 1332 2484
rect 998 2482 1004 2483
rect 352 2467 354 2482
rect 408 2467 410 2482
rect 472 2467 474 2482
rect 536 2467 538 2482
rect 600 2467 602 2482
rect 664 2467 666 2482
rect 728 2467 730 2482
rect 792 2467 794 2482
rect 856 2467 858 2482
rect 928 2467 930 2482
rect 1000 2467 1002 2482
rect 1328 2467 1330 2483
rect 1366 2480 1372 2481
rect 2582 2480 2588 2481
rect 1366 2476 1367 2480
rect 1371 2476 1372 2480
rect 1366 2475 1372 2476
rect 1534 2479 1540 2480
rect 1534 2475 1535 2479
rect 1539 2475 1540 2479
rect 111 2466 115 2467
rect 111 2461 115 2462
rect 271 2466 275 2467
rect 271 2461 275 2462
rect 335 2466 339 2467
rect 335 2461 339 2462
rect 351 2466 355 2467
rect 351 2461 355 2462
rect 399 2466 403 2467
rect 399 2461 403 2462
rect 407 2466 411 2467
rect 407 2461 411 2462
rect 471 2466 475 2467
rect 471 2461 475 2462
rect 535 2466 539 2467
rect 535 2461 539 2462
rect 551 2466 555 2467
rect 551 2461 555 2462
rect 599 2466 603 2467
rect 599 2461 603 2462
rect 631 2466 635 2467
rect 631 2461 635 2462
rect 663 2466 667 2467
rect 663 2461 667 2462
rect 711 2466 715 2467
rect 711 2461 715 2462
rect 727 2466 731 2467
rect 727 2461 731 2462
rect 783 2466 787 2467
rect 783 2461 787 2462
rect 791 2466 795 2467
rect 791 2461 795 2462
rect 855 2466 859 2467
rect 855 2461 859 2462
rect 863 2466 867 2467
rect 863 2461 867 2462
rect 927 2466 931 2467
rect 927 2461 931 2462
rect 943 2466 947 2467
rect 943 2461 947 2462
rect 999 2466 1003 2467
rect 999 2461 1003 2462
rect 1023 2466 1027 2467
rect 1023 2461 1027 2462
rect 1327 2466 1331 2467
rect 1368 2463 1370 2475
rect 1534 2474 1540 2475
rect 1614 2479 1620 2480
rect 1614 2475 1615 2479
rect 1619 2475 1620 2479
rect 1614 2474 1620 2475
rect 1702 2479 1708 2480
rect 1702 2475 1703 2479
rect 1707 2475 1708 2479
rect 1702 2474 1708 2475
rect 1790 2479 1796 2480
rect 1790 2475 1791 2479
rect 1795 2475 1796 2479
rect 1790 2474 1796 2475
rect 1886 2479 1892 2480
rect 1886 2475 1887 2479
rect 1891 2475 1892 2479
rect 1886 2474 1892 2475
rect 1982 2479 1988 2480
rect 1982 2475 1983 2479
rect 1987 2475 1988 2479
rect 1982 2474 1988 2475
rect 2078 2479 2084 2480
rect 2078 2475 2079 2479
rect 2083 2475 2084 2479
rect 2078 2474 2084 2475
rect 2174 2479 2180 2480
rect 2174 2475 2175 2479
rect 2179 2475 2180 2479
rect 2174 2474 2180 2475
rect 2278 2479 2284 2480
rect 2278 2475 2279 2479
rect 2283 2475 2284 2479
rect 2278 2474 2284 2475
rect 2382 2479 2388 2480
rect 2382 2475 2383 2479
rect 2387 2475 2388 2479
rect 2582 2476 2583 2480
rect 2587 2476 2588 2480
rect 2582 2475 2588 2476
rect 2382 2474 2388 2475
rect 1536 2463 1538 2474
rect 1616 2463 1618 2474
rect 1704 2463 1706 2474
rect 1792 2463 1794 2474
rect 1888 2463 1890 2474
rect 1984 2463 1986 2474
rect 2080 2463 2082 2474
rect 2176 2463 2178 2474
rect 2280 2463 2282 2474
rect 2384 2463 2386 2474
rect 2584 2463 2586 2475
rect 1327 2461 1331 2462
rect 1367 2462 1371 2463
rect 112 2449 114 2461
rect 272 2450 274 2461
rect 336 2450 338 2461
rect 400 2450 402 2461
rect 472 2450 474 2461
rect 552 2450 554 2461
rect 632 2450 634 2461
rect 712 2450 714 2461
rect 784 2450 786 2461
rect 864 2450 866 2461
rect 944 2450 946 2461
rect 1024 2450 1026 2461
rect 270 2449 276 2450
rect 110 2448 116 2449
rect 110 2444 111 2448
rect 115 2444 116 2448
rect 270 2445 271 2449
rect 275 2445 276 2449
rect 270 2444 276 2445
rect 334 2449 340 2450
rect 334 2445 335 2449
rect 339 2445 340 2449
rect 334 2444 340 2445
rect 398 2449 404 2450
rect 398 2445 399 2449
rect 403 2445 404 2449
rect 398 2444 404 2445
rect 470 2449 476 2450
rect 470 2445 471 2449
rect 475 2445 476 2449
rect 470 2444 476 2445
rect 550 2449 556 2450
rect 550 2445 551 2449
rect 555 2445 556 2449
rect 550 2444 556 2445
rect 630 2449 636 2450
rect 630 2445 631 2449
rect 635 2445 636 2449
rect 630 2444 636 2445
rect 710 2449 716 2450
rect 710 2445 711 2449
rect 715 2445 716 2449
rect 710 2444 716 2445
rect 782 2449 788 2450
rect 782 2445 783 2449
rect 787 2445 788 2449
rect 782 2444 788 2445
rect 862 2449 868 2450
rect 862 2445 863 2449
rect 867 2445 868 2449
rect 862 2444 868 2445
rect 942 2449 948 2450
rect 942 2445 943 2449
rect 947 2445 948 2449
rect 942 2444 948 2445
rect 1022 2449 1028 2450
rect 1328 2449 1330 2461
rect 1367 2457 1371 2458
rect 1535 2462 1539 2463
rect 1535 2457 1539 2458
rect 1615 2462 1619 2463
rect 1615 2457 1619 2458
rect 1647 2462 1651 2463
rect 1647 2457 1651 2458
rect 1703 2462 1707 2463
rect 1703 2457 1707 2458
rect 1767 2462 1771 2463
rect 1767 2457 1771 2458
rect 1791 2462 1795 2463
rect 1791 2457 1795 2458
rect 1839 2462 1843 2463
rect 1839 2457 1843 2458
rect 1887 2462 1891 2463
rect 1887 2457 1891 2458
rect 1911 2462 1915 2463
rect 1911 2457 1915 2458
rect 1983 2462 1987 2463
rect 1983 2457 1987 2458
rect 1991 2462 1995 2463
rect 1991 2457 1995 2458
rect 2079 2462 2083 2463
rect 2079 2457 2083 2458
rect 2167 2462 2171 2463
rect 2167 2457 2171 2458
rect 2175 2462 2179 2463
rect 2175 2457 2179 2458
rect 2263 2462 2267 2463
rect 2263 2457 2267 2458
rect 2279 2462 2283 2463
rect 2279 2457 2283 2458
rect 2359 2462 2363 2463
rect 2359 2457 2363 2458
rect 2383 2462 2387 2463
rect 2383 2457 2387 2458
rect 2455 2462 2459 2463
rect 2455 2457 2459 2458
rect 2527 2462 2531 2463
rect 2527 2457 2531 2458
rect 2583 2462 2587 2463
rect 2583 2457 2587 2458
rect 1022 2445 1023 2449
rect 1027 2445 1028 2449
rect 1022 2444 1028 2445
rect 1326 2448 1332 2449
rect 1326 2444 1327 2448
rect 1331 2444 1332 2448
rect 1368 2445 1370 2457
rect 1648 2446 1650 2457
rect 1704 2446 1706 2457
rect 1768 2446 1770 2457
rect 1840 2446 1842 2457
rect 1912 2446 1914 2457
rect 1992 2446 1994 2457
rect 2080 2446 2082 2457
rect 2168 2446 2170 2457
rect 2264 2446 2266 2457
rect 2360 2446 2362 2457
rect 2456 2446 2458 2457
rect 2528 2446 2530 2457
rect 1646 2445 1652 2446
rect 110 2443 116 2444
rect 1326 2443 1332 2444
rect 1366 2444 1372 2445
rect 1366 2440 1367 2444
rect 1371 2440 1372 2444
rect 1646 2441 1647 2445
rect 1651 2441 1652 2445
rect 1646 2440 1652 2441
rect 1702 2445 1708 2446
rect 1702 2441 1703 2445
rect 1707 2441 1708 2445
rect 1702 2440 1708 2441
rect 1766 2445 1772 2446
rect 1766 2441 1767 2445
rect 1771 2441 1772 2445
rect 1766 2440 1772 2441
rect 1838 2445 1844 2446
rect 1838 2441 1839 2445
rect 1843 2441 1844 2445
rect 1838 2440 1844 2441
rect 1910 2445 1916 2446
rect 1910 2441 1911 2445
rect 1915 2441 1916 2445
rect 1910 2440 1916 2441
rect 1990 2445 1996 2446
rect 1990 2441 1991 2445
rect 1995 2441 1996 2445
rect 1990 2440 1996 2441
rect 2078 2445 2084 2446
rect 2078 2441 2079 2445
rect 2083 2441 2084 2445
rect 2078 2440 2084 2441
rect 2166 2445 2172 2446
rect 2166 2441 2167 2445
rect 2171 2441 2172 2445
rect 2166 2440 2172 2441
rect 2262 2445 2268 2446
rect 2262 2441 2263 2445
rect 2267 2441 2268 2445
rect 2262 2440 2268 2441
rect 2358 2445 2364 2446
rect 2358 2441 2359 2445
rect 2363 2441 2364 2445
rect 2358 2440 2364 2441
rect 2454 2445 2460 2446
rect 2454 2441 2455 2445
rect 2459 2441 2460 2445
rect 2454 2440 2460 2441
rect 2526 2445 2532 2446
rect 2584 2445 2586 2457
rect 2526 2441 2527 2445
rect 2531 2441 2532 2445
rect 2526 2440 2532 2441
rect 2582 2444 2588 2445
rect 2582 2440 2583 2444
rect 2587 2440 2588 2444
rect 1366 2439 1372 2440
rect 2582 2439 2588 2440
rect 110 2431 116 2432
rect 110 2427 111 2431
rect 115 2427 116 2431
rect 110 2426 116 2427
rect 1326 2431 1332 2432
rect 1326 2427 1327 2431
rect 1331 2427 1332 2431
rect 1326 2426 1332 2427
rect 1366 2427 1372 2428
rect 112 2407 114 2426
rect 286 2422 292 2423
rect 286 2418 287 2422
rect 291 2418 292 2422
rect 286 2417 292 2418
rect 350 2422 356 2423
rect 350 2418 351 2422
rect 355 2418 356 2422
rect 350 2417 356 2418
rect 414 2422 420 2423
rect 414 2418 415 2422
rect 419 2418 420 2422
rect 414 2417 420 2418
rect 486 2422 492 2423
rect 486 2418 487 2422
rect 491 2418 492 2422
rect 486 2417 492 2418
rect 566 2422 572 2423
rect 566 2418 567 2422
rect 571 2418 572 2422
rect 566 2417 572 2418
rect 646 2422 652 2423
rect 646 2418 647 2422
rect 651 2418 652 2422
rect 646 2417 652 2418
rect 726 2422 732 2423
rect 726 2418 727 2422
rect 731 2418 732 2422
rect 726 2417 732 2418
rect 798 2422 804 2423
rect 798 2418 799 2422
rect 803 2418 804 2422
rect 798 2417 804 2418
rect 878 2422 884 2423
rect 878 2418 879 2422
rect 883 2418 884 2422
rect 878 2417 884 2418
rect 958 2422 964 2423
rect 958 2418 959 2422
rect 963 2418 964 2422
rect 958 2417 964 2418
rect 1038 2422 1044 2423
rect 1038 2418 1039 2422
rect 1043 2418 1044 2422
rect 1038 2417 1044 2418
rect 288 2407 290 2417
rect 352 2407 354 2417
rect 416 2407 418 2417
rect 488 2407 490 2417
rect 568 2407 570 2417
rect 648 2407 650 2417
rect 728 2407 730 2417
rect 800 2407 802 2417
rect 880 2407 882 2417
rect 960 2407 962 2417
rect 1040 2407 1042 2417
rect 1328 2407 1330 2426
rect 1366 2423 1367 2427
rect 1371 2423 1372 2427
rect 1366 2422 1372 2423
rect 2582 2427 2588 2428
rect 2582 2423 2583 2427
rect 2587 2423 2588 2427
rect 2582 2422 2588 2423
rect 111 2406 115 2407
rect 111 2401 115 2402
rect 247 2406 251 2407
rect 247 2401 251 2402
rect 287 2406 291 2407
rect 287 2401 291 2402
rect 335 2406 339 2407
rect 335 2401 339 2402
rect 351 2406 355 2407
rect 351 2401 355 2402
rect 415 2406 419 2407
rect 415 2401 419 2402
rect 431 2406 435 2407
rect 431 2401 435 2402
rect 487 2406 491 2407
rect 487 2401 491 2402
rect 527 2406 531 2407
rect 527 2401 531 2402
rect 567 2406 571 2407
rect 567 2401 571 2402
rect 631 2406 635 2407
rect 631 2401 635 2402
rect 647 2406 651 2407
rect 647 2401 651 2402
rect 727 2406 731 2407
rect 727 2401 731 2402
rect 799 2406 803 2407
rect 799 2401 803 2402
rect 823 2406 827 2407
rect 823 2401 827 2402
rect 879 2406 883 2407
rect 879 2401 883 2402
rect 919 2406 923 2407
rect 919 2401 923 2402
rect 959 2406 963 2407
rect 959 2401 963 2402
rect 1015 2406 1019 2407
rect 1015 2401 1019 2402
rect 1039 2406 1043 2407
rect 1039 2401 1043 2402
rect 1111 2406 1115 2407
rect 1111 2401 1115 2402
rect 1327 2406 1331 2407
rect 1368 2403 1370 2422
rect 1662 2418 1668 2419
rect 1662 2414 1663 2418
rect 1667 2414 1668 2418
rect 1662 2413 1668 2414
rect 1718 2418 1724 2419
rect 1718 2414 1719 2418
rect 1723 2414 1724 2418
rect 1718 2413 1724 2414
rect 1782 2418 1788 2419
rect 1782 2414 1783 2418
rect 1787 2414 1788 2418
rect 1782 2413 1788 2414
rect 1854 2418 1860 2419
rect 1854 2414 1855 2418
rect 1859 2414 1860 2418
rect 1854 2413 1860 2414
rect 1926 2418 1932 2419
rect 1926 2414 1927 2418
rect 1931 2414 1932 2418
rect 1926 2413 1932 2414
rect 2006 2418 2012 2419
rect 2006 2414 2007 2418
rect 2011 2414 2012 2418
rect 2006 2413 2012 2414
rect 2094 2418 2100 2419
rect 2094 2414 2095 2418
rect 2099 2414 2100 2418
rect 2094 2413 2100 2414
rect 2182 2418 2188 2419
rect 2182 2414 2183 2418
rect 2187 2414 2188 2418
rect 2182 2413 2188 2414
rect 2278 2418 2284 2419
rect 2278 2414 2279 2418
rect 2283 2414 2284 2418
rect 2278 2413 2284 2414
rect 2374 2418 2380 2419
rect 2374 2414 2375 2418
rect 2379 2414 2380 2418
rect 2374 2413 2380 2414
rect 2470 2418 2476 2419
rect 2470 2414 2471 2418
rect 2475 2414 2476 2418
rect 2470 2413 2476 2414
rect 2542 2418 2548 2419
rect 2542 2414 2543 2418
rect 2547 2414 2548 2418
rect 2542 2413 2548 2414
rect 1664 2403 1666 2413
rect 1720 2403 1722 2413
rect 1784 2403 1786 2413
rect 1856 2403 1858 2413
rect 1928 2403 1930 2413
rect 2008 2403 2010 2413
rect 2096 2403 2098 2413
rect 2184 2403 2186 2413
rect 2280 2403 2282 2413
rect 2376 2403 2378 2413
rect 2472 2403 2474 2413
rect 2544 2403 2546 2413
rect 2584 2403 2586 2422
rect 1327 2401 1331 2402
rect 1367 2402 1371 2403
rect 112 2386 114 2401
rect 248 2395 250 2401
rect 336 2395 338 2401
rect 432 2395 434 2401
rect 528 2395 530 2401
rect 632 2395 634 2401
rect 728 2395 730 2401
rect 824 2395 826 2401
rect 920 2395 922 2401
rect 1016 2395 1018 2401
rect 1112 2395 1114 2401
rect 246 2394 252 2395
rect 246 2390 247 2394
rect 251 2390 252 2394
rect 246 2389 252 2390
rect 334 2394 340 2395
rect 334 2390 335 2394
rect 339 2390 340 2394
rect 334 2389 340 2390
rect 430 2394 436 2395
rect 430 2390 431 2394
rect 435 2390 436 2394
rect 430 2389 436 2390
rect 526 2394 532 2395
rect 526 2390 527 2394
rect 531 2390 532 2394
rect 526 2389 532 2390
rect 630 2394 636 2395
rect 630 2390 631 2394
rect 635 2390 636 2394
rect 630 2389 636 2390
rect 726 2394 732 2395
rect 726 2390 727 2394
rect 731 2390 732 2394
rect 726 2389 732 2390
rect 822 2394 828 2395
rect 822 2390 823 2394
rect 827 2390 828 2394
rect 822 2389 828 2390
rect 918 2394 924 2395
rect 918 2390 919 2394
rect 923 2390 924 2394
rect 918 2389 924 2390
rect 1014 2394 1020 2395
rect 1014 2390 1015 2394
rect 1019 2390 1020 2394
rect 1014 2389 1020 2390
rect 1110 2394 1116 2395
rect 1110 2390 1111 2394
rect 1115 2390 1116 2394
rect 1110 2389 1116 2390
rect 1328 2386 1330 2401
rect 1367 2397 1371 2398
rect 1455 2402 1459 2403
rect 1455 2397 1459 2398
rect 1559 2402 1563 2403
rect 1559 2397 1563 2398
rect 1663 2402 1667 2403
rect 1663 2397 1667 2398
rect 1719 2402 1723 2403
rect 1719 2397 1723 2398
rect 1759 2402 1763 2403
rect 1759 2397 1763 2398
rect 1783 2402 1787 2403
rect 1783 2397 1787 2398
rect 1855 2402 1859 2403
rect 1855 2397 1859 2398
rect 1927 2402 1931 2403
rect 1927 2397 1931 2398
rect 1943 2402 1947 2403
rect 1943 2397 1947 2398
rect 2007 2402 2011 2403
rect 2007 2397 2011 2398
rect 2039 2402 2043 2403
rect 2039 2397 2043 2398
rect 2095 2402 2099 2403
rect 2095 2397 2099 2398
rect 2135 2402 2139 2403
rect 2135 2397 2139 2398
rect 2183 2402 2187 2403
rect 2183 2397 2187 2398
rect 2231 2402 2235 2403
rect 2231 2397 2235 2398
rect 2279 2402 2283 2403
rect 2279 2397 2283 2398
rect 2335 2402 2339 2403
rect 2335 2397 2339 2398
rect 2375 2402 2379 2403
rect 2375 2397 2379 2398
rect 2447 2402 2451 2403
rect 2447 2397 2451 2398
rect 2471 2402 2475 2403
rect 2471 2397 2475 2398
rect 2543 2402 2547 2403
rect 2543 2397 2547 2398
rect 2583 2402 2587 2403
rect 2583 2397 2587 2398
rect 110 2385 116 2386
rect 110 2381 111 2385
rect 115 2381 116 2385
rect 110 2380 116 2381
rect 1326 2385 1332 2386
rect 1326 2381 1327 2385
rect 1331 2381 1332 2385
rect 1368 2382 1370 2397
rect 1456 2391 1458 2397
rect 1560 2391 1562 2397
rect 1664 2391 1666 2397
rect 1760 2391 1762 2397
rect 1856 2391 1858 2397
rect 1944 2391 1946 2397
rect 2040 2391 2042 2397
rect 2136 2391 2138 2397
rect 2232 2391 2234 2397
rect 2336 2391 2338 2397
rect 2448 2391 2450 2397
rect 2544 2391 2546 2397
rect 1454 2390 1460 2391
rect 1454 2386 1455 2390
rect 1459 2386 1460 2390
rect 1454 2385 1460 2386
rect 1558 2390 1564 2391
rect 1558 2386 1559 2390
rect 1563 2386 1564 2390
rect 1558 2385 1564 2386
rect 1662 2390 1668 2391
rect 1662 2386 1663 2390
rect 1667 2386 1668 2390
rect 1662 2385 1668 2386
rect 1758 2390 1764 2391
rect 1758 2386 1759 2390
rect 1763 2386 1764 2390
rect 1758 2385 1764 2386
rect 1854 2390 1860 2391
rect 1854 2386 1855 2390
rect 1859 2386 1860 2390
rect 1854 2385 1860 2386
rect 1942 2390 1948 2391
rect 1942 2386 1943 2390
rect 1947 2386 1948 2390
rect 1942 2385 1948 2386
rect 2038 2390 2044 2391
rect 2038 2386 2039 2390
rect 2043 2386 2044 2390
rect 2038 2385 2044 2386
rect 2134 2390 2140 2391
rect 2134 2386 2135 2390
rect 2139 2386 2140 2390
rect 2134 2385 2140 2386
rect 2230 2390 2236 2391
rect 2230 2386 2231 2390
rect 2235 2386 2236 2390
rect 2230 2385 2236 2386
rect 2334 2390 2340 2391
rect 2334 2386 2335 2390
rect 2339 2386 2340 2390
rect 2334 2385 2340 2386
rect 2446 2390 2452 2391
rect 2446 2386 2447 2390
rect 2451 2386 2452 2390
rect 2446 2385 2452 2386
rect 2542 2390 2548 2391
rect 2542 2386 2543 2390
rect 2547 2386 2548 2390
rect 2542 2385 2548 2386
rect 2584 2382 2586 2397
rect 1326 2380 1332 2381
rect 1366 2381 1372 2382
rect 1366 2377 1367 2381
rect 1371 2377 1372 2381
rect 1366 2376 1372 2377
rect 2582 2381 2588 2382
rect 2582 2377 2583 2381
rect 2587 2377 2588 2381
rect 2582 2376 2588 2377
rect 110 2368 116 2369
rect 1326 2368 1332 2369
rect 110 2364 111 2368
rect 115 2364 116 2368
rect 110 2363 116 2364
rect 230 2367 236 2368
rect 230 2363 231 2367
rect 235 2363 236 2367
rect 112 2351 114 2363
rect 230 2362 236 2363
rect 318 2367 324 2368
rect 318 2363 319 2367
rect 323 2363 324 2367
rect 318 2362 324 2363
rect 414 2367 420 2368
rect 414 2363 415 2367
rect 419 2363 420 2367
rect 414 2362 420 2363
rect 510 2367 516 2368
rect 510 2363 511 2367
rect 515 2363 516 2367
rect 510 2362 516 2363
rect 614 2367 620 2368
rect 614 2363 615 2367
rect 619 2363 620 2367
rect 614 2362 620 2363
rect 710 2367 716 2368
rect 710 2363 711 2367
rect 715 2363 716 2367
rect 710 2362 716 2363
rect 806 2367 812 2368
rect 806 2363 807 2367
rect 811 2363 812 2367
rect 806 2362 812 2363
rect 902 2367 908 2368
rect 902 2363 903 2367
rect 907 2363 908 2367
rect 902 2362 908 2363
rect 998 2367 1004 2368
rect 998 2363 999 2367
rect 1003 2363 1004 2367
rect 998 2362 1004 2363
rect 1094 2367 1100 2368
rect 1094 2363 1095 2367
rect 1099 2363 1100 2367
rect 1326 2364 1327 2368
rect 1331 2364 1332 2368
rect 1326 2363 1332 2364
rect 1366 2364 1372 2365
rect 2582 2364 2588 2365
rect 1094 2362 1100 2363
rect 232 2351 234 2362
rect 320 2351 322 2362
rect 416 2351 418 2362
rect 512 2351 514 2362
rect 616 2351 618 2362
rect 712 2351 714 2362
rect 808 2351 810 2362
rect 904 2351 906 2362
rect 1000 2351 1002 2362
rect 1096 2351 1098 2362
rect 1328 2351 1330 2363
rect 1366 2360 1367 2364
rect 1371 2360 1372 2364
rect 1366 2359 1372 2360
rect 1438 2363 1444 2364
rect 1438 2359 1439 2363
rect 1443 2359 1444 2363
rect 111 2350 115 2351
rect 111 2345 115 2346
rect 159 2350 163 2351
rect 159 2345 163 2346
rect 231 2350 235 2351
rect 231 2345 235 2346
rect 263 2350 267 2351
rect 263 2345 267 2346
rect 319 2350 323 2351
rect 319 2345 323 2346
rect 375 2350 379 2351
rect 375 2345 379 2346
rect 415 2350 419 2351
rect 415 2345 419 2346
rect 487 2350 491 2351
rect 487 2345 491 2346
rect 511 2350 515 2351
rect 511 2345 515 2346
rect 599 2350 603 2351
rect 599 2345 603 2346
rect 615 2350 619 2351
rect 615 2345 619 2346
rect 711 2350 715 2351
rect 711 2345 715 2346
rect 807 2350 811 2351
rect 807 2345 811 2346
rect 815 2350 819 2351
rect 815 2345 819 2346
rect 903 2350 907 2351
rect 903 2345 907 2346
rect 911 2350 915 2351
rect 911 2345 915 2346
rect 999 2350 1003 2351
rect 999 2345 1003 2346
rect 1007 2350 1011 2351
rect 1007 2345 1011 2346
rect 1095 2350 1099 2351
rect 1095 2345 1099 2346
rect 1103 2350 1107 2351
rect 1103 2345 1107 2346
rect 1199 2350 1203 2351
rect 1199 2345 1203 2346
rect 1327 2350 1331 2351
rect 1368 2347 1370 2359
rect 1438 2358 1444 2359
rect 1542 2363 1548 2364
rect 1542 2359 1543 2363
rect 1547 2359 1548 2363
rect 1542 2358 1548 2359
rect 1646 2363 1652 2364
rect 1646 2359 1647 2363
rect 1651 2359 1652 2363
rect 1646 2358 1652 2359
rect 1742 2363 1748 2364
rect 1742 2359 1743 2363
rect 1747 2359 1748 2363
rect 1742 2358 1748 2359
rect 1838 2363 1844 2364
rect 1838 2359 1839 2363
rect 1843 2359 1844 2363
rect 1838 2358 1844 2359
rect 1926 2363 1932 2364
rect 1926 2359 1927 2363
rect 1931 2359 1932 2363
rect 1926 2358 1932 2359
rect 2022 2363 2028 2364
rect 2022 2359 2023 2363
rect 2027 2359 2028 2363
rect 2022 2358 2028 2359
rect 2118 2363 2124 2364
rect 2118 2359 2119 2363
rect 2123 2359 2124 2363
rect 2118 2358 2124 2359
rect 2214 2363 2220 2364
rect 2214 2359 2215 2363
rect 2219 2359 2220 2363
rect 2214 2358 2220 2359
rect 2318 2363 2324 2364
rect 2318 2359 2319 2363
rect 2323 2359 2324 2363
rect 2318 2358 2324 2359
rect 2430 2363 2436 2364
rect 2430 2359 2431 2363
rect 2435 2359 2436 2363
rect 2430 2358 2436 2359
rect 2526 2363 2532 2364
rect 2526 2359 2527 2363
rect 2531 2359 2532 2363
rect 2582 2360 2583 2364
rect 2587 2360 2588 2364
rect 2582 2359 2588 2360
rect 2526 2358 2532 2359
rect 1440 2347 1442 2358
rect 1544 2347 1546 2358
rect 1648 2347 1650 2358
rect 1744 2347 1746 2358
rect 1840 2347 1842 2358
rect 1928 2347 1930 2358
rect 2024 2347 2026 2358
rect 2120 2347 2122 2358
rect 2216 2347 2218 2358
rect 2320 2347 2322 2358
rect 2432 2347 2434 2358
rect 2528 2347 2530 2358
rect 2584 2347 2586 2359
rect 1327 2345 1331 2346
rect 1367 2346 1371 2347
rect 112 2333 114 2345
rect 160 2334 162 2345
rect 264 2334 266 2345
rect 376 2334 378 2345
rect 488 2334 490 2345
rect 600 2334 602 2345
rect 712 2334 714 2345
rect 816 2334 818 2345
rect 912 2334 914 2345
rect 1008 2334 1010 2345
rect 1104 2334 1106 2345
rect 1200 2334 1202 2345
rect 158 2333 164 2334
rect 110 2332 116 2333
rect 110 2328 111 2332
rect 115 2328 116 2332
rect 158 2329 159 2333
rect 163 2329 164 2333
rect 158 2328 164 2329
rect 262 2333 268 2334
rect 262 2329 263 2333
rect 267 2329 268 2333
rect 262 2328 268 2329
rect 374 2333 380 2334
rect 374 2329 375 2333
rect 379 2329 380 2333
rect 374 2328 380 2329
rect 486 2333 492 2334
rect 486 2329 487 2333
rect 491 2329 492 2333
rect 486 2328 492 2329
rect 598 2333 604 2334
rect 598 2329 599 2333
rect 603 2329 604 2333
rect 598 2328 604 2329
rect 710 2333 716 2334
rect 710 2329 711 2333
rect 715 2329 716 2333
rect 710 2328 716 2329
rect 814 2333 820 2334
rect 814 2329 815 2333
rect 819 2329 820 2333
rect 814 2328 820 2329
rect 910 2333 916 2334
rect 910 2329 911 2333
rect 915 2329 916 2333
rect 910 2328 916 2329
rect 1006 2333 1012 2334
rect 1006 2329 1007 2333
rect 1011 2329 1012 2333
rect 1006 2328 1012 2329
rect 1102 2333 1108 2334
rect 1102 2329 1103 2333
rect 1107 2329 1108 2333
rect 1102 2328 1108 2329
rect 1198 2333 1204 2334
rect 1328 2333 1330 2345
rect 1367 2341 1371 2342
rect 1399 2346 1403 2347
rect 1399 2341 1403 2342
rect 1439 2346 1443 2347
rect 1439 2341 1443 2342
rect 1455 2346 1459 2347
rect 1455 2341 1459 2342
rect 1511 2346 1515 2347
rect 1511 2341 1515 2342
rect 1543 2346 1547 2347
rect 1543 2341 1547 2342
rect 1567 2346 1571 2347
rect 1567 2341 1571 2342
rect 1639 2346 1643 2347
rect 1639 2341 1643 2342
rect 1647 2346 1651 2347
rect 1647 2341 1651 2342
rect 1727 2346 1731 2347
rect 1727 2341 1731 2342
rect 1743 2346 1747 2347
rect 1743 2341 1747 2342
rect 1823 2346 1827 2347
rect 1823 2341 1827 2342
rect 1839 2346 1843 2347
rect 1839 2341 1843 2342
rect 1927 2346 1931 2347
rect 1927 2341 1931 2342
rect 1943 2346 1947 2347
rect 1943 2341 1947 2342
rect 2023 2346 2027 2347
rect 2023 2341 2027 2342
rect 2079 2346 2083 2347
rect 2079 2341 2083 2342
rect 2119 2346 2123 2347
rect 2119 2341 2123 2342
rect 2215 2346 2219 2347
rect 2215 2341 2219 2342
rect 2223 2346 2227 2347
rect 2223 2341 2227 2342
rect 2319 2346 2323 2347
rect 2319 2341 2323 2342
rect 2383 2346 2387 2347
rect 2383 2341 2387 2342
rect 2431 2346 2435 2347
rect 2431 2341 2435 2342
rect 2527 2346 2531 2347
rect 2527 2341 2531 2342
rect 2583 2346 2587 2347
rect 2583 2341 2587 2342
rect 1198 2329 1199 2333
rect 1203 2329 1204 2333
rect 1198 2328 1204 2329
rect 1326 2332 1332 2333
rect 1326 2328 1327 2332
rect 1331 2328 1332 2332
rect 1368 2329 1370 2341
rect 1400 2330 1402 2341
rect 1456 2330 1458 2341
rect 1512 2330 1514 2341
rect 1568 2330 1570 2341
rect 1640 2330 1642 2341
rect 1728 2330 1730 2341
rect 1824 2330 1826 2341
rect 1944 2330 1946 2341
rect 2080 2330 2082 2341
rect 2224 2330 2226 2341
rect 2384 2330 2386 2341
rect 2528 2330 2530 2341
rect 1398 2329 1404 2330
rect 110 2327 116 2328
rect 1326 2327 1332 2328
rect 1366 2328 1372 2329
rect 1366 2324 1367 2328
rect 1371 2324 1372 2328
rect 1398 2325 1399 2329
rect 1403 2325 1404 2329
rect 1398 2324 1404 2325
rect 1454 2329 1460 2330
rect 1454 2325 1455 2329
rect 1459 2325 1460 2329
rect 1454 2324 1460 2325
rect 1510 2329 1516 2330
rect 1510 2325 1511 2329
rect 1515 2325 1516 2329
rect 1510 2324 1516 2325
rect 1566 2329 1572 2330
rect 1566 2325 1567 2329
rect 1571 2325 1572 2329
rect 1566 2324 1572 2325
rect 1638 2329 1644 2330
rect 1638 2325 1639 2329
rect 1643 2325 1644 2329
rect 1638 2324 1644 2325
rect 1726 2329 1732 2330
rect 1726 2325 1727 2329
rect 1731 2325 1732 2329
rect 1726 2324 1732 2325
rect 1822 2329 1828 2330
rect 1822 2325 1823 2329
rect 1827 2325 1828 2329
rect 1822 2324 1828 2325
rect 1942 2329 1948 2330
rect 1942 2325 1943 2329
rect 1947 2325 1948 2329
rect 1942 2324 1948 2325
rect 2078 2329 2084 2330
rect 2078 2325 2079 2329
rect 2083 2325 2084 2329
rect 2078 2324 2084 2325
rect 2222 2329 2228 2330
rect 2222 2325 2223 2329
rect 2227 2325 2228 2329
rect 2222 2324 2228 2325
rect 2382 2329 2388 2330
rect 2382 2325 2383 2329
rect 2387 2325 2388 2329
rect 2382 2324 2388 2325
rect 2526 2329 2532 2330
rect 2584 2329 2586 2341
rect 2526 2325 2527 2329
rect 2531 2325 2532 2329
rect 2526 2324 2532 2325
rect 2582 2328 2588 2329
rect 2582 2324 2583 2328
rect 2587 2324 2588 2328
rect 1366 2323 1372 2324
rect 2582 2323 2588 2324
rect 110 2315 116 2316
rect 110 2311 111 2315
rect 115 2311 116 2315
rect 110 2310 116 2311
rect 1326 2315 1332 2316
rect 1326 2311 1327 2315
rect 1331 2311 1332 2315
rect 1326 2310 1332 2311
rect 1366 2311 1372 2312
rect 112 2291 114 2310
rect 174 2306 180 2307
rect 174 2302 175 2306
rect 179 2302 180 2306
rect 174 2301 180 2302
rect 278 2306 284 2307
rect 278 2302 279 2306
rect 283 2302 284 2306
rect 278 2301 284 2302
rect 390 2306 396 2307
rect 390 2302 391 2306
rect 395 2302 396 2306
rect 390 2301 396 2302
rect 502 2306 508 2307
rect 502 2302 503 2306
rect 507 2302 508 2306
rect 502 2301 508 2302
rect 614 2306 620 2307
rect 614 2302 615 2306
rect 619 2302 620 2306
rect 614 2301 620 2302
rect 726 2306 732 2307
rect 726 2302 727 2306
rect 731 2302 732 2306
rect 726 2301 732 2302
rect 830 2306 836 2307
rect 830 2302 831 2306
rect 835 2302 836 2306
rect 830 2301 836 2302
rect 926 2306 932 2307
rect 926 2302 927 2306
rect 931 2302 932 2306
rect 926 2301 932 2302
rect 1022 2306 1028 2307
rect 1022 2302 1023 2306
rect 1027 2302 1028 2306
rect 1022 2301 1028 2302
rect 1118 2306 1124 2307
rect 1118 2302 1119 2306
rect 1123 2302 1124 2306
rect 1118 2301 1124 2302
rect 1214 2306 1220 2307
rect 1214 2302 1215 2306
rect 1219 2302 1220 2306
rect 1214 2301 1220 2302
rect 176 2291 178 2301
rect 280 2291 282 2301
rect 392 2291 394 2301
rect 504 2291 506 2301
rect 616 2291 618 2301
rect 728 2291 730 2301
rect 832 2291 834 2301
rect 928 2291 930 2301
rect 1024 2291 1026 2301
rect 1120 2291 1122 2301
rect 1216 2291 1218 2301
rect 1328 2291 1330 2310
rect 1366 2307 1367 2311
rect 1371 2307 1372 2311
rect 1366 2306 1372 2307
rect 2582 2311 2588 2312
rect 2582 2307 2583 2311
rect 2587 2307 2588 2311
rect 2582 2306 2588 2307
rect 111 2290 115 2291
rect 111 2285 115 2286
rect 159 2290 163 2291
rect 159 2285 163 2286
rect 175 2290 179 2291
rect 175 2285 179 2286
rect 247 2290 251 2291
rect 247 2285 251 2286
rect 279 2290 283 2291
rect 279 2285 283 2286
rect 375 2290 379 2291
rect 375 2285 379 2286
rect 391 2290 395 2291
rect 391 2285 395 2286
rect 503 2290 507 2291
rect 503 2285 507 2286
rect 511 2290 515 2291
rect 511 2285 515 2286
rect 615 2290 619 2291
rect 615 2285 619 2286
rect 639 2290 643 2291
rect 639 2285 643 2286
rect 727 2290 731 2291
rect 727 2285 731 2286
rect 767 2290 771 2291
rect 767 2285 771 2286
rect 831 2290 835 2291
rect 831 2285 835 2286
rect 887 2290 891 2291
rect 887 2285 891 2286
rect 927 2290 931 2291
rect 927 2285 931 2286
rect 999 2290 1003 2291
rect 999 2285 1003 2286
rect 1023 2290 1027 2291
rect 1023 2285 1027 2286
rect 1103 2290 1107 2291
rect 1103 2285 1107 2286
rect 1119 2290 1123 2291
rect 1119 2285 1123 2286
rect 1207 2290 1211 2291
rect 1207 2285 1211 2286
rect 1215 2290 1219 2291
rect 1215 2285 1219 2286
rect 1287 2290 1291 2291
rect 1287 2285 1291 2286
rect 1327 2290 1331 2291
rect 1327 2285 1331 2286
rect 112 2270 114 2285
rect 160 2279 162 2285
rect 248 2279 250 2285
rect 376 2279 378 2285
rect 512 2279 514 2285
rect 640 2279 642 2285
rect 768 2279 770 2285
rect 888 2279 890 2285
rect 1000 2279 1002 2285
rect 1104 2279 1106 2285
rect 1208 2279 1210 2285
rect 1288 2279 1290 2285
rect 158 2278 164 2279
rect 158 2274 159 2278
rect 163 2274 164 2278
rect 158 2273 164 2274
rect 246 2278 252 2279
rect 246 2274 247 2278
rect 251 2274 252 2278
rect 246 2273 252 2274
rect 374 2278 380 2279
rect 374 2274 375 2278
rect 379 2274 380 2278
rect 374 2273 380 2274
rect 510 2278 516 2279
rect 510 2274 511 2278
rect 515 2274 516 2278
rect 510 2273 516 2274
rect 638 2278 644 2279
rect 638 2274 639 2278
rect 643 2274 644 2278
rect 638 2273 644 2274
rect 766 2278 772 2279
rect 766 2274 767 2278
rect 771 2274 772 2278
rect 766 2273 772 2274
rect 886 2278 892 2279
rect 886 2274 887 2278
rect 891 2274 892 2278
rect 886 2273 892 2274
rect 998 2278 1004 2279
rect 998 2274 999 2278
rect 1003 2274 1004 2278
rect 998 2273 1004 2274
rect 1102 2278 1108 2279
rect 1102 2274 1103 2278
rect 1107 2274 1108 2278
rect 1102 2273 1108 2274
rect 1206 2278 1212 2279
rect 1206 2274 1207 2278
rect 1211 2274 1212 2278
rect 1206 2273 1212 2274
rect 1286 2278 1292 2279
rect 1286 2274 1287 2278
rect 1291 2274 1292 2278
rect 1286 2273 1292 2274
rect 1328 2270 1330 2285
rect 1368 2283 1370 2306
rect 1414 2302 1420 2303
rect 1414 2298 1415 2302
rect 1419 2298 1420 2302
rect 1414 2297 1420 2298
rect 1470 2302 1476 2303
rect 1470 2298 1471 2302
rect 1475 2298 1476 2302
rect 1470 2297 1476 2298
rect 1526 2302 1532 2303
rect 1526 2298 1527 2302
rect 1531 2298 1532 2302
rect 1526 2297 1532 2298
rect 1582 2302 1588 2303
rect 1582 2298 1583 2302
rect 1587 2298 1588 2302
rect 1582 2297 1588 2298
rect 1654 2302 1660 2303
rect 1654 2298 1655 2302
rect 1659 2298 1660 2302
rect 1654 2297 1660 2298
rect 1742 2302 1748 2303
rect 1742 2298 1743 2302
rect 1747 2298 1748 2302
rect 1742 2297 1748 2298
rect 1838 2302 1844 2303
rect 1838 2298 1839 2302
rect 1843 2298 1844 2302
rect 1838 2297 1844 2298
rect 1958 2302 1964 2303
rect 1958 2298 1959 2302
rect 1963 2298 1964 2302
rect 1958 2297 1964 2298
rect 2094 2302 2100 2303
rect 2094 2298 2095 2302
rect 2099 2298 2100 2302
rect 2094 2297 2100 2298
rect 2238 2302 2244 2303
rect 2238 2298 2239 2302
rect 2243 2298 2244 2302
rect 2238 2297 2244 2298
rect 2398 2302 2404 2303
rect 2398 2298 2399 2302
rect 2403 2298 2404 2302
rect 2398 2297 2404 2298
rect 2542 2302 2548 2303
rect 2542 2298 2543 2302
rect 2547 2298 2548 2302
rect 2542 2297 2548 2298
rect 1416 2283 1418 2297
rect 1472 2283 1474 2297
rect 1528 2283 1530 2297
rect 1584 2283 1586 2297
rect 1656 2283 1658 2297
rect 1744 2283 1746 2297
rect 1840 2283 1842 2297
rect 1960 2283 1962 2297
rect 2096 2283 2098 2297
rect 2240 2283 2242 2297
rect 2400 2283 2402 2297
rect 2544 2283 2546 2297
rect 2584 2283 2586 2306
rect 1367 2282 1371 2283
rect 1367 2277 1371 2278
rect 1415 2282 1419 2283
rect 1415 2277 1419 2278
rect 1471 2282 1475 2283
rect 1471 2277 1475 2278
rect 1495 2282 1499 2283
rect 1495 2277 1499 2278
rect 1527 2282 1531 2283
rect 1527 2277 1531 2278
rect 1583 2282 1587 2283
rect 1583 2277 1587 2278
rect 1615 2282 1619 2283
rect 1615 2277 1619 2278
rect 1655 2282 1659 2283
rect 1655 2277 1659 2278
rect 1735 2282 1739 2283
rect 1735 2277 1739 2278
rect 1743 2282 1747 2283
rect 1743 2277 1747 2278
rect 1839 2282 1843 2283
rect 1839 2277 1843 2278
rect 1855 2282 1859 2283
rect 1855 2277 1859 2278
rect 1959 2282 1963 2283
rect 1959 2277 1963 2278
rect 1967 2282 1971 2283
rect 1967 2277 1971 2278
rect 2071 2282 2075 2283
rect 2071 2277 2075 2278
rect 2095 2282 2099 2283
rect 2095 2277 2099 2278
rect 2167 2282 2171 2283
rect 2167 2277 2171 2278
rect 2239 2282 2243 2283
rect 2239 2277 2243 2278
rect 2255 2282 2259 2283
rect 2255 2277 2259 2278
rect 2335 2282 2339 2283
rect 2335 2277 2339 2278
rect 2399 2282 2403 2283
rect 2399 2277 2403 2278
rect 2407 2282 2411 2283
rect 2407 2277 2411 2278
rect 2487 2282 2491 2283
rect 2487 2277 2491 2278
rect 2543 2282 2547 2283
rect 2543 2277 2547 2278
rect 2583 2282 2587 2283
rect 2583 2277 2587 2278
rect 110 2269 116 2270
rect 110 2265 111 2269
rect 115 2265 116 2269
rect 110 2264 116 2265
rect 1326 2269 1332 2270
rect 1326 2265 1327 2269
rect 1331 2265 1332 2269
rect 1326 2264 1332 2265
rect 1368 2262 1370 2277
rect 1416 2271 1418 2277
rect 1496 2271 1498 2277
rect 1616 2271 1618 2277
rect 1736 2271 1738 2277
rect 1856 2271 1858 2277
rect 1968 2271 1970 2277
rect 2072 2271 2074 2277
rect 2168 2271 2170 2277
rect 2256 2271 2258 2277
rect 2336 2271 2338 2277
rect 2408 2271 2410 2277
rect 2488 2271 2490 2277
rect 2544 2271 2546 2277
rect 1414 2270 1420 2271
rect 1414 2266 1415 2270
rect 1419 2266 1420 2270
rect 1414 2265 1420 2266
rect 1494 2270 1500 2271
rect 1494 2266 1495 2270
rect 1499 2266 1500 2270
rect 1494 2265 1500 2266
rect 1614 2270 1620 2271
rect 1614 2266 1615 2270
rect 1619 2266 1620 2270
rect 1614 2265 1620 2266
rect 1734 2270 1740 2271
rect 1734 2266 1735 2270
rect 1739 2266 1740 2270
rect 1734 2265 1740 2266
rect 1854 2270 1860 2271
rect 1854 2266 1855 2270
rect 1859 2266 1860 2270
rect 1854 2265 1860 2266
rect 1966 2270 1972 2271
rect 1966 2266 1967 2270
rect 1971 2266 1972 2270
rect 1966 2265 1972 2266
rect 2070 2270 2076 2271
rect 2070 2266 2071 2270
rect 2075 2266 2076 2270
rect 2070 2265 2076 2266
rect 2166 2270 2172 2271
rect 2166 2266 2167 2270
rect 2171 2266 2172 2270
rect 2166 2265 2172 2266
rect 2254 2270 2260 2271
rect 2254 2266 2255 2270
rect 2259 2266 2260 2270
rect 2254 2265 2260 2266
rect 2334 2270 2340 2271
rect 2334 2266 2335 2270
rect 2339 2266 2340 2270
rect 2334 2265 2340 2266
rect 2406 2270 2412 2271
rect 2406 2266 2407 2270
rect 2411 2266 2412 2270
rect 2406 2265 2412 2266
rect 2486 2270 2492 2271
rect 2486 2266 2487 2270
rect 2491 2266 2492 2270
rect 2486 2265 2492 2266
rect 2542 2270 2548 2271
rect 2542 2266 2543 2270
rect 2547 2266 2548 2270
rect 2542 2265 2548 2266
rect 2584 2262 2586 2277
rect 1366 2261 1372 2262
rect 1366 2257 1367 2261
rect 1371 2257 1372 2261
rect 1366 2256 1372 2257
rect 2582 2261 2588 2262
rect 2582 2257 2583 2261
rect 2587 2257 2588 2261
rect 2582 2256 2588 2257
rect 110 2252 116 2253
rect 1326 2252 1332 2253
rect 110 2248 111 2252
rect 115 2248 116 2252
rect 110 2247 116 2248
rect 142 2251 148 2252
rect 142 2247 143 2251
rect 147 2247 148 2251
rect 112 2227 114 2247
rect 142 2246 148 2247
rect 230 2251 236 2252
rect 230 2247 231 2251
rect 235 2247 236 2251
rect 230 2246 236 2247
rect 358 2251 364 2252
rect 358 2247 359 2251
rect 363 2247 364 2251
rect 358 2246 364 2247
rect 494 2251 500 2252
rect 494 2247 495 2251
rect 499 2247 500 2251
rect 494 2246 500 2247
rect 622 2251 628 2252
rect 622 2247 623 2251
rect 627 2247 628 2251
rect 622 2246 628 2247
rect 750 2251 756 2252
rect 750 2247 751 2251
rect 755 2247 756 2251
rect 750 2246 756 2247
rect 870 2251 876 2252
rect 870 2247 871 2251
rect 875 2247 876 2251
rect 870 2246 876 2247
rect 982 2251 988 2252
rect 982 2247 983 2251
rect 987 2247 988 2251
rect 982 2246 988 2247
rect 1086 2251 1092 2252
rect 1086 2247 1087 2251
rect 1091 2247 1092 2251
rect 1086 2246 1092 2247
rect 1190 2251 1196 2252
rect 1190 2247 1191 2251
rect 1195 2247 1196 2251
rect 1190 2246 1196 2247
rect 1270 2251 1276 2252
rect 1270 2247 1271 2251
rect 1275 2247 1276 2251
rect 1326 2248 1327 2252
rect 1331 2248 1332 2252
rect 1326 2247 1332 2248
rect 1270 2246 1276 2247
rect 144 2227 146 2246
rect 232 2227 234 2246
rect 360 2227 362 2246
rect 496 2227 498 2246
rect 624 2227 626 2246
rect 752 2227 754 2246
rect 872 2227 874 2246
rect 984 2227 986 2246
rect 1088 2227 1090 2246
rect 1192 2227 1194 2246
rect 1272 2227 1274 2246
rect 1328 2227 1330 2247
rect 1366 2244 1372 2245
rect 2582 2244 2588 2245
rect 1366 2240 1367 2244
rect 1371 2240 1372 2244
rect 1366 2239 1372 2240
rect 1398 2243 1404 2244
rect 1398 2239 1399 2243
rect 1403 2239 1404 2243
rect 111 2226 115 2227
rect 111 2221 115 2222
rect 143 2226 147 2227
rect 143 2221 147 2222
rect 231 2226 235 2227
rect 231 2221 235 2222
rect 359 2226 363 2227
rect 359 2221 363 2222
rect 495 2226 499 2227
rect 495 2221 499 2222
rect 623 2226 627 2227
rect 623 2221 627 2222
rect 751 2226 755 2227
rect 751 2221 755 2222
rect 871 2226 875 2227
rect 871 2221 875 2222
rect 983 2226 987 2227
rect 983 2221 987 2222
rect 1087 2226 1091 2227
rect 1087 2221 1091 2222
rect 1191 2226 1195 2227
rect 1191 2221 1195 2222
rect 1271 2226 1275 2227
rect 1271 2221 1275 2222
rect 1327 2226 1331 2227
rect 1327 2221 1331 2222
rect 112 2209 114 2221
rect 144 2210 146 2221
rect 232 2210 234 2221
rect 360 2210 362 2221
rect 496 2210 498 2221
rect 624 2210 626 2221
rect 752 2210 754 2221
rect 872 2210 874 2221
rect 984 2210 986 2221
rect 1088 2210 1090 2221
rect 1192 2210 1194 2221
rect 1272 2210 1274 2221
rect 142 2209 148 2210
rect 110 2208 116 2209
rect 110 2204 111 2208
rect 115 2204 116 2208
rect 142 2205 143 2209
rect 147 2205 148 2209
rect 142 2204 148 2205
rect 230 2209 236 2210
rect 230 2205 231 2209
rect 235 2205 236 2209
rect 230 2204 236 2205
rect 358 2209 364 2210
rect 358 2205 359 2209
rect 363 2205 364 2209
rect 358 2204 364 2205
rect 494 2209 500 2210
rect 494 2205 495 2209
rect 499 2205 500 2209
rect 494 2204 500 2205
rect 622 2209 628 2210
rect 622 2205 623 2209
rect 627 2205 628 2209
rect 622 2204 628 2205
rect 750 2209 756 2210
rect 750 2205 751 2209
rect 755 2205 756 2209
rect 750 2204 756 2205
rect 870 2209 876 2210
rect 870 2205 871 2209
rect 875 2205 876 2209
rect 870 2204 876 2205
rect 982 2209 988 2210
rect 982 2205 983 2209
rect 987 2205 988 2209
rect 982 2204 988 2205
rect 1086 2209 1092 2210
rect 1086 2205 1087 2209
rect 1091 2205 1092 2209
rect 1086 2204 1092 2205
rect 1190 2209 1196 2210
rect 1190 2205 1191 2209
rect 1195 2205 1196 2209
rect 1190 2204 1196 2205
rect 1270 2209 1276 2210
rect 1328 2209 1330 2221
rect 1368 2215 1370 2239
rect 1398 2238 1404 2239
rect 1478 2243 1484 2244
rect 1478 2239 1479 2243
rect 1483 2239 1484 2243
rect 1478 2238 1484 2239
rect 1598 2243 1604 2244
rect 1598 2239 1599 2243
rect 1603 2239 1604 2243
rect 1598 2238 1604 2239
rect 1718 2243 1724 2244
rect 1718 2239 1719 2243
rect 1723 2239 1724 2243
rect 1718 2238 1724 2239
rect 1838 2243 1844 2244
rect 1838 2239 1839 2243
rect 1843 2239 1844 2243
rect 1838 2238 1844 2239
rect 1950 2243 1956 2244
rect 1950 2239 1951 2243
rect 1955 2239 1956 2243
rect 1950 2238 1956 2239
rect 2054 2243 2060 2244
rect 2054 2239 2055 2243
rect 2059 2239 2060 2243
rect 2054 2238 2060 2239
rect 2150 2243 2156 2244
rect 2150 2239 2151 2243
rect 2155 2239 2156 2243
rect 2150 2238 2156 2239
rect 2238 2243 2244 2244
rect 2238 2239 2239 2243
rect 2243 2239 2244 2243
rect 2238 2238 2244 2239
rect 2318 2243 2324 2244
rect 2318 2239 2319 2243
rect 2323 2239 2324 2243
rect 2318 2238 2324 2239
rect 2390 2243 2396 2244
rect 2390 2239 2391 2243
rect 2395 2239 2396 2243
rect 2390 2238 2396 2239
rect 2470 2243 2476 2244
rect 2470 2239 2471 2243
rect 2475 2239 2476 2243
rect 2470 2238 2476 2239
rect 2526 2243 2532 2244
rect 2526 2239 2527 2243
rect 2531 2239 2532 2243
rect 2582 2240 2583 2244
rect 2587 2240 2588 2244
rect 2582 2239 2588 2240
rect 2526 2238 2532 2239
rect 1400 2215 1402 2238
rect 1480 2215 1482 2238
rect 1600 2215 1602 2238
rect 1720 2215 1722 2238
rect 1840 2215 1842 2238
rect 1952 2215 1954 2238
rect 2056 2215 2058 2238
rect 2152 2215 2154 2238
rect 2240 2215 2242 2238
rect 2320 2215 2322 2238
rect 2392 2215 2394 2238
rect 2472 2215 2474 2238
rect 2528 2215 2530 2238
rect 2584 2215 2586 2239
rect 1367 2214 1371 2215
rect 1367 2209 1371 2210
rect 1399 2214 1403 2215
rect 1399 2209 1403 2210
rect 1455 2214 1459 2215
rect 1455 2209 1459 2210
rect 1479 2214 1483 2215
rect 1479 2209 1483 2210
rect 1535 2214 1539 2215
rect 1535 2209 1539 2210
rect 1599 2214 1603 2215
rect 1599 2209 1603 2210
rect 1631 2214 1635 2215
rect 1631 2209 1635 2210
rect 1719 2214 1723 2215
rect 1719 2209 1723 2210
rect 1743 2214 1747 2215
rect 1743 2209 1747 2210
rect 1839 2214 1843 2215
rect 1839 2209 1843 2210
rect 1863 2214 1867 2215
rect 1863 2209 1867 2210
rect 1951 2214 1955 2215
rect 1951 2209 1955 2210
rect 1983 2214 1987 2215
rect 1983 2209 1987 2210
rect 2055 2214 2059 2215
rect 2055 2209 2059 2210
rect 2095 2214 2099 2215
rect 2095 2209 2099 2210
rect 2151 2214 2155 2215
rect 2151 2209 2155 2210
rect 2207 2214 2211 2215
rect 2207 2209 2211 2210
rect 2239 2214 2243 2215
rect 2239 2209 2243 2210
rect 2311 2214 2315 2215
rect 2311 2209 2315 2210
rect 2319 2214 2323 2215
rect 2319 2209 2323 2210
rect 2391 2214 2395 2215
rect 2391 2209 2395 2210
rect 2423 2214 2427 2215
rect 2423 2209 2427 2210
rect 2471 2214 2475 2215
rect 2471 2209 2475 2210
rect 2527 2214 2531 2215
rect 2527 2209 2531 2210
rect 2583 2214 2587 2215
rect 2583 2209 2587 2210
rect 1270 2205 1271 2209
rect 1275 2205 1276 2209
rect 1270 2204 1276 2205
rect 1326 2208 1332 2209
rect 1326 2204 1327 2208
rect 1331 2204 1332 2208
rect 110 2203 116 2204
rect 1326 2203 1332 2204
rect 1368 2197 1370 2209
rect 1456 2198 1458 2209
rect 1536 2198 1538 2209
rect 1632 2198 1634 2209
rect 1744 2198 1746 2209
rect 1864 2198 1866 2209
rect 1984 2198 1986 2209
rect 2096 2198 2098 2209
rect 2208 2198 2210 2209
rect 2312 2198 2314 2209
rect 2424 2198 2426 2209
rect 2528 2198 2530 2209
rect 1454 2197 1460 2198
rect 1366 2196 1372 2197
rect 1366 2192 1367 2196
rect 1371 2192 1372 2196
rect 1454 2193 1455 2197
rect 1459 2193 1460 2197
rect 1454 2192 1460 2193
rect 1534 2197 1540 2198
rect 1534 2193 1535 2197
rect 1539 2193 1540 2197
rect 1534 2192 1540 2193
rect 1630 2197 1636 2198
rect 1630 2193 1631 2197
rect 1635 2193 1636 2197
rect 1630 2192 1636 2193
rect 1742 2197 1748 2198
rect 1742 2193 1743 2197
rect 1747 2193 1748 2197
rect 1742 2192 1748 2193
rect 1862 2197 1868 2198
rect 1862 2193 1863 2197
rect 1867 2193 1868 2197
rect 1862 2192 1868 2193
rect 1982 2197 1988 2198
rect 1982 2193 1983 2197
rect 1987 2193 1988 2197
rect 1982 2192 1988 2193
rect 2094 2197 2100 2198
rect 2094 2193 2095 2197
rect 2099 2193 2100 2197
rect 2094 2192 2100 2193
rect 2206 2197 2212 2198
rect 2206 2193 2207 2197
rect 2211 2193 2212 2197
rect 2206 2192 2212 2193
rect 2310 2197 2316 2198
rect 2310 2193 2311 2197
rect 2315 2193 2316 2197
rect 2310 2192 2316 2193
rect 2422 2197 2428 2198
rect 2422 2193 2423 2197
rect 2427 2193 2428 2197
rect 2422 2192 2428 2193
rect 2526 2197 2532 2198
rect 2584 2197 2586 2209
rect 2526 2193 2527 2197
rect 2531 2193 2532 2197
rect 2526 2192 2532 2193
rect 2582 2196 2588 2197
rect 2582 2192 2583 2196
rect 2587 2192 2588 2196
rect 110 2191 116 2192
rect 110 2187 111 2191
rect 115 2187 116 2191
rect 110 2186 116 2187
rect 1326 2191 1332 2192
rect 1366 2191 1372 2192
rect 2582 2191 2588 2192
rect 1326 2187 1327 2191
rect 1331 2187 1332 2191
rect 1326 2186 1332 2187
rect 112 2167 114 2186
rect 158 2182 164 2183
rect 158 2178 159 2182
rect 163 2178 164 2182
rect 158 2177 164 2178
rect 246 2182 252 2183
rect 246 2178 247 2182
rect 251 2178 252 2182
rect 246 2177 252 2178
rect 374 2182 380 2183
rect 374 2178 375 2182
rect 379 2178 380 2182
rect 374 2177 380 2178
rect 510 2182 516 2183
rect 510 2178 511 2182
rect 515 2178 516 2182
rect 510 2177 516 2178
rect 638 2182 644 2183
rect 638 2178 639 2182
rect 643 2178 644 2182
rect 638 2177 644 2178
rect 766 2182 772 2183
rect 766 2178 767 2182
rect 771 2178 772 2182
rect 766 2177 772 2178
rect 886 2182 892 2183
rect 886 2178 887 2182
rect 891 2178 892 2182
rect 886 2177 892 2178
rect 998 2182 1004 2183
rect 998 2178 999 2182
rect 1003 2178 1004 2182
rect 998 2177 1004 2178
rect 1102 2182 1108 2183
rect 1102 2178 1103 2182
rect 1107 2178 1108 2182
rect 1102 2177 1108 2178
rect 1206 2182 1212 2183
rect 1206 2178 1207 2182
rect 1211 2178 1212 2182
rect 1206 2177 1212 2178
rect 1286 2182 1292 2183
rect 1286 2178 1287 2182
rect 1291 2178 1292 2182
rect 1286 2177 1292 2178
rect 160 2167 162 2177
rect 248 2167 250 2177
rect 376 2167 378 2177
rect 512 2167 514 2177
rect 640 2167 642 2177
rect 768 2167 770 2177
rect 888 2167 890 2177
rect 1000 2167 1002 2177
rect 1104 2167 1106 2177
rect 1208 2167 1210 2177
rect 1288 2167 1290 2177
rect 1328 2167 1330 2186
rect 1366 2179 1372 2180
rect 1366 2175 1367 2179
rect 1371 2175 1372 2179
rect 1366 2174 1372 2175
rect 2582 2179 2588 2180
rect 2582 2175 2583 2179
rect 2587 2175 2588 2179
rect 2582 2174 2588 2175
rect 111 2166 115 2167
rect 111 2161 115 2162
rect 159 2166 163 2167
rect 159 2161 163 2162
rect 215 2166 219 2167
rect 215 2161 219 2162
rect 247 2166 251 2167
rect 247 2161 251 2162
rect 311 2166 315 2167
rect 311 2161 315 2162
rect 375 2166 379 2167
rect 375 2161 379 2162
rect 423 2166 427 2167
rect 423 2161 427 2162
rect 511 2166 515 2167
rect 511 2161 515 2162
rect 543 2166 547 2167
rect 543 2161 547 2162
rect 639 2166 643 2167
rect 639 2161 643 2162
rect 663 2166 667 2167
rect 663 2161 667 2162
rect 767 2166 771 2167
rect 767 2161 771 2162
rect 775 2166 779 2167
rect 775 2161 779 2162
rect 879 2166 883 2167
rect 879 2161 883 2162
rect 887 2166 891 2167
rect 887 2161 891 2162
rect 975 2166 979 2167
rect 975 2161 979 2162
rect 999 2166 1003 2167
rect 999 2161 1003 2162
rect 1071 2166 1075 2167
rect 1071 2161 1075 2162
rect 1103 2166 1107 2167
rect 1103 2161 1107 2162
rect 1167 2166 1171 2167
rect 1167 2161 1171 2162
rect 1207 2166 1211 2167
rect 1207 2161 1211 2162
rect 1271 2166 1275 2167
rect 1271 2161 1275 2162
rect 1287 2166 1291 2167
rect 1287 2161 1291 2162
rect 1327 2166 1331 2167
rect 1327 2161 1331 2162
rect 112 2146 114 2161
rect 160 2155 162 2161
rect 216 2155 218 2161
rect 312 2155 314 2161
rect 424 2155 426 2161
rect 544 2155 546 2161
rect 664 2155 666 2161
rect 776 2155 778 2161
rect 880 2155 882 2161
rect 976 2155 978 2161
rect 1072 2155 1074 2161
rect 1168 2155 1170 2161
rect 1272 2155 1274 2161
rect 158 2154 164 2155
rect 158 2150 159 2154
rect 163 2150 164 2154
rect 158 2149 164 2150
rect 214 2154 220 2155
rect 214 2150 215 2154
rect 219 2150 220 2154
rect 214 2149 220 2150
rect 310 2154 316 2155
rect 310 2150 311 2154
rect 315 2150 316 2154
rect 310 2149 316 2150
rect 422 2154 428 2155
rect 422 2150 423 2154
rect 427 2150 428 2154
rect 422 2149 428 2150
rect 542 2154 548 2155
rect 542 2150 543 2154
rect 547 2150 548 2154
rect 542 2149 548 2150
rect 662 2154 668 2155
rect 662 2150 663 2154
rect 667 2150 668 2154
rect 662 2149 668 2150
rect 774 2154 780 2155
rect 774 2150 775 2154
rect 779 2150 780 2154
rect 774 2149 780 2150
rect 878 2154 884 2155
rect 878 2150 879 2154
rect 883 2150 884 2154
rect 878 2149 884 2150
rect 974 2154 980 2155
rect 974 2150 975 2154
rect 979 2150 980 2154
rect 974 2149 980 2150
rect 1070 2154 1076 2155
rect 1070 2150 1071 2154
rect 1075 2150 1076 2154
rect 1070 2149 1076 2150
rect 1166 2154 1172 2155
rect 1166 2150 1167 2154
rect 1171 2150 1172 2154
rect 1166 2149 1172 2150
rect 1270 2154 1276 2155
rect 1270 2150 1271 2154
rect 1275 2150 1276 2154
rect 1270 2149 1276 2150
rect 1328 2146 1330 2161
rect 1368 2159 1370 2174
rect 1470 2170 1476 2171
rect 1470 2166 1471 2170
rect 1475 2166 1476 2170
rect 1470 2165 1476 2166
rect 1550 2170 1556 2171
rect 1550 2166 1551 2170
rect 1555 2166 1556 2170
rect 1550 2165 1556 2166
rect 1646 2170 1652 2171
rect 1646 2166 1647 2170
rect 1651 2166 1652 2170
rect 1646 2165 1652 2166
rect 1758 2170 1764 2171
rect 1758 2166 1759 2170
rect 1763 2166 1764 2170
rect 1758 2165 1764 2166
rect 1878 2170 1884 2171
rect 1878 2166 1879 2170
rect 1883 2166 1884 2170
rect 1878 2165 1884 2166
rect 1998 2170 2004 2171
rect 1998 2166 1999 2170
rect 2003 2166 2004 2170
rect 1998 2165 2004 2166
rect 2110 2170 2116 2171
rect 2110 2166 2111 2170
rect 2115 2166 2116 2170
rect 2110 2165 2116 2166
rect 2222 2170 2228 2171
rect 2222 2166 2223 2170
rect 2227 2166 2228 2170
rect 2222 2165 2228 2166
rect 2326 2170 2332 2171
rect 2326 2166 2327 2170
rect 2331 2166 2332 2170
rect 2326 2165 2332 2166
rect 2438 2170 2444 2171
rect 2438 2166 2439 2170
rect 2443 2166 2444 2170
rect 2438 2165 2444 2166
rect 2542 2170 2548 2171
rect 2542 2166 2543 2170
rect 2547 2166 2548 2170
rect 2542 2165 2548 2166
rect 1472 2159 1474 2165
rect 1552 2159 1554 2165
rect 1648 2159 1650 2165
rect 1760 2159 1762 2165
rect 1880 2159 1882 2165
rect 2000 2159 2002 2165
rect 2112 2159 2114 2165
rect 2224 2159 2226 2165
rect 2328 2159 2330 2165
rect 2440 2159 2442 2165
rect 2544 2159 2546 2165
rect 2584 2159 2586 2174
rect 1367 2158 1371 2159
rect 1367 2153 1371 2154
rect 1471 2158 1475 2159
rect 1471 2153 1475 2154
rect 1535 2158 1539 2159
rect 1535 2153 1539 2154
rect 1551 2158 1555 2159
rect 1551 2153 1555 2154
rect 1631 2158 1635 2159
rect 1631 2153 1635 2154
rect 1647 2158 1651 2159
rect 1647 2153 1651 2154
rect 1735 2158 1739 2159
rect 1735 2153 1739 2154
rect 1759 2158 1763 2159
rect 1759 2153 1763 2154
rect 1839 2158 1843 2159
rect 1839 2153 1843 2154
rect 1879 2158 1883 2159
rect 1879 2153 1883 2154
rect 1951 2158 1955 2159
rect 1951 2153 1955 2154
rect 1999 2158 2003 2159
rect 1999 2153 2003 2154
rect 2055 2158 2059 2159
rect 2055 2153 2059 2154
rect 2111 2158 2115 2159
rect 2111 2153 2115 2154
rect 2159 2158 2163 2159
rect 2159 2153 2163 2154
rect 2223 2158 2227 2159
rect 2223 2153 2227 2154
rect 2263 2158 2267 2159
rect 2263 2153 2267 2154
rect 2327 2158 2331 2159
rect 2327 2153 2331 2154
rect 2359 2158 2363 2159
rect 2359 2153 2363 2154
rect 2439 2158 2443 2159
rect 2439 2153 2443 2154
rect 2463 2158 2467 2159
rect 2463 2153 2467 2154
rect 2543 2158 2547 2159
rect 2543 2153 2547 2154
rect 2583 2158 2587 2159
rect 2583 2153 2587 2154
rect 110 2145 116 2146
rect 110 2141 111 2145
rect 115 2141 116 2145
rect 110 2140 116 2141
rect 1326 2145 1332 2146
rect 1326 2141 1327 2145
rect 1331 2141 1332 2145
rect 1326 2140 1332 2141
rect 1368 2138 1370 2153
rect 1536 2147 1538 2153
rect 1632 2147 1634 2153
rect 1736 2147 1738 2153
rect 1840 2147 1842 2153
rect 1952 2147 1954 2153
rect 2056 2147 2058 2153
rect 2160 2147 2162 2153
rect 2264 2147 2266 2153
rect 2360 2147 2362 2153
rect 2464 2147 2466 2153
rect 2544 2147 2546 2153
rect 1534 2146 1540 2147
rect 1534 2142 1535 2146
rect 1539 2142 1540 2146
rect 1534 2141 1540 2142
rect 1630 2146 1636 2147
rect 1630 2142 1631 2146
rect 1635 2142 1636 2146
rect 1630 2141 1636 2142
rect 1734 2146 1740 2147
rect 1734 2142 1735 2146
rect 1739 2142 1740 2146
rect 1734 2141 1740 2142
rect 1838 2146 1844 2147
rect 1838 2142 1839 2146
rect 1843 2142 1844 2146
rect 1838 2141 1844 2142
rect 1950 2146 1956 2147
rect 1950 2142 1951 2146
rect 1955 2142 1956 2146
rect 1950 2141 1956 2142
rect 2054 2146 2060 2147
rect 2054 2142 2055 2146
rect 2059 2142 2060 2146
rect 2054 2141 2060 2142
rect 2158 2146 2164 2147
rect 2158 2142 2159 2146
rect 2163 2142 2164 2146
rect 2158 2141 2164 2142
rect 2262 2146 2268 2147
rect 2262 2142 2263 2146
rect 2267 2142 2268 2146
rect 2262 2141 2268 2142
rect 2358 2146 2364 2147
rect 2358 2142 2359 2146
rect 2363 2142 2364 2146
rect 2358 2141 2364 2142
rect 2462 2146 2468 2147
rect 2462 2142 2463 2146
rect 2467 2142 2468 2146
rect 2462 2141 2468 2142
rect 2542 2146 2548 2147
rect 2542 2142 2543 2146
rect 2547 2142 2548 2146
rect 2542 2141 2548 2142
rect 2584 2138 2586 2153
rect 1366 2137 1372 2138
rect 1366 2133 1367 2137
rect 1371 2133 1372 2137
rect 1366 2132 1372 2133
rect 2582 2137 2588 2138
rect 2582 2133 2583 2137
rect 2587 2133 2588 2137
rect 2582 2132 2588 2133
rect 110 2128 116 2129
rect 1326 2128 1332 2129
rect 110 2124 111 2128
rect 115 2124 116 2128
rect 110 2123 116 2124
rect 142 2127 148 2128
rect 142 2123 143 2127
rect 147 2123 148 2127
rect 112 2103 114 2123
rect 142 2122 148 2123
rect 198 2127 204 2128
rect 198 2123 199 2127
rect 203 2123 204 2127
rect 198 2122 204 2123
rect 294 2127 300 2128
rect 294 2123 295 2127
rect 299 2123 300 2127
rect 294 2122 300 2123
rect 406 2127 412 2128
rect 406 2123 407 2127
rect 411 2123 412 2127
rect 406 2122 412 2123
rect 526 2127 532 2128
rect 526 2123 527 2127
rect 531 2123 532 2127
rect 526 2122 532 2123
rect 646 2127 652 2128
rect 646 2123 647 2127
rect 651 2123 652 2127
rect 646 2122 652 2123
rect 758 2127 764 2128
rect 758 2123 759 2127
rect 763 2123 764 2127
rect 758 2122 764 2123
rect 862 2127 868 2128
rect 862 2123 863 2127
rect 867 2123 868 2127
rect 862 2122 868 2123
rect 958 2127 964 2128
rect 958 2123 959 2127
rect 963 2123 964 2127
rect 958 2122 964 2123
rect 1054 2127 1060 2128
rect 1054 2123 1055 2127
rect 1059 2123 1060 2127
rect 1054 2122 1060 2123
rect 1150 2127 1156 2128
rect 1150 2123 1151 2127
rect 1155 2123 1156 2127
rect 1150 2122 1156 2123
rect 1254 2127 1260 2128
rect 1254 2123 1255 2127
rect 1259 2123 1260 2127
rect 1326 2124 1327 2128
rect 1331 2124 1332 2128
rect 1326 2123 1332 2124
rect 1254 2122 1260 2123
rect 144 2103 146 2122
rect 200 2103 202 2122
rect 296 2103 298 2122
rect 408 2103 410 2122
rect 528 2103 530 2122
rect 648 2103 650 2122
rect 760 2103 762 2122
rect 864 2103 866 2122
rect 960 2103 962 2122
rect 1056 2103 1058 2122
rect 1152 2103 1154 2122
rect 1256 2103 1258 2122
rect 1328 2103 1330 2123
rect 1366 2120 1372 2121
rect 2582 2120 2588 2121
rect 1366 2116 1367 2120
rect 1371 2116 1372 2120
rect 1366 2115 1372 2116
rect 1518 2119 1524 2120
rect 1518 2115 1519 2119
rect 1523 2115 1524 2119
rect 1368 2103 1370 2115
rect 1518 2114 1524 2115
rect 1614 2119 1620 2120
rect 1614 2115 1615 2119
rect 1619 2115 1620 2119
rect 1614 2114 1620 2115
rect 1718 2119 1724 2120
rect 1718 2115 1719 2119
rect 1723 2115 1724 2119
rect 1718 2114 1724 2115
rect 1822 2119 1828 2120
rect 1822 2115 1823 2119
rect 1827 2115 1828 2119
rect 1822 2114 1828 2115
rect 1934 2119 1940 2120
rect 1934 2115 1935 2119
rect 1939 2115 1940 2119
rect 1934 2114 1940 2115
rect 2038 2119 2044 2120
rect 2038 2115 2039 2119
rect 2043 2115 2044 2119
rect 2038 2114 2044 2115
rect 2142 2119 2148 2120
rect 2142 2115 2143 2119
rect 2147 2115 2148 2119
rect 2142 2114 2148 2115
rect 2246 2119 2252 2120
rect 2246 2115 2247 2119
rect 2251 2115 2252 2119
rect 2246 2114 2252 2115
rect 2342 2119 2348 2120
rect 2342 2115 2343 2119
rect 2347 2115 2348 2119
rect 2342 2114 2348 2115
rect 2446 2119 2452 2120
rect 2446 2115 2447 2119
rect 2451 2115 2452 2119
rect 2446 2114 2452 2115
rect 2526 2119 2532 2120
rect 2526 2115 2527 2119
rect 2531 2115 2532 2119
rect 2582 2116 2583 2120
rect 2587 2116 2588 2120
rect 2582 2115 2588 2116
rect 2526 2114 2532 2115
rect 1520 2103 1522 2114
rect 1616 2103 1618 2114
rect 1720 2103 1722 2114
rect 1824 2103 1826 2114
rect 1936 2103 1938 2114
rect 2040 2103 2042 2114
rect 2144 2103 2146 2114
rect 2248 2103 2250 2114
rect 2344 2103 2346 2114
rect 2448 2103 2450 2114
rect 2528 2103 2530 2114
rect 2584 2103 2586 2115
rect 111 2102 115 2103
rect 111 2097 115 2098
rect 143 2102 147 2103
rect 143 2097 147 2098
rect 199 2102 203 2103
rect 199 2097 203 2098
rect 263 2102 267 2103
rect 263 2097 267 2098
rect 295 2102 299 2103
rect 295 2097 299 2098
rect 327 2102 331 2103
rect 327 2097 331 2098
rect 399 2102 403 2103
rect 399 2097 403 2098
rect 407 2102 411 2103
rect 407 2097 411 2098
rect 479 2102 483 2103
rect 479 2097 483 2098
rect 527 2102 531 2103
rect 527 2097 531 2098
rect 567 2102 571 2103
rect 567 2097 571 2098
rect 647 2102 651 2103
rect 647 2097 651 2098
rect 655 2102 659 2103
rect 655 2097 659 2098
rect 735 2102 739 2103
rect 735 2097 739 2098
rect 759 2102 763 2103
rect 759 2097 763 2098
rect 815 2102 819 2103
rect 815 2097 819 2098
rect 863 2102 867 2103
rect 863 2097 867 2098
rect 887 2102 891 2103
rect 887 2097 891 2098
rect 959 2102 963 2103
rect 959 2097 963 2098
rect 967 2102 971 2103
rect 967 2097 971 2098
rect 1047 2102 1051 2103
rect 1047 2097 1051 2098
rect 1055 2102 1059 2103
rect 1055 2097 1059 2098
rect 1127 2102 1131 2103
rect 1127 2097 1131 2098
rect 1151 2102 1155 2103
rect 1151 2097 1155 2098
rect 1255 2102 1259 2103
rect 1255 2097 1259 2098
rect 1327 2102 1331 2103
rect 1327 2097 1331 2098
rect 1367 2102 1371 2103
rect 1367 2097 1371 2098
rect 1431 2102 1435 2103
rect 1431 2097 1435 2098
rect 1519 2102 1523 2103
rect 1519 2097 1523 2098
rect 1535 2102 1539 2103
rect 1535 2097 1539 2098
rect 1615 2102 1619 2103
rect 1615 2097 1619 2098
rect 1647 2102 1651 2103
rect 1647 2097 1651 2098
rect 1719 2102 1723 2103
rect 1719 2097 1723 2098
rect 1759 2102 1763 2103
rect 1759 2097 1763 2098
rect 1823 2102 1827 2103
rect 1823 2097 1827 2098
rect 1863 2102 1867 2103
rect 1863 2097 1867 2098
rect 1935 2102 1939 2103
rect 1935 2097 1939 2098
rect 1967 2102 1971 2103
rect 1967 2097 1971 2098
rect 2039 2102 2043 2103
rect 2039 2097 2043 2098
rect 2071 2102 2075 2103
rect 2071 2097 2075 2098
rect 2143 2102 2147 2103
rect 2143 2097 2147 2098
rect 2175 2102 2179 2103
rect 2175 2097 2179 2098
rect 2247 2102 2251 2103
rect 2247 2097 2251 2098
rect 2271 2102 2275 2103
rect 2271 2097 2275 2098
rect 2343 2102 2347 2103
rect 2343 2097 2347 2098
rect 2359 2102 2363 2103
rect 2359 2097 2363 2098
rect 2447 2102 2451 2103
rect 2447 2097 2451 2098
rect 2455 2102 2459 2103
rect 2455 2097 2459 2098
rect 2527 2102 2531 2103
rect 2527 2097 2531 2098
rect 2583 2102 2587 2103
rect 2583 2097 2587 2098
rect 112 2085 114 2097
rect 264 2086 266 2097
rect 328 2086 330 2097
rect 400 2086 402 2097
rect 480 2086 482 2097
rect 568 2086 570 2097
rect 656 2086 658 2097
rect 736 2086 738 2097
rect 816 2086 818 2097
rect 888 2086 890 2097
rect 968 2086 970 2097
rect 1048 2086 1050 2097
rect 1128 2086 1130 2097
rect 262 2085 268 2086
rect 110 2084 116 2085
rect 110 2080 111 2084
rect 115 2080 116 2084
rect 262 2081 263 2085
rect 267 2081 268 2085
rect 262 2080 268 2081
rect 326 2085 332 2086
rect 326 2081 327 2085
rect 331 2081 332 2085
rect 326 2080 332 2081
rect 398 2085 404 2086
rect 398 2081 399 2085
rect 403 2081 404 2085
rect 398 2080 404 2081
rect 478 2085 484 2086
rect 478 2081 479 2085
rect 483 2081 484 2085
rect 478 2080 484 2081
rect 566 2085 572 2086
rect 566 2081 567 2085
rect 571 2081 572 2085
rect 566 2080 572 2081
rect 654 2085 660 2086
rect 654 2081 655 2085
rect 659 2081 660 2085
rect 654 2080 660 2081
rect 734 2085 740 2086
rect 734 2081 735 2085
rect 739 2081 740 2085
rect 734 2080 740 2081
rect 814 2085 820 2086
rect 814 2081 815 2085
rect 819 2081 820 2085
rect 814 2080 820 2081
rect 886 2085 892 2086
rect 886 2081 887 2085
rect 891 2081 892 2085
rect 886 2080 892 2081
rect 966 2085 972 2086
rect 966 2081 967 2085
rect 971 2081 972 2085
rect 966 2080 972 2081
rect 1046 2085 1052 2086
rect 1046 2081 1047 2085
rect 1051 2081 1052 2085
rect 1046 2080 1052 2081
rect 1126 2085 1132 2086
rect 1328 2085 1330 2097
rect 1368 2085 1370 2097
rect 1432 2086 1434 2097
rect 1536 2086 1538 2097
rect 1648 2086 1650 2097
rect 1760 2086 1762 2097
rect 1864 2086 1866 2097
rect 1968 2086 1970 2097
rect 2072 2086 2074 2097
rect 2176 2086 2178 2097
rect 2272 2086 2274 2097
rect 2360 2086 2362 2097
rect 2456 2086 2458 2097
rect 2528 2086 2530 2097
rect 1430 2085 1436 2086
rect 1126 2081 1127 2085
rect 1131 2081 1132 2085
rect 1126 2080 1132 2081
rect 1326 2084 1332 2085
rect 1326 2080 1327 2084
rect 1331 2080 1332 2084
rect 110 2079 116 2080
rect 1326 2079 1332 2080
rect 1366 2084 1372 2085
rect 1366 2080 1367 2084
rect 1371 2080 1372 2084
rect 1430 2081 1431 2085
rect 1435 2081 1436 2085
rect 1430 2080 1436 2081
rect 1534 2085 1540 2086
rect 1534 2081 1535 2085
rect 1539 2081 1540 2085
rect 1534 2080 1540 2081
rect 1646 2085 1652 2086
rect 1646 2081 1647 2085
rect 1651 2081 1652 2085
rect 1646 2080 1652 2081
rect 1758 2085 1764 2086
rect 1758 2081 1759 2085
rect 1763 2081 1764 2085
rect 1758 2080 1764 2081
rect 1862 2085 1868 2086
rect 1862 2081 1863 2085
rect 1867 2081 1868 2085
rect 1862 2080 1868 2081
rect 1966 2085 1972 2086
rect 1966 2081 1967 2085
rect 1971 2081 1972 2085
rect 1966 2080 1972 2081
rect 2070 2085 2076 2086
rect 2070 2081 2071 2085
rect 2075 2081 2076 2085
rect 2070 2080 2076 2081
rect 2174 2085 2180 2086
rect 2174 2081 2175 2085
rect 2179 2081 2180 2085
rect 2174 2080 2180 2081
rect 2270 2085 2276 2086
rect 2270 2081 2271 2085
rect 2275 2081 2276 2085
rect 2270 2080 2276 2081
rect 2358 2085 2364 2086
rect 2358 2081 2359 2085
rect 2363 2081 2364 2085
rect 2358 2080 2364 2081
rect 2454 2085 2460 2086
rect 2454 2081 2455 2085
rect 2459 2081 2460 2085
rect 2454 2080 2460 2081
rect 2526 2085 2532 2086
rect 2584 2085 2586 2097
rect 2526 2081 2527 2085
rect 2531 2081 2532 2085
rect 2526 2080 2532 2081
rect 2582 2084 2588 2085
rect 2582 2080 2583 2084
rect 2587 2080 2588 2084
rect 1366 2079 1372 2080
rect 2582 2079 2588 2080
rect 110 2067 116 2068
rect 110 2063 111 2067
rect 115 2063 116 2067
rect 110 2062 116 2063
rect 1326 2067 1332 2068
rect 1326 2063 1327 2067
rect 1331 2063 1332 2067
rect 1326 2062 1332 2063
rect 1366 2067 1372 2068
rect 1366 2063 1367 2067
rect 1371 2063 1372 2067
rect 1366 2062 1372 2063
rect 2582 2067 2588 2068
rect 2582 2063 2583 2067
rect 2587 2063 2588 2067
rect 2582 2062 2588 2063
rect 112 2039 114 2062
rect 278 2058 284 2059
rect 278 2054 279 2058
rect 283 2054 284 2058
rect 278 2053 284 2054
rect 342 2058 348 2059
rect 342 2054 343 2058
rect 347 2054 348 2058
rect 342 2053 348 2054
rect 414 2058 420 2059
rect 414 2054 415 2058
rect 419 2054 420 2058
rect 414 2053 420 2054
rect 494 2058 500 2059
rect 494 2054 495 2058
rect 499 2054 500 2058
rect 494 2053 500 2054
rect 582 2058 588 2059
rect 582 2054 583 2058
rect 587 2054 588 2058
rect 582 2053 588 2054
rect 670 2058 676 2059
rect 670 2054 671 2058
rect 675 2054 676 2058
rect 670 2053 676 2054
rect 750 2058 756 2059
rect 750 2054 751 2058
rect 755 2054 756 2058
rect 750 2053 756 2054
rect 830 2058 836 2059
rect 830 2054 831 2058
rect 835 2054 836 2058
rect 830 2053 836 2054
rect 902 2058 908 2059
rect 902 2054 903 2058
rect 907 2054 908 2058
rect 902 2053 908 2054
rect 982 2058 988 2059
rect 982 2054 983 2058
rect 987 2054 988 2058
rect 982 2053 988 2054
rect 1062 2058 1068 2059
rect 1062 2054 1063 2058
rect 1067 2054 1068 2058
rect 1062 2053 1068 2054
rect 1142 2058 1148 2059
rect 1142 2054 1143 2058
rect 1147 2054 1148 2058
rect 1142 2053 1148 2054
rect 280 2039 282 2053
rect 344 2039 346 2053
rect 416 2039 418 2053
rect 496 2039 498 2053
rect 584 2039 586 2053
rect 672 2039 674 2053
rect 752 2039 754 2053
rect 832 2039 834 2053
rect 904 2039 906 2053
rect 984 2039 986 2053
rect 1064 2039 1066 2053
rect 1144 2039 1146 2053
rect 1328 2039 1330 2062
rect 1368 2047 1370 2062
rect 1446 2058 1452 2059
rect 1446 2054 1447 2058
rect 1451 2054 1452 2058
rect 1446 2053 1452 2054
rect 1550 2058 1556 2059
rect 1550 2054 1551 2058
rect 1555 2054 1556 2058
rect 1550 2053 1556 2054
rect 1662 2058 1668 2059
rect 1662 2054 1663 2058
rect 1667 2054 1668 2058
rect 1662 2053 1668 2054
rect 1774 2058 1780 2059
rect 1774 2054 1775 2058
rect 1779 2054 1780 2058
rect 1774 2053 1780 2054
rect 1878 2058 1884 2059
rect 1878 2054 1879 2058
rect 1883 2054 1884 2058
rect 1878 2053 1884 2054
rect 1982 2058 1988 2059
rect 1982 2054 1983 2058
rect 1987 2054 1988 2058
rect 1982 2053 1988 2054
rect 2086 2058 2092 2059
rect 2086 2054 2087 2058
rect 2091 2054 2092 2058
rect 2086 2053 2092 2054
rect 2190 2058 2196 2059
rect 2190 2054 2191 2058
rect 2195 2054 2196 2058
rect 2190 2053 2196 2054
rect 2286 2058 2292 2059
rect 2286 2054 2287 2058
rect 2291 2054 2292 2058
rect 2286 2053 2292 2054
rect 2374 2058 2380 2059
rect 2374 2054 2375 2058
rect 2379 2054 2380 2058
rect 2374 2053 2380 2054
rect 2470 2058 2476 2059
rect 2470 2054 2471 2058
rect 2475 2054 2476 2058
rect 2470 2053 2476 2054
rect 2542 2058 2548 2059
rect 2542 2054 2543 2058
rect 2547 2054 2548 2058
rect 2542 2053 2548 2054
rect 1448 2047 1450 2053
rect 1552 2047 1554 2053
rect 1664 2047 1666 2053
rect 1776 2047 1778 2053
rect 1880 2047 1882 2053
rect 1984 2047 1986 2053
rect 2088 2047 2090 2053
rect 2192 2047 2194 2053
rect 2288 2047 2290 2053
rect 2376 2047 2378 2053
rect 2472 2047 2474 2053
rect 2544 2047 2546 2053
rect 2584 2047 2586 2062
rect 1367 2046 1371 2047
rect 1367 2041 1371 2042
rect 1415 2046 1419 2047
rect 1415 2041 1419 2042
rect 1447 2046 1451 2047
rect 1447 2041 1451 2042
rect 1503 2046 1507 2047
rect 1503 2041 1507 2042
rect 1551 2046 1555 2047
rect 1551 2041 1555 2042
rect 1607 2046 1611 2047
rect 1607 2041 1611 2042
rect 1663 2046 1667 2047
rect 1663 2041 1667 2042
rect 1711 2046 1715 2047
rect 1711 2041 1715 2042
rect 1775 2046 1779 2047
rect 1775 2041 1779 2042
rect 1807 2046 1811 2047
rect 1807 2041 1811 2042
rect 1879 2046 1883 2047
rect 1879 2041 1883 2042
rect 1903 2046 1907 2047
rect 1903 2041 1907 2042
rect 1983 2046 1987 2047
rect 1983 2041 1987 2042
rect 2007 2046 2011 2047
rect 2007 2041 2011 2042
rect 2087 2046 2091 2047
rect 2087 2041 2091 2042
rect 2111 2046 2115 2047
rect 2111 2041 2115 2042
rect 2191 2046 2195 2047
rect 2191 2041 2195 2042
rect 2215 2046 2219 2047
rect 2215 2041 2219 2042
rect 2287 2046 2291 2047
rect 2287 2041 2291 2042
rect 2327 2046 2331 2047
rect 2327 2041 2331 2042
rect 2375 2046 2379 2047
rect 2375 2041 2379 2042
rect 2447 2046 2451 2047
rect 2447 2041 2451 2042
rect 2471 2046 2475 2047
rect 2471 2041 2475 2042
rect 2543 2046 2547 2047
rect 2543 2041 2547 2042
rect 2583 2046 2587 2047
rect 2583 2041 2587 2042
rect 111 2038 115 2039
rect 111 2033 115 2034
rect 279 2038 283 2039
rect 279 2033 283 2034
rect 343 2038 347 2039
rect 343 2033 347 2034
rect 415 2038 419 2039
rect 415 2033 419 2034
rect 471 2038 475 2039
rect 471 2033 475 2034
rect 495 2038 499 2039
rect 495 2033 499 2034
rect 527 2038 531 2039
rect 527 2033 531 2034
rect 583 2038 587 2039
rect 583 2033 587 2034
rect 639 2038 643 2039
rect 639 2033 643 2034
rect 671 2038 675 2039
rect 671 2033 675 2034
rect 695 2038 699 2039
rect 695 2033 699 2034
rect 751 2038 755 2039
rect 751 2033 755 2034
rect 807 2038 811 2039
rect 807 2033 811 2034
rect 831 2038 835 2039
rect 831 2033 835 2034
rect 863 2038 867 2039
rect 863 2033 867 2034
rect 903 2038 907 2039
rect 903 2033 907 2034
rect 919 2038 923 2039
rect 919 2033 923 2034
rect 975 2038 979 2039
rect 975 2033 979 2034
rect 983 2038 987 2039
rect 983 2033 987 2034
rect 1031 2038 1035 2039
rect 1031 2033 1035 2034
rect 1063 2038 1067 2039
rect 1063 2033 1067 2034
rect 1143 2038 1147 2039
rect 1143 2033 1147 2034
rect 1327 2038 1331 2039
rect 1327 2033 1331 2034
rect 112 2018 114 2033
rect 416 2027 418 2033
rect 472 2027 474 2033
rect 528 2027 530 2033
rect 584 2027 586 2033
rect 640 2027 642 2033
rect 696 2027 698 2033
rect 752 2027 754 2033
rect 808 2027 810 2033
rect 864 2027 866 2033
rect 920 2027 922 2033
rect 976 2027 978 2033
rect 1032 2027 1034 2033
rect 414 2026 420 2027
rect 414 2022 415 2026
rect 419 2022 420 2026
rect 414 2021 420 2022
rect 470 2026 476 2027
rect 470 2022 471 2026
rect 475 2022 476 2026
rect 470 2021 476 2022
rect 526 2026 532 2027
rect 526 2022 527 2026
rect 531 2022 532 2026
rect 526 2021 532 2022
rect 582 2026 588 2027
rect 582 2022 583 2026
rect 587 2022 588 2026
rect 582 2021 588 2022
rect 638 2026 644 2027
rect 638 2022 639 2026
rect 643 2022 644 2026
rect 638 2021 644 2022
rect 694 2026 700 2027
rect 694 2022 695 2026
rect 699 2022 700 2026
rect 694 2021 700 2022
rect 750 2026 756 2027
rect 750 2022 751 2026
rect 755 2022 756 2026
rect 750 2021 756 2022
rect 806 2026 812 2027
rect 806 2022 807 2026
rect 811 2022 812 2026
rect 806 2021 812 2022
rect 862 2026 868 2027
rect 862 2022 863 2026
rect 867 2022 868 2026
rect 862 2021 868 2022
rect 918 2026 924 2027
rect 918 2022 919 2026
rect 923 2022 924 2026
rect 918 2021 924 2022
rect 974 2026 980 2027
rect 974 2022 975 2026
rect 979 2022 980 2026
rect 974 2021 980 2022
rect 1030 2026 1036 2027
rect 1030 2022 1031 2026
rect 1035 2022 1036 2026
rect 1030 2021 1036 2022
rect 1328 2018 1330 2033
rect 1368 2026 1370 2041
rect 1416 2035 1418 2041
rect 1504 2035 1506 2041
rect 1608 2035 1610 2041
rect 1712 2035 1714 2041
rect 1808 2035 1810 2041
rect 1904 2035 1906 2041
rect 2008 2035 2010 2041
rect 2112 2035 2114 2041
rect 2216 2035 2218 2041
rect 2328 2035 2330 2041
rect 2448 2035 2450 2041
rect 2544 2035 2546 2041
rect 1414 2034 1420 2035
rect 1414 2030 1415 2034
rect 1419 2030 1420 2034
rect 1414 2029 1420 2030
rect 1502 2034 1508 2035
rect 1502 2030 1503 2034
rect 1507 2030 1508 2034
rect 1502 2029 1508 2030
rect 1606 2034 1612 2035
rect 1606 2030 1607 2034
rect 1611 2030 1612 2034
rect 1606 2029 1612 2030
rect 1710 2034 1716 2035
rect 1710 2030 1711 2034
rect 1715 2030 1716 2034
rect 1710 2029 1716 2030
rect 1806 2034 1812 2035
rect 1806 2030 1807 2034
rect 1811 2030 1812 2034
rect 1806 2029 1812 2030
rect 1902 2034 1908 2035
rect 1902 2030 1903 2034
rect 1907 2030 1908 2034
rect 1902 2029 1908 2030
rect 2006 2034 2012 2035
rect 2006 2030 2007 2034
rect 2011 2030 2012 2034
rect 2006 2029 2012 2030
rect 2110 2034 2116 2035
rect 2110 2030 2111 2034
rect 2115 2030 2116 2034
rect 2110 2029 2116 2030
rect 2214 2034 2220 2035
rect 2214 2030 2215 2034
rect 2219 2030 2220 2034
rect 2214 2029 2220 2030
rect 2326 2034 2332 2035
rect 2326 2030 2327 2034
rect 2331 2030 2332 2034
rect 2326 2029 2332 2030
rect 2446 2034 2452 2035
rect 2446 2030 2447 2034
rect 2451 2030 2452 2034
rect 2446 2029 2452 2030
rect 2542 2034 2548 2035
rect 2542 2030 2543 2034
rect 2547 2030 2548 2034
rect 2542 2029 2548 2030
rect 2584 2026 2586 2041
rect 1366 2025 1372 2026
rect 1366 2021 1367 2025
rect 1371 2021 1372 2025
rect 1366 2020 1372 2021
rect 2582 2025 2588 2026
rect 2582 2021 2583 2025
rect 2587 2021 2588 2025
rect 2582 2020 2588 2021
rect 110 2017 116 2018
rect 110 2013 111 2017
rect 115 2013 116 2017
rect 110 2012 116 2013
rect 1326 2017 1332 2018
rect 1326 2013 1327 2017
rect 1331 2013 1332 2017
rect 1326 2012 1332 2013
rect 1366 2008 1372 2009
rect 2582 2008 2588 2009
rect 1366 2004 1367 2008
rect 1371 2004 1372 2008
rect 1366 2003 1372 2004
rect 1398 2007 1404 2008
rect 1398 2003 1399 2007
rect 1403 2003 1404 2007
rect 110 2000 116 2001
rect 1326 2000 1332 2001
rect 110 1996 111 2000
rect 115 1996 116 2000
rect 110 1995 116 1996
rect 398 1999 404 2000
rect 398 1995 399 1999
rect 403 1995 404 1999
rect 112 1979 114 1995
rect 398 1994 404 1995
rect 454 1999 460 2000
rect 454 1995 455 1999
rect 459 1995 460 1999
rect 454 1994 460 1995
rect 510 1999 516 2000
rect 510 1995 511 1999
rect 515 1995 516 1999
rect 510 1994 516 1995
rect 566 1999 572 2000
rect 566 1995 567 1999
rect 571 1995 572 1999
rect 566 1994 572 1995
rect 622 1999 628 2000
rect 622 1995 623 1999
rect 627 1995 628 1999
rect 622 1994 628 1995
rect 678 1999 684 2000
rect 678 1995 679 1999
rect 683 1995 684 1999
rect 678 1994 684 1995
rect 734 1999 740 2000
rect 734 1995 735 1999
rect 739 1995 740 1999
rect 734 1994 740 1995
rect 790 1999 796 2000
rect 790 1995 791 1999
rect 795 1995 796 1999
rect 790 1994 796 1995
rect 846 1999 852 2000
rect 846 1995 847 1999
rect 851 1995 852 1999
rect 846 1994 852 1995
rect 902 1999 908 2000
rect 902 1995 903 1999
rect 907 1995 908 1999
rect 902 1994 908 1995
rect 958 1999 964 2000
rect 958 1995 959 1999
rect 963 1995 964 1999
rect 958 1994 964 1995
rect 1014 1999 1020 2000
rect 1014 1995 1015 1999
rect 1019 1995 1020 1999
rect 1326 1996 1327 2000
rect 1331 1996 1332 2000
rect 1326 1995 1332 1996
rect 1014 1994 1020 1995
rect 400 1979 402 1994
rect 456 1979 458 1994
rect 512 1979 514 1994
rect 568 1979 570 1994
rect 624 1979 626 1994
rect 680 1979 682 1994
rect 736 1979 738 1994
rect 792 1979 794 1994
rect 848 1979 850 1994
rect 904 1979 906 1994
rect 960 1979 962 1994
rect 1016 1979 1018 1994
rect 1328 1979 1330 1995
rect 1368 1991 1370 2003
rect 1398 2002 1404 2003
rect 1486 2007 1492 2008
rect 1486 2003 1487 2007
rect 1491 2003 1492 2007
rect 1486 2002 1492 2003
rect 1590 2007 1596 2008
rect 1590 2003 1591 2007
rect 1595 2003 1596 2007
rect 1590 2002 1596 2003
rect 1694 2007 1700 2008
rect 1694 2003 1695 2007
rect 1699 2003 1700 2007
rect 1694 2002 1700 2003
rect 1790 2007 1796 2008
rect 1790 2003 1791 2007
rect 1795 2003 1796 2007
rect 1790 2002 1796 2003
rect 1886 2007 1892 2008
rect 1886 2003 1887 2007
rect 1891 2003 1892 2007
rect 1886 2002 1892 2003
rect 1990 2007 1996 2008
rect 1990 2003 1991 2007
rect 1995 2003 1996 2007
rect 1990 2002 1996 2003
rect 2094 2007 2100 2008
rect 2094 2003 2095 2007
rect 2099 2003 2100 2007
rect 2094 2002 2100 2003
rect 2198 2007 2204 2008
rect 2198 2003 2199 2007
rect 2203 2003 2204 2007
rect 2198 2002 2204 2003
rect 2310 2007 2316 2008
rect 2310 2003 2311 2007
rect 2315 2003 2316 2007
rect 2310 2002 2316 2003
rect 2430 2007 2436 2008
rect 2430 2003 2431 2007
rect 2435 2003 2436 2007
rect 2430 2002 2436 2003
rect 2526 2007 2532 2008
rect 2526 2003 2527 2007
rect 2531 2003 2532 2007
rect 2582 2004 2583 2008
rect 2587 2004 2588 2008
rect 2582 2003 2588 2004
rect 2526 2002 2532 2003
rect 1400 1991 1402 2002
rect 1488 1991 1490 2002
rect 1592 1991 1594 2002
rect 1696 1991 1698 2002
rect 1792 1991 1794 2002
rect 1888 1991 1890 2002
rect 1992 1991 1994 2002
rect 2096 1991 2098 2002
rect 2200 1991 2202 2002
rect 2312 1991 2314 2002
rect 2432 1991 2434 2002
rect 2528 1991 2530 2002
rect 2584 1991 2586 2003
rect 1367 1990 1371 1991
rect 1367 1985 1371 1986
rect 1399 1990 1403 1991
rect 1399 1985 1403 1986
rect 1479 1990 1483 1991
rect 1479 1985 1483 1986
rect 1487 1990 1491 1991
rect 1487 1985 1491 1986
rect 1583 1990 1587 1991
rect 1583 1985 1587 1986
rect 1591 1990 1595 1991
rect 1591 1985 1595 1986
rect 1679 1990 1683 1991
rect 1679 1985 1683 1986
rect 1695 1990 1699 1991
rect 1695 1985 1699 1986
rect 1767 1990 1771 1991
rect 1767 1985 1771 1986
rect 1791 1990 1795 1991
rect 1791 1985 1795 1986
rect 1847 1990 1851 1991
rect 1847 1985 1851 1986
rect 1887 1990 1891 1991
rect 1887 1985 1891 1986
rect 1927 1990 1931 1991
rect 1927 1985 1931 1986
rect 1991 1990 1995 1991
rect 1991 1985 1995 1986
rect 2007 1990 2011 1991
rect 2007 1985 2011 1986
rect 2087 1990 2091 1991
rect 2087 1985 2091 1986
rect 2095 1990 2099 1991
rect 2095 1985 2099 1986
rect 2199 1990 2203 1991
rect 2199 1985 2203 1986
rect 2311 1990 2315 1991
rect 2311 1985 2315 1986
rect 2431 1990 2435 1991
rect 2431 1985 2435 1986
rect 2527 1990 2531 1991
rect 2527 1985 2531 1986
rect 2583 1990 2587 1991
rect 2583 1985 2587 1986
rect 111 1978 115 1979
rect 111 1973 115 1974
rect 335 1978 339 1979
rect 335 1973 339 1974
rect 391 1978 395 1979
rect 391 1973 395 1974
rect 399 1978 403 1979
rect 399 1973 403 1974
rect 447 1978 451 1979
rect 447 1973 451 1974
rect 455 1978 459 1979
rect 455 1973 459 1974
rect 503 1978 507 1979
rect 503 1973 507 1974
rect 511 1978 515 1979
rect 511 1973 515 1974
rect 567 1978 571 1979
rect 567 1973 571 1974
rect 623 1978 627 1979
rect 623 1973 627 1974
rect 647 1978 651 1979
rect 647 1973 651 1974
rect 679 1978 683 1979
rect 679 1973 683 1974
rect 735 1978 739 1979
rect 735 1973 739 1974
rect 743 1978 747 1979
rect 743 1973 747 1974
rect 791 1978 795 1979
rect 791 1973 795 1974
rect 847 1978 851 1979
rect 847 1973 851 1974
rect 863 1978 867 1979
rect 863 1973 867 1974
rect 903 1978 907 1979
rect 903 1973 907 1974
rect 959 1978 963 1979
rect 959 1973 963 1974
rect 999 1978 1003 1979
rect 999 1973 1003 1974
rect 1015 1978 1019 1979
rect 1015 1973 1019 1974
rect 1143 1978 1147 1979
rect 1143 1973 1147 1974
rect 1271 1978 1275 1979
rect 1271 1973 1275 1974
rect 1327 1978 1331 1979
rect 1327 1973 1331 1974
rect 1368 1973 1370 1985
rect 1400 1974 1402 1985
rect 1480 1974 1482 1985
rect 1584 1974 1586 1985
rect 1680 1974 1682 1985
rect 1768 1974 1770 1985
rect 1848 1974 1850 1985
rect 1928 1974 1930 1985
rect 2008 1974 2010 1985
rect 2088 1974 2090 1985
rect 1398 1973 1404 1974
rect 112 1961 114 1973
rect 336 1962 338 1973
rect 392 1962 394 1973
rect 448 1962 450 1973
rect 504 1962 506 1973
rect 568 1962 570 1973
rect 648 1962 650 1973
rect 744 1962 746 1973
rect 864 1962 866 1973
rect 1000 1962 1002 1973
rect 1144 1962 1146 1973
rect 1272 1962 1274 1973
rect 334 1961 340 1962
rect 110 1960 116 1961
rect 110 1956 111 1960
rect 115 1956 116 1960
rect 334 1957 335 1961
rect 339 1957 340 1961
rect 334 1956 340 1957
rect 390 1961 396 1962
rect 390 1957 391 1961
rect 395 1957 396 1961
rect 390 1956 396 1957
rect 446 1961 452 1962
rect 446 1957 447 1961
rect 451 1957 452 1961
rect 446 1956 452 1957
rect 502 1961 508 1962
rect 502 1957 503 1961
rect 507 1957 508 1961
rect 502 1956 508 1957
rect 566 1961 572 1962
rect 566 1957 567 1961
rect 571 1957 572 1961
rect 566 1956 572 1957
rect 646 1961 652 1962
rect 646 1957 647 1961
rect 651 1957 652 1961
rect 646 1956 652 1957
rect 742 1961 748 1962
rect 742 1957 743 1961
rect 747 1957 748 1961
rect 742 1956 748 1957
rect 862 1961 868 1962
rect 862 1957 863 1961
rect 867 1957 868 1961
rect 862 1956 868 1957
rect 998 1961 1004 1962
rect 998 1957 999 1961
rect 1003 1957 1004 1961
rect 998 1956 1004 1957
rect 1142 1961 1148 1962
rect 1142 1957 1143 1961
rect 1147 1957 1148 1961
rect 1142 1956 1148 1957
rect 1270 1961 1276 1962
rect 1328 1961 1330 1973
rect 1366 1972 1372 1973
rect 1366 1968 1367 1972
rect 1371 1968 1372 1972
rect 1398 1969 1399 1973
rect 1403 1969 1404 1973
rect 1398 1968 1404 1969
rect 1478 1973 1484 1974
rect 1478 1969 1479 1973
rect 1483 1969 1484 1973
rect 1478 1968 1484 1969
rect 1582 1973 1588 1974
rect 1582 1969 1583 1973
rect 1587 1969 1588 1973
rect 1582 1968 1588 1969
rect 1678 1973 1684 1974
rect 1678 1969 1679 1973
rect 1683 1969 1684 1973
rect 1678 1968 1684 1969
rect 1766 1973 1772 1974
rect 1766 1969 1767 1973
rect 1771 1969 1772 1973
rect 1766 1968 1772 1969
rect 1846 1973 1852 1974
rect 1846 1969 1847 1973
rect 1851 1969 1852 1973
rect 1846 1968 1852 1969
rect 1926 1973 1932 1974
rect 1926 1969 1927 1973
rect 1931 1969 1932 1973
rect 1926 1968 1932 1969
rect 2006 1973 2012 1974
rect 2006 1969 2007 1973
rect 2011 1969 2012 1973
rect 2006 1968 2012 1969
rect 2086 1973 2092 1974
rect 2584 1973 2586 1985
rect 2086 1969 2087 1973
rect 2091 1969 2092 1973
rect 2086 1968 2092 1969
rect 2582 1972 2588 1973
rect 2582 1968 2583 1972
rect 2587 1968 2588 1972
rect 1366 1967 1372 1968
rect 2582 1967 2588 1968
rect 1270 1957 1271 1961
rect 1275 1957 1276 1961
rect 1270 1956 1276 1957
rect 1326 1960 1332 1961
rect 1326 1956 1327 1960
rect 1331 1956 1332 1960
rect 110 1955 116 1956
rect 1326 1955 1332 1956
rect 1366 1955 1372 1956
rect 1366 1951 1367 1955
rect 1371 1951 1372 1955
rect 1366 1950 1372 1951
rect 2582 1955 2588 1956
rect 2582 1951 2583 1955
rect 2587 1951 2588 1955
rect 2582 1950 2588 1951
rect 110 1943 116 1944
rect 110 1939 111 1943
rect 115 1939 116 1943
rect 110 1938 116 1939
rect 1326 1943 1332 1944
rect 1326 1939 1327 1943
rect 1331 1939 1332 1943
rect 1326 1938 1332 1939
rect 112 1923 114 1938
rect 350 1934 356 1935
rect 350 1930 351 1934
rect 355 1930 356 1934
rect 350 1929 356 1930
rect 406 1934 412 1935
rect 406 1930 407 1934
rect 411 1930 412 1934
rect 406 1929 412 1930
rect 462 1934 468 1935
rect 462 1930 463 1934
rect 467 1930 468 1934
rect 462 1929 468 1930
rect 518 1934 524 1935
rect 518 1930 519 1934
rect 523 1930 524 1934
rect 518 1929 524 1930
rect 582 1934 588 1935
rect 582 1930 583 1934
rect 587 1930 588 1934
rect 582 1929 588 1930
rect 662 1934 668 1935
rect 662 1930 663 1934
rect 667 1930 668 1934
rect 662 1929 668 1930
rect 758 1934 764 1935
rect 758 1930 759 1934
rect 763 1930 764 1934
rect 758 1929 764 1930
rect 878 1934 884 1935
rect 878 1930 879 1934
rect 883 1930 884 1934
rect 878 1929 884 1930
rect 1014 1934 1020 1935
rect 1014 1930 1015 1934
rect 1019 1930 1020 1934
rect 1014 1929 1020 1930
rect 1158 1934 1164 1935
rect 1158 1930 1159 1934
rect 1163 1930 1164 1934
rect 1158 1929 1164 1930
rect 1286 1934 1292 1935
rect 1286 1930 1287 1934
rect 1291 1930 1292 1934
rect 1286 1929 1292 1930
rect 352 1923 354 1929
rect 408 1923 410 1929
rect 464 1923 466 1929
rect 520 1923 522 1929
rect 584 1923 586 1929
rect 664 1923 666 1929
rect 760 1923 762 1929
rect 880 1923 882 1929
rect 1016 1923 1018 1929
rect 1160 1923 1162 1929
rect 1288 1923 1290 1929
rect 1328 1923 1330 1938
rect 1368 1931 1370 1950
rect 1414 1946 1420 1947
rect 1414 1942 1415 1946
rect 1419 1942 1420 1946
rect 1414 1941 1420 1942
rect 1494 1946 1500 1947
rect 1494 1942 1495 1946
rect 1499 1942 1500 1946
rect 1494 1941 1500 1942
rect 1598 1946 1604 1947
rect 1598 1942 1599 1946
rect 1603 1942 1604 1946
rect 1598 1941 1604 1942
rect 1694 1946 1700 1947
rect 1694 1942 1695 1946
rect 1699 1942 1700 1946
rect 1694 1941 1700 1942
rect 1782 1946 1788 1947
rect 1782 1942 1783 1946
rect 1787 1942 1788 1946
rect 1782 1941 1788 1942
rect 1862 1946 1868 1947
rect 1862 1942 1863 1946
rect 1867 1942 1868 1946
rect 1862 1941 1868 1942
rect 1942 1946 1948 1947
rect 1942 1942 1943 1946
rect 1947 1942 1948 1946
rect 1942 1941 1948 1942
rect 2022 1946 2028 1947
rect 2022 1942 2023 1946
rect 2027 1942 2028 1946
rect 2022 1941 2028 1942
rect 2102 1946 2108 1947
rect 2102 1942 2103 1946
rect 2107 1942 2108 1946
rect 2102 1941 2108 1942
rect 1416 1931 1418 1941
rect 1496 1931 1498 1941
rect 1600 1931 1602 1941
rect 1696 1931 1698 1941
rect 1784 1931 1786 1941
rect 1864 1931 1866 1941
rect 1944 1931 1946 1941
rect 2024 1931 2026 1941
rect 2104 1931 2106 1941
rect 2584 1931 2586 1950
rect 1367 1930 1371 1931
rect 1367 1925 1371 1926
rect 1415 1930 1419 1931
rect 1415 1925 1419 1926
rect 1495 1930 1499 1931
rect 1495 1925 1499 1926
rect 1599 1930 1603 1931
rect 1599 1925 1603 1926
rect 1695 1930 1699 1931
rect 1695 1925 1699 1926
rect 1719 1930 1723 1931
rect 1719 1925 1723 1926
rect 1775 1930 1779 1931
rect 1775 1925 1779 1926
rect 1783 1930 1787 1931
rect 1783 1925 1787 1926
rect 1831 1930 1835 1931
rect 1831 1925 1835 1926
rect 1863 1930 1867 1931
rect 1863 1925 1867 1926
rect 1887 1930 1891 1931
rect 1887 1925 1891 1926
rect 1943 1930 1947 1931
rect 1943 1925 1947 1926
rect 1999 1930 2003 1931
rect 1999 1925 2003 1926
rect 2023 1930 2027 1931
rect 2023 1925 2027 1926
rect 2055 1930 2059 1931
rect 2055 1925 2059 1926
rect 2103 1930 2107 1931
rect 2103 1925 2107 1926
rect 2119 1930 2123 1931
rect 2119 1925 2123 1926
rect 2583 1930 2587 1931
rect 2583 1925 2587 1926
rect 111 1922 115 1923
rect 111 1917 115 1918
rect 159 1922 163 1923
rect 159 1917 163 1918
rect 231 1922 235 1923
rect 231 1917 235 1918
rect 327 1922 331 1923
rect 327 1917 331 1918
rect 351 1922 355 1923
rect 351 1917 355 1918
rect 407 1922 411 1923
rect 407 1917 411 1918
rect 431 1922 435 1923
rect 431 1917 435 1918
rect 463 1922 467 1923
rect 463 1917 467 1918
rect 519 1922 523 1923
rect 519 1917 523 1918
rect 543 1922 547 1923
rect 543 1917 547 1918
rect 583 1922 587 1923
rect 583 1917 587 1918
rect 655 1922 659 1923
rect 655 1917 659 1918
rect 663 1922 667 1923
rect 663 1917 667 1918
rect 759 1922 763 1923
rect 759 1917 763 1918
rect 767 1922 771 1923
rect 767 1917 771 1918
rect 879 1922 883 1923
rect 879 1917 883 1918
rect 983 1922 987 1923
rect 983 1917 987 1918
rect 1015 1922 1019 1923
rect 1015 1917 1019 1918
rect 1087 1922 1091 1923
rect 1087 1917 1091 1918
rect 1159 1922 1163 1923
rect 1159 1917 1163 1918
rect 1199 1922 1203 1923
rect 1199 1917 1203 1918
rect 1287 1922 1291 1923
rect 1287 1917 1291 1918
rect 1327 1922 1331 1923
rect 1327 1917 1331 1918
rect 112 1902 114 1917
rect 160 1911 162 1917
rect 232 1911 234 1917
rect 328 1911 330 1917
rect 432 1911 434 1917
rect 544 1911 546 1917
rect 656 1911 658 1917
rect 768 1911 770 1917
rect 880 1911 882 1917
rect 984 1911 986 1917
rect 1088 1911 1090 1917
rect 1200 1911 1202 1917
rect 1288 1911 1290 1917
rect 158 1910 164 1911
rect 158 1906 159 1910
rect 163 1906 164 1910
rect 158 1905 164 1906
rect 230 1910 236 1911
rect 230 1906 231 1910
rect 235 1906 236 1910
rect 230 1905 236 1906
rect 326 1910 332 1911
rect 326 1906 327 1910
rect 331 1906 332 1910
rect 326 1905 332 1906
rect 430 1910 436 1911
rect 430 1906 431 1910
rect 435 1906 436 1910
rect 430 1905 436 1906
rect 542 1910 548 1911
rect 542 1906 543 1910
rect 547 1906 548 1910
rect 542 1905 548 1906
rect 654 1910 660 1911
rect 654 1906 655 1910
rect 659 1906 660 1910
rect 654 1905 660 1906
rect 766 1910 772 1911
rect 766 1906 767 1910
rect 771 1906 772 1910
rect 766 1905 772 1906
rect 878 1910 884 1911
rect 878 1906 879 1910
rect 883 1906 884 1910
rect 878 1905 884 1906
rect 982 1910 988 1911
rect 982 1906 983 1910
rect 987 1906 988 1910
rect 982 1905 988 1906
rect 1086 1910 1092 1911
rect 1086 1906 1087 1910
rect 1091 1906 1092 1910
rect 1086 1905 1092 1906
rect 1198 1910 1204 1911
rect 1198 1906 1199 1910
rect 1203 1906 1204 1910
rect 1198 1905 1204 1906
rect 1286 1910 1292 1911
rect 1286 1906 1287 1910
rect 1291 1906 1292 1910
rect 1286 1905 1292 1906
rect 1328 1902 1330 1917
rect 1368 1910 1370 1925
rect 1720 1919 1722 1925
rect 1776 1919 1778 1925
rect 1832 1919 1834 1925
rect 1888 1919 1890 1925
rect 1944 1919 1946 1925
rect 2000 1919 2002 1925
rect 2056 1919 2058 1925
rect 2120 1919 2122 1925
rect 1718 1918 1724 1919
rect 1718 1914 1719 1918
rect 1723 1914 1724 1918
rect 1718 1913 1724 1914
rect 1774 1918 1780 1919
rect 1774 1914 1775 1918
rect 1779 1914 1780 1918
rect 1774 1913 1780 1914
rect 1830 1918 1836 1919
rect 1830 1914 1831 1918
rect 1835 1914 1836 1918
rect 1830 1913 1836 1914
rect 1886 1918 1892 1919
rect 1886 1914 1887 1918
rect 1891 1914 1892 1918
rect 1886 1913 1892 1914
rect 1942 1918 1948 1919
rect 1942 1914 1943 1918
rect 1947 1914 1948 1918
rect 1942 1913 1948 1914
rect 1998 1918 2004 1919
rect 1998 1914 1999 1918
rect 2003 1914 2004 1918
rect 1998 1913 2004 1914
rect 2054 1918 2060 1919
rect 2054 1914 2055 1918
rect 2059 1914 2060 1918
rect 2054 1913 2060 1914
rect 2118 1918 2124 1919
rect 2118 1914 2119 1918
rect 2123 1914 2124 1918
rect 2118 1913 2124 1914
rect 2584 1910 2586 1925
rect 1366 1909 1372 1910
rect 1366 1905 1367 1909
rect 1371 1905 1372 1909
rect 1366 1904 1372 1905
rect 2582 1909 2588 1910
rect 2582 1905 2583 1909
rect 2587 1905 2588 1909
rect 2582 1904 2588 1905
rect 110 1901 116 1902
rect 110 1897 111 1901
rect 115 1897 116 1901
rect 110 1896 116 1897
rect 1326 1901 1332 1902
rect 1326 1897 1327 1901
rect 1331 1897 1332 1901
rect 1326 1896 1332 1897
rect 1366 1892 1372 1893
rect 2582 1892 2588 1893
rect 1366 1888 1367 1892
rect 1371 1888 1372 1892
rect 1366 1887 1372 1888
rect 1702 1891 1708 1892
rect 1702 1887 1703 1891
rect 1707 1887 1708 1891
rect 110 1884 116 1885
rect 1326 1884 1332 1885
rect 110 1880 111 1884
rect 115 1880 116 1884
rect 110 1879 116 1880
rect 142 1883 148 1884
rect 142 1879 143 1883
rect 147 1879 148 1883
rect 112 1859 114 1879
rect 142 1878 148 1879
rect 214 1883 220 1884
rect 214 1879 215 1883
rect 219 1879 220 1883
rect 214 1878 220 1879
rect 310 1883 316 1884
rect 310 1879 311 1883
rect 315 1879 316 1883
rect 310 1878 316 1879
rect 414 1883 420 1884
rect 414 1879 415 1883
rect 419 1879 420 1883
rect 414 1878 420 1879
rect 526 1883 532 1884
rect 526 1879 527 1883
rect 531 1879 532 1883
rect 526 1878 532 1879
rect 638 1883 644 1884
rect 638 1879 639 1883
rect 643 1879 644 1883
rect 638 1878 644 1879
rect 750 1883 756 1884
rect 750 1879 751 1883
rect 755 1879 756 1883
rect 750 1878 756 1879
rect 862 1883 868 1884
rect 862 1879 863 1883
rect 867 1879 868 1883
rect 862 1878 868 1879
rect 966 1883 972 1884
rect 966 1879 967 1883
rect 971 1879 972 1883
rect 966 1878 972 1879
rect 1070 1883 1076 1884
rect 1070 1879 1071 1883
rect 1075 1879 1076 1883
rect 1070 1878 1076 1879
rect 1182 1883 1188 1884
rect 1182 1879 1183 1883
rect 1187 1879 1188 1883
rect 1182 1878 1188 1879
rect 1270 1883 1276 1884
rect 1270 1879 1271 1883
rect 1275 1879 1276 1883
rect 1326 1880 1327 1884
rect 1331 1880 1332 1884
rect 1326 1879 1332 1880
rect 1270 1878 1276 1879
rect 144 1859 146 1878
rect 216 1859 218 1878
rect 312 1859 314 1878
rect 416 1859 418 1878
rect 528 1859 530 1878
rect 640 1859 642 1878
rect 752 1859 754 1878
rect 864 1859 866 1878
rect 968 1859 970 1878
rect 1072 1859 1074 1878
rect 1184 1859 1186 1878
rect 1272 1859 1274 1878
rect 1328 1859 1330 1879
rect 1368 1871 1370 1887
rect 1702 1886 1708 1887
rect 1758 1891 1764 1892
rect 1758 1887 1759 1891
rect 1763 1887 1764 1891
rect 1758 1886 1764 1887
rect 1814 1891 1820 1892
rect 1814 1887 1815 1891
rect 1819 1887 1820 1891
rect 1814 1886 1820 1887
rect 1870 1891 1876 1892
rect 1870 1887 1871 1891
rect 1875 1887 1876 1891
rect 1870 1886 1876 1887
rect 1926 1891 1932 1892
rect 1926 1887 1927 1891
rect 1931 1887 1932 1891
rect 1926 1886 1932 1887
rect 1982 1891 1988 1892
rect 1982 1887 1983 1891
rect 1987 1887 1988 1891
rect 1982 1886 1988 1887
rect 2038 1891 2044 1892
rect 2038 1887 2039 1891
rect 2043 1887 2044 1891
rect 2038 1886 2044 1887
rect 2102 1891 2108 1892
rect 2102 1887 2103 1891
rect 2107 1887 2108 1891
rect 2582 1888 2583 1892
rect 2587 1888 2588 1892
rect 2582 1887 2588 1888
rect 2102 1886 2108 1887
rect 1704 1871 1706 1886
rect 1760 1871 1762 1886
rect 1816 1871 1818 1886
rect 1872 1871 1874 1886
rect 1928 1871 1930 1886
rect 1984 1871 1986 1886
rect 2040 1871 2042 1886
rect 2104 1871 2106 1886
rect 2584 1871 2586 1887
rect 1367 1870 1371 1871
rect 1367 1865 1371 1866
rect 1399 1870 1403 1871
rect 1399 1865 1403 1866
rect 1463 1870 1467 1871
rect 1463 1865 1467 1866
rect 1559 1870 1563 1871
rect 1559 1865 1563 1866
rect 1655 1870 1659 1871
rect 1655 1865 1659 1866
rect 1703 1870 1707 1871
rect 1703 1865 1707 1866
rect 1743 1870 1747 1871
rect 1743 1865 1747 1866
rect 1759 1870 1763 1871
rect 1759 1865 1763 1866
rect 1815 1870 1819 1871
rect 1815 1865 1819 1866
rect 1831 1870 1835 1871
rect 1831 1865 1835 1866
rect 1871 1870 1875 1871
rect 1871 1865 1875 1866
rect 1919 1870 1923 1871
rect 1919 1865 1923 1866
rect 1927 1870 1931 1871
rect 1927 1865 1931 1866
rect 1983 1870 1987 1871
rect 1983 1865 1987 1866
rect 2007 1870 2011 1871
rect 2007 1865 2011 1866
rect 2039 1870 2043 1871
rect 2039 1865 2043 1866
rect 2095 1870 2099 1871
rect 2095 1865 2099 1866
rect 2103 1870 2107 1871
rect 2103 1865 2107 1866
rect 2183 1870 2187 1871
rect 2183 1865 2187 1866
rect 2583 1870 2587 1871
rect 2583 1865 2587 1866
rect 111 1858 115 1859
rect 111 1853 115 1854
rect 143 1858 147 1859
rect 143 1853 147 1854
rect 199 1858 203 1859
rect 199 1853 203 1854
rect 215 1858 219 1859
rect 215 1853 219 1854
rect 263 1858 267 1859
rect 263 1853 267 1854
rect 311 1858 315 1859
rect 311 1853 315 1854
rect 351 1858 355 1859
rect 351 1853 355 1854
rect 415 1858 419 1859
rect 415 1853 419 1854
rect 439 1858 443 1859
rect 439 1853 443 1854
rect 527 1858 531 1859
rect 527 1853 531 1854
rect 535 1858 539 1859
rect 535 1853 539 1854
rect 623 1858 627 1859
rect 623 1853 627 1854
rect 639 1858 643 1859
rect 639 1853 643 1854
rect 711 1858 715 1859
rect 711 1853 715 1854
rect 751 1858 755 1859
rect 751 1853 755 1854
rect 791 1858 795 1859
rect 791 1853 795 1854
rect 863 1858 867 1859
rect 863 1853 867 1854
rect 871 1858 875 1859
rect 871 1853 875 1854
rect 951 1858 955 1859
rect 951 1853 955 1854
rect 967 1858 971 1859
rect 967 1853 971 1854
rect 1039 1858 1043 1859
rect 1039 1853 1043 1854
rect 1071 1858 1075 1859
rect 1071 1853 1075 1854
rect 1183 1858 1187 1859
rect 1183 1853 1187 1854
rect 1271 1858 1275 1859
rect 1271 1853 1275 1854
rect 1327 1858 1331 1859
rect 1327 1853 1331 1854
rect 1368 1853 1370 1865
rect 1400 1854 1402 1865
rect 1464 1854 1466 1865
rect 1560 1854 1562 1865
rect 1656 1854 1658 1865
rect 1744 1854 1746 1865
rect 1832 1854 1834 1865
rect 1920 1854 1922 1865
rect 2008 1854 2010 1865
rect 2096 1854 2098 1865
rect 2184 1854 2186 1865
rect 1398 1853 1404 1854
rect 112 1841 114 1853
rect 144 1842 146 1853
rect 200 1842 202 1853
rect 264 1842 266 1853
rect 352 1842 354 1853
rect 440 1842 442 1853
rect 536 1842 538 1853
rect 624 1842 626 1853
rect 712 1842 714 1853
rect 792 1842 794 1853
rect 872 1842 874 1853
rect 952 1842 954 1853
rect 1040 1842 1042 1853
rect 142 1841 148 1842
rect 110 1840 116 1841
rect 110 1836 111 1840
rect 115 1836 116 1840
rect 142 1837 143 1841
rect 147 1837 148 1841
rect 142 1836 148 1837
rect 198 1841 204 1842
rect 198 1837 199 1841
rect 203 1837 204 1841
rect 198 1836 204 1837
rect 262 1841 268 1842
rect 262 1837 263 1841
rect 267 1837 268 1841
rect 262 1836 268 1837
rect 350 1841 356 1842
rect 350 1837 351 1841
rect 355 1837 356 1841
rect 350 1836 356 1837
rect 438 1841 444 1842
rect 438 1837 439 1841
rect 443 1837 444 1841
rect 438 1836 444 1837
rect 534 1841 540 1842
rect 534 1837 535 1841
rect 539 1837 540 1841
rect 534 1836 540 1837
rect 622 1841 628 1842
rect 622 1837 623 1841
rect 627 1837 628 1841
rect 622 1836 628 1837
rect 710 1841 716 1842
rect 710 1837 711 1841
rect 715 1837 716 1841
rect 710 1836 716 1837
rect 790 1841 796 1842
rect 790 1837 791 1841
rect 795 1837 796 1841
rect 790 1836 796 1837
rect 870 1841 876 1842
rect 870 1837 871 1841
rect 875 1837 876 1841
rect 870 1836 876 1837
rect 950 1841 956 1842
rect 950 1837 951 1841
rect 955 1837 956 1841
rect 950 1836 956 1837
rect 1038 1841 1044 1842
rect 1328 1841 1330 1853
rect 1366 1852 1372 1853
rect 1366 1848 1367 1852
rect 1371 1848 1372 1852
rect 1398 1849 1399 1853
rect 1403 1849 1404 1853
rect 1398 1848 1404 1849
rect 1462 1853 1468 1854
rect 1462 1849 1463 1853
rect 1467 1849 1468 1853
rect 1462 1848 1468 1849
rect 1558 1853 1564 1854
rect 1558 1849 1559 1853
rect 1563 1849 1564 1853
rect 1558 1848 1564 1849
rect 1654 1853 1660 1854
rect 1654 1849 1655 1853
rect 1659 1849 1660 1853
rect 1654 1848 1660 1849
rect 1742 1853 1748 1854
rect 1742 1849 1743 1853
rect 1747 1849 1748 1853
rect 1742 1848 1748 1849
rect 1830 1853 1836 1854
rect 1830 1849 1831 1853
rect 1835 1849 1836 1853
rect 1830 1848 1836 1849
rect 1918 1853 1924 1854
rect 1918 1849 1919 1853
rect 1923 1849 1924 1853
rect 1918 1848 1924 1849
rect 2006 1853 2012 1854
rect 2006 1849 2007 1853
rect 2011 1849 2012 1853
rect 2006 1848 2012 1849
rect 2094 1853 2100 1854
rect 2094 1849 2095 1853
rect 2099 1849 2100 1853
rect 2094 1848 2100 1849
rect 2182 1853 2188 1854
rect 2584 1853 2586 1865
rect 2182 1849 2183 1853
rect 2187 1849 2188 1853
rect 2182 1848 2188 1849
rect 2582 1852 2588 1853
rect 2582 1848 2583 1852
rect 2587 1848 2588 1852
rect 1366 1847 1372 1848
rect 2582 1847 2588 1848
rect 1038 1837 1039 1841
rect 1043 1837 1044 1841
rect 1038 1836 1044 1837
rect 1326 1840 1332 1841
rect 1326 1836 1327 1840
rect 1331 1836 1332 1840
rect 110 1835 116 1836
rect 1326 1835 1332 1836
rect 1366 1835 1372 1836
rect 1366 1831 1367 1835
rect 1371 1831 1372 1835
rect 1366 1830 1372 1831
rect 2582 1835 2588 1836
rect 2582 1831 2583 1835
rect 2587 1831 2588 1835
rect 2582 1830 2588 1831
rect 110 1823 116 1824
rect 110 1819 111 1823
rect 115 1819 116 1823
rect 110 1818 116 1819
rect 1326 1823 1332 1824
rect 1326 1819 1327 1823
rect 1331 1819 1332 1823
rect 1326 1818 1332 1819
rect 112 1799 114 1818
rect 158 1814 164 1815
rect 158 1810 159 1814
rect 163 1810 164 1814
rect 158 1809 164 1810
rect 214 1814 220 1815
rect 214 1810 215 1814
rect 219 1810 220 1814
rect 214 1809 220 1810
rect 278 1814 284 1815
rect 278 1810 279 1814
rect 283 1810 284 1814
rect 278 1809 284 1810
rect 366 1814 372 1815
rect 366 1810 367 1814
rect 371 1810 372 1814
rect 366 1809 372 1810
rect 454 1814 460 1815
rect 454 1810 455 1814
rect 459 1810 460 1814
rect 454 1809 460 1810
rect 550 1814 556 1815
rect 550 1810 551 1814
rect 555 1810 556 1814
rect 550 1809 556 1810
rect 638 1814 644 1815
rect 638 1810 639 1814
rect 643 1810 644 1814
rect 638 1809 644 1810
rect 726 1814 732 1815
rect 726 1810 727 1814
rect 731 1810 732 1814
rect 726 1809 732 1810
rect 806 1814 812 1815
rect 806 1810 807 1814
rect 811 1810 812 1814
rect 806 1809 812 1810
rect 886 1814 892 1815
rect 886 1810 887 1814
rect 891 1810 892 1814
rect 886 1809 892 1810
rect 966 1814 972 1815
rect 966 1810 967 1814
rect 971 1810 972 1814
rect 966 1809 972 1810
rect 1054 1814 1060 1815
rect 1054 1810 1055 1814
rect 1059 1810 1060 1814
rect 1054 1809 1060 1810
rect 160 1799 162 1809
rect 216 1799 218 1809
rect 280 1799 282 1809
rect 368 1799 370 1809
rect 456 1799 458 1809
rect 552 1799 554 1809
rect 640 1799 642 1809
rect 728 1799 730 1809
rect 808 1799 810 1809
rect 888 1799 890 1809
rect 968 1799 970 1809
rect 1056 1799 1058 1809
rect 1328 1799 1330 1818
rect 1368 1815 1370 1830
rect 1414 1826 1420 1827
rect 1414 1822 1415 1826
rect 1419 1822 1420 1826
rect 1414 1821 1420 1822
rect 1478 1826 1484 1827
rect 1478 1822 1479 1826
rect 1483 1822 1484 1826
rect 1478 1821 1484 1822
rect 1574 1826 1580 1827
rect 1574 1822 1575 1826
rect 1579 1822 1580 1826
rect 1574 1821 1580 1822
rect 1670 1826 1676 1827
rect 1670 1822 1671 1826
rect 1675 1822 1676 1826
rect 1670 1821 1676 1822
rect 1758 1826 1764 1827
rect 1758 1822 1759 1826
rect 1763 1822 1764 1826
rect 1758 1821 1764 1822
rect 1846 1826 1852 1827
rect 1846 1822 1847 1826
rect 1851 1822 1852 1826
rect 1846 1821 1852 1822
rect 1934 1826 1940 1827
rect 1934 1822 1935 1826
rect 1939 1822 1940 1826
rect 1934 1821 1940 1822
rect 2022 1826 2028 1827
rect 2022 1822 2023 1826
rect 2027 1822 2028 1826
rect 2022 1821 2028 1822
rect 2110 1826 2116 1827
rect 2110 1822 2111 1826
rect 2115 1822 2116 1826
rect 2110 1821 2116 1822
rect 2198 1826 2204 1827
rect 2198 1822 2199 1826
rect 2203 1822 2204 1826
rect 2198 1821 2204 1822
rect 1416 1815 1418 1821
rect 1480 1815 1482 1821
rect 1576 1815 1578 1821
rect 1672 1815 1674 1821
rect 1760 1815 1762 1821
rect 1848 1815 1850 1821
rect 1936 1815 1938 1821
rect 2024 1815 2026 1821
rect 2112 1815 2114 1821
rect 2200 1815 2202 1821
rect 2584 1815 2586 1830
rect 1367 1814 1371 1815
rect 1367 1809 1371 1810
rect 1415 1814 1419 1815
rect 1415 1809 1419 1810
rect 1479 1814 1483 1815
rect 1479 1809 1483 1810
rect 1511 1814 1515 1815
rect 1511 1809 1515 1810
rect 1575 1814 1579 1815
rect 1575 1809 1579 1810
rect 1623 1814 1627 1815
rect 1623 1809 1627 1810
rect 1671 1814 1675 1815
rect 1671 1809 1675 1810
rect 1735 1814 1739 1815
rect 1735 1809 1739 1810
rect 1759 1814 1763 1815
rect 1759 1809 1763 1810
rect 1839 1814 1843 1815
rect 1839 1809 1843 1810
rect 1847 1814 1851 1815
rect 1847 1809 1851 1810
rect 1935 1814 1939 1815
rect 1935 1809 1939 1810
rect 1951 1814 1955 1815
rect 1951 1809 1955 1810
rect 2023 1814 2027 1815
rect 2023 1809 2027 1810
rect 2063 1814 2067 1815
rect 2063 1809 2067 1810
rect 2111 1814 2115 1815
rect 2111 1809 2115 1810
rect 2183 1814 2187 1815
rect 2183 1809 2187 1810
rect 2199 1814 2203 1815
rect 2199 1809 2203 1810
rect 2303 1814 2307 1815
rect 2303 1809 2307 1810
rect 2431 1814 2435 1815
rect 2431 1809 2435 1810
rect 2543 1814 2547 1815
rect 2543 1809 2547 1810
rect 2583 1814 2587 1815
rect 2583 1809 2587 1810
rect 111 1798 115 1799
rect 111 1793 115 1794
rect 159 1798 163 1799
rect 159 1793 163 1794
rect 215 1798 219 1799
rect 215 1793 219 1794
rect 231 1798 235 1799
rect 231 1793 235 1794
rect 279 1798 283 1799
rect 279 1793 283 1794
rect 295 1798 299 1799
rect 295 1793 299 1794
rect 367 1798 371 1799
rect 367 1793 371 1794
rect 447 1798 451 1799
rect 447 1793 451 1794
rect 455 1798 459 1799
rect 455 1793 459 1794
rect 535 1798 539 1799
rect 535 1793 539 1794
rect 551 1798 555 1799
rect 551 1793 555 1794
rect 623 1798 627 1799
rect 623 1793 627 1794
rect 639 1798 643 1799
rect 639 1793 643 1794
rect 711 1798 715 1799
rect 711 1793 715 1794
rect 727 1798 731 1799
rect 727 1793 731 1794
rect 791 1798 795 1799
rect 791 1793 795 1794
rect 807 1798 811 1799
rect 807 1793 811 1794
rect 871 1798 875 1799
rect 871 1793 875 1794
rect 887 1798 891 1799
rect 887 1793 891 1794
rect 951 1798 955 1799
rect 951 1793 955 1794
rect 967 1798 971 1799
rect 967 1793 971 1794
rect 1031 1798 1035 1799
rect 1031 1793 1035 1794
rect 1055 1798 1059 1799
rect 1055 1793 1059 1794
rect 1119 1798 1123 1799
rect 1119 1793 1123 1794
rect 1327 1798 1331 1799
rect 1368 1794 1370 1809
rect 1416 1803 1418 1809
rect 1512 1803 1514 1809
rect 1624 1803 1626 1809
rect 1736 1803 1738 1809
rect 1840 1803 1842 1809
rect 1952 1803 1954 1809
rect 2064 1803 2066 1809
rect 2184 1803 2186 1809
rect 2304 1803 2306 1809
rect 2432 1803 2434 1809
rect 2544 1803 2546 1809
rect 1414 1802 1420 1803
rect 1414 1798 1415 1802
rect 1419 1798 1420 1802
rect 1414 1797 1420 1798
rect 1510 1802 1516 1803
rect 1510 1798 1511 1802
rect 1515 1798 1516 1802
rect 1510 1797 1516 1798
rect 1622 1802 1628 1803
rect 1622 1798 1623 1802
rect 1627 1798 1628 1802
rect 1622 1797 1628 1798
rect 1734 1802 1740 1803
rect 1734 1798 1735 1802
rect 1739 1798 1740 1802
rect 1734 1797 1740 1798
rect 1838 1802 1844 1803
rect 1838 1798 1839 1802
rect 1843 1798 1844 1802
rect 1838 1797 1844 1798
rect 1950 1802 1956 1803
rect 1950 1798 1951 1802
rect 1955 1798 1956 1802
rect 1950 1797 1956 1798
rect 2062 1802 2068 1803
rect 2062 1798 2063 1802
rect 2067 1798 2068 1802
rect 2062 1797 2068 1798
rect 2182 1802 2188 1803
rect 2182 1798 2183 1802
rect 2187 1798 2188 1802
rect 2182 1797 2188 1798
rect 2302 1802 2308 1803
rect 2302 1798 2303 1802
rect 2307 1798 2308 1802
rect 2302 1797 2308 1798
rect 2430 1802 2436 1803
rect 2430 1798 2431 1802
rect 2435 1798 2436 1802
rect 2430 1797 2436 1798
rect 2542 1802 2548 1803
rect 2542 1798 2543 1802
rect 2547 1798 2548 1802
rect 2542 1797 2548 1798
rect 2584 1794 2586 1809
rect 1327 1793 1331 1794
rect 1366 1793 1372 1794
rect 112 1778 114 1793
rect 232 1787 234 1793
rect 296 1787 298 1793
rect 368 1787 370 1793
rect 448 1787 450 1793
rect 536 1787 538 1793
rect 624 1787 626 1793
rect 712 1787 714 1793
rect 792 1787 794 1793
rect 872 1787 874 1793
rect 952 1787 954 1793
rect 1032 1787 1034 1793
rect 1120 1787 1122 1793
rect 230 1786 236 1787
rect 230 1782 231 1786
rect 235 1782 236 1786
rect 230 1781 236 1782
rect 294 1786 300 1787
rect 294 1782 295 1786
rect 299 1782 300 1786
rect 294 1781 300 1782
rect 366 1786 372 1787
rect 366 1782 367 1786
rect 371 1782 372 1786
rect 366 1781 372 1782
rect 446 1786 452 1787
rect 446 1782 447 1786
rect 451 1782 452 1786
rect 446 1781 452 1782
rect 534 1786 540 1787
rect 534 1782 535 1786
rect 539 1782 540 1786
rect 534 1781 540 1782
rect 622 1786 628 1787
rect 622 1782 623 1786
rect 627 1782 628 1786
rect 622 1781 628 1782
rect 710 1786 716 1787
rect 710 1782 711 1786
rect 715 1782 716 1786
rect 710 1781 716 1782
rect 790 1786 796 1787
rect 790 1782 791 1786
rect 795 1782 796 1786
rect 790 1781 796 1782
rect 870 1786 876 1787
rect 870 1782 871 1786
rect 875 1782 876 1786
rect 870 1781 876 1782
rect 950 1786 956 1787
rect 950 1782 951 1786
rect 955 1782 956 1786
rect 950 1781 956 1782
rect 1030 1786 1036 1787
rect 1030 1782 1031 1786
rect 1035 1782 1036 1786
rect 1030 1781 1036 1782
rect 1118 1786 1124 1787
rect 1118 1782 1119 1786
rect 1123 1782 1124 1786
rect 1118 1781 1124 1782
rect 1328 1778 1330 1793
rect 1366 1789 1367 1793
rect 1371 1789 1372 1793
rect 1366 1788 1372 1789
rect 2582 1793 2588 1794
rect 2582 1789 2583 1793
rect 2587 1789 2588 1793
rect 2582 1788 2588 1789
rect 110 1777 116 1778
rect 110 1773 111 1777
rect 115 1773 116 1777
rect 110 1772 116 1773
rect 1326 1777 1332 1778
rect 1326 1773 1327 1777
rect 1331 1773 1332 1777
rect 1326 1772 1332 1773
rect 1366 1776 1372 1777
rect 2582 1776 2588 1777
rect 1366 1772 1367 1776
rect 1371 1772 1372 1776
rect 1366 1771 1372 1772
rect 1398 1775 1404 1776
rect 1398 1771 1399 1775
rect 1403 1771 1404 1775
rect 110 1760 116 1761
rect 1326 1760 1332 1761
rect 110 1756 111 1760
rect 115 1756 116 1760
rect 110 1755 116 1756
rect 214 1759 220 1760
rect 214 1755 215 1759
rect 219 1755 220 1759
rect 112 1739 114 1755
rect 214 1754 220 1755
rect 278 1759 284 1760
rect 278 1755 279 1759
rect 283 1755 284 1759
rect 278 1754 284 1755
rect 350 1759 356 1760
rect 350 1755 351 1759
rect 355 1755 356 1759
rect 350 1754 356 1755
rect 430 1759 436 1760
rect 430 1755 431 1759
rect 435 1755 436 1759
rect 430 1754 436 1755
rect 518 1759 524 1760
rect 518 1755 519 1759
rect 523 1755 524 1759
rect 518 1754 524 1755
rect 606 1759 612 1760
rect 606 1755 607 1759
rect 611 1755 612 1759
rect 606 1754 612 1755
rect 694 1759 700 1760
rect 694 1755 695 1759
rect 699 1755 700 1759
rect 694 1754 700 1755
rect 774 1759 780 1760
rect 774 1755 775 1759
rect 779 1755 780 1759
rect 774 1754 780 1755
rect 854 1759 860 1760
rect 854 1755 855 1759
rect 859 1755 860 1759
rect 854 1754 860 1755
rect 934 1759 940 1760
rect 934 1755 935 1759
rect 939 1755 940 1759
rect 934 1754 940 1755
rect 1014 1759 1020 1760
rect 1014 1755 1015 1759
rect 1019 1755 1020 1759
rect 1014 1754 1020 1755
rect 1102 1759 1108 1760
rect 1102 1755 1103 1759
rect 1107 1755 1108 1759
rect 1326 1756 1327 1760
rect 1331 1756 1332 1760
rect 1368 1759 1370 1771
rect 1398 1770 1404 1771
rect 1494 1775 1500 1776
rect 1494 1771 1495 1775
rect 1499 1771 1500 1775
rect 1494 1770 1500 1771
rect 1606 1775 1612 1776
rect 1606 1771 1607 1775
rect 1611 1771 1612 1775
rect 1606 1770 1612 1771
rect 1718 1775 1724 1776
rect 1718 1771 1719 1775
rect 1723 1771 1724 1775
rect 1718 1770 1724 1771
rect 1822 1775 1828 1776
rect 1822 1771 1823 1775
rect 1827 1771 1828 1775
rect 1822 1770 1828 1771
rect 1934 1775 1940 1776
rect 1934 1771 1935 1775
rect 1939 1771 1940 1775
rect 1934 1770 1940 1771
rect 2046 1775 2052 1776
rect 2046 1771 2047 1775
rect 2051 1771 2052 1775
rect 2046 1770 2052 1771
rect 2166 1775 2172 1776
rect 2166 1771 2167 1775
rect 2171 1771 2172 1775
rect 2166 1770 2172 1771
rect 2286 1775 2292 1776
rect 2286 1771 2287 1775
rect 2291 1771 2292 1775
rect 2286 1770 2292 1771
rect 2414 1775 2420 1776
rect 2414 1771 2415 1775
rect 2419 1771 2420 1775
rect 2414 1770 2420 1771
rect 2526 1775 2532 1776
rect 2526 1771 2527 1775
rect 2531 1771 2532 1775
rect 2582 1772 2583 1776
rect 2587 1772 2588 1776
rect 2582 1771 2588 1772
rect 2526 1770 2532 1771
rect 1400 1759 1402 1770
rect 1496 1759 1498 1770
rect 1608 1759 1610 1770
rect 1720 1759 1722 1770
rect 1824 1759 1826 1770
rect 1936 1759 1938 1770
rect 2048 1759 2050 1770
rect 2168 1759 2170 1770
rect 2288 1759 2290 1770
rect 2416 1759 2418 1770
rect 2528 1759 2530 1770
rect 2584 1759 2586 1771
rect 1326 1755 1332 1756
rect 1367 1758 1371 1759
rect 1102 1754 1108 1755
rect 216 1739 218 1754
rect 280 1739 282 1754
rect 352 1739 354 1754
rect 432 1739 434 1754
rect 520 1739 522 1754
rect 608 1739 610 1754
rect 696 1739 698 1754
rect 776 1739 778 1754
rect 856 1739 858 1754
rect 936 1739 938 1754
rect 1016 1739 1018 1754
rect 1104 1739 1106 1754
rect 1328 1739 1330 1755
rect 1367 1753 1371 1754
rect 1399 1758 1403 1759
rect 1399 1753 1403 1754
rect 1439 1758 1443 1759
rect 1439 1753 1443 1754
rect 1495 1758 1499 1759
rect 1495 1753 1499 1754
rect 1519 1758 1523 1759
rect 1519 1753 1523 1754
rect 1607 1758 1611 1759
rect 1607 1753 1611 1754
rect 1615 1758 1619 1759
rect 1615 1753 1619 1754
rect 1719 1758 1723 1759
rect 1719 1753 1723 1754
rect 1823 1758 1827 1759
rect 1823 1753 1827 1754
rect 1927 1758 1931 1759
rect 1927 1753 1931 1754
rect 1935 1758 1939 1759
rect 1935 1753 1939 1754
rect 2023 1758 2027 1759
rect 2023 1753 2027 1754
rect 2047 1758 2051 1759
rect 2047 1753 2051 1754
rect 2119 1758 2123 1759
rect 2119 1753 2123 1754
rect 2167 1758 2171 1759
rect 2167 1753 2171 1754
rect 2207 1758 2211 1759
rect 2207 1753 2211 1754
rect 2287 1758 2291 1759
rect 2287 1753 2291 1754
rect 2375 1758 2379 1759
rect 2375 1753 2379 1754
rect 2415 1758 2419 1759
rect 2415 1753 2419 1754
rect 2463 1758 2467 1759
rect 2463 1753 2467 1754
rect 2527 1758 2531 1759
rect 2527 1753 2531 1754
rect 2583 1758 2587 1759
rect 2583 1753 2587 1754
rect 1368 1741 1370 1753
rect 1440 1742 1442 1753
rect 1520 1742 1522 1753
rect 1616 1742 1618 1753
rect 1720 1742 1722 1753
rect 1824 1742 1826 1753
rect 1928 1742 1930 1753
rect 2024 1742 2026 1753
rect 2120 1742 2122 1753
rect 2208 1742 2210 1753
rect 2288 1742 2290 1753
rect 2376 1742 2378 1753
rect 2464 1742 2466 1753
rect 2528 1742 2530 1753
rect 1438 1741 1444 1742
rect 1366 1740 1372 1741
rect 111 1738 115 1739
rect 111 1733 115 1734
rect 215 1738 219 1739
rect 215 1733 219 1734
rect 279 1738 283 1739
rect 279 1733 283 1734
rect 351 1738 355 1739
rect 351 1733 355 1734
rect 407 1738 411 1739
rect 407 1733 411 1734
rect 431 1738 435 1739
rect 431 1733 435 1734
rect 471 1738 475 1739
rect 471 1733 475 1734
rect 519 1738 523 1739
rect 519 1733 523 1734
rect 551 1738 555 1739
rect 551 1733 555 1734
rect 607 1738 611 1739
rect 607 1733 611 1734
rect 639 1738 643 1739
rect 639 1733 643 1734
rect 695 1738 699 1739
rect 695 1733 699 1734
rect 727 1738 731 1739
rect 727 1733 731 1734
rect 775 1738 779 1739
rect 775 1733 779 1734
rect 823 1738 827 1739
rect 823 1733 827 1734
rect 855 1738 859 1739
rect 855 1733 859 1734
rect 919 1738 923 1739
rect 919 1733 923 1734
rect 935 1738 939 1739
rect 935 1733 939 1734
rect 1015 1738 1019 1739
rect 1015 1733 1019 1734
rect 1103 1738 1107 1739
rect 1103 1733 1107 1734
rect 1111 1738 1115 1739
rect 1111 1733 1115 1734
rect 1207 1738 1211 1739
rect 1207 1733 1211 1734
rect 1327 1738 1331 1739
rect 1366 1736 1367 1740
rect 1371 1736 1372 1740
rect 1438 1737 1439 1741
rect 1443 1737 1444 1741
rect 1438 1736 1444 1737
rect 1518 1741 1524 1742
rect 1518 1737 1519 1741
rect 1523 1737 1524 1741
rect 1518 1736 1524 1737
rect 1614 1741 1620 1742
rect 1614 1737 1615 1741
rect 1619 1737 1620 1741
rect 1614 1736 1620 1737
rect 1718 1741 1724 1742
rect 1718 1737 1719 1741
rect 1723 1737 1724 1741
rect 1718 1736 1724 1737
rect 1822 1741 1828 1742
rect 1822 1737 1823 1741
rect 1827 1737 1828 1741
rect 1822 1736 1828 1737
rect 1926 1741 1932 1742
rect 1926 1737 1927 1741
rect 1931 1737 1932 1741
rect 1926 1736 1932 1737
rect 2022 1741 2028 1742
rect 2022 1737 2023 1741
rect 2027 1737 2028 1741
rect 2022 1736 2028 1737
rect 2118 1741 2124 1742
rect 2118 1737 2119 1741
rect 2123 1737 2124 1741
rect 2118 1736 2124 1737
rect 2206 1741 2212 1742
rect 2206 1737 2207 1741
rect 2211 1737 2212 1741
rect 2206 1736 2212 1737
rect 2286 1741 2292 1742
rect 2286 1737 2287 1741
rect 2291 1737 2292 1741
rect 2286 1736 2292 1737
rect 2374 1741 2380 1742
rect 2374 1737 2375 1741
rect 2379 1737 2380 1741
rect 2374 1736 2380 1737
rect 2462 1741 2468 1742
rect 2462 1737 2463 1741
rect 2467 1737 2468 1741
rect 2462 1736 2468 1737
rect 2526 1741 2532 1742
rect 2584 1741 2586 1753
rect 2526 1737 2527 1741
rect 2531 1737 2532 1741
rect 2526 1736 2532 1737
rect 2582 1740 2588 1741
rect 2582 1736 2583 1740
rect 2587 1736 2588 1740
rect 1366 1735 1372 1736
rect 2582 1735 2588 1736
rect 1327 1733 1331 1734
rect 112 1721 114 1733
rect 352 1722 354 1733
rect 408 1722 410 1733
rect 472 1722 474 1733
rect 552 1722 554 1733
rect 640 1722 642 1733
rect 728 1722 730 1733
rect 824 1722 826 1733
rect 920 1722 922 1733
rect 1016 1722 1018 1733
rect 1112 1722 1114 1733
rect 1208 1722 1210 1733
rect 350 1721 356 1722
rect 110 1720 116 1721
rect 110 1716 111 1720
rect 115 1716 116 1720
rect 350 1717 351 1721
rect 355 1717 356 1721
rect 350 1716 356 1717
rect 406 1721 412 1722
rect 406 1717 407 1721
rect 411 1717 412 1721
rect 406 1716 412 1717
rect 470 1721 476 1722
rect 470 1717 471 1721
rect 475 1717 476 1721
rect 470 1716 476 1717
rect 550 1721 556 1722
rect 550 1717 551 1721
rect 555 1717 556 1721
rect 550 1716 556 1717
rect 638 1721 644 1722
rect 638 1717 639 1721
rect 643 1717 644 1721
rect 638 1716 644 1717
rect 726 1721 732 1722
rect 726 1717 727 1721
rect 731 1717 732 1721
rect 726 1716 732 1717
rect 822 1721 828 1722
rect 822 1717 823 1721
rect 827 1717 828 1721
rect 822 1716 828 1717
rect 918 1721 924 1722
rect 918 1717 919 1721
rect 923 1717 924 1721
rect 918 1716 924 1717
rect 1014 1721 1020 1722
rect 1014 1717 1015 1721
rect 1019 1717 1020 1721
rect 1014 1716 1020 1717
rect 1110 1721 1116 1722
rect 1110 1717 1111 1721
rect 1115 1717 1116 1721
rect 1110 1716 1116 1717
rect 1206 1721 1212 1722
rect 1328 1721 1330 1733
rect 1366 1723 1372 1724
rect 1206 1717 1207 1721
rect 1211 1717 1212 1721
rect 1206 1716 1212 1717
rect 1326 1720 1332 1721
rect 1326 1716 1327 1720
rect 1331 1716 1332 1720
rect 1366 1719 1367 1723
rect 1371 1719 1372 1723
rect 1366 1718 1372 1719
rect 2582 1723 2588 1724
rect 2582 1719 2583 1723
rect 2587 1719 2588 1723
rect 2582 1718 2588 1719
rect 110 1715 116 1716
rect 1326 1715 1332 1716
rect 110 1703 116 1704
rect 110 1699 111 1703
rect 115 1699 116 1703
rect 110 1698 116 1699
rect 1326 1703 1332 1704
rect 1326 1699 1327 1703
rect 1331 1699 1332 1703
rect 1326 1698 1332 1699
rect 112 1679 114 1698
rect 366 1694 372 1695
rect 366 1690 367 1694
rect 371 1690 372 1694
rect 366 1689 372 1690
rect 422 1694 428 1695
rect 422 1690 423 1694
rect 427 1690 428 1694
rect 422 1689 428 1690
rect 486 1694 492 1695
rect 486 1690 487 1694
rect 491 1690 492 1694
rect 486 1689 492 1690
rect 566 1694 572 1695
rect 566 1690 567 1694
rect 571 1690 572 1694
rect 566 1689 572 1690
rect 654 1694 660 1695
rect 654 1690 655 1694
rect 659 1690 660 1694
rect 654 1689 660 1690
rect 742 1694 748 1695
rect 742 1690 743 1694
rect 747 1690 748 1694
rect 742 1689 748 1690
rect 838 1694 844 1695
rect 838 1690 839 1694
rect 843 1690 844 1694
rect 838 1689 844 1690
rect 934 1694 940 1695
rect 934 1690 935 1694
rect 939 1690 940 1694
rect 934 1689 940 1690
rect 1030 1694 1036 1695
rect 1030 1690 1031 1694
rect 1035 1690 1036 1694
rect 1030 1689 1036 1690
rect 1126 1694 1132 1695
rect 1126 1690 1127 1694
rect 1131 1690 1132 1694
rect 1126 1689 1132 1690
rect 1222 1694 1228 1695
rect 1222 1690 1223 1694
rect 1227 1690 1228 1694
rect 1222 1689 1228 1690
rect 368 1679 370 1689
rect 424 1679 426 1689
rect 488 1679 490 1689
rect 568 1679 570 1689
rect 656 1679 658 1689
rect 744 1679 746 1689
rect 840 1679 842 1689
rect 936 1679 938 1689
rect 1032 1679 1034 1689
rect 1128 1679 1130 1689
rect 1224 1679 1226 1689
rect 1328 1679 1330 1698
rect 1368 1691 1370 1718
rect 1454 1714 1460 1715
rect 1454 1710 1455 1714
rect 1459 1710 1460 1714
rect 1454 1709 1460 1710
rect 1534 1714 1540 1715
rect 1534 1710 1535 1714
rect 1539 1710 1540 1714
rect 1534 1709 1540 1710
rect 1630 1714 1636 1715
rect 1630 1710 1631 1714
rect 1635 1710 1636 1714
rect 1630 1709 1636 1710
rect 1734 1714 1740 1715
rect 1734 1710 1735 1714
rect 1739 1710 1740 1714
rect 1734 1709 1740 1710
rect 1838 1714 1844 1715
rect 1838 1710 1839 1714
rect 1843 1710 1844 1714
rect 1838 1709 1844 1710
rect 1942 1714 1948 1715
rect 1942 1710 1943 1714
rect 1947 1710 1948 1714
rect 1942 1709 1948 1710
rect 2038 1714 2044 1715
rect 2038 1710 2039 1714
rect 2043 1710 2044 1714
rect 2038 1709 2044 1710
rect 2134 1714 2140 1715
rect 2134 1710 2135 1714
rect 2139 1710 2140 1714
rect 2134 1709 2140 1710
rect 2222 1714 2228 1715
rect 2222 1710 2223 1714
rect 2227 1710 2228 1714
rect 2222 1709 2228 1710
rect 2302 1714 2308 1715
rect 2302 1710 2303 1714
rect 2307 1710 2308 1714
rect 2302 1709 2308 1710
rect 2390 1714 2396 1715
rect 2390 1710 2391 1714
rect 2395 1710 2396 1714
rect 2390 1709 2396 1710
rect 2478 1714 2484 1715
rect 2478 1710 2479 1714
rect 2483 1710 2484 1714
rect 2478 1709 2484 1710
rect 2542 1714 2548 1715
rect 2542 1710 2543 1714
rect 2547 1710 2548 1714
rect 2542 1709 2548 1710
rect 1456 1691 1458 1709
rect 1536 1691 1538 1709
rect 1632 1691 1634 1709
rect 1736 1691 1738 1709
rect 1840 1691 1842 1709
rect 1944 1691 1946 1709
rect 2040 1691 2042 1709
rect 2136 1691 2138 1709
rect 2224 1691 2226 1709
rect 2304 1691 2306 1709
rect 2392 1691 2394 1709
rect 2480 1691 2482 1709
rect 2544 1691 2546 1709
rect 2584 1691 2586 1718
rect 1367 1690 1371 1691
rect 1367 1685 1371 1686
rect 1455 1690 1459 1691
rect 1455 1685 1459 1686
rect 1535 1690 1539 1691
rect 1535 1685 1539 1686
rect 1559 1690 1563 1691
rect 1559 1685 1563 1686
rect 1631 1690 1635 1691
rect 1631 1685 1635 1686
rect 1711 1690 1715 1691
rect 1711 1685 1715 1686
rect 1735 1690 1739 1691
rect 1735 1685 1739 1686
rect 1799 1690 1803 1691
rect 1799 1685 1803 1686
rect 1839 1690 1843 1691
rect 1839 1685 1843 1686
rect 1887 1690 1891 1691
rect 1887 1685 1891 1686
rect 1943 1690 1947 1691
rect 1943 1685 1947 1686
rect 1975 1690 1979 1691
rect 1975 1685 1979 1686
rect 2039 1690 2043 1691
rect 2039 1685 2043 1686
rect 2063 1690 2067 1691
rect 2063 1685 2067 1686
rect 2135 1690 2139 1691
rect 2135 1685 2139 1686
rect 2143 1690 2147 1691
rect 2143 1685 2147 1686
rect 2215 1690 2219 1691
rect 2215 1685 2219 1686
rect 2223 1690 2227 1691
rect 2223 1685 2227 1686
rect 2287 1690 2291 1691
rect 2287 1685 2291 1686
rect 2303 1690 2307 1691
rect 2303 1685 2307 1686
rect 2351 1690 2355 1691
rect 2351 1685 2355 1686
rect 2391 1690 2395 1691
rect 2391 1685 2395 1686
rect 2423 1690 2427 1691
rect 2423 1685 2427 1686
rect 2479 1690 2483 1691
rect 2479 1685 2483 1686
rect 2487 1690 2491 1691
rect 2487 1685 2491 1686
rect 2543 1690 2547 1691
rect 2543 1685 2547 1686
rect 2583 1690 2587 1691
rect 2583 1685 2587 1686
rect 111 1678 115 1679
rect 111 1673 115 1674
rect 367 1678 371 1679
rect 367 1673 371 1674
rect 399 1678 403 1679
rect 399 1673 403 1674
rect 423 1678 427 1679
rect 423 1673 427 1674
rect 455 1678 459 1679
rect 455 1673 459 1674
rect 487 1678 491 1679
rect 487 1673 491 1674
rect 511 1678 515 1679
rect 511 1673 515 1674
rect 567 1678 571 1679
rect 567 1673 571 1674
rect 575 1678 579 1679
rect 575 1673 579 1674
rect 647 1678 651 1679
rect 647 1673 651 1674
rect 655 1678 659 1679
rect 655 1673 659 1674
rect 727 1678 731 1679
rect 727 1673 731 1674
rect 743 1678 747 1679
rect 743 1673 747 1674
rect 807 1678 811 1679
rect 807 1673 811 1674
rect 839 1678 843 1679
rect 839 1673 843 1674
rect 887 1678 891 1679
rect 887 1673 891 1674
rect 935 1678 939 1679
rect 935 1673 939 1674
rect 967 1678 971 1679
rect 967 1673 971 1674
rect 1031 1678 1035 1679
rect 1031 1673 1035 1674
rect 1047 1678 1051 1679
rect 1047 1673 1051 1674
rect 1127 1678 1131 1679
rect 1127 1673 1131 1674
rect 1135 1678 1139 1679
rect 1135 1673 1139 1674
rect 1223 1678 1227 1679
rect 1223 1673 1227 1674
rect 1287 1678 1291 1679
rect 1287 1673 1291 1674
rect 1327 1678 1331 1679
rect 1327 1673 1331 1674
rect 112 1658 114 1673
rect 400 1667 402 1673
rect 456 1667 458 1673
rect 512 1667 514 1673
rect 576 1667 578 1673
rect 648 1667 650 1673
rect 728 1667 730 1673
rect 808 1667 810 1673
rect 888 1667 890 1673
rect 968 1667 970 1673
rect 1048 1667 1050 1673
rect 1136 1667 1138 1673
rect 1224 1667 1226 1673
rect 1288 1667 1290 1673
rect 398 1666 404 1667
rect 398 1662 399 1666
rect 403 1662 404 1666
rect 398 1661 404 1662
rect 454 1666 460 1667
rect 454 1662 455 1666
rect 459 1662 460 1666
rect 454 1661 460 1662
rect 510 1666 516 1667
rect 510 1662 511 1666
rect 515 1662 516 1666
rect 510 1661 516 1662
rect 574 1666 580 1667
rect 574 1662 575 1666
rect 579 1662 580 1666
rect 574 1661 580 1662
rect 646 1666 652 1667
rect 646 1662 647 1666
rect 651 1662 652 1666
rect 646 1661 652 1662
rect 726 1666 732 1667
rect 726 1662 727 1666
rect 731 1662 732 1666
rect 726 1661 732 1662
rect 806 1666 812 1667
rect 806 1662 807 1666
rect 811 1662 812 1666
rect 806 1661 812 1662
rect 886 1666 892 1667
rect 886 1662 887 1666
rect 891 1662 892 1666
rect 886 1661 892 1662
rect 966 1666 972 1667
rect 966 1662 967 1666
rect 971 1662 972 1666
rect 966 1661 972 1662
rect 1046 1666 1052 1667
rect 1046 1662 1047 1666
rect 1051 1662 1052 1666
rect 1046 1661 1052 1662
rect 1134 1666 1140 1667
rect 1134 1662 1135 1666
rect 1139 1662 1140 1666
rect 1134 1661 1140 1662
rect 1222 1666 1228 1667
rect 1222 1662 1223 1666
rect 1227 1662 1228 1666
rect 1222 1661 1228 1662
rect 1286 1666 1292 1667
rect 1286 1662 1287 1666
rect 1291 1662 1292 1666
rect 1286 1661 1292 1662
rect 1328 1658 1330 1673
rect 1368 1670 1370 1685
rect 1560 1679 1562 1685
rect 1632 1679 1634 1685
rect 1712 1679 1714 1685
rect 1800 1679 1802 1685
rect 1888 1679 1890 1685
rect 1976 1679 1978 1685
rect 2064 1679 2066 1685
rect 2144 1679 2146 1685
rect 2216 1679 2218 1685
rect 2288 1679 2290 1685
rect 2352 1679 2354 1685
rect 2424 1679 2426 1685
rect 2488 1679 2490 1685
rect 2544 1679 2546 1685
rect 1558 1678 1564 1679
rect 1558 1674 1559 1678
rect 1563 1674 1564 1678
rect 1558 1673 1564 1674
rect 1630 1678 1636 1679
rect 1630 1674 1631 1678
rect 1635 1674 1636 1678
rect 1630 1673 1636 1674
rect 1710 1678 1716 1679
rect 1710 1674 1711 1678
rect 1715 1674 1716 1678
rect 1710 1673 1716 1674
rect 1798 1678 1804 1679
rect 1798 1674 1799 1678
rect 1803 1674 1804 1678
rect 1798 1673 1804 1674
rect 1886 1678 1892 1679
rect 1886 1674 1887 1678
rect 1891 1674 1892 1678
rect 1886 1673 1892 1674
rect 1974 1678 1980 1679
rect 1974 1674 1975 1678
rect 1979 1674 1980 1678
rect 1974 1673 1980 1674
rect 2062 1678 2068 1679
rect 2062 1674 2063 1678
rect 2067 1674 2068 1678
rect 2062 1673 2068 1674
rect 2142 1678 2148 1679
rect 2142 1674 2143 1678
rect 2147 1674 2148 1678
rect 2142 1673 2148 1674
rect 2214 1678 2220 1679
rect 2214 1674 2215 1678
rect 2219 1674 2220 1678
rect 2214 1673 2220 1674
rect 2286 1678 2292 1679
rect 2286 1674 2287 1678
rect 2291 1674 2292 1678
rect 2286 1673 2292 1674
rect 2350 1678 2356 1679
rect 2350 1674 2351 1678
rect 2355 1674 2356 1678
rect 2350 1673 2356 1674
rect 2422 1678 2428 1679
rect 2422 1674 2423 1678
rect 2427 1674 2428 1678
rect 2422 1673 2428 1674
rect 2486 1678 2492 1679
rect 2486 1674 2487 1678
rect 2491 1674 2492 1678
rect 2486 1673 2492 1674
rect 2542 1678 2548 1679
rect 2542 1674 2543 1678
rect 2547 1674 2548 1678
rect 2542 1673 2548 1674
rect 2584 1670 2586 1685
rect 1366 1669 1372 1670
rect 1366 1665 1367 1669
rect 1371 1665 1372 1669
rect 1366 1664 1372 1665
rect 2582 1669 2588 1670
rect 2582 1665 2583 1669
rect 2587 1665 2588 1669
rect 2582 1664 2588 1665
rect 110 1657 116 1658
rect 110 1653 111 1657
rect 115 1653 116 1657
rect 110 1652 116 1653
rect 1326 1657 1332 1658
rect 1326 1653 1327 1657
rect 1331 1653 1332 1657
rect 1326 1652 1332 1653
rect 1366 1652 1372 1653
rect 2582 1652 2588 1653
rect 1366 1648 1367 1652
rect 1371 1648 1372 1652
rect 1366 1647 1372 1648
rect 1542 1651 1548 1652
rect 1542 1647 1543 1651
rect 1547 1647 1548 1651
rect 110 1640 116 1641
rect 1326 1640 1332 1641
rect 110 1636 111 1640
rect 115 1636 116 1640
rect 110 1635 116 1636
rect 382 1639 388 1640
rect 382 1635 383 1639
rect 387 1635 388 1639
rect 112 1607 114 1635
rect 382 1634 388 1635
rect 438 1639 444 1640
rect 438 1635 439 1639
rect 443 1635 444 1639
rect 438 1634 444 1635
rect 494 1639 500 1640
rect 494 1635 495 1639
rect 499 1635 500 1639
rect 494 1634 500 1635
rect 558 1639 564 1640
rect 558 1635 559 1639
rect 563 1635 564 1639
rect 558 1634 564 1635
rect 630 1639 636 1640
rect 630 1635 631 1639
rect 635 1635 636 1639
rect 630 1634 636 1635
rect 710 1639 716 1640
rect 710 1635 711 1639
rect 715 1635 716 1639
rect 710 1634 716 1635
rect 790 1639 796 1640
rect 790 1635 791 1639
rect 795 1635 796 1639
rect 790 1634 796 1635
rect 870 1639 876 1640
rect 870 1635 871 1639
rect 875 1635 876 1639
rect 870 1634 876 1635
rect 950 1639 956 1640
rect 950 1635 951 1639
rect 955 1635 956 1639
rect 950 1634 956 1635
rect 1030 1639 1036 1640
rect 1030 1635 1031 1639
rect 1035 1635 1036 1639
rect 1030 1634 1036 1635
rect 1118 1639 1124 1640
rect 1118 1635 1119 1639
rect 1123 1635 1124 1639
rect 1118 1634 1124 1635
rect 1206 1639 1212 1640
rect 1206 1635 1207 1639
rect 1211 1635 1212 1639
rect 1206 1634 1212 1635
rect 1270 1639 1276 1640
rect 1270 1635 1271 1639
rect 1275 1635 1276 1639
rect 1326 1636 1327 1640
rect 1331 1636 1332 1640
rect 1326 1635 1332 1636
rect 1270 1634 1276 1635
rect 384 1607 386 1634
rect 440 1607 442 1634
rect 496 1607 498 1634
rect 560 1607 562 1634
rect 632 1607 634 1634
rect 712 1607 714 1634
rect 792 1607 794 1634
rect 872 1607 874 1634
rect 952 1607 954 1634
rect 1032 1607 1034 1634
rect 1120 1607 1122 1634
rect 1208 1607 1210 1634
rect 1272 1607 1274 1634
rect 1328 1607 1330 1635
rect 1368 1623 1370 1647
rect 1542 1646 1548 1647
rect 1614 1651 1620 1652
rect 1614 1647 1615 1651
rect 1619 1647 1620 1651
rect 1614 1646 1620 1647
rect 1694 1651 1700 1652
rect 1694 1647 1695 1651
rect 1699 1647 1700 1651
rect 1694 1646 1700 1647
rect 1782 1651 1788 1652
rect 1782 1647 1783 1651
rect 1787 1647 1788 1651
rect 1782 1646 1788 1647
rect 1870 1651 1876 1652
rect 1870 1647 1871 1651
rect 1875 1647 1876 1651
rect 1870 1646 1876 1647
rect 1958 1651 1964 1652
rect 1958 1647 1959 1651
rect 1963 1647 1964 1651
rect 1958 1646 1964 1647
rect 2046 1651 2052 1652
rect 2046 1647 2047 1651
rect 2051 1647 2052 1651
rect 2046 1646 2052 1647
rect 2126 1651 2132 1652
rect 2126 1647 2127 1651
rect 2131 1647 2132 1651
rect 2126 1646 2132 1647
rect 2198 1651 2204 1652
rect 2198 1647 2199 1651
rect 2203 1647 2204 1651
rect 2198 1646 2204 1647
rect 2270 1651 2276 1652
rect 2270 1647 2271 1651
rect 2275 1647 2276 1651
rect 2270 1646 2276 1647
rect 2334 1651 2340 1652
rect 2334 1647 2335 1651
rect 2339 1647 2340 1651
rect 2334 1646 2340 1647
rect 2406 1651 2412 1652
rect 2406 1647 2407 1651
rect 2411 1647 2412 1651
rect 2406 1646 2412 1647
rect 2470 1651 2476 1652
rect 2470 1647 2471 1651
rect 2475 1647 2476 1651
rect 2470 1646 2476 1647
rect 2526 1651 2532 1652
rect 2526 1647 2527 1651
rect 2531 1647 2532 1651
rect 2582 1648 2583 1652
rect 2587 1648 2588 1652
rect 2582 1647 2588 1648
rect 2526 1646 2532 1647
rect 1544 1623 1546 1646
rect 1616 1623 1618 1646
rect 1696 1623 1698 1646
rect 1784 1623 1786 1646
rect 1872 1623 1874 1646
rect 1960 1623 1962 1646
rect 2048 1623 2050 1646
rect 2128 1623 2130 1646
rect 2200 1623 2202 1646
rect 2272 1623 2274 1646
rect 2336 1623 2338 1646
rect 2408 1623 2410 1646
rect 2472 1623 2474 1646
rect 2528 1623 2530 1646
rect 2584 1623 2586 1647
rect 1367 1622 1371 1623
rect 1367 1617 1371 1618
rect 1543 1622 1547 1623
rect 1543 1617 1547 1618
rect 1575 1622 1579 1623
rect 1575 1617 1579 1618
rect 1615 1622 1619 1623
rect 1615 1617 1619 1618
rect 1631 1622 1635 1623
rect 1631 1617 1635 1618
rect 1687 1622 1691 1623
rect 1687 1617 1691 1618
rect 1695 1622 1699 1623
rect 1695 1617 1699 1618
rect 1751 1622 1755 1623
rect 1751 1617 1755 1618
rect 1783 1622 1787 1623
rect 1783 1617 1787 1618
rect 1831 1622 1835 1623
rect 1831 1617 1835 1618
rect 1871 1622 1875 1623
rect 1871 1617 1875 1618
rect 1919 1622 1923 1623
rect 1919 1617 1923 1618
rect 1959 1622 1963 1623
rect 1959 1617 1963 1618
rect 2007 1622 2011 1623
rect 2007 1617 2011 1618
rect 2047 1622 2051 1623
rect 2047 1617 2051 1618
rect 2103 1622 2107 1623
rect 2103 1617 2107 1618
rect 2127 1622 2131 1623
rect 2127 1617 2131 1618
rect 2199 1622 2203 1623
rect 2199 1617 2203 1618
rect 2207 1622 2211 1623
rect 2207 1617 2211 1618
rect 2271 1622 2275 1623
rect 2271 1617 2275 1618
rect 2319 1622 2323 1623
rect 2319 1617 2323 1618
rect 2335 1622 2339 1623
rect 2335 1617 2339 1618
rect 2407 1622 2411 1623
rect 2407 1617 2411 1618
rect 2431 1622 2435 1623
rect 2431 1617 2435 1618
rect 2471 1622 2475 1623
rect 2471 1617 2475 1618
rect 2527 1622 2531 1623
rect 2527 1617 2531 1618
rect 2583 1622 2587 1623
rect 2583 1617 2587 1618
rect 111 1606 115 1607
rect 111 1601 115 1602
rect 287 1606 291 1607
rect 287 1601 291 1602
rect 367 1606 371 1607
rect 367 1601 371 1602
rect 383 1606 387 1607
rect 383 1601 387 1602
rect 439 1606 443 1607
rect 439 1601 443 1602
rect 455 1606 459 1607
rect 455 1601 459 1602
rect 495 1606 499 1607
rect 495 1601 499 1602
rect 551 1606 555 1607
rect 551 1601 555 1602
rect 559 1606 563 1607
rect 559 1601 563 1602
rect 631 1606 635 1607
rect 631 1601 635 1602
rect 647 1606 651 1607
rect 647 1601 651 1602
rect 711 1606 715 1607
rect 711 1601 715 1602
rect 735 1606 739 1607
rect 735 1601 739 1602
rect 791 1606 795 1607
rect 791 1601 795 1602
rect 823 1606 827 1607
rect 823 1601 827 1602
rect 871 1606 875 1607
rect 871 1601 875 1602
rect 903 1606 907 1607
rect 903 1601 907 1602
rect 951 1606 955 1607
rect 951 1601 955 1602
rect 983 1606 987 1607
rect 983 1601 987 1602
rect 1031 1606 1035 1607
rect 1031 1601 1035 1602
rect 1063 1606 1067 1607
rect 1063 1601 1067 1602
rect 1119 1606 1123 1607
rect 1119 1601 1123 1602
rect 1151 1606 1155 1607
rect 1151 1601 1155 1602
rect 1207 1606 1211 1607
rect 1207 1601 1211 1602
rect 1271 1606 1275 1607
rect 1271 1601 1275 1602
rect 1327 1606 1331 1607
rect 1368 1605 1370 1617
rect 1576 1606 1578 1617
rect 1632 1606 1634 1617
rect 1688 1606 1690 1617
rect 1752 1606 1754 1617
rect 1832 1606 1834 1617
rect 1920 1606 1922 1617
rect 2008 1606 2010 1617
rect 2104 1606 2106 1617
rect 2208 1606 2210 1617
rect 2320 1606 2322 1617
rect 2432 1606 2434 1617
rect 2528 1606 2530 1617
rect 1574 1605 1580 1606
rect 1327 1601 1331 1602
rect 1366 1604 1372 1605
rect 112 1589 114 1601
rect 288 1590 290 1601
rect 368 1590 370 1601
rect 456 1590 458 1601
rect 552 1590 554 1601
rect 648 1590 650 1601
rect 736 1590 738 1601
rect 824 1590 826 1601
rect 904 1590 906 1601
rect 984 1590 986 1601
rect 1064 1590 1066 1601
rect 1152 1590 1154 1601
rect 286 1589 292 1590
rect 110 1588 116 1589
rect 110 1584 111 1588
rect 115 1584 116 1588
rect 286 1585 287 1589
rect 291 1585 292 1589
rect 286 1584 292 1585
rect 366 1589 372 1590
rect 366 1585 367 1589
rect 371 1585 372 1589
rect 366 1584 372 1585
rect 454 1589 460 1590
rect 454 1585 455 1589
rect 459 1585 460 1589
rect 454 1584 460 1585
rect 550 1589 556 1590
rect 550 1585 551 1589
rect 555 1585 556 1589
rect 550 1584 556 1585
rect 646 1589 652 1590
rect 646 1585 647 1589
rect 651 1585 652 1589
rect 646 1584 652 1585
rect 734 1589 740 1590
rect 734 1585 735 1589
rect 739 1585 740 1589
rect 734 1584 740 1585
rect 822 1589 828 1590
rect 822 1585 823 1589
rect 827 1585 828 1589
rect 822 1584 828 1585
rect 902 1589 908 1590
rect 902 1585 903 1589
rect 907 1585 908 1589
rect 902 1584 908 1585
rect 982 1589 988 1590
rect 982 1585 983 1589
rect 987 1585 988 1589
rect 982 1584 988 1585
rect 1062 1589 1068 1590
rect 1062 1585 1063 1589
rect 1067 1585 1068 1589
rect 1062 1584 1068 1585
rect 1150 1589 1156 1590
rect 1328 1589 1330 1601
rect 1366 1600 1367 1604
rect 1371 1600 1372 1604
rect 1574 1601 1575 1605
rect 1579 1601 1580 1605
rect 1574 1600 1580 1601
rect 1630 1605 1636 1606
rect 1630 1601 1631 1605
rect 1635 1601 1636 1605
rect 1630 1600 1636 1601
rect 1686 1605 1692 1606
rect 1686 1601 1687 1605
rect 1691 1601 1692 1605
rect 1686 1600 1692 1601
rect 1750 1605 1756 1606
rect 1750 1601 1751 1605
rect 1755 1601 1756 1605
rect 1750 1600 1756 1601
rect 1830 1605 1836 1606
rect 1830 1601 1831 1605
rect 1835 1601 1836 1605
rect 1830 1600 1836 1601
rect 1918 1605 1924 1606
rect 1918 1601 1919 1605
rect 1923 1601 1924 1605
rect 1918 1600 1924 1601
rect 2006 1605 2012 1606
rect 2006 1601 2007 1605
rect 2011 1601 2012 1605
rect 2006 1600 2012 1601
rect 2102 1605 2108 1606
rect 2102 1601 2103 1605
rect 2107 1601 2108 1605
rect 2102 1600 2108 1601
rect 2206 1605 2212 1606
rect 2206 1601 2207 1605
rect 2211 1601 2212 1605
rect 2206 1600 2212 1601
rect 2318 1605 2324 1606
rect 2318 1601 2319 1605
rect 2323 1601 2324 1605
rect 2318 1600 2324 1601
rect 2430 1605 2436 1606
rect 2430 1601 2431 1605
rect 2435 1601 2436 1605
rect 2430 1600 2436 1601
rect 2526 1605 2532 1606
rect 2584 1605 2586 1617
rect 2526 1601 2527 1605
rect 2531 1601 2532 1605
rect 2526 1600 2532 1601
rect 2582 1604 2588 1605
rect 2582 1600 2583 1604
rect 2587 1600 2588 1604
rect 1366 1599 1372 1600
rect 2582 1599 2588 1600
rect 1150 1585 1151 1589
rect 1155 1585 1156 1589
rect 1150 1584 1156 1585
rect 1326 1588 1332 1589
rect 1326 1584 1327 1588
rect 1331 1584 1332 1588
rect 110 1583 116 1584
rect 1326 1583 1332 1584
rect 1366 1587 1372 1588
rect 1366 1583 1367 1587
rect 1371 1583 1372 1587
rect 1366 1582 1372 1583
rect 2582 1587 2588 1588
rect 2582 1583 2583 1587
rect 2587 1583 2588 1587
rect 2582 1582 2588 1583
rect 110 1571 116 1572
rect 110 1567 111 1571
rect 115 1567 116 1571
rect 110 1566 116 1567
rect 1326 1571 1332 1572
rect 1326 1567 1327 1571
rect 1331 1567 1332 1571
rect 1326 1566 1332 1567
rect 112 1551 114 1566
rect 302 1562 308 1563
rect 302 1558 303 1562
rect 307 1558 308 1562
rect 302 1557 308 1558
rect 382 1562 388 1563
rect 382 1558 383 1562
rect 387 1558 388 1562
rect 382 1557 388 1558
rect 470 1562 476 1563
rect 470 1558 471 1562
rect 475 1558 476 1562
rect 470 1557 476 1558
rect 566 1562 572 1563
rect 566 1558 567 1562
rect 571 1558 572 1562
rect 566 1557 572 1558
rect 662 1562 668 1563
rect 662 1558 663 1562
rect 667 1558 668 1562
rect 662 1557 668 1558
rect 750 1562 756 1563
rect 750 1558 751 1562
rect 755 1558 756 1562
rect 750 1557 756 1558
rect 838 1562 844 1563
rect 838 1558 839 1562
rect 843 1558 844 1562
rect 838 1557 844 1558
rect 918 1562 924 1563
rect 918 1558 919 1562
rect 923 1558 924 1562
rect 918 1557 924 1558
rect 998 1562 1004 1563
rect 998 1558 999 1562
rect 1003 1558 1004 1562
rect 998 1557 1004 1558
rect 1078 1562 1084 1563
rect 1078 1558 1079 1562
rect 1083 1558 1084 1562
rect 1078 1557 1084 1558
rect 1166 1562 1172 1563
rect 1166 1558 1167 1562
rect 1171 1558 1172 1562
rect 1166 1557 1172 1558
rect 304 1551 306 1557
rect 384 1551 386 1557
rect 472 1551 474 1557
rect 568 1551 570 1557
rect 664 1551 666 1557
rect 752 1551 754 1557
rect 840 1551 842 1557
rect 920 1551 922 1557
rect 1000 1551 1002 1557
rect 1080 1551 1082 1557
rect 1168 1551 1170 1557
rect 1328 1551 1330 1566
rect 1368 1563 1370 1582
rect 1590 1578 1596 1579
rect 1590 1574 1591 1578
rect 1595 1574 1596 1578
rect 1590 1573 1596 1574
rect 1646 1578 1652 1579
rect 1646 1574 1647 1578
rect 1651 1574 1652 1578
rect 1646 1573 1652 1574
rect 1702 1578 1708 1579
rect 1702 1574 1703 1578
rect 1707 1574 1708 1578
rect 1702 1573 1708 1574
rect 1766 1578 1772 1579
rect 1766 1574 1767 1578
rect 1771 1574 1772 1578
rect 1766 1573 1772 1574
rect 1846 1578 1852 1579
rect 1846 1574 1847 1578
rect 1851 1574 1852 1578
rect 1846 1573 1852 1574
rect 1934 1578 1940 1579
rect 1934 1574 1935 1578
rect 1939 1574 1940 1578
rect 1934 1573 1940 1574
rect 2022 1578 2028 1579
rect 2022 1574 2023 1578
rect 2027 1574 2028 1578
rect 2022 1573 2028 1574
rect 2118 1578 2124 1579
rect 2118 1574 2119 1578
rect 2123 1574 2124 1578
rect 2118 1573 2124 1574
rect 2222 1578 2228 1579
rect 2222 1574 2223 1578
rect 2227 1574 2228 1578
rect 2222 1573 2228 1574
rect 2334 1578 2340 1579
rect 2334 1574 2335 1578
rect 2339 1574 2340 1578
rect 2334 1573 2340 1574
rect 2446 1578 2452 1579
rect 2446 1574 2447 1578
rect 2451 1574 2452 1578
rect 2446 1573 2452 1574
rect 2542 1578 2548 1579
rect 2542 1574 2543 1578
rect 2547 1574 2548 1578
rect 2542 1573 2548 1574
rect 1592 1563 1594 1573
rect 1648 1563 1650 1573
rect 1704 1563 1706 1573
rect 1768 1563 1770 1573
rect 1848 1563 1850 1573
rect 1936 1563 1938 1573
rect 2024 1563 2026 1573
rect 2120 1563 2122 1573
rect 2224 1563 2226 1573
rect 2336 1563 2338 1573
rect 2448 1563 2450 1573
rect 2544 1563 2546 1573
rect 2584 1563 2586 1582
rect 1367 1562 1371 1563
rect 1367 1557 1371 1558
rect 1591 1562 1595 1563
rect 1591 1557 1595 1558
rect 1647 1562 1651 1563
rect 1647 1557 1651 1558
rect 1679 1562 1683 1563
rect 1679 1557 1683 1558
rect 1703 1562 1707 1563
rect 1703 1557 1707 1558
rect 1735 1562 1739 1563
rect 1735 1557 1739 1558
rect 1767 1562 1771 1563
rect 1767 1557 1771 1558
rect 1791 1562 1795 1563
rect 1791 1557 1795 1558
rect 1847 1562 1851 1563
rect 1847 1557 1851 1558
rect 1855 1562 1859 1563
rect 1855 1557 1859 1558
rect 1927 1562 1931 1563
rect 1927 1557 1931 1558
rect 1935 1562 1939 1563
rect 1935 1557 1939 1558
rect 2007 1562 2011 1563
rect 2007 1557 2011 1558
rect 2023 1562 2027 1563
rect 2023 1557 2027 1558
rect 2087 1562 2091 1563
rect 2087 1557 2091 1558
rect 2119 1562 2123 1563
rect 2119 1557 2123 1558
rect 2167 1562 2171 1563
rect 2167 1557 2171 1558
rect 2223 1562 2227 1563
rect 2223 1557 2227 1558
rect 2247 1562 2251 1563
rect 2247 1557 2251 1558
rect 2327 1562 2331 1563
rect 2327 1557 2331 1558
rect 2335 1562 2339 1563
rect 2335 1557 2339 1558
rect 2407 1562 2411 1563
rect 2407 1557 2411 1558
rect 2447 1562 2451 1563
rect 2447 1557 2451 1558
rect 2487 1562 2491 1563
rect 2487 1557 2491 1558
rect 2543 1562 2547 1563
rect 2543 1557 2547 1558
rect 2583 1562 2587 1563
rect 2583 1557 2587 1558
rect 111 1550 115 1551
rect 111 1545 115 1546
rect 279 1550 283 1551
rect 279 1545 283 1546
rect 303 1550 307 1551
rect 303 1545 307 1546
rect 335 1550 339 1551
rect 335 1545 339 1546
rect 383 1550 387 1551
rect 383 1545 387 1546
rect 399 1550 403 1551
rect 399 1545 403 1546
rect 471 1550 475 1551
rect 471 1545 475 1546
rect 543 1550 547 1551
rect 543 1545 547 1546
rect 567 1550 571 1551
rect 567 1545 571 1546
rect 615 1550 619 1551
rect 615 1545 619 1546
rect 663 1550 667 1551
rect 663 1545 667 1546
rect 687 1550 691 1551
rect 687 1545 691 1546
rect 751 1550 755 1551
rect 751 1545 755 1546
rect 759 1550 763 1551
rect 759 1545 763 1546
rect 831 1550 835 1551
rect 831 1545 835 1546
rect 839 1550 843 1551
rect 839 1545 843 1546
rect 903 1550 907 1551
rect 903 1545 907 1546
rect 919 1550 923 1551
rect 919 1545 923 1546
rect 975 1550 979 1551
rect 975 1545 979 1546
rect 999 1550 1003 1551
rect 999 1545 1003 1546
rect 1055 1550 1059 1551
rect 1055 1545 1059 1546
rect 1079 1550 1083 1551
rect 1079 1545 1083 1546
rect 1167 1550 1171 1551
rect 1167 1545 1171 1546
rect 1327 1550 1331 1551
rect 1327 1545 1331 1546
rect 112 1530 114 1545
rect 280 1539 282 1545
rect 336 1539 338 1545
rect 400 1539 402 1545
rect 472 1539 474 1545
rect 544 1539 546 1545
rect 616 1539 618 1545
rect 688 1539 690 1545
rect 760 1539 762 1545
rect 832 1539 834 1545
rect 904 1539 906 1545
rect 976 1539 978 1545
rect 1056 1539 1058 1545
rect 278 1538 284 1539
rect 278 1534 279 1538
rect 283 1534 284 1538
rect 278 1533 284 1534
rect 334 1538 340 1539
rect 334 1534 335 1538
rect 339 1534 340 1538
rect 334 1533 340 1534
rect 398 1538 404 1539
rect 398 1534 399 1538
rect 403 1534 404 1538
rect 398 1533 404 1534
rect 470 1538 476 1539
rect 470 1534 471 1538
rect 475 1534 476 1538
rect 470 1533 476 1534
rect 542 1538 548 1539
rect 542 1534 543 1538
rect 547 1534 548 1538
rect 542 1533 548 1534
rect 614 1538 620 1539
rect 614 1534 615 1538
rect 619 1534 620 1538
rect 614 1533 620 1534
rect 686 1538 692 1539
rect 686 1534 687 1538
rect 691 1534 692 1538
rect 686 1533 692 1534
rect 758 1538 764 1539
rect 758 1534 759 1538
rect 763 1534 764 1538
rect 758 1533 764 1534
rect 830 1538 836 1539
rect 830 1534 831 1538
rect 835 1534 836 1538
rect 830 1533 836 1534
rect 902 1538 908 1539
rect 902 1534 903 1538
rect 907 1534 908 1538
rect 902 1533 908 1534
rect 974 1538 980 1539
rect 974 1534 975 1538
rect 979 1534 980 1538
rect 974 1533 980 1534
rect 1054 1538 1060 1539
rect 1054 1534 1055 1538
rect 1059 1534 1060 1538
rect 1054 1533 1060 1534
rect 1328 1530 1330 1545
rect 1368 1542 1370 1557
rect 1680 1551 1682 1557
rect 1736 1551 1738 1557
rect 1792 1551 1794 1557
rect 1856 1551 1858 1557
rect 1928 1551 1930 1557
rect 2008 1551 2010 1557
rect 2088 1551 2090 1557
rect 2168 1551 2170 1557
rect 2248 1551 2250 1557
rect 2328 1551 2330 1557
rect 2408 1551 2410 1557
rect 2488 1551 2490 1557
rect 2544 1551 2546 1557
rect 1678 1550 1684 1551
rect 1678 1546 1679 1550
rect 1683 1546 1684 1550
rect 1678 1545 1684 1546
rect 1734 1550 1740 1551
rect 1734 1546 1735 1550
rect 1739 1546 1740 1550
rect 1734 1545 1740 1546
rect 1790 1550 1796 1551
rect 1790 1546 1791 1550
rect 1795 1546 1796 1550
rect 1790 1545 1796 1546
rect 1854 1550 1860 1551
rect 1854 1546 1855 1550
rect 1859 1546 1860 1550
rect 1854 1545 1860 1546
rect 1926 1550 1932 1551
rect 1926 1546 1927 1550
rect 1931 1546 1932 1550
rect 1926 1545 1932 1546
rect 2006 1550 2012 1551
rect 2006 1546 2007 1550
rect 2011 1546 2012 1550
rect 2006 1545 2012 1546
rect 2086 1550 2092 1551
rect 2086 1546 2087 1550
rect 2091 1546 2092 1550
rect 2086 1545 2092 1546
rect 2166 1550 2172 1551
rect 2166 1546 2167 1550
rect 2171 1546 2172 1550
rect 2166 1545 2172 1546
rect 2246 1550 2252 1551
rect 2246 1546 2247 1550
rect 2251 1546 2252 1550
rect 2246 1545 2252 1546
rect 2326 1550 2332 1551
rect 2326 1546 2327 1550
rect 2331 1546 2332 1550
rect 2326 1545 2332 1546
rect 2406 1550 2412 1551
rect 2406 1546 2407 1550
rect 2411 1546 2412 1550
rect 2406 1545 2412 1546
rect 2486 1550 2492 1551
rect 2486 1546 2487 1550
rect 2491 1546 2492 1550
rect 2486 1545 2492 1546
rect 2542 1550 2548 1551
rect 2542 1546 2543 1550
rect 2547 1546 2548 1550
rect 2542 1545 2548 1546
rect 2584 1542 2586 1557
rect 1366 1541 1372 1542
rect 1366 1537 1367 1541
rect 1371 1537 1372 1541
rect 1366 1536 1372 1537
rect 2582 1541 2588 1542
rect 2582 1537 2583 1541
rect 2587 1537 2588 1541
rect 2582 1536 2588 1537
rect 110 1529 116 1530
rect 110 1525 111 1529
rect 115 1525 116 1529
rect 110 1524 116 1525
rect 1326 1529 1332 1530
rect 1326 1525 1327 1529
rect 1331 1525 1332 1529
rect 1326 1524 1332 1525
rect 1366 1524 1372 1525
rect 2582 1524 2588 1525
rect 1366 1520 1367 1524
rect 1371 1520 1372 1524
rect 1366 1519 1372 1520
rect 1662 1523 1668 1524
rect 1662 1519 1663 1523
rect 1667 1519 1668 1523
rect 110 1512 116 1513
rect 1326 1512 1332 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 110 1507 116 1508
rect 262 1511 268 1512
rect 262 1507 263 1511
rect 267 1507 268 1511
rect 112 1491 114 1507
rect 262 1506 268 1507
rect 318 1511 324 1512
rect 318 1507 319 1511
rect 323 1507 324 1511
rect 318 1506 324 1507
rect 382 1511 388 1512
rect 382 1507 383 1511
rect 387 1507 388 1511
rect 382 1506 388 1507
rect 454 1511 460 1512
rect 454 1507 455 1511
rect 459 1507 460 1511
rect 454 1506 460 1507
rect 526 1511 532 1512
rect 526 1507 527 1511
rect 531 1507 532 1511
rect 526 1506 532 1507
rect 598 1511 604 1512
rect 598 1507 599 1511
rect 603 1507 604 1511
rect 598 1506 604 1507
rect 670 1511 676 1512
rect 670 1507 671 1511
rect 675 1507 676 1511
rect 670 1506 676 1507
rect 742 1511 748 1512
rect 742 1507 743 1511
rect 747 1507 748 1511
rect 742 1506 748 1507
rect 814 1511 820 1512
rect 814 1507 815 1511
rect 819 1507 820 1511
rect 814 1506 820 1507
rect 886 1511 892 1512
rect 886 1507 887 1511
rect 891 1507 892 1511
rect 886 1506 892 1507
rect 958 1511 964 1512
rect 958 1507 959 1511
rect 963 1507 964 1511
rect 958 1506 964 1507
rect 1038 1511 1044 1512
rect 1038 1507 1039 1511
rect 1043 1507 1044 1511
rect 1326 1508 1327 1512
rect 1331 1508 1332 1512
rect 1326 1507 1332 1508
rect 1038 1506 1044 1507
rect 264 1491 266 1506
rect 320 1491 322 1506
rect 384 1491 386 1506
rect 456 1491 458 1506
rect 528 1491 530 1506
rect 600 1491 602 1506
rect 672 1491 674 1506
rect 744 1491 746 1506
rect 816 1491 818 1506
rect 888 1491 890 1506
rect 960 1491 962 1506
rect 1040 1491 1042 1506
rect 1328 1491 1330 1507
rect 1368 1499 1370 1519
rect 1662 1518 1668 1519
rect 1718 1523 1724 1524
rect 1718 1519 1719 1523
rect 1723 1519 1724 1523
rect 1718 1518 1724 1519
rect 1774 1523 1780 1524
rect 1774 1519 1775 1523
rect 1779 1519 1780 1523
rect 1774 1518 1780 1519
rect 1838 1523 1844 1524
rect 1838 1519 1839 1523
rect 1843 1519 1844 1523
rect 1838 1518 1844 1519
rect 1910 1523 1916 1524
rect 1910 1519 1911 1523
rect 1915 1519 1916 1523
rect 1910 1518 1916 1519
rect 1990 1523 1996 1524
rect 1990 1519 1991 1523
rect 1995 1519 1996 1523
rect 1990 1518 1996 1519
rect 2070 1523 2076 1524
rect 2070 1519 2071 1523
rect 2075 1519 2076 1523
rect 2070 1518 2076 1519
rect 2150 1523 2156 1524
rect 2150 1519 2151 1523
rect 2155 1519 2156 1523
rect 2150 1518 2156 1519
rect 2230 1523 2236 1524
rect 2230 1519 2231 1523
rect 2235 1519 2236 1523
rect 2230 1518 2236 1519
rect 2310 1523 2316 1524
rect 2310 1519 2311 1523
rect 2315 1519 2316 1523
rect 2310 1518 2316 1519
rect 2390 1523 2396 1524
rect 2390 1519 2391 1523
rect 2395 1519 2396 1523
rect 2390 1518 2396 1519
rect 2470 1523 2476 1524
rect 2470 1519 2471 1523
rect 2475 1519 2476 1523
rect 2470 1518 2476 1519
rect 2526 1523 2532 1524
rect 2526 1519 2527 1523
rect 2531 1519 2532 1523
rect 2582 1520 2583 1524
rect 2587 1520 2588 1524
rect 2582 1519 2588 1520
rect 2526 1518 2532 1519
rect 1664 1499 1666 1518
rect 1720 1499 1722 1518
rect 1776 1499 1778 1518
rect 1840 1499 1842 1518
rect 1912 1499 1914 1518
rect 1992 1499 1994 1518
rect 2072 1499 2074 1518
rect 2152 1499 2154 1518
rect 2232 1499 2234 1518
rect 2312 1499 2314 1518
rect 2392 1499 2394 1518
rect 2472 1499 2474 1518
rect 2528 1499 2530 1518
rect 2584 1499 2586 1519
rect 1367 1498 1371 1499
rect 1367 1493 1371 1494
rect 1519 1498 1523 1499
rect 1519 1493 1523 1494
rect 1575 1498 1579 1499
rect 1575 1493 1579 1494
rect 1647 1498 1651 1499
rect 1647 1493 1651 1494
rect 1663 1498 1667 1499
rect 1663 1493 1667 1494
rect 1719 1498 1723 1499
rect 1719 1493 1723 1494
rect 1727 1498 1731 1499
rect 1727 1493 1731 1494
rect 1775 1498 1779 1499
rect 1775 1493 1779 1494
rect 1807 1498 1811 1499
rect 1807 1493 1811 1494
rect 1839 1498 1843 1499
rect 1839 1493 1843 1494
rect 1895 1498 1899 1499
rect 1895 1493 1899 1494
rect 1911 1498 1915 1499
rect 1911 1493 1915 1494
rect 1983 1498 1987 1499
rect 1983 1493 1987 1494
rect 1991 1498 1995 1499
rect 1991 1493 1995 1494
rect 2071 1498 2075 1499
rect 2071 1493 2075 1494
rect 2151 1498 2155 1499
rect 2151 1493 2155 1494
rect 2231 1498 2235 1499
rect 2231 1493 2235 1494
rect 2311 1498 2315 1499
rect 2311 1493 2315 1494
rect 2391 1498 2395 1499
rect 2391 1493 2395 1494
rect 2471 1498 2475 1499
rect 2471 1493 2475 1494
rect 2527 1498 2531 1499
rect 2527 1493 2531 1494
rect 2583 1498 2587 1499
rect 2583 1493 2587 1494
rect 111 1490 115 1491
rect 111 1485 115 1486
rect 199 1490 203 1491
rect 199 1485 203 1486
rect 263 1490 267 1491
rect 263 1485 267 1486
rect 287 1490 291 1491
rect 287 1485 291 1486
rect 319 1490 323 1491
rect 319 1485 323 1486
rect 383 1490 387 1491
rect 383 1485 387 1486
rect 455 1490 459 1491
rect 455 1485 459 1486
rect 487 1490 491 1491
rect 487 1485 491 1486
rect 527 1490 531 1491
rect 527 1485 531 1486
rect 583 1490 587 1491
rect 583 1485 587 1486
rect 599 1490 603 1491
rect 599 1485 603 1486
rect 671 1490 675 1491
rect 671 1485 675 1486
rect 679 1490 683 1491
rect 679 1485 683 1486
rect 743 1490 747 1491
rect 743 1485 747 1486
rect 775 1490 779 1491
rect 775 1485 779 1486
rect 815 1490 819 1491
rect 815 1485 819 1486
rect 863 1490 867 1491
rect 863 1485 867 1486
rect 887 1490 891 1491
rect 887 1485 891 1486
rect 951 1490 955 1491
rect 951 1485 955 1486
rect 959 1490 963 1491
rect 959 1485 963 1486
rect 1039 1490 1043 1491
rect 1039 1485 1043 1486
rect 1135 1490 1139 1491
rect 1135 1485 1139 1486
rect 1327 1490 1331 1491
rect 1327 1485 1331 1486
rect 112 1473 114 1485
rect 200 1474 202 1485
rect 288 1474 290 1485
rect 384 1474 386 1485
rect 488 1474 490 1485
rect 584 1474 586 1485
rect 680 1474 682 1485
rect 776 1474 778 1485
rect 864 1474 866 1485
rect 952 1474 954 1485
rect 1040 1474 1042 1485
rect 1136 1474 1138 1485
rect 198 1473 204 1474
rect 110 1472 116 1473
rect 110 1468 111 1472
rect 115 1468 116 1472
rect 198 1469 199 1473
rect 203 1469 204 1473
rect 198 1468 204 1469
rect 286 1473 292 1474
rect 286 1469 287 1473
rect 291 1469 292 1473
rect 286 1468 292 1469
rect 382 1473 388 1474
rect 382 1469 383 1473
rect 387 1469 388 1473
rect 382 1468 388 1469
rect 486 1473 492 1474
rect 486 1469 487 1473
rect 491 1469 492 1473
rect 486 1468 492 1469
rect 582 1473 588 1474
rect 582 1469 583 1473
rect 587 1469 588 1473
rect 582 1468 588 1469
rect 678 1473 684 1474
rect 678 1469 679 1473
rect 683 1469 684 1473
rect 678 1468 684 1469
rect 774 1473 780 1474
rect 774 1469 775 1473
rect 779 1469 780 1473
rect 774 1468 780 1469
rect 862 1473 868 1474
rect 862 1469 863 1473
rect 867 1469 868 1473
rect 862 1468 868 1469
rect 950 1473 956 1474
rect 950 1469 951 1473
rect 955 1469 956 1473
rect 950 1468 956 1469
rect 1038 1473 1044 1474
rect 1038 1469 1039 1473
rect 1043 1469 1044 1473
rect 1038 1468 1044 1469
rect 1134 1473 1140 1474
rect 1328 1473 1330 1485
rect 1368 1481 1370 1493
rect 1520 1482 1522 1493
rect 1576 1482 1578 1493
rect 1648 1482 1650 1493
rect 1728 1482 1730 1493
rect 1808 1482 1810 1493
rect 1896 1482 1898 1493
rect 1984 1482 1986 1493
rect 2072 1482 2074 1493
rect 2152 1482 2154 1493
rect 2232 1482 2234 1493
rect 2312 1482 2314 1493
rect 2392 1482 2394 1493
rect 2472 1482 2474 1493
rect 2528 1482 2530 1493
rect 1518 1481 1524 1482
rect 1366 1480 1372 1481
rect 1366 1476 1367 1480
rect 1371 1476 1372 1480
rect 1518 1477 1519 1481
rect 1523 1477 1524 1481
rect 1518 1476 1524 1477
rect 1574 1481 1580 1482
rect 1574 1477 1575 1481
rect 1579 1477 1580 1481
rect 1574 1476 1580 1477
rect 1646 1481 1652 1482
rect 1646 1477 1647 1481
rect 1651 1477 1652 1481
rect 1646 1476 1652 1477
rect 1726 1481 1732 1482
rect 1726 1477 1727 1481
rect 1731 1477 1732 1481
rect 1726 1476 1732 1477
rect 1806 1481 1812 1482
rect 1806 1477 1807 1481
rect 1811 1477 1812 1481
rect 1806 1476 1812 1477
rect 1894 1481 1900 1482
rect 1894 1477 1895 1481
rect 1899 1477 1900 1481
rect 1894 1476 1900 1477
rect 1982 1481 1988 1482
rect 1982 1477 1983 1481
rect 1987 1477 1988 1481
rect 1982 1476 1988 1477
rect 2070 1481 2076 1482
rect 2070 1477 2071 1481
rect 2075 1477 2076 1481
rect 2070 1476 2076 1477
rect 2150 1481 2156 1482
rect 2150 1477 2151 1481
rect 2155 1477 2156 1481
rect 2150 1476 2156 1477
rect 2230 1481 2236 1482
rect 2230 1477 2231 1481
rect 2235 1477 2236 1481
rect 2230 1476 2236 1477
rect 2310 1481 2316 1482
rect 2310 1477 2311 1481
rect 2315 1477 2316 1481
rect 2310 1476 2316 1477
rect 2390 1481 2396 1482
rect 2390 1477 2391 1481
rect 2395 1477 2396 1481
rect 2390 1476 2396 1477
rect 2470 1481 2476 1482
rect 2470 1477 2471 1481
rect 2475 1477 2476 1481
rect 2470 1476 2476 1477
rect 2526 1481 2532 1482
rect 2584 1481 2586 1493
rect 2526 1477 2527 1481
rect 2531 1477 2532 1481
rect 2526 1476 2532 1477
rect 2582 1480 2588 1481
rect 2582 1476 2583 1480
rect 2587 1476 2588 1480
rect 1366 1475 1372 1476
rect 2582 1475 2588 1476
rect 1134 1469 1135 1473
rect 1139 1469 1140 1473
rect 1134 1468 1140 1469
rect 1326 1472 1332 1473
rect 1326 1468 1327 1472
rect 1331 1468 1332 1472
rect 110 1467 116 1468
rect 1326 1467 1332 1468
rect 1366 1463 1372 1464
rect 1366 1459 1367 1463
rect 1371 1459 1372 1463
rect 1366 1458 1372 1459
rect 2582 1463 2588 1464
rect 2582 1459 2583 1463
rect 2587 1459 2588 1463
rect 2582 1458 2588 1459
rect 110 1455 116 1456
rect 110 1451 111 1455
rect 115 1451 116 1455
rect 110 1450 116 1451
rect 1326 1455 1332 1456
rect 1326 1451 1327 1455
rect 1331 1451 1332 1455
rect 1326 1450 1332 1451
rect 112 1431 114 1450
rect 214 1446 220 1447
rect 214 1442 215 1446
rect 219 1442 220 1446
rect 214 1441 220 1442
rect 302 1446 308 1447
rect 302 1442 303 1446
rect 307 1442 308 1446
rect 302 1441 308 1442
rect 398 1446 404 1447
rect 398 1442 399 1446
rect 403 1442 404 1446
rect 398 1441 404 1442
rect 502 1446 508 1447
rect 502 1442 503 1446
rect 507 1442 508 1446
rect 502 1441 508 1442
rect 598 1446 604 1447
rect 598 1442 599 1446
rect 603 1442 604 1446
rect 598 1441 604 1442
rect 694 1446 700 1447
rect 694 1442 695 1446
rect 699 1442 700 1446
rect 694 1441 700 1442
rect 790 1446 796 1447
rect 790 1442 791 1446
rect 795 1442 796 1446
rect 790 1441 796 1442
rect 878 1446 884 1447
rect 878 1442 879 1446
rect 883 1442 884 1446
rect 878 1441 884 1442
rect 966 1446 972 1447
rect 966 1442 967 1446
rect 971 1442 972 1446
rect 966 1441 972 1442
rect 1054 1446 1060 1447
rect 1054 1442 1055 1446
rect 1059 1442 1060 1446
rect 1054 1441 1060 1442
rect 1150 1446 1156 1447
rect 1150 1442 1151 1446
rect 1155 1442 1156 1446
rect 1150 1441 1156 1442
rect 216 1431 218 1441
rect 304 1431 306 1441
rect 400 1431 402 1441
rect 504 1431 506 1441
rect 600 1431 602 1441
rect 696 1431 698 1441
rect 792 1431 794 1441
rect 880 1431 882 1441
rect 968 1431 970 1441
rect 1056 1431 1058 1441
rect 1152 1431 1154 1441
rect 1328 1431 1330 1450
rect 1368 1435 1370 1458
rect 1534 1454 1540 1455
rect 1534 1450 1535 1454
rect 1539 1450 1540 1454
rect 1534 1449 1540 1450
rect 1590 1454 1596 1455
rect 1590 1450 1591 1454
rect 1595 1450 1596 1454
rect 1590 1449 1596 1450
rect 1662 1454 1668 1455
rect 1662 1450 1663 1454
rect 1667 1450 1668 1454
rect 1662 1449 1668 1450
rect 1742 1454 1748 1455
rect 1742 1450 1743 1454
rect 1747 1450 1748 1454
rect 1742 1449 1748 1450
rect 1822 1454 1828 1455
rect 1822 1450 1823 1454
rect 1827 1450 1828 1454
rect 1822 1449 1828 1450
rect 1910 1454 1916 1455
rect 1910 1450 1911 1454
rect 1915 1450 1916 1454
rect 1910 1449 1916 1450
rect 1998 1454 2004 1455
rect 1998 1450 1999 1454
rect 2003 1450 2004 1454
rect 1998 1449 2004 1450
rect 2086 1454 2092 1455
rect 2086 1450 2087 1454
rect 2091 1450 2092 1454
rect 2086 1449 2092 1450
rect 2166 1454 2172 1455
rect 2166 1450 2167 1454
rect 2171 1450 2172 1454
rect 2166 1449 2172 1450
rect 2246 1454 2252 1455
rect 2246 1450 2247 1454
rect 2251 1450 2252 1454
rect 2246 1449 2252 1450
rect 2326 1454 2332 1455
rect 2326 1450 2327 1454
rect 2331 1450 2332 1454
rect 2326 1449 2332 1450
rect 2406 1454 2412 1455
rect 2406 1450 2407 1454
rect 2411 1450 2412 1454
rect 2406 1449 2412 1450
rect 2486 1454 2492 1455
rect 2486 1450 2487 1454
rect 2491 1450 2492 1454
rect 2486 1449 2492 1450
rect 2542 1454 2548 1455
rect 2542 1450 2543 1454
rect 2547 1450 2548 1454
rect 2542 1449 2548 1450
rect 1536 1435 1538 1449
rect 1592 1435 1594 1449
rect 1664 1435 1666 1449
rect 1744 1435 1746 1449
rect 1824 1435 1826 1449
rect 1912 1435 1914 1449
rect 2000 1435 2002 1449
rect 2088 1435 2090 1449
rect 2168 1435 2170 1449
rect 2248 1435 2250 1449
rect 2328 1435 2330 1449
rect 2408 1435 2410 1449
rect 2488 1435 2490 1449
rect 2544 1435 2546 1449
rect 2584 1435 2586 1458
rect 1367 1434 1371 1435
rect 111 1430 115 1431
rect 111 1425 115 1426
rect 159 1430 163 1431
rect 159 1425 163 1426
rect 215 1430 219 1431
rect 215 1425 219 1426
rect 247 1430 251 1431
rect 247 1425 251 1426
rect 303 1430 307 1431
rect 303 1425 307 1426
rect 343 1430 347 1431
rect 343 1425 347 1426
rect 399 1430 403 1431
rect 399 1425 403 1426
rect 447 1430 451 1431
rect 447 1425 451 1426
rect 503 1430 507 1431
rect 503 1425 507 1426
rect 551 1430 555 1431
rect 551 1425 555 1426
rect 599 1430 603 1431
rect 599 1425 603 1426
rect 663 1430 667 1431
rect 663 1425 667 1426
rect 695 1430 699 1431
rect 695 1425 699 1426
rect 767 1430 771 1431
rect 767 1425 771 1426
rect 791 1430 795 1431
rect 791 1425 795 1426
rect 879 1430 883 1431
rect 879 1425 883 1426
rect 967 1430 971 1431
rect 967 1425 971 1426
rect 991 1430 995 1431
rect 991 1425 995 1426
rect 1055 1430 1059 1431
rect 1055 1425 1059 1426
rect 1103 1430 1107 1431
rect 1103 1425 1107 1426
rect 1151 1430 1155 1431
rect 1151 1425 1155 1426
rect 1215 1430 1219 1431
rect 1215 1425 1219 1426
rect 1327 1430 1331 1431
rect 1367 1429 1371 1430
rect 1415 1434 1419 1435
rect 1415 1429 1419 1430
rect 1471 1434 1475 1435
rect 1471 1429 1475 1430
rect 1535 1434 1539 1435
rect 1535 1429 1539 1430
rect 1591 1434 1595 1435
rect 1591 1429 1595 1430
rect 1623 1434 1627 1435
rect 1623 1429 1627 1430
rect 1663 1434 1667 1435
rect 1663 1429 1667 1430
rect 1719 1434 1723 1435
rect 1719 1429 1723 1430
rect 1743 1434 1747 1435
rect 1743 1429 1747 1430
rect 1823 1434 1827 1435
rect 1823 1429 1827 1430
rect 1911 1434 1915 1435
rect 1911 1429 1915 1430
rect 1927 1434 1931 1435
rect 1927 1429 1931 1430
rect 1999 1434 2003 1435
rect 1999 1429 2003 1430
rect 2023 1434 2027 1435
rect 2023 1429 2027 1430
rect 2087 1434 2091 1435
rect 2087 1429 2091 1430
rect 2119 1434 2123 1435
rect 2119 1429 2123 1430
rect 2167 1434 2171 1435
rect 2167 1429 2171 1430
rect 2215 1434 2219 1435
rect 2215 1429 2219 1430
rect 2247 1434 2251 1435
rect 2247 1429 2251 1430
rect 2303 1434 2307 1435
rect 2303 1429 2307 1430
rect 2327 1434 2331 1435
rect 2327 1429 2331 1430
rect 2391 1434 2395 1435
rect 2391 1429 2395 1430
rect 2407 1434 2411 1435
rect 2407 1429 2411 1430
rect 2479 1434 2483 1435
rect 2479 1429 2483 1430
rect 2487 1434 2491 1435
rect 2487 1429 2491 1430
rect 2543 1434 2547 1435
rect 2543 1429 2547 1430
rect 2583 1434 2587 1435
rect 2583 1429 2587 1430
rect 1327 1425 1331 1426
rect 112 1410 114 1425
rect 160 1419 162 1425
rect 248 1419 250 1425
rect 344 1419 346 1425
rect 448 1419 450 1425
rect 552 1419 554 1425
rect 664 1419 666 1425
rect 768 1419 770 1425
rect 880 1419 882 1425
rect 992 1419 994 1425
rect 1104 1419 1106 1425
rect 1216 1419 1218 1425
rect 158 1418 164 1419
rect 158 1414 159 1418
rect 163 1414 164 1418
rect 158 1413 164 1414
rect 246 1418 252 1419
rect 246 1414 247 1418
rect 251 1414 252 1418
rect 246 1413 252 1414
rect 342 1418 348 1419
rect 342 1414 343 1418
rect 347 1414 348 1418
rect 342 1413 348 1414
rect 446 1418 452 1419
rect 446 1414 447 1418
rect 451 1414 452 1418
rect 446 1413 452 1414
rect 550 1418 556 1419
rect 550 1414 551 1418
rect 555 1414 556 1418
rect 550 1413 556 1414
rect 662 1418 668 1419
rect 662 1414 663 1418
rect 667 1414 668 1418
rect 662 1413 668 1414
rect 766 1418 772 1419
rect 766 1414 767 1418
rect 771 1414 772 1418
rect 766 1413 772 1414
rect 878 1418 884 1419
rect 878 1414 879 1418
rect 883 1414 884 1418
rect 878 1413 884 1414
rect 990 1418 996 1419
rect 990 1414 991 1418
rect 995 1414 996 1418
rect 990 1413 996 1414
rect 1102 1418 1108 1419
rect 1102 1414 1103 1418
rect 1107 1414 1108 1418
rect 1102 1413 1108 1414
rect 1214 1418 1220 1419
rect 1214 1414 1215 1418
rect 1219 1414 1220 1418
rect 1214 1413 1220 1414
rect 1328 1410 1330 1425
rect 1368 1414 1370 1429
rect 1416 1423 1418 1429
rect 1472 1423 1474 1429
rect 1536 1423 1538 1429
rect 1624 1423 1626 1429
rect 1720 1423 1722 1429
rect 1824 1423 1826 1429
rect 1928 1423 1930 1429
rect 2024 1423 2026 1429
rect 2120 1423 2122 1429
rect 2216 1423 2218 1429
rect 2304 1423 2306 1429
rect 2392 1423 2394 1429
rect 2480 1423 2482 1429
rect 2544 1423 2546 1429
rect 1414 1422 1420 1423
rect 1414 1418 1415 1422
rect 1419 1418 1420 1422
rect 1414 1417 1420 1418
rect 1470 1422 1476 1423
rect 1470 1418 1471 1422
rect 1475 1418 1476 1422
rect 1470 1417 1476 1418
rect 1534 1422 1540 1423
rect 1534 1418 1535 1422
rect 1539 1418 1540 1422
rect 1534 1417 1540 1418
rect 1622 1422 1628 1423
rect 1622 1418 1623 1422
rect 1627 1418 1628 1422
rect 1622 1417 1628 1418
rect 1718 1422 1724 1423
rect 1718 1418 1719 1422
rect 1723 1418 1724 1422
rect 1718 1417 1724 1418
rect 1822 1422 1828 1423
rect 1822 1418 1823 1422
rect 1827 1418 1828 1422
rect 1822 1417 1828 1418
rect 1926 1422 1932 1423
rect 1926 1418 1927 1422
rect 1931 1418 1932 1422
rect 1926 1417 1932 1418
rect 2022 1422 2028 1423
rect 2022 1418 2023 1422
rect 2027 1418 2028 1422
rect 2022 1417 2028 1418
rect 2118 1422 2124 1423
rect 2118 1418 2119 1422
rect 2123 1418 2124 1422
rect 2118 1417 2124 1418
rect 2214 1422 2220 1423
rect 2214 1418 2215 1422
rect 2219 1418 2220 1422
rect 2214 1417 2220 1418
rect 2302 1422 2308 1423
rect 2302 1418 2303 1422
rect 2307 1418 2308 1422
rect 2302 1417 2308 1418
rect 2390 1422 2396 1423
rect 2390 1418 2391 1422
rect 2395 1418 2396 1422
rect 2390 1417 2396 1418
rect 2478 1422 2484 1423
rect 2478 1418 2479 1422
rect 2483 1418 2484 1422
rect 2478 1417 2484 1418
rect 2542 1422 2548 1423
rect 2542 1418 2543 1422
rect 2547 1418 2548 1422
rect 2542 1417 2548 1418
rect 2584 1414 2586 1429
rect 1366 1413 1372 1414
rect 110 1409 116 1410
rect 110 1405 111 1409
rect 115 1405 116 1409
rect 110 1404 116 1405
rect 1326 1409 1332 1410
rect 1326 1405 1327 1409
rect 1331 1405 1332 1409
rect 1366 1409 1367 1413
rect 1371 1409 1372 1413
rect 1366 1408 1372 1409
rect 2582 1413 2588 1414
rect 2582 1409 2583 1413
rect 2587 1409 2588 1413
rect 2582 1408 2588 1409
rect 1326 1404 1332 1405
rect 1366 1396 1372 1397
rect 2582 1396 2588 1397
rect 110 1392 116 1393
rect 1326 1392 1332 1393
rect 110 1388 111 1392
rect 115 1388 116 1392
rect 110 1387 116 1388
rect 142 1391 148 1392
rect 142 1387 143 1391
rect 147 1387 148 1391
rect 112 1375 114 1387
rect 142 1386 148 1387
rect 230 1391 236 1392
rect 230 1387 231 1391
rect 235 1387 236 1391
rect 230 1386 236 1387
rect 326 1391 332 1392
rect 326 1387 327 1391
rect 331 1387 332 1391
rect 326 1386 332 1387
rect 430 1391 436 1392
rect 430 1387 431 1391
rect 435 1387 436 1391
rect 430 1386 436 1387
rect 534 1391 540 1392
rect 534 1387 535 1391
rect 539 1387 540 1391
rect 534 1386 540 1387
rect 646 1391 652 1392
rect 646 1387 647 1391
rect 651 1387 652 1391
rect 646 1386 652 1387
rect 750 1391 756 1392
rect 750 1387 751 1391
rect 755 1387 756 1391
rect 750 1386 756 1387
rect 862 1391 868 1392
rect 862 1387 863 1391
rect 867 1387 868 1391
rect 862 1386 868 1387
rect 974 1391 980 1392
rect 974 1387 975 1391
rect 979 1387 980 1391
rect 974 1386 980 1387
rect 1086 1391 1092 1392
rect 1086 1387 1087 1391
rect 1091 1387 1092 1391
rect 1086 1386 1092 1387
rect 1198 1391 1204 1392
rect 1198 1387 1199 1391
rect 1203 1387 1204 1391
rect 1326 1388 1327 1392
rect 1331 1388 1332 1392
rect 1366 1392 1367 1396
rect 1371 1392 1372 1396
rect 1366 1391 1372 1392
rect 1398 1395 1404 1396
rect 1398 1391 1399 1395
rect 1403 1391 1404 1395
rect 1326 1387 1332 1388
rect 1198 1386 1204 1387
rect 144 1375 146 1386
rect 232 1375 234 1386
rect 328 1375 330 1386
rect 432 1375 434 1386
rect 536 1375 538 1386
rect 648 1375 650 1386
rect 752 1375 754 1386
rect 864 1375 866 1386
rect 976 1375 978 1386
rect 1088 1375 1090 1386
rect 1200 1375 1202 1386
rect 1328 1375 1330 1387
rect 111 1374 115 1375
rect 111 1369 115 1370
rect 143 1374 147 1375
rect 143 1369 147 1370
rect 207 1374 211 1375
rect 207 1369 211 1370
rect 231 1374 235 1375
rect 231 1369 235 1370
rect 295 1374 299 1375
rect 295 1369 299 1370
rect 327 1374 331 1375
rect 327 1369 331 1370
rect 399 1374 403 1375
rect 399 1369 403 1370
rect 431 1374 435 1375
rect 431 1369 435 1370
rect 511 1374 515 1375
rect 511 1369 515 1370
rect 535 1374 539 1375
rect 535 1369 539 1370
rect 623 1374 627 1375
rect 623 1369 627 1370
rect 647 1374 651 1375
rect 647 1369 651 1370
rect 735 1374 739 1375
rect 735 1369 739 1370
rect 751 1374 755 1375
rect 751 1369 755 1370
rect 847 1374 851 1375
rect 847 1369 851 1370
rect 863 1374 867 1375
rect 863 1369 867 1370
rect 959 1374 963 1375
rect 959 1369 963 1370
rect 975 1374 979 1375
rect 975 1369 979 1370
rect 1071 1374 1075 1375
rect 1071 1369 1075 1370
rect 1087 1374 1091 1375
rect 1087 1369 1091 1370
rect 1183 1374 1187 1375
rect 1183 1369 1187 1370
rect 1199 1374 1203 1375
rect 1199 1369 1203 1370
rect 1271 1374 1275 1375
rect 1271 1369 1275 1370
rect 1327 1374 1331 1375
rect 1368 1371 1370 1391
rect 1398 1390 1404 1391
rect 1454 1395 1460 1396
rect 1454 1391 1455 1395
rect 1459 1391 1460 1395
rect 1454 1390 1460 1391
rect 1518 1395 1524 1396
rect 1518 1391 1519 1395
rect 1523 1391 1524 1395
rect 1518 1390 1524 1391
rect 1606 1395 1612 1396
rect 1606 1391 1607 1395
rect 1611 1391 1612 1395
rect 1606 1390 1612 1391
rect 1702 1395 1708 1396
rect 1702 1391 1703 1395
rect 1707 1391 1708 1395
rect 1702 1390 1708 1391
rect 1806 1395 1812 1396
rect 1806 1391 1807 1395
rect 1811 1391 1812 1395
rect 1806 1390 1812 1391
rect 1910 1395 1916 1396
rect 1910 1391 1911 1395
rect 1915 1391 1916 1395
rect 1910 1390 1916 1391
rect 2006 1395 2012 1396
rect 2006 1391 2007 1395
rect 2011 1391 2012 1395
rect 2006 1390 2012 1391
rect 2102 1395 2108 1396
rect 2102 1391 2103 1395
rect 2107 1391 2108 1395
rect 2102 1390 2108 1391
rect 2198 1395 2204 1396
rect 2198 1391 2199 1395
rect 2203 1391 2204 1395
rect 2198 1390 2204 1391
rect 2286 1395 2292 1396
rect 2286 1391 2287 1395
rect 2291 1391 2292 1395
rect 2286 1390 2292 1391
rect 2374 1395 2380 1396
rect 2374 1391 2375 1395
rect 2379 1391 2380 1395
rect 2374 1390 2380 1391
rect 2462 1395 2468 1396
rect 2462 1391 2463 1395
rect 2467 1391 2468 1395
rect 2462 1390 2468 1391
rect 2526 1395 2532 1396
rect 2526 1391 2527 1395
rect 2531 1391 2532 1395
rect 2582 1392 2583 1396
rect 2587 1392 2588 1396
rect 2582 1391 2588 1392
rect 2526 1390 2532 1391
rect 1400 1371 1402 1390
rect 1456 1371 1458 1390
rect 1520 1371 1522 1390
rect 1608 1371 1610 1390
rect 1704 1371 1706 1390
rect 1808 1371 1810 1390
rect 1912 1371 1914 1390
rect 2008 1371 2010 1390
rect 2104 1371 2106 1390
rect 2200 1371 2202 1390
rect 2288 1371 2290 1390
rect 2376 1371 2378 1390
rect 2464 1371 2466 1390
rect 2528 1371 2530 1390
rect 2584 1371 2586 1391
rect 1327 1369 1331 1370
rect 1367 1370 1371 1371
rect 112 1357 114 1369
rect 144 1358 146 1369
rect 208 1358 210 1369
rect 296 1358 298 1369
rect 400 1358 402 1369
rect 512 1358 514 1369
rect 624 1358 626 1369
rect 736 1358 738 1369
rect 848 1358 850 1369
rect 960 1358 962 1369
rect 1072 1358 1074 1369
rect 1184 1358 1186 1369
rect 1272 1358 1274 1369
rect 142 1357 148 1358
rect 110 1356 116 1357
rect 110 1352 111 1356
rect 115 1352 116 1356
rect 142 1353 143 1357
rect 147 1353 148 1357
rect 142 1352 148 1353
rect 206 1357 212 1358
rect 206 1353 207 1357
rect 211 1353 212 1357
rect 206 1352 212 1353
rect 294 1357 300 1358
rect 294 1353 295 1357
rect 299 1353 300 1357
rect 294 1352 300 1353
rect 398 1357 404 1358
rect 398 1353 399 1357
rect 403 1353 404 1357
rect 398 1352 404 1353
rect 510 1357 516 1358
rect 510 1353 511 1357
rect 515 1353 516 1357
rect 510 1352 516 1353
rect 622 1357 628 1358
rect 622 1353 623 1357
rect 627 1353 628 1357
rect 622 1352 628 1353
rect 734 1357 740 1358
rect 734 1353 735 1357
rect 739 1353 740 1357
rect 734 1352 740 1353
rect 846 1357 852 1358
rect 846 1353 847 1357
rect 851 1353 852 1357
rect 846 1352 852 1353
rect 958 1357 964 1358
rect 958 1353 959 1357
rect 963 1353 964 1357
rect 958 1352 964 1353
rect 1070 1357 1076 1358
rect 1070 1353 1071 1357
rect 1075 1353 1076 1357
rect 1070 1352 1076 1353
rect 1182 1357 1188 1358
rect 1182 1353 1183 1357
rect 1187 1353 1188 1357
rect 1182 1352 1188 1353
rect 1270 1357 1276 1358
rect 1328 1357 1330 1369
rect 1367 1365 1371 1366
rect 1399 1370 1403 1371
rect 1399 1365 1403 1366
rect 1455 1370 1459 1371
rect 1455 1365 1459 1366
rect 1519 1370 1523 1371
rect 1519 1365 1523 1366
rect 1543 1370 1547 1371
rect 1543 1365 1547 1366
rect 1607 1370 1611 1371
rect 1607 1365 1611 1366
rect 1631 1370 1635 1371
rect 1631 1365 1635 1366
rect 1703 1370 1707 1371
rect 1703 1365 1707 1366
rect 1719 1370 1723 1371
rect 1719 1365 1723 1366
rect 1807 1370 1811 1371
rect 1807 1365 1811 1366
rect 1887 1370 1891 1371
rect 1887 1365 1891 1366
rect 1911 1370 1915 1371
rect 1911 1365 1915 1366
rect 1967 1370 1971 1371
rect 1967 1365 1971 1366
rect 2007 1370 2011 1371
rect 2007 1365 2011 1366
rect 2047 1370 2051 1371
rect 2047 1365 2051 1366
rect 2103 1370 2107 1371
rect 2103 1365 2107 1366
rect 2127 1370 2131 1371
rect 2127 1365 2131 1366
rect 2199 1370 2203 1371
rect 2199 1365 2203 1366
rect 2207 1370 2211 1371
rect 2207 1365 2211 1366
rect 2287 1370 2291 1371
rect 2287 1365 2291 1366
rect 2375 1370 2379 1371
rect 2375 1365 2379 1366
rect 2463 1370 2467 1371
rect 2463 1365 2467 1366
rect 2527 1370 2531 1371
rect 2527 1365 2531 1366
rect 2583 1370 2587 1371
rect 2583 1365 2587 1366
rect 1270 1353 1271 1357
rect 1275 1353 1276 1357
rect 1270 1352 1276 1353
rect 1326 1356 1332 1357
rect 1326 1352 1327 1356
rect 1331 1352 1332 1356
rect 1368 1353 1370 1365
rect 1400 1354 1402 1365
rect 1456 1354 1458 1365
rect 1544 1354 1546 1365
rect 1632 1354 1634 1365
rect 1720 1354 1722 1365
rect 1808 1354 1810 1365
rect 1888 1354 1890 1365
rect 1968 1354 1970 1365
rect 2048 1354 2050 1365
rect 2128 1354 2130 1365
rect 2208 1354 2210 1365
rect 1398 1353 1404 1354
rect 110 1351 116 1352
rect 1326 1351 1332 1352
rect 1366 1352 1372 1353
rect 1366 1348 1367 1352
rect 1371 1348 1372 1352
rect 1398 1349 1399 1353
rect 1403 1349 1404 1353
rect 1398 1348 1404 1349
rect 1454 1353 1460 1354
rect 1454 1349 1455 1353
rect 1459 1349 1460 1353
rect 1454 1348 1460 1349
rect 1542 1353 1548 1354
rect 1542 1349 1543 1353
rect 1547 1349 1548 1353
rect 1542 1348 1548 1349
rect 1630 1353 1636 1354
rect 1630 1349 1631 1353
rect 1635 1349 1636 1353
rect 1630 1348 1636 1349
rect 1718 1353 1724 1354
rect 1718 1349 1719 1353
rect 1723 1349 1724 1353
rect 1718 1348 1724 1349
rect 1806 1353 1812 1354
rect 1806 1349 1807 1353
rect 1811 1349 1812 1353
rect 1806 1348 1812 1349
rect 1886 1353 1892 1354
rect 1886 1349 1887 1353
rect 1891 1349 1892 1353
rect 1886 1348 1892 1349
rect 1966 1353 1972 1354
rect 1966 1349 1967 1353
rect 1971 1349 1972 1353
rect 1966 1348 1972 1349
rect 2046 1353 2052 1354
rect 2046 1349 2047 1353
rect 2051 1349 2052 1353
rect 2046 1348 2052 1349
rect 2126 1353 2132 1354
rect 2126 1349 2127 1353
rect 2131 1349 2132 1353
rect 2126 1348 2132 1349
rect 2206 1353 2212 1354
rect 2584 1353 2586 1365
rect 2206 1349 2207 1353
rect 2211 1349 2212 1353
rect 2206 1348 2212 1349
rect 2582 1352 2588 1353
rect 2582 1348 2583 1352
rect 2587 1348 2588 1352
rect 1366 1347 1372 1348
rect 2582 1347 2588 1348
rect 110 1339 116 1340
rect 110 1335 111 1339
rect 115 1335 116 1339
rect 110 1334 116 1335
rect 1326 1339 1332 1340
rect 1326 1335 1327 1339
rect 1331 1335 1332 1339
rect 1326 1334 1332 1335
rect 1366 1335 1372 1336
rect 112 1319 114 1334
rect 158 1330 164 1331
rect 158 1326 159 1330
rect 163 1326 164 1330
rect 158 1325 164 1326
rect 222 1330 228 1331
rect 222 1326 223 1330
rect 227 1326 228 1330
rect 222 1325 228 1326
rect 310 1330 316 1331
rect 310 1326 311 1330
rect 315 1326 316 1330
rect 310 1325 316 1326
rect 414 1330 420 1331
rect 414 1326 415 1330
rect 419 1326 420 1330
rect 414 1325 420 1326
rect 526 1330 532 1331
rect 526 1326 527 1330
rect 531 1326 532 1330
rect 526 1325 532 1326
rect 638 1330 644 1331
rect 638 1326 639 1330
rect 643 1326 644 1330
rect 638 1325 644 1326
rect 750 1330 756 1331
rect 750 1326 751 1330
rect 755 1326 756 1330
rect 750 1325 756 1326
rect 862 1330 868 1331
rect 862 1326 863 1330
rect 867 1326 868 1330
rect 862 1325 868 1326
rect 974 1330 980 1331
rect 974 1326 975 1330
rect 979 1326 980 1330
rect 974 1325 980 1326
rect 1086 1330 1092 1331
rect 1086 1326 1087 1330
rect 1091 1326 1092 1330
rect 1086 1325 1092 1326
rect 1198 1330 1204 1331
rect 1198 1326 1199 1330
rect 1203 1326 1204 1330
rect 1198 1325 1204 1326
rect 1286 1330 1292 1331
rect 1286 1326 1287 1330
rect 1291 1326 1292 1330
rect 1286 1325 1292 1326
rect 160 1319 162 1325
rect 224 1319 226 1325
rect 312 1319 314 1325
rect 416 1319 418 1325
rect 528 1319 530 1325
rect 640 1319 642 1325
rect 752 1319 754 1325
rect 864 1319 866 1325
rect 976 1319 978 1325
rect 1088 1319 1090 1325
rect 1200 1319 1202 1325
rect 1288 1319 1290 1325
rect 1328 1319 1330 1334
rect 1366 1331 1367 1335
rect 1371 1331 1372 1335
rect 1366 1330 1372 1331
rect 2582 1335 2588 1336
rect 2582 1331 2583 1335
rect 2587 1331 2588 1335
rect 2582 1330 2588 1331
rect 111 1318 115 1319
rect 111 1313 115 1314
rect 159 1318 163 1319
rect 159 1313 163 1314
rect 223 1318 227 1319
rect 223 1313 227 1314
rect 231 1318 235 1319
rect 231 1313 235 1314
rect 311 1318 315 1319
rect 311 1313 315 1314
rect 327 1318 331 1319
rect 327 1313 331 1314
rect 415 1318 419 1319
rect 415 1313 419 1314
rect 431 1318 435 1319
rect 431 1313 435 1314
rect 527 1318 531 1319
rect 527 1313 531 1314
rect 535 1318 539 1319
rect 535 1313 539 1314
rect 631 1318 635 1319
rect 631 1313 635 1314
rect 639 1318 643 1319
rect 639 1313 643 1314
rect 727 1318 731 1319
rect 727 1313 731 1314
rect 751 1318 755 1319
rect 751 1313 755 1314
rect 823 1318 827 1319
rect 823 1313 827 1314
rect 863 1318 867 1319
rect 863 1313 867 1314
rect 911 1318 915 1319
rect 911 1313 915 1314
rect 975 1318 979 1319
rect 975 1313 979 1314
rect 991 1318 995 1319
rect 991 1313 995 1314
rect 1071 1318 1075 1319
rect 1071 1313 1075 1314
rect 1087 1318 1091 1319
rect 1087 1313 1091 1314
rect 1151 1318 1155 1319
rect 1151 1313 1155 1314
rect 1199 1318 1203 1319
rect 1199 1313 1203 1314
rect 1231 1318 1235 1319
rect 1231 1313 1235 1314
rect 1287 1318 1291 1319
rect 1287 1313 1291 1314
rect 1327 1318 1331 1319
rect 1327 1313 1331 1314
rect 112 1298 114 1313
rect 160 1307 162 1313
rect 232 1307 234 1313
rect 328 1307 330 1313
rect 432 1307 434 1313
rect 536 1307 538 1313
rect 632 1307 634 1313
rect 728 1307 730 1313
rect 824 1307 826 1313
rect 912 1307 914 1313
rect 992 1307 994 1313
rect 1072 1307 1074 1313
rect 1152 1307 1154 1313
rect 1232 1307 1234 1313
rect 1288 1307 1290 1313
rect 158 1306 164 1307
rect 158 1302 159 1306
rect 163 1302 164 1306
rect 158 1301 164 1302
rect 230 1306 236 1307
rect 230 1302 231 1306
rect 235 1302 236 1306
rect 230 1301 236 1302
rect 326 1306 332 1307
rect 326 1302 327 1306
rect 331 1302 332 1306
rect 326 1301 332 1302
rect 430 1306 436 1307
rect 430 1302 431 1306
rect 435 1302 436 1306
rect 430 1301 436 1302
rect 534 1306 540 1307
rect 534 1302 535 1306
rect 539 1302 540 1306
rect 534 1301 540 1302
rect 630 1306 636 1307
rect 630 1302 631 1306
rect 635 1302 636 1306
rect 630 1301 636 1302
rect 726 1306 732 1307
rect 726 1302 727 1306
rect 731 1302 732 1306
rect 726 1301 732 1302
rect 822 1306 828 1307
rect 822 1302 823 1306
rect 827 1302 828 1306
rect 822 1301 828 1302
rect 910 1306 916 1307
rect 910 1302 911 1306
rect 915 1302 916 1306
rect 910 1301 916 1302
rect 990 1306 996 1307
rect 990 1302 991 1306
rect 995 1302 996 1306
rect 990 1301 996 1302
rect 1070 1306 1076 1307
rect 1070 1302 1071 1306
rect 1075 1302 1076 1306
rect 1070 1301 1076 1302
rect 1150 1306 1156 1307
rect 1150 1302 1151 1306
rect 1155 1302 1156 1306
rect 1150 1301 1156 1302
rect 1230 1306 1236 1307
rect 1230 1302 1231 1306
rect 1235 1302 1236 1306
rect 1230 1301 1236 1302
rect 1286 1306 1292 1307
rect 1286 1302 1287 1306
rect 1291 1302 1292 1306
rect 1286 1301 1292 1302
rect 1328 1298 1330 1313
rect 1368 1311 1370 1330
rect 1414 1326 1420 1327
rect 1414 1322 1415 1326
rect 1419 1322 1420 1326
rect 1414 1321 1420 1322
rect 1470 1326 1476 1327
rect 1470 1322 1471 1326
rect 1475 1322 1476 1326
rect 1470 1321 1476 1322
rect 1558 1326 1564 1327
rect 1558 1322 1559 1326
rect 1563 1322 1564 1326
rect 1558 1321 1564 1322
rect 1646 1326 1652 1327
rect 1646 1322 1647 1326
rect 1651 1322 1652 1326
rect 1646 1321 1652 1322
rect 1734 1326 1740 1327
rect 1734 1322 1735 1326
rect 1739 1322 1740 1326
rect 1734 1321 1740 1322
rect 1822 1326 1828 1327
rect 1822 1322 1823 1326
rect 1827 1322 1828 1326
rect 1822 1321 1828 1322
rect 1902 1326 1908 1327
rect 1902 1322 1903 1326
rect 1907 1322 1908 1326
rect 1902 1321 1908 1322
rect 1982 1326 1988 1327
rect 1982 1322 1983 1326
rect 1987 1322 1988 1326
rect 1982 1321 1988 1322
rect 2062 1326 2068 1327
rect 2062 1322 2063 1326
rect 2067 1322 2068 1326
rect 2062 1321 2068 1322
rect 2142 1326 2148 1327
rect 2142 1322 2143 1326
rect 2147 1322 2148 1326
rect 2142 1321 2148 1322
rect 2222 1326 2228 1327
rect 2222 1322 2223 1326
rect 2227 1322 2228 1326
rect 2222 1321 2228 1322
rect 1416 1311 1418 1321
rect 1472 1311 1474 1321
rect 1560 1311 1562 1321
rect 1648 1311 1650 1321
rect 1736 1311 1738 1321
rect 1824 1311 1826 1321
rect 1904 1311 1906 1321
rect 1984 1311 1986 1321
rect 2064 1311 2066 1321
rect 2144 1311 2146 1321
rect 2224 1311 2226 1321
rect 2584 1311 2586 1330
rect 1367 1310 1371 1311
rect 1367 1305 1371 1306
rect 1415 1310 1419 1311
rect 1415 1305 1419 1306
rect 1471 1310 1475 1311
rect 1471 1305 1475 1306
rect 1559 1310 1563 1311
rect 1559 1305 1563 1306
rect 1647 1310 1651 1311
rect 1647 1305 1651 1306
rect 1671 1310 1675 1311
rect 1671 1305 1675 1306
rect 1735 1310 1739 1311
rect 1735 1305 1739 1306
rect 1767 1310 1771 1311
rect 1767 1305 1771 1306
rect 1823 1310 1827 1311
rect 1823 1305 1827 1306
rect 1863 1310 1867 1311
rect 1863 1305 1867 1306
rect 1903 1310 1907 1311
rect 1903 1305 1907 1306
rect 1959 1310 1963 1311
rect 1959 1305 1963 1306
rect 1983 1310 1987 1311
rect 1983 1305 1987 1306
rect 2047 1310 2051 1311
rect 2047 1305 2051 1306
rect 2063 1310 2067 1311
rect 2063 1305 2067 1306
rect 2135 1310 2139 1311
rect 2135 1305 2139 1306
rect 2143 1310 2147 1311
rect 2143 1305 2147 1306
rect 2223 1310 2227 1311
rect 2223 1305 2227 1306
rect 2231 1310 2235 1311
rect 2231 1305 2235 1306
rect 2583 1310 2587 1311
rect 2583 1305 2587 1306
rect 110 1297 116 1298
rect 110 1293 111 1297
rect 115 1293 116 1297
rect 110 1292 116 1293
rect 1326 1297 1332 1298
rect 1326 1293 1327 1297
rect 1331 1293 1332 1297
rect 1326 1292 1332 1293
rect 1368 1290 1370 1305
rect 1672 1299 1674 1305
rect 1768 1299 1770 1305
rect 1864 1299 1866 1305
rect 1960 1299 1962 1305
rect 2048 1299 2050 1305
rect 2136 1299 2138 1305
rect 2232 1299 2234 1305
rect 1670 1298 1676 1299
rect 1670 1294 1671 1298
rect 1675 1294 1676 1298
rect 1670 1293 1676 1294
rect 1766 1298 1772 1299
rect 1766 1294 1767 1298
rect 1771 1294 1772 1298
rect 1766 1293 1772 1294
rect 1862 1298 1868 1299
rect 1862 1294 1863 1298
rect 1867 1294 1868 1298
rect 1862 1293 1868 1294
rect 1958 1298 1964 1299
rect 1958 1294 1959 1298
rect 1963 1294 1964 1298
rect 1958 1293 1964 1294
rect 2046 1298 2052 1299
rect 2046 1294 2047 1298
rect 2051 1294 2052 1298
rect 2046 1293 2052 1294
rect 2134 1298 2140 1299
rect 2134 1294 2135 1298
rect 2139 1294 2140 1298
rect 2134 1293 2140 1294
rect 2230 1298 2236 1299
rect 2230 1294 2231 1298
rect 2235 1294 2236 1298
rect 2230 1293 2236 1294
rect 2584 1290 2586 1305
rect 1366 1289 1372 1290
rect 1366 1285 1367 1289
rect 1371 1285 1372 1289
rect 1366 1284 1372 1285
rect 2582 1289 2588 1290
rect 2582 1285 2583 1289
rect 2587 1285 2588 1289
rect 2582 1284 2588 1285
rect 110 1280 116 1281
rect 1326 1280 1332 1281
rect 110 1276 111 1280
rect 115 1276 116 1280
rect 110 1275 116 1276
rect 142 1279 148 1280
rect 142 1275 143 1279
rect 147 1275 148 1279
rect 112 1251 114 1275
rect 142 1274 148 1275
rect 214 1279 220 1280
rect 214 1275 215 1279
rect 219 1275 220 1279
rect 214 1274 220 1275
rect 310 1279 316 1280
rect 310 1275 311 1279
rect 315 1275 316 1279
rect 310 1274 316 1275
rect 414 1279 420 1280
rect 414 1275 415 1279
rect 419 1275 420 1279
rect 414 1274 420 1275
rect 518 1279 524 1280
rect 518 1275 519 1279
rect 523 1275 524 1279
rect 518 1274 524 1275
rect 614 1279 620 1280
rect 614 1275 615 1279
rect 619 1275 620 1279
rect 614 1274 620 1275
rect 710 1279 716 1280
rect 710 1275 711 1279
rect 715 1275 716 1279
rect 710 1274 716 1275
rect 806 1279 812 1280
rect 806 1275 807 1279
rect 811 1275 812 1279
rect 806 1274 812 1275
rect 894 1279 900 1280
rect 894 1275 895 1279
rect 899 1275 900 1279
rect 894 1274 900 1275
rect 974 1279 980 1280
rect 974 1275 975 1279
rect 979 1275 980 1279
rect 974 1274 980 1275
rect 1054 1279 1060 1280
rect 1054 1275 1055 1279
rect 1059 1275 1060 1279
rect 1054 1274 1060 1275
rect 1134 1279 1140 1280
rect 1134 1275 1135 1279
rect 1139 1275 1140 1279
rect 1134 1274 1140 1275
rect 1214 1279 1220 1280
rect 1214 1275 1215 1279
rect 1219 1275 1220 1279
rect 1214 1274 1220 1275
rect 1270 1279 1276 1280
rect 1270 1275 1271 1279
rect 1275 1275 1276 1279
rect 1326 1276 1327 1280
rect 1331 1276 1332 1280
rect 1326 1275 1332 1276
rect 1270 1274 1276 1275
rect 144 1251 146 1274
rect 216 1251 218 1274
rect 312 1251 314 1274
rect 416 1251 418 1274
rect 520 1251 522 1274
rect 616 1251 618 1274
rect 712 1251 714 1274
rect 808 1251 810 1274
rect 896 1251 898 1274
rect 976 1251 978 1274
rect 1056 1251 1058 1274
rect 1136 1251 1138 1274
rect 1216 1251 1218 1274
rect 1272 1251 1274 1274
rect 1328 1251 1330 1275
rect 1366 1272 1372 1273
rect 2582 1272 2588 1273
rect 1366 1268 1367 1272
rect 1371 1268 1372 1272
rect 1366 1267 1372 1268
rect 1654 1271 1660 1272
rect 1654 1267 1655 1271
rect 1659 1267 1660 1271
rect 1368 1255 1370 1267
rect 1654 1266 1660 1267
rect 1750 1271 1756 1272
rect 1750 1267 1751 1271
rect 1755 1267 1756 1271
rect 1750 1266 1756 1267
rect 1846 1271 1852 1272
rect 1846 1267 1847 1271
rect 1851 1267 1852 1271
rect 1846 1266 1852 1267
rect 1942 1271 1948 1272
rect 1942 1267 1943 1271
rect 1947 1267 1948 1271
rect 1942 1266 1948 1267
rect 2030 1271 2036 1272
rect 2030 1267 2031 1271
rect 2035 1267 2036 1271
rect 2030 1266 2036 1267
rect 2118 1271 2124 1272
rect 2118 1267 2119 1271
rect 2123 1267 2124 1271
rect 2118 1266 2124 1267
rect 2214 1271 2220 1272
rect 2214 1267 2215 1271
rect 2219 1267 2220 1271
rect 2582 1268 2583 1272
rect 2587 1268 2588 1272
rect 2582 1267 2588 1268
rect 2214 1266 2220 1267
rect 1656 1255 1658 1266
rect 1752 1255 1754 1266
rect 1848 1255 1850 1266
rect 1944 1255 1946 1266
rect 2032 1255 2034 1266
rect 2120 1255 2122 1266
rect 2216 1255 2218 1266
rect 2584 1255 2586 1267
rect 1367 1254 1371 1255
rect 111 1250 115 1251
rect 111 1245 115 1246
rect 143 1250 147 1251
rect 143 1245 147 1246
rect 199 1250 203 1251
rect 199 1245 203 1246
rect 215 1250 219 1251
rect 215 1245 219 1246
rect 279 1250 283 1251
rect 279 1245 283 1246
rect 311 1250 315 1251
rect 311 1245 315 1246
rect 359 1250 363 1251
rect 359 1245 363 1246
rect 415 1250 419 1251
rect 415 1245 419 1246
rect 439 1250 443 1251
rect 439 1245 443 1246
rect 519 1250 523 1251
rect 519 1245 523 1246
rect 599 1250 603 1251
rect 599 1245 603 1246
rect 615 1250 619 1251
rect 615 1245 619 1246
rect 671 1250 675 1251
rect 671 1245 675 1246
rect 711 1250 715 1251
rect 711 1245 715 1246
rect 743 1250 747 1251
rect 743 1245 747 1246
rect 807 1250 811 1251
rect 807 1245 811 1246
rect 815 1250 819 1251
rect 815 1245 819 1246
rect 895 1250 899 1251
rect 895 1245 899 1246
rect 975 1250 979 1251
rect 975 1245 979 1246
rect 1055 1250 1059 1251
rect 1055 1245 1059 1246
rect 1135 1250 1139 1251
rect 1135 1245 1139 1246
rect 1215 1250 1219 1251
rect 1215 1245 1219 1246
rect 1271 1250 1275 1251
rect 1271 1245 1275 1246
rect 1327 1250 1331 1251
rect 1367 1249 1371 1250
rect 1495 1254 1499 1255
rect 1495 1249 1499 1250
rect 1559 1254 1563 1255
rect 1559 1249 1563 1250
rect 1623 1254 1627 1255
rect 1623 1249 1627 1250
rect 1655 1254 1659 1255
rect 1655 1249 1659 1250
rect 1687 1254 1691 1255
rect 1687 1249 1691 1250
rect 1751 1254 1755 1255
rect 1751 1249 1755 1250
rect 1759 1254 1763 1255
rect 1759 1249 1763 1250
rect 1823 1254 1827 1255
rect 1823 1249 1827 1250
rect 1847 1254 1851 1255
rect 1847 1249 1851 1250
rect 1887 1254 1891 1255
rect 1887 1249 1891 1250
rect 1943 1254 1947 1255
rect 1943 1249 1947 1250
rect 1951 1254 1955 1255
rect 1951 1249 1955 1250
rect 2015 1254 2019 1255
rect 2015 1249 2019 1250
rect 2031 1254 2035 1255
rect 2031 1249 2035 1250
rect 2079 1254 2083 1255
rect 2079 1249 2083 1250
rect 2119 1254 2123 1255
rect 2119 1249 2123 1250
rect 2151 1254 2155 1255
rect 2151 1249 2155 1250
rect 2215 1254 2219 1255
rect 2215 1249 2219 1250
rect 2223 1254 2227 1255
rect 2223 1249 2227 1250
rect 2295 1254 2299 1255
rect 2295 1249 2299 1250
rect 2583 1254 2587 1255
rect 2583 1249 2587 1250
rect 1327 1245 1331 1246
rect 112 1233 114 1245
rect 144 1234 146 1245
rect 200 1234 202 1245
rect 280 1234 282 1245
rect 360 1234 362 1245
rect 440 1234 442 1245
rect 520 1234 522 1245
rect 600 1234 602 1245
rect 672 1234 674 1245
rect 744 1234 746 1245
rect 816 1234 818 1245
rect 896 1234 898 1245
rect 142 1233 148 1234
rect 110 1232 116 1233
rect 110 1228 111 1232
rect 115 1228 116 1232
rect 142 1229 143 1233
rect 147 1229 148 1233
rect 142 1228 148 1229
rect 198 1233 204 1234
rect 198 1229 199 1233
rect 203 1229 204 1233
rect 198 1228 204 1229
rect 278 1233 284 1234
rect 278 1229 279 1233
rect 283 1229 284 1233
rect 278 1228 284 1229
rect 358 1233 364 1234
rect 358 1229 359 1233
rect 363 1229 364 1233
rect 358 1228 364 1229
rect 438 1233 444 1234
rect 438 1229 439 1233
rect 443 1229 444 1233
rect 438 1228 444 1229
rect 518 1233 524 1234
rect 518 1229 519 1233
rect 523 1229 524 1233
rect 518 1228 524 1229
rect 598 1233 604 1234
rect 598 1229 599 1233
rect 603 1229 604 1233
rect 598 1228 604 1229
rect 670 1233 676 1234
rect 670 1229 671 1233
rect 675 1229 676 1233
rect 670 1228 676 1229
rect 742 1233 748 1234
rect 742 1229 743 1233
rect 747 1229 748 1233
rect 742 1228 748 1229
rect 814 1233 820 1234
rect 814 1229 815 1233
rect 819 1229 820 1233
rect 814 1228 820 1229
rect 894 1233 900 1234
rect 1328 1233 1330 1245
rect 1368 1237 1370 1249
rect 1496 1238 1498 1249
rect 1560 1238 1562 1249
rect 1624 1238 1626 1249
rect 1688 1238 1690 1249
rect 1760 1238 1762 1249
rect 1824 1238 1826 1249
rect 1888 1238 1890 1249
rect 1952 1238 1954 1249
rect 2016 1238 2018 1249
rect 2080 1238 2082 1249
rect 2152 1238 2154 1249
rect 2224 1238 2226 1249
rect 2296 1238 2298 1249
rect 1494 1237 1500 1238
rect 1366 1236 1372 1237
rect 894 1229 895 1233
rect 899 1229 900 1233
rect 894 1228 900 1229
rect 1326 1232 1332 1233
rect 1326 1228 1327 1232
rect 1331 1228 1332 1232
rect 1366 1232 1367 1236
rect 1371 1232 1372 1236
rect 1494 1233 1495 1237
rect 1499 1233 1500 1237
rect 1494 1232 1500 1233
rect 1558 1237 1564 1238
rect 1558 1233 1559 1237
rect 1563 1233 1564 1237
rect 1558 1232 1564 1233
rect 1622 1237 1628 1238
rect 1622 1233 1623 1237
rect 1627 1233 1628 1237
rect 1622 1232 1628 1233
rect 1686 1237 1692 1238
rect 1686 1233 1687 1237
rect 1691 1233 1692 1237
rect 1686 1232 1692 1233
rect 1758 1237 1764 1238
rect 1758 1233 1759 1237
rect 1763 1233 1764 1237
rect 1758 1232 1764 1233
rect 1822 1237 1828 1238
rect 1822 1233 1823 1237
rect 1827 1233 1828 1237
rect 1822 1232 1828 1233
rect 1886 1237 1892 1238
rect 1886 1233 1887 1237
rect 1891 1233 1892 1237
rect 1886 1232 1892 1233
rect 1950 1237 1956 1238
rect 1950 1233 1951 1237
rect 1955 1233 1956 1237
rect 1950 1232 1956 1233
rect 2014 1237 2020 1238
rect 2014 1233 2015 1237
rect 2019 1233 2020 1237
rect 2014 1232 2020 1233
rect 2078 1237 2084 1238
rect 2078 1233 2079 1237
rect 2083 1233 2084 1237
rect 2078 1232 2084 1233
rect 2150 1237 2156 1238
rect 2150 1233 2151 1237
rect 2155 1233 2156 1237
rect 2150 1232 2156 1233
rect 2222 1237 2228 1238
rect 2222 1233 2223 1237
rect 2227 1233 2228 1237
rect 2222 1232 2228 1233
rect 2294 1237 2300 1238
rect 2584 1237 2586 1249
rect 2294 1233 2295 1237
rect 2299 1233 2300 1237
rect 2294 1232 2300 1233
rect 2582 1236 2588 1237
rect 2582 1232 2583 1236
rect 2587 1232 2588 1236
rect 1366 1231 1372 1232
rect 2582 1231 2588 1232
rect 110 1227 116 1228
rect 1326 1227 1332 1228
rect 1366 1219 1372 1220
rect 110 1215 116 1216
rect 110 1211 111 1215
rect 115 1211 116 1215
rect 110 1210 116 1211
rect 1326 1215 1332 1216
rect 1326 1211 1327 1215
rect 1331 1211 1332 1215
rect 1366 1215 1367 1219
rect 1371 1215 1372 1219
rect 1366 1214 1372 1215
rect 2582 1219 2588 1220
rect 2582 1215 2583 1219
rect 2587 1215 2588 1219
rect 2582 1214 2588 1215
rect 1326 1210 1332 1211
rect 112 1191 114 1210
rect 158 1206 164 1207
rect 158 1202 159 1206
rect 163 1202 164 1206
rect 158 1201 164 1202
rect 214 1206 220 1207
rect 214 1202 215 1206
rect 219 1202 220 1206
rect 214 1201 220 1202
rect 294 1206 300 1207
rect 294 1202 295 1206
rect 299 1202 300 1206
rect 294 1201 300 1202
rect 374 1206 380 1207
rect 374 1202 375 1206
rect 379 1202 380 1206
rect 374 1201 380 1202
rect 454 1206 460 1207
rect 454 1202 455 1206
rect 459 1202 460 1206
rect 454 1201 460 1202
rect 534 1206 540 1207
rect 534 1202 535 1206
rect 539 1202 540 1206
rect 534 1201 540 1202
rect 614 1206 620 1207
rect 614 1202 615 1206
rect 619 1202 620 1206
rect 614 1201 620 1202
rect 686 1206 692 1207
rect 686 1202 687 1206
rect 691 1202 692 1206
rect 686 1201 692 1202
rect 758 1206 764 1207
rect 758 1202 759 1206
rect 763 1202 764 1206
rect 758 1201 764 1202
rect 830 1206 836 1207
rect 830 1202 831 1206
rect 835 1202 836 1206
rect 830 1201 836 1202
rect 910 1206 916 1207
rect 910 1202 911 1206
rect 915 1202 916 1206
rect 910 1201 916 1202
rect 160 1191 162 1201
rect 216 1191 218 1201
rect 296 1191 298 1201
rect 376 1191 378 1201
rect 456 1191 458 1201
rect 536 1191 538 1201
rect 616 1191 618 1201
rect 688 1191 690 1201
rect 760 1191 762 1201
rect 832 1191 834 1201
rect 912 1191 914 1201
rect 1328 1191 1330 1210
rect 1368 1191 1370 1214
rect 1510 1210 1516 1211
rect 1510 1206 1511 1210
rect 1515 1206 1516 1210
rect 1510 1205 1516 1206
rect 1574 1210 1580 1211
rect 1574 1206 1575 1210
rect 1579 1206 1580 1210
rect 1574 1205 1580 1206
rect 1638 1210 1644 1211
rect 1638 1206 1639 1210
rect 1643 1206 1644 1210
rect 1638 1205 1644 1206
rect 1702 1210 1708 1211
rect 1702 1206 1703 1210
rect 1707 1206 1708 1210
rect 1702 1205 1708 1206
rect 1774 1210 1780 1211
rect 1774 1206 1775 1210
rect 1779 1206 1780 1210
rect 1774 1205 1780 1206
rect 1838 1210 1844 1211
rect 1838 1206 1839 1210
rect 1843 1206 1844 1210
rect 1838 1205 1844 1206
rect 1902 1210 1908 1211
rect 1902 1206 1903 1210
rect 1907 1206 1908 1210
rect 1902 1205 1908 1206
rect 1966 1210 1972 1211
rect 1966 1206 1967 1210
rect 1971 1206 1972 1210
rect 1966 1205 1972 1206
rect 2030 1210 2036 1211
rect 2030 1206 2031 1210
rect 2035 1206 2036 1210
rect 2030 1205 2036 1206
rect 2094 1210 2100 1211
rect 2094 1206 2095 1210
rect 2099 1206 2100 1210
rect 2094 1205 2100 1206
rect 2166 1210 2172 1211
rect 2166 1206 2167 1210
rect 2171 1206 2172 1210
rect 2166 1205 2172 1206
rect 2238 1210 2244 1211
rect 2238 1206 2239 1210
rect 2243 1206 2244 1210
rect 2238 1205 2244 1206
rect 2310 1210 2316 1211
rect 2310 1206 2311 1210
rect 2315 1206 2316 1210
rect 2310 1205 2316 1206
rect 1512 1191 1514 1205
rect 1576 1191 1578 1205
rect 1640 1191 1642 1205
rect 1704 1191 1706 1205
rect 1776 1191 1778 1205
rect 1840 1191 1842 1205
rect 1904 1191 1906 1205
rect 1968 1191 1970 1205
rect 2032 1191 2034 1205
rect 2096 1191 2098 1205
rect 2168 1191 2170 1205
rect 2240 1191 2242 1205
rect 2312 1191 2314 1205
rect 2584 1191 2586 1214
rect 111 1190 115 1191
rect 111 1185 115 1186
rect 159 1190 163 1191
rect 159 1185 163 1186
rect 215 1190 219 1191
rect 215 1185 219 1186
rect 239 1190 243 1191
rect 239 1185 243 1186
rect 295 1190 299 1191
rect 295 1185 299 1186
rect 327 1190 331 1191
rect 327 1185 331 1186
rect 375 1190 379 1191
rect 375 1185 379 1186
rect 423 1190 427 1191
rect 423 1185 427 1186
rect 455 1190 459 1191
rect 455 1185 459 1186
rect 511 1190 515 1191
rect 511 1185 515 1186
rect 535 1190 539 1191
rect 535 1185 539 1186
rect 599 1190 603 1191
rect 599 1185 603 1186
rect 615 1190 619 1191
rect 615 1185 619 1186
rect 687 1190 691 1191
rect 687 1185 691 1186
rect 759 1190 763 1191
rect 759 1185 763 1186
rect 767 1190 771 1191
rect 767 1185 771 1186
rect 831 1190 835 1191
rect 831 1185 835 1186
rect 839 1190 843 1191
rect 839 1185 843 1186
rect 911 1190 915 1191
rect 911 1185 915 1186
rect 983 1190 987 1191
rect 983 1185 987 1186
rect 1063 1190 1067 1191
rect 1063 1185 1067 1186
rect 1327 1190 1331 1191
rect 1327 1185 1331 1186
rect 1367 1190 1371 1191
rect 1367 1185 1371 1186
rect 1415 1190 1419 1191
rect 1415 1185 1419 1186
rect 1503 1190 1507 1191
rect 1503 1185 1507 1186
rect 1511 1190 1515 1191
rect 1511 1185 1515 1186
rect 1575 1190 1579 1191
rect 1575 1185 1579 1186
rect 1599 1190 1603 1191
rect 1599 1185 1603 1186
rect 1639 1190 1643 1191
rect 1639 1185 1643 1186
rect 1703 1190 1707 1191
rect 1703 1185 1707 1186
rect 1775 1190 1779 1191
rect 1775 1185 1779 1186
rect 1807 1190 1811 1191
rect 1807 1185 1811 1186
rect 1839 1190 1843 1191
rect 1839 1185 1843 1186
rect 1903 1190 1907 1191
rect 1903 1185 1907 1186
rect 1911 1190 1915 1191
rect 1911 1185 1915 1186
rect 1967 1190 1971 1191
rect 1967 1185 1971 1186
rect 2015 1190 2019 1191
rect 2015 1185 2019 1186
rect 2031 1190 2035 1191
rect 2031 1185 2035 1186
rect 2095 1190 2099 1191
rect 2095 1185 2099 1186
rect 2111 1190 2115 1191
rect 2111 1185 2115 1186
rect 2167 1190 2171 1191
rect 2167 1185 2171 1186
rect 2207 1190 2211 1191
rect 2207 1185 2211 1186
rect 2239 1190 2243 1191
rect 2239 1185 2243 1186
rect 2303 1190 2307 1191
rect 2303 1185 2307 1186
rect 2311 1190 2315 1191
rect 2311 1185 2315 1186
rect 2399 1190 2403 1191
rect 2399 1185 2403 1186
rect 2583 1190 2587 1191
rect 2583 1185 2587 1186
rect 112 1170 114 1185
rect 160 1179 162 1185
rect 240 1179 242 1185
rect 328 1179 330 1185
rect 424 1179 426 1185
rect 512 1179 514 1185
rect 600 1179 602 1185
rect 688 1179 690 1185
rect 768 1179 770 1185
rect 840 1179 842 1185
rect 912 1179 914 1185
rect 984 1179 986 1185
rect 1064 1179 1066 1185
rect 158 1178 164 1179
rect 158 1174 159 1178
rect 163 1174 164 1178
rect 158 1173 164 1174
rect 238 1178 244 1179
rect 238 1174 239 1178
rect 243 1174 244 1178
rect 238 1173 244 1174
rect 326 1178 332 1179
rect 326 1174 327 1178
rect 331 1174 332 1178
rect 326 1173 332 1174
rect 422 1178 428 1179
rect 422 1174 423 1178
rect 427 1174 428 1178
rect 422 1173 428 1174
rect 510 1178 516 1179
rect 510 1174 511 1178
rect 515 1174 516 1178
rect 510 1173 516 1174
rect 598 1178 604 1179
rect 598 1174 599 1178
rect 603 1174 604 1178
rect 598 1173 604 1174
rect 686 1178 692 1179
rect 686 1174 687 1178
rect 691 1174 692 1178
rect 686 1173 692 1174
rect 766 1178 772 1179
rect 766 1174 767 1178
rect 771 1174 772 1178
rect 766 1173 772 1174
rect 838 1178 844 1179
rect 838 1174 839 1178
rect 843 1174 844 1178
rect 838 1173 844 1174
rect 910 1178 916 1179
rect 910 1174 911 1178
rect 915 1174 916 1178
rect 910 1173 916 1174
rect 982 1178 988 1179
rect 982 1174 983 1178
rect 987 1174 988 1178
rect 982 1173 988 1174
rect 1062 1178 1068 1179
rect 1062 1174 1063 1178
rect 1067 1174 1068 1178
rect 1062 1173 1068 1174
rect 1328 1170 1330 1185
rect 1368 1170 1370 1185
rect 1416 1179 1418 1185
rect 1504 1179 1506 1185
rect 1600 1179 1602 1185
rect 1704 1179 1706 1185
rect 1808 1179 1810 1185
rect 1912 1179 1914 1185
rect 2016 1179 2018 1185
rect 2112 1179 2114 1185
rect 2208 1179 2210 1185
rect 2304 1179 2306 1185
rect 2400 1179 2402 1185
rect 1414 1178 1420 1179
rect 1414 1174 1415 1178
rect 1419 1174 1420 1178
rect 1414 1173 1420 1174
rect 1502 1178 1508 1179
rect 1502 1174 1503 1178
rect 1507 1174 1508 1178
rect 1502 1173 1508 1174
rect 1598 1178 1604 1179
rect 1598 1174 1599 1178
rect 1603 1174 1604 1178
rect 1598 1173 1604 1174
rect 1702 1178 1708 1179
rect 1702 1174 1703 1178
rect 1707 1174 1708 1178
rect 1702 1173 1708 1174
rect 1806 1178 1812 1179
rect 1806 1174 1807 1178
rect 1811 1174 1812 1178
rect 1806 1173 1812 1174
rect 1910 1178 1916 1179
rect 1910 1174 1911 1178
rect 1915 1174 1916 1178
rect 1910 1173 1916 1174
rect 2014 1178 2020 1179
rect 2014 1174 2015 1178
rect 2019 1174 2020 1178
rect 2014 1173 2020 1174
rect 2110 1178 2116 1179
rect 2110 1174 2111 1178
rect 2115 1174 2116 1178
rect 2110 1173 2116 1174
rect 2206 1178 2212 1179
rect 2206 1174 2207 1178
rect 2211 1174 2212 1178
rect 2206 1173 2212 1174
rect 2302 1178 2308 1179
rect 2302 1174 2303 1178
rect 2307 1174 2308 1178
rect 2302 1173 2308 1174
rect 2398 1178 2404 1179
rect 2398 1174 2399 1178
rect 2403 1174 2404 1178
rect 2398 1173 2404 1174
rect 2584 1170 2586 1185
rect 110 1169 116 1170
rect 110 1165 111 1169
rect 115 1165 116 1169
rect 110 1164 116 1165
rect 1326 1169 1332 1170
rect 1326 1165 1327 1169
rect 1331 1165 1332 1169
rect 1326 1164 1332 1165
rect 1366 1169 1372 1170
rect 1366 1165 1367 1169
rect 1371 1165 1372 1169
rect 1366 1164 1372 1165
rect 2582 1169 2588 1170
rect 2582 1165 2583 1169
rect 2587 1165 2588 1169
rect 2582 1164 2588 1165
rect 110 1152 116 1153
rect 1326 1152 1332 1153
rect 110 1148 111 1152
rect 115 1148 116 1152
rect 110 1147 116 1148
rect 142 1151 148 1152
rect 142 1147 143 1151
rect 147 1147 148 1151
rect 112 1127 114 1147
rect 142 1146 148 1147
rect 222 1151 228 1152
rect 222 1147 223 1151
rect 227 1147 228 1151
rect 222 1146 228 1147
rect 310 1151 316 1152
rect 310 1147 311 1151
rect 315 1147 316 1151
rect 310 1146 316 1147
rect 406 1151 412 1152
rect 406 1147 407 1151
rect 411 1147 412 1151
rect 406 1146 412 1147
rect 494 1151 500 1152
rect 494 1147 495 1151
rect 499 1147 500 1151
rect 494 1146 500 1147
rect 582 1151 588 1152
rect 582 1147 583 1151
rect 587 1147 588 1151
rect 582 1146 588 1147
rect 670 1151 676 1152
rect 670 1147 671 1151
rect 675 1147 676 1151
rect 670 1146 676 1147
rect 750 1151 756 1152
rect 750 1147 751 1151
rect 755 1147 756 1151
rect 750 1146 756 1147
rect 822 1151 828 1152
rect 822 1147 823 1151
rect 827 1147 828 1151
rect 822 1146 828 1147
rect 894 1151 900 1152
rect 894 1147 895 1151
rect 899 1147 900 1151
rect 894 1146 900 1147
rect 966 1151 972 1152
rect 966 1147 967 1151
rect 971 1147 972 1151
rect 966 1146 972 1147
rect 1046 1151 1052 1152
rect 1046 1147 1047 1151
rect 1051 1147 1052 1151
rect 1326 1148 1327 1152
rect 1331 1148 1332 1152
rect 1326 1147 1332 1148
rect 1366 1152 1372 1153
rect 2582 1152 2588 1153
rect 1366 1148 1367 1152
rect 1371 1148 1372 1152
rect 1366 1147 1372 1148
rect 1398 1151 1404 1152
rect 1398 1147 1399 1151
rect 1403 1147 1404 1151
rect 1046 1146 1052 1147
rect 144 1127 146 1146
rect 224 1127 226 1146
rect 312 1127 314 1146
rect 408 1127 410 1146
rect 496 1127 498 1146
rect 584 1127 586 1146
rect 672 1127 674 1146
rect 752 1127 754 1146
rect 824 1127 826 1146
rect 896 1127 898 1146
rect 968 1127 970 1146
rect 1048 1127 1050 1146
rect 1328 1127 1330 1147
rect 1368 1131 1370 1147
rect 1398 1146 1404 1147
rect 1486 1151 1492 1152
rect 1486 1147 1487 1151
rect 1491 1147 1492 1151
rect 1486 1146 1492 1147
rect 1582 1151 1588 1152
rect 1582 1147 1583 1151
rect 1587 1147 1588 1151
rect 1582 1146 1588 1147
rect 1686 1151 1692 1152
rect 1686 1147 1687 1151
rect 1691 1147 1692 1151
rect 1686 1146 1692 1147
rect 1790 1151 1796 1152
rect 1790 1147 1791 1151
rect 1795 1147 1796 1151
rect 1790 1146 1796 1147
rect 1894 1151 1900 1152
rect 1894 1147 1895 1151
rect 1899 1147 1900 1151
rect 1894 1146 1900 1147
rect 1998 1151 2004 1152
rect 1998 1147 1999 1151
rect 2003 1147 2004 1151
rect 1998 1146 2004 1147
rect 2094 1151 2100 1152
rect 2094 1147 2095 1151
rect 2099 1147 2100 1151
rect 2094 1146 2100 1147
rect 2190 1151 2196 1152
rect 2190 1147 2191 1151
rect 2195 1147 2196 1151
rect 2190 1146 2196 1147
rect 2286 1151 2292 1152
rect 2286 1147 2287 1151
rect 2291 1147 2292 1151
rect 2286 1146 2292 1147
rect 2382 1151 2388 1152
rect 2382 1147 2383 1151
rect 2387 1147 2388 1151
rect 2582 1148 2583 1152
rect 2587 1148 2588 1152
rect 2582 1147 2588 1148
rect 2382 1146 2388 1147
rect 1400 1131 1402 1146
rect 1488 1131 1490 1146
rect 1584 1131 1586 1146
rect 1688 1131 1690 1146
rect 1792 1131 1794 1146
rect 1896 1131 1898 1146
rect 2000 1131 2002 1146
rect 2096 1131 2098 1146
rect 2192 1131 2194 1146
rect 2288 1131 2290 1146
rect 2384 1131 2386 1146
rect 2584 1131 2586 1147
rect 1367 1130 1371 1131
rect 111 1126 115 1127
rect 111 1121 115 1122
rect 143 1126 147 1127
rect 143 1121 147 1122
rect 223 1126 227 1127
rect 223 1121 227 1122
rect 311 1126 315 1127
rect 311 1121 315 1122
rect 319 1126 323 1127
rect 319 1121 323 1122
rect 407 1126 411 1127
rect 407 1121 411 1122
rect 423 1126 427 1127
rect 423 1121 427 1122
rect 495 1126 499 1127
rect 495 1121 499 1122
rect 527 1126 531 1127
rect 527 1121 531 1122
rect 583 1126 587 1127
rect 583 1121 587 1122
rect 631 1126 635 1127
rect 631 1121 635 1122
rect 671 1126 675 1127
rect 671 1121 675 1122
rect 727 1126 731 1127
rect 727 1121 731 1122
rect 751 1126 755 1127
rect 751 1121 755 1122
rect 823 1126 827 1127
rect 823 1121 827 1122
rect 895 1126 899 1127
rect 895 1121 899 1122
rect 911 1126 915 1127
rect 911 1121 915 1122
rect 967 1126 971 1127
rect 967 1121 971 1122
rect 991 1126 995 1127
rect 991 1121 995 1122
rect 1047 1126 1051 1127
rect 1047 1121 1051 1122
rect 1079 1126 1083 1127
rect 1079 1121 1083 1122
rect 1167 1126 1171 1127
rect 1167 1121 1171 1122
rect 1327 1126 1331 1127
rect 1367 1125 1371 1126
rect 1399 1130 1403 1131
rect 1399 1125 1403 1126
rect 1479 1130 1483 1131
rect 1479 1125 1483 1126
rect 1487 1130 1491 1131
rect 1487 1125 1491 1126
rect 1583 1130 1587 1131
rect 1583 1125 1587 1126
rect 1687 1130 1691 1131
rect 1687 1125 1691 1126
rect 1791 1130 1795 1131
rect 1791 1125 1795 1126
rect 1887 1130 1891 1131
rect 1887 1125 1891 1126
rect 1895 1130 1899 1131
rect 1895 1125 1899 1126
rect 1975 1130 1979 1131
rect 1975 1125 1979 1126
rect 1999 1130 2003 1131
rect 1999 1125 2003 1126
rect 2063 1130 2067 1131
rect 2063 1125 2067 1126
rect 2095 1130 2099 1131
rect 2095 1125 2099 1126
rect 2143 1130 2147 1131
rect 2143 1125 2147 1126
rect 2191 1130 2195 1131
rect 2191 1125 2195 1126
rect 2215 1130 2219 1131
rect 2215 1125 2219 1126
rect 2279 1130 2283 1131
rect 2279 1125 2283 1126
rect 2287 1130 2291 1131
rect 2287 1125 2291 1126
rect 2343 1130 2347 1131
rect 2343 1125 2347 1126
rect 2383 1130 2387 1131
rect 2383 1125 2387 1126
rect 2407 1130 2411 1131
rect 2407 1125 2411 1126
rect 2471 1130 2475 1131
rect 2471 1125 2475 1126
rect 2527 1130 2531 1131
rect 2527 1125 2531 1126
rect 2583 1130 2587 1131
rect 2583 1125 2587 1126
rect 1327 1121 1331 1122
rect 112 1109 114 1121
rect 224 1110 226 1121
rect 320 1110 322 1121
rect 424 1110 426 1121
rect 528 1110 530 1121
rect 632 1110 634 1121
rect 728 1110 730 1121
rect 824 1110 826 1121
rect 912 1110 914 1121
rect 992 1110 994 1121
rect 1080 1110 1082 1121
rect 1168 1110 1170 1121
rect 222 1109 228 1110
rect 110 1108 116 1109
rect 110 1104 111 1108
rect 115 1104 116 1108
rect 222 1105 223 1109
rect 227 1105 228 1109
rect 222 1104 228 1105
rect 318 1109 324 1110
rect 318 1105 319 1109
rect 323 1105 324 1109
rect 318 1104 324 1105
rect 422 1109 428 1110
rect 422 1105 423 1109
rect 427 1105 428 1109
rect 422 1104 428 1105
rect 526 1109 532 1110
rect 526 1105 527 1109
rect 531 1105 532 1109
rect 526 1104 532 1105
rect 630 1109 636 1110
rect 630 1105 631 1109
rect 635 1105 636 1109
rect 630 1104 636 1105
rect 726 1109 732 1110
rect 726 1105 727 1109
rect 731 1105 732 1109
rect 726 1104 732 1105
rect 822 1109 828 1110
rect 822 1105 823 1109
rect 827 1105 828 1109
rect 822 1104 828 1105
rect 910 1109 916 1110
rect 910 1105 911 1109
rect 915 1105 916 1109
rect 910 1104 916 1105
rect 990 1109 996 1110
rect 990 1105 991 1109
rect 995 1105 996 1109
rect 990 1104 996 1105
rect 1078 1109 1084 1110
rect 1078 1105 1079 1109
rect 1083 1105 1084 1109
rect 1078 1104 1084 1105
rect 1166 1109 1172 1110
rect 1328 1109 1330 1121
rect 1368 1113 1370 1125
rect 1400 1114 1402 1125
rect 1480 1114 1482 1125
rect 1584 1114 1586 1125
rect 1688 1114 1690 1125
rect 1792 1114 1794 1125
rect 1888 1114 1890 1125
rect 1976 1114 1978 1125
rect 2064 1114 2066 1125
rect 2144 1114 2146 1125
rect 2216 1114 2218 1125
rect 2280 1114 2282 1125
rect 2344 1114 2346 1125
rect 2408 1114 2410 1125
rect 2472 1114 2474 1125
rect 2528 1114 2530 1125
rect 1398 1113 1404 1114
rect 1366 1112 1372 1113
rect 1166 1105 1167 1109
rect 1171 1105 1172 1109
rect 1166 1104 1172 1105
rect 1326 1108 1332 1109
rect 1326 1104 1327 1108
rect 1331 1104 1332 1108
rect 1366 1108 1367 1112
rect 1371 1108 1372 1112
rect 1398 1109 1399 1113
rect 1403 1109 1404 1113
rect 1398 1108 1404 1109
rect 1478 1113 1484 1114
rect 1478 1109 1479 1113
rect 1483 1109 1484 1113
rect 1478 1108 1484 1109
rect 1582 1113 1588 1114
rect 1582 1109 1583 1113
rect 1587 1109 1588 1113
rect 1582 1108 1588 1109
rect 1686 1113 1692 1114
rect 1686 1109 1687 1113
rect 1691 1109 1692 1113
rect 1686 1108 1692 1109
rect 1790 1113 1796 1114
rect 1790 1109 1791 1113
rect 1795 1109 1796 1113
rect 1790 1108 1796 1109
rect 1886 1113 1892 1114
rect 1886 1109 1887 1113
rect 1891 1109 1892 1113
rect 1886 1108 1892 1109
rect 1974 1113 1980 1114
rect 1974 1109 1975 1113
rect 1979 1109 1980 1113
rect 1974 1108 1980 1109
rect 2062 1113 2068 1114
rect 2062 1109 2063 1113
rect 2067 1109 2068 1113
rect 2062 1108 2068 1109
rect 2142 1113 2148 1114
rect 2142 1109 2143 1113
rect 2147 1109 2148 1113
rect 2142 1108 2148 1109
rect 2214 1113 2220 1114
rect 2214 1109 2215 1113
rect 2219 1109 2220 1113
rect 2214 1108 2220 1109
rect 2278 1113 2284 1114
rect 2278 1109 2279 1113
rect 2283 1109 2284 1113
rect 2278 1108 2284 1109
rect 2342 1113 2348 1114
rect 2342 1109 2343 1113
rect 2347 1109 2348 1113
rect 2342 1108 2348 1109
rect 2406 1113 2412 1114
rect 2406 1109 2407 1113
rect 2411 1109 2412 1113
rect 2406 1108 2412 1109
rect 2470 1113 2476 1114
rect 2470 1109 2471 1113
rect 2475 1109 2476 1113
rect 2470 1108 2476 1109
rect 2526 1113 2532 1114
rect 2584 1113 2586 1125
rect 2526 1109 2527 1113
rect 2531 1109 2532 1113
rect 2526 1108 2532 1109
rect 2582 1112 2588 1113
rect 2582 1108 2583 1112
rect 2587 1108 2588 1112
rect 1366 1107 1372 1108
rect 2582 1107 2588 1108
rect 110 1103 116 1104
rect 1326 1103 1332 1104
rect 1366 1095 1372 1096
rect 110 1091 116 1092
rect 110 1087 111 1091
rect 115 1087 116 1091
rect 110 1086 116 1087
rect 1326 1091 1332 1092
rect 1326 1087 1327 1091
rect 1331 1087 1332 1091
rect 1366 1091 1367 1095
rect 1371 1091 1372 1095
rect 1366 1090 1372 1091
rect 2582 1095 2588 1096
rect 2582 1091 2583 1095
rect 2587 1091 2588 1095
rect 2582 1090 2588 1091
rect 1326 1086 1332 1087
rect 112 1067 114 1086
rect 238 1082 244 1083
rect 238 1078 239 1082
rect 243 1078 244 1082
rect 238 1077 244 1078
rect 334 1082 340 1083
rect 334 1078 335 1082
rect 339 1078 340 1082
rect 334 1077 340 1078
rect 438 1082 444 1083
rect 438 1078 439 1082
rect 443 1078 444 1082
rect 438 1077 444 1078
rect 542 1082 548 1083
rect 542 1078 543 1082
rect 547 1078 548 1082
rect 542 1077 548 1078
rect 646 1082 652 1083
rect 646 1078 647 1082
rect 651 1078 652 1082
rect 646 1077 652 1078
rect 742 1082 748 1083
rect 742 1078 743 1082
rect 747 1078 748 1082
rect 742 1077 748 1078
rect 838 1082 844 1083
rect 838 1078 839 1082
rect 843 1078 844 1082
rect 838 1077 844 1078
rect 926 1082 932 1083
rect 926 1078 927 1082
rect 931 1078 932 1082
rect 926 1077 932 1078
rect 1006 1082 1012 1083
rect 1006 1078 1007 1082
rect 1011 1078 1012 1082
rect 1006 1077 1012 1078
rect 1094 1082 1100 1083
rect 1094 1078 1095 1082
rect 1099 1078 1100 1082
rect 1094 1077 1100 1078
rect 1182 1082 1188 1083
rect 1182 1078 1183 1082
rect 1187 1078 1188 1082
rect 1182 1077 1188 1078
rect 240 1067 242 1077
rect 336 1067 338 1077
rect 440 1067 442 1077
rect 544 1067 546 1077
rect 648 1067 650 1077
rect 744 1067 746 1077
rect 840 1067 842 1077
rect 928 1067 930 1077
rect 1008 1067 1010 1077
rect 1096 1067 1098 1077
rect 1184 1067 1186 1077
rect 1328 1067 1330 1086
rect 1368 1071 1370 1090
rect 1414 1086 1420 1087
rect 1414 1082 1415 1086
rect 1419 1082 1420 1086
rect 1414 1081 1420 1082
rect 1494 1086 1500 1087
rect 1494 1082 1495 1086
rect 1499 1082 1500 1086
rect 1494 1081 1500 1082
rect 1598 1086 1604 1087
rect 1598 1082 1599 1086
rect 1603 1082 1604 1086
rect 1598 1081 1604 1082
rect 1702 1086 1708 1087
rect 1702 1082 1703 1086
rect 1707 1082 1708 1086
rect 1702 1081 1708 1082
rect 1806 1086 1812 1087
rect 1806 1082 1807 1086
rect 1811 1082 1812 1086
rect 1806 1081 1812 1082
rect 1902 1086 1908 1087
rect 1902 1082 1903 1086
rect 1907 1082 1908 1086
rect 1902 1081 1908 1082
rect 1990 1086 1996 1087
rect 1990 1082 1991 1086
rect 1995 1082 1996 1086
rect 1990 1081 1996 1082
rect 2078 1086 2084 1087
rect 2078 1082 2079 1086
rect 2083 1082 2084 1086
rect 2078 1081 2084 1082
rect 2158 1086 2164 1087
rect 2158 1082 2159 1086
rect 2163 1082 2164 1086
rect 2158 1081 2164 1082
rect 2230 1086 2236 1087
rect 2230 1082 2231 1086
rect 2235 1082 2236 1086
rect 2230 1081 2236 1082
rect 2294 1086 2300 1087
rect 2294 1082 2295 1086
rect 2299 1082 2300 1086
rect 2294 1081 2300 1082
rect 2358 1086 2364 1087
rect 2358 1082 2359 1086
rect 2363 1082 2364 1086
rect 2358 1081 2364 1082
rect 2422 1086 2428 1087
rect 2422 1082 2423 1086
rect 2427 1082 2428 1086
rect 2422 1081 2428 1082
rect 2486 1086 2492 1087
rect 2486 1082 2487 1086
rect 2491 1082 2492 1086
rect 2486 1081 2492 1082
rect 2542 1086 2548 1087
rect 2542 1082 2543 1086
rect 2547 1082 2548 1086
rect 2542 1081 2548 1082
rect 1416 1071 1418 1081
rect 1496 1071 1498 1081
rect 1600 1071 1602 1081
rect 1704 1071 1706 1081
rect 1808 1071 1810 1081
rect 1904 1071 1906 1081
rect 1992 1071 1994 1081
rect 2080 1071 2082 1081
rect 2160 1071 2162 1081
rect 2232 1071 2234 1081
rect 2296 1071 2298 1081
rect 2360 1071 2362 1081
rect 2424 1071 2426 1081
rect 2488 1071 2490 1081
rect 2544 1071 2546 1081
rect 2584 1071 2586 1090
rect 1367 1070 1371 1071
rect 111 1066 115 1067
rect 111 1061 115 1062
rect 239 1066 243 1067
rect 239 1061 243 1062
rect 311 1066 315 1067
rect 311 1061 315 1062
rect 335 1066 339 1067
rect 335 1061 339 1062
rect 367 1066 371 1067
rect 367 1061 371 1062
rect 439 1066 443 1067
rect 439 1061 443 1062
rect 519 1066 523 1067
rect 519 1061 523 1062
rect 543 1066 547 1067
rect 543 1061 547 1062
rect 607 1066 611 1067
rect 607 1061 611 1062
rect 647 1066 651 1067
rect 647 1061 651 1062
rect 703 1066 707 1067
rect 703 1061 707 1062
rect 743 1066 747 1067
rect 743 1061 747 1062
rect 799 1066 803 1067
rect 799 1061 803 1062
rect 839 1066 843 1067
rect 839 1061 843 1062
rect 887 1066 891 1067
rect 887 1061 891 1062
rect 927 1066 931 1067
rect 927 1061 931 1062
rect 975 1066 979 1067
rect 975 1061 979 1062
rect 1007 1066 1011 1067
rect 1007 1061 1011 1062
rect 1055 1066 1059 1067
rect 1055 1061 1059 1062
rect 1095 1066 1099 1067
rect 1095 1061 1099 1062
rect 1135 1066 1139 1067
rect 1135 1061 1139 1062
rect 1183 1066 1187 1067
rect 1183 1061 1187 1062
rect 1223 1066 1227 1067
rect 1223 1061 1227 1062
rect 1287 1066 1291 1067
rect 1287 1061 1291 1062
rect 1327 1066 1331 1067
rect 1367 1065 1371 1066
rect 1415 1070 1419 1071
rect 1415 1065 1419 1066
rect 1471 1070 1475 1071
rect 1471 1065 1475 1066
rect 1495 1070 1499 1071
rect 1495 1065 1499 1066
rect 1535 1070 1539 1071
rect 1535 1065 1539 1066
rect 1599 1070 1603 1071
rect 1599 1065 1603 1066
rect 1623 1070 1627 1071
rect 1623 1065 1627 1066
rect 1703 1070 1707 1071
rect 1703 1065 1707 1066
rect 1727 1070 1731 1071
rect 1727 1065 1731 1066
rect 1807 1070 1811 1071
rect 1807 1065 1811 1066
rect 1839 1070 1843 1071
rect 1839 1065 1843 1066
rect 1903 1070 1907 1071
rect 1903 1065 1907 1066
rect 1951 1070 1955 1071
rect 1951 1065 1955 1066
rect 1991 1070 1995 1071
rect 1991 1065 1995 1066
rect 2063 1070 2067 1071
rect 2063 1065 2067 1066
rect 2079 1070 2083 1071
rect 2079 1065 2083 1066
rect 2159 1070 2163 1071
rect 2159 1065 2163 1066
rect 2167 1070 2171 1071
rect 2167 1065 2171 1066
rect 2231 1070 2235 1071
rect 2231 1065 2235 1066
rect 2271 1070 2275 1071
rect 2271 1065 2275 1066
rect 2295 1070 2299 1071
rect 2295 1065 2299 1066
rect 2359 1070 2363 1071
rect 2359 1065 2363 1066
rect 2367 1070 2371 1071
rect 2367 1065 2371 1066
rect 2423 1070 2427 1071
rect 2423 1065 2427 1066
rect 2463 1070 2467 1071
rect 2463 1065 2467 1066
rect 2487 1070 2491 1071
rect 2487 1065 2491 1066
rect 2543 1070 2547 1071
rect 2543 1065 2547 1066
rect 2583 1070 2587 1071
rect 2583 1065 2587 1066
rect 1327 1061 1331 1062
rect 112 1046 114 1061
rect 312 1055 314 1061
rect 368 1055 370 1061
rect 440 1055 442 1061
rect 520 1055 522 1061
rect 608 1055 610 1061
rect 704 1055 706 1061
rect 800 1055 802 1061
rect 888 1055 890 1061
rect 976 1055 978 1061
rect 1056 1055 1058 1061
rect 1136 1055 1138 1061
rect 1224 1055 1226 1061
rect 1288 1055 1290 1061
rect 310 1054 316 1055
rect 310 1050 311 1054
rect 315 1050 316 1054
rect 310 1049 316 1050
rect 366 1054 372 1055
rect 366 1050 367 1054
rect 371 1050 372 1054
rect 366 1049 372 1050
rect 438 1054 444 1055
rect 438 1050 439 1054
rect 443 1050 444 1054
rect 438 1049 444 1050
rect 518 1054 524 1055
rect 518 1050 519 1054
rect 523 1050 524 1054
rect 518 1049 524 1050
rect 606 1054 612 1055
rect 606 1050 607 1054
rect 611 1050 612 1054
rect 606 1049 612 1050
rect 702 1054 708 1055
rect 702 1050 703 1054
rect 707 1050 708 1054
rect 702 1049 708 1050
rect 798 1054 804 1055
rect 798 1050 799 1054
rect 803 1050 804 1054
rect 798 1049 804 1050
rect 886 1054 892 1055
rect 886 1050 887 1054
rect 891 1050 892 1054
rect 886 1049 892 1050
rect 974 1054 980 1055
rect 974 1050 975 1054
rect 979 1050 980 1054
rect 974 1049 980 1050
rect 1054 1054 1060 1055
rect 1054 1050 1055 1054
rect 1059 1050 1060 1054
rect 1054 1049 1060 1050
rect 1134 1054 1140 1055
rect 1134 1050 1135 1054
rect 1139 1050 1140 1054
rect 1134 1049 1140 1050
rect 1222 1054 1228 1055
rect 1222 1050 1223 1054
rect 1227 1050 1228 1054
rect 1222 1049 1228 1050
rect 1286 1054 1292 1055
rect 1286 1050 1287 1054
rect 1291 1050 1292 1054
rect 1286 1049 1292 1050
rect 1328 1046 1330 1061
rect 1368 1050 1370 1065
rect 1416 1059 1418 1065
rect 1472 1059 1474 1065
rect 1536 1059 1538 1065
rect 1624 1059 1626 1065
rect 1728 1059 1730 1065
rect 1840 1059 1842 1065
rect 1952 1059 1954 1065
rect 2064 1059 2066 1065
rect 2168 1059 2170 1065
rect 2272 1059 2274 1065
rect 2368 1059 2370 1065
rect 2464 1059 2466 1065
rect 2544 1059 2546 1065
rect 1414 1058 1420 1059
rect 1414 1054 1415 1058
rect 1419 1054 1420 1058
rect 1414 1053 1420 1054
rect 1470 1058 1476 1059
rect 1470 1054 1471 1058
rect 1475 1054 1476 1058
rect 1470 1053 1476 1054
rect 1534 1058 1540 1059
rect 1534 1054 1535 1058
rect 1539 1054 1540 1058
rect 1534 1053 1540 1054
rect 1622 1058 1628 1059
rect 1622 1054 1623 1058
rect 1627 1054 1628 1058
rect 1622 1053 1628 1054
rect 1726 1058 1732 1059
rect 1726 1054 1727 1058
rect 1731 1054 1732 1058
rect 1726 1053 1732 1054
rect 1838 1058 1844 1059
rect 1838 1054 1839 1058
rect 1843 1054 1844 1058
rect 1838 1053 1844 1054
rect 1950 1058 1956 1059
rect 1950 1054 1951 1058
rect 1955 1054 1956 1058
rect 1950 1053 1956 1054
rect 2062 1058 2068 1059
rect 2062 1054 2063 1058
rect 2067 1054 2068 1058
rect 2062 1053 2068 1054
rect 2166 1058 2172 1059
rect 2166 1054 2167 1058
rect 2171 1054 2172 1058
rect 2166 1053 2172 1054
rect 2270 1058 2276 1059
rect 2270 1054 2271 1058
rect 2275 1054 2276 1058
rect 2270 1053 2276 1054
rect 2366 1058 2372 1059
rect 2366 1054 2367 1058
rect 2371 1054 2372 1058
rect 2366 1053 2372 1054
rect 2462 1058 2468 1059
rect 2462 1054 2463 1058
rect 2467 1054 2468 1058
rect 2462 1053 2468 1054
rect 2542 1058 2548 1059
rect 2542 1054 2543 1058
rect 2547 1054 2548 1058
rect 2542 1053 2548 1054
rect 2584 1050 2586 1065
rect 1366 1049 1372 1050
rect 110 1045 116 1046
rect 110 1041 111 1045
rect 115 1041 116 1045
rect 110 1040 116 1041
rect 1326 1045 1332 1046
rect 1326 1041 1327 1045
rect 1331 1041 1332 1045
rect 1366 1045 1367 1049
rect 1371 1045 1372 1049
rect 1366 1044 1372 1045
rect 2582 1049 2588 1050
rect 2582 1045 2583 1049
rect 2587 1045 2588 1049
rect 2582 1044 2588 1045
rect 1326 1040 1332 1041
rect 1366 1032 1372 1033
rect 2582 1032 2588 1033
rect 110 1028 116 1029
rect 1326 1028 1332 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 110 1023 116 1024
rect 294 1027 300 1028
rect 294 1023 295 1027
rect 299 1023 300 1027
rect 112 1007 114 1023
rect 294 1022 300 1023
rect 350 1027 356 1028
rect 350 1023 351 1027
rect 355 1023 356 1027
rect 350 1022 356 1023
rect 422 1027 428 1028
rect 422 1023 423 1027
rect 427 1023 428 1027
rect 422 1022 428 1023
rect 502 1027 508 1028
rect 502 1023 503 1027
rect 507 1023 508 1027
rect 502 1022 508 1023
rect 590 1027 596 1028
rect 590 1023 591 1027
rect 595 1023 596 1027
rect 590 1022 596 1023
rect 686 1027 692 1028
rect 686 1023 687 1027
rect 691 1023 692 1027
rect 686 1022 692 1023
rect 782 1027 788 1028
rect 782 1023 783 1027
rect 787 1023 788 1027
rect 782 1022 788 1023
rect 870 1027 876 1028
rect 870 1023 871 1027
rect 875 1023 876 1027
rect 870 1022 876 1023
rect 958 1027 964 1028
rect 958 1023 959 1027
rect 963 1023 964 1027
rect 958 1022 964 1023
rect 1038 1027 1044 1028
rect 1038 1023 1039 1027
rect 1043 1023 1044 1027
rect 1038 1022 1044 1023
rect 1118 1027 1124 1028
rect 1118 1023 1119 1027
rect 1123 1023 1124 1027
rect 1118 1022 1124 1023
rect 1206 1027 1212 1028
rect 1206 1023 1207 1027
rect 1211 1023 1212 1027
rect 1206 1022 1212 1023
rect 1270 1027 1276 1028
rect 1270 1023 1271 1027
rect 1275 1023 1276 1027
rect 1326 1024 1327 1028
rect 1331 1024 1332 1028
rect 1366 1028 1367 1032
rect 1371 1028 1372 1032
rect 1366 1027 1372 1028
rect 1398 1031 1404 1032
rect 1398 1027 1399 1031
rect 1403 1027 1404 1031
rect 1326 1023 1332 1024
rect 1270 1022 1276 1023
rect 296 1007 298 1022
rect 352 1007 354 1022
rect 424 1007 426 1022
rect 504 1007 506 1022
rect 592 1007 594 1022
rect 688 1007 690 1022
rect 784 1007 786 1022
rect 872 1007 874 1022
rect 960 1007 962 1022
rect 1040 1007 1042 1022
rect 1120 1007 1122 1022
rect 1208 1007 1210 1022
rect 1272 1007 1274 1022
rect 1328 1007 1330 1023
rect 111 1006 115 1007
rect 111 1001 115 1002
rect 295 1006 299 1007
rect 295 1001 299 1002
rect 351 1006 355 1007
rect 351 1001 355 1002
rect 415 1006 419 1007
rect 415 1001 419 1002
rect 423 1006 427 1007
rect 423 1001 427 1002
rect 471 1006 475 1007
rect 471 1001 475 1002
rect 503 1006 507 1007
rect 503 1001 507 1002
rect 527 1006 531 1007
rect 527 1001 531 1002
rect 591 1006 595 1007
rect 591 1001 595 1002
rect 655 1006 659 1007
rect 655 1001 659 1002
rect 687 1006 691 1007
rect 687 1001 691 1002
rect 719 1006 723 1007
rect 719 1001 723 1002
rect 783 1006 787 1007
rect 783 1001 787 1002
rect 847 1006 851 1007
rect 847 1001 851 1002
rect 871 1006 875 1007
rect 871 1001 875 1002
rect 911 1006 915 1007
rect 911 1001 915 1002
rect 959 1006 963 1007
rect 959 1001 963 1002
rect 975 1006 979 1007
rect 975 1001 979 1002
rect 1039 1006 1043 1007
rect 1039 1001 1043 1002
rect 1103 1006 1107 1007
rect 1103 1001 1107 1002
rect 1119 1006 1123 1007
rect 1119 1001 1123 1002
rect 1159 1006 1163 1007
rect 1159 1001 1163 1002
rect 1207 1006 1211 1007
rect 1207 1001 1211 1002
rect 1215 1006 1219 1007
rect 1215 1001 1219 1002
rect 1271 1006 1275 1007
rect 1271 1001 1275 1002
rect 1327 1006 1331 1007
rect 1327 1001 1331 1002
rect 112 989 114 1001
rect 416 990 418 1001
rect 472 990 474 1001
rect 528 990 530 1001
rect 592 990 594 1001
rect 656 990 658 1001
rect 720 990 722 1001
rect 784 990 786 1001
rect 848 990 850 1001
rect 912 990 914 1001
rect 976 990 978 1001
rect 1040 990 1042 1001
rect 1104 990 1106 1001
rect 1160 990 1162 1001
rect 1216 990 1218 1001
rect 1272 990 1274 1001
rect 414 989 420 990
rect 110 988 116 989
rect 110 984 111 988
rect 115 984 116 988
rect 414 985 415 989
rect 419 985 420 989
rect 414 984 420 985
rect 470 989 476 990
rect 470 985 471 989
rect 475 985 476 989
rect 470 984 476 985
rect 526 989 532 990
rect 526 985 527 989
rect 531 985 532 989
rect 526 984 532 985
rect 590 989 596 990
rect 590 985 591 989
rect 595 985 596 989
rect 590 984 596 985
rect 654 989 660 990
rect 654 985 655 989
rect 659 985 660 989
rect 654 984 660 985
rect 718 989 724 990
rect 718 985 719 989
rect 723 985 724 989
rect 718 984 724 985
rect 782 989 788 990
rect 782 985 783 989
rect 787 985 788 989
rect 782 984 788 985
rect 846 989 852 990
rect 846 985 847 989
rect 851 985 852 989
rect 846 984 852 985
rect 910 989 916 990
rect 910 985 911 989
rect 915 985 916 989
rect 910 984 916 985
rect 974 989 980 990
rect 974 985 975 989
rect 979 985 980 989
rect 974 984 980 985
rect 1038 989 1044 990
rect 1038 985 1039 989
rect 1043 985 1044 989
rect 1038 984 1044 985
rect 1102 989 1108 990
rect 1102 985 1103 989
rect 1107 985 1108 989
rect 1102 984 1108 985
rect 1158 989 1164 990
rect 1158 985 1159 989
rect 1163 985 1164 989
rect 1158 984 1164 985
rect 1214 989 1220 990
rect 1214 985 1215 989
rect 1219 985 1220 989
rect 1214 984 1220 985
rect 1270 989 1276 990
rect 1328 989 1330 1001
rect 1368 999 1370 1027
rect 1398 1026 1404 1027
rect 1454 1031 1460 1032
rect 1454 1027 1455 1031
rect 1459 1027 1460 1031
rect 1454 1026 1460 1027
rect 1518 1031 1524 1032
rect 1518 1027 1519 1031
rect 1523 1027 1524 1031
rect 1518 1026 1524 1027
rect 1606 1031 1612 1032
rect 1606 1027 1607 1031
rect 1611 1027 1612 1031
rect 1606 1026 1612 1027
rect 1710 1031 1716 1032
rect 1710 1027 1711 1031
rect 1715 1027 1716 1031
rect 1710 1026 1716 1027
rect 1822 1031 1828 1032
rect 1822 1027 1823 1031
rect 1827 1027 1828 1031
rect 1822 1026 1828 1027
rect 1934 1031 1940 1032
rect 1934 1027 1935 1031
rect 1939 1027 1940 1031
rect 1934 1026 1940 1027
rect 2046 1031 2052 1032
rect 2046 1027 2047 1031
rect 2051 1027 2052 1031
rect 2046 1026 2052 1027
rect 2150 1031 2156 1032
rect 2150 1027 2151 1031
rect 2155 1027 2156 1031
rect 2150 1026 2156 1027
rect 2254 1031 2260 1032
rect 2254 1027 2255 1031
rect 2259 1027 2260 1031
rect 2254 1026 2260 1027
rect 2350 1031 2356 1032
rect 2350 1027 2351 1031
rect 2355 1027 2356 1031
rect 2350 1026 2356 1027
rect 2446 1031 2452 1032
rect 2446 1027 2447 1031
rect 2451 1027 2452 1031
rect 2446 1026 2452 1027
rect 2526 1031 2532 1032
rect 2526 1027 2527 1031
rect 2531 1027 2532 1031
rect 2582 1028 2583 1032
rect 2587 1028 2588 1032
rect 2582 1027 2588 1028
rect 2526 1026 2532 1027
rect 1400 999 1402 1026
rect 1456 999 1458 1026
rect 1520 999 1522 1026
rect 1608 999 1610 1026
rect 1712 999 1714 1026
rect 1824 999 1826 1026
rect 1936 999 1938 1026
rect 2048 999 2050 1026
rect 2152 999 2154 1026
rect 2256 999 2258 1026
rect 2352 999 2354 1026
rect 2448 999 2450 1026
rect 2528 999 2530 1026
rect 2584 999 2586 1027
rect 1367 998 1371 999
rect 1367 993 1371 994
rect 1399 998 1403 999
rect 1399 993 1403 994
rect 1455 998 1459 999
rect 1455 993 1459 994
rect 1511 998 1515 999
rect 1511 993 1515 994
rect 1519 998 1523 999
rect 1519 993 1523 994
rect 1567 998 1571 999
rect 1567 993 1571 994
rect 1607 998 1611 999
rect 1607 993 1611 994
rect 1639 998 1643 999
rect 1639 993 1643 994
rect 1711 998 1715 999
rect 1711 993 1715 994
rect 1719 998 1723 999
rect 1719 993 1723 994
rect 1807 998 1811 999
rect 1807 993 1811 994
rect 1823 998 1827 999
rect 1823 993 1827 994
rect 1903 998 1907 999
rect 1903 993 1907 994
rect 1935 998 1939 999
rect 1935 993 1939 994
rect 2015 998 2019 999
rect 2015 993 2019 994
rect 2047 998 2051 999
rect 2047 993 2051 994
rect 2143 998 2147 999
rect 2143 993 2147 994
rect 2151 998 2155 999
rect 2151 993 2155 994
rect 2255 998 2259 999
rect 2255 993 2259 994
rect 2271 998 2275 999
rect 2271 993 2275 994
rect 2351 998 2355 999
rect 2351 993 2355 994
rect 2407 998 2411 999
rect 2407 993 2411 994
rect 2447 998 2451 999
rect 2447 993 2451 994
rect 2527 998 2531 999
rect 2527 993 2531 994
rect 2583 998 2587 999
rect 2583 993 2587 994
rect 1270 985 1271 989
rect 1275 985 1276 989
rect 1270 984 1276 985
rect 1326 988 1332 989
rect 1326 984 1327 988
rect 1331 984 1332 988
rect 110 983 116 984
rect 1326 983 1332 984
rect 1368 981 1370 993
rect 1400 982 1402 993
rect 1456 982 1458 993
rect 1512 982 1514 993
rect 1568 982 1570 993
rect 1640 982 1642 993
rect 1720 982 1722 993
rect 1808 982 1810 993
rect 1904 982 1906 993
rect 2016 982 2018 993
rect 2144 982 2146 993
rect 2272 982 2274 993
rect 2408 982 2410 993
rect 2528 982 2530 993
rect 1398 981 1404 982
rect 1366 980 1372 981
rect 1366 976 1367 980
rect 1371 976 1372 980
rect 1398 977 1399 981
rect 1403 977 1404 981
rect 1398 976 1404 977
rect 1454 981 1460 982
rect 1454 977 1455 981
rect 1459 977 1460 981
rect 1454 976 1460 977
rect 1510 981 1516 982
rect 1510 977 1511 981
rect 1515 977 1516 981
rect 1510 976 1516 977
rect 1566 981 1572 982
rect 1566 977 1567 981
rect 1571 977 1572 981
rect 1566 976 1572 977
rect 1638 981 1644 982
rect 1638 977 1639 981
rect 1643 977 1644 981
rect 1638 976 1644 977
rect 1718 981 1724 982
rect 1718 977 1719 981
rect 1723 977 1724 981
rect 1718 976 1724 977
rect 1806 981 1812 982
rect 1806 977 1807 981
rect 1811 977 1812 981
rect 1806 976 1812 977
rect 1902 981 1908 982
rect 1902 977 1903 981
rect 1907 977 1908 981
rect 1902 976 1908 977
rect 2014 981 2020 982
rect 2014 977 2015 981
rect 2019 977 2020 981
rect 2014 976 2020 977
rect 2142 981 2148 982
rect 2142 977 2143 981
rect 2147 977 2148 981
rect 2142 976 2148 977
rect 2270 981 2276 982
rect 2270 977 2271 981
rect 2275 977 2276 981
rect 2270 976 2276 977
rect 2406 981 2412 982
rect 2406 977 2407 981
rect 2411 977 2412 981
rect 2406 976 2412 977
rect 2526 981 2532 982
rect 2584 981 2586 993
rect 2526 977 2527 981
rect 2531 977 2532 981
rect 2526 976 2532 977
rect 2582 980 2588 981
rect 2582 976 2583 980
rect 2587 976 2588 980
rect 1366 975 1372 976
rect 2582 975 2588 976
rect 110 971 116 972
rect 110 967 111 971
rect 115 967 116 971
rect 110 966 116 967
rect 1326 971 1332 972
rect 1326 967 1327 971
rect 1331 967 1332 971
rect 1326 966 1332 967
rect 112 947 114 966
rect 430 962 436 963
rect 430 958 431 962
rect 435 958 436 962
rect 430 957 436 958
rect 486 962 492 963
rect 486 958 487 962
rect 491 958 492 962
rect 486 957 492 958
rect 542 962 548 963
rect 542 958 543 962
rect 547 958 548 962
rect 542 957 548 958
rect 606 962 612 963
rect 606 958 607 962
rect 611 958 612 962
rect 606 957 612 958
rect 670 962 676 963
rect 670 958 671 962
rect 675 958 676 962
rect 670 957 676 958
rect 734 962 740 963
rect 734 958 735 962
rect 739 958 740 962
rect 734 957 740 958
rect 798 962 804 963
rect 798 958 799 962
rect 803 958 804 962
rect 798 957 804 958
rect 862 962 868 963
rect 862 958 863 962
rect 867 958 868 962
rect 862 957 868 958
rect 926 962 932 963
rect 926 958 927 962
rect 931 958 932 962
rect 926 957 932 958
rect 990 962 996 963
rect 990 958 991 962
rect 995 958 996 962
rect 990 957 996 958
rect 1054 962 1060 963
rect 1054 958 1055 962
rect 1059 958 1060 962
rect 1054 957 1060 958
rect 1118 962 1124 963
rect 1118 958 1119 962
rect 1123 958 1124 962
rect 1118 957 1124 958
rect 1174 962 1180 963
rect 1174 958 1175 962
rect 1179 958 1180 962
rect 1174 957 1180 958
rect 1230 962 1236 963
rect 1230 958 1231 962
rect 1235 958 1236 962
rect 1230 957 1236 958
rect 1286 962 1292 963
rect 1286 958 1287 962
rect 1291 958 1292 962
rect 1286 957 1292 958
rect 432 947 434 957
rect 488 947 490 957
rect 544 947 546 957
rect 608 947 610 957
rect 672 947 674 957
rect 736 947 738 957
rect 800 947 802 957
rect 864 947 866 957
rect 928 947 930 957
rect 992 947 994 957
rect 1056 947 1058 957
rect 1120 947 1122 957
rect 1176 947 1178 957
rect 1232 947 1234 957
rect 1288 947 1290 957
rect 1328 947 1330 966
rect 1366 963 1372 964
rect 1366 959 1367 963
rect 1371 959 1372 963
rect 1366 958 1372 959
rect 2582 963 2588 964
rect 2582 959 2583 963
rect 2587 959 2588 963
rect 2582 958 2588 959
rect 111 946 115 947
rect 111 941 115 942
rect 423 946 427 947
rect 423 941 427 942
rect 431 946 435 947
rect 431 941 435 942
rect 479 946 483 947
rect 479 941 483 942
rect 487 946 491 947
rect 487 941 491 942
rect 535 946 539 947
rect 535 941 539 942
rect 543 946 547 947
rect 543 941 547 942
rect 591 946 595 947
rect 591 941 595 942
rect 607 946 611 947
rect 607 941 611 942
rect 647 946 651 947
rect 647 941 651 942
rect 671 946 675 947
rect 671 941 675 942
rect 703 946 707 947
rect 703 941 707 942
rect 735 946 739 947
rect 735 941 739 942
rect 759 946 763 947
rect 759 941 763 942
rect 799 946 803 947
rect 799 941 803 942
rect 815 946 819 947
rect 815 941 819 942
rect 863 946 867 947
rect 863 941 867 942
rect 927 946 931 947
rect 927 941 931 942
rect 991 946 995 947
rect 991 941 995 942
rect 1055 946 1059 947
rect 1055 941 1059 942
rect 1119 946 1123 947
rect 1119 941 1123 942
rect 1175 946 1179 947
rect 1175 941 1179 942
rect 1231 946 1235 947
rect 1231 941 1235 942
rect 1287 946 1291 947
rect 1287 941 1291 942
rect 1327 946 1331 947
rect 1327 941 1331 942
rect 112 926 114 941
rect 424 935 426 941
rect 480 935 482 941
rect 536 935 538 941
rect 592 935 594 941
rect 648 935 650 941
rect 704 935 706 941
rect 760 935 762 941
rect 816 935 818 941
rect 422 934 428 935
rect 422 930 423 934
rect 427 930 428 934
rect 422 929 428 930
rect 478 934 484 935
rect 478 930 479 934
rect 483 930 484 934
rect 478 929 484 930
rect 534 934 540 935
rect 534 930 535 934
rect 539 930 540 934
rect 534 929 540 930
rect 590 934 596 935
rect 590 930 591 934
rect 595 930 596 934
rect 590 929 596 930
rect 646 934 652 935
rect 646 930 647 934
rect 651 930 652 934
rect 646 929 652 930
rect 702 934 708 935
rect 702 930 703 934
rect 707 930 708 934
rect 702 929 708 930
rect 758 934 764 935
rect 758 930 759 934
rect 763 930 764 934
rect 758 929 764 930
rect 814 934 820 935
rect 814 930 815 934
rect 819 930 820 934
rect 814 929 820 930
rect 1328 926 1330 941
rect 1368 935 1370 958
rect 1414 954 1420 955
rect 1414 950 1415 954
rect 1419 950 1420 954
rect 1414 949 1420 950
rect 1470 954 1476 955
rect 1470 950 1471 954
rect 1475 950 1476 954
rect 1470 949 1476 950
rect 1526 954 1532 955
rect 1526 950 1527 954
rect 1531 950 1532 954
rect 1526 949 1532 950
rect 1582 954 1588 955
rect 1582 950 1583 954
rect 1587 950 1588 954
rect 1582 949 1588 950
rect 1654 954 1660 955
rect 1654 950 1655 954
rect 1659 950 1660 954
rect 1654 949 1660 950
rect 1734 954 1740 955
rect 1734 950 1735 954
rect 1739 950 1740 954
rect 1734 949 1740 950
rect 1822 954 1828 955
rect 1822 950 1823 954
rect 1827 950 1828 954
rect 1822 949 1828 950
rect 1918 954 1924 955
rect 1918 950 1919 954
rect 1923 950 1924 954
rect 1918 949 1924 950
rect 2030 954 2036 955
rect 2030 950 2031 954
rect 2035 950 2036 954
rect 2030 949 2036 950
rect 2158 954 2164 955
rect 2158 950 2159 954
rect 2163 950 2164 954
rect 2158 949 2164 950
rect 2286 954 2292 955
rect 2286 950 2287 954
rect 2291 950 2292 954
rect 2286 949 2292 950
rect 2422 954 2428 955
rect 2422 950 2423 954
rect 2427 950 2428 954
rect 2422 949 2428 950
rect 2542 954 2548 955
rect 2542 950 2543 954
rect 2547 950 2548 954
rect 2542 949 2548 950
rect 1416 935 1418 949
rect 1472 935 1474 949
rect 1528 935 1530 949
rect 1584 935 1586 949
rect 1656 935 1658 949
rect 1736 935 1738 949
rect 1824 935 1826 949
rect 1920 935 1922 949
rect 2032 935 2034 949
rect 2160 935 2162 949
rect 2288 935 2290 949
rect 2424 935 2426 949
rect 2544 935 2546 949
rect 2584 935 2586 958
rect 1367 934 1371 935
rect 1367 929 1371 930
rect 1415 934 1419 935
rect 1415 929 1419 930
rect 1471 934 1475 935
rect 1471 929 1475 930
rect 1527 934 1531 935
rect 1527 929 1531 930
rect 1583 934 1587 935
rect 1583 929 1587 930
rect 1615 934 1619 935
rect 1615 929 1619 930
rect 1655 934 1659 935
rect 1655 929 1659 930
rect 1711 934 1715 935
rect 1711 929 1715 930
rect 1735 934 1739 935
rect 1735 929 1739 930
rect 1823 934 1827 935
rect 1823 929 1827 930
rect 1919 934 1923 935
rect 1919 929 1923 930
rect 1943 934 1947 935
rect 1943 929 1947 930
rect 2031 934 2035 935
rect 2031 929 2035 930
rect 2063 934 2067 935
rect 2063 929 2067 930
rect 2159 934 2163 935
rect 2159 929 2163 930
rect 2183 934 2187 935
rect 2183 929 2187 930
rect 2287 934 2291 935
rect 2287 929 2291 930
rect 2311 934 2315 935
rect 2311 929 2315 930
rect 2423 934 2427 935
rect 2423 929 2427 930
rect 2439 934 2443 935
rect 2439 929 2443 930
rect 2543 934 2547 935
rect 2543 929 2547 930
rect 2583 934 2587 935
rect 2583 929 2587 930
rect 110 925 116 926
rect 110 921 111 925
rect 115 921 116 925
rect 110 920 116 921
rect 1326 925 1332 926
rect 1326 921 1327 925
rect 1331 921 1332 925
rect 1326 920 1332 921
rect 1368 914 1370 929
rect 1416 923 1418 929
rect 1472 923 1474 929
rect 1528 923 1530 929
rect 1616 923 1618 929
rect 1712 923 1714 929
rect 1824 923 1826 929
rect 1944 923 1946 929
rect 2064 923 2066 929
rect 2184 923 2186 929
rect 2312 923 2314 929
rect 2440 923 2442 929
rect 2544 923 2546 929
rect 1414 922 1420 923
rect 1414 918 1415 922
rect 1419 918 1420 922
rect 1414 917 1420 918
rect 1470 922 1476 923
rect 1470 918 1471 922
rect 1475 918 1476 922
rect 1470 917 1476 918
rect 1526 922 1532 923
rect 1526 918 1527 922
rect 1531 918 1532 922
rect 1526 917 1532 918
rect 1614 922 1620 923
rect 1614 918 1615 922
rect 1619 918 1620 922
rect 1614 917 1620 918
rect 1710 922 1716 923
rect 1710 918 1711 922
rect 1715 918 1716 922
rect 1710 917 1716 918
rect 1822 922 1828 923
rect 1822 918 1823 922
rect 1827 918 1828 922
rect 1822 917 1828 918
rect 1942 922 1948 923
rect 1942 918 1943 922
rect 1947 918 1948 922
rect 1942 917 1948 918
rect 2062 922 2068 923
rect 2062 918 2063 922
rect 2067 918 2068 922
rect 2062 917 2068 918
rect 2182 922 2188 923
rect 2182 918 2183 922
rect 2187 918 2188 922
rect 2182 917 2188 918
rect 2310 922 2316 923
rect 2310 918 2311 922
rect 2315 918 2316 922
rect 2310 917 2316 918
rect 2438 922 2444 923
rect 2438 918 2439 922
rect 2443 918 2444 922
rect 2438 917 2444 918
rect 2542 922 2548 923
rect 2542 918 2543 922
rect 2547 918 2548 922
rect 2542 917 2548 918
rect 2584 914 2586 929
rect 1366 913 1372 914
rect 1366 909 1367 913
rect 1371 909 1372 913
rect 110 908 116 909
rect 1326 908 1332 909
rect 1366 908 1372 909
rect 2582 913 2588 914
rect 2582 909 2583 913
rect 2587 909 2588 913
rect 2582 908 2588 909
rect 110 904 111 908
rect 115 904 116 908
rect 110 903 116 904
rect 406 907 412 908
rect 406 903 407 907
rect 411 903 412 907
rect 112 891 114 903
rect 406 902 412 903
rect 462 907 468 908
rect 462 903 463 907
rect 467 903 468 907
rect 462 902 468 903
rect 518 907 524 908
rect 518 903 519 907
rect 523 903 524 907
rect 518 902 524 903
rect 574 907 580 908
rect 574 903 575 907
rect 579 903 580 907
rect 574 902 580 903
rect 630 907 636 908
rect 630 903 631 907
rect 635 903 636 907
rect 630 902 636 903
rect 686 907 692 908
rect 686 903 687 907
rect 691 903 692 907
rect 686 902 692 903
rect 742 907 748 908
rect 742 903 743 907
rect 747 903 748 907
rect 742 902 748 903
rect 798 907 804 908
rect 798 903 799 907
rect 803 903 804 907
rect 1326 904 1327 908
rect 1331 904 1332 908
rect 1326 903 1332 904
rect 798 902 804 903
rect 408 891 410 902
rect 464 891 466 902
rect 520 891 522 902
rect 576 891 578 902
rect 632 891 634 902
rect 688 891 690 902
rect 744 891 746 902
rect 800 891 802 902
rect 1328 891 1330 903
rect 1366 896 1372 897
rect 2582 896 2588 897
rect 1366 892 1367 896
rect 1371 892 1372 896
rect 1366 891 1372 892
rect 1398 895 1404 896
rect 1398 891 1399 895
rect 1403 891 1404 895
rect 111 890 115 891
rect 111 885 115 886
rect 279 890 283 891
rect 279 885 283 886
rect 335 890 339 891
rect 335 885 339 886
rect 391 890 395 891
rect 391 885 395 886
rect 407 890 411 891
rect 407 885 411 886
rect 455 890 459 891
rect 455 885 459 886
rect 463 890 467 891
rect 463 885 467 886
rect 519 890 523 891
rect 519 885 523 886
rect 575 890 579 891
rect 575 885 579 886
rect 583 890 587 891
rect 583 885 587 886
rect 631 890 635 891
rect 631 885 635 886
rect 647 890 651 891
rect 647 885 651 886
rect 687 890 691 891
rect 687 885 691 886
rect 711 890 715 891
rect 711 885 715 886
rect 743 890 747 891
rect 743 885 747 886
rect 775 890 779 891
rect 775 885 779 886
rect 799 890 803 891
rect 799 885 803 886
rect 847 890 851 891
rect 847 885 851 886
rect 919 890 923 891
rect 919 885 923 886
rect 1327 890 1331 891
rect 1327 885 1331 886
rect 112 873 114 885
rect 280 874 282 885
rect 336 874 338 885
rect 392 874 394 885
rect 456 874 458 885
rect 520 874 522 885
rect 584 874 586 885
rect 648 874 650 885
rect 712 874 714 885
rect 776 874 778 885
rect 848 874 850 885
rect 920 874 922 885
rect 278 873 284 874
rect 110 872 116 873
rect 110 868 111 872
rect 115 868 116 872
rect 278 869 279 873
rect 283 869 284 873
rect 278 868 284 869
rect 334 873 340 874
rect 334 869 335 873
rect 339 869 340 873
rect 334 868 340 869
rect 390 873 396 874
rect 390 869 391 873
rect 395 869 396 873
rect 390 868 396 869
rect 454 873 460 874
rect 454 869 455 873
rect 459 869 460 873
rect 454 868 460 869
rect 518 873 524 874
rect 518 869 519 873
rect 523 869 524 873
rect 518 868 524 869
rect 582 873 588 874
rect 582 869 583 873
rect 587 869 588 873
rect 582 868 588 869
rect 646 873 652 874
rect 646 869 647 873
rect 651 869 652 873
rect 646 868 652 869
rect 710 873 716 874
rect 710 869 711 873
rect 715 869 716 873
rect 710 868 716 869
rect 774 873 780 874
rect 774 869 775 873
rect 779 869 780 873
rect 774 868 780 869
rect 846 873 852 874
rect 846 869 847 873
rect 851 869 852 873
rect 846 868 852 869
rect 918 873 924 874
rect 1328 873 1330 885
rect 1368 879 1370 891
rect 1398 890 1404 891
rect 1454 895 1460 896
rect 1454 891 1455 895
rect 1459 891 1460 895
rect 1454 890 1460 891
rect 1510 895 1516 896
rect 1510 891 1511 895
rect 1515 891 1516 895
rect 1510 890 1516 891
rect 1598 895 1604 896
rect 1598 891 1599 895
rect 1603 891 1604 895
rect 1598 890 1604 891
rect 1694 895 1700 896
rect 1694 891 1695 895
rect 1699 891 1700 895
rect 1694 890 1700 891
rect 1806 895 1812 896
rect 1806 891 1807 895
rect 1811 891 1812 895
rect 1806 890 1812 891
rect 1926 895 1932 896
rect 1926 891 1927 895
rect 1931 891 1932 895
rect 1926 890 1932 891
rect 2046 895 2052 896
rect 2046 891 2047 895
rect 2051 891 2052 895
rect 2046 890 2052 891
rect 2166 895 2172 896
rect 2166 891 2167 895
rect 2171 891 2172 895
rect 2166 890 2172 891
rect 2294 895 2300 896
rect 2294 891 2295 895
rect 2299 891 2300 895
rect 2294 890 2300 891
rect 2422 895 2428 896
rect 2422 891 2423 895
rect 2427 891 2428 895
rect 2422 890 2428 891
rect 2526 895 2532 896
rect 2526 891 2527 895
rect 2531 891 2532 895
rect 2582 892 2583 896
rect 2587 892 2588 896
rect 2582 891 2588 892
rect 2526 890 2532 891
rect 1400 879 1402 890
rect 1456 879 1458 890
rect 1512 879 1514 890
rect 1600 879 1602 890
rect 1696 879 1698 890
rect 1808 879 1810 890
rect 1928 879 1930 890
rect 2048 879 2050 890
rect 2168 879 2170 890
rect 2296 879 2298 890
rect 2424 879 2426 890
rect 2528 879 2530 890
rect 2584 879 2586 891
rect 1367 878 1371 879
rect 1367 873 1371 874
rect 1399 878 1403 879
rect 1399 873 1403 874
rect 1455 878 1459 879
rect 1455 873 1459 874
rect 1471 878 1475 879
rect 1471 873 1475 874
rect 1511 878 1515 879
rect 1511 873 1515 874
rect 1551 878 1555 879
rect 1551 873 1555 874
rect 1599 878 1603 879
rect 1599 873 1603 874
rect 1639 878 1643 879
rect 1639 873 1643 874
rect 1695 878 1699 879
rect 1695 873 1699 874
rect 1727 878 1731 879
rect 1727 873 1731 874
rect 1807 878 1811 879
rect 1807 873 1811 874
rect 1815 878 1819 879
rect 1815 873 1819 874
rect 1903 878 1907 879
rect 1903 873 1907 874
rect 1927 878 1931 879
rect 1927 873 1931 874
rect 1991 878 1995 879
rect 1991 873 1995 874
rect 2047 878 2051 879
rect 2047 873 2051 874
rect 2071 878 2075 879
rect 2071 873 2075 874
rect 2143 878 2147 879
rect 2143 873 2147 874
rect 2167 878 2171 879
rect 2167 873 2171 874
rect 2215 878 2219 879
rect 2215 873 2219 874
rect 2279 878 2283 879
rect 2279 873 2283 874
rect 2295 878 2299 879
rect 2295 873 2299 874
rect 2343 878 2347 879
rect 2343 873 2347 874
rect 2407 878 2411 879
rect 2407 873 2411 874
rect 2423 878 2427 879
rect 2423 873 2427 874
rect 2471 878 2475 879
rect 2471 873 2475 874
rect 2527 878 2531 879
rect 2527 873 2531 874
rect 2583 878 2587 879
rect 2583 873 2587 874
rect 918 869 919 873
rect 923 869 924 873
rect 918 868 924 869
rect 1326 872 1332 873
rect 1326 868 1327 872
rect 1331 868 1332 872
rect 110 867 116 868
rect 1326 867 1332 868
rect 1368 861 1370 873
rect 1472 862 1474 873
rect 1552 862 1554 873
rect 1640 862 1642 873
rect 1728 862 1730 873
rect 1816 862 1818 873
rect 1904 862 1906 873
rect 1992 862 1994 873
rect 2072 862 2074 873
rect 2144 862 2146 873
rect 2216 862 2218 873
rect 2280 862 2282 873
rect 2344 862 2346 873
rect 2408 862 2410 873
rect 2472 862 2474 873
rect 2528 862 2530 873
rect 1470 861 1476 862
rect 1366 860 1372 861
rect 1366 856 1367 860
rect 1371 856 1372 860
rect 1470 857 1471 861
rect 1475 857 1476 861
rect 1470 856 1476 857
rect 1550 861 1556 862
rect 1550 857 1551 861
rect 1555 857 1556 861
rect 1550 856 1556 857
rect 1638 861 1644 862
rect 1638 857 1639 861
rect 1643 857 1644 861
rect 1638 856 1644 857
rect 1726 861 1732 862
rect 1726 857 1727 861
rect 1731 857 1732 861
rect 1726 856 1732 857
rect 1814 861 1820 862
rect 1814 857 1815 861
rect 1819 857 1820 861
rect 1814 856 1820 857
rect 1902 861 1908 862
rect 1902 857 1903 861
rect 1907 857 1908 861
rect 1902 856 1908 857
rect 1990 861 1996 862
rect 1990 857 1991 861
rect 1995 857 1996 861
rect 1990 856 1996 857
rect 2070 861 2076 862
rect 2070 857 2071 861
rect 2075 857 2076 861
rect 2070 856 2076 857
rect 2142 861 2148 862
rect 2142 857 2143 861
rect 2147 857 2148 861
rect 2142 856 2148 857
rect 2214 861 2220 862
rect 2214 857 2215 861
rect 2219 857 2220 861
rect 2214 856 2220 857
rect 2278 861 2284 862
rect 2278 857 2279 861
rect 2283 857 2284 861
rect 2278 856 2284 857
rect 2342 861 2348 862
rect 2342 857 2343 861
rect 2347 857 2348 861
rect 2342 856 2348 857
rect 2406 861 2412 862
rect 2406 857 2407 861
rect 2411 857 2412 861
rect 2406 856 2412 857
rect 2470 861 2476 862
rect 2470 857 2471 861
rect 2475 857 2476 861
rect 2470 856 2476 857
rect 2526 861 2532 862
rect 2584 861 2586 873
rect 2526 857 2527 861
rect 2531 857 2532 861
rect 2526 856 2532 857
rect 2582 860 2588 861
rect 2582 856 2583 860
rect 2587 856 2588 860
rect 110 855 116 856
rect 110 851 111 855
rect 115 851 116 855
rect 110 850 116 851
rect 1326 855 1332 856
rect 1366 855 1372 856
rect 2582 855 2588 856
rect 1326 851 1327 855
rect 1331 851 1332 855
rect 1326 850 1332 851
rect 112 827 114 850
rect 294 846 300 847
rect 294 842 295 846
rect 299 842 300 846
rect 294 841 300 842
rect 350 846 356 847
rect 350 842 351 846
rect 355 842 356 846
rect 350 841 356 842
rect 406 846 412 847
rect 406 842 407 846
rect 411 842 412 846
rect 406 841 412 842
rect 470 846 476 847
rect 470 842 471 846
rect 475 842 476 846
rect 470 841 476 842
rect 534 846 540 847
rect 534 842 535 846
rect 539 842 540 846
rect 534 841 540 842
rect 598 846 604 847
rect 598 842 599 846
rect 603 842 604 846
rect 598 841 604 842
rect 662 846 668 847
rect 662 842 663 846
rect 667 842 668 846
rect 662 841 668 842
rect 726 846 732 847
rect 726 842 727 846
rect 731 842 732 846
rect 726 841 732 842
rect 790 846 796 847
rect 790 842 791 846
rect 795 842 796 846
rect 790 841 796 842
rect 862 846 868 847
rect 862 842 863 846
rect 867 842 868 846
rect 862 841 868 842
rect 934 846 940 847
rect 934 842 935 846
rect 939 842 940 846
rect 934 841 940 842
rect 296 827 298 841
rect 352 827 354 841
rect 408 827 410 841
rect 472 827 474 841
rect 536 827 538 841
rect 600 827 602 841
rect 664 827 666 841
rect 728 827 730 841
rect 792 827 794 841
rect 864 827 866 841
rect 936 827 938 841
rect 1328 827 1330 850
rect 1366 843 1372 844
rect 1366 839 1367 843
rect 1371 839 1372 843
rect 1366 838 1372 839
rect 2582 843 2588 844
rect 2582 839 2583 843
rect 2587 839 2588 843
rect 2582 838 2588 839
rect 111 826 115 827
rect 111 821 115 822
rect 167 826 171 827
rect 167 821 171 822
rect 231 826 235 827
rect 231 821 235 822
rect 295 826 299 827
rect 295 821 299 822
rect 311 826 315 827
rect 311 821 315 822
rect 351 826 355 827
rect 351 821 355 822
rect 399 826 403 827
rect 399 821 403 822
rect 407 826 411 827
rect 407 821 411 822
rect 471 826 475 827
rect 471 821 475 822
rect 487 826 491 827
rect 487 821 491 822
rect 535 826 539 827
rect 535 821 539 822
rect 583 826 587 827
rect 583 821 587 822
rect 599 826 603 827
rect 599 821 603 822
rect 663 826 667 827
rect 663 821 667 822
rect 671 826 675 827
rect 671 821 675 822
rect 727 826 731 827
rect 727 821 731 822
rect 759 826 763 827
rect 759 821 763 822
rect 791 826 795 827
rect 791 821 795 822
rect 839 826 843 827
rect 839 821 843 822
rect 863 826 867 827
rect 863 821 867 822
rect 919 826 923 827
rect 919 821 923 822
rect 935 826 939 827
rect 935 821 939 822
rect 1007 826 1011 827
rect 1007 821 1011 822
rect 1095 826 1099 827
rect 1095 821 1099 822
rect 1327 826 1331 827
rect 1327 821 1331 822
rect 112 806 114 821
rect 168 815 170 821
rect 232 815 234 821
rect 312 815 314 821
rect 400 815 402 821
rect 488 815 490 821
rect 584 815 586 821
rect 672 815 674 821
rect 760 815 762 821
rect 840 815 842 821
rect 920 815 922 821
rect 1008 815 1010 821
rect 1096 815 1098 821
rect 166 814 172 815
rect 166 810 167 814
rect 171 810 172 814
rect 166 809 172 810
rect 230 814 236 815
rect 230 810 231 814
rect 235 810 236 814
rect 230 809 236 810
rect 310 814 316 815
rect 310 810 311 814
rect 315 810 316 814
rect 310 809 316 810
rect 398 814 404 815
rect 398 810 399 814
rect 403 810 404 814
rect 398 809 404 810
rect 486 814 492 815
rect 486 810 487 814
rect 491 810 492 814
rect 486 809 492 810
rect 582 814 588 815
rect 582 810 583 814
rect 587 810 588 814
rect 582 809 588 810
rect 670 814 676 815
rect 670 810 671 814
rect 675 810 676 814
rect 670 809 676 810
rect 758 814 764 815
rect 758 810 759 814
rect 763 810 764 814
rect 758 809 764 810
rect 838 814 844 815
rect 838 810 839 814
rect 843 810 844 814
rect 838 809 844 810
rect 918 814 924 815
rect 918 810 919 814
rect 923 810 924 814
rect 918 809 924 810
rect 1006 814 1012 815
rect 1006 810 1007 814
rect 1011 810 1012 814
rect 1006 809 1012 810
rect 1094 814 1100 815
rect 1094 810 1095 814
rect 1099 810 1100 814
rect 1094 809 1100 810
rect 1328 806 1330 821
rect 1368 815 1370 838
rect 1486 834 1492 835
rect 1486 830 1487 834
rect 1491 830 1492 834
rect 1486 829 1492 830
rect 1566 834 1572 835
rect 1566 830 1567 834
rect 1571 830 1572 834
rect 1566 829 1572 830
rect 1654 834 1660 835
rect 1654 830 1655 834
rect 1659 830 1660 834
rect 1654 829 1660 830
rect 1742 834 1748 835
rect 1742 830 1743 834
rect 1747 830 1748 834
rect 1742 829 1748 830
rect 1830 834 1836 835
rect 1830 830 1831 834
rect 1835 830 1836 834
rect 1830 829 1836 830
rect 1918 834 1924 835
rect 1918 830 1919 834
rect 1923 830 1924 834
rect 1918 829 1924 830
rect 2006 834 2012 835
rect 2006 830 2007 834
rect 2011 830 2012 834
rect 2006 829 2012 830
rect 2086 834 2092 835
rect 2086 830 2087 834
rect 2091 830 2092 834
rect 2086 829 2092 830
rect 2158 834 2164 835
rect 2158 830 2159 834
rect 2163 830 2164 834
rect 2158 829 2164 830
rect 2230 834 2236 835
rect 2230 830 2231 834
rect 2235 830 2236 834
rect 2230 829 2236 830
rect 2294 834 2300 835
rect 2294 830 2295 834
rect 2299 830 2300 834
rect 2294 829 2300 830
rect 2358 834 2364 835
rect 2358 830 2359 834
rect 2363 830 2364 834
rect 2358 829 2364 830
rect 2422 834 2428 835
rect 2422 830 2423 834
rect 2427 830 2428 834
rect 2422 829 2428 830
rect 2486 834 2492 835
rect 2486 830 2487 834
rect 2491 830 2492 834
rect 2486 829 2492 830
rect 2542 834 2548 835
rect 2542 830 2543 834
rect 2547 830 2548 834
rect 2542 829 2548 830
rect 1488 815 1490 829
rect 1568 815 1570 829
rect 1656 815 1658 829
rect 1744 815 1746 829
rect 1832 815 1834 829
rect 1920 815 1922 829
rect 2008 815 2010 829
rect 2088 815 2090 829
rect 2160 815 2162 829
rect 2232 815 2234 829
rect 2296 815 2298 829
rect 2360 815 2362 829
rect 2424 815 2426 829
rect 2488 815 2490 829
rect 2544 815 2546 829
rect 2584 815 2586 838
rect 1367 814 1371 815
rect 1367 809 1371 810
rect 1487 814 1491 815
rect 1487 809 1491 810
rect 1567 814 1571 815
rect 1567 809 1571 810
rect 1631 814 1635 815
rect 1631 809 1635 810
rect 1655 814 1659 815
rect 1655 809 1659 810
rect 1687 814 1691 815
rect 1687 809 1691 810
rect 1743 814 1747 815
rect 1743 809 1747 810
rect 1751 814 1755 815
rect 1751 809 1755 810
rect 1823 814 1827 815
rect 1823 809 1827 810
rect 1831 814 1835 815
rect 1831 809 1835 810
rect 1903 814 1907 815
rect 1903 809 1907 810
rect 1919 814 1923 815
rect 1919 809 1923 810
rect 1991 814 1995 815
rect 1991 809 1995 810
rect 2007 814 2011 815
rect 2007 809 2011 810
rect 2071 814 2075 815
rect 2071 809 2075 810
rect 2087 814 2091 815
rect 2087 809 2091 810
rect 2159 814 2163 815
rect 2159 809 2163 810
rect 2231 814 2235 815
rect 2231 809 2235 810
rect 2247 814 2251 815
rect 2247 809 2251 810
rect 2295 814 2299 815
rect 2295 809 2299 810
rect 2335 814 2339 815
rect 2335 809 2339 810
rect 2359 814 2363 815
rect 2359 809 2363 810
rect 2423 814 2427 815
rect 2423 809 2427 810
rect 2487 814 2491 815
rect 2487 809 2491 810
rect 2543 814 2547 815
rect 2543 809 2547 810
rect 2583 814 2587 815
rect 2583 809 2587 810
rect 110 805 116 806
rect 110 801 111 805
rect 115 801 116 805
rect 110 800 116 801
rect 1326 805 1332 806
rect 1326 801 1327 805
rect 1331 801 1332 805
rect 1326 800 1332 801
rect 1368 794 1370 809
rect 1632 803 1634 809
rect 1688 803 1690 809
rect 1752 803 1754 809
rect 1824 803 1826 809
rect 1904 803 1906 809
rect 1992 803 1994 809
rect 2072 803 2074 809
rect 2160 803 2162 809
rect 2248 803 2250 809
rect 2336 803 2338 809
rect 2424 803 2426 809
rect 1630 802 1636 803
rect 1630 798 1631 802
rect 1635 798 1636 802
rect 1630 797 1636 798
rect 1686 802 1692 803
rect 1686 798 1687 802
rect 1691 798 1692 802
rect 1686 797 1692 798
rect 1750 802 1756 803
rect 1750 798 1751 802
rect 1755 798 1756 802
rect 1750 797 1756 798
rect 1822 802 1828 803
rect 1822 798 1823 802
rect 1827 798 1828 802
rect 1822 797 1828 798
rect 1902 802 1908 803
rect 1902 798 1903 802
rect 1907 798 1908 802
rect 1902 797 1908 798
rect 1990 802 1996 803
rect 1990 798 1991 802
rect 1995 798 1996 802
rect 1990 797 1996 798
rect 2070 802 2076 803
rect 2070 798 2071 802
rect 2075 798 2076 802
rect 2070 797 2076 798
rect 2158 802 2164 803
rect 2158 798 2159 802
rect 2163 798 2164 802
rect 2158 797 2164 798
rect 2246 802 2252 803
rect 2246 798 2247 802
rect 2251 798 2252 802
rect 2246 797 2252 798
rect 2334 802 2340 803
rect 2334 798 2335 802
rect 2339 798 2340 802
rect 2334 797 2340 798
rect 2422 802 2428 803
rect 2422 798 2423 802
rect 2427 798 2428 802
rect 2422 797 2428 798
rect 2584 794 2586 809
rect 1366 793 1372 794
rect 1366 789 1367 793
rect 1371 789 1372 793
rect 110 788 116 789
rect 1326 788 1332 789
rect 1366 788 1372 789
rect 2582 793 2588 794
rect 2582 789 2583 793
rect 2587 789 2588 793
rect 2582 788 2588 789
rect 110 784 111 788
rect 115 784 116 788
rect 110 783 116 784
rect 150 787 156 788
rect 150 783 151 787
rect 155 783 156 787
rect 112 763 114 783
rect 150 782 156 783
rect 214 787 220 788
rect 214 783 215 787
rect 219 783 220 787
rect 214 782 220 783
rect 294 787 300 788
rect 294 783 295 787
rect 299 783 300 787
rect 294 782 300 783
rect 382 787 388 788
rect 382 783 383 787
rect 387 783 388 787
rect 382 782 388 783
rect 470 787 476 788
rect 470 783 471 787
rect 475 783 476 787
rect 470 782 476 783
rect 566 787 572 788
rect 566 783 567 787
rect 571 783 572 787
rect 566 782 572 783
rect 654 787 660 788
rect 654 783 655 787
rect 659 783 660 787
rect 654 782 660 783
rect 742 787 748 788
rect 742 783 743 787
rect 747 783 748 787
rect 742 782 748 783
rect 822 787 828 788
rect 822 783 823 787
rect 827 783 828 787
rect 822 782 828 783
rect 902 787 908 788
rect 902 783 903 787
rect 907 783 908 787
rect 902 782 908 783
rect 990 787 996 788
rect 990 783 991 787
rect 995 783 996 787
rect 990 782 996 783
rect 1078 787 1084 788
rect 1078 783 1079 787
rect 1083 783 1084 787
rect 1326 784 1327 788
rect 1331 784 1332 788
rect 1326 783 1332 784
rect 1078 782 1084 783
rect 152 763 154 782
rect 216 763 218 782
rect 296 763 298 782
rect 384 763 386 782
rect 472 763 474 782
rect 568 763 570 782
rect 656 763 658 782
rect 744 763 746 782
rect 824 763 826 782
rect 904 763 906 782
rect 992 763 994 782
rect 1080 763 1082 782
rect 1328 763 1330 783
rect 1366 776 1372 777
rect 2582 776 2588 777
rect 1366 772 1367 776
rect 1371 772 1372 776
rect 1366 771 1372 772
rect 1614 775 1620 776
rect 1614 771 1615 775
rect 1619 771 1620 775
rect 111 762 115 763
rect 111 757 115 758
rect 143 762 147 763
rect 143 757 147 758
rect 151 762 155 763
rect 151 757 155 758
rect 199 762 203 763
rect 199 757 203 758
rect 215 762 219 763
rect 215 757 219 758
rect 279 762 283 763
rect 279 757 283 758
rect 295 762 299 763
rect 295 757 299 758
rect 383 762 387 763
rect 383 757 387 758
rect 471 762 475 763
rect 471 757 475 758
rect 487 762 491 763
rect 487 757 491 758
rect 567 762 571 763
rect 567 757 571 758
rect 599 762 603 763
rect 599 757 603 758
rect 655 762 659 763
rect 655 757 659 758
rect 703 762 707 763
rect 703 757 707 758
rect 743 762 747 763
rect 743 757 747 758
rect 807 762 811 763
rect 807 757 811 758
rect 823 762 827 763
rect 823 757 827 758
rect 903 762 907 763
rect 903 757 907 758
rect 991 762 995 763
rect 991 757 995 758
rect 1079 762 1083 763
rect 1079 757 1083 758
rect 1175 762 1179 763
rect 1175 757 1179 758
rect 1327 762 1331 763
rect 1327 757 1331 758
rect 112 745 114 757
rect 144 746 146 757
rect 200 746 202 757
rect 280 746 282 757
rect 384 746 386 757
rect 488 746 490 757
rect 600 746 602 757
rect 704 746 706 757
rect 808 746 810 757
rect 904 746 906 757
rect 992 746 994 757
rect 1080 746 1082 757
rect 1176 746 1178 757
rect 142 745 148 746
rect 110 744 116 745
rect 110 740 111 744
rect 115 740 116 744
rect 142 741 143 745
rect 147 741 148 745
rect 142 740 148 741
rect 198 745 204 746
rect 198 741 199 745
rect 203 741 204 745
rect 198 740 204 741
rect 278 745 284 746
rect 278 741 279 745
rect 283 741 284 745
rect 278 740 284 741
rect 382 745 388 746
rect 382 741 383 745
rect 387 741 388 745
rect 382 740 388 741
rect 486 745 492 746
rect 486 741 487 745
rect 491 741 492 745
rect 486 740 492 741
rect 598 745 604 746
rect 598 741 599 745
rect 603 741 604 745
rect 598 740 604 741
rect 702 745 708 746
rect 702 741 703 745
rect 707 741 708 745
rect 702 740 708 741
rect 806 745 812 746
rect 806 741 807 745
rect 811 741 812 745
rect 806 740 812 741
rect 902 745 908 746
rect 902 741 903 745
rect 907 741 908 745
rect 902 740 908 741
rect 990 745 996 746
rect 990 741 991 745
rect 995 741 996 745
rect 990 740 996 741
rect 1078 745 1084 746
rect 1078 741 1079 745
rect 1083 741 1084 745
rect 1078 740 1084 741
rect 1174 745 1180 746
rect 1328 745 1330 757
rect 1368 755 1370 771
rect 1614 770 1620 771
rect 1670 775 1676 776
rect 1670 771 1671 775
rect 1675 771 1676 775
rect 1670 770 1676 771
rect 1734 775 1740 776
rect 1734 771 1735 775
rect 1739 771 1740 775
rect 1734 770 1740 771
rect 1806 775 1812 776
rect 1806 771 1807 775
rect 1811 771 1812 775
rect 1806 770 1812 771
rect 1886 775 1892 776
rect 1886 771 1887 775
rect 1891 771 1892 775
rect 1886 770 1892 771
rect 1974 775 1980 776
rect 1974 771 1975 775
rect 1979 771 1980 775
rect 1974 770 1980 771
rect 2054 775 2060 776
rect 2054 771 2055 775
rect 2059 771 2060 775
rect 2054 770 2060 771
rect 2142 775 2148 776
rect 2142 771 2143 775
rect 2147 771 2148 775
rect 2142 770 2148 771
rect 2230 775 2236 776
rect 2230 771 2231 775
rect 2235 771 2236 775
rect 2230 770 2236 771
rect 2318 775 2324 776
rect 2318 771 2319 775
rect 2323 771 2324 775
rect 2318 770 2324 771
rect 2406 775 2412 776
rect 2406 771 2407 775
rect 2411 771 2412 775
rect 2582 772 2583 776
rect 2587 772 2588 776
rect 2582 771 2588 772
rect 2406 770 2412 771
rect 1616 755 1618 770
rect 1672 755 1674 770
rect 1736 755 1738 770
rect 1808 755 1810 770
rect 1888 755 1890 770
rect 1976 755 1978 770
rect 2056 755 2058 770
rect 2144 755 2146 770
rect 2232 755 2234 770
rect 2320 755 2322 770
rect 2408 755 2410 770
rect 2584 755 2586 771
rect 1367 754 1371 755
rect 1367 749 1371 750
rect 1567 754 1571 755
rect 1567 749 1571 750
rect 1615 754 1619 755
rect 1615 749 1619 750
rect 1623 754 1627 755
rect 1623 749 1627 750
rect 1671 754 1675 755
rect 1671 749 1675 750
rect 1687 754 1691 755
rect 1687 749 1691 750
rect 1735 754 1739 755
rect 1735 749 1739 750
rect 1759 754 1763 755
rect 1759 749 1763 750
rect 1807 754 1811 755
rect 1807 749 1811 750
rect 1839 754 1843 755
rect 1839 749 1843 750
rect 1887 754 1891 755
rect 1887 749 1891 750
rect 1919 754 1923 755
rect 1919 749 1923 750
rect 1975 754 1979 755
rect 1975 749 1979 750
rect 1999 754 2003 755
rect 1999 749 2003 750
rect 2055 754 2059 755
rect 2055 749 2059 750
rect 2079 754 2083 755
rect 2079 749 2083 750
rect 2143 754 2147 755
rect 2143 749 2147 750
rect 2159 754 2163 755
rect 2159 749 2163 750
rect 2231 754 2235 755
rect 2231 749 2235 750
rect 2247 754 2251 755
rect 2247 749 2251 750
rect 2319 754 2323 755
rect 2319 749 2323 750
rect 2335 754 2339 755
rect 2335 749 2339 750
rect 2407 754 2411 755
rect 2407 749 2411 750
rect 2583 754 2587 755
rect 2583 749 2587 750
rect 1174 741 1175 745
rect 1179 741 1180 745
rect 1174 740 1180 741
rect 1326 744 1332 745
rect 1326 740 1327 744
rect 1331 740 1332 744
rect 110 739 116 740
rect 1326 739 1332 740
rect 1368 737 1370 749
rect 1568 738 1570 749
rect 1624 738 1626 749
rect 1688 738 1690 749
rect 1760 738 1762 749
rect 1840 738 1842 749
rect 1920 738 1922 749
rect 2000 738 2002 749
rect 2080 738 2082 749
rect 2160 738 2162 749
rect 2248 738 2250 749
rect 2336 738 2338 749
rect 1566 737 1572 738
rect 1366 736 1372 737
rect 1366 732 1367 736
rect 1371 732 1372 736
rect 1566 733 1567 737
rect 1571 733 1572 737
rect 1566 732 1572 733
rect 1622 737 1628 738
rect 1622 733 1623 737
rect 1627 733 1628 737
rect 1622 732 1628 733
rect 1686 737 1692 738
rect 1686 733 1687 737
rect 1691 733 1692 737
rect 1686 732 1692 733
rect 1758 737 1764 738
rect 1758 733 1759 737
rect 1763 733 1764 737
rect 1758 732 1764 733
rect 1838 737 1844 738
rect 1838 733 1839 737
rect 1843 733 1844 737
rect 1838 732 1844 733
rect 1918 737 1924 738
rect 1918 733 1919 737
rect 1923 733 1924 737
rect 1918 732 1924 733
rect 1998 737 2004 738
rect 1998 733 1999 737
rect 2003 733 2004 737
rect 1998 732 2004 733
rect 2078 737 2084 738
rect 2078 733 2079 737
rect 2083 733 2084 737
rect 2078 732 2084 733
rect 2158 737 2164 738
rect 2158 733 2159 737
rect 2163 733 2164 737
rect 2158 732 2164 733
rect 2246 737 2252 738
rect 2246 733 2247 737
rect 2251 733 2252 737
rect 2246 732 2252 733
rect 2334 737 2340 738
rect 2584 737 2586 749
rect 2334 733 2335 737
rect 2339 733 2340 737
rect 2334 732 2340 733
rect 2582 736 2588 737
rect 2582 732 2583 736
rect 2587 732 2588 736
rect 1366 731 1372 732
rect 2582 731 2588 732
rect 110 727 116 728
rect 110 723 111 727
rect 115 723 116 727
rect 110 722 116 723
rect 1326 727 1332 728
rect 1326 723 1327 727
rect 1331 723 1332 727
rect 1326 722 1332 723
rect 112 703 114 722
rect 158 718 164 719
rect 158 714 159 718
rect 163 714 164 718
rect 158 713 164 714
rect 214 718 220 719
rect 214 714 215 718
rect 219 714 220 718
rect 214 713 220 714
rect 294 718 300 719
rect 294 714 295 718
rect 299 714 300 718
rect 294 713 300 714
rect 398 718 404 719
rect 398 714 399 718
rect 403 714 404 718
rect 398 713 404 714
rect 502 718 508 719
rect 502 714 503 718
rect 507 714 508 718
rect 502 713 508 714
rect 614 718 620 719
rect 614 714 615 718
rect 619 714 620 718
rect 614 713 620 714
rect 718 718 724 719
rect 718 714 719 718
rect 723 714 724 718
rect 718 713 724 714
rect 822 718 828 719
rect 822 714 823 718
rect 827 714 828 718
rect 822 713 828 714
rect 918 718 924 719
rect 918 714 919 718
rect 923 714 924 718
rect 918 713 924 714
rect 1006 718 1012 719
rect 1006 714 1007 718
rect 1011 714 1012 718
rect 1006 713 1012 714
rect 1094 718 1100 719
rect 1094 714 1095 718
rect 1099 714 1100 718
rect 1094 713 1100 714
rect 1190 718 1196 719
rect 1190 714 1191 718
rect 1195 714 1196 718
rect 1190 713 1196 714
rect 160 703 162 713
rect 216 703 218 713
rect 296 703 298 713
rect 400 703 402 713
rect 504 703 506 713
rect 616 703 618 713
rect 720 703 722 713
rect 824 703 826 713
rect 920 703 922 713
rect 1008 703 1010 713
rect 1096 703 1098 713
rect 1192 703 1194 713
rect 1328 703 1330 722
rect 1366 719 1372 720
rect 1366 715 1367 719
rect 1371 715 1372 719
rect 1366 714 1372 715
rect 2582 719 2588 720
rect 2582 715 2583 719
rect 2587 715 2588 719
rect 2582 714 2588 715
rect 111 702 115 703
rect 111 697 115 698
rect 159 702 163 703
rect 159 697 163 698
rect 215 702 219 703
rect 215 697 219 698
rect 279 702 283 703
rect 279 697 283 698
rect 295 702 299 703
rect 295 697 299 698
rect 359 702 363 703
rect 359 697 363 698
rect 399 702 403 703
rect 399 697 403 698
rect 447 702 451 703
rect 447 697 451 698
rect 503 702 507 703
rect 503 697 507 698
rect 535 702 539 703
rect 535 697 539 698
rect 615 702 619 703
rect 615 697 619 698
rect 623 702 627 703
rect 623 697 627 698
rect 711 702 715 703
rect 711 697 715 698
rect 719 702 723 703
rect 719 697 723 698
rect 791 702 795 703
rect 791 697 795 698
rect 823 702 827 703
rect 823 697 827 698
rect 871 702 875 703
rect 871 697 875 698
rect 919 702 923 703
rect 919 697 923 698
rect 951 702 955 703
rect 951 697 955 698
rect 1007 702 1011 703
rect 1007 697 1011 698
rect 1039 702 1043 703
rect 1039 697 1043 698
rect 1095 702 1099 703
rect 1095 697 1099 698
rect 1191 702 1195 703
rect 1191 697 1195 698
rect 1327 702 1331 703
rect 1327 697 1331 698
rect 112 682 114 697
rect 160 691 162 697
rect 216 691 218 697
rect 280 691 282 697
rect 360 691 362 697
rect 448 691 450 697
rect 536 691 538 697
rect 624 691 626 697
rect 712 691 714 697
rect 792 691 794 697
rect 872 691 874 697
rect 952 691 954 697
rect 1040 691 1042 697
rect 158 690 164 691
rect 158 686 159 690
rect 163 686 164 690
rect 158 685 164 686
rect 214 690 220 691
rect 214 686 215 690
rect 219 686 220 690
rect 214 685 220 686
rect 278 690 284 691
rect 278 686 279 690
rect 283 686 284 690
rect 278 685 284 686
rect 358 690 364 691
rect 358 686 359 690
rect 363 686 364 690
rect 358 685 364 686
rect 446 690 452 691
rect 446 686 447 690
rect 451 686 452 690
rect 446 685 452 686
rect 534 690 540 691
rect 534 686 535 690
rect 539 686 540 690
rect 534 685 540 686
rect 622 690 628 691
rect 622 686 623 690
rect 627 686 628 690
rect 622 685 628 686
rect 710 690 716 691
rect 710 686 711 690
rect 715 686 716 690
rect 710 685 716 686
rect 790 690 796 691
rect 790 686 791 690
rect 795 686 796 690
rect 790 685 796 686
rect 870 690 876 691
rect 870 686 871 690
rect 875 686 876 690
rect 870 685 876 686
rect 950 690 956 691
rect 950 686 951 690
rect 955 686 956 690
rect 950 685 956 686
rect 1038 690 1044 691
rect 1038 686 1039 690
rect 1043 686 1044 690
rect 1038 685 1044 686
rect 1328 682 1330 697
rect 1368 695 1370 714
rect 1582 710 1588 711
rect 1582 706 1583 710
rect 1587 706 1588 710
rect 1582 705 1588 706
rect 1638 710 1644 711
rect 1638 706 1639 710
rect 1643 706 1644 710
rect 1638 705 1644 706
rect 1702 710 1708 711
rect 1702 706 1703 710
rect 1707 706 1708 710
rect 1702 705 1708 706
rect 1774 710 1780 711
rect 1774 706 1775 710
rect 1779 706 1780 710
rect 1774 705 1780 706
rect 1854 710 1860 711
rect 1854 706 1855 710
rect 1859 706 1860 710
rect 1854 705 1860 706
rect 1934 710 1940 711
rect 1934 706 1935 710
rect 1939 706 1940 710
rect 1934 705 1940 706
rect 2014 710 2020 711
rect 2014 706 2015 710
rect 2019 706 2020 710
rect 2014 705 2020 706
rect 2094 710 2100 711
rect 2094 706 2095 710
rect 2099 706 2100 710
rect 2094 705 2100 706
rect 2174 710 2180 711
rect 2174 706 2175 710
rect 2179 706 2180 710
rect 2174 705 2180 706
rect 2262 710 2268 711
rect 2262 706 2263 710
rect 2267 706 2268 710
rect 2262 705 2268 706
rect 2350 710 2356 711
rect 2350 706 2351 710
rect 2355 706 2356 710
rect 2350 705 2356 706
rect 1584 695 1586 705
rect 1640 695 1642 705
rect 1704 695 1706 705
rect 1776 695 1778 705
rect 1856 695 1858 705
rect 1936 695 1938 705
rect 2016 695 2018 705
rect 2096 695 2098 705
rect 2176 695 2178 705
rect 2264 695 2266 705
rect 2352 695 2354 705
rect 2584 695 2586 714
rect 1367 694 1371 695
rect 1367 689 1371 690
rect 1415 694 1419 695
rect 1415 689 1419 690
rect 1511 694 1515 695
rect 1511 689 1515 690
rect 1583 694 1587 695
rect 1583 689 1587 690
rect 1615 694 1619 695
rect 1615 689 1619 690
rect 1639 694 1643 695
rect 1639 689 1643 690
rect 1703 694 1707 695
rect 1703 689 1707 690
rect 1719 694 1723 695
rect 1719 689 1723 690
rect 1775 694 1779 695
rect 1775 689 1779 690
rect 1823 694 1827 695
rect 1823 689 1827 690
rect 1855 694 1859 695
rect 1855 689 1859 690
rect 1927 694 1931 695
rect 1927 689 1931 690
rect 1935 694 1939 695
rect 1935 689 1939 690
rect 2015 694 2019 695
rect 2015 689 2019 690
rect 2023 694 2027 695
rect 2023 689 2027 690
rect 2095 694 2099 695
rect 2095 689 2099 690
rect 2119 694 2123 695
rect 2119 689 2123 690
rect 2175 694 2179 695
rect 2175 689 2179 690
rect 2207 694 2211 695
rect 2207 689 2211 690
rect 2263 694 2267 695
rect 2263 689 2267 690
rect 2295 694 2299 695
rect 2295 689 2299 690
rect 2351 694 2355 695
rect 2351 689 2355 690
rect 2391 694 2395 695
rect 2391 689 2395 690
rect 2583 694 2587 695
rect 2583 689 2587 690
rect 110 681 116 682
rect 110 677 111 681
rect 115 677 116 681
rect 110 676 116 677
rect 1326 681 1332 682
rect 1326 677 1327 681
rect 1331 677 1332 681
rect 1326 676 1332 677
rect 1368 674 1370 689
rect 1416 683 1418 689
rect 1512 683 1514 689
rect 1616 683 1618 689
rect 1720 683 1722 689
rect 1824 683 1826 689
rect 1928 683 1930 689
rect 2024 683 2026 689
rect 2120 683 2122 689
rect 2208 683 2210 689
rect 2296 683 2298 689
rect 2392 683 2394 689
rect 1414 682 1420 683
rect 1414 678 1415 682
rect 1419 678 1420 682
rect 1414 677 1420 678
rect 1510 682 1516 683
rect 1510 678 1511 682
rect 1515 678 1516 682
rect 1510 677 1516 678
rect 1614 682 1620 683
rect 1614 678 1615 682
rect 1619 678 1620 682
rect 1614 677 1620 678
rect 1718 682 1724 683
rect 1718 678 1719 682
rect 1723 678 1724 682
rect 1718 677 1724 678
rect 1822 682 1828 683
rect 1822 678 1823 682
rect 1827 678 1828 682
rect 1822 677 1828 678
rect 1926 682 1932 683
rect 1926 678 1927 682
rect 1931 678 1932 682
rect 1926 677 1932 678
rect 2022 682 2028 683
rect 2022 678 2023 682
rect 2027 678 2028 682
rect 2022 677 2028 678
rect 2118 682 2124 683
rect 2118 678 2119 682
rect 2123 678 2124 682
rect 2118 677 2124 678
rect 2206 682 2212 683
rect 2206 678 2207 682
rect 2211 678 2212 682
rect 2206 677 2212 678
rect 2294 682 2300 683
rect 2294 678 2295 682
rect 2299 678 2300 682
rect 2294 677 2300 678
rect 2390 682 2396 683
rect 2390 678 2391 682
rect 2395 678 2396 682
rect 2390 677 2396 678
rect 2584 674 2586 689
rect 1366 673 1372 674
rect 1366 669 1367 673
rect 1371 669 1372 673
rect 1366 668 1372 669
rect 2582 673 2588 674
rect 2582 669 2583 673
rect 2587 669 2588 673
rect 2582 668 2588 669
rect 110 664 116 665
rect 1326 664 1332 665
rect 110 660 111 664
rect 115 660 116 664
rect 110 659 116 660
rect 142 663 148 664
rect 142 659 143 663
rect 147 659 148 663
rect 112 639 114 659
rect 142 658 148 659
rect 198 663 204 664
rect 198 659 199 663
rect 203 659 204 663
rect 198 658 204 659
rect 262 663 268 664
rect 262 659 263 663
rect 267 659 268 663
rect 262 658 268 659
rect 342 663 348 664
rect 342 659 343 663
rect 347 659 348 663
rect 342 658 348 659
rect 430 663 436 664
rect 430 659 431 663
rect 435 659 436 663
rect 430 658 436 659
rect 518 663 524 664
rect 518 659 519 663
rect 523 659 524 663
rect 518 658 524 659
rect 606 663 612 664
rect 606 659 607 663
rect 611 659 612 663
rect 606 658 612 659
rect 694 663 700 664
rect 694 659 695 663
rect 699 659 700 663
rect 694 658 700 659
rect 774 663 780 664
rect 774 659 775 663
rect 779 659 780 663
rect 774 658 780 659
rect 854 663 860 664
rect 854 659 855 663
rect 859 659 860 663
rect 854 658 860 659
rect 934 663 940 664
rect 934 659 935 663
rect 939 659 940 663
rect 934 658 940 659
rect 1022 663 1028 664
rect 1022 659 1023 663
rect 1027 659 1028 663
rect 1326 660 1327 664
rect 1331 660 1332 664
rect 1326 659 1332 660
rect 1022 658 1028 659
rect 144 639 146 658
rect 200 639 202 658
rect 264 639 266 658
rect 344 639 346 658
rect 432 639 434 658
rect 520 639 522 658
rect 608 639 610 658
rect 696 639 698 658
rect 776 639 778 658
rect 856 639 858 658
rect 936 639 938 658
rect 1024 639 1026 658
rect 1328 639 1330 659
rect 1366 656 1372 657
rect 2582 656 2588 657
rect 1366 652 1367 656
rect 1371 652 1372 656
rect 1366 651 1372 652
rect 1398 655 1404 656
rect 1398 651 1399 655
rect 1403 651 1404 655
rect 1368 639 1370 651
rect 1398 650 1404 651
rect 1494 655 1500 656
rect 1494 651 1495 655
rect 1499 651 1500 655
rect 1494 650 1500 651
rect 1598 655 1604 656
rect 1598 651 1599 655
rect 1603 651 1604 655
rect 1598 650 1604 651
rect 1702 655 1708 656
rect 1702 651 1703 655
rect 1707 651 1708 655
rect 1702 650 1708 651
rect 1806 655 1812 656
rect 1806 651 1807 655
rect 1811 651 1812 655
rect 1806 650 1812 651
rect 1910 655 1916 656
rect 1910 651 1911 655
rect 1915 651 1916 655
rect 1910 650 1916 651
rect 2006 655 2012 656
rect 2006 651 2007 655
rect 2011 651 2012 655
rect 2006 650 2012 651
rect 2102 655 2108 656
rect 2102 651 2103 655
rect 2107 651 2108 655
rect 2102 650 2108 651
rect 2190 655 2196 656
rect 2190 651 2191 655
rect 2195 651 2196 655
rect 2190 650 2196 651
rect 2278 655 2284 656
rect 2278 651 2279 655
rect 2283 651 2284 655
rect 2278 650 2284 651
rect 2374 655 2380 656
rect 2374 651 2375 655
rect 2379 651 2380 655
rect 2582 652 2583 656
rect 2587 652 2588 656
rect 2582 651 2588 652
rect 2374 650 2380 651
rect 1400 639 1402 650
rect 1496 639 1498 650
rect 1600 639 1602 650
rect 1704 639 1706 650
rect 1808 639 1810 650
rect 1912 639 1914 650
rect 2008 639 2010 650
rect 2104 639 2106 650
rect 2192 639 2194 650
rect 2280 639 2282 650
rect 2376 639 2378 650
rect 2584 639 2586 651
rect 111 638 115 639
rect 111 633 115 634
rect 143 638 147 639
rect 143 633 147 634
rect 199 638 203 639
rect 199 633 203 634
rect 255 638 259 639
rect 255 633 259 634
rect 263 638 267 639
rect 263 633 267 634
rect 311 638 315 639
rect 311 633 315 634
rect 343 638 347 639
rect 343 633 347 634
rect 391 638 395 639
rect 391 633 395 634
rect 431 638 435 639
rect 431 633 435 634
rect 479 638 483 639
rect 479 633 483 634
rect 519 638 523 639
rect 519 633 523 634
rect 575 638 579 639
rect 575 633 579 634
rect 607 638 611 639
rect 607 633 611 634
rect 679 638 683 639
rect 679 633 683 634
rect 695 638 699 639
rect 695 633 699 634
rect 775 638 779 639
rect 775 633 779 634
rect 783 638 787 639
rect 783 633 787 634
rect 855 638 859 639
rect 855 633 859 634
rect 887 638 891 639
rect 887 633 891 634
rect 935 638 939 639
rect 935 633 939 634
rect 991 638 995 639
rect 991 633 995 634
rect 1023 638 1027 639
rect 1023 633 1027 634
rect 1087 638 1091 639
rect 1087 633 1091 634
rect 1191 638 1195 639
rect 1191 633 1195 634
rect 1271 638 1275 639
rect 1271 633 1275 634
rect 1327 638 1331 639
rect 1327 633 1331 634
rect 1367 638 1371 639
rect 1367 633 1371 634
rect 1399 638 1403 639
rect 1399 633 1403 634
rect 1495 638 1499 639
rect 1495 633 1499 634
rect 1511 638 1515 639
rect 1511 633 1515 634
rect 1599 638 1603 639
rect 1599 633 1603 634
rect 1647 638 1651 639
rect 1647 633 1651 634
rect 1703 638 1707 639
rect 1703 633 1707 634
rect 1783 638 1787 639
rect 1783 633 1787 634
rect 1807 638 1811 639
rect 1807 633 1811 634
rect 1911 638 1915 639
rect 1911 633 1915 634
rect 2007 638 2011 639
rect 2007 633 2011 634
rect 2039 638 2043 639
rect 2039 633 2043 634
rect 2103 638 2107 639
rect 2103 633 2107 634
rect 2159 638 2163 639
rect 2159 633 2163 634
rect 2191 638 2195 639
rect 2191 633 2195 634
rect 2279 638 2283 639
rect 2279 633 2283 634
rect 2375 638 2379 639
rect 2375 633 2379 634
rect 2407 638 2411 639
rect 2407 633 2411 634
rect 2583 638 2587 639
rect 2583 633 2587 634
rect 112 621 114 633
rect 144 622 146 633
rect 200 622 202 633
rect 256 622 258 633
rect 312 622 314 633
rect 392 622 394 633
rect 480 622 482 633
rect 576 622 578 633
rect 680 622 682 633
rect 784 622 786 633
rect 888 622 890 633
rect 992 622 994 633
rect 1088 622 1090 633
rect 1192 622 1194 633
rect 1272 622 1274 633
rect 142 621 148 622
rect 110 620 116 621
rect 110 616 111 620
rect 115 616 116 620
rect 142 617 143 621
rect 147 617 148 621
rect 142 616 148 617
rect 198 621 204 622
rect 198 617 199 621
rect 203 617 204 621
rect 198 616 204 617
rect 254 621 260 622
rect 254 617 255 621
rect 259 617 260 621
rect 254 616 260 617
rect 310 621 316 622
rect 310 617 311 621
rect 315 617 316 621
rect 310 616 316 617
rect 390 621 396 622
rect 390 617 391 621
rect 395 617 396 621
rect 390 616 396 617
rect 478 621 484 622
rect 478 617 479 621
rect 483 617 484 621
rect 478 616 484 617
rect 574 621 580 622
rect 574 617 575 621
rect 579 617 580 621
rect 574 616 580 617
rect 678 621 684 622
rect 678 617 679 621
rect 683 617 684 621
rect 678 616 684 617
rect 782 621 788 622
rect 782 617 783 621
rect 787 617 788 621
rect 782 616 788 617
rect 886 621 892 622
rect 886 617 887 621
rect 891 617 892 621
rect 886 616 892 617
rect 990 621 996 622
rect 990 617 991 621
rect 995 617 996 621
rect 990 616 996 617
rect 1086 621 1092 622
rect 1086 617 1087 621
rect 1091 617 1092 621
rect 1086 616 1092 617
rect 1190 621 1196 622
rect 1190 617 1191 621
rect 1195 617 1196 621
rect 1190 616 1196 617
rect 1270 621 1276 622
rect 1328 621 1330 633
rect 1368 621 1370 633
rect 1400 622 1402 633
rect 1512 622 1514 633
rect 1648 622 1650 633
rect 1784 622 1786 633
rect 1912 622 1914 633
rect 2040 622 2042 633
rect 2160 622 2162 633
rect 2280 622 2282 633
rect 2408 622 2410 633
rect 1398 621 1404 622
rect 1270 617 1271 621
rect 1275 617 1276 621
rect 1270 616 1276 617
rect 1326 620 1332 621
rect 1326 616 1327 620
rect 1331 616 1332 620
rect 110 615 116 616
rect 1326 615 1332 616
rect 1366 620 1372 621
rect 1366 616 1367 620
rect 1371 616 1372 620
rect 1398 617 1399 621
rect 1403 617 1404 621
rect 1398 616 1404 617
rect 1510 621 1516 622
rect 1510 617 1511 621
rect 1515 617 1516 621
rect 1510 616 1516 617
rect 1646 621 1652 622
rect 1646 617 1647 621
rect 1651 617 1652 621
rect 1646 616 1652 617
rect 1782 621 1788 622
rect 1782 617 1783 621
rect 1787 617 1788 621
rect 1782 616 1788 617
rect 1910 621 1916 622
rect 1910 617 1911 621
rect 1915 617 1916 621
rect 1910 616 1916 617
rect 2038 621 2044 622
rect 2038 617 2039 621
rect 2043 617 2044 621
rect 2038 616 2044 617
rect 2158 621 2164 622
rect 2158 617 2159 621
rect 2163 617 2164 621
rect 2158 616 2164 617
rect 2278 621 2284 622
rect 2278 617 2279 621
rect 2283 617 2284 621
rect 2278 616 2284 617
rect 2406 621 2412 622
rect 2584 621 2586 633
rect 2406 617 2407 621
rect 2411 617 2412 621
rect 2406 616 2412 617
rect 2582 620 2588 621
rect 2582 616 2583 620
rect 2587 616 2588 620
rect 1366 615 1372 616
rect 2582 615 2588 616
rect 110 603 116 604
rect 110 599 111 603
rect 115 599 116 603
rect 110 598 116 599
rect 1326 603 1332 604
rect 1326 599 1327 603
rect 1331 599 1332 603
rect 1326 598 1332 599
rect 1366 603 1372 604
rect 1366 599 1367 603
rect 1371 599 1372 603
rect 1366 598 1372 599
rect 2582 603 2588 604
rect 2582 599 2583 603
rect 2587 599 2588 603
rect 2582 598 2588 599
rect 112 579 114 598
rect 158 594 164 595
rect 158 590 159 594
rect 163 590 164 594
rect 158 589 164 590
rect 214 594 220 595
rect 214 590 215 594
rect 219 590 220 594
rect 214 589 220 590
rect 270 594 276 595
rect 270 590 271 594
rect 275 590 276 594
rect 270 589 276 590
rect 326 594 332 595
rect 326 590 327 594
rect 331 590 332 594
rect 326 589 332 590
rect 406 594 412 595
rect 406 590 407 594
rect 411 590 412 594
rect 406 589 412 590
rect 494 594 500 595
rect 494 590 495 594
rect 499 590 500 594
rect 494 589 500 590
rect 590 594 596 595
rect 590 590 591 594
rect 595 590 596 594
rect 590 589 596 590
rect 694 594 700 595
rect 694 590 695 594
rect 699 590 700 594
rect 694 589 700 590
rect 798 594 804 595
rect 798 590 799 594
rect 803 590 804 594
rect 798 589 804 590
rect 902 594 908 595
rect 902 590 903 594
rect 907 590 908 594
rect 902 589 908 590
rect 1006 594 1012 595
rect 1006 590 1007 594
rect 1011 590 1012 594
rect 1006 589 1012 590
rect 1102 594 1108 595
rect 1102 590 1103 594
rect 1107 590 1108 594
rect 1102 589 1108 590
rect 1206 594 1212 595
rect 1206 590 1207 594
rect 1211 590 1212 594
rect 1206 589 1212 590
rect 1286 594 1292 595
rect 1286 590 1287 594
rect 1291 590 1292 594
rect 1286 589 1292 590
rect 160 579 162 589
rect 216 579 218 589
rect 272 579 274 589
rect 328 579 330 589
rect 408 579 410 589
rect 496 579 498 589
rect 592 579 594 589
rect 696 579 698 589
rect 800 579 802 589
rect 904 579 906 589
rect 1008 579 1010 589
rect 1104 579 1106 589
rect 1208 579 1210 589
rect 1288 579 1290 589
rect 1328 579 1330 598
rect 111 578 115 579
rect 111 573 115 574
rect 159 578 163 579
rect 159 573 163 574
rect 199 578 203 579
rect 199 573 203 574
rect 215 578 219 579
rect 215 573 219 574
rect 263 578 267 579
rect 263 573 267 574
rect 271 578 275 579
rect 271 573 275 574
rect 327 578 331 579
rect 327 573 331 574
rect 335 578 339 579
rect 335 573 339 574
rect 407 578 411 579
rect 407 573 411 574
rect 415 578 419 579
rect 415 573 419 574
rect 495 578 499 579
rect 495 573 499 574
rect 511 578 515 579
rect 511 573 515 574
rect 591 578 595 579
rect 591 573 595 574
rect 615 578 619 579
rect 615 573 619 574
rect 695 578 699 579
rect 695 573 699 574
rect 719 578 723 579
rect 719 573 723 574
rect 799 578 803 579
rect 799 573 803 574
rect 831 578 835 579
rect 831 573 835 574
rect 903 578 907 579
rect 903 573 907 574
rect 943 578 947 579
rect 943 573 947 574
rect 1007 578 1011 579
rect 1007 573 1011 574
rect 1063 578 1067 579
rect 1063 573 1067 574
rect 1103 578 1107 579
rect 1103 573 1107 574
rect 1183 578 1187 579
rect 1183 573 1187 574
rect 1207 578 1211 579
rect 1207 573 1211 574
rect 1287 578 1291 579
rect 1287 573 1291 574
rect 1327 578 1331 579
rect 1368 575 1370 598
rect 1414 594 1420 595
rect 1414 590 1415 594
rect 1419 590 1420 594
rect 1414 589 1420 590
rect 1526 594 1532 595
rect 1526 590 1527 594
rect 1531 590 1532 594
rect 1526 589 1532 590
rect 1662 594 1668 595
rect 1662 590 1663 594
rect 1667 590 1668 594
rect 1662 589 1668 590
rect 1798 594 1804 595
rect 1798 590 1799 594
rect 1803 590 1804 594
rect 1798 589 1804 590
rect 1926 594 1932 595
rect 1926 590 1927 594
rect 1931 590 1932 594
rect 1926 589 1932 590
rect 2054 594 2060 595
rect 2054 590 2055 594
rect 2059 590 2060 594
rect 2054 589 2060 590
rect 2174 594 2180 595
rect 2174 590 2175 594
rect 2179 590 2180 594
rect 2174 589 2180 590
rect 2294 594 2300 595
rect 2294 590 2295 594
rect 2299 590 2300 594
rect 2294 589 2300 590
rect 2422 594 2428 595
rect 2422 590 2423 594
rect 2427 590 2428 594
rect 2422 589 2428 590
rect 1416 575 1418 589
rect 1528 575 1530 589
rect 1664 575 1666 589
rect 1800 575 1802 589
rect 1928 575 1930 589
rect 2056 575 2058 589
rect 2176 575 2178 589
rect 2296 575 2298 589
rect 2424 575 2426 589
rect 2584 575 2586 598
rect 1327 573 1331 574
rect 1367 574 1371 575
rect 112 558 114 573
rect 200 567 202 573
rect 264 567 266 573
rect 336 567 338 573
rect 416 567 418 573
rect 512 567 514 573
rect 616 567 618 573
rect 720 567 722 573
rect 832 567 834 573
rect 944 567 946 573
rect 1064 567 1066 573
rect 1184 567 1186 573
rect 1288 567 1290 573
rect 198 566 204 567
rect 198 562 199 566
rect 203 562 204 566
rect 198 561 204 562
rect 262 566 268 567
rect 262 562 263 566
rect 267 562 268 566
rect 262 561 268 562
rect 334 566 340 567
rect 334 562 335 566
rect 339 562 340 566
rect 334 561 340 562
rect 414 566 420 567
rect 414 562 415 566
rect 419 562 420 566
rect 414 561 420 562
rect 510 566 516 567
rect 510 562 511 566
rect 515 562 516 566
rect 510 561 516 562
rect 614 566 620 567
rect 614 562 615 566
rect 619 562 620 566
rect 614 561 620 562
rect 718 566 724 567
rect 718 562 719 566
rect 723 562 724 566
rect 718 561 724 562
rect 830 566 836 567
rect 830 562 831 566
rect 835 562 836 566
rect 830 561 836 562
rect 942 566 948 567
rect 942 562 943 566
rect 947 562 948 566
rect 942 561 948 562
rect 1062 566 1068 567
rect 1062 562 1063 566
rect 1067 562 1068 566
rect 1062 561 1068 562
rect 1182 566 1188 567
rect 1182 562 1183 566
rect 1187 562 1188 566
rect 1182 561 1188 562
rect 1286 566 1292 567
rect 1286 562 1287 566
rect 1291 562 1292 566
rect 1286 561 1292 562
rect 1328 558 1330 573
rect 1367 569 1371 570
rect 1415 574 1419 575
rect 1415 569 1419 570
rect 1471 574 1475 575
rect 1471 569 1475 570
rect 1527 574 1531 575
rect 1527 569 1531 570
rect 1551 574 1555 575
rect 1551 569 1555 570
rect 1647 574 1651 575
rect 1647 569 1651 570
rect 1663 574 1667 575
rect 1663 569 1667 570
rect 1751 574 1755 575
rect 1751 569 1755 570
rect 1799 574 1803 575
rect 1799 569 1803 570
rect 1855 574 1859 575
rect 1855 569 1859 570
rect 1927 574 1931 575
rect 1927 569 1931 570
rect 1959 574 1963 575
rect 1959 569 1963 570
rect 2055 574 2059 575
rect 2055 569 2059 570
rect 2151 574 2155 575
rect 2151 569 2155 570
rect 2175 574 2179 575
rect 2175 569 2179 570
rect 2239 574 2243 575
rect 2239 569 2243 570
rect 2295 574 2299 575
rect 2295 569 2299 570
rect 2319 574 2323 575
rect 2319 569 2323 570
rect 2399 574 2403 575
rect 2399 569 2403 570
rect 2423 574 2427 575
rect 2423 569 2427 570
rect 2479 574 2483 575
rect 2479 569 2483 570
rect 2543 574 2547 575
rect 2543 569 2547 570
rect 2583 574 2587 575
rect 2583 569 2587 570
rect 110 557 116 558
rect 110 553 111 557
rect 115 553 116 557
rect 110 552 116 553
rect 1326 557 1332 558
rect 1326 553 1327 557
rect 1331 553 1332 557
rect 1368 554 1370 569
rect 1416 563 1418 569
rect 1472 563 1474 569
rect 1552 563 1554 569
rect 1648 563 1650 569
rect 1752 563 1754 569
rect 1856 563 1858 569
rect 1960 563 1962 569
rect 2056 563 2058 569
rect 2152 563 2154 569
rect 2240 563 2242 569
rect 2320 563 2322 569
rect 2400 563 2402 569
rect 2480 563 2482 569
rect 2544 563 2546 569
rect 1414 562 1420 563
rect 1414 558 1415 562
rect 1419 558 1420 562
rect 1414 557 1420 558
rect 1470 562 1476 563
rect 1470 558 1471 562
rect 1475 558 1476 562
rect 1470 557 1476 558
rect 1550 562 1556 563
rect 1550 558 1551 562
rect 1555 558 1556 562
rect 1550 557 1556 558
rect 1646 562 1652 563
rect 1646 558 1647 562
rect 1651 558 1652 562
rect 1646 557 1652 558
rect 1750 562 1756 563
rect 1750 558 1751 562
rect 1755 558 1756 562
rect 1750 557 1756 558
rect 1854 562 1860 563
rect 1854 558 1855 562
rect 1859 558 1860 562
rect 1854 557 1860 558
rect 1958 562 1964 563
rect 1958 558 1959 562
rect 1963 558 1964 562
rect 1958 557 1964 558
rect 2054 562 2060 563
rect 2054 558 2055 562
rect 2059 558 2060 562
rect 2054 557 2060 558
rect 2150 562 2156 563
rect 2150 558 2151 562
rect 2155 558 2156 562
rect 2150 557 2156 558
rect 2238 562 2244 563
rect 2238 558 2239 562
rect 2243 558 2244 562
rect 2238 557 2244 558
rect 2318 562 2324 563
rect 2318 558 2319 562
rect 2323 558 2324 562
rect 2318 557 2324 558
rect 2398 562 2404 563
rect 2398 558 2399 562
rect 2403 558 2404 562
rect 2398 557 2404 558
rect 2478 562 2484 563
rect 2478 558 2479 562
rect 2483 558 2484 562
rect 2478 557 2484 558
rect 2542 562 2548 563
rect 2542 558 2543 562
rect 2547 558 2548 562
rect 2542 557 2548 558
rect 2584 554 2586 569
rect 1326 552 1332 553
rect 1366 553 1372 554
rect 1366 549 1367 553
rect 1371 549 1372 553
rect 1366 548 1372 549
rect 2582 553 2588 554
rect 2582 549 2583 553
rect 2587 549 2588 553
rect 2582 548 2588 549
rect 110 540 116 541
rect 1326 540 1332 541
rect 110 536 111 540
rect 115 536 116 540
rect 110 535 116 536
rect 182 539 188 540
rect 182 535 183 539
rect 187 535 188 539
rect 112 515 114 535
rect 182 534 188 535
rect 246 539 252 540
rect 246 535 247 539
rect 251 535 252 539
rect 246 534 252 535
rect 318 539 324 540
rect 318 535 319 539
rect 323 535 324 539
rect 318 534 324 535
rect 398 539 404 540
rect 398 535 399 539
rect 403 535 404 539
rect 398 534 404 535
rect 494 539 500 540
rect 494 535 495 539
rect 499 535 500 539
rect 494 534 500 535
rect 598 539 604 540
rect 598 535 599 539
rect 603 535 604 539
rect 598 534 604 535
rect 702 539 708 540
rect 702 535 703 539
rect 707 535 708 539
rect 702 534 708 535
rect 814 539 820 540
rect 814 535 815 539
rect 819 535 820 539
rect 814 534 820 535
rect 926 539 932 540
rect 926 535 927 539
rect 931 535 932 539
rect 926 534 932 535
rect 1046 539 1052 540
rect 1046 535 1047 539
rect 1051 535 1052 539
rect 1046 534 1052 535
rect 1166 539 1172 540
rect 1166 535 1167 539
rect 1171 535 1172 539
rect 1166 534 1172 535
rect 1270 539 1276 540
rect 1270 535 1271 539
rect 1275 535 1276 539
rect 1326 536 1327 540
rect 1331 536 1332 540
rect 1326 535 1332 536
rect 1366 536 1372 537
rect 2582 536 2588 537
rect 1270 534 1276 535
rect 184 515 186 534
rect 248 515 250 534
rect 320 515 322 534
rect 400 515 402 534
rect 496 515 498 534
rect 600 515 602 534
rect 704 515 706 534
rect 816 515 818 534
rect 928 515 930 534
rect 1048 515 1050 534
rect 1168 515 1170 534
rect 1272 515 1274 534
rect 1328 515 1330 535
rect 1366 532 1367 536
rect 1371 532 1372 536
rect 1366 531 1372 532
rect 1398 535 1404 536
rect 1398 531 1399 535
rect 1403 531 1404 535
rect 1368 519 1370 531
rect 1398 530 1404 531
rect 1454 535 1460 536
rect 1454 531 1455 535
rect 1459 531 1460 535
rect 1454 530 1460 531
rect 1534 535 1540 536
rect 1534 531 1535 535
rect 1539 531 1540 535
rect 1534 530 1540 531
rect 1630 535 1636 536
rect 1630 531 1631 535
rect 1635 531 1636 535
rect 1630 530 1636 531
rect 1734 535 1740 536
rect 1734 531 1735 535
rect 1739 531 1740 535
rect 1734 530 1740 531
rect 1838 535 1844 536
rect 1838 531 1839 535
rect 1843 531 1844 535
rect 1838 530 1844 531
rect 1942 535 1948 536
rect 1942 531 1943 535
rect 1947 531 1948 535
rect 1942 530 1948 531
rect 2038 535 2044 536
rect 2038 531 2039 535
rect 2043 531 2044 535
rect 2038 530 2044 531
rect 2134 535 2140 536
rect 2134 531 2135 535
rect 2139 531 2140 535
rect 2134 530 2140 531
rect 2222 535 2228 536
rect 2222 531 2223 535
rect 2227 531 2228 535
rect 2222 530 2228 531
rect 2302 535 2308 536
rect 2302 531 2303 535
rect 2307 531 2308 535
rect 2302 530 2308 531
rect 2382 535 2388 536
rect 2382 531 2383 535
rect 2387 531 2388 535
rect 2382 530 2388 531
rect 2462 535 2468 536
rect 2462 531 2463 535
rect 2467 531 2468 535
rect 2462 530 2468 531
rect 2526 535 2532 536
rect 2526 531 2527 535
rect 2531 531 2532 535
rect 2582 532 2583 536
rect 2587 532 2588 536
rect 2582 531 2588 532
rect 2526 530 2532 531
rect 1400 519 1402 530
rect 1456 519 1458 530
rect 1536 519 1538 530
rect 1632 519 1634 530
rect 1736 519 1738 530
rect 1840 519 1842 530
rect 1944 519 1946 530
rect 2040 519 2042 530
rect 2136 519 2138 530
rect 2224 519 2226 530
rect 2304 519 2306 530
rect 2384 519 2386 530
rect 2464 519 2466 530
rect 2528 519 2530 530
rect 2584 519 2586 531
rect 1367 518 1371 519
rect 111 514 115 515
rect 111 509 115 510
rect 183 514 187 515
rect 183 509 187 510
rect 247 514 251 515
rect 247 509 251 510
rect 303 514 307 515
rect 303 509 307 510
rect 319 514 323 515
rect 319 509 323 510
rect 359 514 363 515
rect 359 509 363 510
rect 399 514 403 515
rect 399 509 403 510
rect 423 514 427 515
rect 423 509 427 510
rect 495 514 499 515
rect 495 509 499 510
rect 575 514 579 515
rect 575 509 579 510
rect 599 514 603 515
rect 599 509 603 510
rect 647 514 651 515
rect 647 509 651 510
rect 703 514 707 515
rect 703 509 707 510
rect 719 514 723 515
rect 719 509 723 510
rect 791 514 795 515
rect 791 509 795 510
rect 815 514 819 515
rect 815 509 819 510
rect 863 514 867 515
rect 863 509 867 510
rect 927 514 931 515
rect 927 509 931 510
rect 935 514 939 515
rect 935 509 939 510
rect 1007 514 1011 515
rect 1007 509 1011 510
rect 1047 514 1051 515
rect 1047 509 1051 510
rect 1087 514 1091 515
rect 1087 509 1091 510
rect 1167 514 1171 515
rect 1167 509 1171 510
rect 1271 514 1275 515
rect 1271 509 1275 510
rect 1327 514 1331 515
rect 1367 513 1371 514
rect 1399 518 1403 519
rect 1399 513 1403 514
rect 1455 518 1459 519
rect 1455 513 1459 514
rect 1535 518 1539 519
rect 1535 513 1539 514
rect 1599 518 1603 519
rect 1599 513 1603 514
rect 1631 518 1635 519
rect 1631 513 1635 514
rect 1671 518 1675 519
rect 1671 513 1675 514
rect 1735 518 1739 519
rect 1735 513 1739 514
rect 1751 518 1755 519
rect 1751 513 1755 514
rect 1839 518 1843 519
rect 1839 513 1843 514
rect 1927 518 1931 519
rect 1927 513 1931 514
rect 1943 518 1947 519
rect 1943 513 1947 514
rect 2015 518 2019 519
rect 2015 513 2019 514
rect 2039 518 2043 519
rect 2039 513 2043 514
rect 2095 518 2099 519
rect 2095 513 2099 514
rect 2135 518 2139 519
rect 2135 513 2139 514
rect 2175 518 2179 519
rect 2175 513 2179 514
rect 2223 518 2227 519
rect 2223 513 2227 514
rect 2255 518 2259 519
rect 2255 513 2259 514
rect 2303 518 2307 519
rect 2303 513 2307 514
rect 2327 518 2331 519
rect 2327 513 2331 514
rect 2383 518 2387 519
rect 2383 513 2387 514
rect 2399 518 2403 519
rect 2399 513 2403 514
rect 2463 518 2467 519
rect 2463 513 2467 514
rect 2471 518 2475 519
rect 2471 513 2475 514
rect 2527 518 2531 519
rect 2527 513 2531 514
rect 2583 518 2587 519
rect 2583 513 2587 514
rect 1327 509 1331 510
rect 112 497 114 509
rect 304 498 306 509
rect 360 498 362 509
rect 424 498 426 509
rect 496 498 498 509
rect 576 498 578 509
rect 648 498 650 509
rect 720 498 722 509
rect 792 498 794 509
rect 864 498 866 509
rect 936 498 938 509
rect 1008 498 1010 509
rect 1088 498 1090 509
rect 302 497 308 498
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 302 493 303 497
rect 307 493 308 497
rect 302 492 308 493
rect 358 497 364 498
rect 358 493 359 497
rect 363 493 364 497
rect 358 492 364 493
rect 422 497 428 498
rect 422 493 423 497
rect 427 493 428 497
rect 422 492 428 493
rect 494 497 500 498
rect 494 493 495 497
rect 499 493 500 497
rect 494 492 500 493
rect 574 497 580 498
rect 574 493 575 497
rect 579 493 580 497
rect 574 492 580 493
rect 646 497 652 498
rect 646 493 647 497
rect 651 493 652 497
rect 646 492 652 493
rect 718 497 724 498
rect 718 493 719 497
rect 723 493 724 497
rect 718 492 724 493
rect 790 497 796 498
rect 790 493 791 497
rect 795 493 796 497
rect 790 492 796 493
rect 862 497 868 498
rect 862 493 863 497
rect 867 493 868 497
rect 862 492 868 493
rect 934 497 940 498
rect 934 493 935 497
rect 939 493 940 497
rect 934 492 940 493
rect 1006 497 1012 498
rect 1006 493 1007 497
rect 1011 493 1012 497
rect 1006 492 1012 493
rect 1086 497 1092 498
rect 1328 497 1330 509
rect 1368 501 1370 513
rect 1536 502 1538 513
rect 1600 502 1602 513
rect 1672 502 1674 513
rect 1752 502 1754 513
rect 1840 502 1842 513
rect 1928 502 1930 513
rect 2016 502 2018 513
rect 2096 502 2098 513
rect 2176 502 2178 513
rect 2256 502 2258 513
rect 2328 502 2330 513
rect 2400 502 2402 513
rect 2472 502 2474 513
rect 2528 502 2530 513
rect 1534 501 1540 502
rect 1366 500 1372 501
rect 1086 493 1087 497
rect 1091 493 1092 497
rect 1086 492 1092 493
rect 1326 496 1332 497
rect 1326 492 1327 496
rect 1331 492 1332 496
rect 1366 496 1367 500
rect 1371 496 1372 500
rect 1534 497 1535 501
rect 1539 497 1540 501
rect 1534 496 1540 497
rect 1598 501 1604 502
rect 1598 497 1599 501
rect 1603 497 1604 501
rect 1598 496 1604 497
rect 1670 501 1676 502
rect 1670 497 1671 501
rect 1675 497 1676 501
rect 1670 496 1676 497
rect 1750 501 1756 502
rect 1750 497 1751 501
rect 1755 497 1756 501
rect 1750 496 1756 497
rect 1838 501 1844 502
rect 1838 497 1839 501
rect 1843 497 1844 501
rect 1838 496 1844 497
rect 1926 501 1932 502
rect 1926 497 1927 501
rect 1931 497 1932 501
rect 1926 496 1932 497
rect 2014 501 2020 502
rect 2014 497 2015 501
rect 2019 497 2020 501
rect 2014 496 2020 497
rect 2094 501 2100 502
rect 2094 497 2095 501
rect 2099 497 2100 501
rect 2094 496 2100 497
rect 2174 501 2180 502
rect 2174 497 2175 501
rect 2179 497 2180 501
rect 2174 496 2180 497
rect 2254 501 2260 502
rect 2254 497 2255 501
rect 2259 497 2260 501
rect 2254 496 2260 497
rect 2326 501 2332 502
rect 2326 497 2327 501
rect 2331 497 2332 501
rect 2326 496 2332 497
rect 2398 501 2404 502
rect 2398 497 2399 501
rect 2403 497 2404 501
rect 2398 496 2404 497
rect 2470 501 2476 502
rect 2470 497 2471 501
rect 2475 497 2476 501
rect 2470 496 2476 497
rect 2526 501 2532 502
rect 2584 501 2586 513
rect 2526 497 2527 501
rect 2531 497 2532 501
rect 2526 496 2532 497
rect 2582 500 2588 501
rect 2582 496 2583 500
rect 2587 496 2588 500
rect 1366 495 1372 496
rect 2582 495 2588 496
rect 110 491 116 492
rect 1326 491 1332 492
rect 1366 483 1372 484
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 110 474 116 475
rect 1326 479 1332 480
rect 1326 475 1327 479
rect 1331 475 1332 479
rect 1366 479 1367 483
rect 1371 479 1372 483
rect 1366 478 1372 479
rect 2582 483 2588 484
rect 2582 479 2583 483
rect 2587 479 2588 483
rect 2582 478 2588 479
rect 1326 474 1332 475
rect 112 455 114 474
rect 318 470 324 471
rect 318 466 319 470
rect 323 466 324 470
rect 318 465 324 466
rect 374 470 380 471
rect 374 466 375 470
rect 379 466 380 470
rect 374 465 380 466
rect 438 470 444 471
rect 438 466 439 470
rect 443 466 444 470
rect 438 465 444 466
rect 510 470 516 471
rect 510 466 511 470
rect 515 466 516 470
rect 510 465 516 466
rect 590 470 596 471
rect 590 466 591 470
rect 595 466 596 470
rect 590 465 596 466
rect 662 470 668 471
rect 662 466 663 470
rect 667 466 668 470
rect 662 465 668 466
rect 734 470 740 471
rect 734 466 735 470
rect 739 466 740 470
rect 734 465 740 466
rect 806 470 812 471
rect 806 466 807 470
rect 811 466 812 470
rect 806 465 812 466
rect 878 470 884 471
rect 878 466 879 470
rect 883 466 884 470
rect 878 465 884 466
rect 950 470 956 471
rect 950 466 951 470
rect 955 466 956 470
rect 950 465 956 466
rect 1022 470 1028 471
rect 1022 466 1023 470
rect 1027 466 1028 470
rect 1022 465 1028 466
rect 1102 470 1108 471
rect 1102 466 1103 470
rect 1107 466 1108 470
rect 1102 465 1108 466
rect 320 455 322 465
rect 376 455 378 465
rect 440 455 442 465
rect 512 455 514 465
rect 592 455 594 465
rect 664 455 666 465
rect 736 455 738 465
rect 808 455 810 465
rect 880 455 882 465
rect 952 455 954 465
rect 1024 455 1026 465
rect 1104 455 1106 465
rect 1328 455 1330 474
rect 1368 455 1370 478
rect 1550 474 1556 475
rect 1550 470 1551 474
rect 1555 470 1556 474
rect 1550 469 1556 470
rect 1614 474 1620 475
rect 1614 470 1615 474
rect 1619 470 1620 474
rect 1614 469 1620 470
rect 1686 474 1692 475
rect 1686 470 1687 474
rect 1691 470 1692 474
rect 1686 469 1692 470
rect 1766 474 1772 475
rect 1766 470 1767 474
rect 1771 470 1772 474
rect 1766 469 1772 470
rect 1854 474 1860 475
rect 1854 470 1855 474
rect 1859 470 1860 474
rect 1854 469 1860 470
rect 1942 474 1948 475
rect 1942 470 1943 474
rect 1947 470 1948 474
rect 1942 469 1948 470
rect 2030 474 2036 475
rect 2030 470 2031 474
rect 2035 470 2036 474
rect 2030 469 2036 470
rect 2110 474 2116 475
rect 2110 470 2111 474
rect 2115 470 2116 474
rect 2110 469 2116 470
rect 2190 474 2196 475
rect 2190 470 2191 474
rect 2195 470 2196 474
rect 2190 469 2196 470
rect 2270 474 2276 475
rect 2270 470 2271 474
rect 2275 470 2276 474
rect 2270 469 2276 470
rect 2342 474 2348 475
rect 2342 470 2343 474
rect 2347 470 2348 474
rect 2342 469 2348 470
rect 2414 474 2420 475
rect 2414 470 2415 474
rect 2419 470 2420 474
rect 2414 469 2420 470
rect 2486 474 2492 475
rect 2486 470 2487 474
rect 2491 470 2492 474
rect 2486 469 2492 470
rect 2542 474 2548 475
rect 2542 470 2543 474
rect 2547 470 2548 474
rect 2542 469 2548 470
rect 1552 455 1554 469
rect 1616 455 1618 469
rect 1688 455 1690 469
rect 1768 455 1770 469
rect 1856 455 1858 469
rect 1944 455 1946 469
rect 2032 455 2034 469
rect 2112 455 2114 469
rect 2192 455 2194 469
rect 2272 455 2274 469
rect 2344 455 2346 469
rect 2416 455 2418 469
rect 2488 455 2490 469
rect 2544 455 2546 469
rect 2584 455 2586 478
rect 111 454 115 455
rect 111 449 115 450
rect 319 454 323 455
rect 319 449 323 450
rect 375 454 379 455
rect 375 449 379 450
rect 439 454 443 455
rect 439 449 443 450
rect 455 454 459 455
rect 455 449 459 450
rect 511 454 515 455
rect 511 449 515 450
rect 575 454 579 455
rect 575 449 579 450
rect 591 454 595 455
rect 591 449 595 450
rect 647 454 651 455
rect 647 449 651 450
rect 663 454 667 455
rect 663 449 667 450
rect 727 454 731 455
rect 727 449 731 450
rect 735 454 739 455
rect 735 449 739 450
rect 799 454 803 455
rect 799 449 803 450
rect 807 454 811 455
rect 807 449 811 450
rect 871 454 875 455
rect 871 449 875 450
rect 879 454 883 455
rect 879 449 883 450
rect 943 454 947 455
rect 943 449 947 450
rect 951 454 955 455
rect 951 449 955 450
rect 1015 454 1019 455
rect 1015 449 1019 450
rect 1023 454 1027 455
rect 1023 449 1027 450
rect 1087 454 1091 455
rect 1087 449 1091 450
rect 1103 454 1107 455
rect 1103 449 1107 450
rect 1159 454 1163 455
rect 1159 449 1163 450
rect 1239 454 1243 455
rect 1239 449 1243 450
rect 1327 454 1331 455
rect 1327 449 1331 450
rect 1367 454 1371 455
rect 1367 449 1371 450
rect 1551 454 1555 455
rect 1551 449 1555 450
rect 1615 454 1619 455
rect 1615 449 1619 450
rect 1647 454 1651 455
rect 1647 449 1651 450
rect 1687 454 1691 455
rect 1687 449 1691 450
rect 1703 454 1707 455
rect 1703 449 1707 450
rect 1759 454 1763 455
rect 1759 449 1763 450
rect 1767 454 1771 455
rect 1767 449 1771 450
rect 1815 454 1819 455
rect 1815 449 1819 450
rect 1855 454 1859 455
rect 1855 449 1859 450
rect 1871 454 1875 455
rect 1871 449 1875 450
rect 1927 454 1931 455
rect 1927 449 1931 450
rect 1943 454 1947 455
rect 1943 449 1947 450
rect 1999 454 2003 455
rect 1999 449 2003 450
rect 2031 454 2035 455
rect 2031 449 2035 450
rect 2087 454 2091 455
rect 2087 449 2091 450
rect 2111 454 2115 455
rect 2111 449 2115 450
rect 2191 454 2195 455
rect 2191 449 2195 450
rect 2271 454 2275 455
rect 2271 449 2275 450
rect 2311 454 2315 455
rect 2311 449 2315 450
rect 2343 454 2347 455
rect 2343 449 2347 450
rect 2415 454 2419 455
rect 2415 449 2419 450
rect 2439 454 2443 455
rect 2439 449 2443 450
rect 2487 454 2491 455
rect 2487 449 2491 450
rect 2543 454 2547 455
rect 2543 449 2547 450
rect 2583 454 2587 455
rect 2583 449 2587 450
rect 112 434 114 449
rect 456 443 458 449
rect 512 443 514 449
rect 576 443 578 449
rect 648 443 650 449
rect 728 443 730 449
rect 800 443 802 449
rect 872 443 874 449
rect 944 443 946 449
rect 1016 443 1018 449
rect 1088 443 1090 449
rect 1160 443 1162 449
rect 1240 443 1242 449
rect 454 442 460 443
rect 454 438 455 442
rect 459 438 460 442
rect 454 437 460 438
rect 510 442 516 443
rect 510 438 511 442
rect 515 438 516 442
rect 510 437 516 438
rect 574 442 580 443
rect 574 438 575 442
rect 579 438 580 442
rect 574 437 580 438
rect 646 442 652 443
rect 646 438 647 442
rect 651 438 652 442
rect 646 437 652 438
rect 726 442 732 443
rect 726 438 727 442
rect 731 438 732 442
rect 726 437 732 438
rect 798 442 804 443
rect 798 438 799 442
rect 803 438 804 442
rect 798 437 804 438
rect 870 442 876 443
rect 870 438 871 442
rect 875 438 876 442
rect 870 437 876 438
rect 942 442 948 443
rect 942 438 943 442
rect 947 438 948 442
rect 942 437 948 438
rect 1014 442 1020 443
rect 1014 438 1015 442
rect 1019 438 1020 442
rect 1014 437 1020 438
rect 1086 442 1092 443
rect 1086 438 1087 442
rect 1091 438 1092 442
rect 1086 437 1092 438
rect 1158 442 1164 443
rect 1158 438 1159 442
rect 1163 438 1164 442
rect 1158 437 1164 438
rect 1238 442 1244 443
rect 1238 438 1239 442
rect 1243 438 1244 442
rect 1238 437 1244 438
rect 1328 434 1330 449
rect 1368 434 1370 449
rect 1648 443 1650 449
rect 1704 443 1706 449
rect 1760 443 1762 449
rect 1816 443 1818 449
rect 1872 443 1874 449
rect 1928 443 1930 449
rect 2000 443 2002 449
rect 2088 443 2090 449
rect 2192 443 2194 449
rect 2312 443 2314 449
rect 2440 443 2442 449
rect 2544 443 2546 449
rect 1646 442 1652 443
rect 1646 438 1647 442
rect 1651 438 1652 442
rect 1646 437 1652 438
rect 1702 442 1708 443
rect 1702 438 1703 442
rect 1707 438 1708 442
rect 1702 437 1708 438
rect 1758 442 1764 443
rect 1758 438 1759 442
rect 1763 438 1764 442
rect 1758 437 1764 438
rect 1814 442 1820 443
rect 1814 438 1815 442
rect 1819 438 1820 442
rect 1814 437 1820 438
rect 1870 442 1876 443
rect 1870 438 1871 442
rect 1875 438 1876 442
rect 1870 437 1876 438
rect 1926 442 1932 443
rect 1926 438 1927 442
rect 1931 438 1932 442
rect 1926 437 1932 438
rect 1998 442 2004 443
rect 1998 438 1999 442
rect 2003 438 2004 442
rect 1998 437 2004 438
rect 2086 442 2092 443
rect 2086 438 2087 442
rect 2091 438 2092 442
rect 2086 437 2092 438
rect 2190 442 2196 443
rect 2190 438 2191 442
rect 2195 438 2196 442
rect 2190 437 2196 438
rect 2310 442 2316 443
rect 2310 438 2311 442
rect 2315 438 2316 442
rect 2310 437 2316 438
rect 2438 442 2444 443
rect 2438 438 2439 442
rect 2443 438 2444 442
rect 2438 437 2444 438
rect 2542 442 2548 443
rect 2542 438 2543 442
rect 2547 438 2548 442
rect 2542 437 2548 438
rect 2584 434 2586 449
rect 110 433 116 434
rect 110 429 111 433
rect 115 429 116 433
rect 110 428 116 429
rect 1326 433 1332 434
rect 1326 429 1327 433
rect 1331 429 1332 433
rect 1326 428 1332 429
rect 1366 433 1372 434
rect 1366 429 1367 433
rect 1371 429 1372 433
rect 1366 428 1372 429
rect 2582 433 2588 434
rect 2582 429 2583 433
rect 2587 429 2588 433
rect 2582 428 2588 429
rect 110 416 116 417
rect 1326 416 1332 417
rect 110 412 111 416
rect 115 412 116 416
rect 110 411 116 412
rect 438 415 444 416
rect 438 411 439 415
rect 443 411 444 415
rect 112 395 114 411
rect 438 410 444 411
rect 494 415 500 416
rect 494 411 495 415
rect 499 411 500 415
rect 494 410 500 411
rect 558 415 564 416
rect 558 411 559 415
rect 563 411 564 415
rect 558 410 564 411
rect 630 415 636 416
rect 630 411 631 415
rect 635 411 636 415
rect 630 410 636 411
rect 710 415 716 416
rect 710 411 711 415
rect 715 411 716 415
rect 710 410 716 411
rect 782 415 788 416
rect 782 411 783 415
rect 787 411 788 415
rect 782 410 788 411
rect 854 415 860 416
rect 854 411 855 415
rect 859 411 860 415
rect 854 410 860 411
rect 926 415 932 416
rect 926 411 927 415
rect 931 411 932 415
rect 926 410 932 411
rect 998 415 1004 416
rect 998 411 999 415
rect 1003 411 1004 415
rect 998 410 1004 411
rect 1070 415 1076 416
rect 1070 411 1071 415
rect 1075 411 1076 415
rect 1070 410 1076 411
rect 1142 415 1148 416
rect 1142 411 1143 415
rect 1147 411 1148 415
rect 1142 410 1148 411
rect 1222 415 1228 416
rect 1222 411 1223 415
rect 1227 411 1228 415
rect 1326 412 1327 416
rect 1331 412 1332 416
rect 1326 411 1332 412
rect 1366 416 1372 417
rect 2582 416 2588 417
rect 1366 412 1367 416
rect 1371 412 1372 416
rect 1366 411 1372 412
rect 1630 415 1636 416
rect 1630 411 1631 415
rect 1635 411 1636 415
rect 1222 410 1228 411
rect 440 395 442 410
rect 496 395 498 410
rect 560 395 562 410
rect 632 395 634 410
rect 712 395 714 410
rect 784 395 786 410
rect 856 395 858 410
rect 928 395 930 410
rect 1000 395 1002 410
rect 1072 395 1074 410
rect 1144 395 1146 410
rect 1224 395 1226 410
rect 1328 395 1330 411
rect 1368 399 1370 411
rect 1630 410 1636 411
rect 1686 415 1692 416
rect 1686 411 1687 415
rect 1691 411 1692 415
rect 1686 410 1692 411
rect 1742 415 1748 416
rect 1742 411 1743 415
rect 1747 411 1748 415
rect 1742 410 1748 411
rect 1798 415 1804 416
rect 1798 411 1799 415
rect 1803 411 1804 415
rect 1798 410 1804 411
rect 1854 415 1860 416
rect 1854 411 1855 415
rect 1859 411 1860 415
rect 1854 410 1860 411
rect 1910 415 1916 416
rect 1910 411 1911 415
rect 1915 411 1916 415
rect 1910 410 1916 411
rect 1982 415 1988 416
rect 1982 411 1983 415
rect 1987 411 1988 415
rect 1982 410 1988 411
rect 2070 415 2076 416
rect 2070 411 2071 415
rect 2075 411 2076 415
rect 2070 410 2076 411
rect 2174 415 2180 416
rect 2174 411 2175 415
rect 2179 411 2180 415
rect 2174 410 2180 411
rect 2294 415 2300 416
rect 2294 411 2295 415
rect 2299 411 2300 415
rect 2294 410 2300 411
rect 2422 415 2428 416
rect 2422 411 2423 415
rect 2427 411 2428 415
rect 2422 410 2428 411
rect 2526 415 2532 416
rect 2526 411 2527 415
rect 2531 411 2532 415
rect 2582 412 2583 416
rect 2587 412 2588 416
rect 2582 411 2588 412
rect 2526 410 2532 411
rect 1632 399 1634 410
rect 1688 399 1690 410
rect 1744 399 1746 410
rect 1800 399 1802 410
rect 1856 399 1858 410
rect 1912 399 1914 410
rect 1984 399 1986 410
rect 2072 399 2074 410
rect 2176 399 2178 410
rect 2296 399 2298 410
rect 2424 399 2426 410
rect 2528 399 2530 410
rect 2584 399 2586 411
rect 1367 398 1371 399
rect 111 394 115 395
rect 111 389 115 390
rect 415 394 419 395
rect 415 389 419 390
rect 439 394 443 395
rect 439 389 443 390
rect 471 394 475 395
rect 471 389 475 390
rect 495 394 499 395
rect 495 389 499 390
rect 535 394 539 395
rect 535 389 539 390
rect 559 394 563 395
rect 559 389 563 390
rect 607 394 611 395
rect 607 389 611 390
rect 631 394 635 395
rect 631 389 635 390
rect 687 394 691 395
rect 687 389 691 390
rect 711 394 715 395
rect 711 389 715 390
rect 767 394 771 395
rect 767 389 771 390
rect 783 394 787 395
rect 783 389 787 390
rect 847 394 851 395
rect 847 389 851 390
rect 855 394 859 395
rect 855 389 859 390
rect 927 394 931 395
rect 927 389 931 390
rect 999 394 1003 395
rect 999 389 1003 390
rect 1007 394 1011 395
rect 1007 389 1011 390
rect 1071 394 1075 395
rect 1071 389 1075 390
rect 1087 394 1091 395
rect 1087 389 1091 390
rect 1143 394 1147 395
rect 1143 389 1147 390
rect 1175 394 1179 395
rect 1175 389 1179 390
rect 1223 394 1227 395
rect 1223 389 1227 390
rect 1263 394 1267 395
rect 1263 389 1267 390
rect 1327 394 1331 395
rect 1367 393 1371 394
rect 1631 398 1635 399
rect 1631 393 1635 394
rect 1655 398 1659 399
rect 1655 393 1659 394
rect 1687 398 1691 399
rect 1687 393 1691 394
rect 1711 398 1715 399
rect 1711 393 1715 394
rect 1743 398 1747 399
rect 1743 393 1747 394
rect 1767 398 1771 399
rect 1767 393 1771 394
rect 1799 398 1803 399
rect 1799 393 1803 394
rect 1823 398 1827 399
rect 1823 393 1827 394
rect 1855 398 1859 399
rect 1855 393 1859 394
rect 1879 398 1883 399
rect 1879 393 1883 394
rect 1911 398 1915 399
rect 1911 393 1915 394
rect 1951 398 1955 399
rect 1951 393 1955 394
rect 1983 398 1987 399
rect 1983 393 1987 394
rect 2039 398 2043 399
rect 2039 393 2043 394
rect 2071 398 2075 399
rect 2071 393 2075 394
rect 2151 398 2155 399
rect 2151 393 2155 394
rect 2175 398 2179 399
rect 2175 393 2179 394
rect 2279 398 2283 399
rect 2279 393 2283 394
rect 2295 398 2299 399
rect 2295 393 2299 394
rect 2415 398 2419 399
rect 2415 393 2419 394
rect 2423 398 2427 399
rect 2423 393 2427 394
rect 2527 398 2531 399
rect 2527 393 2531 394
rect 2583 398 2587 399
rect 2583 393 2587 394
rect 1327 389 1331 390
rect 112 377 114 389
rect 416 378 418 389
rect 472 378 474 389
rect 536 378 538 389
rect 608 378 610 389
rect 688 378 690 389
rect 768 378 770 389
rect 848 378 850 389
rect 928 378 930 389
rect 1008 378 1010 389
rect 1088 378 1090 389
rect 1176 378 1178 389
rect 1264 378 1266 389
rect 414 377 420 378
rect 110 376 116 377
rect 110 372 111 376
rect 115 372 116 376
rect 414 373 415 377
rect 419 373 420 377
rect 414 372 420 373
rect 470 377 476 378
rect 470 373 471 377
rect 475 373 476 377
rect 470 372 476 373
rect 534 377 540 378
rect 534 373 535 377
rect 539 373 540 377
rect 534 372 540 373
rect 606 377 612 378
rect 606 373 607 377
rect 611 373 612 377
rect 606 372 612 373
rect 686 377 692 378
rect 686 373 687 377
rect 691 373 692 377
rect 686 372 692 373
rect 766 377 772 378
rect 766 373 767 377
rect 771 373 772 377
rect 766 372 772 373
rect 846 377 852 378
rect 846 373 847 377
rect 851 373 852 377
rect 846 372 852 373
rect 926 377 932 378
rect 926 373 927 377
rect 931 373 932 377
rect 926 372 932 373
rect 1006 377 1012 378
rect 1006 373 1007 377
rect 1011 373 1012 377
rect 1006 372 1012 373
rect 1086 377 1092 378
rect 1086 373 1087 377
rect 1091 373 1092 377
rect 1086 372 1092 373
rect 1174 377 1180 378
rect 1174 373 1175 377
rect 1179 373 1180 377
rect 1174 372 1180 373
rect 1262 377 1268 378
rect 1328 377 1330 389
rect 1368 381 1370 393
rect 1656 382 1658 393
rect 1712 382 1714 393
rect 1768 382 1770 393
rect 1824 382 1826 393
rect 1880 382 1882 393
rect 1952 382 1954 393
rect 2040 382 2042 393
rect 2152 382 2154 393
rect 2280 382 2282 393
rect 2416 382 2418 393
rect 2528 382 2530 393
rect 1654 381 1660 382
rect 1366 380 1372 381
rect 1262 373 1263 377
rect 1267 373 1268 377
rect 1262 372 1268 373
rect 1326 376 1332 377
rect 1326 372 1327 376
rect 1331 372 1332 376
rect 1366 376 1367 380
rect 1371 376 1372 380
rect 1654 377 1655 381
rect 1659 377 1660 381
rect 1654 376 1660 377
rect 1710 381 1716 382
rect 1710 377 1711 381
rect 1715 377 1716 381
rect 1710 376 1716 377
rect 1766 381 1772 382
rect 1766 377 1767 381
rect 1771 377 1772 381
rect 1766 376 1772 377
rect 1822 381 1828 382
rect 1822 377 1823 381
rect 1827 377 1828 381
rect 1822 376 1828 377
rect 1878 381 1884 382
rect 1878 377 1879 381
rect 1883 377 1884 381
rect 1878 376 1884 377
rect 1950 381 1956 382
rect 1950 377 1951 381
rect 1955 377 1956 381
rect 1950 376 1956 377
rect 2038 381 2044 382
rect 2038 377 2039 381
rect 2043 377 2044 381
rect 2038 376 2044 377
rect 2150 381 2156 382
rect 2150 377 2151 381
rect 2155 377 2156 381
rect 2150 376 2156 377
rect 2278 381 2284 382
rect 2278 377 2279 381
rect 2283 377 2284 381
rect 2278 376 2284 377
rect 2414 381 2420 382
rect 2414 377 2415 381
rect 2419 377 2420 381
rect 2414 376 2420 377
rect 2526 381 2532 382
rect 2584 381 2586 393
rect 2526 377 2527 381
rect 2531 377 2532 381
rect 2526 376 2532 377
rect 2582 380 2588 381
rect 2582 376 2583 380
rect 2587 376 2588 380
rect 1366 375 1372 376
rect 2582 375 2588 376
rect 110 371 116 372
rect 1326 371 1332 372
rect 1366 363 1372 364
rect 110 359 116 360
rect 110 355 111 359
rect 115 355 116 359
rect 110 354 116 355
rect 1326 359 1332 360
rect 1326 355 1327 359
rect 1331 355 1332 359
rect 1366 359 1367 363
rect 1371 359 1372 363
rect 1366 358 1372 359
rect 2582 363 2588 364
rect 2582 359 2583 363
rect 2587 359 2588 363
rect 2582 358 2588 359
rect 1326 354 1332 355
rect 112 335 114 354
rect 430 350 436 351
rect 430 346 431 350
rect 435 346 436 350
rect 430 345 436 346
rect 486 350 492 351
rect 486 346 487 350
rect 491 346 492 350
rect 486 345 492 346
rect 550 350 556 351
rect 550 346 551 350
rect 555 346 556 350
rect 550 345 556 346
rect 622 350 628 351
rect 622 346 623 350
rect 627 346 628 350
rect 622 345 628 346
rect 702 350 708 351
rect 702 346 703 350
rect 707 346 708 350
rect 702 345 708 346
rect 782 350 788 351
rect 782 346 783 350
rect 787 346 788 350
rect 782 345 788 346
rect 862 350 868 351
rect 862 346 863 350
rect 867 346 868 350
rect 862 345 868 346
rect 942 350 948 351
rect 942 346 943 350
rect 947 346 948 350
rect 942 345 948 346
rect 1022 350 1028 351
rect 1022 346 1023 350
rect 1027 346 1028 350
rect 1022 345 1028 346
rect 1102 350 1108 351
rect 1102 346 1103 350
rect 1107 346 1108 350
rect 1102 345 1108 346
rect 1190 350 1196 351
rect 1190 346 1191 350
rect 1195 346 1196 350
rect 1190 345 1196 346
rect 1278 350 1284 351
rect 1278 346 1279 350
rect 1283 346 1284 350
rect 1278 345 1284 346
rect 432 335 434 345
rect 488 335 490 345
rect 552 335 554 345
rect 624 335 626 345
rect 704 335 706 345
rect 784 335 786 345
rect 864 335 866 345
rect 944 335 946 345
rect 1024 335 1026 345
rect 1104 335 1106 345
rect 1192 335 1194 345
rect 1280 335 1282 345
rect 1328 335 1330 354
rect 1368 335 1370 358
rect 1670 354 1676 355
rect 1670 350 1671 354
rect 1675 350 1676 354
rect 1670 349 1676 350
rect 1726 354 1732 355
rect 1726 350 1727 354
rect 1731 350 1732 354
rect 1726 349 1732 350
rect 1782 354 1788 355
rect 1782 350 1783 354
rect 1787 350 1788 354
rect 1782 349 1788 350
rect 1838 354 1844 355
rect 1838 350 1839 354
rect 1843 350 1844 354
rect 1838 349 1844 350
rect 1894 354 1900 355
rect 1894 350 1895 354
rect 1899 350 1900 354
rect 1894 349 1900 350
rect 1966 354 1972 355
rect 1966 350 1967 354
rect 1971 350 1972 354
rect 1966 349 1972 350
rect 2054 354 2060 355
rect 2054 350 2055 354
rect 2059 350 2060 354
rect 2054 349 2060 350
rect 2166 354 2172 355
rect 2166 350 2167 354
rect 2171 350 2172 354
rect 2166 349 2172 350
rect 2294 354 2300 355
rect 2294 350 2295 354
rect 2299 350 2300 354
rect 2294 349 2300 350
rect 2430 354 2436 355
rect 2430 350 2431 354
rect 2435 350 2436 354
rect 2430 349 2436 350
rect 2542 354 2548 355
rect 2542 350 2543 354
rect 2547 350 2548 354
rect 2542 349 2548 350
rect 1672 335 1674 349
rect 1728 335 1730 349
rect 1784 335 1786 349
rect 1840 335 1842 349
rect 1896 335 1898 349
rect 1968 335 1970 349
rect 2056 335 2058 349
rect 2168 335 2170 349
rect 2296 335 2298 349
rect 2432 335 2434 349
rect 2544 335 2546 349
rect 2584 335 2586 358
rect 111 334 115 335
rect 111 329 115 330
rect 431 334 435 335
rect 431 329 435 330
rect 463 334 467 335
rect 463 329 467 330
rect 487 334 491 335
rect 487 329 491 330
rect 519 334 523 335
rect 519 329 523 330
rect 551 334 555 335
rect 551 329 555 330
rect 575 334 579 335
rect 575 329 579 330
rect 623 334 627 335
rect 623 329 627 330
rect 631 334 635 335
rect 631 329 635 330
rect 695 334 699 335
rect 695 329 699 330
rect 703 334 707 335
rect 703 329 707 330
rect 767 334 771 335
rect 767 329 771 330
rect 783 334 787 335
rect 783 329 787 330
rect 847 334 851 335
rect 847 329 851 330
rect 863 334 867 335
rect 863 329 867 330
rect 927 334 931 335
rect 927 329 931 330
rect 943 334 947 335
rect 943 329 947 330
rect 1015 334 1019 335
rect 1015 329 1019 330
rect 1023 334 1027 335
rect 1023 329 1027 330
rect 1103 334 1107 335
rect 1103 329 1107 330
rect 1111 334 1115 335
rect 1111 329 1115 330
rect 1191 334 1195 335
rect 1191 329 1195 330
rect 1215 334 1219 335
rect 1215 329 1219 330
rect 1279 334 1283 335
rect 1279 329 1283 330
rect 1327 334 1331 335
rect 1327 329 1331 330
rect 1367 334 1371 335
rect 1367 329 1371 330
rect 1631 334 1635 335
rect 1631 329 1635 330
rect 1671 334 1675 335
rect 1671 329 1675 330
rect 1687 334 1691 335
rect 1687 329 1691 330
rect 1727 334 1731 335
rect 1727 329 1731 330
rect 1743 334 1747 335
rect 1743 329 1747 330
rect 1783 334 1787 335
rect 1783 329 1787 330
rect 1807 334 1811 335
rect 1807 329 1811 330
rect 1839 334 1843 335
rect 1839 329 1843 330
rect 1887 334 1891 335
rect 1887 329 1891 330
rect 1895 334 1899 335
rect 1895 329 1899 330
rect 1967 334 1971 335
rect 1967 329 1971 330
rect 2055 334 2059 335
rect 2055 329 2059 330
rect 2143 334 2147 335
rect 2143 329 2147 330
rect 2167 334 2171 335
rect 2167 329 2171 330
rect 2231 334 2235 335
rect 2231 329 2235 330
rect 2295 334 2299 335
rect 2295 329 2299 330
rect 2311 334 2315 335
rect 2311 329 2315 330
rect 2391 334 2395 335
rect 2391 329 2395 330
rect 2431 334 2435 335
rect 2431 329 2435 330
rect 2479 334 2483 335
rect 2479 329 2483 330
rect 2543 334 2547 335
rect 2543 329 2547 330
rect 2583 334 2587 335
rect 2583 329 2587 330
rect 112 314 114 329
rect 464 323 466 329
rect 520 323 522 329
rect 576 323 578 329
rect 632 323 634 329
rect 696 323 698 329
rect 768 323 770 329
rect 848 323 850 329
rect 928 323 930 329
rect 1016 323 1018 329
rect 1112 323 1114 329
rect 1216 323 1218 329
rect 462 322 468 323
rect 462 318 463 322
rect 467 318 468 322
rect 462 317 468 318
rect 518 322 524 323
rect 518 318 519 322
rect 523 318 524 322
rect 518 317 524 318
rect 574 322 580 323
rect 574 318 575 322
rect 579 318 580 322
rect 574 317 580 318
rect 630 322 636 323
rect 630 318 631 322
rect 635 318 636 322
rect 630 317 636 318
rect 694 322 700 323
rect 694 318 695 322
rect 699 318 700 322
rect 694 317 700 318
rect 766 322 772 323
rect 766 318 767 322
rect 771 318 772 322
rect 766 317 772 318
rect 846 322 852 323
rect 846 318 847 322
rect 851 318 852 322
rect 846 317 852 318
rect 926 322 932 323
rect 926 318 927 322
rect 931 318 932 322
rect 926 317 932 318
rect 1014 322 1020 323
rect 1014 318 1015 322
rect 1019 318 1020 322
rect 1014 317 1020 318
rect 1110 322 1116 323
rect 1110 318 1111 322
rect 1115 318 1116 322
rect 1110 317 1116 318
rect 1214 322 1220 323
rect 1214 318 1215 322
rect 1219 318 1220 322
rect 1214 317 1220 318
rect 1328 314 1330 329
rect 1368 314 1370 329
rect 1632 323 1634 329
rect 1688 323 1690 329
rect 1744 323 1746 329
rect 1808 323 1810 329
rect 1888 323 1890 329
rect 1968 323 1970 329
rect 2056 323 2058 329
rect 2144 323 2146 329
rect 2232 323 2234 329
rect 2312 323 2314 329
rect 2392 323 2394 329
rect 2480 323 2482 329
rect 2544 323 2546 329
rect 1630 322 1636 323
rect 1630 318 1631 322
rect 1635 318 1636 322
rect 1630 317 1636 318
rect 1686 322 1692 323
rect 1686 318 1687 322
rect 1691 318 1692 322
rect 1686 317 1692 318
rect 1742 322 1748 323
rect 1742 318 1743 322
rect 1747 318 1748 322
rect 1742 317 1748 318
rect 1806 322 1812 323
rect 1806 318 1807 322
rect 1811 318 1812 322
rect 1806 317 1812 318
rect 1886 322 1892 323
rect 1886 318 1887 322
rect 1891 318 1892 322
rect 1886 317 1892 318
rect 1966 322 1972 323
rect 1966 318 1967 322
rect 1971 318 1972 322
rect 1966 317 1972 318
rect 2054 322 2060 323
rect 2054 318 2055 322
rect 2059 318 2060 322
rect 2054 317 2060 318
rect 2142 322 2148 323
rect 2142 318 2143 322
rect 2147 318 2148 322
rect 2142 317 2148 318
rect 2230 322 2236 323
rect 2230 318 2231 322
rect 2235 318 2236 322
rect 2230 317 2236 318
rect 2310 322 2316 323
rect 2310 318 2311 322
rect 2315 318 2316 322
rect 2310 317 2316 318
rect 2390 322 2396 323
rect 2390 318 2391 322
rect 2395 318 2396 322
rect 2390 317 2396 318
rect 2478 322 2484 323
rect 2478 318 2479 322
rect 2483 318 2484 322
rect 2478 317 2484 318
rect 2542 322 2548 323
rect 2542 318 2543 322
rect 2547 318 2548 322
rect 2542 317 2548 318
rect 2584 314 2586 329
rect 110 313 116 314
rect 110 309 111 313
rect 115 309 116 313
rect 110 308 116 309
rect 1326 313 1332 314
rect 1326 309 1327 313
rect 1331 309 1332 313
rect 1326 308 1332 309
rect 1366 313 1372 314
rect 1366 309 1367 313
rect 1371 309 1372 313
rect 1366 308 1372 309
rect 2582 313 2588 314
rect 2582 309 2583 313
rect 2587 309 2588 313
rect 2582 308 2588 309
rect 110 296 116 297
rect 1326 296 1332 297
rect 110 292 111 296
rect 115 292 116 296
rect 110 291 116 292
rect 446 295 452 296
rect 446 291 447 295
rect 451 291 452 295
rect 112 275 114 291
rect 446 290 452 291
rect 502 295 508 296
rect 502 291 503 295
rect 507 291 508 295
rect 502 290 508 291
rect 558 295 564 296
rect 558 291 559 295
rect 563 291 564 295
rect 558 290 564 291
rect 614 295 620 296
rect 614 291 615 295
rect 619 291 620 295
rect 614 290 620 291
rect 678 295 684 296
rect 678 291 679 295
rect 683 291 684 295
rect 678 290 684 291
rect 750 295 756 296
rect 750 291 751 295
rect 755 291 756 295
rect 750 290 756 291
rect 830 295 836 296
rect 830 291 831 295
rect 835 291 836 295
rect 830 290 836 291
rect 910 295 916 296
rect 910 291 911 295
rect 915 291 916 295
rect 910 290 916 291
rect 998 295 1004 296
rect 998 291 999 295
rect 1003 291 1004 295
rect 998 290 1004 291
rect 1094 295 1100 296
rect 1094 291 1095 295
rect 1099 291 1100 295
rect 1094 290 1100 291
rect 1198 295 1204 296
rect 1198 291 1199 295
rect 1203 291 1204 295
rect 1326 292 1327 296
rect 1331 292 1332 296
rect 1326 291 1332 292
rect 1366 296 1372 297
rect 2582 296 2588 297
rect 1366 292 1367 296
rect 1371 292 1372 296
rect 1366 291 1372 292
rect 1614 295 1620 296
rect 1614 291 1615 295
rect 1619 291 1620 295
rect 1198 290 1204 291
rect 448 275 450 290
rect 504 275 506 290
rect 560 275 562 290
rect 616 275 618 290
rect 680 275 682 290
rect 752 275 754 290
rect 832 275 834 290
rect 912 275 914 290
rect 1000 275 1002 290
rect 1096 275 1098 290
rect 1200 275 1202 290
rect 1328 275 1330 291
rect 1368 279 1370 291
rect 1614 290 1620 291
rect 1670 295 1676 296
rect 1670 291 1671 295
rect 1675 291 1676 295
rect 1670 290 1676 291
rect 1726 295 1732 296
rect 1726 291 1727 295
rect 1731 291 1732 295
rect 1726 290 1732 291
rect 1790 295 1796 296
rect 1790 291 1791 295
rect 1795 291 1796 295
rect 1790 290 1796 291
rect 1870 295 1876 296
rect 1870 291 1871 295
rect 1875 291 1876 295
rect 1870 290 1876 291
rect 1950 295 1956 296
rect 1950 291 1951 295
rect 1955 291 1956 295
rect 1950 290 1956 291
rect 2038 295 2044 296
rect 2038 291 2039 295
rect 2043 291 2044 295
rect 2038 290 2044 291
rect 2126 295 2132 296
rect 2126 291 2127 295
rect 2131 291 2132 295
rect 2126 290 2132 291
rect 2214 295 2220 296
rect 2214 291 2215 295
rect 2219 291 2220 295
rect 2214 290 2220 291
rect 2294 295 2300 296
rect 2294 291 2295 295
rect 2299 291 2300 295
rect 2294 290 2300 291
rect 2374 295 2380 296
rect 2374 291 2375 295
rect 2379 291 2380 295
rect 2374 290 2380 291
rect 2462 295 2468 296
rect 2462 291 2463 295
rect 2467 291 2468 295
rect 2462 290 2468 291
rect 2526 295 2532 296
rect 2526 291 2527 295
rect 2531 291 2532 295
rect 2582 292 2583 296
rect 2587 292 2588 296
rect 2582 291 2588 292
rect 2526 290 2532 291
rect 1616 279 1618 290
rect 1672 279 1674 290
rect 1728 279 1730 290
rect 1792 279 1794 290
rect 1872 279 1874 290
rect 1952 279 1954 290
rect 2040 279 2042 290
rect 2128 279 2130 290
rect 2216 279 2218 290
rect 2296 279 2298 290
rect 2376 279 2378 290
rect 2464 279 2466 290
rect 2528 279 2530 290
rect 2584 279 2586 291
rect 1367 278 1371 279
rect 111 274 115 275
rect 111 269 115 270
rect 287 274 291 275
rect 287 269 291 270
rect 359 274 363 275
rect 359 269 363 270
rect 439 274 443 275
rect 439 269 443 270
rect 447 274 451 275
rect 447 269 451 270
rect 503 274 507 275
rect 503 269 507 270
rect 527 274 531 275
rect 527 269 531 270
rect 559 274 563 275
rect 559 269 563 270
rect 615 274 619 275
rect 615 269 619 270
rect 623 274 627 275
rect 623 269 627 270
rect 679 274 683 275
rect 679 269 683 270
rect 719 274 723 275
rect 719 269 723 270
rect 751 274 755 275
rect 751 269 755 270
rect 823 274 827 275
rect 823 269 827 270
rect 831 274 835 275
rect 831 269 835 270
rect 911 274 915 275
rect 911 269 915 270
rect 927 274 931 275
rect 927 269 931 270
rect 999 274 1003 275
rect 999 269 1003 270
rect 1031 274 1035 275
rect 1031 269 1035 270
rect 1095 274 1099 275
rect 1095 269 1099 270
rect 1143 274 1147 275
rect 1143 269 1147 270
rect 1199 274 1203 275
rect 1199 269 1203 270
rect 1255 274 1259 275
rect 1255 269 1259 270
rect 1327 274 1331 275
rect 1367 273 1371 274
rect 1535 278 1539 279
rect 1535 273 1539 274
rect 1607 278 1611 279
rect 1607 273 1611 274
rect 1615 278 1619 279
rect 1615 273 1619 274
rect 1671 278 1675 279
rect 1671 273 1675 274
rect 1687 278 1691 279
rect 1687 273 1691 274
rect 1727 278 1731 279
rect 1727 273 1731 274
rect 1775 278 1779 279
rect 1775 273 1779 274
rect 1791 278 1795 279
rect 1791 273 1795 274
rect 1863 278 1867 279
rect 1863 273 1867 274
rect 1871 278 1875 279
rect 1871 273 1875 274
rect 1951 278 1955 279
rect 1951 273 1955 274
rect 2039 278 2043 279
rect 2039 273 2043 274
rect 2119 278 2123 279
rect 2119 273 2123 274
rect 2127 278 2131 279
rect 2127 273 2131 274
rect 2199 278 2203 279
rect 2199 273 2203 274
rect 2215 278 2219 279
rect 2215 273 2219 274
rect 2271 278 2275 279
rect 2271 273 2275 274
rect 2295 278 2299 279
rect 2295 273 2299 274
rect 2335 278 2339 279
rect 2335 273 2339 274
rect 2375 278 2379 279
rect 2375 273 2379 274
rect 2407 278 2411 279
rect 2407 273 2411 274
rect 2463 278 2467 279
rect 2463 273 2467 274
rect 2471 278 2475 279
rect 2471 273 2475 274
rect 2527 278 2531 279
rect 2527 273 2531 274
rect 2583 278 2587 279
rect 2583 273 2587 274
rect 1327 269 1331 270
rect 112 257 114 269
rect 288 258 290 269
rect 360 258 362 269
rect 440 258 442 269
rect 528 258 530 269
rect 624 258 626 269
rect 720 258 722 269
rect 824 258 826 269
rect 928 258 930 269
rect 1032 258 1034 269
rect 1144 258 1146 269
rect 1256 258 1258 269
rect 286 257 292 258
rect 110 256 116 257
rect 110 252 111 256
rect 115 252 116 256
rect 286 253 287 257
rect 291 253 292 257
rect 286 252 292 253
rect 358 257 364 258
rect 358 253 359 257
rect 363 253 364 257
rect 358 252 364 253
rect 438 257 444 258
rect 438 253 439 257
rect 443 253 444 257
rect 438 252 444 253
rect 526 257 532 258
rect 526 253 527 257
rect 531 253 532 257
rect 526 252 532 253
rect 622 257 628 258
rect 622 253 623 257
rect 627 253 628 257
rect 622 252 628 253
rect 718 257 724 258
rect 718 253 719 257
rect 723 253 724 257
rect 718 252 724 253
rect 822 257 828 258
rect 822 253 823 257
rect 827 253 828 257
rect 822 252 828 253
rect 926 257 932 258
rect 926 253 927 257
rect 931 253 932 257
rect 926 252 932 253
rect 1030 257 1036 258
rect 1030 253 1031 257
rect 1035 253 1036 257
rect 1030 252 1036 253
rect 1142 257 1148 258
rect 1142 253 1143 257
rect 1147 253 1148 257
rect 1142 252 1148 253
rect 1254 257 1260 258
rect 1328 257 1330 269
rect 1368 261 1370 273
rect 1536 262 1538 273
rect 1608 262 1610 273
rect 1688 262 1690 273
rect 1776 262 1778 273
rect 1864 262 1866 273
rect 1952 262 1954 273
rect 2040 262 2042 273
rect 2120 262 2122 273
rect 2200 262 2202 273
rect 2272 262 2274 273
rect 2336 262 2338 273
rect 2408 262 2410 273
rect 2472 262 2474 273
rect 2528 262 2530 273
rect 1534 261 1540 262
rect 1366 260 1372 261
rect 1254 253 1255 257
rect 1259 253 1260 257
rect 1254 252 1260 253
rect 1326 256 1332 257
rect 1326 252 1327 256
rect 1331 252 1332 256
rect 1366 256 1367 260
rect 1371 256 1372 260
rect 1534 257 1535 261
rect 1539 257 1540 261
rect 1534 256 1540 257
rect 1606 261 1612 262
rect 1606 257 1607 261
rect 1611 257 1612 261
rect 1606 256 1612 257
rect 1686 261 1692 262
rect 1686 257 1687 261
rect 1691 257 1692 261
rect 1686 256 1692 257
rect 1774 261 1780 262
rect 1774 257 1775 261
rect 1779 257 1780 261
rect 1774 256 1780 257
rect 1862 261 1868 262
rect 1862 257 1863 261
rect 1867 257 1868 261
rect 1862 256 1868 257
rect 1950 261 1956 262
rect 1950 257 1951 261
rect 1955 257 1956 261
rect 1950 256 1956 257
rect 2038 261 2044 262
rect 2038 257 2039 261
rect 2043 257 2044 261
rect 2038 256 2044 257
rect 2118 261 2124 262
rect 2118 257 2119 261
rect 2123 257 2124 261
rect 2118 256 2124 257
rect 2198 261 2204 262
rect 2198 257 2199 261
rect 2203 257 2204 261
rect 2198 256 2204 257
rect 2270 261 2276 262
rect 2270 257 2271 261
rect 2275 257 2276 261
rect 2270 256 2276 257
rect 2334 261 2340 262
rect 2334 257 2335 261
rect 2339 257 2340 261
rect 2334 256 2340 257
rect 2406 261 2412 262
rect 2406 257 2407 261
rect 2411 257 2412 261
rect 2406 256 2412 257
rect 2470 261 2476 262
rect 2470 257 2471 261
rect 2475 257 2476 261
rect 2470 256 2476 257
rect 2526 261 2532 262
rect 2584 261 2586 273
rect 2526 257 2527 261
rect 2531 257 2532 261
rect 2526 256 2532 257
rect 2582 260 2588 261
rect 2582 256 2583 260
rect 2587 256 2588 260
rect 1366 255 1372 256
rect 2582 255 2588 256
rect 110 251 116 252
rect 1326 251 1332 252
rect 1366 243 1372 244
rect 110 239 116 240
rect 110 235 111 239
rect 115 235 116 239
rect 110 234 116 235
rect 1326 239 1332 240
rect 1326 235 1327 239
rect 1331 235 1332 239
rect 1366 239 1367 243
rect 1371 239 1372 243
rect 1366 238 1372 239
rect 2582 243 2588 244
rect 2582 239 2583 243
rect 2587 239 2588 243
rect 2582 238 2588 239
rect 1326 234 1332 235
rect 112 219 114 234
rect 302 230 308 231
rect 302 226 303 230
rect 307 226 308 230
rect 302 225 308 226
rect 374 230 380 231
rect 374 226 375 230
rect 379 226 380 230
rect 374 225 380 226
rect 454 230 460 231
rect 454 226 455 230
rect 459 226 460 230
rect 454 225 460 226
rect 542 230 548 231
rect 542 226 543 230
rect 547 226 548 230
rect 542 225 548 226
rect 638 230 644 231
rect 638 226 639 230
rect 643 226 644 230
rect 638 225 644 226
rect 734 230 740 231
rect 734 226 735 230
rect 739 226 740 230
rect 734 225 740 226
rect 838 230 844 231
rect 838 226 839 230
rect 843 226 844 230
rect 838 225 844 226
rect 942 230 948 231
rect 942 226 943 230
rect 947 226 948 230
rect 942 225 948 226
rect 1046 230 1052 231
rect 1046 226 1047 230
rect 1051 226 1052 230
rect 1046 225 1052 226
rect 1158 230 1164 231
rect 1158 226 1159 230
rect 1163 226 1164 230
rect 1158 225 1164 226
rect 1270 230 1276 231
rect 1270 226 1271 230
rect 1275 226 1276 230
rect 1270 225 1276 226
rect 304 219 306 225
rect 376 219 378 225
rect 456 219 458 225
rect 544 219 546 225
rect 640 219 642 225
rect 736 219 738 225
rect 840 219 842 225
rect 944 219 946 225
rect 1048 219 1050 225
rect 1160 219 1162 225
rect 1272 219 1274 225
rect 1328 219 1330 234
rect 1368 223 1370 238
rect 1550 234 1556 235
rect 1550 230 1551 234
rect 1555 230 1556 234
rect 1550 229 1556 230
rect 1622 234 1628 235
rect 1622 230 1623 234
rect 1627 230 1628 234
rect 1622 229 1628 230
rect 1702 234 1708 235
rect 1702 230 1703 234
rect 1707 230 1708 234
rect 1702 229 1708 230
rect 1790 234 1796 235
rect 1790 230 1791 234
rect 1795 230 1796 234
rect 1790 229 1796 230
rect 1878 234 1884 235
rect 1878 230 1879 234
rect 1883 230 1884 234
rect 1878 229 1884 230
rect 1966 234 1972 235
rect 1966 230 1967 234
rect 1971 230 1972 234
rect 1966 229 1972 230
rect 2054 234 2060 235
rect 2054 230 2055 234
rect 2059 230 2060 234
rect 2054 229 2060 230
rect 2134 234 2140 235
rect 2134 230 2135 234
rect 2139 230 2140 234
rect 2134 229 2140 230
rect 2214 234 2220 235
rect 2214 230 2215 234
rect 2219 230 2220 234
rect 2214 229 2220 230
rect 2286 234 2292 235
rect 2286 230 2287 234
rect 2291 230 2292 234
rect 2286 229 2292 230
rect 2350 234 2356 235
rect 2350 230 2351 234
rect 2355 230 2356 234
rect 2350 229 2356 230
rect 2422 234 2428 235
rect 2422 230 2423 234
rect 2427 230 2428 234
rect 2422 229 2428 230
rect 2486 234 2492 235
rect 2486 230 2487 234
rect 2491 230 2492 234
rect 2486 229 2492 230
rect 2542 234 2548 235
rect 2542 230 2543 234
rect 2547 230 2548 234
rect 2542 229 2548 230
rect 1552 223 1554 229
rect 1624 223 1626 229
rect 1704 223 1706 229
rect 1792 223 1794 229
rect 1880 223 1882 229
rect 1968 223 1970 229
rect 2056 223 2058 229
rect 2136 223 2138 229
rect 2216 223 2218 229
rect 2288 223 2290 229
rect 2352 223 2354 229
rect 2424 223 2426 229
rect 2488 223 2490 229
rect 2544 223 2546 229
rect 2584 223 2586 238
rect 1367 222 1371 223
rect 111 218 115 219
rect 111 213 115 214
rect 199 218 203 219
rect 199 213 203 214
rect 271 218 275 219
rect 271 213 275 214
rect 303 218 307 219
rect 303 213 307 214
rect 359 218 363 219
rect 359 213 363 214
rect 375 218 379 219
rect 375 213 379 214
rect 455 218 459 219
rect 455 213 459 214
rect 463 218 467 219
rect 463 213 467 214
rect 543 218 547 219
rect 543 213 547 214
rect 567 218 571 219
rect 567 213 571 214
rect 639 218 643 219
rect 639 213 643 214
rect 679 218 683 219
rect 679 213 683 214
rect 735 218 739 219
rect 735 213 739 214
rect 791 218 795 219
rect 791 213 795 214
rect 839 218 843 219
rect 839 213 843 214
rect 911 218 915 219
rect 911 213 915 214
rect 943 218 947 219
rect 943 213 947 214
rect 1031 218 1035 219
rect 1031 213 1035 214
rect 1047 218 1051 219
rect 1047 213 1051 214
rect 1151 218 1155 219
rect 1151 213 1155 214
rect 1159 218 1163 219
rect 1159 213 1163 214
rect 1271 218 1275 219
rect 1271 213 1275 214
rect 1327 218 1331 219
rect 1367 217 1371 218
rect 1415 222 1419 223
rect 1415 217 1419 218
rect 1479 222 1483 223
rect 1479 217 1483 218
rect 1551 222 1555 223
rect 1551 217 1555 218
rect 1559 222 1563 223
rect 1559 217 1563 218
rect 1623 222 1627 223
rect 1623 217 1627 218
rect 1655 222 1659 223
rect 1655 217 1659 218
rect 1703 222 1707 223
rect 1703 217 1707 218
rect 1751 222 1755 223
rect 1751 217 1755 218
rect 1791 222 1795 223
rect 1791 217 1795 218
rect 1855 222 1859 223
rect 1855 217 1859 218
rect 1879 222 1883 223
rect 1879 217 1883 218
rect 1959 222 1963 223
rect 1959 217 1963 218
rect 1967 222 1971 223
rect 1967 217 1971 218
rect 2055 222 2059 223
rect 2055 217 2059 218
rect 2063 222 2067 223
rect 2063 217 2067 218
rect 2135 222 2139 223
rect 2135 217 2139 218
rect 2167 222 2171 223
rect 2167 217 2171 218
rect 2215 222 2219 223
rect 2215 217 2219 218
rect 2263 222 2267 223
rect 2263 217 2267 218
rect 2287 222 2291 223
rect 2287 217 2291 218
rect 2351 222 2355 223
rect 2351 217 2355 218
rect 2359 222 2363 223
rect 2359 217 2363 218
rect 2423 222 2427 223
rect 2423 217 2427 218
rect 2463 222 2467 223
rect 2463 217 2467 218
rect 2487 222 2491 223
rect 2487 217 2491 218
rect 2543 222 2547 223
rect 2543 217 2547 218
rect 2583 222 2587 223
rect 2583 217 2587 218
rect 1327 213 1331 214
rect 112 198 114 213
rect 200 207 202 213
rect 272 207 274 213
rect 360 207 362 213
rect 464 207 466 213
rect 568 207 570 213
rect 680 207 682 213
rect 792 207 794 213
rect 912 207 914 213
rect 1032 207 1034 213
rect 1152 207 1154 213
rect 1272 207 1274 213
rect 198 206 204 207
rect 198 202 199 206
rect 203 202 204 206
rect 198 201 204 202
rect 270 206 276 207
rect 270 202 271 206
rect 275 202 276 206
rect 270 201 276 202
rect 358 206 364 207
rect 358 202 359 206
rect 363 202 364 206
rect 358 201 364 202
rect 462 206 468 207
rect 462 202 463 206
rect 467 202 468 206
rect 462 201 468 202
rect 566 206 572 207
rect 566 202 567 206
rect 571 202 572 206
rect 566 201 572 202
rect 678 206 684 207
rect 678 202 679 206
rect 683 202 684 206
rect 678 201 684 202
rect 790 206 796 207
rect 790 202 791 206
rect 795 202 796 206
rect 790 201 796 202
rect 910 206 916 207
rect 910 202 911 206
rect 915 202 916 206
rect 910 201 916 202
rect 1030 206 1036 207
rect 1030 202 1031 206
rect 1035 202 1036 206
rect 1030 201 1036 202
rect 1150 206 1156 207
rect 1150 202 1151 206
rect 1155 202 1156 206
rect 1150 201 1156 202
rect 1270 206 1276 207
rect 1270 202 1271 206
rect 1275 202 1276 206
rect 1270 201 1276 202
rect 1328 198 1330 213
rect 1368 202 1370 217
rect 1416 211 1418 217
rect 1480 211 1482 217
rect 1560 211 1562 217
rect 1656 211 1658 217
rect 1752 211 1754 217
rect 1856 211 1858 217
rect 1960 211 1962 217
rect 2064 211 2066 217
rect 2168 211 2170 217
rect 2264 211 2266 217
rect 2360 211 2362 217
rect 2464 211 2466 217
rect 2544 211 2546 217
rect 1414 210 1420 211
rect 1414 206 1415 210
rect 1419 206 1420 210
rect 1414 205 1420 206
rect 1478 210 1484 211
rect 1478 206 1479 210
rect 1483 206 1484 210
rect 1478 205 1484 206
rect 1558 210 1564 211
rect 1558 206 1559 210
rect 1563 206 1564 210
rect 1558 205 1564 206
rect 1654 210 1660 211
rect 1654 206 1655 210
rect 1659 206 1660 210
rect 1654 205 1660 206
rect 1750 210 1756 211
rect 1750 206 1751 210
rect 1755 206 1756 210
rect 1750 205 1756 206
rect 1854 210 1860 211
rect 1854 206 1855 210
rect 1859 206 1860 210
rect 1854 205 1860 206
rect 1958 210 1964 211
rect 1958 206 1959 210
rect 1963 206 1964 210
rect 1958 205 1964 206
rect 2062 210 2068 211
rect 2062 206 2063 210
rect 2067 206 2068 210
rect 2062 205 2068 206
rect 2166 210 2172 211
rect 2166 206 2167 210
rect 2171 206 2172 210
rect 2166 205 2172 206
rect 2262 210 2268 211
rect 2262 206 2263 210
rect 2267 206 2268 210
rect 2262 205 2268 206
rect 2358 210 2364 211
rect 2358 206 2359 210
rect 2363 206 2364 210
rect 2358 205 2364 206
rect 2462 210 2468 211
rect 2462 206 2463 210
rect 2467 206 2468 210
rect 2462 205 2468 206
rect 2542 210 2548 211
rect 2542 206 2543 210
rect 2547 206 2548 210
rect 2542 205 2548 206
rect 2584 202 2586 217
rect 1366 201 1372 202
rect 110 197 116 198
rect 110 193 111 197
rect 115 193 116 197
rect 110 192 116 193
rect 1326 197 1332 198
rect 1326 193 1327 197
rect 1331 193 1332 197
rect 1366 197 1367 201
rect 1371 197 1372 201
rect 1366 196 1372 197
rect 2582 201 2588 202
rect 2582 197 2583 201
rect 2587 197 2588 201
rect 2582 196 2588 197
rect 1326 192 1332 193
rect 1366 184 1372 185
rect 2582 184 2588 185
rect 110 180 116 181
rect 1326 180 1332 181
rect 110 176 111 180
rect 115 176 116 180
rect 110 175 116 176
rect 182 179 188 180
rect 182 175 183 179
rect 187 175 188 179
rect 112 139 114 175
rect 182 174 188 175
rect 254 179 260 180
rect 254 175 255 179
rect 259 175 260 179
rect 254 174 260 175
rect 342 179 348 180
rect 342 175 343 179
rect 347 175 348 179
rect 342 174 348 175
rect 446 179 452 180
rect 446 175 447 179
rect 451 175 452 179
rect 446 174 452 175
rect 550 179 556 180
rect 550 175 551 179
rect 555 175 556 179
rect 550 174 556 175
rect 662 179 668 180
rect 662 175 663 179
rect 667 175 668 179
rect 662 174 668 175
rect 774 179 780 180
rect 774 175 775 179
rect 779 175 780 179
rect 774 174 780 175
rect 894 179 900 180
rect 894 175 895 179
rect 899 175 900 179
rect 894 174 900 175
rect 1014 179 1020 180
rect 1014 175 1015 179
rect 1019 175 1020 179
rect 1014 174 1020 175
rect 1134 179 1140 180
rect 1134 175 1135 179
rect 1139 175 1140 179
rect 1134 174 1140 175
rect 1254 179 1260 180
rect 1254 175 1255 179
rect 1259 175 1260 179
rect 1326 176 1327 180
rect 1331 176 1332 180
rect 1366 180 1367 184
rect 1371 180 1372 184
rect 1366 179 1372 180
rect 1398 183 1404 184
rect 1398 179 1399 183
rect 1403 179 1404 183
rect 1326 175 1332 176
rect 1254 174 1260 175
rect 184 139 186 174
rect 256 139 258 174
rect 344 139 346 174
rect 448 139 450 174
rect 552 139 554 174
rect 664 139 666 174
rect 776 139 778 174
rect 896 139 898 174
rect 1016 139 1018 174
rect 1136 139 1138 174
rect 1256 139 1258 174
rect 1328 139 1330 175
rect 1368 151 1370 179
rect 1398 178 1404 179
rect 1462 183 1468 184
rect 1462 179 1463 183
rect 1467 179 1468 183
rect 1462 178 1468 179
rect 1542 183 1548 184
rect 1542 179 1543 183
rect 1547 179 1548 183
rect 1542 178 1548 179
rect 1638 183 1644 184
rect 1638 179 1639 183
rect 1643 179 1644 183
rect 1638 178 1644 179
rect 1734 183 1740 184
rect 1734 179 1735 183
rect 1739 179 1740 183
rect 1734 178 1740 179
rect 1838 183 1844 184
rect 1838 179 1839 183
rect 1843 179 1844 183
rect 1838 178 1844 179
rect 1942 183 1948 184
rect 1942 179 1943 183
rect 1947 179 1948 183
rect 1942 178 1948 179
rect 2046 183 2052 184
rect 2046 179 2047 183
rect 2051 179 2052 183
rect 2046 178 2052 179
rect 2150 183 2156 184
rect 2150 179 2151 183
rect 2155 179 2156 183
rect 2150 178 2156 179
rect 2246 183 2252 184
rect 2246 179 2247 183
rect 2251 179 2252 183
rect 2246 178 2252 179
rect 2342 183 2348 184
rect 2342 179 2343 183
rect 2347 179 2348 183
rect 2342 178 2348 179
rect 2446 183 2452 184
rect 2446 179 2447 183
rect 2451 179 2452 183
rect 2446 178 2452 179
rect 2526 183 2532 184
rect 2526 179 2527 183
rect 2531 179 2532 183
rect 2582 180 2583 184
rect 2587 180 2588 184
rect 2582 179 2588 180
rect 2526 178 2532 179
rect 1400 151 1402 178
rect 1464 151 1466 178
rect 1544 151 1546 178
rect 1640 151 1642 178
rect 1736 151 1738 178
rect 1840 151 1842 178
rect 1944 151 1946 178
rect 2048 151 2050 178
rect 2152 151 2154 178
rect 2248 151 2250 178
rect 2344 151 2346 178
rect 2448 151 2450 178
rect 2528 151 2530 178
rect 2584 151 2586 179
rect 1367 150 1371 151
rect 1367 145 1371 146
rect 1399 150 1403 151
rect 1399 145 1403 146
rect 1455 150 1459 151
rect 1455 145 1459 146
rect 1463 150 1467 151
rect 1463 145 1467 146
rect 1511 150 1515 151
rect 1511 145 1515 146
rect 1543 150 1547 151
rect 1543 145 1547 146
rect 1567 150 1571 151
rect 1567 145 1571 146
rect 1631 150 1635 151
rect 1631 145 1635 146
rect 1639 150 1643 151
rect 1639 145 1643 146
rect 1711 150 1715 151
rect 1711 145 1715 146
rect 1735 150 1739 151
rect 1735 145 1739 146
rect 1791 150 1795 151
rect 1791 145 1795 146
rect 1839 150 1843 151
rect 1839 145 1843 146
rect 1871 150 1875 151
rect 1871 145 1875 146
rect 1943 150 1947 151
rect 1943 145 1947 146
rect 2015 150 2019 151
rect 2015 145 2019 146
rect 2047 150 2051 151
rect 2047 145 2051 146
rect 2079 150 2083 151
rect 2079 145 2083 146
rect 2143 150 2147 151
rect 2143 145 2147 146
rect 2151 150 2155 151
rect 2151 145 2155 146
rect 2207 150 2211 151
rect 2207 145 2211 146
rect 2247 150 2251 151
rect 2247 145 2251 146
rect 2271 150 2275 151
rect 2271 145 2275 146
rect 2343 150 2347 151
rect 2343 145 2347 146
rect 2415 150 2419 151
rect 2415 145 2419 146
rect 2447 150 2451 151
rect 2447 145 2451 146
rect 2527 150 2531 151
rect 2527 145 2531 146
rect 2583 150 2587 151
rect 2583 145 2587 146
rect 111 138 115 139
rect 111 133 115 134
rect 143 138 147 139
rect 143 133 147 134
rect 183 138 187 139
rect 183 133 187 134
rect 199 138 203 139
rect 199 133 203 134
rect 255 138 259 139
rect 255 133 259 134
rect 311 138 315 139
rect 311 133 315 134
rect 343 138 347 139
rect 343 133 347 134
rect 367 138 371 139
rect 367 133 371 134
rect 423 138 427 139
rect 423 133 427 134
rect 447 138 451 139
rect 447 133 451 134
rect 479 138 483 139
rect 479 133 483 134
rect 535 138 539 139
rect 535 133 539 134
rect 551 138 555 139
rect 551 133 555 134
rect 591 138 595 139
rect 591 133 595 134
rect 647 138 651 139
rect 647 133 651 134
rect 663 138 667 139
rect 663 133 667 134
rect 703 138 707 139
rect 703 133 707 134
rect 759 138 763 139
rect 759 133 763 134
rect 775 138 779 139
rect 775 133 779 134
rect 823 138 827 139
rect 823 133 827 134
rect 887 138 891 139
rect 887 133 891 134
rect 895 138 899 139
rect 895 133 899 134
rect 951 138 955 139
rect 951 133 955 134
rect 1015 138 1019 139
rect 1015 133 1019 134
rect 1079 138 1083 139
rect 1079 133 1083 134
rect 1135 138 1139 139
rect 1135 133 1139 134
rect 1151 138 1155 139
rect 1151 133 1155 134
rect 1215 138 1219 139
rect 1215 133 1219 134
rect 1255 138 1259 139
rect 1255 133 1259 134
rect 1271 138 1275 139
rect 1271 133 1275 134
rect 1327 138 1331 139
rect 1327 133 1331 134
rect 1368 133 1370 145
rect 1400 134 1402 145
rect 1456 134 1458 145
rect 1512 134 1514 145
rect 1568 134 1570 145
rect 1632 134 1634 145
rect 1712 134 1714 145
rect 1792 134 1794 145
rect 1872 134 1874 145
rect 1944 134 1946 145
rect 2016 134 2018 145
rect 2080 134 2082 145
rect 2144 134 2146 145
rect 2208 134 2210 145
rect 2272 134 2274 145
rect 2344 134 2346 145
rect 2416 134 2418 145
rect 1398 133 1404 134
rect 112 121 114 133
rect 144 122 146 133
rect 200 122 202 133
rect 256 122 258 133
rect 312 122 314 133
rect 368 122 370 133
rect 424 122 426 133
rect 480 122 482 133
rect 536 122 538 133
rect 592 122 594 133
rect 648 122 650 133
rect 704 122 706 133
rect 760 122 762 133
rect 824 122 826 133
rect 888 122 890 133
rect 952 122 954 133
rect 1016 122 1018 133
rect 1080 122 1082 133
rect 1152 122 1154 133
rect 1216 122 1218 133
rect 1272 122 1274 133
rect 142 121 148 122
rect 110 120 116 121
rect 110 116 111 120
rect 115 116 116 120
rect 142 117 143 121
rect 147 117 148 121
rect 142 116 148 117
rect 198 121 204 122
rect 198 117 199 121
rect 203 117 204 121
rect 198 116 204 117
rect 254 121 260 122
rect 254 117 255 121
rect 259 117 260 121
rect 254 116 260 117
rect 310 121 316 122
rect 310 117 311 121
rect 315 117 316 121
rect 310 116 316 117
rect 366 121 372 122
rect 366 117 367 121
rect 371 117 372 121
rect 366 116 372 117
rect 422 121 428 122
rect 422 117 423 121
rect 427 117 428 121
rect 422 116 428 117
rect 478 121 484 122
rect 478 117 479 121
rect 483 117 484 121
rect 478 116 484 117
rect 534 121 540 122
rect 534 117 535 121
rect 539 117 540 121
rect 534 116 540 117
rect 590 121 596 122
rect 590 117 591 121
rect 595 117 596 121
rect 590 116 596 117
rect 646 121 652 122
rect 646 117 647 121
rect 651 117 652 121
rect 646 116 652 117
rect 702 121 708 122
rect 702 117 703 121
rect 707 117 708 121
rect 702 116 708 117
rect 758 121 764 122
rect 758 117 759 121
rect 763 117 764 121
rect 758 116 764 117
rect 822 121 828 122
rect 822 117 823 121
rect 827 117 828 121
rect 822 116 828 117
rect 886 121 892 122
rect 886 117 887 121
rect 891 117 892 121
rect 886 116 892 117
rect 950 121 956 122
rect 950 117 951 121
rect 955 117 956 121
rect 950 116 956 117
rect 1014 121 1020 122
rect 1014 117 1015 121
rect 1019 117 1020 121
rect 1014 116 1020 117
rect 1078 121 1084 122
rect 1078 117 1079 121
rect 1083 117 1084 121
rect 1078 116 1084 117
rect 1150 121 1156 122
rect 1150 117 1151 121
rect 1155 117 1156 121
rect 1150 116 1156 117
rect 1214 121 1220 122
rect 1214 117 1215 121
rect 1219 117 1220 121
rect 1214 116 1220 117
rect 1270 121 1276 122
rect 1328 121 1330 133
rect 1366 132 1372 133
rect 1366 128 1367 132
rect 1371 128 1372 132
rect 1398 129 1399 133
rect 1403 129 1404 133
rect 1398 128 1404 129
rect 1454 133 1460 134
rect 1454 129 1455 133
rect 1459 129 1460 133
rect 1454 128 1460 129
rect 1510 133 1516 134
rect 1510 129 1511 133
rect 1515 129 1516 133
rect 1510 128 1516 129
rect 1566 133 1572 134
rect 1566 129 1567 133
rect 1571 129 1572 133
rect 1566 128 1572 129
rect 1630 133 1636 134
rect 1630 129 1631 133
rect 1635 129 1636 133
rect 1630 128 1636 129
rect 1710 133 1716 134
rect 1710 129 1711 133
rect 1715 129 1716 133
rect 1710 128 1716 129
rect 1790 133 1796 134
rect 1790 129 1791 133
rect 1795 129 1796 133
rect 1790 128 1796 129
rect 1870 133 1876 134
rect 1870 129 1871 133
rect 1875 129 1876 133
rect 1870 128 1876 129
rect 1942 133 1948 134
rect 1942 129 1943 133
rect 1947 129 1948 133
rect 1942 128 1948 129
rect 2014 133 2020 134
rect 2014 129 2015 133
rect 2019 129 2020 133
rect 2014 128 2020 129
rect 2078 133 2084 134
rect 2078 129 2079 133
rect 2083 129 2084 133
rect 2078 128 2084 129
rect 2142 133 2148 134
rect 2142 129 2143 133
rect 2147 129 2148 133
rect 2142 128 2148 129
rect 2206 133 2212 134
rect 2206 129 2207 133
rect 2211 129 2212 133
rect 2206 128 2212 129
rect 2270 133 2276 134
rect 2270 129 2271 133
rect 2275 129 2276 133
rect 2270 128 2276 129
rect 2342 133 2348 134
rect 2342 129 2343 133
rect 2347 129 2348 133
rect 2342 128 2348 129
rect 2414 133 2420 134
rect 2584 133 2586 145
rect 2414 129 2415 133
rect 2419 129 2420 133
rect 2414 128 2420 129
rect 2582 132 2588 133
rect 2582 128 2583 132
rect 2587 128 2588 132
rect 1366 127 1372 128
rect 2582 127 2588 128
rect 1270 117 1271 121
rect 1275 117 1276 121
rect 1270 116 1276 117
rect 1326 120 1332 121
rect 1326 116 1327 120
rect 1331 116 1332 120
rect 110 115 116 116
rect 1326 115 1332 116
rect 1366 115 1372 116
rect 1366 111 1367 115
rect 1371 111 1372 115
rect 1366 110 1372 111
rect 2582 115 2588 116
rect 2582 111 2583 115
rect 2587 111 2588 115
rect 2582 110 2588 111
rect 110 103 116 104
rect 110 99 111 103
rect 115 99 116 103
rect 110 98 116 99
rect 1326 103 1332 104
rect 1326 99 1327 103
rect 1331 99 1332 103
rect 1326 98 1332 99
rect 112 83 114 98
rect 158 94 164 95
rect 158 90 159 94
rect 163 90 164 94
rect 158 89 164 90
rect 214 94 220 95
rect 214 90 215 94
rect 219 90 220 94
rect 214 89 220 90
rect 270 94 276 95
rect 270 90 271 94
rect 275 90 276 94
rect 270 89 276 90
rect 326 94 332 95
rect 326 90 327 94
rect 331 90 332 94
rect 326 89 332 90
rect 382 94 388 95
rect 382 90 383 94
rect 387 90 388 94
rect 382 89 388 90
rect 438 94 444 95
rect 438 90 439 94
rect 443 90 444 94
rect 438 89 444 90
rect 494 94 500 95
rect 494 90 495 94
rect 499 90 500 94
rect 494 89 500 90
rect 550 94 556 95
rect 550 90 551 94
rect 555 90 556 94
rect 550 89 556 90
rect 606 94 612 95
rect 606 90 607 94
rect 611 90 612 94
rect 606 89 612 90
rect 662 94 668 95
rect 662 90 663 94
rect 667 90 668 94
rect 662 89 668 90
rect 718 94 724 95
rect 718 90 719 94
rect 723 90 724 94
rect 718 89 724 90
rect 774 94 780 95
rect 774 90 775 94
rect 779 90 780 94
rect 774 89 780 90
rect 838 94 844 95
rect 838 90 839 94
rect 843 90 844 94
rect 838 89 844 90
rect 902 94 908 95
rect 902 90 903 94
rect 907 90 908 94
rect 902 89 908 90
rect 966 94 972 95
rect 966 90 967 94
rect 971 90 972 94
rect 966 89 972 90
rect 1030 94 1036 95
rect 1030 90 1031 94
rect 1035 90 1036 94
rect 1030 89 1036 90
rect 1094 94 1100 95
rect 1094 90 1095 94
rect 1099 90 1100 94
rect 1094 89 1100 90
rect 1166 94 1172 95
rect 1166 90 1167 94
rect 1171 90 1172 94
rect 1166 89 1172 90
rect 1230 94 1236 95
rect 1230 90 1231 94
rect 1235 90 1236 94
rect 1230 89 1236 90
rect 1286 94 1292 95
rect 1286 90 1287 94
rect 1291 90 1292 94
rect 1286 89 1292 90
rect 160 83 162 89
rect 216 83 218 89
rect 272 83 274 89
rect 328 83 330 89
rect 384 83 386 89
rect 440 83 442 89
rect 496 83 498 89
rect 552 83 554 89
rect 608 83 610 89
rect 664 83 666 89
rect 720 83 722 89
rect 776 83 778 89
rect 840 83 842 89
rect 904 83 906 89
rect 968 83 970 89
rect 1032 83 1034 89
rect 1096 83 1098 89
rect 1168 83 1170 89
rect 1232 83 1234 89
rect 1288 83 1290 89
rect 1328 83 1330 98
rect 1368 95 1370 110
rect 1414 106 1420 107
rect 1414 102 1415 106
rect 1419 102 1420 106
rect 1414 101 1420 102
rect 1470 106 1476 107
rect 1470 102 1471 106
rect 1475 102 1476 106
rect 1470 101 1476 102
rect 1526 106 1532 107
rect 1526 102 1527 106
rect 1531 102 1532 106
rect 1526 101 1532 102
rect 1582 106 1588 107
rect 1582 102 1583 106
rect 1587 102 1588 106
rect 1582 101 1588 102
rect 1646 106 1652 107
rect 1646 102 1647 106
rect 1651 102 1652 106
rect 1646 101 1652 102
rect 1726 106 1732 107
rect 1726 102 1727 106
rect 1731 102 1732 106
rect 1726 101 1732 102
rect 1806 106 1812 107
rect 1806 102 1807 106
rect 1811 102 1812 106
rect 1806 101 1812 102
rect 1886 106 1892 107
rect 1886 102 1887 106
rect 1891 102 1892 106
rect 1886 101 1892 102
rect 1958 106 1964 107
rect 1958 102 1959 106
rect 1963 102 1964 106
rect 1958 101 1964 102
rect 2030 106 2036 107
rect 2030 102 2031 106
rect 2035 102 2036 106
rect 2030 101 2036 102
rect 2094 106 2100 107
rect 2094 102 2095 106
rect 2099 102 2100 106
rect 2094 101 2100 102
rect 2158 106 2164 107
rect 2158 102 2159 106
rect 2163 102 2164 106
rect 2158 101 2164 102
rect 2222 106 2228 107
rect 2222 102 2223 106
rect 2227 102 2228 106
rect 2222 101 2228 102
rect 2286 106 2292 107
rect 2286 102 2287 106
rect 2291 102 2292 106
rect 2286 101 2292 102
rect 2358 106 2364 107
rect 2358 102 2359 106
rect 2363 102 2364 106
rect 2358 101 2364 102
rect 2430 106 2436 107
rect 2430 102 2431 106
rect 2435 102 2436 106
rect 2430 101 2436 102
rect 1416 95 1418 101
rect 1472 95 1474 101
rect 1528 95 1530 101
rect 1584 95 1586 101
rect 1648 95 1650 101
rect 1728 95 1730 101
rect 1808 95 1810 101
rect 1888 95 1890 101
rect 1960 95 1962 101
rect 2032 95 2034 101
rect 2096 95 2098 101
rect 2160 95 2162 101
rect 2224 95 2226 101
rect 2288 95 2290 101
rect 2360 95 2362 101
rect 2432 95 2434 101
rect 2584 95 2586 110
rect 1367 94 1371 95
rect 1367 89 1371 90
rect 1415 94 1419 95
rect 1415 89 1419 90
rect 1471 94 1475 95
rect 1471 89 1475 90
rect 1527 94 1531 95
rect 1527 89 1531 90
rect 1583 94 1587 95
rect 1583 89 1587 90
rect 1647 94 1651 95
rect 1647 89 1651 90
rect 1727 94 1731 95
rect 1727 89 1731 90
rect 1807 94 1811 95
rect 1807 89 1811 90
rect 1887 94 1891 95
rect 1887 89 1891 90
rect 1959 94 1963 95
rect 1959 89 1963 90
rect 2031 94 2035 95
rect 2031 89 2035 90
rect 2095 94 2099 95
rect 2095 89 2099 90
rect 2159 94 2163 95
rect 2159 89 2163 90
rect 2223 94 2227 95
rect 2223 89 2227 90
rect 2287 94 2291 95
rect 2287 89 2291 90
rect 2359 94 2363 95
rect 2359 89 2363 90
rect 2431 94 2435 95
rect 2431 89 2435 90
rect 2583 94 2587 95
rect 2583 89 2587 90
rect 111 82 115 83
rect 111 77 115 78
rect 159 82 163 83
rect 159 77 163 78
rect 215 82 219 83
rect 215 77 219 78
rect 271 82 275 83
rect 271 77 275 78
rect 327 82 331 83
rect 327 77 331 78
rect 383 82 387 83
rect 383 77 387 78
rect 439 82 443 83
rect 439 77 443 78
rect 495 82 499 83
rect 495 77 499 78
rect 551 82 555 83
rect 551 77 555 78
rect 607 82 611 83
rect 607 77 611 78
rect 663 82 667 83
rect 663 77 667 78
rect 719 82 723 83
rect 719 77 723 78
rect 775 82 779 83
rect 775 77 779 78
rect 839 82 843 83
rect 839 77 843 78
rect 903 82 907 83
rect 903 77 907 78
rect 967 82 971 83
rect 967 77 971 78
rect 1031 82 1035 83
rect 1031 77 1035 78
rect 1095 82 1099 83
rect 1095 77 1099 78
rect 1167 82 1171 83
rect 1167 77 1171 78
rect 1231 82 1235 83
rect 1231 77 1235 78
rect 1287 82 1291 83
rect 1287 77 1291 78
rect 1327 82 1331 83
rect 1327 77 1331 78
<< m4c >>
rect 111 2638 115 2642
rect 551 2638 555 2642
rect 607 2638 611 2642
rect 663 2638 667 2642
rect 719 2638 723 2642
rect 775 2638 779 2642
rect 1327 2638 1331 2642
rect 1367 2634 1371 2638
rect 1551 2634 1555 2638
rect 1607 2634 1611 2638
rect 1663 2634 1667 2638
rect 1719 2634 1723 2638
rect 1775 2634 1779 2638
rect 1831 2634 1835 2638
rect 1887 2634 1891 2638
rect 1943 2634 1947 2638
rect 1999 2634 2003 2638
rect 2055 2634 2059 2638
rect 2111 2634 2115 2638
rect 2167 2634 2171 2638
rect 2583 2634 2587 2638
rect 111 2582 115 2586
rect 215 2582 219 2586
rect 271 2582 275 2586
rect 327 2582 331 2586
rect 383 2582 387 2586
rect 439 2582 443 2586
rect 495 2582 499 2586
rect 535 2582 539 2586
rect 551 2582 555 2586
rect 591 2582 595 2586
rect 607 2582 611 2586
rect 647 2582 651 2586
rect 663 2582 667 2586
rect 703 2582 707 2586
rect 719 2582 723 2586
rect 759 2582 763 2586
rect 775 2582 779 2586
rect 831 2582 835 2586
rect 887 2582 891 2586
rect 943 2582 947 2586
rect 999 2582 1003 2586
rect 1055 2582 1059 2586
rect 1111 2582 1115 2586
rect 1327 2582 1331 2586
rect 1367 2578 1371 2582
rect 1439 2578 1443 2582
rect 1535 2578 1539 2582
rect 1543 2578 1547 2582
rect 1591 2578 1595 2582
rect 1647 2578 1651 2582
rect 1655 2578 1659 2582
rect 1703 2578 1707 2582
rect 1759 2578 1763 2582
rect 1767 2578 1771 2582
rect 1815 2578 1819 2582
rect 1871 2578 1875 2582
rect 1879 2578 1883 2582
rect 1927 2578 1931 2582
rect 1983 2578 1987 2582
rect 1991 2578 1995 2582
rect 2039 2578 2043 2582
rect 2095 2578 2099 2582
rect 2111 2578 2115 2582
rect 2151 2578 2155 2582
rect 2231 2578 2235 2582
rect 2351 2578 2355 2582
rect 2583 2578 2587 2582
rect 111 2522 115 2526
rect 231 2522 235 2526
rect 287 2522 291 2526
rect 343 2522 347 2526
rect 367 2522 371 2526
rect 399 2522 403 2526
rect 423 2522 427 2526
rect 455 2522 459 2526
rect 487 2522 491 2526
rect 511 2522 515 2526
rect 551 2522 555 2526
rect 567 2522 571 2526
rect 615 2522 619 2526
rect 623 2522 627 2526
rect 679 2522 683 2526
rect 735 2522 739 2526
rect 743 2522 747 2526
rect 791 2522 795 2526
rect 807 2522 811 2526
rect 847 2522 851 2526
rect 871 2522 875 2526
rect 903 2522 907 2526
rect 943 2522 947 2526
rect 959 2522 963 2526
rect 1015 2522 1019 2526
rect 1071 2522 1075 2526
rect 1127 2522 1131 2526
rect 1327 2522 1331 2526
rect 1367 2514 1371 2518
rect 1455 2514 1459 2518
rect 1551 2514 1555 2518
rect 1559 2514 1563 2518
rect 1631 2514 1635 2518
rect 1671 2514 1675 2518
rect 1719 2514 1723 2518
rect 1783 2514 1787 2518
rect 1807 2514 1811 2518
rect 1895 2514 1899 2518
rect 1903 2514 1907 2518
rect 1999 2514 2003 2518
rect 2007 2514 2011 2518
rect 2095 2514 2099 2518
rect 2127 2514 2131 2518
rect 2191 2514 2195 2518
rect 2247 2514 2251 2518
rect 2295 2514 2299 2518
rect 2367 2514 2371 2518
rect 2399 2514 2403 2518
rect 2583 2514 2587 2518
rect 111 2462 115 2466
rect 271 2462 275 2466
rect 335 2462 339 2466
rect 351 2462 355 2466
rect 399 2462 403 2466
rect 407 2462 411 2466
rect 471 2462 475 2466
rect 535 2462 539 2466
rect 551 2462 555 2466
rect 599 2462 603 2466
rect 631 2462 635 2466
rect 663 2462 667 2466
rect 711 2462 715 2466
rect 727 2462 731 2466
rect 783 2462 787 2466
rect 791 2462 795 2466
rect 855 2462 859 2466
rect 863 2462 867 2466
rect 927 2462 931 2466
rect 943 2462 947 2466
rect 999 2462 1003 2466
rect 1023 2462 1027 2466
rect 1327 2462 1331 2466
rect 1367 2458 1371 2462
rect 1535 2458 1539 2462
rect 1615 2458 1619 2462
rect 1647 2458 1651 2462
rect 1703 2458 1707 2462
rect 1767 2458 1771 2462
rect 1791 2458 1795 2462
rect 1839 2458 1843 2462
rect 1887 2458 1891 2462
rect 1911 2458 1915 2462
rect 1983 2458 1987 2462
rect 1991 2458 1995 2462
rect 2079 2458 2083 2462
rect 2167 2458 2171 2462
rect 2175 2458 2179 2462
rect 2263 2458 2267 2462
rect 2279 2458 2283 2462
rect 2359 2458 2363 2462
rect 2383 2458 2387 2462
rect 2455 2458 2459 2462
rect 2527 2458 2531 2462
rect 2583 2458 2587 2462
rect 111 2402 115 2406
rect 247 2402 251 2406
rect 287 2402 291 2406
rect 335 2402 339 2406
rect 351 2402 355 2406
rect 415 2402 419 2406
rect 431 2402 435 2406
rect 487 2402 491 2406
rect 527 2402 531 2406
rect 567 2402 571 2406
rect 631 2402 635 2406
rect 647 2402 651 2406
rect 727 2402 731 2406
rect 799 2402 803 2406
rect 823 2402 827 2406
rect 879 2402 883 2406
rect 919 2402 923 2406
rect 959 2402 963 2406
rect 1015 2402 1019 2406
rect 1039 2402 1043 2406
rect 1111 2402 1115 2406
rect 1327 2402 1331 2406
rect 1367 2398 1371 2402
rect 1455 2398 1459 2402
rect 1559 2398 1563 2402
rect 1663 2398 1667 2402
rect 1719 2398 1723 2402
rect 1759 2398 1763 2402
rect 1783 2398 1787 2402
rect 1855 2398 1859 2402
rect 1927 2398 1931 2402
rect 1943 2398 1947 2402
rect 2007 2398 2011 2402
rect 2039 2398 2043 2402
rect 2095 2398 2099 2402
rect 2135 2398 2139 2402
rect 2183 2398 2187 2402
rect 2231 2398 2235 2402
rect 2279 2398 2283 2402
rect 2335 2398 2339 2402
rect 2375 2398 2379 2402
rect 2447 2398 2451 2402
rect 2471 2398 2475 2402
rect 2543 2398 2547 2402
rect 2583 2398 2587 2402
rect 111 2346 115 2350
rect 159 2346 163 2350
rect 231 2346 235 2350
rect 263 2346 267 2350
rect 319 2346 323 2350
rect 375 2346 379 2350
rect 415 2346 419 2350
rect 487 2346 491 2350
rect 511 2346 515 2350
rect 599 2346 603 2350
rect 615 2346 619 2350
rect 711 2346 715 2350
rect 807 2346 811 2350
rect 815 2346 819 2350
rect 903 2346 907 2350
rect 911 2346 915 2350
rect 999 2346 1003 2350
rect 1007 2346 1011 2350
rect 1095 2346 1099 2350
rect 1103 2346 1107 2350
rect 1199 2346 1203 2350
rect 1327 2346 1331 2350
rect 1367 2342 1371 2346
rect 1399 2342 1403 2346
rect 1439 2342 1443 2346
rect 1455 2342 1459 2346
rect 1511 2342 1515 2346
rect 1543 2342 1547 2346
rect 1567 2342 1571 2346
rect 1639 2342 1643 2346
rect 1647 2342 1651 2346
rect 1727 2342 1731 2346
rect 1743 2342 1747 2346
rect 1823 2342 1827 2346
rect 1839 2342 1843 2346
rect 1927 2342 1931 2346
rect 1943 2342 1947 2346
rect 2023 2342 2027 2346
rect 2079 2342 2083 2346
rect 2119 2342 2123 2346
rect 2215 2342 2219 2346
rect 2223 2342 2227 2346
rect 2319 2342 2323 2346
rect 2383 2342 2387 2346
rect 2431 2342 2435 2346
rect 2527 2342 2531 2346
rect 2583 2342 2587 2346
rect 111 2286 115 2290
rect 159 2286 163 2290
rect 175 2286 179 2290
rect 247 2286 251 2290
rect 279 2286 283 2290
rect 375 2286 379 2290
rect 391 2286 395 2290
rect 503 2286 507 2290
rect 511 2286 515 2290
rect 615 2286 619 2290
rect 639 2286 643 2290
rect 727 2286 731 2290
rect 767 2286 771 2290
rect 831 2286 835 2290
rect 887 2286 891 2290
rect 927 2286 931 2290
rect 999 2286 1003 2290
rect 1023 2286 1027 2290
rect 1103 2286 1107 2290
rect 1119 2286 1123 2290
rect 1207 2286 1211 2290
rect 1215 2286 1219 2290
rect 1287 2286 1291 2290
rect 1327 2286 1331 2290
rect 1367 2278 1371 2282
rect 1415 2278 1419 2282
rect 1471 2278 1475 2282
rect 1495 2278 1499 2282
rect 1527 2278 1531 2282
rect 1583 2278 1587 2282
rect 1615 2278 1619 2282
rect 1655 2278 1659 2282
rect 1735 2278 1739 2282
rect 1743 2278 1747 2282
rect 1839 2278 1843 2282
rect 1855 2278 1859 2282
rect 1959 2278 1963 2282
rect 1967 2278 1971 2282
rect 2071 2278 2075 2282
rect 2095 2278 2099 2282
rect 2167 2278 2171 2282
rect 2239 2278 2243 2282
rect 2255 2278 2259 2282
rect 2335 2278 2339 2282
rect 2399 2278 2403 2282
rect 2407 2278 2411 2282
rect 2487 2278 2491 2282
rect 2543 2278 2547 2282
rect 2583 2278 2587 2282
rect 111 2222 115 2226
rect 143 2222 147 2226
rect 231 2222 235 2226
rect 359 2222 363 2226
rect 495 2222 499 2226
rect 623 2222 627 2226
rect 751 2222 755 2226
rect 871 2222 875 2226
rect 983 2222 987 2226
rect 1087 2222 1091 2226
rect 1191 2222 1195 2226
rect 1271 2222 1275 2226
rect 1327 2222 1331 2226
rect 1367 2210 1371 2214
rect 1399 2210 1403 2214
rect 1455 2210 1459 2214
rect 1479 2210 1483 2214
rect 1535 2210 1539 2214
rect 1599 2210 1603 2214
rect 1631 2210 1635 2214
rect 1719 2210 1723 2214
rect 1743 2210 1747 2214
rect 1839 2210 1843 2214
rect 1863 2210 1867 2214
rect 1951 2210 1955 2214
rect 1983 2210 1987 2214
rect 2055 2210 2059 2214
rect 2095 2210 2099 2214
rect 2151 2210 2155 2214
rect 2207 2210 2211 2214
rect 2239 2210 2243 2214
rect 2311 2210 2315 2214
rect 2319 2210 2323 2214
rect 2391 2210 2395 2214
rect 2423 2210 2427 2214
rect 2471 2210 2475 2214
rect 2527 2210 2531 2214
rect 2583 2210 2587 2214
rect 111 2162 115 2166
rect 159 2162 163 2166
rect 215 2162 219 2166
rect 247 2162 251 2166
rect 311 2162 315 2166
rect 375 2162 379 2166
rect 423 2162 427 2166
rect 511 2162 515 2166
rect 543 2162 547 2166
rect 639 2162 643 2166
rect 663 2162 667 2166
rect 767 2162 771 2166
rect 775 2162 779 2166
rect 879 2162 883 2166
rect 887 2162 891 2166
rect 975 2162 979 2166
rect 999 2162 1003 2166
rect 1071 2162 1075 2166
rect 1103 2162 1107 2166
rect 1167 2162 1171 2166
rect 1207 2162 1211 2166
rect 1271 2162 1275 2166
rect 1287 2162 1291 2166
rect 1327 2162 1331 2166
rect 1367 2154 1371 2158
rect 1471 2154 1475 2158
rect 1535 2154 1539 2158
rect 1551 2154 1555 2158
rect 1631 2154 1635 2158
rect 1647 2154 1651 2158
rect 1735 2154 1739 2158
rect 1759 2154 1763 2158
rect 1839 2154 1843 2158
rect 1879 2154 1883 2158
rect 1951 2154 1955 2158
rect 1999 2154 2003 2158
rect 2055 2154 2059 2158
rect 2111 2154 2115 2158
rect 2159 2154 2163 2158
rect 2223 2154 2227 2158
rect 2263 2154 2267 2158
rect 2327 2154 2331 2158
rect 2359 2154 2363 2158
rect 2439 2154 2443 2158
rect 2463 2154 2467 2158
rect 2543 2154 2547 2158
rect 2583 2154 2587 2158
rect 111 2098 115 2102
rect 143 2098 147 2102
rect 199 2098 203 2102
rect 263 2098 267 2102
rect 295 2098 299 2102
rect 327 2098 331 2102
rect 399 2098 403 2102
rect 407 2098 411 2102
rect 479 2098 483 2102
rect 527 2098 531 2102
rect 567 2098 571 2102
rect 647 2098 651 2102
rect 655 2098 659 2102
rect 735 2098 739 2102
rect 759 2098 763 2102
rect 815 2098 819 2102
rect 863 2098 867 2102
rect 887 2098 891 2102
rect 959 2098 963 2102
rect 967 2098 971 2102
rect 1047 2098 1051 2102
rect 1055 2098 1059 2102
rect 1127 2098 1131 2102
rect 1151 2098 1155 2102
rect 1255 2098 1259 2102
rect 1327 2098 1331 2102
rect 1367 2098 1371 2102
rect 1431 2098 1435 2102
rect 1519 2098 1523 2102
rect 1535 2098 1539 2102
rect 1615 2098 1619 2102
rect 1647 2098 1651 2102
rect 1719 2098 1723 2102
rect 1759 2098 1763 2102
rect 1823 2098 1827 2102
rect 1863 2098 1867 2102
rect 1935 2098 1939 2102
rect 1967 2098 1971 2102
rect 2039 2098 2043 2102
rect 2071 2098 2075 2102
rect 2143 2098 2147 2102
rect 2175 2098 2179 2102
rect 2247 2098 2251 2102
rect 2271 2098 2275 2102
rect 2343 2098 2347 2102
rect 2359 2098 2363 2102
rect 2447 2098 2451 2102
rect 2455 2098 2459 2102
rect 2527 2098 2531 2102
rect 2583 2098 2587 2102
rect 1367 2042 1371 2046
rect 1415 2042 1419 2046
rect 1447 2042 1451 2046
rect 1503 2042 1507 2046
rect 1551 2042 1555 2046
rect 1607 2042 1611 2046
rect 1663 2042 1667 2046
rect 1711 2042 1715 2046
rect 1775 2042 1779 2046
rect 1807 2042 1811 2046
rect 1879 2042 1883 2046
rect 1903 2042 1907 2046
rect 1983 2042 1987 2046
rect 2007 2042 2011 2046
rect 2087 2042 2091 2046
rect 2111 2042 2115 2046
rect 2191 2042 2195 2046
rect 2215 2042 2219 2046
rect 2287 2042 2291 2046
rect 2327 2042 2331 2046
rect 2375 2042 2379 2046
rect 2447 2042 2451 2046
rect 2471 2042 2475 2046
rect 2543 2042 2547 2046
rect 2583 2042 2587 2046
rect 111 2034 115 2038
rect 279 2034 283 2038
rect 343 2034 347 2038
rect 415 2034 419 2038
rect 471 2034 475 2038
rect 495 2034 499 2038
rect 527 2034 531 2038
rect 583 2034 587 2038
rect 639 2034 643 2038
rect 671 2034 675 2038
rect 695 2034 699 2038
rect 751 2034 755 2038
rect 807 2034 811 2038
rect 831 2034 835 2038
rect 863 2034 867 2038
rect 903 2034 907 2038
rect 919 2034 923 2038
rect 975 2034 979 2038
rect 983 2034 987 2038
rect 1031 2034 1035 2038
rect 1063 2034 1067 2038
rect 1143 2034 1147 2038
rect 1327 2034 1331 2038
rect 1367 1986 1371 1990
rect 1399 1986 1403 1990
rect 1479 1986 1483 1990
rect 1487 1986 1491 1990
rect 1583 1986 1587 1990
rect 1591 1986 1595 1990
rect 1679 1986 1683 1990
rect 1695 1986 1699 1990
rect 1767 1986 1771 1990
rect 1791 1986 1795 1990
rect 1847 1986 1851 1990
rect 1887 1986 1891 1990
rect 1927 1986 1931 1990
rect 1991 1986 1995 1990
rect 2007 1986 2011 1990
rect 2087 1986 2091 1990
rect 2095 1986 2099 1990
rect 2199 1986 2203 1990
rect 2311 1986 2315 1990
rect 2431 1986 2435 1990
rect 2527 1986 2531 1990
rect 2583 1986 2587 1990
rect 111 1974 115 1978
rect 335 1974 339 1978
rect 391 1974 395 1978
rect 399 1974 403 1978
rect 447 1974 451 1978
rect 455 1974 459 1978
rect 503 1974 507 1978
rect 511 1974 515 1978
rect 567 1974 571 1978
rect 623 1974 627 1978
rect 647 1974 651 1978
rect 679 1974 683 1978
rect 735 1974 739 1978
rect 743 1974 747 1978
rect 791 1974 795 1978
rect 847 1974 851 1978
rect 863 1974 867 1978
rect 903 1974 907 1978
rect 959 1974 963 1978
rect 999 1974 1003 1978
rect 1015 1974 1019 1978
rect 1143 1974 1147 1978
rect 1271 1974 1275 1978
rect 1327 1974 1331 1978
rect 1367 1926 1371 1930
rect 1415 1926 1419 1930
rect 1495 1926 1499 1930
rect 1599 1926 1603 1930
rect 1695 1926 1699 1930
rect 1719 1926 1723 1930
rect 1775 1926 1779 1930
rect 1783 1926 1787 1930
rect 1831 1926 1835 1930
rect 1863 1926 1867 1930
rect 1887 1926 1891 1930
rect 1943 1926 1947 1930
rect 1999 1926 2003 1930
rect 2023 1926 2027 1930
rect 2055 1926 2059 1930
rect 2103 1926 2107 1930
rect 2119 1926 2123 1930
rect 2583 1926 2587 1930
rect 111 1918 115 1922
rect 159 1918 163 1922
rect 231 1918 235 1922
rect 327 1918 331 1922
rect 351 1918 355 1922
rect 407 1918 411 1922
rect 431 1918 435 1922
rect 463 1918 467 1922
rect 519 1918 523 1922
rect 543 1918 547 1922
rect 583 1918 587 1922
rect 655 1918 659 1922
rect 663 1918 667 1922
rect 759 1918 763 1922
rect 767 1918 771 1922
rect 879 1918 883 1922
rect 983 1918 987 1922
rect 1015 1918 1019 1922
rect 1087 1918 1091 1922
rect 1159 1918 1163 1922
rect 1199 1918 1203 1922
rect 1287 1918 1291 1922
rect 1327 1918 1331 1922
rect 1367 1866 1371 1870
rect 1399 1866 1403 1870
rect 1463 1866 1467 1870
rect 1559 1866 1563 1870
rect 1655 1866 1659 1870
rect 1703 1866 1707 1870
rect 1743 1866 1747 1870
rect 1759 1866 1763 1870
rect 1815 1866 1819 1870
rect 1831 1866 1835 1870
rect 1871 1866 1875 1870
rect 1919 1866 1923 1870
rect 1927 1866 1931 1870
rect 1983 1866 1987 1870
rect 2007 1866 2011 1870
rect 2039 1866 2043 1870
rect 2095 1866 2099 1870
rect 2103 1866 2107 1870
rect 2183 1866 2187 1870
rect 2583 1866 2587 1870
rect 111 1854 115 1858
rect 143 1854 147 1858
rect 199 1854 203 1858
rect 215 1854 219 1858
rect 263 1854 267 1858
rect 311 1854 315 1858
rect 351 1854 355 1858
rect 415 1854 419 1858
rect 439 1854 443 1858
rect 527 1854 531 1858
rect 535 1854 539 1858
rect 623 1854 627 1858
rect 639 1854 643 1858
rect 711 1854 715 1858
rect 751 1854 755 1858
rect 791 1854 795 1858
rect 863 1854 867 1858
rect 871 1854 875 1858
rect 951 1854 955 1858
rect 967 1854 971 1858
rect 1039 1854 1043 1858
rect 1071 1854 1075 1858
rect 1183 1854 1187 1858
rect 1271 1854 1275 1858
rect 1327 1854 1331 1858
rect 1367 1810 1371 1814
rect 1415 1810 1419 1814
rect 1479 1810 1483 1814
rect 1511 1810 1515 1814
rect 1575 1810 1579 1814
rect 1623 1810 1627 1814
rect 1671 1810 1675 1814
rect 1735 1810 1739 1814
rect 1759 1810 1763 1814
rect 1839 1810 1843 1814
rect 1847 1810 1851 1814
rect 1935 1810 1939 1814
rect 1951 1810 1955 1814
rect 2023 1810 2027 1814
rect 2063 1810 2067 1814
rect 2111 1810 2115 1814
rect 2183 1810 2187 1814
rect 2199 1810 2203 1814
rect 2303 1810 2307 1814
rect 2431 1810 2435 1814
rect 2543 1810 2547 1814
rect 2583 1810 2587 1814
rect 111 1794 115 1798
rect 159 1794 163 1798
rect 215 1794 219 1798
rect 231 1794 235 1798
rect 279 1794 283 1798
rect 295 1794 299 1798
rect 367 1794 371 1798
rect 447 1794 451 1798
rect 455 1794 459 1798
rect 535 1794 539 1798
rect 551 1794 555 1798
rect 623 1794 627 1798
rect 639 1794 643 1798
rect 711 1794 715 1798
rect 727 1794 731 1798
rect 791 1794 795 1798
rect 807 1794 811 1798
rect 871 1794 875 1798
rect 887 1794 891 1798
rect 951 1794 955 1798
rect 967 1794 971 1798
rect 1031 1794 1035 1798
rect 1055 1794 1059 1798
rect 1119 1794 1123 1798
rect 1327 1794 1331 1798
rect 1367 1754 1371 1758
rect 1399 1754 1403 1758
rect 1439 1754 1443 1758
rect 1495 1754 1499 1758
rect 1519 1754 1523 1758
rect 1607 1754 1611 1758
rect 1615 1754 1619 1758
rect 1719 1754 1723 1758
rect 1823 1754 1827 1758
rect 1927 1754 1931 1758
rect 1935 1754 1939 1758
rect 2023 1754 2027 1758
rect 2047 1754 2051 1758
rect 2119 1754 2123 1758
rect 2167 1754 2171 1758
rect 2207 1754 2211 1758
rect 2287 1754 2291 1758
rect 2375 1754 2379 1758
rect 2415 1754 2419 1758
rect 2463 1754 2467 1758
rect 2527 1754 2531 1758
rect 2583 1754 2587 1758
rect 111 1734 115 1738
rect 215 1734 219 1738
rect 279 1734 283 1738
rect 351 1734 355 1738
rect 407 1734 411 1738
rect 431 1734 435 1738
rect 471 1734 475 1738
rect 519 1734 523 1738
rect 551 1734 555 1738
rect 607 1734 611 1738
rect 639 1734 643 1738
rect 695 1734 699 1738
rect 727 1734 731 1738
rect 775 1734 779 1738
rect 823 1734 827 1738
rect 855 1734 859 1738
rect 919 1734 923 1738
rect 935 1734 939 1738
rect 1015 1734 1019 1738
rect 1103 1734 1107 1738
rect 1111 1734 1115 1738
rect 1207 1734 1211 1738
rect 1327 1734 1331 1738
rect 1367 1686 1371 1690
rect 1455 1686 1459 1690
rect 1535 1686 1539 1690
rect 1559 1686 1563 1690
rect 1631 1686 1635 1690
rect 1711 1686 1715 1690
rect 1735 1686 1739 1690
rect 1799 1686 1803 1690
rect 1839 1686 1843 1690
rect 1887 1686 1891 1690
rect 1943 1686 1947 1690
rect 1975 1686 1979 1690
rect 2039 1686 2043 1690
rect 2063 1686 2067 1690
rect 2135 1686 2139 1690
rect 2143 1686 2147 1690
rect 2215 1686 2219 1690
rect 2223 1686 2227 1690
rect 2287 1686 2291 1690
rect 2303 1686 2307 1690
rect 2351 1686 2355 1690
rect 2391 1686 2395 1690
rect 2423 1686 2427 1690
rect 2479 1686 2483 1690
rect 2487 1686 2491 1690
rect 2543 1686 2547 1690
rect 2583 1686 2587 1690
rect 111 1674 115 1678
rect 367 1674 371 1678
rect 399 1674 403 1678
rect 423 1674 427 1678
rect 455 1674 459 1678
rect 487 1674 491 1678
rect 511 1674 515 1678
rect 567 1674 571 1678
rect 575 1674 579 1678
rect 647 1674 651 1678
rect 655 1674 659 1678
rect 727 1674 731 1678
rect 743 1674 747 1678
rect 807 1674 811 1678
rect 839 1674 843 1678
rect 887 1674 891 1678
rect 935 1674 939 1678
rect 967 1674 971 1678
rect 1031 1674 1035 1678
rect 1047 1674 1051 1678
rect 1127 1674 1131 1678
rect 1135 1674 1139 1678
rect 1223 1674 1227 1678
rect 1287 1674 1291 1678
rect 1327 1674 1331 1678
rect 1367 1618 1371 1622
rect 1543 1618 1547 1622
rect 1575 1618 1579 1622
rect 1615 1618 1619 1622
rect 1631 1618 1635 1622
rect 1687 1618 1691 1622
rect 1695 1618 1699 1622
rect 1751 1618 1755 1622
rect 1783 1618 1787 1622
rect 1831 1618 1835 1622
rect 1871 1618 1875 1622
rect 1919 1618 1923 1622
rect 1959 1618 1963 1622
rect 2007 1618 2011 1622
rect 2047 1618 2051 1622
rect 2103 1618 2107 1622
rect 2127 1618 2131 1622
rect 2199 1618 2203 1622
rect 2207 1618 2211 1622
rect 2271 1618 2275 1622
rect 2319 1618 2323 1622
rect 2335 1618 2339 1622
rect 2407 1618 2411 1622
rect 2431 1618 2435 1622
rect 2471 1618 2475 1622
rect 2527 1618 2531 1622
rect 2583 1618 2587 1622
rect 111 1602 115 1606
rect 287 1602 291 1606
rect 367 1602 371 1606
rect 383 1602 387 1606
rect 439 1602 443 1606
rect 455 1602 459 1606
rect 495 1602 499 1606
rect 551 1602 555 1606
rect 559 1602 563 1606
rect 631 1602 635 1606
rect 647 1602 651 1606
rect 711 1602 715 1606
rect 735 1602 739 1606
rect 791 1602 795 1606
rect 823 1602 827 1606
rect 871 1602 875 1606
rect 903 1602 907 1606
rect 951 1602 955 1606
rect 983 1602 987 1606
rect 1031 1602 1035 1606
rect 1063 1602 1067 1606
rect 1119 1602 1123 1606
rect 1151 1602 1155 1606
rect 1207 1602 1211 1606
rect 1271 1602 1275 1606
rect 1327 1602 1331 1606
rect 1367 1558 1371 1562
rect 1591 1558 1595 1562
rect 1647 1558 1651 1562
rect 1679 1558 1683 1562
rect 1703 1558 1707 1562
rect 1735 1558 1739 1562
rect 1767 1558 1771 1562
rect 1791 1558 1795 1562
rect 1847 1558 1851 1562
rect 1855 1558 1859 1562
rect 1927 1558 1931 1562
rect 1935 1558 1939 1562
rect 2007 1558 2011 1562
rect 2023 1558 2027 1562
rect 2087 1558 2091 1562
rect 2119 1558 2123 1562
rect 2167 1558 2171 1562
rect 2223 1558 2227 1562
rect 2247 1558 2251 1562
rect 2327 1558 2331 1562
rect 2335 1558 2339 1562
rect 2407 1558 2411 1562
rect 2447 1558 2451 1562
rect 2487 1558 2491 1562
rect 2543 1558 2547 1562
rect 2583 1558 2587 1562
rect 111 1546 115 1550
rect 279 1546 283 1550
rect 303 1546 307 1550
rect 335 1546 339 1550
rect 383 1546 387 1550
rect 399 1546 403 1550
rect 471 1546 475 1550
rect 543 1546 547 1550
rect 567 1546 571 1550
rect 615 1546 619 1550
rect 663 1546 667 1550
rect 687 1546 691 1550
rect 751 1546 755 1550
rect 759 1546 763 1550
rect 831 1546 835 1550
rect 839 1546 843 1550
rect 903 1546 907 1550
rect 919 1546 923 1550
rect 975 1546 979 1550
rect 999 1546 1003 1550
rect 1055 1546 1059 1550
rect 1079 1546 1083 1550
rect 1167 1546 1171 1550
rect 1327 1546 1331 1550
rect 1367 1494 1371 1498
rect 1519 1494 1523 1498
rect 1575 1494 1579 1498
rect 1647 1494 1651 1498
rect 1663 1494 1667 1498
rect 1719 1494 1723 1498
rect 1727 1494 1731 1498
rect 1775 1494 1779 1498
rect 1807 1494 1811 1498
rect 1839 1494 1843 1498
rect 1895 1494 1899 1498
rect 1911 1494 1915 1498
rect 1983 1494 1987 1498
rect 1991 1494 1995 1498
rect 2071 1494 2075 1498
rect 2151 1494 2155 1498
rect 2231 1494 2235 1498
rect 2311 1494 2315 1498
rect 2391 1494 2395 1498
rect 2471 1494 2475 1498
rect 2527 1494 2531 1498
rect 2583 1494 2587 1498
rect 111 1486 115 1490
rect 199 1486 203 1490
rect 263 1486 267 1490
rect 287 1486 291 1490
rect 319 1486 323 1490
rect 383 1486 387 1490
rect 455 1486 459 1490
rect 487 1486 491 1490
rect 527 1486 531 1490
rect 583 1486 587 1490
rect 599 1486 603 1490
rect 671 1486 675 1490
rect 679 1486 683 1490
rect 743 1486 747 1490
rect 775 1486 779 1490
rect 815 1486 819 1490
rect 863 1486 867 1490
rect 887 1486 891 1490
rect 951 1486 955 1490
rect 959 1486 963 1490
rect 1039 1486 1043 1490
rect 1135 1486 1139 1490
rect 1327 1486 1331 1490
rect 111 1426 115 1430
rect 159 1426 163 1430
rect 215 1426 219 1430
rect 247 1426 251 1430
rect 303 1426 307 1430
rect 343 1426 347 1430
rect 399 1426 403 1430
rect 447 1426 451 1430
rect 503 1426 507 1430
rect 551 1426 555 1430
rect 599 1426 603 1430
rect 663 1426 667 1430
rect 695 1426 699 1430
rect 767 1426 771 1430
rect 791 1426 795 1430
rect 879 1426 883 1430
rect 967 1426 971 1430
rect 991 1426 995 1430
rect 1055 1426 1059 1430
rect 1103 1426 1107 1430
rect 1151 1426 1155 1430
rect 1215 1426 1219 1430
rect 1327 1426 1331 1430
rect 1367 1430 1371 1434
rect 1415 1430 1419 1434
rect 1471 1430 1475 1434
rect 1535 1430 1539 1434
rect 1591 1430 1595 1434
rect 1623 1430 1627 1434
rect 1663 1430 1667 1434
rect 1719 1430 1723 1434
rect 1743 1430 1747 1434
rect 1823 1430 1827 1434
rect 1911 1430 1915 1434
rect 1927 1430 1931 1434
rect 1999 1430 2003 1434
rect 2023 1430 2027 1434
rect 2087 1430 2091 1434
rect 2119 1430 2123 1434
rect 2167 1430 2171 1434
rect 2215 1430 2219 1434
rect 2247 1430 2251 1434
rect 2303 1430 2307 1434
rect 2327 1430 2331 1434
rect 2391 1430 2395 1434
rect 2407 1430 2411 1434
rect 2479 1430 2483 1434
rect 2487 1430 2491 1434
rect 2543 1430 2547 1434
rect 2583 1430 2587 1434
rect 111 1370 115 1374
rect 143 1370 147 1374
rect 207 1370 211 1374
rect 231 1370 235 1374
rect 295 1370 299 1374
rect 327 1370 331 1374
rect 399 1370 403 1374
rect 431 1370 435 1374
rect 511 1370 515 1374
rect 535 1370 539 1374
rect 623 1370 627 1374
rect 647 1370 651 1374
rect 735 1370 739 1374
rect 751 1370 755 1374
rect 847 1370 851 1374
rect 863 1370 867 1374
rect 959 1370 963 1374
rect 975 1370 979 1374
rect 1071 1370 1075 1374
rect 1087 1370 1091 1374
rect 1183 1370 1187 1374
rect 1199 1370 1203 1374
rect 1271 1370 1275 1374
rect 1327 1370 1331 1374
rect 1367 1366 1371 1370
rect 1399 1366 1403 1370
rect 1455 1366 1459 1370
rect 1519 1366 1523 1370
rect 1543 1366 1547 1370
rect 1607 1366 1611 1370
rect 1631 1366 1635 1370
rect 1703 1366 1707 1370
rect 1719 1366 1723 1370
rect 1807 1366 1811 1370
rect 1887 1366 1891 1370
rect 1911 1366 1915 1370
rect 1967 1366 1971 1370
rect 2007 1366 2011 1370
rect 2047 1366 2051 1370
rect 2103 1366 2107 1370
rect 2127 1366 2131 1370
rect 2199 1366 2203 1370
rect 2207 1366 2211 1370
rect 2287 1366 2291 1370
rect 2375 1366 2379 1370
rect 2463 1366 2467 1370
rect 2527 1366 2531 1370
rect 2583 1366 2587 1370
rect 111 1314 115 1318
rect 159 1314 163 1318
rect 223 1314 227 1318
rect 231 1314 235 1318
rect 311 1314 315 1318
rect 327 1314 331 1318
rect 415 1314 419 1318
rect 431 1314 435 1318
rect 527 1314 531 1318
rect 535 1314 539 1318
rect 631 1314 635 1318
rect 639 1314 643 1318
rect 727 1314 731 1318
rect 751 1314 755 1318
rect 823 1314 827 1318
rect 863 1314 867 1318
rect 911 1314 915 1318
rect 975 1314 979 1318
rect 991 1314 995 1318
rect 1071 1314 1075 1318
rect 1087 1314 1091 1318
rect 1151 1314 1155 1318
rect 1199 1314 1203 1318
rect 1231 1314 1235 1318
rect 1287 1314 1291 1318
rect 1327 1314 1331 1318
rect 1367 1306 1371 1310
rect 1415 1306 1419 1310
rect 1471 1306 1475 1310
rect 1559 1306 1563 1310
rect 1647 1306 1651 1310
rect 1671 1306 1675 1310
rect 1735 1306 1739 1310
rect 1767 1306 1771 1310
rect 1823 1306 1827 1310
rect 1863 1306 1867 1310
rect 1903 1306 1907 1310
rect 1959 1306 1963 1310
rect 1983 1306 1987 1310
rect 2047 1306 2051 1310
rect 2063 1306 2067 1310
rect 2135 1306 2139 1310
rect 2143 1306 2147 1310
rect 2223 1306 2227 1310
rect 2231 1306 2235 1310
rect 2583 1306 2587 1310
rect 111 1246 115 1250
rect 143 1246 147 1250
rect 199 1246 203 1250
rect 215 1246 219 1250
rect 279 1246 283 1250
rect 311 1246 315 1250
rect 359 1246 363 1250
rect 415 1246 419 1250
rect 439 1246 443 1250
rect 519 1246 523 1250
rect 599 1246 603 1250
rect 615 1246 619 1250
rect 671 1246 675 1250
rect 711 1246 715 1250
rect 743 1246 747 1250
rect 807 1246 811 1250
rect 815 1246 819 1250
rect 895 1246 899 1250
rect 975 1246 979 1250
rect 1055 1246 1059 1250
rect 1135 1246 1139 1250
rect 1215 1246 1219 1250
rect 1271 1246 1275 1250
rect 1327 1246 1331 1250
rect 1367 1250 1371 1254
rect 1495 1250 1499 1254
rect 1559 1250 1563 1254
rect 1623 1250 1627 1254
rect 1655 1250 1659 1254
rect 1687 1250 1691 1254
rect 1751 1250 1755 1254
rect 1759 1250 1763 1254
rect 1823 1250 1827 1254
rect 1847 1250 1851 1254
rect 1887 1250 1891 1254
rect 1943 1250 1947 1254
rect 1951 1250 1955 1254
rect 2015 1250 2019 1254
rect 2031 1250 2035 1254
rect 2079 1250 2083 1254
rect 2119 1250 2123 1254
rect 2151 1250 2155 1254
rect 2215 1250 2219 1254
rect 2223 1250 2227 1254
rect 2295 1250 2299 1254
rect 2583 1250 2587 1254
rect 111 1186 115 1190
rect 159 1186 163 1190
rect 215 1186 219 1190
rect 239 1186 243 1190
rect 295 1186 299 1190
rect 327 1186 331 1190
rect 375 1186 379 1190
rect 423 1186 427 1190
rect 455 1186 459 1190
rect 511 1186 515 1190
rect 535 1186 539 1190
rect 599 1186 603 1190
rect 615 1186 619 1190
rect 687 1186 691 1190
rect 759 1186 763 1190
rect 767 1186 771 1190
rect 831 1186 835 1190
rect 839 1186 843 1190
rect 911 1186 915 1190
rect 983 1186 987 1190
rect 1063 1186 1067 1190
rect 1327 1186 1331 1190
rect 1367 1186 1371 1190
rect 1415 1186 1419 1190
rect 1503 1186 1507 1190
rect 1511 1186 1515 1190
rect 1575 1186 1579 1190
rect 1599 1186 1603 1190
rect 1639 1186 1643 1190
rect 1703 1186 1707 1190
rect 1775 1186 1779 1190
rect 1807 1186 1811 1190
rect 1839 1186 1843 1190
rect 1903 1186 1907 1190
rect 1911 1186 1915 1190
rect 1967 1186 1971 1190
rect 2015 1186 2019 1190
rect 2031 1186 2035 1190
rect 2095 1186 2099 1190
rect 2111 1186 2115 1190
rect 2167 1186 2171 1190
rect 2207 1186 2211 1190
rect 2239 1186 2243 1190
rect 2303 1186 2307 1190
rect 2311 1186 2315 1190
rect 2399 1186 2403 1190
rect 2583 1186 2587 1190
rect 111 1122 115 1126
rect 143 1122 147 1126
rect 223 1122 227 1126
rect 311 1122 315 1126
rect 319 1122 323 1126
rect 407 1122 411 1126
rect 423 1122 427 1126
rect 495 1122 499 1126
rect 527 1122 531 1126
rect 583 1122 587 1126
rect 631 1122 635 1126
rect 671 1122 675 1126
rect 727 1122 731 1126
rect 751 1122 755 1126
rect 823 1122 827 1126
rect 895 1122 899 1126
rect 911 1122 915 1126
rect 967 1122 971 1126
rect 991 1122 995 1126
rect 1047 1122 1051 1126
rect 1079 1122 1083 1126
rect 1167 1122 1171 1126
rect 1327 1122 1331 1126
rect 1367 1126 1371 1130
rect 1399 1126 1403 1130
rect 1479 1126 1483 1130
rect 1487 1126 1491 1130
rect 1583 1126 1587 1130
rect 1687 1126 1691 1130
rect 1791 1126 1795 1130
rect 1887 1126 1891 1130
rect 1895 1126 1899 1130
rect 1975 1126 1979 1130
rect 1999 1126 2003 1130
rect 2063 1126 2067 1130
rect 2095 1126 2099 1130
rect 2143 1126 2147 1130
rect 2191 1126 2195 1130
rect 2215 1126 2219 1130
rect 2279 1126 2283 1130
rect 2287 1126 2291 1130
rect 2343 1126 2347 1130
rect 2383 1126 2387 1130
rect 2407 1126 2411 1130
rect 2471 1126 2475 1130
rect 2527 1126 2531 1130
rect 2583 1126 2587 1130
rect 111 1062 115 1066
rect 239 1062 243 1066
rect 311 1062 315 1066
rect 335 1062 339 1066
rect 367 1062 371 1066
rect 439 1062 443 1066
rect 519 1062 523 1066
rect 543 1062 547 1066
rect 607 1062 611 1066
rect 647 1062 651 1066
rect 703 1062 707 1066
rect 743 1062 747 1066
rect 799 1062 803 1066
rect 839 1062 843 1066
rect 887 1062 891 1066
rect 927 1062 931 1066
rect 975 1062 979 1066
rect 1007 1062 1011 1066
rect 1055 1062 1059 1066
rect 1095 1062 1099 1066
rect 1135 1062 1139 1066
rect 1183 1062 1187 1066
rect 1223 1062 1227 1066
rect 1287 1062 1291 1066
rect 1327 1062 1331 1066
rect 1367 1066 1371 1070
rect 1415 1066 1419 1070
rect 1471 1066 1475 1070
rect 1495 1066 1499 1070
rect 1535 1066 1539 1070
rect 1599 1066 1603 1070
rect 1623 1066 1627 1070
rect 1703 1066 1707 1070
rect 1727 1066 1731 1070
rect 1807 1066 1811 1070
rect 1839 1066 1843 1070
rect 1903 1066 1907 1070
rect 1951 1066 1955 1070
rect 1991 1066 1995 1070
rect 2063 1066 2067 1070
rect 2079 1066 2083 1070
rect 2159 1066 2163 1070
rect 2167 1066 2171 1070
rect 2231 1066 2235 1070
rect 2271 1066 2275 1070
rect 2295 1066 2299 1070
rect 2359 1066 2363 1070
rect 2367 1066 2371 1070
rect 2423 1066 2427 1070
rect 2463 1066 2467 1070
rect 2487 1066 2491 1070
rect 2543 1066 2547 1070
rect 2583 1066 2587 1070
rect 111 1002 115 1006
rect 295 1002 299 1006
rect 351 1002 355 1006
rect 415 1002 419 1006
rect 423 1002 427 1006
rect 471 1002 475 1006
rect 503 1002 507 1006
rect 527 1002 531 1006
rect 591 1002 595 1006
rect 655 1002 659 1006
rect 687 1002 691 1006
rect 719 1002 723 1006
rect 783 1002 787 1006
rect 847 1002 851 1006
rect 871 1002 875 1006
rect 911 1002 915 1006
rect 959 1002 963 1006
rect 975 1002 979 1006
rect 1039 1002 1043 1006
rect 1103 1002 1107 1006
rect 1119 1002 1123 1006
rect 1159 1002 1163 1006
rect 1207 1002 1211 1006
rect 1215 1002 1219 1006
rect 1271 1002 1275 1006
rect 1327 1002 1331 1006
rect 1367 994 1371 998
rect 1399 994 1403 998
rect 1455 994 1459 998
rect 1511 994 1515 998
rect 1519 994 1523 998
rect 1567 994 1571 998
rect 1607 994 1611 998
rect 1639 994 1643 998
rect 1711 994 1715 998
rect 1719 994 1723 998
rect 1807 994 1811 998
rect 1823 994 1827 998
rect 1903 994 1907 998
rect 1935 994 1939 998
rect 2015 994 2019 998
rect 2047 994 2051 998
rect 2143 994 2147 998
rect 2151 994 2155 998
rect 2255 994 2259 998
rect 2271 994 2275 998
rect 2351 994 2355 998
rect 2407 994 2411 998
rect 2447 994 2451 998
rect 2527 994 2531 998
rect 2583 994 2587 998
rect 111 942 115 946
rect 423 942 427 946
rect 431 942 435 946
rect 479 942 483 946
rect 487 942 491 946
rect 535 942 539 946
rect 543 942 547 946
rect 591 942 595 946
rect 607 942 611 946
rect 647 942 651 946
rect 671 942 675 946
rect 703 942 707 946
rect 735 942 739 946
rect 759 942 763 946
rect 799 942 803 946
rect 815 942 819 946
rect 863 942 867 946
rect 927 942 931 946
rect 991 942 995 946
rect 1055 942 1059 946
rect 1119 942 1123 946
rect 1175 942 1179 946
rect 1231 942 1235 946
rect 1287 942 1291 946
rect 1327 942 1331 946
rect 1367 930 1371 934
rect 1415 930 1419 934
rect 1471 930 1475 934
rect 1527 930 1531 934
rect 1583 930 1587 934
rect 1615 930 1619 934
rect 1655 930 1659 934
rect 1711 930 1715 934
rect 1735 930 1739 934
rect 1823 930 1827 934
rect 1919 930 1923 934
rect 1943 930 1947 934
rect 2031 930 2035 934
rect 2063 930 2067 934
rect 2159 930 2163 934
rect 2183 930 2187 934
rect 2287 930 2291 934
rect 2311 930 2315 934
rect 2423 930 2427 934
rect 2439 930 2443 934
rect 2543 930 2547 934
rect 2583 930 2587 934
rect 111 886 115 890
rect 279 886 283 890
rect 335 886 339 890
rect 391 886 395 890
rect 407 886 411 890
rect 455 886 459 890
rect 463 886 467 890
rect 519 886 523 890
rect 575 886 579 890
rect 583 886 587 890
rect 631 886 635 890
rect 647 886 651 890
rect 687 886 691 890
rect 711 886 715 890
rect 743 886 747 890
rect 775 886 779 890
rect 799 886 803 890
rect 847 886 851 890
rect 919 886 923 890
rect 1327 886 1331 890
rect 1367 874 1371 878
rect 1399 874 1403 878
rect 1455 874 1459 878
rect 1471 874 1475 878
rect 1511 874 1515 878
rect 1551 874 1555 878
rect 1599 874 1603 878
rect 1639 874 1643 878
rect 1695 874 1699 878
rect 1727 874 1731 878
rect 1807 874 1811 878
rect 1815 874 1819 878
rect 1903 874 1907 878
rect 1927 874 1931 878
rect 1991 874 1995 878
rect 2047 874 2051 878
rect 2071 874 2075 878
rect 2143 874 2147 878
rect 2167 874 2171 878
rect 2215 874 2219 878
rect 2279 874 2283 878
rect 2295 874 2299 878
rect 2343 874 2347 878
rect 2407 874 2411 878
rect 2423 874 2427 878
rect 2471 874 2475 878
rect 2527 874 2531 878
rect 2583 874 2587 878
rect 111 822 115 826
rect 167 822 171 826
rect 231 822 235 826
rect 295 822 299 826
rect 311 822 315 826
rect 351 822 355 826
rect 399 822 403 826
rect 407 822 411 826
rect 471 822 475 826
rect 487 822 491 826
rect 535 822 539 826
rect 583 822 587 826
rect 599 822 603 826
rect 663 822 667 826
rect 671 822 675 826
rect 727 822 731 826
rect 759 822 763 826
rect 791 822 795 826
rect 839 822 843 826
rect 863 822 867 826
rect 919 822 923 826
rect 935 822 939 826
rect 1007 822 1011 826
rect 1095 822 1099 826
rect 1327 822 1331 826
rect 1367 810 1371 814
rect 1487 810 1491 814
rect 1567 810 1571 814
rect 1631 810 1635 814
rect 1655 810 1659 814
rect 1687 810 1691 814
rect 1743 810 1747 814
rect 1751 810 1755 814
rect 1823 810 1827 814
rect 1831 810 1835 814
rect 1903 810 1907 814
rect 1919 810 1923 814
rect 1991 810 1995 814
rect 2007 810 2011 814
rect 2071 810 2075 814
rect 2087 810 2091 814
rect 2159 810 2163 814
rect 2231 810 2235 814
rect 2247 810 2251 814
rect 2295 810 2299 814
rect 2335 810 2339 814
rect 2359 810 2363 814
rect 2423 810 2427 814
rect 2487 810 2491 814
rect 2543 810 2547 814
rect 2583 810 2587 814
rect 111 758 115 762
rect 143 758 147 762
rect 151 758 155 762
rect 199 758 203 762
rect 215 758 219 762
rect 279 758 283 762
rect 295 758 299 762
rect 383 758 387 762
rect 471 758 475 762
rect 487 758 491 762
rect 567 758 571 762
rect 599 758 603 762
rect 655 758 659 762
rect 703 758 707 762
rect 743 758 747 762
rect 807 758 811 762
rect 823 758 827 762
rect 903 758 907 762
rect 991 758 995 762
rect 1079 758 1083 762
rect 1175 758 1179 762
rect 1327 758 1331 762
rect 1367 750 1371 754
rect 1567 750 1571 754
rect 1615 750 1619 754
rect 1623 750 1627 754
rect 1671 750 1675 754
rect 1687 750 1691 754
rect 1735 750 1739 754
rect 1759 750 1763 754
rect 1807 750 1811 754
rect 1839 750 1843 754
rect 1887 750 1891 754
rect 1919 750 1923 754
rect 1975 750 1979 754
rect 1999 750 2003 754
rect 2055 750 2059 754
rect 2079 750 2083 754
rect 2143 750 2147 754
rect 2159 750 2163 754
rect 2231 750 2235 754
rect 2247 750 2251 754
rect 2319 750 2323 754
rect 2335 750 2339 754
rect 2407 750 2411 754
rect 2583 750 2587 754
rect 111 698 115 702
rect 159 698 163 702
rect 215 698 219 702
rect 279 698 283 702
rect 295 698 299 702
rect 359 698 363 702
rect 399 698 403 702
rect 447 698 451 702
rect 503 698 507 702
rect 535 698 539 702
rect 615 698 619 702
rect 623 698 627 702
rect 711 698 715 702
rect 719 698 723 702
rect 791 698 795 702
rect 823 698 827 702
rect 871 698 875 702
rect 919 698 923 702
rect 951 698 955 702
rect 1007 698 1011 702
rect 1039 698 1043 702
rect 1095 698 1099 702
rect 1191 698 1195 702
rect 1327 698 1331 702
rect 1367 690 1371 694
rect 1415 690 1419 694
rect 1511 690 1515 694
rect 1583 690 1587 694
rect 1615 690 1619 694
rect 1639 690 1643 694
rect 1703 690 1707 694
rect 1719 690 1723 694
rect 1775 690 1779 694
rect 1823 690 1827 694
rect 1855 690 1859 694
rect 1927 690 1931 694
rect 1935 690 1939 694
rect 2015 690 2019 694
rect 2023 690 2027 694
rect 2095 690 2099 694
rect 2119 690 2123 694
rect 2175 690 2179 694
rect 2207 690 2211 694
rect 2263 690 2267 694
rect 2295 690 2299 694
rect 2351 690 2355 694
rect 2391 690 2395 694
rect 2583 690 2587 694
rect 111 634 115 638
rect 143 634 147 638
rect 199 634 203 638
rect 255 634 259 638
rect 263 634 267 638
rect 311 634 315 638
rect 343 634 347 638
rect 391 634 395 638
rect 431 634 435 638
rect 479 634 483 638
rect 519 634 523 638
rect 575 634 579 638
rect 607 634 611 638
rect 679 634 683 638
rect 695 634 699 638
rect 775 634 779 638
rect 783 634 787 638
rect 855 634 859 638
rect 887 634 891 638
rect 935 634 939 638
rect 991 634 995 638
rect 1023 634 1027 638
rect 1087 634 1091 638
rect 1191 634 1195 638
rect 1271 634 1275 638
rect 1327 634 1331 638
rect 1367 634 1371 638
rect 1399 634 1403 638
rect 1495 634 1499 638
rect 1511 634 1515 638
rect 1599 634 1603 638
rect 1647 634 1651 638
rect 1703 634 1707 638
rect 1783 634 1787 638
rect 1807 634 1811 638
rect 1911 634 1915 638
rect 2007 634 2011 638
rect 2039 634 2043 638
rect 2103 634 2107 638
rect 2159 634 2163 638
rect 2191 634 2195 638
rect 2279 634 2283 638
rect 2375 634 2379 638
rect 2407 634 2411 638
rect 2583 634 2587 638
rect 111 574 115 578
rect 159 574 163 578
rect 199 574 203 578
rect 215 574 219 578
rect 263 574 267 578
rect 271 574 275 578
rect 327 574 331 578
rect 335 574 339 578
rect 407 574 411 578
rect 415 574 419 578
rect 495 574 499 578
rect 511 574 515 578
rect 591 574 595 578
rect 615 574 619 578
rect 695 574 699 578
rect 719 574 723 578
rect 799 574 803 578
rect 831 574 835 578
rect 903 574 907 578
rect 943 574 947 578
rect 1007 574 1011 578
rect 1063 574 1067 578
rect 1103 574 1107 578
rect 1183 574 1187 578
rect 1207 574 1211 578
rect 1287 574 1291 578
rect 1327 574 1331 578
rect 1367 570 1371 574
rect 1415 570 1419 574
rect 1471 570 1475 574
rect 1527 570 1531 574
rect 1551 570 1555 574
rect 1647 570 1651 574
rect 1663 570 1667 574
rect 1751 570 1755 574
rect 1799 570 1803 574
rect 1855 570 1859 574
rect 1927 570 1931 574
rect 1959 570 1963 574
rect 2055 570 2059 574
rect 2151 570 2155 574
rect 2175 570 2179 574
rect 2239 570 2243 574
rect 2295 570 2299 574
rect 2319 570 2323 574
rect 2399 570 2403 574
rect 2423 570 2427 574
rect 2479 570 2483 574
rect 2543 570 2547 574
rect 2583 570 2587 574
rect 111 510 115 514
rect 183 510 187 514
rect 247 510 251 514
rect 303 510 307 514
rect 319 510 323 514
rect 359 510 363 514
rect 399 510 403 514
rect 423 510 427 514
rect 495 510 499 514
rect 575 510 579 514
rect 599 510 603 514
rect 647 510 651 514
rect 703 510 707 514
rect 719 510 723 514
rect 791 510 795 514
rect 815 510 819 514
rect 863 510 867 514
rect 927 510 931 514
rect 935 510 939 514
rect 1007 510 1011 514
rect 1047 510 1051 514
rect 1087 510 1091 514
rect 1167 510 1171 514
rect 1271 510 1275 514
rect 1327 510 1331 514
rect 1367 514 1371 518
rect 1399 514 1403 518
rect 1455 514 1459 518
rect 1535 514 1539 518
rect 1599 514 1603 518
rect 1631 514 1635 518
rect 1671 514 1675 518
rect 1735 514 1739 518
rect 1751 514 1755 518
rect 1839 514 1843 518
rect 1927 514 1931 518
rect 1943 514 1947 518
rect 2015 514 2019 518
rect 2039 514 2043 518
rect 2095 514 2099 518
rect 2135 514 2139 518
rect 2175 514 2179 518
rect 2223 514 2227 518
rect 2255 514 2259 518
rect 2303 514 2307 518
rect 2327 514 2331 518
rect 2383 514 2387 518
rect 2399 514 2403 518
rect 2463 514 2467 518
rect 2471 514 2475 518
rect 2527 514 2531 518
rect 2583 514 2587 518
rect 111 450 115 454
rect 319 450 323 454
rect 375 450 379 454
rect 439 450 443 454
rect 455 450 459 454
rect 511 450 515 454
rect 575 450 579 454
rect 591 450 595 454
rect 647 450 651 454
rect 663 450 667 454
rect 727 450 731 454
rect 735 450 739 454
rect 799 450 803 454
rect 807 450 811 454
rect 871 450 875 454
rect 879 450 883 454
rect 943 450 947 454
rect 951 450 955 454
rect 1015 450 1019 454
rect 1023 450 1027 454
rect 1087 450 1091 454
rect 1103 450 1107 454
rect 1159 450 1163 454
rect 1239 450 1243 454
rect 1327 450 1331 454
rect 1367 450 1371 454
rect 1551 450 1555 454
rect 1615 450 1619 454
rect 1647 450 1651 454
rect 1687 450 1691 454
rect 1703 450 1707 454
rect 1759 450 1763 454
rect 1767 450 1771 454
rect 1815 450 1819 454
rect 1855 450 1859 454
rect 1871 450 1875 454
rect 1927 450 1931 454
rect 1943 450 1947 454
rect 1999 450 2003 454
rect 2031 450 2035 454
rect 2087 450 2091 454
rect 2111 450 2115 454
rect 2191 450 2195 454
rect 2271 450 2275 454
rect 2311 450 2315 454
rect 2343 450 2347 454
rect 2415 450 2419 454
rect 2439 450 2443 454
rect 2487 450 2491 454
rect 2543 450 2547 454
rect 2583 450 2587 454
rect 111 390 115 394
rect 415 390 419 394
rect 439 390 443 394
rect 471 390 475 394
rect 495 390 499 394
rect 535 390 539 394
rect 559 390 563 394
rect 607 390 611 394
rect 631 390 635 394
rect 687 390 691 394
rect 711 390 715 394
rect 767 390 771 394
rect 783 390 787 394
rect 847 390 851 394
rect 855 390 859 394
rect 927 390 931 394
rect 999 390 1003 394
rect 1007 390 1011 394
rect 1071 390 1075 394
rect 1087 390 1091 394
rect 1143 390 1147 394
rect 1175 390 1179 394
rect 1223 390 1227 394
rect 1263 390 1267 394
rect 1327 390 1331 394
rect 1367 394 1371 398
rect 1631 394 1635 398
rect 1655 394 1659 398
rect 1687 394 1691 398
rect 1711 394 1715 398
rect 1743 394 1747 398
rect 1767 394 1771 398
rect 1799 394 1803 398
rect 1823 394 1827 398
rect 1855 394 1859 398
rect 1879 394 1883 398
rect 1911 394 1915 398
rect 1951 394 1955 398
rect 1983 394 1987 398
rect 2039 394 2043 398
rect 2071 394 2075 398
rect 2151 394 2155 398
rect 2175 394 2179 398
rect 2279 394 2283 398
rect 2295 394 2299 398
rect 2415 394 2419 398
rect 2423 394 2427 398
rect 2527 394 2531 398
rect 2583 394 2587 398
rect 111 330 115 334
rect 431 330 435 334
rect 463 330 467 334
rect 487 330 491 334
rect 519 330 523 334
rect 551 330 555 334
rect 575 330 579 334
rect 623 330 627 334
rect 631 330 635 334
rect 695 330 699 334
rect 703 330 707 334
rect 767 330 771 334
rect 783 330 787 334
rect 847 330 851 334
rect 863 330 867 334
rect 927 330 931 334
rect 943 330 947 334
rect 1015 330 1019 334
rect 1023 330 1027 334
rect 1103 330 1107 334
rect 1111 330 1115 334
rect 1191 330 1195 334
rect 1215 330 1219 334
rect 1279 330 1283 334
rect 1327 330 1331 334
rect 1367 330 1371 334
rect 1631 330 1635 334
rect 1671 330 1675 334
rect 1687 330 1691 334
rect 1727 330 1731 334
rect 1743 330 1747 334
rect 1783 330 1787 334
rect 1807 330 1811 334
rect 1839 330 1843 334
rect 1887 330 1891 334
rect 1895 330 1899 334
rect 1967 330 1971 334
rect 2055 330 2059 334
rect 2143 330 2147 334
rect 2167 330 2171 334
rect 2231 330 2235 334
rect 2295 330 2299 334
rect 2311 330 2315 334
rect 2391 330 2395 334
rect 2431 330 2435 334
rect 2479 330 2483 334
rect 2543 330 2547 334
rect 2583 330 2587 334
rect 111 270 115 274
rect 287 270 291 274
rect 359 270 363 274
rect 439 270 443 274
rect 447 270 451 274
rect 503 270 507 274
rect 527 270 531 274
rect 559 270 563 274
rect 615 270 619 274
rect 623 270 627 274
rect 679 270 683 274
rect 719 270 723 274
rect 751 270 755 274
rect 823 270 827 274
rect 831 270 835 274
rect 911 270 915 274
rect 927 270 931 274
rect 999 270 1003 274
rect 1031 270 1035 274
rect 1095 270 1099 274
rect 1143 270 1147 274
rect 1199 270 1203 274
rect 1255 270 1259 274
rect 1327 270 1331 274
rect 1367 274 1371 278
rect 1535 274 1539 278
rect 1607 274 1611 278
rect 1615 274 1619 278
rect 1671 274 1675 278
rect 1687 274 1691 278
rect 1727 274 1731 278
rect 1775 274 1779 278
rect 1791 274 1795 278
rect 1863 274 1867 278
rect 1871 274 1875 278
rect 1951 274 1955 278
rect 2039 274 2043 278
rect 2119 274 2123 278
rect 2127 274 2131 278
rect 2199 274 2203 278
rect 2215 274 2219 278
rect 2271 274 2275 278
rect 2295 274 2299 278
rect 2335 274 2339 278
rect 2375 274 2379 278
rect 2407 274 2411 278
rect 2463 274 2467 278
rect 2471 274 2475 278
rect 2527 274 2531 278
rect 2583 274 2587 278
rect 111 214 115 218
rect 199 214 203 218
rect 271 214 275 218
rect 303 214 307 218
rect 359 214 363 218
rect 375 214 379 218
rect 455 214 459 218
rect 463 214 467 218
rect 543 214 547 218
rect 567 214 571 218
rect 639 214 643 218
rect 679 214 683 218
rect 735 214 739 218
rect 791 214 795 218
rect 839 214 843 218
rect 911 214 915 218
rect 943 214 947 218
rect 1031 214 1035 218
rect 1047 214 1051 218
rect 1151 214 1155 218
rect 1159 214 1163 218
rect 1271 214 1275 218
rect 1327 214 1331 218
rect 1367 218 1371 222
rect 1415 218 1419 222
rect 1479 218 1483 222
rect 1551 218 1555 222
rect 1559 218 1563 222
rect 1623 218 1627 222
rect 1655 218 1659 222
rect 1703 218 1707 222
rect 1751 218 1755 222
rect 1791 218 1795 222
rect 1855 218 1859 222
rect 1879 218 1883 222
rect 1959 218 1963 222
rect 1967 218 1971 222
rect 2055 218 2059 222
rect 2063 218 2067 222
rect 2135 218 2139 222
rect 2167 218 2171 222
rect 2215 218 2219 222
rect 2263 218 2267 222
rect 2287 218 2291 222
rect 2351 218 2355 222
rect 2359 218 2363 222
rect 2423 218 2427 222
rect 2463 218 2467 222
rect 2487 218 2491 222
rect 2543 218 2547 222
rect 2583 218 2587 222
rect 1367 146 1371 150
rect 1399 146 1403 150
rect 1455 146 1459 150
rect 1463 146 1467 150
rect 1511 146 1515 150
rect 1543 146 1547 150
rect 1567 146 1571 150
rect 1631 146 1635 150
rect 1639 146 1643 150
rect 1711 146 1715 150
rect 1735 146 1739 150
rect 1791 146 1795 150
rect 1839 146 1843 150
rect 1871 146 1875 150
rect 1943 146 1947 150
rect 2015 146 2019 150
rect 2047 146 2051 150
rect 2079 146 2083 150
rect 2143 146 2147 150
rect 2151 146 2155 150
rect 2207 146 2211 150
rect 2247 146 2251 150
rect 2271 146 2275 150
rect 2343 146 2347 150
rect 2415 146 2419 150
rect 2447 146 2451 150
rect 2527 146 2531 150
rect 2583 146 2587 150
rect 111 134 115 138
rect 143 134 147 138
rect 183 134 187 138
rect 199 134 203 138
rect 255 134 259 138
rect 311 134 315 138
rect 343 134 347 138
rect 367 134 371 138
rect 423 134 427 138
rect 447 134 451 138
rect 479 134 483 138
rect 535 134 539 138
rect 551 134 555 138
rect 591 134 595 138
rect 647 134 651 138
rect 663 134 667 138
rect 703 134 707 138
rect 759 134 763 138
rect 775 134 779 138
rect 823 134 827 138
rect 887 134 891 138
rect 895 134 899 138
rect 951 134 955 138
rect 1015 134 1019 138
rect 1079 134 1083 138
rect 1135 134 1139 138
rect 1151 134 1155 138
rect 1215 134 1219 138
rect 1255 134 1259 138
rect 1271 134 1275 138
rect 1327 134 1331 138
rect 1367 90 1371 94
rect 1415 90 1419 94
rect 1471 90 1475 94
rect 1527 90 1531 94
rect 1583 90 1587 94
rect 1647 90 1651 94
rect 1727 90 1731 94
rect 1807 90 1811 94
rect 1887 90 1891 94
rect 1959 90 1963 94
rect 2031 90 2035 94
rect 2095 90 2099 94
rect 2159 90 2163 94
rect 2223 90 2227 94
rect 2287 90 2291 94
rect 2359 90 2363 94
rect 2431 90 2435 94
rect 2583 90 2587 94
rect 111 78 115 82
rect 159 78 163 82
rect 215 78 219 82
rect 271 78 275 82
rect 327 78 331 82
rect 383 78 387 82
rect 439 78 443 82
rect 495 78 499 82
rect 551 78 555 82
rect 607 78 611 82
rect 663 78 667 82
rect 719 78 723 82
rect 775 78 779 82
rect 839 78 843 82
rect 903 78 907 82
rect 967 78 971 82
rect 1031 78 1035 82
rect 1095 78 1099 82
rect 1167 78 1171 82
rect 1231 78 1235 82
rect 1287 78 1291 82
rect 1327 78 1331 82
<< m4 >>
rect 84 2637 85 2643
rect 91 2642 1339 2643
rect 91 2638 111 2642
rect 115 2638 551 2642
rect 555 2638 607 2642
rect 611 2638 663 2642
rect 667 2638 719 2642
rect 723 2638 775 2642
rect 779 2638 1327 2642
rect 1331 2638 1339 2642
rect 91 2637 1339 2638
rect 1345 2639 1346 2643
rect 1345 2638 2618 2639
rect 1345 2637 1367 2638
rect 1338 2634 1367 2637
rect 1371 2634 1551 2638
rect 1555 2634 1607 2638
rect 1611 2634 1663 2638
rect 1667 2634 1719 2638
rect 1723 2634 1775 2638
rect 1779 2634 1831 2638
rect 1835 2634 1887 2638
rect 1891 2634 1943 2638
rect 1947 2634 1999 2638
rect 2003 2634 2055 2638
rect 2059 2634 2111 2638
rect 2115 2634 2167 2638
rect 2171 2634 2583 2638
rect 2587 2634 2618 2638
rect 1338 2633 2618 2634
rect 96 2581 97 2587
rect 103 2586 1351 2587
rect 103 2582 111 2586
rect 115 2582 215 2586
rect 219 2582 271 2586
rect 275 2582 327 2586
rect 331 2582 383 2586
rect 387 2582 439 2586
rect 443 2582 495 2586
rect 499 2582 535 2586
rect 539 2582 551 2586
rect 555 2582 591 2586
rect 595 2582 607 2586
rect 611 2582 647 2586
rect 651 2582 663 2586
rect 667 2582 703 2586
rect 707 2582 719 2586
rect 723 2582 759 2586
rect 763 2582 775 2586
rect 779 2582 831 2586
rect 835 2582 887 2586
rect 891 2582 943 2586
rect 947 2582 999 2586
rect 1003 2582 1055 2586
rect 1059 2582 1111 2586
rect 1115 2582 1327 2586
rect 1331 2582 1351 2586
rect 103 2581 1351 2582
rect 1357 2583 1358 2587
rect 1357 2582 2630 2583
rect 1357 2581 1367 2582
rect 1350 2578 1367 2581
rect 1371 2578 1439 2582
rect 1443 2578 1535 2582
rect 1539 2578 1543 2582
rect 1547 2578 1591 2582
rect 1595 2578 1647 2582
rect 1651 2578 1655 2582
rect 1659 2578 1703 2582
rect 1707 2578 1759 2582
rect 1763 2578 1767 2582
rect 1771 2578 1815 2582
rect 1819 2578 1871 2582
rect 1875 2578 1879 2582
rect 1883 2578 1927 2582
rect 1931 2578 1983 2582
rect 1987 2578 1991 2582
rect 1995 2578 2039 2582
rect 2043 2578 2095 2582
rect 2099 2578 2111 2582
rect 2115 2578 2151 2582
rect 2155 2578 2231 2582
rect 2235 2578 2351 2582
rect 2355 2578 2583 2582
rect 2587 2578 2630 2582
rect 1350 2577 2630 2578
rect 84 2521 85 2527
rect 91 2526 1339 2527
rect 91 2522 111 2526
rect 115 2522 231 2526
rect 235 2522 287 2526
rect 291 2522 343 2526
rect 347 2522 367 2526
rect 371 2522 399 2526
rect 403 2522 423 2526
rect 427 2522 455 2526
rect 459 2522 487 2526
rect 491 2522 511 2526
rect 515 2522 551 2526
rect 555 2522 567 2526
rect 571 2522 615 2526
rect 619 2522 623 2526
rect 627 2522 679 2526
rect 683 2522 735 2526
rect 739 2522 743 2526
rect 747 2522 791 2526
rect 795 2522 807 2526
rect 811 2522 847 2526
rect 851 2522 871 2526
rect 875 2522 903 2526
rect 907 2522 943 2526
rect 947 2522 959 2526
rect 963 2522 1015 2526
rect 1019 2522 1071 2526
rect 1075 2522 1127 2526
rect 1131 2522 1327 2526
rect 1331 2522 1339 2526
rect 91 2521 1339 2522
rect 1345 2521 1346 2527
rect 1338 2519 1346 2521
rect 1338 2513 1339 2519
rect 1345 2518 2611 2519
rect 1345 2514 1367 2518
rect 1371 2514 1455 2518
rect 1459 2514 1551 2518
rect 1555 2514 1559 2518
rect 1563 2514 1631 2518
rect 1635 2514 1671 2518
rect 1675 2514 1719 2518
rect 1723 2514 1783 2518
rect 1787 2514 1807 2518
rect 1811 2514 1895 2518
rect 1899 2514 1903 2518
rect 1907 2514 1999 2518
rect 2003 2514 2007 2518
rect 2011 2514 2095 2518
rect 2099 2514 2127 2518
rect 2131 2514 2191 2518
rect 2195 2514 2247 2518
rect 2251 2514 2295 2518
rect 2299 2514 2367 2518
rect 2371 2514 2399 2518
rect 2403 2514 2583 2518
rect 2587 2514 2611 2518
rect 1345 2513 2611 2514
rect 2617 2513 2618 2519
rect 96 2461 97 2467
rect 103 2466 1351 2467
rect 103 2462 111 2466
rect 115 2462 271 2466
rect 275 2462 335 2466
rect 339 2462 351 2466
rect 355 2462 399 2466
rect 403 2462 407 2466
rect 411 2462 471 2466
rect 475 2462 535 2466
rect 539 2462 551 2466
rect 555 2462 599 2466
rect 603 2462 631 2466
rect 635 2462 663 2466
rect 667 2462 711 2466
rect 715 2462 727 2466
rect 731 2462 783 2466
rect 787 2462 791 2466
rect 795 2462 855 2466
rect 859 2462 863 2466
rect 867 2462 927 2466
rect 931 2462 943 2466
rect 947 2462 999 2466
rect 1003 2462 1023 2466
rect 1027 2462 1327 2466
rect 1331 2462 1351 2466
rect 103 2461 1351 2462
rect 1357 2463 1358 2467
rect 1357 2462 2630 2463
rect 1357 2461 1367 2462
rect 1350 2458 1367 2461
rect 1371 2458 1535 2462
rect 1539 2458 1615 2462
rect 1619 2458 1647 2462
rect 1651 2458 1703 2462
rect 1707 2458 1767 2462
rect 1771 2458 1791 2462
rect 1795 2458 1839 2462
rect 1843 2458 1887 2462
rect 1891 2458 1911 2462
rect 1915 2458 1983 2462
rect 1987 2458 1991 2462
rect 1995 2458 2079 2462
rect 2083 2458 2167 2462
rect 2171 2458 2175 2462
rect 2179 2458 2263 2462
rect 2267 2458 2279 2462
rect 2283 2458 2359 2462
rect 2363 2458 2383 2462
rect 2387 2458 2455 2462
rect 2459 2458 2527 2462
rect 2531 2458 2583 2462
rect 2587 2458 2630 2462
rect 1350 2457 2630 2458
rect 84 2401 85 2407
rect 91 2406 1339 2407
rect 91 2402 111 2406
rect 115 2402 247 2406
rect 251 2402 287 2406
rect 291 2402 335 2406
rect 339 2402 351 2406
rect 355 2402 415 2406
rect 419 2402 431 2406
rect 435 2402 487 2406
rect 491 2402 527 2406
rect 531 2402 567 2406
rect 571 2402 631 2406
rect 635 2402 647 2406
rect 651 2402 727 2406
rect 731 2402 799 2406
rect 803 2402 823 2406
rect 827 2402 879 2406
rect 883 2402 919 2406
rect 923 2402 959 2406
rect 963 2402 1015 2406
rect 1019 2402 1039 2406
rect 1043 2402 1111 2406
rect 1115 2402 1327 2406
rect 1331 2402 1339 2406
rect 91 2401 1339 2402
rect 1345 2403 1346 2407
rect 1345 2402 2618 2403
rect 1345 2401 1367 2402
rect 1338 2398 1367 2401
rect 1371 2398 1455 2402
rect 1459 2398 1559 2402
rect 1563 2398 1663 2402
rect 1667 2398 1719 2402
rect 1723 2398 1759 2402
rect 1763 2398 1783 2402
rect 1787 2398 1855 2402
rect 1859 2398 1927 2402
rect 1931 2398 1943 2402
rect 1947 2398 2007 2402
rect 2011 2398 2039 2402
rect 2043 2398 2095 2402
rect 2099 2398 2135 2402
rect 2139 2398 2183 2402
rect 2187 2398 2231 2402
rect 2235 2398 2279 2402
rect 2283 2398 2335 2402
rect 2339 2398 2375 2402
rect 2379 2398 2447 2402
rect 2451 2398 2471 2402
rect 2475 2398 2543 2402
rect 2547 2398 2583 2402
rect 2587 2398 2618 2402
rect 1338 2397 2618 2398
rect 96 2345 97 2351
rect 103 2350 1351 2351
rect 103 2346 111 2350
rect 115 2346 159 2350
rect 163 2346 231 2350
rect 235 2346 263 2350
rect 267 2346 319 2350
rect 323 2346 375 2350
rect 379 2346 415 2350
rect 419 2346 487 2350
rect 491 2346 511 2350
rect 515 2346 599 2350
rect 603 2346 615 2350
rect 619 2346 711 2350
rect 715 2346 807 2350
rect 811 2346 815 2350
rect 819 2346 903 2350
rect 907 2346 911 2350
rect 915 2346 999 2350
rect 1003 2346 1007 2350
rect 1011 2346 1095 2350
rect 1099 2346 1103 2350
rect 1107 2346 1199 2350
rect 1203 2346 1327 2350
rect 1331 2346 1351 2350
rect 103 2345 1351 2346
rect 1357 2347 1358 2351
rect 1357 2346 2630 2347
rect 1357 2345 1367 2346
rect 1350 2342 1367 2345
rect 1371 2342 1399 2346
rect 1403 2342 1439 2346
rect 1443 2342 1455 2346
rect 1459 2342 1511 2346
rect 1515 2342 1543 2346
rect 1547 2342 1567 2346
rect 1571 2342 1639 2346
rect 1643 2342 1647 2346
rect 1651 2342 1727 2346
rect 1731 2342 1743 2346
rect 1747 2342 1823 2346
rect 1827 2342 1839 2346
rect 1843 2342 1927 2346
rect 1931 2342 1943 2346
rect 1947 2342 2023 2346
rect 2027 2342 2079 2346
rect 2083 2342 2119 2346
rect 2123 2342 2215 2346
rect 2219 2342 2223 2346
rect 2227 2342 2319 2346
rect 2323 2342 2383 2346
rect 2387 2342 2431 2346
rect 2435 2342 2527 2346
rect 2531 2342 2583 2346
rect 2587 2342 2630 2346
rect 1350 2341 2630 2342
rect 84 2285 85 2291
rect 91 2290 1339 2291
rect 91 2286 111 2290
rect 115 2286 159 2290
rect 163 2286 175 2290
rect 179 2286 247 2290
rect 251 2286 279 2290
rect 283 2286 375 2290
rect 379 2286 391 2290
rect 395 2286 503 2290
rect 507 2286 511 2290
rect 515 2286 615 2290
rect 619 2286 639 2290
rect 643 2286 727 2290
rect 731 2286 767 2290
rect 771 2286 831 2290
rect 835 2286 887 2290
rect 891 2286 927 2290
rect 931 2286 999 2290
rect 1003 2286 1023 2290
rect 1027 2286 1103 2290
rect 1107 2286 1119 2290
rect 1123 2286 1207 2290
rect 1211 2286 1215 2290
rect 1219 2286 1287 2290
rect 1291 2286 1327 2290
rect 1331 2286 1339 2290
rect 91 2285 1339 2286
rect 1345 2285 1346 2291
rect 1338 2283 1346 2285
rect 1338 2277 1339 2283
rect 1345 2282 2611 2283
rect 1345 2278 1367 2282
rect 1371 2278 1415 2282
rect 1419 2278 1471 2282
rect 1475 2278 1495 2282
rect 1499 2278 1527 2282
rect 1531 2278 1583 2282
rect 1587 2278 1615 2282
rect 1619 2278 1655 2282
rect 1659 2278 1735 2282
rect 1739 2278 1743 2282
rect 1747 2278 1839 2282
rect 1843 2278 1855 2282
rect 1859 2278 1959 2282
rect 1963 2278 1967 2282
rect 1971 2278 2071 2282
rect 2075 2278 2095 2282
rect 2099 2278 2167 2282
rect 2171 2278 2239 2282
rect 2243 2278 2255 2282
rect 2259 2278 2335 2282
rect 2339 2278 2399 2282
rect 2403 2278 2407 2282
rect 2411 2278 2487 2282
rect 2491 2278 2543 2282
rect 2547 2278 2583 2282
rect 2587 2278 2611 2282
rect 1345 2277 2611 2278
rect 2617 2277 2618 2283
rect 96 2221 97 2227
rect 103 2226 1351 2227
rect 103 2222 111 2226
rect 115 2222 143 2226
rect 147 2222 231 2226
rect 235 2222 359 2226
rect 363 2222 495 2226
rect 499 2222 623 2226
rect 627 2222 751 2226
rect 755 2222 871 2226
rect 875 2222 983 2226
rect 987 2222 1087 2226
rect 1091 2222 1191 2226
rect 1195 2222 1271 2226
rect 1275 2222 1327 2226
rect 1331 2222 1351 2226
rect 103 2221 1351 2222
rect 1357 2221 1358 2227
rect 1350 2209 1351 2215
rect 1357 2214 2623 2215
rect 1357 2210 1367 2214
rect 1371 2210 1399 2214
rect 1403 2210 1455 2214
rect 1459 2210 1479 2214
rect 1483 2210 1535 2214
rect 1539 2210 1599 2214
rect 1603 2210 1631 2214
rect 1635 2210 1719 2214
rect 1723 2210 1743 2214
rect 1747 2210 1839 2214
rect 1843 2210 1863 2214
rect 1867 2210 1951 2214
rect 1955 2210 1983 2214
rect 1987 2210 2055 2214
rect 2059 2210 2095 2214
rect 2099 2210 2151 2214
rect 2155 2210 2207 2214
rect 2211 2210 2239 2214
rect 2243 2210 2311 2214
rect 2315 2210 2319 2214
rect 2323 2210 2391 2214
rect 2395 2210 2423 2214
rect 2427 2210 2471 2214
rect 2475 2210 2527 2214
rect 2531 2210 2583 2214
rect 2587 2210 2623 2214
rect 1357 2209 2623 2210
rect 2629 2209 2630 2215
rect 84 2161 85 2167
rect 91 2166 1339 2167
rect 91 2162 111 2166
rect 115 2162 159 2166
rect 163 2162 215 2166
rect 219 2162 247 2166
rect 251 2162 311 2166
rect 315 2162 375 2166
rect 379 2162 423 2166
rect 427 2162 511 2166
rect 515 2162 543 2166
rect 547 2162 639 2166
rect 643 2162 663 2166
rect 667 2162 767 2166
rect 771 2162 775 2166
rect 779 2162 879 2166
rect 883 2162 887 2166
rect 891 2162 975 2166
rect 979 2162 999 2166
rect 1003 2162 1071 2166
rect 1075 2162 1103 2166
rect 1107 2162 1167 2166
rect 1171 2162 1207 2166
rect 1211 2162 1271 2166
rect 1275 2162 1287 2166
rect 1291 2162 1327 2166
rect 1331 2162 1339 2166
rect 91 2161 1339 2162
rect 1345 2161 1346 2167
rect 1338 2159 1346 2161
rect 1338 2153 1339 2159
rect 1345 2158 2611 2159
rect 1345 2154 1367 2158
rect 1371 2154 1471 2158
rect 1475 2154 1535 2158
rect 1539 2154 1551 2158
rect 1555 2154 1631 2158
rect 1635 2154 1647 2158
rect 1651 2154 1735 2158
rect 1739 2154 1759 2158
rect 1763 2154 1839 2158
rect 1843 2154 1879 2158
rect 1883 2154 1951 2158
rect 1955 2154 1999 2158
rect 2003 2154 2055 2158
rect 2059 2154 2111 2158
rect 2115 2154 2159 2158
rect 2163 2154 2223 2158
rect 2227 2154 2263 2158
rect 2267 2154 2327 2158
rect 2331 2154 2359 2158
rect 2363 2154 2439 2158
rect 2443 2154 2463 2158
rect 2467 2154 2543 2158
rect 2547 2154 2583 2158
rect 2587 2154 2611 2158
rect 1345 2153 2611 2154
rect 2617 2153 2618 2159
rect 96 2097 97 2103
rect 103 2102 1351 2103
rect 103 2098 111 2102
rect 115 2098 143 2102
rect 147 2098 199 2102
rect 203 2098 263 2102
rect 267 2098 295 2102
rect 299 2098 327 2102
rect 331 2098 399 2102
rect 403 2098 407 2102
rect 411 2098 479 2102
rect 483 2098 527 2102
rect 531 2098 567 2102
rect 571 2098 647 2102
rect 651 2098 655 2102
rect 659 2098 735 2102
rect 739 2098 759 2102
rect 763 2098 815 2102
rect 819 2098 863 2102
rect 867 2098 887 2102
rect 891 2098 959 2102
rect 963 2098 967 2102
rect 971 2098 1047 2102
rect 1051 2098 1055 2102
rect 1059 2098 1127 2102
rect 1131 2098 1151 2102
rect 1155 2098 1255 2102
rect 1259 2098 1327 2102
rect 1331 2098 1351 2102
rect 103 2097 1351 2098
rect 1357 2102 2630 2103
rect 1357 2098 1367 2102
rect 1371 2098 1431 2102
rect 1435 2098 1519 2102
rect 1523 2098 1535 2102
rect 1539 2098 1615 2102
rect 1619 2098 1647 2102
rect 1651 2098 1719 2102
rect 1723 2098 1759 2102
rect 1763 2098 1823 2102
rect 1827 2098 1863 2102
rect 1867 2098 1935 2102
rect 1939 2098 1967 2102
rect 1971 2098 2039 2102
rect 2043 2098 2071 2102
rect 2075 2098 2143 2102
rect 2147 2098 2175 2102
rect 2179 2098 2247 2102
rect 2251 2098 2271 2102
rect 2275 2098 2343 2102
rect 2347 2098 2359 2102
rect 2363 2098 2447 2102
rect 2451 2098 2455 2102
rect 2459 2098 2527 2102
rect 2531 2098 2583 2102
rect 2587 2098 2630 2102
rect 1357 2097 2630 2098
rect 1338 2041 1339 2047
rect 1345 2046 2611 2047
rect 1345 2042 1367 2046
rect 1371 2042 1415 2046
rect 1419 2042 1447 2046
rect 1451 2042 1503 2046
rect 1507 2042 1551 2046
rect 1555 2042 1607 2046
rect 1611 2042 1663 2046
rect 1667 2042 1711 2046
rect 1715 2042 1775 2046
rect 1779 2042 1807 2046
rect 1811 2042 1879 2046
rect 1883 2042 1903 2046
rect 1907 2042 1983 2046
rect 1987 2042 2007 2046
rect 2011 2042 2087 2046
rect 2091 2042 2111 2046
rect 2115 2042 2191 2046
rect 2195 2042 2215 2046
rect 2219 2042 2287 2046
rect 2291 2042 2327 2046
rect 2331 2042 2375 2046
rect 2379 2042 2447 2046
rect 2451 2042 2471 2046
rect 2475 2042 2543 2046
rect 2547 2042 2583 2046
rect 2587 2042 2611 2046
rect 1345 2041 2611 2042
rect 2617 2041 2618 2047
rect 1338 2039 1346 2041
rect 84 2033 85 2039
rect 91 2038 1339 2039
rect 91 2034 111 2038
rect 115 2034 279 2038
rect 283 2034 343 2038
rect 347 2034 415 2038
rect 419 2034 471 2038
rect 475 2034 495 2038
rect 499 2034 527 2038
rect 531 2034 583 2038
rect 587 2034 639 2038
rect 643 2034 671 2038
rect 675 2034 695 2038
rect 699 2034 751 2038
rect 755 2034 807 2038
rect 811 2034 831 2038
rect 835 2034 863 2038
rect 867 2034 903 2038
rect 907 2034 919 2038
rect 923 2034 975 2038
rect 979 2034 983 2038
rect 987 2034 1031 2038
rect 1035 2034 1063 2038
rect 1067 2034 1143 2038
rect 1147 2034 1327 2038
rect 1331 2034 1339 2038
rect 91 2033 1339 2034
rect 1345 2033 1346 2039
rect 1350 1985 1351 1991
rect 1357 1990 2623 1991
rect 1357 1986 1367 1990
rect 1371 1986 1399 1990
rect 1403 1986 1479 1990
rect 1483 1986 1487 1990
rect 1491 1986 1583 1990
rect 1587 1986 1591 1990
rect 1595 1986 1679 1990
rect 1683 1986 1695 1990
rect 1699 1986 1767 1990
rect 1771 1986 1791 1990
rect 1795 1986 1847 1990
rect 1851 1986 1887 1990
rect 1891 1986 1927 1990
rect 1931 1986 1991 1990
rect 1995 1986 2007 1990
rect 2011 1986 2087 1990
rect 2091 1986 2095 1990
rect 2099 1986 2199 1990
rect 2203 1986 2311 1990
rect 2315 1986 2431 1990
rect 2435 1986 2527 1990
rect 2531 1986 2583 1990
rect 2587 1986 2623 1990
rect 1357 1985 2623 1986
rect 2629 1985 2630 1991
rect 96 1973 97 1979
rect 103 1978 1351 1979
rect 103 1974 111 1978
rect 115 1974 335 1978
rect 339 1974 391 1978
rect 395 1974 399 1978
rect 403 1974 447 1978
rect 451 1974 455 1978
rect 459 1974 503 1978
rect 507 1974 511 1978
rect 515 1974 567 1978
rect 571 1974 623 1978
rect 627 1974 647 1978
rect 651 1974 679 1978
rect 683 1974 735 1978
rect 739 1974 743 1978
rect 747 1974 791 1978
rect 795 1974 847 1978
rect 851 1974 863 1978
rect 867 1974 903 1978
rect 907 1974 959 1978
rect 963 1974 999 1978
rect 1003 1974 1015 1978
rect 1019 1974 1143 1978
rect 1147 1974 1271 1978
rect 1275 1974 1327 1978
rect 1331 1974 1351 1978
rect 103 1973 1351 1974
rect 1357 1973 1358 1979
rect 1338 1925 1339 1931
rect 1345 1930 2611 1931
rect 1345 1926 1367 1930
rect 1371 1926 1415 1930
rect 1419 1926 1495 1930
rect 1499 1926 1599 1930
rect 1603 1926 1695 1930
rect 1699 1926 1719 1930
rect 1723 1926 1775 1930
rect 1779 1926 1783 1930
rect 1787 1926 1831 1930
rect 1835 1926 1863 1930
rect 1867 1926 1887 1930
rect 1891 1926 1943 1930
rect 1947 1926 1999 1930
rect 2003 1926 2023 1930
rect 2027 1926 2055 1930
rect 2059 1926 2103 1930
rect 2107 1926 2119 1930
rect 2123 1926 2583 1930
rect 2587 1926 2611 1930
rect 1345 1925 2611 1926
rect 2617 1925 2618 1931
rect 1338 1923 1346 1925
rect 84 1917 85 1923
rect 91 1922 1339 1923
rect 91 1918 111 1922
rect 115 1918 159 1922
rect 163 1918 231 1922
rect 235 1918 327 1922
rect 331 1918 351 1922
rect 355 1918 407 1922
rect 411 1918 431 1922
rect 435 1918 463 1922
rect 467 1918 519 1922
rect 523 1918 543 1922
rect 547 1918 583 1922
rect 587 1918 655 1922
rect 659 1918 663 1922
rect 667 1918 759 1922
rect 763 1918 767 1922
rect 771 1918 879 1922
rect 883 1918 983 1922
rect 987 1918 1015 1922
rect 1019 1918 1087 1922
rect 1091 1918 1159 1922
rect 1163 1918 1199 1922
rect 1203 1918 1287 1922
rect 1291 1918 1327 1922
rect 1331 1918 1339 1922
rect 91 1917 1339 1918
rect 1345 1917 1346 1923
rect 1350 1865 1351 1871
rect 1357 1870 2623 1871
rect 1357 1866 1367 1870
rect 1371 1866 1399 1870
rect 1403 1866 1463 1870
rect 1467 1866 1559 1870
rect 1563 1866 1655 1870
rect 1659 1866 1703 1870
rect 1707 1866 1743 1870
rect 1747 1866 1759 1870
rect 1763 1866 1815 1870
rect 1819 1866 1831 1870
rect 1835 1866 1871 1870
rect 1875 1866 1919 1870
rect 1923 1866 1927 1870
rect 1931 1866 1983 1870
rect 1987 1866 2007 1870
rect 2011 1866 2039 1870
rect 2043 1866 2095 1870
rect 2099 1866 2103 1870
rect 2107 1866 2183 1870
rect 2187 1866 2583 1870
rect 2587 1866 2623 1870
rect 1357 1865 2623 1866
rect 2629 1865 2630 1871
rect 96 1853 97 1859
rect 103 1858 1351 1859
rect 103 1854 111 1858
rect 115 1854 143 1858
rect 147 1854 199 1858
rect 203 1854 215 1858
rect 219 1854 263 1858
rect 267 1854 311 1858
rect 315 1854 351 1858
rect 355 1854 415 1858
rect 419 1854 439 1858
rect 443 1854 527 1858
rect 531 1854 535 1858
rect 539 1854 623 1858
rect 627 1854 639 1858
rect 643 1854 711 1858
rect 715 1854 751 1858
rect 755 1854 791 1858
rect 795 1854 863 1858
rect 867 1854 871 1858
rect 875 1854 951 1858
rect 955 1854 967 1858
rect 971 1854 1039 1858
rect 1043 1854 1071 1858
rect 1075 1854 1183 1858
rect 1187 1854 1271 1858
rect 1275 1854 1327 1858
rect 1331 1854 1351 1858
rect 103 1853 1351 1854
rect 1357 1853 1358 1859
rect 1338 1809 1339 1815
rect 1345 1814 2611 1815
rect 1345 1810 1367 1814
rect 1371 1810 1415 1814
rect 1419 1810 1479 1814
rect 1483 1810 1511 1814
rect 1515 1810 1575 1814
rect 1579 1810 1623 1814
rect 1627 1810 1671 1814
rect 1675 1810 1735 1814
rect 1739 1810 1759 1814
rect 1763 1810 1839 1814
rect 1843 1810 1847 1814
rect 1851 1810 1935 1814
rect 1939 1810 1951 1814
rect 1955 1810 2023 1814
rect 2027 1810 2063 1814
rect 2067 1810 2111 1814
rect 2115 1810 2183 1814
rect 2187 1810 2199 1814
rect 2203 1810 2303 1814
rect 2307 1810 2431 1814
rect 2435 1810 2543 1814
rect 2547 1810 2583 1814
rect 2587 1810 2611 1814
rect 1345 1809 2611 1810
rect 2617 1809 2618 1815
rect 84 1793 85 1799
rect 91 1798 1339 1799
rect 91 1794 111 1798
rect 115 1794 159 1798
rect 163 1794 215 1798
rect 219 1794 231 1798
rect 235 1794 279 1798
rect 283 1794 295 1798
rect 299 1794 367 1798
rect 371 1794 447 1798
rect 451 1794 455 1798
rect 459 1794 535 1798
rect 539 1794 551 1798
rect 555 1794 623 1798
rect 627 1794 639 1798
rect 643 1794 711 1798
rect 715 1794 727 1798
rect 731 1794 791 1798
rect 795 1794 807 1798
rect 811 1794 871 1798
rect 875 1794 887 1798
rect 891 1794 951 1798
rect 955 1794 967 1798
rect 971 1794 1031 1798
rect 1035 1794 1055 1798
rect 1059 1794 1119 1798
rect 1123 1794 1327 1798
rect 1331 1794 1339 1798
rect 91 1793 1339 1794
rect 1345 1793 1346 1799
rect 1350 1753 1351 1759
rect 1357 1758 2623 1759
rect 1357 1754 1367 1758
rect 1371 1754 1399 1758
rect 1403 1754 1439 1758
rect 1443 1754 1495 1758
rect 1499 1754 1519 1758
rect 1523 1754 1607 1758
rect 1611 1754 1615 1758
rect 1619 1754 1719 1758
rect 1723 1754 1823 1758
rect 1827 1754 1927 1758
rect 1931 1754 1935 1758
rect 1939 1754 2023 1758
rect 2027 1754 2047 1758
rect 2051 1754 2119 1758
rect 2123 1754 2167 1758
rect 2171 1754 2207 1758
rect 2211 1754 2287 1758
rect 2291 1754 2375 1758
rect 2379 1754 2415 1758
rect 2419 1754 2463 1758
rect 2467 1754 2527 1758
rect 2531 1754 2583 1758
rect 2587 1754 2623 1758
rect 1357 1753 2623 1754
rect 2629 1753 2630 1759
rect 96 1733 97 1739
rect 103 1738 1351 1739
rect 103 1734 111 1738
rect 115 1734 215 1738
rect 219 1734 279 1738
rect 283 1734 351 1738
rect 355 1734 407 1738
rect 411 1734 431 1738
rect 435 1734 471 1738
rect 475 1734 519 1738
rect 523 1734 551 1738
rect 555 1734 607 1738
rect 611 1734 639 1738
rect 643 1734 695 1738
rect 699 1734 727 1738
rect 731 1734 775 1738
rect 779 1734 823 1738
rect 827 1734 855 1738
rect 859 1734 919 1738
rect 923 1734 935 1738
rect 939 1734 1015 1738
rect 1019 1734 1103 1738
rect 1107 1734 1111 1738
rect 1115 1734 1207 1738
rect 1211 1734 1327 1738
rect 1331 1734 1351 1738
rect 103 1733 1351 1734
rect 1357 1733 1358 1739
rect 1338 1685 1339 1691
rect 1345 1690 2611 1691
rect 1345 1686 1367 1690
rect 1371 1686 1455 1690
rect 1459 1686 1535 1690
rect 1539 1686 1559 1690
rect 1563 1686 1631 1690
rect 1635 1686 1711 1690
rect 1715 1686 1735 1690
rect 1739 1686 1799 1690
rect 1803 1686 1839 1690
rect 1843 1686 1887 1690
rect 1891 1686 1943 1690
rect 1947 1686 1975 1690
rect 1979 1686 2039 1690
rect 2043 1686 2063 1690
rect 2067 1686 2135 1690
rect 2139 1686 2143 1690
rect 2147 1686 2215 1690
rect 2219 1686 2223 1690
rect 2227 1686 2287 1690
rect 2291 1686 2303 1690
rect 2307 1686 2351 1690
rect 2355 1686 2391 1690
rect 2395 1686 2423 1690
rect 2427 1686 2479 1690
rect 2483 1686 2487 1690
rect 2491 1686 2543 1690
rect 2547 1686 2583 1690
rect 2587 1686 2611 1690
rect 1345 1685 2611 1686
rect 2617 1685 2618 1691
rect 84 1673 85 1679
rect 91 1678 1339 1679
rect 91 1674 111 1678
rect 115 1674 367 1678
rect 371 1674 399 1678
rect 403 1674 423 1678
rect 427 1674 455 1678
rect 459 1674 487 1678
rect 491 1674 511 1678
rect 515 1674 567 1678
rect 571 1674 575 1678
rect 579 1674 647 1678
rect 651 1674 655 1678
rect 659 1674 727 1678
rect 731 1674 743 1678
rect 747 1674 807 1678
rect 811 1674 839 1678
rect 843 1674 887 1678
rect 891 1674 935 1678
rect 939 1674 967 1678
rect 971 1674 1031 1678
rect 1035 1674 1047 1678
rect 1051 1674 1127 1678
rect 1131 1674 1135 1678
rect 1139 1674 1223 1678
rect 1227 1674 1287 1678
rect 1291 1674 1327 1678
rect 1331 1674 1339 1678
rect 91 1673 1339 1674
rect 1345 1673 1346 1679
rect 1350 1617 1351 1623
rect 1357 1622 2623 1623
rect 1357 1618 1367 1622
rect 1371 1618 1543 1622
rect 1547 1618 1575 1622
rect 1579 1618 1615 1622
rect 1619 1618 1631 1622
rect 1635 1618 1687 1622
rect 1691 1618 1695 1622
rect 1699 1618 1751 1622
rect 1755 1618 1783 1622
rect 1787 1618 1831 1622
rect 1835 1618 1871 1622
rect 1875 1618 1919 1622
rect 1923 1618 1959 1622
rect 1963 1618 2007 1622
rect 2011 1618 2047 1622
rect 2051 1618 2103 1622
rect 2107 1618 2127 1622
rect 2131 1618 2199 1622
rect 2203 1618 2207 1622
rect 2211 1618 2271 1622
rect 2275 1618 2319 1622
rect 2323 1618 2335 1622
rect 2339 1618 2407 1622
rect 2411 1618 2431 1622
rect 2435 1618 2471 1622
rect 2475 1618 2527 1622
rect 2531 1618 2583 1622
rect 2587 1618 2623 1622
rect 1357 1617 2623 1618
rect 2629 1617 2630 1623
rect 96 1601 97 1607
rect 103 1606 1351 1607
rect 103 1602 111 1606
rect 115 1602 287 1606
rect 291 1602 367 1606
rect 371 1602 383 1606
rect 387 1602 439 1606
rect 443 1602 455 1606
rect 459 1602 495 1606
rect 499 1602 551 1606
rect 555 1602 559 1606
rect 563 1602 631 1606
rect 635 1602 647 1606
rect 651 1602 711 1606
rect 715 1602 735 1606
rect 739 1602 791 1606
rect 795 1602 823 1606
rect 827 1602 871 1606
rect 875 1602 903 1606
rect 907 1602 951 1606
rect 955 1602 983 1606
rect 987 1602 1031 1606
rect 1035 1602 1063 1606
rect 1067 1602 1119 1606
rect 1123 1602 1151 1606
rect 1155 1602 1207 1606
rect 1211 1602 1271 1606
rect 1275 1602 1327 1606
rect 1331 1602 1351 1606
rect 103 1601 1351 1602
rect 1357 1601 1358 1607
rect 1338 1557 1339 1563
rect 1345 1562 2611 1563
rect 1345 1558 1367 1562
rect 1371 1558 1591 1562
rect 1595 1558 1647 1562
rect 1651 1558 1679 1562
rect 1683 1558 1703 1562
rect 1707 1558 1735 1562
rect 1739 1558 1767 1562
rect 1771 1558 1791 1562
rect 1795 1558 1847 1562
rect 1851 1558 1855 1562
rect 1859 1558 1927 1562
rect 1931 1558 1935 1562
rect 1939 1558 2007 1562
rect 2011 1558 2023 1562
rect 2027 1558 2087 1562
rect 2091 1558 2119 1562
rect 2123 1558 2167 1562
rect 2171 1558 2223 1562
rect 2227 1558 2247 1562
rect 2251 1558 2327 1562
rect 2331 1558 2335 1562
rect 2339 1558 2407 1562
rect 2411 1558 2447 1562
rect 2451 1558 2487 1562
rect 2491 1558 2543 1562
rect 2547 1558 2583 1562
rect 2587 1558 2611 1562
rect 1345 1557 2611 1558
rect 2617 1557 2618 1563
rect 84 1545 85 1551
rect 91 1550 1339 1551
rect 91 1546 111 1550
rect 115 1546 279 1550
rect 283 1546 303 1550
rect 307 1546 335 1550
rect 339 1546 383 1550
rect 387 1546 399 1550
rect 403 1546 471 1550
rect 475 1546 543 1550
rect 547 1546 567 1550
rect 571 1546 615 1550
rect 619 1546 663 1550
rect 667 1546 687 1550
rect 691 1546 751 1550
rect 755 1546 759 1550
rect 763 1546 831 1550
rect 835 1546 839 1550
rect 843 1546 903 1550
rect 907 1546 919 1550
rect 923 1546 975 1550
rect 979 1546 999 1550
rect 1003 1546 1055 1550
rect 1059 1546 1079 1550
rect 1083 1546 1167 1550
rect 1171 1546 1327 1550
rect 1331 1546 1339 1550
rect 91 1545 1339 1546
rect 1345 1545 1346 1551
rect 1350 1493 1351 1499
rect 1357 1498 2623 1499
rect 1357 1494 1367 1498
rect 1371 1494 1519 1498
rect 1523 1494 1575 1498
rect 1579 1494 1647 1498
rect 1651 1494 1663 1498
rect 1667 1494 1719 1498
rect 1723 1494 1727 1498
rect 1731 1494 1775 1498
rect 1779 1494 1807 1498
rect 1811 1494 1839 1498
rect 1843 1494 1895 1498
rect 1899 1494 1911 1498
rect 1915 1494 1983 1498
rect 1987 1494 1991 1498
rect 1995 1494 2071 1498
rect 2075 1494 2151 1498
rect 2155 1494 2231 1498
rect 2235 1494 2311 1498
rect 2315 1494 2391 1498
rect 2395 1494 2471 1498
rect 2475 1494 2527 1498
rect 2531 1494 2583 1498
rect 2587 1494 2623 1498
rect 1357 1493 2623 1494
rect 2629 1493 2630 1499
rect 1350 1491 1358 1493
rect 96 1485 97 1491
rect 103 1490 1351 1491
rect 103 1486 111 1490
rect 115 1486 199 1490
rect 203 1486 263 1490
rect 267 1486 287 1490
rect 291 1486 319 1490
rect 323 1486 383 1490
rect 387 1486 455 1490
rect 459 1486 487 1490
rect 491 1486 527 1490
rect 531 1486 583 1490
rect 587 1486 599 1490
rect 603 1486 671 1490
rect 675 1486 679 1490
rect 683 1486 743 1490
rect 747 1486 775 1490
rect 779 1486 815 1490
rect 819 1486 863 1490
rect 867 1486 887 1490
rect 891 1486 951 1490
rect 955 1486 959 1490
rect 963 1486 1039 1490
rect 1043 1486 1135 1490
rect 1139 1486 1327 1490
rect 1331 1486 1351 1490
rect 103 1485 1351 1486
rect 1357 1485 1358 1491
rect 1338 1434 2618 1435
rect 1338 1431 1367 1434
rect 84 1425 85 1431
rect 91 1430 1339 1431
rect 91 1426 111 1430
rect 115 1426 159 1430
rect 163 1426 215 1430
rect 219 1426 247 1430
rect 251 1426 303 1430
rect 307 1426 343 1430
rect 347 1426 399 1430
rect 403 1426 447 1430
rect 451 1426 503 1430
rect 507 1426 551 1430
rect 555 1426 599 1430
rect 603 1426 663 1430
rect 667 1426 695 1430
rect 699 1426 767 1430
rect 771 1426 791 1430
rect 795 1426 879 1430
rect 883 1426 967 1430
rect 971 1426 991 1430
rect 995 1426 1055 1430
rect 1059 1426 1103 1430
rect 1107 1426 1151 1430
rect 1155 1426 1215 1430
rect 1219 1426 1327 1430
rect 1331 1426 1339 1430
rect 91 1425 1339 1426
rect 1345 1430 1367 1431
rect 1371 1430 1415 1434
rect 1419 1430 1471 1434
rect 1475 1430 1535 1434
rect 1539 1430 1591 1434
rect 1595 1430 1623 1434
rect 1627 1430 1663 1434
rect 1667 1430 1719 1434
rect 1723 1430 1743 1434
rect 1747 1430 1823 1434
rect 1827 1430 1911 1434
rect 1915 1430 1927 1434
rect 1931 1430 1999 1434
rect 2003 1430 2023 1434
rect 2027 1430 2087 1434
rect 2091 1430 2119 1434
rect 2123 1430 2167 1434
rect 2171 1430 2215 1434
rect 2219 1430 2247 1434
rect 2251 1430 2303 1434
rect 2307 1430 2327 1434
rect 2331 1430 2391 1434
rect 2395 1430 2407 1434
rect 2411 1430 2479 1434
rect 2483 1430 2487 1434
rect 2491 1430 2543 1434
rect 2547 1430 2583 1434
rect 2587 1430 2618 1434
rect 1345 1429 2618 1430
rect 1345 1425 1346 1429
rect 96 1369 97 1375
rect 103 1374 1351 1375
rect 103 1370 111 1374
rect 115 1370 143 1374
rect 147 1370 207 1374
rect 211 1370 231 1374
rect 235 1370 295 1374
rect 299 1370 327 1374
rect 331 1370 399 1374
rect 403 1370 431 1374
rect 435 1370 511 1374
rect 515 1370 535 1374
rect 539 1370 623 1374
rect 627 1370 647 1374
rect 651 1370 735 1374
rect 739 1370 751 1374
rect 755 1370 847 1374
rect 851 1370 863 1374
rect 867 1370 959 1374
rect 963 1370 975 1374
rect 979 1370 1071 1374
rect 1075 1370 1087 1374
rect 1091 1370 1183 1374
rect 1187 1370 1199 1374
rect 1203 1370 1271 1374
rect 1275 1370 1327 1374
rect 1331 1370 1351 1374
rect 103 1369 1351 1370
rect 1357 1371 1358 1375
rect 1357 1370 2630 1371
rect 1357 1369 1367 1370
rect 1350 1366 1367 1369
rect 1371 1366 1399 1370
rect 1403 1366 1455 1370
rect 1459 1366 1519 1370
rect 1523 1366 1543 1370
rect 1547 1366 1607 1370
rect 1611 1366 1631 1370
rect 1635 1366 1703 1370
rect 1707 1366 1719 1370
rect 1723 1366 1807 1370
rect 1811 1366 1887 1370
rect 1891 1366 1911 1370
rect 1915 1366 1967 1370
rect 1971 1366 2007 1370
rect 2011 1366 2047 1370
rect 2051 1366 2103 1370
rect 2107 1366 2127 1370
rect 2131 1366 2199 1370
rect 2203 1366 2207 1370
rect 2211 1366 2287 1370
rect 2291 1366 2375 1370
rect 2379 1366 2463 1370
rect 2467 1366 2527 1370
rect 2531 1366 2583 1370
rect 2587 1366 2630 1370
rect 1350 1365 2630 1366
rect 84 1313 85 1319
rect 91 1318 1339 1319
rect 91 1314 111 1318
rect 115 1314 159 1318
rect 163 1314 223 1318
rect 227 1314 231 1318
rect 235 1314 311 1318
rect 315 1314 327 1318
rect 331 1314 415 1318
rect 419 1314 431 1318
rect 435 1314 527 1318
rect 531 1314 535 1318
rect 539 1314 631 1318
rect 635 1314 639 1318
rect 643 1314 727 1318
rect 731 1314 751 1318
rect 755 1314 823 1318
rect 827 1314 863 1318
rect 867 1314 911 1318
rect 915 1314 975 1318
rect 979 1314 991 1318
rect 995 1314 1071 1318
rect 1075 1314 1087 1318
rect 1091 1314 1151 1318
rect 1155 1314 1199 1318
rect 1203 1314 1231 1318
rect 1235 1314 1287 1318
rect 1291 1314 1327 1318
rect 1331 1314 1339 1318
rect 91 1313 1339 1314
rect 1345 1313 1346 1319
rect 1338 1311 1346 1313
rect 1338 1305 1339 1311
rect 1345 1310 2611 1311
rect 1345 1306 1367 1310
rect 1371 1306 1415 1310
rect 1419 1306 1471 1310
rect 1475 1306 1559 1310
rect 1563 1306 1647 1310
rect 1651 1306 1671 1310
rect 1675 1306 1735 1310
rect 1739 1306 1767 1310
rect 1771 1306 1823 1310
rect 1827 1306 1863 1310
rect 1867 1306 1903 1310
rect 1907 1306 1959 1310
rect 1963 1306 1983 1310
rect 1987 1306 2047 1310
rect 2051 1306 2063 1310
rect 2067 1306 2135 1310
rect 2139 1306 2143 1310
rect 2147 1306 2223 1310
rect 2227 1306 2231 1310
rect 2235 1306 2583 1310
rect 2587 1306 2611 1310
rect 1345 1305 2611 1306
rect 2617 1305 2618 1311
rect 1350 1254 2630 1255
rect 1350 1251 1367 1254
rect 96 1245 97 1251
rect 103 1250 1351 1251
rect 103 1246 111 1250
rect 115 1246 143 1250
rect 147 1246 199 1250
rect 203 1246 215 1250
rect 219 1246 279 1250
rect 283 1246 311 1250
rect 315 1246 359 1250
rect 363 1246 415 1250
rect 419 1246 439 1250
rect 443 1246 519 1250
rect 523 1246 599 1250
rect 603 1246 615 1250
rect 619 1246 671 1250
rect 675 1246 711 1250
rect 715 1246 743 1250
rect 747 1246 807 1250
rect 811 1246 815 1250
rect 819 1246 895 1250
rect 899 1246 975 1250
rect 979 1246 1055 1250
rect 1059 1246 1135 1250
rect 1139 1246 1215 1250
rect 1219 1246 1271 1250
rect 1275 1246 1327 1250
rect 1331 1246 1351 1250
rect 103 1245 1351 1246
rect 1357 1250 1367 1251
rect 1371 1250 1495 1254
rect 1499 1250 1559 1254
rect 1563 1250 1623 1254
rect 1627 1250 1655 1254
rect 1659 1250 1687 1254
rect 1691 1250 1751 1254
rect 1755 1250 1759 1254
rect 1763 1250 1823 1254
rect 1827 1250 1847 1254
rect 1851 1250 1887 1254
rect 1891 1250 1943 1254
rect 1947 1250 1951 1254
rect 1955 1250 2015 1254
rect 2019 1250 2031 1254
rect 2035 1250 2079 1254
rect 2083 1250 2119 1254
rect 2123 1250 2151 1254
rect 2155 1250 2215 1254
rect 2219 1250 2223 1254
rect 2227 1250 2295 1254
rect 2299 1250 2583 1254
rect 2587 1250 2630 1254
rect 1357 1249 2630 1250
rect 1357 1245 1358 1249
rect 84 1185 85 1191
rect 91 1190 1339 1191
rect 91 1186 111 1190
rect 115 1186 159 1190
rect 163 1186 215 1190
rect 219 1186 239 1190
rect 243 1186 295 1190
rect 299 1186 327 1190
rect 331 1186 375 1190
rect 379 1186 423 1190
rect 427 1186 455 1190
rect 459 1186 511 1190
rect 515 1186 535 1190
rect 539 1186 599 1190
rect 603 1186 615 1190
rect 619 1186 687 1190
rect 691 1186 759 1190
rect 763 1186 767 1190
rect 771 1186 831 1190
rect 835 1186 839 1190
rect 843 1186 911 1190
rect 915 1186 983 1190
rect 987 1186 1063 1190
rect 1067 1186 1327 1190
rect 1331 1186 1339 1190
rect 91 1185 1339 1186
rect 1345 1190 2618 1191
rect 1345 1186 1367 1190
rect 1371 1186 1415 1190
rect 1419 1186 1503 1190
rect 1507 1186 1511 1190
rect 1515 1186 1575 1190
rect 1579 1186 1599 1190
rect 1603 1186 1639 1190
rect 1643 1186 1703 1190
rect 1707 1186 1775 1190
rect 1779 1186 1807 1190
rect 1811 1186 1839 1190
rect 1843 1186 1903 1190
rect 1907 1186 1911 1190
rect 1915 1186 1967 1190
rect 1971 1186 2015 1190
rect 2019 1186 2031 1190
rect 2035 1186 2095 1190
rect 2099 1186 2111 1190
rect 2115 1186 2167 1190
rect 2171 1186 2207 1190
rect 2211 1186 2239 1190
rect 2243 1186 2303 1190
rect 2307 1186 2311 1190
rect 2315 1186 2399 1190
rect 2403 1186 2583 1190
rect 2587 1186 2618 1190
rect 1345 1185 2618 1186
rect 1350 1130 2630 1131
rect 1350 1127 1367 1130
rect 96 1121 97 1127
rect 103 1126 1351 1127
rect 103 1122 111 1126
rect 115 1122 143 1126
rect 147 1122 223 1126
rect 227 1122 311 1126
rect 315 1122 319 1126
rect 323 1122 407 1126
rect 411 1122 423 1126
rect 427 1122 495 1126
rect 499 1122 527 1126
rect 531 1122 583 1126
rect 587 1122 631 1126
rect 635 1122 671 1126
rect 675 1122 727 1126
rect 731 1122 751 1126
rect 755 1122 823 1126
rect 827 1122 895 1126
rect 899 1122 911 1126
rect 915 1122 967 1126
rect 971 1122 991 1126
rect 995 1122 1047 1126
rect 1051 1122 1079 1126
rect 1083 1122 1167 1126
rect 1171 1122 1327 1126
rect 1331 1122 1351 1126
rect 103 1121 1351 1122
rect 1357 1126 1367 1127
rect 1371 1126 1399 1130
rect 1403 1126 1479 1130
rect 1483 1126 1487 1130
rect 1491 1126 1583 1130
rect 1587 1126 1687 1130
rect 1691 1126 1791 1130
rect 1795 1126 1887 1130
rect 1891 1126 1895 1130
rect 1899 1126 1975 1130
rect 1979 1126 1999 1130
rect 2003 1126 2063 1130
rect 2067 1126 2095 1130
rect 2099 1126 2143 1130
rect 2147 1126 2191 1130
rect 2195 1126 2215 1130
rect 2219 1126 2279 1130
rect 2283 1126 2287 1130
rect 2291 1126 2343 1130
rect 2347 1126 2383 1130
rect 2387 1126 2407 1130
rect 2411 1126 2471 1130
rect 2475 1126 2527 1130
rect 2531 1126 2583 1130
rect 2587 1126 2630 1130
rect 1357 1125 2630 1126
rect 1357 1121 1358 1125
rect 1338 1070 2618 1071
rect 1338 1067 1367 1070
rect 84 1061 85 1067
rect 91 1066 1339 1067
rect 91 1062 111 1066
rect 115 1062 239 1066
rect 243 1062 311 1066
rect 315 1062 335 1066
rect 339 1062 367 1066
rect 371 1062 439 1066
rect 443 1062 519 1066
rect 523 1062 543 1066
rect 547 1062 607 1066
rect 611 1062 647 1066
rect 651 1062 703 1066
rect 707 1062 743 1066
rect 747 1062 799 1066
rect 803 1062 839 1066
rect 843 1062 887 1066
rect 891 1062 927 1066
rect 931 1062 975 1066
rect 979 1062 1007 1066
rect 1011 1062 1055 1066
rect 1059 1062 1095 1066
rect 1099 1062 1135 1066
rect 1139 1062 1183 1066
rect 1187 1062 1223 1066
rect 1227 1062 1287 1066
rect 1291 1062 1327 1066
rect 1331 1062 1339 1066
rect 91 1061 1339 1062
rect 1345 1066 1367 1067
rect 1371 1066 1415 1070
rect 1419 1066 1471 1070
rect 1475 1066 1495 1070
rect 1499 1066 1535 1070
rect 1539 1066 1599 1070
rect 1603 1066 1623 1070
rect 1627 1066 1703 1070
rect 1707 1066 1727 1070
rect 1731 1066 1807 1070
rect 1811 1066 1839 1070
rect 1843 1066 1903 1070
rect 1907 1066 1951 1070
rect 1955 1066 1991 1070
rect 1995 1066 2063 1070
rect 2067 1066 2079 1070
rect 2083 1066 2159 1070
rect 2163 1066 2167 1070
rect 2171 1066 2231 1070
rect 2235 1066 2271 1070
rect 2275 1066 2295 1070
rect 2299 1066 2359 1070
rect 2363 1066 2367 1070
rect 2371 1066 2423 1070
rect 2427 1066 2463 1070
rect 2467 1066 2487 1070
rect 2491 1066 2543 1070
rect 2547 1066 2583 1070
rect 2587 1066 2618 1070
rect 1345 1065 2618 1066
rect 1345 1061 1346 1065
rect 96 1001 97 1007
rect 103 1006 1351 1007
rect 103 1002 111 1006
rect 115 1002 295 1006
rect 299 1002 351 1006
rect 355 1002 415 1006
rect 419 1002 423 1006
rect 427 1002 471 1006
rect 475 1002 503 1006
rect 507 1002 527 1006
rect 531 1002 591 1006
rect 595 1002 655 1006
rect 659 1002 687 1006
rect 691 1002 719 1006
rect 723 1002 783 1006
rect 787 1002 847 1006
rect 851 1002 871 1006
rect 875 1002 911 1006
rect 915 1002 959 1006
rect 963 1002 975 1006
rect 979 1002 1039 1006
rect 1043 1002 1103 1006
rect 1107 1002 1119 1006
rect 1123 1002 1159 1006
rect 1163 1002 1207 1006
rect 1211 1002 1215 1006
rect 1219 1002 1271 1006
rect 1275 1002 1327 1006
rect 1331 1002 1351 1006
rect 103 1001 1351 1002
rect 1357 1001 1358 1007
rect 1350 999 1358 1001
rect 1350 993 1351 999
rect 1357 998 2623 999
rect 1357 994 1367 998
rect 1371 994 1399 998
rect 1403 994 1455 998
rect 1459 994 1511 998
rect 1515 994 1519 998
rect 1523 994 1567 998
rect 1571 994 1607 998
rect 1611 994 1639 998
rect 1643 994 1711 998
rect 1715 994 1719 998
rect 1723 994 1807 998
rect 1811 994 1823 998
rect 1827 994 1903 998
rect 1907 994 1935 998
rect 1939 994 2015 998
rect 2019 994 2047 998
rect 2051 994 2143 998
rect 2147 994 2151 998
rect 2155 994 2255 998
rect 2259 994 2271 998
rect 2275 994 2351 998
rect 2355 994 2407 998
rect 2411 994 2447 998
rect 2451 994 2527 998
rect 2531 994 2583 998
rect 2587 994 2623 998
rect 1357 993 2623 994
rect 2629 993 2630 999
rect 84 941 85 947
rect 91 946 1339 947
rect 91 942 111 946
rect 115 942 423 946
rect 427 942 431 946
rect 435 942 479 946
rect 483 942 487 946
rect 491 942 535 946
rect 539 942 543 946
rect 547 942 591 946
rect 595 942 607 946
rect 611 942 647 946
rect 651 942 671 946
rect 675 942 703 946
rect 707 942 735 946
rect 739 942 759 946
rect 763 942 799 946
rect 803 942 815 946
rect 819 942 863 946
rect 867 942 927 946
rect 931 942 991 946
rect 995 942 1055 946
rect 1059 942 1119 946
rect 1123 942 1175 946
rect 1179 942 1231 946
rect 1235 942 1287 946
rect 1291 942 1327 946
rect 1331 942 1339 946
rect 91 941 1339 942
rect 1345 941 1346 947
rect 1338 929 1339 935
rect 1345 934 2611 935
rect 1345 930 1367 934
rect 1371 930 1415 934
rect 1419 930 1471 934
rect 1475 930 1527 934
rect 1531 930 1583 934
rect 1587 930 1615 934
rect 1619 930 1655 934
rect 1659 930 1711 934
rect 1715 930 1735 934
rect 1739 930 1823 934
rect 1827 930 1919 934
rect 1923 930 1943 934
rect 1947 930 2031 934
rect 2035 930 2063 934
rect 2067 930 2159 934
rect 2163 930 2183 934
rect 2187 930 2287 934
rect 2291 930 2311 934
rect 2315 930 2423 934
rect 2427 930 2439 934
rect 2443 930 2543 934
rect 2547 930 2583 934
rect 2587 930 2611 934
rect 1345 929 2611 930
rect 2617 929 2618 935
rect 96 885 97 891
rect 103 890 1351 891
rect 103 886 111 890
rect 115 886 279 890
rect 283 886 335 890
rect 339 886 391 890
rect 395 886 407 890
rect 411 886 455 890
rect 459 886 463 890
rect 467 886 519 890
rect 523 886 575 890
rect 579 886 583 890
rect 587 886 631 890
rect 635 886 647 890
rect 651 886 687 890
rect 691 886 711 890
rect 715 886 743 890
rect 747 886 775 890
rect 779 886 799 890
rect 803 886 847 890
rect 851 886 919 890
rect 923 886 1327 890
rect 1331 886 1351 890
rect 103 885 1351 886
rect 1357 885 1358 891
rect 1350 873 1351 879
rect 1357 878 2623 879
rect 1357 874 1367 878
rect 1371 874 1399 878
rect 1403 874 1455 878
rect 1459 874 1471 878
rect 1475 874 1511 878
rect 1515 874 1551 878
rect 1555 874 1599 878
rect 1603 874 1639 878
rect 1643 874 1695 878
rect 1699 874 1727 878
rect 1731 874 1807 878
rect 1811 874 1815 878
rect 1819 874 1903 878
rect 1907 874 1927 878
rect 1931 874 1991 878
rect 1995 874 2047 878
rect 2051 874 2071 878
rect 2075 874 2143 878
rect 2147 874 2167 878
rect 2171 874 2215 878
rect 2219 874 2279 878
rect 2283 874 2295 878
rect 2299 874 2343 878
rect 2347 874 2407 878
rect 2411 874 2423 878
rect 2427 874 2471 878
rect 2475 874 2527 878
rect 2531 874 2583 878
rect 2587 874 2623 878
rect 1357 873 2623 874
rect 2629 873 2630 879
rect 84 821 85 827
rect 91 826 1339 827
rect 91 822 111 826
rect 115 822 167 826
rect 171 822 231 826
rect 235 822 295 826
rect 299 822 311 826
rect 315 822 351 826
rect 355 822 399 826
rect 403 822 407 826
rect 411 822 471 826
rect 475 822 487 826
rect 491 822 535 826
rect 539 822 583 826
rect 587 822 599 826
rect 603 822 663 826
rect 667 822 671 826
rect 675 822 727 826
rect 731 822 759 826
rect 763 822 791 826
rect 795 822 839 826
rect 843 822 863 826
rect 867 822 919 826
rect 923 822 935 826
rect 939 822 1007 826
rect 1011 822 1095 826
rect 1099 822 1327 826
rect 1331 822 1339 826
rect 91 821 1339 822
rect 1345 821 1346 827
rect 1338 809 1339 815
rect 1345 814 2611 815
rect 1345 810 1367 814
rect 1371 810 1487 814
rect 1491 810 1567 814
rect 1571 810 1631 814
rect 1635 810 1655 814
rect 1659 810 1687 814
rect 1691 810 1743 814
rect 1747 810 1751 814
rect 1755 810 1823 814
rect 1827 810 1831 814
rect 1835 810 1903 814
rect 1907 810 1919 814
rect 1923 810 1991 814
rect 1995 810 2007 814
rect 2011 810 2071 814
rect 2075 810 2087 814
rect 2091 810 2159 814
rect 2163 810 2231 814
rect 2235 810 2247 814
rect 2251 810 2295 814
rect 2299 810 2335 814
rect 2339 810 2359 814
rect 2363 810 2423 814
rect 2427 810 2487 814
rect 2491 810 2543 814
rect 2547 810 2583 814
rect 2587 810 2611 814
rect 1345 809 2611 810
rect 2617 809 2618 815
rect 96 757 97 763
rect 103 762 1351 763
rect 103 758 111 762
rect 115 758 143 762
rect 147 758 151 762
rect 155 758 199 762
rect 203 758 215 762
rect 219 758 279 762
rect 283 758 295 762
rect 299 758 383 762
rect 387 758 471 762
rect 475 758 487 762
rect 491 758 567 762
rect 571 758 599 762
rect 603 758 655 762
rect 659 758 703 762
rect 707 758 743 762
rect 747 758 807 762
rect 811 758 823 762
rect 827 758 903 762
rect 907 758 991 762
rect 995 758 1079 762
rect 1083 758 1175 762
rect 1179 758 1327 762
rect 1331 758 1351 762
rect 103 757 1351 758
rect 1357 757 1358 763
rect 1350 755 1358 757
rect 1350 749 1351 755
rect 1357 754 2623 755
rect 1357 750 1367 754
rect 1371 750 1567 754
rect 1571 750 1615 754
rect 1619 750 1623 754
rect 1627 750 1671 754
rect 1675 750 1687 754
rect 1691 750 1735 754
rect 1739 750 1759 754
rect 1763 750 1807 754
rect 1811 750 1839 754
rect 1843 750 1887 754
rect 1891 750 1919 754
rect 1923 750 1975 754
rect 1979 750 1999 754
rect 2003 750 2055 754
rect 2059 750 2079 754
rect 2083 750 2143 754
rect 2147 750 2159 754
rect 2163 750 2231 754
rect 2235 750 2247 754
rect 2251 750 2319 754
rect 2323 750 2335 754
rect 2339 750 2407 754
rect 2411 750 2583 754
rect 2587 750 2623 754
rect 1357 749 2623 750
rect 2629 749 2630 755
rect 84 697 85 703
rect 91 702 1339 703
rect 91 698 111 702
rect 115 698 159 702
rect 163 698 215 702
rect 219 698 279 702
rect 283 698 295 702
rect 299 698 359 702
rect 363 698 399 702
rect 403 698 447 702
rect 451 698 503 702
rect 507 698 535 702
rect 539 698 615 702
rect 619 698 623 702
rect 627 698 711 702
rect 715 698 719 702
rect 723 698 791 702
rect 795 698 823 702
rect 827 698 871 702
rect 875 698 919 702
rect 923 698 951 702
rect 955 698 1007 702
rect 1011 698 1039 702
rect 1043 698 1095 702
rect 1099 698 1191 702
rect 1195 698 1327 702
rect 1331 698 1339 702
rect 91 697 1339 698
rect 1345 697 1346 703
rect 1338 695 1346 697
rect 1338 689 1339 695
rect 1345 694 2611 695
rect 1345 690 1367 694
rect 1371 690 1415 694
rect 1419 690 1511 694
rect 1515 690 1583 694
rect 1587 690 1615 694
rect 1619 690 1639 694
rect 1643 690 1703 694
rect 1707 690 1719 694
rect 1723 690 1775 694
rect 1779 690 1823 694
rect 1827 690 1855 694
rect 1859 690 1927 694
rect 1931 690 1935 694
rect 1939 690 2015 694
rect 2019 690 2023 694
rect 2027 690 2095 694
rect 2099 690 2119 694
rect 2123 690 2175 694
rect 2179 690 2207 694
rect 2211 690 2263 694
rect 2267 690 2295 694
rect 2299 690 2351 694
rect 2355 690 2391 694
rect 2395 690 2583 694
rect 2587 690 2611 694
rect 1345 689 2611 690
rect 2617 689 2618 695
rect 96 633 97 639
rect 103 638 1351 639
rect 103 634 111 638
rect 115 634 143 638
rect 147 634 199 638
rect 203 634 255 638
rect 259 634 263 638
rect 267 634 311 638
rect 315 634 343 638
rect 347 634 391 638
rect 395 634 431 638
rect 435 634 479 638
rect 483 634 519 638
rect 523 634 575 638
rect 579 634 607 638
rect 611 634 679 638
rect 683 634 695 638
rect 699 634 775 638
rect 779 634 783 638
rect 787 634 855 638
rect 859 634 887 638
rect 891 634 935 638
rect 939 634 991 638
rect 995 634 1023 638
rect 1027 634 1087 638
rect 1091 634 1191 638
rect 1195 634 1271 638
rect 1275 634 1327 638
rect 1331 634 1351 638
rect 103 633 1351 634
rect 1357 638 2630 639
rect 1357 634 1367 638
rect 1371 634 1399 638
rect 1403 634 1495 638
rect 1499 634 1511 638
rect 1515 634 1599 638
rect 1603 634 1647 638
rect 1651 634 1703 638
rect 1707 634 1783 638
rect 1787 634 1807 638
rect 1811 634 1911 638
rect 1915 634 2007 638
rect 2011 634 2039 638
rect 2043 634 2103 638
rect 2107 634 2159 638
rect 2163 634 2191 638
rect 2195 634 2279 638
rect 2283 634 2375 638
rect 2379 634 2407 638
rect 2411 634 2583 638
rect 2587 634 2630 638
rect 1357 633 2630 634
rect 84 573 85 579
rect 91 578 1339 579
rect 91 574 111 578
rect 115 574 159 578
rect 163 574 199 578
rect 203 574 215 578
rect 219 574 263 578
rect 267 574 271 578
rect 275 574 327 578
rect 331 574 335 578
rect 339 574 407 578
rect 411 574 415 578
rect 419 574 495 578
rect 499 574 511 578
rect 515 574 591 578
rect 595 574 615 578
rect 619 574 695 578
rect 699 574 719 578
rect 723 574 799 578
rect 803 574 831 578
rect 835 574 903 578
rect 907 574 943 578
rect 947 574 1007 578
rect 1011 574 1063 578
rect 1067 574 1103 578
rect 1107 574 1183 578
rect 1187 574 1207 578
rect 1211 574 1287 578
rect 1291 574 1327 578
rect 1331 574 1339 578
rect 91 573 1339 574
rect 1345 575 1346 579
rect 1345 574 2618 575
rect 1345 573 1367 574
rect 1338 570 1367 573
rect 1371 570 1415 574
rect 1419 570 1471 574
rect 1475 570 1527 574
rect 1531 570 1551 574
rect 1555 570 1647 574
rect 1651 570 1663 574
rect 1667 570 1751 574
rect 1755 570 1799 574
rect 1803 570 1855 574
rect 1859 570 1927 574
rect 1931 570 1959 574
rect 1963 570 2055 574
rect 2059 570 2151 574
rect 2155 570 2175 574
rect 2179 570 2239 574
rect 2243 570 2295 574
rect 2299 570 2319 574
rect 2323 570 2399 574
rect 2403 570 2423 574
rect 2427 570 2479 574
rect 2483 570 2543 574
rect 2547 570 2583 574
rect 2587 570 2618 574
rect 1338 569 2618 570
rect 1350 518 2630 519
rect 1350 515 1367 518
rect 96 509 97 515
rect 103 514 1351 515
rect 103 510 111 514
rect 115 510 183 514
rect 187 510 247 514
rect 251 510 303 514
rect 307 510 319 514
rect 323 510 359 514
rect 363 510 399 514
rect 403 510 423 514
rect 427 510 495 514
rect 499 510 575 514
rect 579 510 599 514
rect 603 510 647 514
rect 651 510 703 514
rect 707 510 719 514
rect 723 510 791 514
rect 795 510 815 514
rect 819 510 863 514
rect 867 510 927 514
rect 931 510 935 514
rect 939 510 1007 514
rect 1011 510 1047 514
rect 1051 510 1087 514
rect 1091 510 1167 514
rect 1171 510 1271 514
rect 1275 510 1327 514
rect 1331 510 1351 514
rect 103 509 1351 510
rect 1357 514 1367 515
rect 1371 514 1399 518
rect 1403 514 1455 518
rect 1459 514 1535 518
rect 1539 514 1599 518
rect 1603 514 1631 518
rect 1635 514 1671 518
rect 1675 514 1735 518
rect 1739 514 1751 518
rect 1755 514 1839 518
rect 1843 514 1927 518
rect 1931 514 1943 518
rect 1947 514 2015 518
rect 2019 514 2039 518
rect 2043 514 2095 518
rect 2099 514 2135 518
rect 2139 514 2175 518
rect 2179 514 2223 518
rect 2227 514 2255 518
rect 2259 514 2303 518
rect 2307 514 2327 518
rect 2331 514 2383 518
rect 2387 514 2399 518
rect 2403 514 2463 518
rect 2467 514 2471 518
rect 2475 514 2527 518
rect 2531 514 2583 518
rect 2587 514 2630 518
rect 1357 513 2630 514
rect 1357 509 1358 513
rect 84 449 85 455
rect 91 454 1339 455
rect 91 450 111 454
rect 115 450 319 454
rect 323 450 375 454
rect 379 450 439 454
rect 443 450 455 454
rect 459 450 511 454
rect 515 450 575 454
rect 579 450 591 454
rect 595 450 647 454
rect 651 450 663 454
rect 667 450 727 454
rect 731 450 735 454
rect 739 450 799 454
rect 803 450 807 454
rect 811 450 871 454
rect 875 450 879 454
rect 883 450 943 454
rect 947 450 951 454
rect 955 450 1015 454
rect 1019 450 1023 454
rect 1027 450 1087 454
rect 1091 450 1103 454
rect 1107 450 1159 454
rect 1163 450 1239 454
rect 1243 450 1327 454
rect 1331 450 1339 454
rect 91 449 1339 450
rect 1345 454 2618 455
rect 1345 450 1367 454
rect 1371 450 1551 454
rect 1555 450 1615 454
rect 1619 450 1647 454
rect 1651 450 1687 454
rect 1691 450 1703 454
rect 1707 450 1759 454
rect 1763 450 1767 454
rect 1771 450 1815 454
rect 1819 450 1855 454
rect 1859 450 1871 454
rect 1875 450 1927 454
rect 1931 450 1943 454
rect 1947 450 1999 454
rect 2003 450 2031 454
rect 2035 450 2087 454
rect 2091 450 2111 454
rect 2115 450 2191 454
rect 2195 450 2271 454
rect 2275 450 2311 454
rect 2315 450 2343 454
rect 2347 450 2415 454
rect 2419 450 2439 454
rect 2443 450 2487 454
rect 2491 450 2543 454
rect 2547 450 2583 454
rect 2587 450 2618 454
rect 1345 449 2618 450
rect 1350 398 2630 399
rect 1350 395 1367 398
rect 96 389 97 395
rect 103 394 1351 395
rect 103 390 111 394
rect 115 390 415 394
rect 419 390 439 394
rect 443 390 471 394
rect 475 390 495 394
rect 499 390 535 394
rect 539 390 559 394
rect 563 390 607 394
rect 611 390 631 394
rect 635 390 687 394
rect 691 390 711 394
rect 715 390 767 394
rect 771 390 783 394
rect 787 390 847 394
rect 851 390 855 394
rect 859 390 927 394
rect 931 390 999 394
rect 1003 390 1007 394
rect 1011 390 1071 394
rect 1075 390 1087 394
rect 1091 390 1143 394
rect 1147 390 1175 394
rect 1179 390 1223 394
rect 1227 390 1263 394
rect 1267 390 1327 394
rect 1331 390 1351 394
rect 103 389 1351 390
rect 1357 394 1367 395
rect 1371 394 1631 398
rect 1635 394 1655 398
rect 1659 394 1687 398
rect 1691 394 1711 398
rect 1715 394 1743 398
rect 1747 394 1767 398
rect 1771 394 1799 398
rect 1803 394 1823 398
rect 1827 394 1855 398
rect 1859 394 1879 398
rect 1883 394 1911 398
rect 1915 394 1951 398
rect 1955 394 1983 398
rect 1987 394 2039 398
rect 2043 394 2071 398
rect 2075 394 2151 398
rect 2155 394 2175 398
rect 2179 394 2279 398
rect 2283 394 2295 398
rect 2299 394 2415 398
rect 2419 394 2423 398
rect 2427 394 2527 398
rect 2531 394 2583 398
rect 2587 394 2630 398
rect 1357 393 2630 394
rect 1357 389 1358 393
rect 84 329 85 335
rect 91 334 1339 335
rect 91 330 111 334
rect 115 330 431 334
rect 435 330 463 334
rect 467 330 487 334
rect 491 330 519 334
rect 523 330 551 334
rect 555 330 575 334
rect 579 330 623 334
rect 627 330 631 334
rect 635 330 695 334
rect 699 330 703 334
rect 707 330 767 334
rect 771 330 783 334
rect 787 330 847 334
rect 851 330 863 334
rect 867 330 927 334
rect 931 330 943 334
rect 947 330 1015 334
rect 1019 330 1023 334
rect 1027 330 1103 334
rect 1107 330 1111 334
rect 1115 330 1191 334
rect 1195 330 1215 334
rect 1219 330 1279 334
rect 1283 330 1327 334
rect 1331 330 1339 334
rect 91 329 1339 330
rect 1345 334 2618 335
rect 1345 330 1367 334
rect 1371 330 1631 334
rect 1635 330 1671 334
rect 1675 330 1687 334
rect 1691 330 1727 334
rect 1731 330 1743 334
rect 1747 330 1783 334
rect 1787 330 1807 334
rect 1811 330 1839 334
rect 1843 330 1887 334
rect 1891 330 1895 334
rect 1899 330 1967 334
rect 1971 330 2055 334
rect 2059 330 2143 334
rect 2147 330 2167 334
rect 2171 330 2231 334
rect 2235 330 2295 334
rect 2299 330 2311 334
rect 2315 330 2391 334
rect 2395 330 2431 334
rect 2435 330 2479 334
rect 2483 330 2543 334
rect 2547 330 2583 334
rect 2587 330 2618 334
rect 1345 329 2618 330
rect 1350 278 2630 279
rect 1350 275 1367 278
rect 96 269 97 275
rect 103 274 1351 275
rect 103 270 111 274
rect 115 270 287 274
rect 291 270 359 274
rect 363 270 439 274
rect 443 270 447 274
rect 451 270 503 274
rect 507 270 527 274
rect 531 270 559 274
rect 563 270 615 274
rect 619 270 623 274
rect 627 270 679 274
rect 683 270 719 274
rect 723 270 751 274
rect 755 270 823 274
rect 827 270 831 274
rect 835 270 911 274
rect 915 270 927 274
rect 931 270 999 274
rect 1003 270 1031 274
rect 1035 270 1095 274
rect 1099 270 1143 274
rect 1147 270 1199 274
rect 1203 270 1255 274
rect 1259 270 1327 274
rect 1331 270 1351 274
rect 103 269 1351 270
rect 1357 274 1367 275
rect 1371 274 1535 278
rect 1539 274 1607 278
rect 1611 274 1615 278
rect 1619 274 1671 278
rect 1675 274 1687 278
rect 1691 274 1727 278
rect 1731 274 1775 278
rect 1779 274 1791 278
rect 1795 274 1863 278
rect 1867 274 1871 278
rect 1875 274 1951 278
rect 1955 274 2039 278
rect 2043 274 2119 278
rect 2123 274 2127 278
rect 2131 274 2199 278
rect 2203 274 2215 278
rect 2219 274 2271 278
rect 2275 274 2295 278
rect 2299 274 2335 278
rect 2339 274 2375 278
rect 2379 274 2407 278
rect 2411 274 2463 278
rect 2467 274 2471 278
rect 2475 274 2527 278
rect 2531 274 2583 278
rect 2587 274 2630 278
rect 1357 273 2630 274
rect 1357 269 1358 273
rect 1338 222 2618 223
rect 1338 219 1367 222
rect 84 213 85 219
rect 91 218 1339 219
rect 91 214 111 218
rect 115 214 199 218
rect 203 214 271 218
rect 275 214 303 218
rect 307 214 359 218
rect 363 214 375 218
rect 379 214 455 218
rect 459 214 463 218
rect 467 214 543 218
rect 547 214 567 218
rect 571 214 639 218
rect 643 214 679 218
rect 683 214 735 218
rect 739 214 791 218
rect 795 214 839 218
rect 843 214 911 218
rect 915 214 943 218
rect 947 214 1031 218
rect 1035 214 1047 218
rect 1051 214 1151 218
rect 1155 214 1159 218
rect 1163 214 1271 218
rect 1275 214 1327 218
rect 1331 214 1339 218
rect 91 213 1339 214
rect 1345 218 1367 219
rect 1371 218 1415 222
rect 1419 218 1479 222
rect 1483 218 1551 222
rect 1555 218 1559 222
rect 1563 218 1623 222
rect 1627 218 1655 222
rect 1659 218 1703 222
rect 1707 218 1751 222
rect 1755 218 1791 222
rect 1795 218 1855 222
rect 1859 218 1879 222
rect 1883 218 1959 222
rect 1963 218 1967 222
rect 1971 218 2055 222
rect 2059 218 2063 222
rect 2067 218 2135 222
rect 2139 218 2167 222
rect 2171 218 2215 222
rect 2219 218 2263 222
rect 2267 218 2287 222
rect 2291 218 2351 222
rect 2355 218 2359 222
rect 2363 218 2423 222
rect 2427 218 2463 222
rect 2467 218 2487 222
rect 2491 218 2543 222
rect 2547 218 2583 222
rect 2587 218 2618 222
rect 1345 217 2618 218
rect 1345 213 1346 217
rect 1350 145 1351 151
rect 1357 150 2623 151
rect 1357 146 1367 150
rect 1371 146 1399 150
rect 1403 146 1455 150
rect 1459 146 1463 150
rect 1467 146 1511 150
rect 1515 146 1543 150
rect 1547 146 1567 150
rect 1571 146 1631 150
rect 1635 146 1639 150
rect 1643 146 1711 150
rect 1715 146 1735 150
rect 1739 146 1791 150
rect 1795 146 1839 150
rect 1843 146 1871 150
rect 1875 146 1943 150
rect 1947 146 2015 150
rect 2019 146 2047 150
rect 2051 146 2079 150
rect 2083 146 2143 150
rect 2147 146 2151 150
rect 2155 146 2207 150
rect 2211 146 2247 150
rect 2251 146 2271 150
rect 2275 146 2343 150
rect 2347 146 2415 150
rect 2419 146 2447 150
rect 2451 146 2527 150
rect 2531 146 2583 150
rect 2587 146 2623 150
rect 1357 145 2623 146
rect 2629 145 2630 151
rect 96 133 97 139
rect 103 138 1351 139
rect 103 134 111 138
rect 115 134 143 138
rect 147 134 183 138
rect 187 134 199 138
rect 203 134 255 138
rect 259 134 311 138
rect 315 134 343 138
rect 347 134 367 138
rect 371 134 423 138
rect 427 134 447 138
rect 451 134 479 138
rect 483 134 535 138
rect 539 134 551 138
rect 555 134 591 138
rect 595 134 647 138
rect 651 134 663 138
rect 667 134 703 138
rect 707 134 759 138
rect 763 134 775 138
rect 779 134 823 138
rect 827 134 887 138
rect 891 134 895 138
rect 899 134 951 138
rect 955 134 1015 138
rect 1019 134 1079 138
rect 1083 134 1135 138
rect 1139 134 1151 138
rect 1155 134 1215 138
rect 1219 134 1255 138
rect 1259 134 1271 138
rect 1275 134 1327 138
rect 1331 134 1351 138
rect 103 133 1351 134
rect 1357 133 1358 139
rect 1338 89 1339 95
rect 1345 94 2611 95
rect 1345 90 1367 94
rect 1371 90 1415 94
rect 1419 90 1471 94
rect 1475 90 1527 94
rect 1531 90 1583 94
rect 1587 90 1647 94
rect 1651 90 1727 94
rect 1731 90 1807 94
rect 1811 90 1887 94
rect 1891 90 1959 94
rect 1963 90 2031 94
rect 2035 90 2095 94
rect 2099 90 2159 94
rect 2163 90 2223 94
rect 2227 90 2287 94
rect 2291 90 2359 94
rect 2363 90 2431 94
rect 2435 90 2583 94
rect 2587 90 2611 94
rect 1345 89 2611 90
rect 2617 89 2618 95
rect 84 77 85 83
rect 91 82 1339 83
rect 91 78 111 82
rect 115 78 159 82
rect 163 78 215 82
rect 219 78 271 82
rect 275 78 327 82
rect 331 78 383 82
rect 387 78 439 82
rect 443 78 495 82
rect 499 78 551 82
rect 555 78 607 82
rect 611 78 663 82
rect 667 78 719 82
rect 723 78 775 82
rect 779 78 839 82
rect 843 78 903 82
rect 907 78 967 82
rect 971 78 1031 82
rect 1035 78 1095 82
rect 1099 78 1167 82
rect 1171 78 1231 82
rect 1235 78 1287 82
rect 1291 78 1327 82
rect 1331 78 1339 82
rect 91 77 1339 78
rect 1345 77 1346 83
<< m5c >>
rect 85 2637 91 2643
rect 1339 2637 1345 2643
rect 97 2581 103 2587
rect 1351 2581 1357 2587
rect 85 2521 91 2527
rect 1339 2521 1345 2527
rect 1339 2513 1345 2519
rect 2611 2513 2617 2519
rect 97 2461 103 2467
rect 1351 2461 1357 2467
rect 85 2401 91 2407
rect 1339 2401 1345 2407
rect 97 2345 103 2351
rect 1351 2345 1357 2351
rect 85 2285 91 2291
rect 1339 2285 1345 2291
rect 1339 2277 1345 2283
rect 2611 2277 2617 2283
rect 97 2221 103 2227
rect 1351 2221 1357 2227
rect 1351 2209 1357 2215
rect 2623 2209 2629 2215
rect 85 2161 91 2167
rect 1339 2161 1345 2167
rect 1339 2153 1345 2159
rect 2611 2153 2617 2159
rect 97 2097 103 2103
rect 1351 2097 1357 2103
rect 1339 2041 1345 2047
rect 2611 2041 2617 2047
rect 85 2033 91 2039
rect 1339 2033 1345 2039
rect 1351 1985 1357 1991
rect 2623 1985 2629 1991
rect 97 1973 103 1979
rect 1351 1973 1357 1979
rect 1339 1925 1345 1931
rect 2611 1925 2617 1931
rect 85 1917 91 1923
rect 1339 1917 1345 1923
rect 1351 1865 1357 1871
rect 2623 1865 2629 1871
rect 97 1853 103 1859
rect 1351 1853 1357 1859
rect 1339 1809 1345 1815
rect 2611 1809 2617 1815
rect 85 1793 91 1799
rect 1339 1793 1345 1799
rect 1351 1753 1357 1759
rect 2623 1753 2629 1759
rect 97 1733 103 1739
rect 1351 1733 1357 1739
rect 1339 1685 1345 1691
rect 2611 1685 2617 1691
rect 85 1673 91 1679
rect 1339 1673 1345 1679
rect 1351 1617 1357 1623
rect 2623 1617 2629 1623
rect 97 1601 103 1607
rect 1351 1601 1357 1607
rect 1339 1557 1345 1563
rect 2611 1557 2617 1563
rect 85 1545 91 1551
rect 1339 1545 1345 1551
rect 1351 1493 1357 1499
rect 2623 1493 2629 1499
rect 97 1485 103 1491
rect 1351 1485 1357 1491
rect 85 1425 91 1431
rect 1339 1425 1345 1431
rect 97 1369 103 1375
rect 1351 1369 1357 1375
rect 85 1313 91 1319
rect 1339 1313 1345 1319
rect 1339 1305 1345 1311
rect 2611 1305 2617 1311
rect 97 1245 103 1251
rect 1351 1245 1357 1251
rect 85 1185 91 1191
rect 1339 1185 1345 1191
rect 97 1121 103 1127
rect 1351 1121 1357 1127
rect 85 1061 91 1067
rect 1339 1061 1345 1067
rect 97 1001 103 1007
rect 1351 1001 1357 1007
rect 1351 993 1357 999
rect 2623 993 2629 999
rect 85 941 91 947
rect 1339 941 1345 947
rect 1339 929 1345 935
rect 2611 929 2617 935
rect 97 885 103 891
rect 1351 885 1357 891
rect 1351 873 1357 879
rect 2623 873 2629 879
rect 85 821 91 827
rect 1339 821 1345 827
rect 1339 809 1345 815
rect 2611 809 2617 815
rect 97 757 103 763
rect 1351 757 1357 763
rect 1351 749 1357 755
rect 2623 749 2629 755
rect 85 697 91 703
rect 1339 697 1345 703
rect 1339 689 1345 695
rect 2611 689 2617 695
rect 97 633 103 639
rect 1351 633 1357 639
rect 85 573 91 579
rect 1339 573 1345 579
rect 97 509 103 515
rect 1351 509 1357 515
rect 85 449 91 455
rect 1339 449 1345 455
rect 97 389 103 395
rect 1351 389 1357 395
rect 85 329 91 335
rect 1339 329 1345 335
rect 97 269 103 275
rect 1351 269 1357 275
rect 85 213 91 219
rect 1339 213 1345 219
rect 1351 145 1357 151
rect 2623 145 2629 151
rect 97 133 103 139
rect 1351 133 1357 139
rect 1339 89 1345 95
rect 2611 89 2617 95
rect 85 77 91 83
rect 1339 77 1345 83
<< m5 >>
rect 84 2643 92 2664
rect 84 2637 85 2643
rect 91 2637 92 2643
rect 84 2527 92 2637
rect 84 2521 85 2527
rect 91 2521 92 2527
rect 84 2407 92 2521
rect 84 2401 85 2407
rect 91 2401 92 2407
rect 84 2291 92 2401
rect 84 2285 85 2291
rect 91 2285 92 2291
rect 84 2167 92 2285
rect 84 2161 85 2167
rect 91 2161 92 2167
rect 84 2039 92 2161
rect 84 2033 85 2039
rect 91 2033 92 2039
rect 84 1923 92 2033
rect 84 1917 85 1923
rect 91 1917 92 1923
rect 84 1799 92 1917
rect 84 1793 85 1799
rect 91 1793 92 1799
rect 84 1679 92 1793
rect 84 1673 85 1679
rect 91 1673 92 1679
rect 84 1551 92 1673
rect 84 1545 85 1551
rect 91 1545 92 1551
rect 84 1431 92 1545
rect 84 1425 85 1431
rect 91 1425 92 1431
rect 84 1319 92 1425
rect 84 1313 85 1319
rect 91 1313 92 1319
rect 84 1191 92 1313
rect 84 1185 85 1191
rect 91 1185 92 1191
rect 84 1067 92 1185
rect 84 1061 85 1067
rect 91 1061 92 1067
rect 84 947 92 1061
rect 84 941 85 947
rect 91 941 92 947
rect 84 827 92 941
rect 84 821 85 827
rect 91 821 92 827
rect 84 703 92 821
rect 84 697 85 703
rect 91 697 92 703
rect 84 579 92 697
rect 84 573 85 579
rect 91 573 92 579
rect 84 455 92 573
rect 84 449 85 455
rect 91 449 92 455
rect 84 335 92 449
rect 84 329 85 335
rect 91 329 92 335
rect 84 219 92 329
rect 84 213 85 219
rect 91 213 92 219
rect 84 83 92 213
rect 84 77 85 83
rect 91 77 92 83
rect 84 72 92 77
rect 96 2587 104 2664
rect 96 2581 97 2587
rect 103 2581 104 2587
rect 96 2467 104 2581
rect 96 2461 97 2467
rect 103 2461 104 2467
rect 96 2351 104 2461
rect 96 2345 97 2351
rect 103 2345 104 2351
rect 96 2227 104 2345
rect 96 2221 97 2227
rect 103 2221 104 2227
rect 96 2103 104 2221
rect 96 2097 97 2103
rect 103 2097 104 2103
rect 96 1979 104 2097
rect 96 1973 97 1979
rect 103 1973 104 1979
rect 96 1859 104 1973
rect 96 1853 97 1859
rect 103 1853 104 1859
rect 96 1739 104 1853
rect 96 1733 97 1739
rect 103 1733 104 1739
rect 96 1607 104 1733
rect 96 1601 97 1607
rect 103 1601 104 1607
rect 96 1491 104 1601
rect 96 1485 97 1491
rect 103 1485 104 1491
rect 96 1375 104 1485
rect 96 1369 97 1375
rect 103 1369 104 1375
rect 96 1251 104 1369
rect 96 1245 97 1251
rect 103 1245 104 1251
rect 96 1127 104 1245
rect 96 1121 97 1127
rect 103 1121 104 1127
rect 96 1007 104 1121
rect 96 1001 97 1007
rect 103 1001 104 1007
rect 96 891 104 1001
rect 96 885 97 891
rect 103 885 104 891
rect 96 763 104 885
rect 96 757 97 763
rect 103 757 104 763
rect 96 639 104 757
rect 96 633 97 639
rect 103 633 104 639
rect 96 515 104 633
rect 96 509 97 515
rect 103 509 104 515
rect 96 395 104 509
rect 96 389 97 395
rect 103 389 104 395
rect 96 275 104 389
rect 96 269 97 275
rect 103 269 104 275
rect 96 139 104 269
rect 96 133 97 139
rect 103 133 104 139
rect 96 72 104 133
rect 1338 2643 1346 2664
rect 1338 2637 1339 2643
rect 1345 2637 1346 2643
rect 1338 2527 1346 2637
rect 1338 2521 1339 2527
rect 1345 2521 1346 2527
rect 1338 2519 1346 2521
rect 1338 2513 1339 2519
rect 1345 2513 1346 2519
rect 1338 2407 1346 2513
rect 1338 2401 1339 2407
rect 1345 2401 1346 2407
rect 1338 2291 1346 2401
rect 1338 2285 1339 2291
rect 1345 2285 1346 2291
rect 1338 2283 1346 2285
rect 1338 2277 1339 2283
rect 1345 2277 1346 2283
rect 1338 2167 1346 2277
rect 1338 2161 1339 2167
rect 1345 2161 1346 2167
rect 1338 2159 1346 2161
rect 1338 2153 1339 2159
rect 1345 2153 1346 2159
rect 1338 2047 1346 2153
rect 1338 2041 1339 2047
rect 1345 2041 1346 2047
rect 1338 2039 1346 2041
rect 1338 2033 1339 2039
rect 1345 2033 1346 2039
rect 1338 1931 1346 2033
rect 1338 1925 1339 1931
rect 1345 1925 1346 1931
rect 1338 1923 1346 1925
rect 1338 1917 1339 1923
rect 1345 1917 1346 1923
rect 1338 1815 1346 1917
rect 1338 1809 1339 1815
rect 1345 1809 1346 1815
rect 1338 1799 1346 1809
rect 1338 1793 1339 1799
rect 1345 1793 1346 1799
rect 1338 1691 1346 1793
rect 1338 1685 1339 1691
rect 1345 1685 1346 1691
rect 1338 1679 1346 1685
rect 1338 1673 1339 1679
rect 1345 1673 1346 1679
rect 1338 1563 1346 1673
rect 1338 1557 1339 1563
rect 1345 1557 1346 1563
rect 1338 1551 1346 1557
rect 1338 1545 1339 1551
rect 1345 1545 1346 1551
rect 1338 1431 1346 1545
rect 1338 1425 1339 1431
rect 1345 1425 1346 1431
rect 1338 1319 1346 1425
rect 1338 1313 1339 1319
rect 1345 1313 1346 1319
rect 1338 1311 1346 1313
rect 1338 1305 1339 1311
rect 1345 1305 1346 1311
rect 1338 1191 1346 1305
rect 1338 1185 1339 1191
rect 1345 1185 1346 1191
rect 1338 1067 1346 1185
rect 1338 1061 1339 1067
rect 1345 1061 1346 1067
rect 1338 947 1346 1061
rect 1338 941 1339 947
rect 1345 941 1346 947
rect 1338 935 1346 941
rect 1338 929 1339 935
rect 1345 929 1346 935
rect 1338 827 1346 929
rect 1338 821 1339 827
rect 1345 821 1346 827
rect 1338 815 1346 821
rect 1338 809 1339 815
rect 1345 809 1346 815
rect 1338 703 1346 809
rect 1338 697 1339 703
rect 1345 697 1346 703
rect 1338 695 1346 697
rect 1338 689 1339 695
rect 1345 689 1346 695
rect 1338 579 1346 689
rect 1338 573 1339 579
rect 1345 573 1346 579
rect 1338 455 1346 573
rect 1338 449 1339 455
rect 1345 449 1346 455
rect 1338 335 1346 449
rect 1338 329 1339 335
rect 1345 329 1346 335
rect 1338 219 1346 329
rect 1338 213 1339 219
rect 1345 213 1346 219
rect 1338 95 1346 213
rect 1338 89 1339 95
rect 1345 89 1346 95
rect 1338 83 1346 89
rect 1338 77 1339 83
rect 1345 77 1346 83
rect 1338 72 1346 77
rect 1350 2587 1358 2664
rect 1350 2581 1351 2587
rect 1357 2581 1358 2587
rect 1350 2467 1358 2581
rect 1350 2461 1351 2467
rect 1357 2461 1358 2467
rect 1350 2351 1358 2461
rect 1350 2345 1351 2351
rect 1357 2345 1358 2351
rect 1350 2227 1358 2345
rect 1350 2221 1351 2227
rect 1357 2221 1358 2227
rect 1350 2215 1358 2221
rect 1350 2209 1351 2215
rect 1357 2209 1358 2215
rect 1350 2103 1358 2209
rect 1350 2097 1351 2103
rect 1357 2097 1358 2103
rect 1350 1991 1358 2097
rect 1350 1985 1351 1991
rect 1357 1985 1358 1991
rect 1350 1979 1358 1985
rect 1350 1973 1351 1979
rect 1357 1973 1358 1979
rect 1350 1871 1358 1973
rect 1350 1865 1351 1871
rect 1357 1865 1358 1871
rect 1350 1859 1358 1865
rect 1350 1853 1351 1859
rect 1357 1853 1358 1859
rect 1350 1759 1358 1853
rect 1350 1753 1351 1759
rect 1357 1753 1358 1759
rect 1350 1739 1358 1753
rect 1350 1733 1351 1739
rect 1357 1733 1358 1739
rect 1350 1623 1358 1733
rect 1350 1617 1351 1623
rect 1357 1617 1358 1623
rect 1350 1607 1358 1617
rect 1350 1601 1351 1607
rect 1357 1601 1358 1607
rect 1350 1499 1358 1601
rect 1350 1493 1351 1499
rect 1357 1493 1358 1499
rect 1350 1491 1358 1493
rect 1350 1485 1351 1491
rect 1357 1485 1358 1491
rect 1350 1375 1358 1485
rect 1350 1369 1351 1375
rect 1357 1369 1358 1375
rect 1350 1251 1358 1369
rect 1350 1245 1351 1251
rect 1357 1245 1358 1251
rect 1350 1127 1358 1245
rect 1350 1121 1351 1127
rect 1357 1121 1358 1127
rect 1350 1007 1358 1121
rect 1350 1001 1351 1007
rect 1357 1001 1358 1007
rect 1350 999 1358 1001
rect 1350 993 1351 999
rect 1357 993 1358 999
rect 1350 891 1358 993
rect 1350 885 1351 891
rect 1357 885 1358 891
rect 1350 879 1358 885
rect 1350 873 1351 879
rect 1357 873 1358 879
rect 1350 763 1358 873
rect 1350 757 1351 763
rect 1357 757 1358 763
rect 1350 755 1358 757
rect 1350 749 1351 755
rect 1357 749 1358 755
rect 1350 639 1358 749
rect 1350 633 1351 639
rect 1357 633 1358 639
rect 1350 515 1358 633
rect 1350 509 1351 515
rect 1357 509 1358 515
rect 1350 395 1358 509
rect 1350 389 1351 395
rect 1357 389 1358 395
rect 1350 275 1358 389
rect 1350 269 1351 275
rect 1357 269 1358 275
rect 1350 151 1358 269
rect 1350 145 1351 151
rect 1357 145 1358 151
rect 1350 139 1358 145
rect 1350 133 1351 139
rect 1357 133 1358 139
rect 1350 72 1358 133
rect 2610 2519 2618 2664
rect 2610 2513 2611 2519
rect 2617 2513 2618 2519
rect 2610 2283 2618 2513
rect 2610 2277 2611 2283
rect 2617 2277 2618 2283
rect 2610 2159 2618 2277
rect 2610 2153 2611 2159
rect 2617 2153 2618 2159
rect 2610 2047 2618 2153
rect 2610 2041 2611 2047
rect 2617 2041 2618 2047
rect 2610 1931 2618 2041
rect 2610 1925 2611 1931
rect 2617 1925 2618 1931
rect 2610 1815 2618 1925
rect 2610 1809 2611 1815
rect 2617 1809 2618 1815
rect 2610 1691 2618 1809
rect 2610 1685 2611 1691
rect 2617 1685 2618 1691
rect 2610 1563 2618 1685
rect 2610 1557 2611 1563
rect 2617 1557 2618 1563
rect 2610 1311 2618 1557
rect 2610 1305 2611 1311
rect 2617 1305 2618 1311
rect 2610 935 2618 1305
rect 2610 929 2611 935
rect 2617 929 2618 935
rect 2610 815 2618 929
rect 2610 809 2611 815
rect 2617 809 2618 815
rect 2610 695 2618 809
rect 2610 689 2611 695
rect 2617 689 2618 695
rect 2610 95 2618 689
rect 2610 89 2611 95
rect 2617 89 2618 95
rect 2610 72 2618 89
rect 2622 2215 2630 2664
rect 2622 2209 2623 2215
rect 2629 2209 2630 2215
rect 2622 1991 2630 2209
rect 2622 1985 2623 1991
rect 2629 1985 2630 1991
rect 2622 1871 2630 1985
rect 2622 1865 2623 1871
rect 2629 1865 2630 1871
rect 2622 1759 2630 1865
rect 2622 1753 2623 1759
rect 2629 1753 2630 1759
rect 2622 1623 2630 1753
rect 2622 1617 2623 1623
rect 2629 1617 2630 1623
rect 2622 1499 2630 1617
rect 2622 1493 2623 1499
rect 2629 1493 2630 1499
rect 2622 999 2630 1493
rect 2622 993 2623 999
rect 2629 993 2630 999
rect 2622 879 2630 993
rect 2622 873 2623 879
rect 2629 873 2630 879
rect 2622 755 2630 873
rect 2622 749 2623 755
rect 2629 749 2630 755
rect 2622 151 2630 749
rect 2622 145 2623 151
rect 2629 145 2630 151
rect 2622 72 2630 145
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__167
timestamp 1731220380
transform 1 0 2576 0 -1 2620
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220380
transform 1 0 1360 0 -1 2620
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220380
transform 1 0 2576 0 1 2540
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220380
transform 1 0 1360 0 1 2540
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220380
transform 1 0 2576 0 -1 2500
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220380
transform 1 0 1360 0 -1 2500
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220380
transform 1 0 2576 0 1 2420
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220380
transform 1 0 1360 0 1 2420
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220380
transform 1 0 2576 0 -1 2384
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220380
transform 1 0 1360 0 -1 2384
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220380
transform 1 0 2576 0 1 2304
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220380
transform 1 0 1360 0 1 2304
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220380
transform 1 0 2576 0 -1 2264
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220380
transform 1 0 1360 0 -1 2264
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220380
transform 1 0 2576 0 1 2172
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220380
transform 1 0 1360 0 1 2172
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220380
transform 1 0 2576 0 -1 2140
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220380
transform 1 0 1360 0 -1 2140
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220380
transform 1 0 2576 0 1 2060
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220380
transform 1 0 1360 0 1 2060
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220380
transform 1 0 2576 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220380
transform 1 0 1360 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220380
transform 1 0 2576 0 1 1948
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220380
transform 1 0 1360 0 1 1948
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220380
transform 1 0 2576 0 -1 1912
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220380
transform 1 0 1360 0 -1 1912
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220380
transform 1 0 2576 0 1 1828
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220380
transform 1 0 1360 0 1 1828
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220380
transform 1 0 2576 0 -1 1796
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220380
transform 1 0 1360 0 -1 1796
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220380
transform 1 0 2576 0 1 1716
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220380
transform 1 0 1360 0 1 1716
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220380
transform 1 0 2576 0 -1 1672
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220380
transform 1 0 1360 0 -1 1672
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220380
transform 1 0 2576 0 1 1580
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220380
transform 1 0 1360 0 1 1580
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220380
transform 1 0 2576 0 -1 1544
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220380
transform 1 0 1360 0 -1 1544
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220380
transform 1 0 2576 0 1 1456
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220380
transform 1 0 1360 0 1 1456
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220380
transform 1 0 2576 0 -1 1416
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220380
transform 1 0 1360 0 -1 1416
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220380
transform 1 0 2576 0 1 1328
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220380
transform 1 0 1360 0 1 1328
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220380
transform 1 0 2576 0 -1 1292
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220380
transform 1 0 1360 0 -1 1292
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220380
transform 1 0 2576 0 1 1212
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220380
transform 1 0 1360 0 1 1212
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220380
transform 1 0 2576 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220380
transform 1 0 1360 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220380
transform 1 0 2576 0 1 1088
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220380
transform 1 0 1360 0 1 1088
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220380
transform 1 0 2576 0 -1 1052
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220380
transform 1 0 1360 0 -1 1052
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220380
transform 1 0 2576 0 1 956
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220380
transform 1 0 1360 0 1 956
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220380
transform 1 0 2576 0 -1 916
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220380
transform 1 0 1360 0 -1 916
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220380
transform 1 0 2576 0 1 836
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220380
transform 1 0 1360 0 1 836
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220380
transform 1 0 2576 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220380
transform 1 0 1360 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220380
transform 1 0 2576 0 1 712
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220380
transform 1 0 1360 0 1 712
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220380
transform 1 0 2576 0 -1 676
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220380
transform 1 0 1360 0 -1 676
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220380
transform 1 0 2576 0 1 596
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220380
transform 1 0 1360 0 1 596
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220380
transform 1 0 2576 0 -1 556
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220380
transform 1 0 1360 0 -1 556
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220380
transform 1 0 2576 0 1 476
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220380
transform 1 0 1360 0 1 476
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220380
transform 1 0 2576 0 -1 436
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220380
transform 1 0 1360 0 -1 436
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220380
transform 1 0 2576 0 1 356
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220380
transform 1 0 1360 0 1 356
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220380
transform 1 0 2576 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220380
transform 1 0 1360 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220380
transform 1 0 2576 0 1 236
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220380
transform 1 0 1360 0 1 236
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220380
transform 1 0 2576 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220380
transform 1 0 1360 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220380
transform 1 0 2576 0 1 108
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220380
transform 1 0 1360 0 1 108
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220380
transform 1 0 1320 0 -1 2624
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220380
transform 1 0 104 0 -1 2624
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220380
transform 1 0 1320 0 1 2544
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220380
transform 1 0 104 0 1 2544
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220380
transform 1 0 1320 0 -1 2508
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220380
transform 1 0 104 0 -1 2508
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220380
transform 1 0 1320 0 1 2424
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220380
transform 1 0 104 0 1 2424
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220380
transform 1 0 1320 0 -1 2388
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220380
transform 1 0 104 0 -1 2388
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220380
transform 1 0 1320 0 1 2308
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220380
transform 1 0 104 0 1 2308
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220380
transform 1 0 1320 0 -1 2272
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220380
transform 1 0 104 0 -1 2272
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220380
transform 1 0 1320 0 1 2184
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220380
transform 1 0 104 0 1 2184
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220380
transform 1 0 1320 0 -1 2148
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220380
transform 1 0 104 0 -1 2148
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220380
transform 1 0 1320 0 1 2060
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220380
transform 1 0 104 0 1 2060
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220380
transform 1 0 1320 0 -1 2020
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220380
transform 1 0 104 0 -1 2020
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220380
transform 1 0 1320 0 1 1936
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220380
transform 1 0 104 0 1 1936
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220380
transform 1 0 1320 0 -1 1904
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220380
transform 1 0 104 0 -1 1904
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220380
transform 1 0 1320 0 1 1816
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220380
transform 1 0 104 0 1 1816
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220380
transform 1 0 1320 0 -1 1780
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220380
transform 1 0 104 0 -1 1780
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220380
transform 1 0 1320 0 1 1696
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220380
transform 1 0 104 0 1 1696
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220380
transform 1 0 1320 0 -1 1660
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220380
transform 1 0 104 0 -1 1660
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220380
transform 1 0 1320 0 1 1564
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220380
transform 1 0 104 0 1 1564
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220380
transform 1 0 1320 0 -1 1532
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220380
transform 1 0 104 0 -1 1532
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220380
transform 1 0 1320 0 1 1448
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220380
transform 1 0 104 0 1 1448
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220380
transform 1 0 1320 0 -1 1412
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220380
transform 1 0 104 0 -1 1412
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220380
transform 1 0 1320 0 1 1332
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220380
transform 1 0 104 0 1 1332
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220380
transform 1 0 1320 0 -1 1300
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220380
transform 1 0 104 0 -1 1300
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220380
transform 1 0 1320 0 1 1208
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220380
transform 1 0 104 0 1 1208
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220380
transform 1 0 1320 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220380
transform 1 0 104 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220380
transform 1 0 1320 0 1 1084
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220380
transform 1 0 104 0 1 1084
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220380
transform 1 0 1320 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220380
transform 1 0 104 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220380
transform 1 0 1320 0 1 964
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220380
transform 1 0 104 0 1 964
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220380
transform 1 0 1320 0 -1 928
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220380
transform 1 0 104 0 -1 928
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220380
transform 1 0 1320 0 1 848
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220380
transform 1 0 104 0 1 848
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220380
transform 1 0 1320 0 -1 808
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220380
transform 1 0 104 0 -1 808
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220380
transform 1 0 1320 0 1 720
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220380
transform 1 0 104 0 1 720
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220380
transform 1 0 1320 0 -1 684
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220380
transform 1 0 104 0 -1 684
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220380
transform 1 0 1320 0 1 596
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220380
transform 1 0 104 0 1 596
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220380
transform 1 0 1320 0 -1 560
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220380
transform 1 0 104 0 -1 560
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220380
transform 1 0 1320 0 1 472
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220380
transform 1 0 104 0 1 472
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220380
transform 1 0 1320 0 -1 436
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220380
transform 1 0 104 0 -1 436
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220380
transform 1 0 1320 0 1 352
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220380
transform 1 0 104 0 1 352
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220380
transform 1 0 1320 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220380
transform 1 0 104 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220380
transform 1 0 1320 0 1 232
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220380
transform 1 0 104 0 1 232
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220380
transform 1 0 1320 0 -1 200
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220380
transform 1 0 104 0 -1 200
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220380
transform 1 0 1320 0 1 96
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220380
transform 1 0 104 0 1 96
box 7 3 12 24
use _0_0std_0_0cells_0_0AND2X1  tst_5999_6
timestamp 1731220380
transform 1 0 2440 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5998_6
timestamp 1731220380
transform 1 0 2512 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5997_6
timestamp 1731220380
transform 1 0 2512 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5996_6
timestamp 1731220380
transform 1 0 2512 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5995_6
timestamp 1731220380
transform 1 0 2512 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5994_6
timestamp 1731220380
transform 1 0 2456 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5993_6
timestamp 1731220380
transform 1 0 2304 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5992_6
timestamp 1731220380
transform 1 0 2224 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5991_6
timestamp 1731220380
transform 1 0 2136 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5990_6
timestamp 1731220380
transform 1 0 2040 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5989_6
timestamp 1731220380
transform 1 0 1936 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5988_6
timestamp 1731220380
transform 1 0 2368 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5987_6
timestamp 1731220380
transform 1 0 2304 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5986_6
timestamp 1731220380
transform 1 0 2200 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5985_6
timestamp 1731220380
transform 1 0 2248 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5984_6
timestamp 1731220380
transform 1 0 2160 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5983_6
timestamp 1731220380
transform 1 0 2064 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5982_6
timestamp 1731220380
transform 1 0 1968 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5981_6
timestamp 1731220380
transform 1 0 2152 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5980_6
timestamp 1731220380
transform 1 0 2064 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5979_6
timestamp 1731220380
transform 1 0 1976 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5978_6
timestamp 1731220380
transform 1 0 1912 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5977_6
timestamp 1731220380
transform 1 0 2008 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5976_6
timestamp 1731220380
transform 1 0 2104 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5975_6
timestamp 1731220380
transform 1 0 2208 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5974_6
timestamp 1731220380
transform 1 0 2064 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5973_6
timestamp 1731220380
transform 1 0 1928 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5972_6
timestamp 1731220380
transform 1 0 1808 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5971_6
timestamp 1731220380
transform 1 0 1824 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5970_6
timestamp 1731220380
transform 1 0 1728 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5969_6
timestamp 1731220380
transform 1 0 1632 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5968_6
timestamp 1731220380
transform 1 0 1528 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5967_6
timestamp 1731220380
transform 1 0 1896 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5966_6
timestamp 1731220380
transform 1 0 1824 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5965_6
timestamp 1731220380
transform 1 0 1752 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5964_6
timestamp 1731220380
transform 1 0 1688 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5963_6
timestamp 1731220380
transform 1 0 1632 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5962_6
timestamp 1731220380
transform 1 0 1872 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5961_6
timestamp 1731220380
transform 1 0 1776 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5960_6
timestamp 1731220380
transform 1 0 1688 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5959_6
timestamp 1731220380
transform 1 0 1600 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5958_6
timestamp 1731220380
transform 1 0 1520 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5957_6
timestamp 1731220380
transform 1 0 1864 0 1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5956_6
timestamp 1731220380
transform 1 0 1752 0 1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5955_6
timestamp 1731220380
transform 1 0 1640 0 1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5954_6
timestamp 1731220380
transform 1 0 1528 0 1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5953_6
timestamp 1731220380
transform 1 0 1424 0 1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5952_6
timestamp 1731220380
transform 1 0 1520 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5951_6
timestamp 1731220380
transform 1 0 1576 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5950_6
timestamp 1731220380
transform 1 0 1632 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5949_6
timestamp 1731220380
transform 1 0 1688 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5948_6
timestamp 1731220380
transform 1 0 1744 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5947_6
timestamp 1731220380
transform 1 0 1800 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5946_6
timestamp 1731220380
transform 1 0 1856 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5945_6
timestamp 1731220380
transform 1 0 1912 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5944_6
timestamp 1731220380
transform 1 0 1968 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5943_6
timestamp 1731220380
transform 1 0 2136 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5942_6
timestamp 1731220380
transform 1 0 2080 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5941_6
timestamp 1731220380
transform 1 0 2024 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5940_6
timestamp 1731220380
transform 1 0 1976 0 1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5939_6
timestamp 1731220380
transform 1 0 2096 0 1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5938_6
timestamp 1731220380
transform 1 0 2216 0 1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5937_6
timestamp 1731220380
transform 1 0 2336 0 1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5936_6
timestamp 1731220380
transform 1 0 2264 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5935_6
timestamp 1731220380
transform 1 0 2368 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5934_6
timestamp 1731220380
transform 1 0 2344 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5933_6
timestamp 1731220380
transform 1 0 2416 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5932_6
timestamp 1731220380
transform 1 0 2376 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5931_6
timestamp 1731220380
transform 1 0 2408 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5930_6
timestamp 1731220380
transform 1 0 2512 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5929_6
timestamp 1731220380
transform 1 0 2512 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5928_6
timestamp 1731220380
transform 1 0 2512 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5927_6
timestamp 1731220380
transform 1 0 2512 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5926_6
timestamp 1731220380
transform 1 0 2416 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5925_6
timestamp 1731220380
transform 1 0 2344 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5924_6
timestamp 1731220380
transform 1 0 2440 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5923_6
timestamp 1731220380
transform 1 0 2432 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5922_6
timestamp 1731220380
transform 1 0 2328 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5921_6
timestamp 1731220380
transform 1 0 2296 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5920_6
timestamp 1731220380
transform 1 0 2192 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5919_6
timestamp 1731220380
transform 1 0 2080 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5918_6
timestamp 1731220380
transform 1 0 2024 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5917_6
timestamp 1731220380
transform 1 0 2128 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5916_6
timestamp 1731220380
transform 1 0 2232 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5915_6
timestamp 1731220380
transform 1 0 2256 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5914_6
timestamp 1731220380
transform 1 0 2160 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5913_6
timestamp 1731220380
transform 1 0 2056 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5912_6
timestamp 1731220380
transform 1 0 1952 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5911_6
timestamp 1731220380
transform 1 0 2296 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5910_6
timestamp 1731220380
transform 1 0 2184 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5909_6
timestamp 1731220380
transform 1 0 2080 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5908_6
timestamp 1731220380
transform 1 0 1976 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5907_6
timestamp 1731220380
transform 1 0 1872 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5906_6
timestamp 1731220380
transform 1 0 2072 0 1 1932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5905_6
timestamp 1731220380
transform 1 0 1992 0 1 1932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5904_6
timestamp 1731220380
transform 1 0 1912 0 1 1932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5903_6
timestamp 1731220380
transform 1 0 1832 0 1 1932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5902_6
timestamp 1731220380
transform 1 0 1800 0 -1 1928
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5901_6
timestamp 1731220380
transform 1 0 1856 0 -1 1928
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5900_6
timestamp 1731220380
transform 1 0 1912 0 -1 1928
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5899_6
timestamp 1731220380
transform 1 0 1968 0 -1 1928
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5898_6
timestamp 1731220380
transform 1 0 2088 0 -1 1928
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5897_6
timestamp 1731220380
transform 1 0 2024 0 -1 1928
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5896_6
timestamp 1731220380
transform 1 0 1992 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5895_6
timestamp 1731220380
transform 1 0 1904 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5894_6
timestamp 1731220380
transform 1 0 1816 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5893_6
timestamp 1731220380
transform 1 0 2168 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5892_6
timestamp 1731220380
transform 1 0 2080 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5891_6
timestamp 1731220380
transform 1 0 2032 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5890_6
timestamp 1731220380
transform 1 0 1920 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5889_6
timestamp 1731220380
transform 1 0 2400 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5888_6
timestamp 1731220380
transform 1 0 2272 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5887_6
timestamp 1731220380
transform 1 0 2152 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5886_6
timestamp 1731220380
transform 1 0 2104 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5885_6
timestamp 1731220380
transform 1 0 2008 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5884_6
timestamp 1731220380
transform 1 0 2360 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5883_6
timestamp 1731220380
transform 1 0 2272 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5882_6
timestamp 1731220380
transform 1 0 2192 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5881_6
timestamp 1731220380
transform 1 0 2184 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5880_6
timestamp 1731220380
transform 1 0 2112 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5879_6
timestamp 1731220380
transform 1 0 2032 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5878_6
timestamp 1731220380
transform 1 0 2256 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5877_6
timestamp 1731220380
transform 1 0 2320 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5876_6
timestamp 1731220380
transform 1 0 2392 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5875_6
timestamp 1731220380
transform 1 0 2456 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5874_6
timestamp 1731220380
transform 1 0 2448 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5873_6
timestamp 1731220380
transform 1 0 2512 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5872_6
timestamp 1731220380
transform 1 0 2512 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5871_6
timestamp 1731220380
transform 1 0 2512 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5870_6
timestamp 1731220380
transform 1 0 2512 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5869_6
timestamp 1731220380
transform 1 0 2512 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5868_6
timestamp 1731220380
transform 1 0 2512 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5867_6
timestamp 1731220380
transform 1 0 2456 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5866_6
timestamp 1731220380
transform 1 0 2512 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5865_6
timestamp 1731220380
transform 1 0 2448 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5864_6
timestamp 1731220380
transform 1 0 2360 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5863_6
timestamp 1731220380
transform 1 0 2272 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5862_6
timestamp 1731220380
transform 1 0 2296 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5861_6
timestamp 1731220380
transform 1 0 2376 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5860_6
timestamp 1731220380
transform 1 0 2376 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5859_6
timestamp 1731220380
transform 1 0 2456 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5858_6
timestamp 1731220380
transform 1 0 2416 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5857_6
timestamp 1731220380
transform 1 0 2304 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5856_6
timestamp 1731220380
transform 1 0 2192 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5855_6
timestamp 1731220380
transform 1 0 2136 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5854_6
timestamp 1731220380
transform 1 0 2216 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5853_6
timestamp 1731220380
transform 1 0 2296 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5852_6
timestamp 1731220380
transform 1 0 2216 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5851_6
timestamp 1731220380
transform 1 0 2136 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5850_6
timestamp 1731220380
transform 1 0 2056 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5849_6
timestamp 1731220380
transform 1 0 1992 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5848_6
timestamp 1731220380
transform 1 0 2088 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5847_6
timestamp 1731220380
transform 1 0 2184 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5846_6
timestamp 1731220380
transform 1 0 2192 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5845_6
timestamp 1731220380
transform 1 0 2112 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5844_6
timestamp 1731220380
transform 1 0 2032 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5843_6
timestamp 1731220380
transform 1 0 1952 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5842_6
timestamp 1731220380
transform 1 0 1928 0 -1 1308
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5841_6
timestamp 1731220380
transform 1 0 2016 0 -1 1308
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5840_6
timestamp 1731220380
transform 1 0 2104 0 -1 1308
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5839_6
timestamp 1731220380
transform 1 0 2200 0 -1 1308
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5838_6
timestamp 1731220380
transform 1 0 2136 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5837_6
timestamp 1731220380
transform 1 0 2064 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5836_6
timestamp 1731220380
transform 1 0 2280 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5835_6
timestamp 1731220380
transform 1 0 2208 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5834_6
timestamp 1731220380
transform 1 0 2176 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5833_6
timestamp 1731220380
transform 1 0 2080 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5832_6
timestamp 1731220380
transform 1 0 2368 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5831_6
timestamp 1731220380
transform 1 0 2272 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5830_6
timestamp 1731220380
transform 1 0 2264 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5829_6
timestamp 1731220380
transform 1 0 2200 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5828_6
timestamp 1731220380
transform 1 0 2128 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5827_6
timestamp 1731220380
transform 1 0 2048 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5826_6
timestamp 1731220380
transform 1 0 2136 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5825_6
timestamp 1731220380
transform 1 0 2240 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5824_6
timestamp 1731220380
transform 1 0 2336 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5823_6
timestamp 1731220380
transform 1 0 2328 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5822_6
timestamp 1731220380
transform 1 0 2392 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5821_6
timestamp 1731220380
transform 1 0 2512 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5820_6
timestamp 1731220380
transform 1 0 2456 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5819_6
timestamp 1731220380
transform 1 0 2432 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5818_6
timestamp 1731220380
transform 1 0 2512 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5817_6
timestamp 1731220380
transform 1 0 2512 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5816_6
timestamp 1731220380
transform 1 0 2392 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5815_6
timestamp 1731220380
transform 1 0 2280 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5814_6
timestamp 1731220380
transform 1 0 2408 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5813_6
timestamp 1731220380
transform 1 0 2512 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5812_6
timestamp 1731220380
transform 1 0 2512 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5811_6
timestamp 1731220380
transform 1 0 2456 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5810_6
timestamp 1731220380
transform 1 0 2392 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5809_6
timestamp 1731220380
transform 1 0 2328 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5808_6
timestamp 1731220380
transform 1 0 2264 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5807_6
timestamp 1731220380
transform 1 0 2200 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5806_6
timestamp 1731220380
transform 1 0 2128 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5805_6
timestamp 1731220380
transform 1 0 2056 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5804_6
timestamp 1731220380
transform 1 0 2392 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5803_6
timestamp 1731220380
transform 1 0 2304 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5802_6
timestamp 1731220380
transform 1 0 2216 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5801_6
timestamp 1731220380
transform 1 0 2128 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5800_6
timestamp 1731220380
transform 1 0 2320 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5799_6
timestamp 1731220380
transform 1 0 2232 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5798_6
timestamp 1731220380
transform 1 0 2144 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5797_6
timestamp 1731220380
transform 1 0 2088 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5796_6
timestamp 1731220380
transform 1 0 2176 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5795_6
timestamp 1731220380
transform 1 0 2264 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5794_6
timestamp 1731220380
transform 1 0 2360 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5793_6
timestamp 1731220380
transform 1 0 2392 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5792_6
timestamp 1731220380
transform 1 0 2264 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5791_6
timestamp 1731220380
transform 1 0 2144 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5790_6
timestamp 1731220380
transform 1 0 2208 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5789_6
timestamp 1731220380
transform 1 0 2288 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5788_6
timestamp 1731220380
transform 1 0 2368 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5787_6
timestamp 1731220380
transform 1 0 2512 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5786_6
timestamp 1731220380
transform 1 0 2448 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5785_6
timestamp 1731220380
transform 1 0 2384 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5784_6
timestamp 1731220380
transform 1 0 2312 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5783_6
timestamp 1731220380
transform 1 0 2240 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5782_6
timestamp 1731220380
transform 1 0 2456 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5781_6
timestamp 1731220380
transform 1 0 2512 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5780_6
timestamp 1731220380
transform 1 0 2512 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5779_6
timestamp 1731220380
transform 1 0 2512 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5778_6
timestamp 1731220380
transform 1 0 2512 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5777_6
timestamp 1731220380
transform 1 0 2448 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5776_6
timestamp 1731220380
transform 1 0 2512 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5775_6
timestamp 1731220380
transform 1 0 2512 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5774_6
timestamp 1731220380
transform 1 0 2432 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5773_6
timestamp 1731220380
transform 1 0 2456 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5772_6
timestamp 1731220380
transform 1 0 2392 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5771_6
timestamp 1731220380
transform 1 0 2360 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5770_6
timestamp 1731220380
transform 1 0 2280 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5769_6
timestamp 1731220380
transform 1 0 2200 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5768_6
timestamp 1731220380
transform 1 0 2320 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5767_6
timestamp 1731220380
transform 1 0 2256 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5766_6
timestamp 1731220380
transform 1 0 2184 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5765_6
timestamp 1731220380
transform 1 0 2104 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5764_6
timestamp 1731220380
transform 1 0 2136 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5763_6
timestamp 1731220380
transform 1 0 2232 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5762_6
timestamp 1731220380
transform 1 0 2328 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5761_6
timestamp 1731220380
transform 1 0 2400 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5760_6
timestamp 1731220380
transform 1 0 2328 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5759_6
timestamp 1731220380
transform 1 0 2256 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5758_6
timestamp 1731220380
transform 1 0 2192 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5757_6
timestamp 1731220380
transform 1 0 2128 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5756_6
timestamp 1731220380
transform 1 0 2064 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5755_6
timestamp 1731220380
transform 1 0 2000 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5754_6
timestamp 1731220380
transform 1 0 1928 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5753_6
timestamp 1731220380
transform 1 0 1856 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5752_6
timestamp 1731220380
transform 1 0 1928 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5751_6
timestamp 1731220380
transform 1 0 2032 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5750_6
timestamp 1731220380
transform 1 0 2024 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5749_6
timestamp 1731220380
transform 1 0 1936 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5748_6
timestamp 1731220380
transform 1 0 2024 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5747_6
timestamp 1731220380
transform 1 0 2112 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5746_6
timestamp 1731220380
transform 1 0 2400 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5745_6
timestamp 1731220380
transform 1 0 2264 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5744_6
timestamp 1731220380
transform 1 0 2136 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5743_6
timestamp 1731220380
transform 1 0 2024 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5742_6
timestamp 1731220380
transform 1 0 1968 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5741_6
timestamp 1731220380
transform 1 0 2056 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5740_6
timestamp 1731220380
transform 1 0 2408 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5739_6
timestamp 1731220380
transform 1 0 2280 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5738_6
timestamp 1731220380
transform 1 0 2160 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5737_6
timestamp 1731220380
transform 1 0 2160 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5736_6
timestamp 1731220380
transform 1 0 2080 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5735_6
timestamp 1731220380
transform 1 0 2000 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5734_6
timestamp 1731220380
transform 1 0 2120 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5733_6
timestamp 1731220380
transform 1 0 2024 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5732_6
timestamp 1731220380
transform 1 0 1928 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5731_6
timestamp 1731220380
transform 1 0 1896 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5730_6
timestamp 1731220380
transform 1 0 2024 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5729_6
timestamp 1731220380
transform 1 0 1992 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5728_6
timestamp 1731220380
transform 1 0 1896 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5727_6
timestamp 1731220380
transform 1 0 1984 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5726_6
timestamp 1731220380
transform 1 0 2064 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5725_6
timestamp 1731220380
transform 1 0 2040 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5724_6
timestamp 1731220380
transform 1 0 1976 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5723_6
timestamp 1731220380
transform 1 0 1888 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5722_6
timestamp 1731220380
transform 1 0 1912 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5721_6
timestamp 1731220380
transform 1 0 2032 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5720_6
timestamp 1731220380
transform 1 0 2152 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5719_6
timestamp 1731220380
transform 1 0 2256 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5718_6
timestamp 1731220380
transform 1 0 2128 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5717_6
timestamp 1731220380
transform 1 0 2000 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5716_6
timestamp 1731220380
transform 1 0 1888 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5715_6
timestamp 1731220380
transform 1 0 1792 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5714_6
timestamp 1731220380
transform 1 0 1920 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5713_6
timestamp 1731220380
transform 1 0 2032 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5712_6
timestamp 1731220380
transform 1 0 1960 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5711_6
timestamp 1731220380
transform 1 0 1872 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5710_6
timestamp 1731220380
transform 1 0 1984 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5709_6
timestamp 1731220380
transform 1 0 2000 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5708_6
timestamp 1731220380
transform 1 0 1936 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5707_6
timestamp 1731220380
transform 1 0 1832 0 -1 1308
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5706_6
timestamp 1731220380
transform 1 0 1792 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5705_6
timestamp 1731220380
transform 1 0 1872 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5704_6
timestamp 1731220380
transform 1 0 1896 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5703_6
timestamp 1731220380
transform 1 0 1968 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5702_6
timestamp 1731220380
transform 1 0 2056 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5701_6
timestamp 1731220380
transform 1 0 2088 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5700_6
timestamp 1731220380
transform 1 0 1992 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5699_6
timestamp 1731220380
transform 1 0 1904 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5698_6
timestamp 1731220380
transform 1 0 1944 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5697_6
timestamp 1731220380
transform 1 0 1856 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5696_6
timestamp 1731220380
transform 1 0 1768 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5695_6
timestamp 1731220380
transform 1 0 1808 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5694_6
timestamp 1731220380
transform 1 0 1912 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5693_6
timestamp 1731220380
transform 1 0 1808 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5692_6
timestamp 1731220380
transform 1 0 1704 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5691_6
timestamp 1731220380
transform 1 0 1728 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5690_6
timestamp 1731220380
transform 1 0 1744 0 -1 1928
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5689_6
timestamp 1731220380
transform 1 0 1688 0 -1 1928
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5688_6
timestamp 1731220380
transform 1 0 1664 0 1 1932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5687_6
timestamp 1731220380
transform 1 0 1568 0 1 1932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5686_6
timestamp 1731220380
transform 1 0 1752 0 1 1932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5685_6
timestamp 1731220380
transform 1 0 1680 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5684_6
timestamp 1731220380
transform 1 0 1776 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5683_6
timestamp 1731220380
transform 1 0 1744 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5682_6
timestamp 1731220380
transform 1 0 1848 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5681_6
timestamp 1731220380
transform 1 0 1808 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5680_6
timestamp 1731220380
transform 1 0 1920 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5679_6
timestamp 1731220380
transform 1 0 1968 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5678_6
timestamp 1731220380
transform 1 0 1848 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5677_6
timestamp 1731220380
transform 1 0 1728 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5676_6
timestamp 1731220380
transform 1 0 1704 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5675_6
timestamp 1731220380
transform 1 0 1824 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5674_6
timestamp 1731220380
transform 1 0 1712 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5673_6
timestamp 1731220380
transform 1 0 1624 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5672_6
timestamp 1731220380
transform 1 0 1552 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5671_6
timestamp 1731220380
transform 1 0 1424 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5670_6
timestamp 1731220380
transform 1 0 1496 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5669_6
timestamp 1731220380
transform 1 0 1440 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5668_6
timestamp 1731220380
transform 1 0 1384 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5667_6
timestamp 1731220380
transform 1 0 1256 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5666_6
timestamp 1731220380
transform 1 0 1384 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5665_6
timestamp 1731220380
transform 1 0 1464 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5664_6
timestamp 1731220380
transform 1 0 1584 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5663_6
timestamp 1731220380
transform 1 0 1616 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5662_6
timestamp 1731220380
transform 1 0 1520 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5661_6
timestamp 1731220380
transform 1 0 1440 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5660_6
timestamp 1731220380
transform 1 0 1504 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5659_6
timestamp 1731220380
transform 1 0 1600 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5658_6
timestamp 1731220380
transform 1 0 1704 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5657_6
timestamp 1731220380
transform 1 0 1632 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5656_6
timestamp 1731220380
transform 1 0 1520 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5655_6
timestamp 1731220380
transform 1 0 1416 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5654_6
timestamp 1731220380
transform 1 0 1384 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5653_6
timestamp 1731220380
transform 1 0 1576 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5652_6
timestamp 1731220380
transform 1 0 1472 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5651_6
timestamp 1731220380
transform 1 0 1464 0 1 1932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5650_6
timestamp 1731220380
transform 1 0 1384 0 1 1932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5649_6
timestamp 1731220380
transform 1 0 1256 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5648_6
timestamp 1731220380
transform 1 0 1168 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5647_6
timestamp 1731220380
transform 1 0 1056 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5646_6
timestamp 1731220380
transform 1 0 1256 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5645_6
timestamp 1731220380
transform 1 0 1384 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5644_6
timestamp 1731220380
transform 1 0 1448 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5643_6
timestamp 1731220380
transform 1 0 1544 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5642_6
timestamp 1731220380
transform 1 0 1640 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5641_6
timestamp 1731220380
transform 1 0 1592 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5640_6
timestamp 1731220380
transform 1 0 1480 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5639_6
timestamp 1731220380
transform 1 0 1384 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5638_6
timestamp 1731220380
transform 1 0 1424 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5637_6
timestamp 1731220380
transform 1 0 1504 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5636_6
timestamp 1731220380
transform 1 0 1600 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5635_6
timestamp 1731220380
transform 1 0 1704 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5634_6
timestamp 1731220380
transform 1 0 1680 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5633_6
timestamp 1731220380
transform 1 0 1600 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5632_6
timestamp 1731220380
transform 1 0 1528 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5631_6
timestamp 1731220380
transform 1 0 1560 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5630_6
timestamp 1731220380
transform 1 0 1616 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5629_6
timestamp 1731220380
transform 1 0 1672 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5628_6
timestamp 1731220380
transform 1 0 1736 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5627_6
timestamp 1731220380
transform 1 0 1816 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5626_6
timestamp 1731220380
transform 1 0 1976 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5625_6
timestamp 1731220380
transform 1 0 1896 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5624_6
timestamp 1731220380
transform 1 0 1824 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5623_6
timestamp 1731220380
transform 1 0 1760 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5622_6
timestamp 1731220380
transform 1 0 1704 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5621_6
timestamp 1731220380
transform 1 0 1648 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5620_6
timestamp 1731220380
transform 1 0 1880 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5619_6
timestamp 1731220380
transform 1 0 1792 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5618_6
timestamp 1731220380
transform 1 0 1712 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5617_6
timestamp 1731220380
transform 1 0 1632 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5616_6
timestamp 1731220380
transform 1 0 1560 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5615_6
timestamp 1731220380
transform 1 0 1504 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5614_6
timestamp 1731220380
transform 1 0 1792 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5613_6
timestamp 1731220380
transform 1 0 1688 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5612_6
timestamp 1731220380
transform 1 0 1592 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5611_6
timestamp 1731220380
transform 1 0 1504 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5610_6
timestamp 1731220380
transform 1 0 1440 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5609_6
timestamp 1731220380
transform 1 0 1384 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5608_6
timestamp 1731220380
transform 1 0 1704 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5607_6
timestamp 1731220380
transform 1 0 1616 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5606_6
timestamp 1731220380
transform 1 0 1528 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5605_6
timestamp 1731220380
transform 1 0 1440 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5604_6
timestamp 1731220380
transform 1 0 1384 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5603_6
timestamp 1731220380
transform 1 0 1256 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5602_6
timestamp 1731220380
transform 1 0 1200 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5601_6
timestamp 1731220380
transform 1 0 1120 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5600_6
timestamp 1731220380
transform 1 0 1040 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5599_6
timestamp 1731220380
transform 1 0 960 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5598_6
timestamp 1731220380
transform 1 0 880 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5597_6
timestamp 1731220380
transform 1 0 1256 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5596_6
timestamp 1731220380
transform 1 0 1168 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5595_6
timestamp 1731220380
transform 1 0 1056 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5594_6
timestamp 1731220380
transform 1 0 944 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5593_6
timestamp 1731220380
transform 1 0 960 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5592_6
timestamp 1731220380
transform 1 0 1072 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5591_6
timestamp 1731220380
transform 1 0 1184 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5590_6
timestamp 1731220380
transform 1 0 1120 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5589_6
timestamp 1731220380
transform 1 0 1024 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5588_6
timestamp 1731220380
transform 1 0 936 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5587_6
timestamp 1731220380
transform 1 0 848 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5586_6
timestamp 1731220380
transform 1 0 872 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5585_6
timestamp 1731220380
transform 1 0 944 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5584_6
timestamp 1731220380
transform 1 0 1024 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5583_6
timestamp 1731220380
transform 1 0 968 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5582_6
timestamp 1731220380
transform 1 0 888 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5581_6
timestamp 1731220380
transform 1 0 1048 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5580_6
timestamp 1731220380
transform 1 0 1136 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5579_6
timestamp 1731220380
transform 1 0 1104 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5578_6
timestamp 1731220380
transform 1 0 1016 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5577_6
timestamp 1731220380
transform 1 0 1256 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5576_6
timestamp 1731220380
transform 1 0 1192 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5575_6
timestamp 1731220380
transform 1 0 1192 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5574_6
timestamp 1731220380
transform 1 0 1096 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5573_6
timestamp 1731220380
transform 1 0 1000 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5572_6
timestamp 1731220380
transform 1 0 1088 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5571_6
timestamp 1731220380
transform 1 0 1000 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5570_6
timestamp 1731220380
transform 1 0 856 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5569_6
timestamp 1731220380
transform 1 0 776 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5568_6
timestamp 1731220380
transform 1 0 696 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5567_6
timestamp 1731220380
transform 1 0 608 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5566_6
timestamp 1731220380
transform 1 0 592 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5565_6
timestamp 1731220380
transform 1 0 760 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5564_6
timestamp 1731220380
transform 1 0 680 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5563_6
timestamp 1731220380
transform 1 0 624 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5562_6
timestamp 1731220380
transform 1 0 712 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5561_6
timestamp 1731220380
transform 1 0 808 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5560_6
timestamp 1731220380
transform 1 0 776 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5559_6
timestamp 1731220380
transform 1 0 696 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5558_6
timestamp 1731220380
transform 1 0 616 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5557_6
timestamp 1731220380
transform 1 0 544 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5556_6
timestamp 1731220380
transform 1 0 480 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5555_6
timestamp 1731220380
transform 1 0 424 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5554_6
timestamp 1731220380
transform 1 0 368 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5553_6
timestamp 1731220380
transform 1 0 536 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5552_6
timestamp 1731220380
transform 1 0 456 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5551_6
timestamp 1731220380
transform 1 0 392 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5550_6
timestamp 1731220380
transform 1 0 336 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5549_6
timestamp 1731220380
transform 1 0 504 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5548_6
timestamp 1731220380
transform 1 0 416 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5547_6
timestamp 1731220380
transform 1 0 336 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5546_6
timestamp 1731220380
transform 1 0 264 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5545_6
timestamp 1731220380
transform 1 0 200 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5544_6
timestamp 1731220380
transform 1 0 520 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5543_6
timestamp 1731220380
transform 1 0 424 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5542_6
timestamp 1731220380
transform 1 0 336 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5541_6
timestamp 1731220380
transform 1 0 248 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5540_6
timestamp 1731220380
transform 1 0 184 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5539_6
timestamp 1731220380
transform 1 0 128 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5538_6
timestamp 1731220380
transform 1 0 128 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5537_6
timestamp 1731220380
transform 1 0 200 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5536_6
timestamp 1731220380
transform 1 0 296 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5535_6
timestamp 1731220380
transform 1 0 400 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5534_6
timestamp 1731220380
transform 1 0 512 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5533_6
timestamp 1731220380
transform 1 0 432 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5532_6
timestamp 1731220380
transform 1 0 376 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5531_6
timestamp 1731220380
transform 1 0 320 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5530_6
timestamp 1731220380
transform 1 0 488 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5529_6
timestamp 1731220380
transform 1 0 552 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5528_6
timestamp 1731220380
transform 1 0 664 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5527_6
timestamp 1731220380
transform 1 0 608 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5526_6
timestamp 1731220380
transform 1 0 552 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5525_6
timestamp 1731220380
transform 1 0 496 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5524_6
timestamp 1731220380
transform 1 0 440 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5523_6
timestamp 1731220380
transform 1 0 384 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5522_6
timestamp 1731220380
transform 1 0 640 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5521_6
timestamp 1731220380
transform 1 0 552 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5520_6
timestamp 1731220380
transform 1 0 464 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5519_6
timestamp 1731220380
transform 1 0 384 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5518_6
timestamp 1731220380
transform 1 0 312 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5517_6
timestamp 1731220380
transform 1 0 248 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5516_6
timestamp 1731220380
transform 1 0 632 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5515_6
timestamp 1731220380
transform 1 0 512 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5514_6
timestamp 1731220380
transform 1 0 392 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5513_6
timestamp 1731220380
transform 1 0 280 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5512_6
timestamp 1731220380
transform 1 0 184 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5511_6
timestamp 1731220380
transform 1 0 128 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5510_6
timestamp 1731220380
transform 1 0 608 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5509_6
timestamp 1731220380
transform 1 0 480 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5508_6
timestamp 1731220380
transform 1 0 344 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5507_6
timestamp 1731220380
transform 1 0 216 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5506_6
timestamp 1731220380
transform 1 0 128 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5505_6
timestamp 1731220380
transform 1 0 128 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5504_6
timestamp 1731220380
transform 1 0 216 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5503_6
timestamp 1731220380
transform 1 0 608 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5502_6
timestamp 1731220380
transform 1 0 480 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5501_6
timestamp 1731220380
transform 1 0 344 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5500_6
timestamp 1731220380
transform 1 0 248 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5499_6
timestamp 1731220380
transform 1 0 144 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5498_6
timestamp 1731220380
transform 1 0 584 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5497_6
timestamp 1731220380
transform 1 0 472 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5496_6
timestamp 1731220380
transform 1 0 360 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5495_6
timestamp 1731220380
transform 1 0 304 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5494_6
timestamp 1731220380
transform 1 0 216 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5493_6
timestamp 1731220380
transform 1 0 600 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5492_6
timestamp 1731220380
transform 1 0 496 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5491_6
timestamp 1731220380
transform 1 0 400 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5490_6
timestamp 1731220380
transform 1 0 384 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5489_6
timestamp 1731220380
transform 1 0 320 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5488_6
timestamp 1731220380
transform 1 0 256 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5487_6
timestamp 1731220380
transform 1 0 456 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5486_6
timestamp 1731220380
transform 1 0 536 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5485_6
timestamp 1731220380
transform 1 0 616 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5484_6
timestamp 1731220380
transform 1 0 584 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5483_6
timestamp 1731220380
transform 1 0 520 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5482_6
timestamp 1731220380
transform 1 0 456 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5481_6
timestamp 1731220380
transform 1 0 392 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5480_6
timestamp 1731220380
transform 1 0 336 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5479_6
timestamp 1731220380
transform 1 0 312 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5478_6
timestamp 1731220380
transform 1 0 256 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5477_6
timestamp 1731220380
transform 1 0 200 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5476_6
timestamp 1731220380
transform 1 0 368 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5475_6
timestamp 1731220380
transform 1 0 424 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5474_6
timestamp 1731220380
transform 1 0 480 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5473_6
timestamp 1731220380
transform 1 0 592 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5472_6
timestamp 1731220380
transform 1 0 536 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5471_6
timestamp 1731220380
transform 1 0 520 0 -1 2640
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5470_6
timestamp 1731220380
transform 1 0 576 0 -1 2640
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5469_6
timestamp 1731220380
transform 1 0 632 0 -1 2640
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5468_6
timestamp 1731220380
transform 1 0 688 0 -1 2640
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5467_6
timestamp 1731220380
transform 1 0 744 0 -1 2640
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5466_6
timestamp 1731220380
transform 1 0 704 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5465_6
timestamp 1731220380
transform 1 0 648 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5464_6
timestamp 1731220380
transform 1 0 760 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5463_6
timestamp 1731220380
transform 1 0 816 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5462_6
timestamp 1731220380
transform 1 0 872 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5461_6
timestamp 1731220380
transform 1 0 928 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5460_6
timestamp 1731220380
transform 1 0 1096 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5459_6
timestamp 1731220380
transform 1 0 1040 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5458_6
timestamp 1731220380
transform 1 0 984 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5457_6
timestamp 1731220380
transform 1 0 776 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5456_6
timestamp 1731220380
transform 1 0 712 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5455_6
timestamp 1731220380
transform 1 0 648 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5454_6
timestamp 1731220380
transform 1 0 840 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5453_6
timestamp 1731220380
transform 1 0 984 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5452_6
timestamp 1731220380
transform 1 0 912 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5451_6
timestamp 1731220380
transform 1 0 848 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5450_6
timestamp 1731220380
transform 1 0 768 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5449_6
timestamp 1731220380
transform 1 0 696 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5448_6
timestamp 1731220380
transform 1 0 1008 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5447_6
timestamp 1731220380
transform 1 0 928 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5446_6
timestamp 1731220380
transform 1 0 888 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5445_6
timestamp 1731220380
transform 1 0 792 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5444_6
timestamp 1731220380
transform 1 0 696 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5443_6
timestamp 1731220380
transform 1 0 1080 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5442_6
timestamp 1731220380
transform 1 0 984 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5441_6
timestamp 1731220380
transform 1 0 896 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5440_6
timestamp 1731220380
transform 1 0 800 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5439_6
timestamp 1731220380
transform 1 0 696 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5438_6
timestamp 1731220380
transform 1 0 1184 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5437_6
timestamp 1731220380
transform 1 0 1088 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5436_6
timestamp 1731220380
transform 1 0 992 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5435_6
timestamp 1731220380
transform 1 0 968 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5434_6
timestamp 1731220380
transform 1 0 856 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5433_6
timestamp 1731220380
transform 1 0 736 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5432_6
timestamp 1731220380
transform 1 0 1072 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5431_6
timestamp 1731220380
transform 1 0 1176 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5430_6
timestamp 1731220380
transform 1 0 1256 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5429_6
timestamp 1731220380
transform 1 0 1176 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5428_6
timestamp 1731220380
transform 1 0 1072 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5427_6
timestamp 1731220380
transform 1 0 968 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5426_6
timestamp 1731220380
transform 1 0 856 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5425_6
timestamp 1731220380
transform 1 0 736 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5424_6
timestamp 1731220380
transform 1 0 1240 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5423_6
timestamp 1731220380
transform 1 0 1136 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5422_6
timestamp 1731220380
transform 1 0 1040 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5421_6
timestamp 1731220380
transform 1 0 944 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5420_6
timestamp 1731220380
transform 1 0 848 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5419_6
timestamp 1731220380
transform 1 0 744 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5418_6
timestamp 1731220380
transform 1 0 1112 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5417_6
timestamp 1731220380
transform 1 0 1032 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5416_6
timestamp 1731220380
transform 1 0 952 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5415_6
timestamp 1731220380
transform 1 0 872 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5414_6
timestamp 1731220380
transform 1 0 800 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5413_6
timestamp 1731220380
transform 1 0 720 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5412_6
timestamp 1731220380
transform 1 0 1000 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5411_6
timestamp 1731220380
transform 1 0 944 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5410_6
timestamp 1731220380
transform 1 0 888 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5409_6
timestamp 1731220380
transform 1 0 832 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5408_6
timestamp 1731220380
transform 1 0 776 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5407_6
timestamp 1731220380
transform 1 0 720 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5406_6
timestamp 1731220380
transform 1 0 1128 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5405_6
timestamp 1731220380
transform 1 0 984 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5404_6
timestamp 1731220380
transform 1 0 848 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5403_6
timestamp 1731220380
transform 1 0 728 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5402_6
timestamp 1731220380
transform 1 0 632 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5401_6
timestamp 1731220380
transform 1 0 624 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5400_6
timestamp 1731220380
transform 1 0 736 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5399_6
timestamp 1731220380
transform 1 0 848 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5398_6
timestamp 1731220380
transform 1 0 952 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5397_6
timestamp 1731220380
transform 1 0 1024 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5396_6
timestamp 1731220380
transform 1 0 936 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5395_6
timestamp 1731220380
transform 1 0 920 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5394_6
timestamp 1731220380
transform 1 0 840 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5393_6
timestamp 1731220380
transform 1 0 904 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5392_6
timestamp 1731220380
transform 1 0 936 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5391_6
timestamp 1731220380
transform 1 0 856 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5390_6
timestamp 1731220380
transform 1 0 808 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5389_6
timestamp 1731220380
transform 1 0 720 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5388_6
timestamp 1731220380
transform 1 0 656 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5387_6
timestamp 1731220380
transform 1 0 728 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5386_6
timestamp 1731220380
transform 1 0 800 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5385_6
timestamp 1731220380
transform 1 0 760 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5384_6
timestamp 1731220380
transform 1 0 664 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5383_6
timestamp 1731220380
transform 1 0 736 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5382_6
timestamp 1731220380
transform 1 0 848 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5381_6
timestamp 1731220380
transform 1 0 832 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5380_6
timestamp 1731220380
transform 1 0 720 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5379_6
timestamp 1731220380
transform 1 0 696 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5378_6
timestamp 1731220380
transform 1 0 600 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5377_6
timestamp 1731220380
transform 1 0 792 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5376_6
timestamp 1731220380
transform 1 0 728 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5375_6
timestamp 1731220380
transform 1 0 656 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5374_6
timestamp 1731220380
transform 1 0 584 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5373_6
timestamp 1731220380
transform 1 0 800 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5372_6
timestamp 1731220380
transform 1 0 880 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5371_6
timestamp 1731220380
transform 1 0 808 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5370_6
timestamp 1731220380
transform 1 0 736 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5369_6
timestamp 1731220380
transform 1 0 656 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5368_6
timestamp 1731220380
transform 1 0 880 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5367_6
timestamp 1731220380
transform 1 0 1032 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5366_6
timestamp 1731220380
transform 1 0 952 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5365_6
timestamp 1731220380
transform 1 0 896 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5364_6
timestamp 1731220380
transform 1 0 808 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5363_6
timestamp 1731220380
transform 1 0 712 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5362_6
timestamp 1731220380
transform 1 0 976 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5361_6
timestamp 1731220380
transform 1 0 1152 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5360_6
timestamp 1731220380
transform 1 0 1064 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5359_6
timestamp 1731220380
transform 1 0 1024 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5358_6
timestamp 1731220380
transform 1 0 944 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5357_6
timestamp 1731220380
transform 1 0 856 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5356_6
timestamp 1731220380
transform 1 0 1192 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5355_6
timestamp 1731220380
transform 1 0 1104 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5354_6
timestamp 1731220380
transform 1 0 896 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5353_6
timestamp 1731220380
transform 1 0 832 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5352_6
timestamp 1731220380
transform 1 0 768 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5351_6
timestamp 1731220380
transform 1 0 960 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5350_6
timestamp 1731220380
transform 1 0 1024 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5349_6
timestamp 1731220380
transform 1 0 1088 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5348_6
timestamp 1731220380
transform 1 0 1144 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5347_6
timestamp 1731220380
transform 1 0 1200 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5346_6
timestamp 1731220380
transform 1 0 1256 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5345_6
timestamp 1731220380
transform 1 0 1256 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5344_6
timestamp 1731220380
transform 1 0 1384 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5343_6
timestamp 1731220380
transform 1 0 1440 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5342_6
timestamp 1731220380
transform 1 0 1464 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5341_6
timestamp 1731220380
transform 1 0 1384 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5340_6
timestamp 1731220380
transform 1 0 1384 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5339_6
timestamp 1731220380
transform 1 0 1472 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5338_6
timestamp 1731220380
transform 1 0 1568 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5337_6
timestamp 1731220380
transform 1 0 1544 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5336_6
timestamp 1731220380
transform 1 0 1480 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5335_6
timestamp 1731220380
transform 1 0 1608 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5334_6
timestamp 1731220380
transform 1 0 1640 0 -1 1308
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5333_6
timestamp 1731220380
transform 1 0 1736 0 -1 1308
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5332_6
timestamp 1731220380
transform 1 0 1744 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5331_6
timestamp 1731220380
transform 1 0 1672 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5330_6
timestamp 1731220380
transform 1 0 1808 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5329_6
timestamp 1731220380
transform 1 0 1872 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5328_6
timestamp 1731220380
transform 1 0 1880 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5327_6
timestamp 1731220380
transform 1 0 1776 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5326_6
timestamp 1731220380
transform 1 0 1672 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5325_6
timestamp 1731220380
transform 1 0 1568 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5324_6
timestamp 1731220380
transform 1 0 1672 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5323_6
timestamp 1731220380
transform 1 0 1776 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5322_6
timestamp 1731220380
transform 1 0 1808 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5321_6
timestamp 1731220380
transform 1 0 1696 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5320_6
timestamp 1731220380
transform 1 0 1592 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5319_6
timestamp 1731220380
transform 1 0 1504 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5318_6
timestamp 1731220380
transform 1 0 1704 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5317_6
timestamp 1731220380
transform 1 0 1624 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5316_6
timestamp 1731220380
transform 1 0 1552 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5315_6
timestamp 1731220380
transform 1 0 1496 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5314_6
timestamp 1731220380
transform 1 0 1440 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5313_6
timestamp 1731220380
transform 1 0 1384 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5312_6
timestamp 1731220380
transform 1 0 1384 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5311_6
timestamp 1731220380
transform 1 0 1440 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5310_6
timestamp 1731220380
transform 1 0 1496 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5309_6
timestamp 1731220380
transform 1 0 1584 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5308_6
timestamp 1731220380
transform 1 0 1792 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5307_6
timestamp 1731220380
transform 1 0 1680 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5306_6
timestamp 1731220380
transform 1 0 1624 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5305_6
timestamp 1731220380
transform 1 0 1536 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5304_6
timestamp 1731220380
transform 1 0 1456 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5303_6
timestamp 1731220380
transform 1 0 1712 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5302_6
timestamp 1731220380
transform 1 0 1800 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5301_6
timestamp 1731220380
transform 1 0 1720 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5300_6
timestamp 1731220380
transform 1 0 1656 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5299_6
timestamp 1731220380
transform 1 0 1600 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5298_6
timestamp 1731220380
transform 1 0 1792 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5297_6
timestamp 1731220380
transform 1 0 1872 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5296_6
timestamp 1731220380
transform 1 0 1960 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5295_6
timestamp 1731220380
transform 1 0 1904 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5294_6
timestamp 1731220380
transform 1 0 1824 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5293_6
timestamp 1731220380
transform 1 0 1744 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5292_6
timestamp 1731220380
transform 1 0 1672 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5291_6
timestamp 1731220380
transform 1 0 1608 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5290_6
timestamp 1731220380
transform 1 0 1552 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5289_6
timestamp 1731220380
transform 1 0 1792 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5288_6
timestamp 1731220380
transform 1 0 1688 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5287_6
timestamp 1731220380
transform 1 0 1584 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5286_6
timestamp 1731220380
transform 1 0 1480 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5285_6
timestamp 1731220380
transform 1 0 1384 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5284_6
timestamp 1731220380
transform 1 0 1768 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5283_6
timestamp 1731220380
transform 1 0 1632 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5282_6
timestamp 1731220380
transform 1 0 1256 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5281_6
timestamp 1731220380
transform 1 0 1176 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5280_6
timestamp 1731220380
transform 1 0 1072 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5279_6
timestamp 1731220380
transform 1 0 976 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5278_6
timestamp 1731220380
transform 1 0 1032 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5277_6
timestamp 1731220380
transform 1 0 1152 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5276_6
timestamp 1731220380
transform 1 0 1256 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5275_6
timestamp 1731220380
transform 1 0 1384 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5274_6
timestamp 1731220380
transform 1 0 1496 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5273_6
timestamp 1731220380
transform 1 0 1440 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5272_6
timestamp 1731220380
transform 1 0 1384 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5271_6
timestamp 1731220380
transform 1 0 1520 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5270_6
timestamp 1731220380
transform 1 0 1616 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5269_6
timestamp 1731220380
transform 1 0 1824 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5268_6
timestamp 1731220380
transform 1 0 1720 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5267_6
timestamp 1731220380
transform 1 0 1656 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5266_6
timestamp 1731220380
transform 1 0 1584 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5265_6
timestamp 1731220380
transform 1 0 1520 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5264_6
timestamp 1731220380
transform 1 0 1912 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5263_6
timestamp 1731220380
transform 1 0 1824 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5262_6
timestamp 1731220380
transform 1 0 1736 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5261_6
timestamp 1731220380
transform 1 0 1728 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5260_6
timestamp 1731220380
transform 1 0 1672 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5259_6
timestamp 1731220380
transform 1 0 1616 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5258_6
timestamp 1731220380
transform 1 0 1784 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5257_6
timestamp 1731220380
transform 1 0 1840 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5256_6
timestamp 1731220380
transform 1 0 1896 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5255_6
timestamp 1731220380
transform 1 0 1936 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5254_6
timestamp 1731220380
transform 1 0 1864 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5253_6
timestamp 1731220380
transform 1 0 1808 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5252_6
timestamp 1731220380
transform 1 0 1752 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5251_6
timestamp 1731220380
transform 1 0 1696 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5250_6
timestamp 1731220380
transform 1 0 1640 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5249_6
timestamp 1731220380
transform 1 0 1936 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5248_6
timestamp 1731220380
transform 1 0 1856 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5247_6
timestamp 1731220380
transform 1 0 1776 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5246_6
timestamp 1731220380
transform 1 0 1712 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5245_6
timestamp 1731220380
transform 1 0 1656 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5244_6
timestamp 1731220380
transform 1 0 1600 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5243_6
timestamp 1731220380
transform 1 0 1848 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5242_6
timestamp 1731220380
transform 1 0 1760 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5241_6
timestamp 1731220380
transform 1 0 1672 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5240_6
timestamp 1731220380
transform 1 0 1592 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5239_6
timestamp 1731220380
transform 1 0 1520 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5238_6
timestamp 1731220380
transform 1 0 1824 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5237_6
timestamp 1731220380
transform 1 0 1720 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5236_6
timestamp 1731220380
transform 1 0 1624 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5235_6
timestamp 1731220380
transform 1 0 1528 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5234_6
timestamp 1731220380
transform 1 0 1448 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5233_6
timestamp 1731220380
transform 1 0 1384 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5232_6
timestamp 1731220380
transform 1 0 1776 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5231_6
timestamp 1731220380
transform 1 0 1696 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5230_6
timestamp 1731220380
transform 1 0 1616 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5229_6
timestamp 1731220380
transform 1 0 1552 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5228_6
timestamp 1731220380
transform 1 0 1496 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5227_6
timestamp 1731220380
transform 1 0 1440 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5226_6
timestamp 1731220380
transform 1 0 1384 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5225_6
timestamp 1731220380
transform 1 0 1256 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5224_6
timestamp 1731220380
transform 1 0 1200 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5223_6
timestamp 1731220380
transform 1 0 1136 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5222_6
timestamp 1731220380
transform 1 0 1240 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5221_6
timestamp 1731220380
transform 1 0 1240 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5220_6
timestamp 1731220380
transform 1 0 1128 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5219_6
timestamp 1731220380
transform 1 0 1184 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5218_6
timestamp 1731220380
transform 1 0 1080 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5217_6
timestamp 1731220380
transform 1 0 992 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5216_6
timestamp 1731220380
transform 1 0 912 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5215_6
timestamp 1731220380
transform 1 0 1072 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5214_6
timestamp 1731220380
transform 1 0 1160 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5213_6
timestamp 1731220380
transform 1 0 1248 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5212_6
timestamp 1731220380
transform 1 0 1208 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5211_6
timestamp 1731220380
transform 1 0 1128 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5210_6
timestamp 1731220380
transform 1 0 1056 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5209_6
timestamp 1731220380
transform 1 0 984 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5208_6
timestamp 1731220380
transform 1 0 912 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5207_6
timestamp 1731220380
transform 1 0 840 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5206_6
timestamp 1731220380
transform 1 0 1072 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5205_6
timestamp 1731220380
transform 1 0 992 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5204_6
timestamp 1731220380
transform 1 0 920 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5203_6
timestamp 1731220380
transform 1 0 848 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5202_6
timestamp 1731220380
transform 1 0 776 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5201_6
timestamp 1731220380
transform 1 0 704 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5200_6
timestamp 1731220380
transform 1 0 688 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5199_6
timestamp 1731220380
transform 1 0 800 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5198_6
timestamp 1731220380
transform 1 0 912 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5197_6
timestamp 1731220380
transform 1 0 872 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5196_6
timestamp 1731220380
transform 1 0 768 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5195_6
timestamp 1731220380
transform 1 0 664 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5194_6
timestamp 1731220380
transform 1 0 560 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5193_6
timestamp 1731220380
transform 1 0 592 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5192_6
timestamp 1731220380
transform 1 0 680 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5191_6
timestamp 1731220380
transform 1 0 760 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5190_6
timestamp 1731220380
transform 1 0 840 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5189_6
timestamp 1731220380
transform 1 0 920 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5188_6
timestamp 1731220380
transform 1 0 1008 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5187_6
timestamp 1731220380
transform 1 0 1160 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5186_6
timestamp 1731220380
transform 1 0 1064 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5185_6
timestamp 1731220380
transform 1 0 976 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5184_6
timestamp 1731220380
transform 1 0 888 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5183_6
timestamp 1731220380
transform 1 0 792 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5182_6
timestamp 1731220380
transform 1 0 688 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5181_6
timestamp 1731220380
transform 1 0 1064 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5180_6
timestamp 1731220380
transform 1 0 976 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5179_6
timestamp 1731220380
transform 1 0 888 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5178_6
timestamp 1731220380
transform 1 0 808 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5177_6
timestamp 1731220380
transform 1 0 728 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5176_6
timestamp 1731220380
transform 1 0 640 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5175_6
timestamp 1731220380
transform 1 0 904 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5174_6
timestamp 1731220380
transform 1 0 832 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5173_6
timestamp 1731220380
transform 1 0 760 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5172_6
timestamp 1731220380
transform 1 0 696 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5171_6
timestamp 1731220380
transform 1 0 632 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5170_6
timestamp 1731220380
transform 1 0 672 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5169_6
timestamp 1731220380
transform 1 0 784 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5168_6
timestamp 1731220380
transform 1 0 728 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5167_6
timestamp 1731220380
transform 1 0 704 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5166_6
timestamp 1731220380
transform 1 0 768 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5165_6
timestamp 1731220380
transform 1 0 672 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5164_6
timestamp 1731220380
transform 1 0 616 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5163_6
timestamp 1731220380
transform 1 0 568 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5162_6
timestamp 1731220380
transform 1 0 480 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5161_6
timestamp 1731220380
transform 1 0 424 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5160_6
timestamp 1731220380
transform 1 0 504 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5159_6
timestamp 1731220380
transform 1 0 504 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5158_6
timestamp 1731220380
transform 1 0 400 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5157_6
timestamp 1731220380
transform 1 0 496 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5156_6
timestamp 1731220380
transform 1 0 608 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5155_6
timestamp 1731220380
transform 1 0 632 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5154_6
timestamp 1731220380
transform 1 0 520 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5153_6
timestamp 1731220380
transform 1 0 416 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5152_6
timestamp 1731220380
transform 1 0 472 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5151_6
timestamp 1731220380
transform 1 0 568 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5150_6
timestamp 1731220380
transform 1 0 512 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5149_6
timestamp 1731220380
transform 1 0 440 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5148_6
timestamp 1731220380
transform 1 0 584 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5147_6
timestamp 1731220380
transform 1 0 632 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5146_6
timestamp 1731220380
transform 1 0 536 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5145_6
timestamp 1731220380
transform 1 0 440 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5144_6
timestamp 1731220380
transform 1 0 352 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5143_6
timestamp 1731220380
transform 1 0 272 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5142_6
timestamp 1731220380
transform 1 0 248 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5141_6
timestamp 1731220380
transform 1 0 304 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5140_6
timestamp 1731220380
transform 1 0 368 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5139_6
timestamp 1731220380
transform 1 0 368 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5138_6
timestamp 1731220380
transform 1 0 272 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5137_6
timestamp 1731220380
transform 1 0 184 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5136_6
timestamp 1731220380
transform 1 0 128 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5135_6
timestamp 1731220380
transform 1 0 216 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5134_6
timestamp 1731220380
transform 1 0 312 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5133_6
timestamp 1731220380
transform 1 0 384 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5132_6
timestamp 1731220380
transform 1 0 280 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5131_6
timestamp 1731220380
transform 1 0 192 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5130_6
timestamp 1731220380
transform 1 0 128 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5129_6
timestamp 1731220380
transform 1 0 128 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5128_6
timestamp 1731220380
transform 1 0 200 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5127_6
timestamp 1731220380
transform 1 0 296 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5126_6
timestamp 1731220380
transform 1 0 264 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5125_6
timestamp 1731220380
transform 1 0 184 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5124_6
timestamp 1731220380
transform 1 0 128 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5123_6
timestamp 1731220380
transform 1 0 344 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5122_6
timestamp 1731220380
transform 1 0 296 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5121_6
timestamp 1731220380
transform 1 0 208 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5120_6
timestamp 1731220380
transform 1 0 128 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5119_6
timestamp 1731220380
transform 1 0 392 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5118_6
timestamp 1731220380
transform 1 0 304 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5117_6
timestamp 1731220380
transform 1 0 208 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5116_6
timestamp 1731220380
transform 1 0 512 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5115_6
timestamp 1731220380
transform 1 0 408 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5114_6
timestamp 1731220380
transform 1 0 408 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5113_6
timestamp 1731220380
transform 1 0 336 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5112_6
timestamp 1731220380
transform 1 0 280 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5111_6
timestamp 1731220380
transform 1 0 488 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5110_6
timestamp 1731220380
transform 1 0 576 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5109_6
timestamp 1731220380
transform 1 0 512 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5108_6
timestamp 1731220380
transform 1 0 456 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5107_6
timestamp 1731220380
transform 1 0 400 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5106_6
timestamp 1731220380
transform 1 0 576 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5105_6
timestamp 1731220380
transform 1 0 640 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5104_6
timestamp 1731220380
transform 1 0 616 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5103_6
timestamp 1731220380
transform 1 0 560 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5102_6
timestamp 1731220380
transform 1 0 504 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5101_6
timestamp 1731220380
transform 1 0 448 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5100_6
timestamp 1731220380
transform 1 0 392 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_599_6
timestamp 1731220380
transform 1 0 568 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_598_6
timestamp 1731220380
transform 1 0 504 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_597_6
timestamp 1731220380
transform 1 0 440 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_596_6
timestamp 1731220380
transform 1 0 376 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_595_6
timestamp 1731220380
transform 1 0 320 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_594_6
timestamp 1731220380
transform 1 0 264 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_593_6
timestamp 1731220380
transform 1 0 552 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_592_6
timestamp 1731220380
transform 1 0 456 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_591_6
timestamp 1731220380
transform 1 0 368 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_590_6
timestamp 1731220380
transform 1 0 280 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_589_6
timestamp 1731220380
transform 1 0 200 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_588_6
timestamp 1731220380
transform 1 0 136 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_587_6
timestamp 1731220380
transform 1 0 584 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_586_6
timestamp 1731220380
transform 1 0 472 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_585_6
timestamp 1731220380
transform 1 0 368 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_584_6
timestamp 1731220380
transform 1 0 264 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_583_6
timestamp 1731220380
transform 1 0 184 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_582_6
timestamp 1731220380
transform 1 0 128 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_581_6
timestamp 1731220380
transform 1 0 328 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_580_6
timestamp 1731220380
transform 1 0 248 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_579_6
timestamp 1731220380
transform 1 0 184 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_578_6
timestamp 1731220380
transform 1 0 128 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_577_6
timestamp 1731220380
transform 1 0 504 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_576_6
timestamp 1731220380
transform 1 0 416 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_575_6
timestamp 1731220380
transform 1 0 240 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_574_6
timestamp 1731220380
transform 1 0 184 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_573_6
timestamp 1731220380
transform 1 0 128 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_572_6
timestamp 1731220380
transform 1 0 296 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_571_6
timestamp 1731220380
transform 1 0 464 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_570_6
timestamp 1731220380
transform 1 0 376 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_569_6
timestamp 1731220380
transform 1 0 304 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_568_6
timestamp 1731220380
transform 1 0 232 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_567_6
timestamp 1731220380
transform 1 0 168 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_566_6
timestamp 1731220380
transform 1 0 384 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_565_6
timestamp 1731220380
transform 1 0 584 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_564_6
timestamp 1731220380
transform 1 0 480 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_563_6
timestamp 1731220380
transform 1 0 408 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_562_6
timestamp 1731220380
transform 1 0 344 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_561_6
timestamp 1731220380
transform 1 0 288 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_560_6
timestamp 1731220380
transform 1 0 480 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_559_6
timestamp 1731220380
transform 1 0 632 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_558_6
timestamp 1731220380
transform 1 0 560 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_557_6
timestamp 1731220380
transform 1 0 544 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_556_6
timestamp 1731220380
transform 1 0 480 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_555_6
timestamp 1731220380
transform 1 0 424 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_554_6
timestamp 1731220380
transform 1 0 616 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_553_6
timestamp 1731220380
transform 1 0 696 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_552_6
timestamp 1731220380
transform 1 0 768 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_551_6
timestamp 1731220380
transform 1 0 752 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_550_6
timestamp 1731220380
transform 1 0 832 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_549_6
timestamp 1731220380
transform 1 0 816 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_548_6
timestamp 1731220380
transform 1 0 736 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_547_6
timestamp 1731220380
transform 1 0 896 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_546_6
timestamp 1731220380
transform 1 0 984 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_545_6
timestamp 1731220380
transform 1 0 912 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_544_6
timestamp 1731220380
transform 1 0 808 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_543_6
timestamp 1731220380
transform 1 0 1016 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_542_6
timestamp 1731220380
transform 1 0 1000 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_541_6
timestamp 1731220380
transform 1 0 880 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_540_6
timestamp 1731220380
transform 1 0 1120 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_539_6
timestamp 1731220380
transform 1 0 1064 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_538_6
timestamp 1731220380
transform 1 0 1000 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_537_6
timestamp 1731220380
transform 1 0 936 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_536_6
timestamp 1731220380
transform 1 0 872 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_535_6
timestamp 1731220380
transform 1 0 808 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_534_6
timestamp 1731220380
transform 1 0 744 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_533_6
timestamp 1731220380
transform 1 0 688 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_532_6
timestamp 1731220380
transform 1 0 632 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_531_6
timestamp 1731220380
transform 1 0 648 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_530_6
timestamp 1731220380
transform 1 0 760 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_529_6
timestamp 1731220380
transform 1 0 704 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_528_6
timestamp 1731220380
transform 1 0 664 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_527_6
timestamp 1731220380
transform 1 0 600 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_526_6
timestamp 1731220380
transform 1 0 544 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_525_6
timestamp 1731220380
transform 1 0 672 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_524_6
timestamp 1731220380
transform 1 0 592 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_523_6
timestamp 1731220380
transform 1 0 520 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_522_6
timestamp 1731220380
transform 1 0 456 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_521_6
timestamp 1731220380
transform 1 0 400 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_520_6
timestamp 1731220380
transform 1 0 432 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_519_6
timestamp 1731220380
transform 1 0 488 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_518_6
timestamp 1731220380
transform 1 0 608 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_517_6
timestamp 1731220380
transform 1 0 512 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_516_6
timestamp 1731220380
transform 1 0 424 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_515_6
timestamp 1731220380
transform 1 0 344 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_514_6
timestamp 1731220380
transform 1 0 272 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_513_6
timestamp 1731220380
transform 1 0 536 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_512_6
timestamp 1731220380
transform 1 0 432 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_511_6
timestamp 1731220380
transform 1 0 328 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_510_6
timestamp 1731220380
transform 1 0 240 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_59_6
timestamp 1731220380
transform 1 0 168 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_58_6
timestamp 1731220380
transform 1 0 576 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_57_6
timestamp 1731220380
transform 1 0 520 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_56_6
timestamp 1731220380
transform 1 0 464 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_55_6
timestamp 1731220380
transform 1 0 408 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_54_6
timestamp 1731220380
transform 1 0 352 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_53_6
timestamp 1731220380
transform 1 0 296 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_52_6
timestamp 1731220380
transform 1 0 240 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_51_6
timestamp 1731220380
transform 1 0 184 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_50_6
timestamp 1731220380
transform 1 0 128 0 1 80
box 8 4 52 52
<< end >>
