magic
tech sky130l
timestamp 1730954142
<< m1 >>
rect 736 1183 740 1259
rect 240 971 244 991
rect 736 971 740 991
rect 1168 951 1172 991
rect 1168 783 1172 831
rect 1168 639 1172 667
rect 216 515 220 619
rect 1168 487 1172 519
rect 1168 359 1172 471
rect 864 219 868 267
rect 288 171 292 215
<< m2c >>
rect 736 1259 740 1263
rect 111 1253 115 1257
rect 111 1235 115 1239
rect 111 1185 115 1189
rect 1183 1253 1187 1257
rect 1183 1235 1187 1239
rect 1183 1185 1187 1189
rect 736 1179 740 1183
rect 111 1167 115 1171
rect 1183 1167 1187 1171
rect 111 1101 115 1105
rect 1183 1101 1187 1105
rect 111 1083 115 1087
rect 1183 1083 1187 1087
rect 111 1017 115 1021
rect 1183 1017 1187 1021
rect 111 999 115 1003
rect 1183 999 1187 1003
rect 240 991 244 995
rect 240 967 244 971
rect 736 991 740 995
rect 736 967 740 971
rect 1168 991 1172 995
rect 1168 947 1172 951
rect 111 933 115 937
rect 1183 933 1187 937
rect 111 915 115 919
rect 1183 915 1187 919
rect 111 857 115 861
rect 1000 859 1004 863
rect 1183 857 1187 861
rect 111 839 115 843
rect 1183 839 1187 843
rect 1168 831 1172 835
rect 1168 779 1172 783
rect 111 765 115 769
rect 1183 765 1187 769
rect 111 747 115 751
rect 1183 747 1187 751
rect 111 693 115 697
rect 1183 693 1187 697
rect 111 675 115 679
rect 1183 675 1187 679
rect 1168 667 1172 671
rect 1168 635 1172 639
rect 216 619 220 623
rect 111 613 115 617
rect 111 595 115 599
rect 111 545 115 549
rect 111 527 115 531
rect 1183 613 1187 617
rect 1183 595 1187 599
rect 1183 545 1187 549
rect 1183 527 1187 531
rect 216 511 220 515
rect 1168 519 1172 523
rect 1168 483 1172 487
rect 1168 471 1172 475
rect 111 461 115 465
rect 111 443 115 447
rect 111 389 115 393
rect 111 371 115 375
rect 1183 461 1187 465
rect 1183 443 1187 447
rect 1183 389 1187 393
rect 1183 371 1187 375
rect 1168 355 1172 359
rect 111 313 115 317
rect 1183 313 1187 317
rect 111 295 115 299
rect 1183 295 1187 299
rect 864 267 868 271
rect 111 241 115 245
rect 111 223 115 227
rect 1183 241 1187 245
rect 1183 223 1187 227
rect 288 215 292 219
rect 864 215 868 219
rect 288 167 292 171
rect 111 137 115 141
rect 1183 137 1187 141
rect 111 119 115 123
rect 1183 119 1187 123
<< m2 >>
rect 662 1275 668 1276
rect 662 1271 663 1275
rect 667 1271 668 1275
rect 662 1270 668 1271
rect 750 1275 756 1276
rect 750 1271 751 1275
rect 755 1271 756 1275
rect 750 1270 756 1271
rect 838 1275 844 1276
rect 838 1271 839 1275
rect 843 1271 844 1275
rect 838 1270 844 1271
rect 926 1275 932 1276
rect 926 1271 927 1275
rect 931 1271 932 1275
rect 926 1270 932 1271
rect 990 1271 996 1272
rect 733 1268 746 1270
rect 821 1268 834 1270
rect 909 1268 922 1270
rect 713 1264 738 1266
rect 744 1265 746 1268
rect 832 1265 834 1268
rect 920 1265 922 1268
rect 990 1267 991 1271
rect 995 1267 996 1271
rect 990 1266 996 1267
rect 735 1263 741 1264
rect 735 1259 736 1263
rect 740 1259 741 1263
rect 735 1258 741 1259
rect 110 1257 116 1258
rect 110 1253 111 1257
rect 115 1253 116 1257
rect 110 1252 116 1253
rect 1182 1257 1188 1258
rect 1182 1253 1183 1257
rect 1187 1253 1188 1257
rect 1182 1252 1188 1253
rect 110 1239 116 1240
rect 110 1235 111 1239
rect 115 1235 116 1239
rect 1182 1239 1188 1240
rect 1182 1235 1183 1239
rect 1187 1235 1188 1239
rect 110 1234 116 1235
rect 666 1234 672 1235
rect 666 1230 667 1234
rect 671 1230 672 1234
rect 666 1229 672 1230
rect 754 1234 760 1235
rect 754 1230 755 1234
rect 759 1230 760 1234
rect 754 1229 760 1230
rect 842 1234 848 1235
rect 842 1230 843 1234
rect 847 1230 848 1234
rect 842 1229 848 1230
rect 930 1234 936 1235
rect 1182 1234 1188 1235
rect 930 1230 931 1234
rect 935 1230 936 1234
rect 930 1229 936 1230
rect 370 1194 376 1195
rect 370 1190 371 1194
rect 375 1190 376 1194
rect 110 1189 116 1190
rect 370 1189 376 1190
rect 458 1194 464 1195
rect 458 1190 459 1194
rect 463 1190 464 1194
rect 458 1189 464 1190
rect 554 1194 560 1195
rect 554 1190 555 1194
rect 559 1190 560 1194
rect 554 1189 560 1190
rect 650 1194 656 1195
rect 650 1190 651 1194
rect 655 1190 656 1194
rect 650 1189 656 1190
rect 754 1194 760 1195
rect 754 1190 755 1194
rect 759 1190 760 1194
rect 754 1189 760 1190
rect 858 1194 864 1195
rect 858 1190 859 1194
rect 863 1190 864 1194
rect 858 1189 864 1190
rect 962 1194 968 1195
rect 962 1190 963 1194
rect 967 1190 968 1194
rect 962 1189 968 1190
rect 1182 1189 1188 1190
rect 110 1185 111 1189
rect 115 1185 116 1189
rect 110 1184 116 1185
rect 1182 1185 1183 1189
rect 1187 1185 1188 1189
rect 1182 1184 1188 1185
rect 735 1183 741 1184
rect 735 1179 736 1183
rect 740 1182 741 1183
rect 740 1180 818 1182
rect 740 1179 741 1180
rect 735 1178 741 1179
rect 814 1179 820 1180
rect 814 1175 815 1179
rect 819 1175 820 1179
rect 814 1174 820 1175
rect 110 1171 116 1172
rect 110 1167 111 1171
rect 115 1167 116 1171
rect 110 1166 116 1167
rect 1182 1171 1188 1172
rect 1182 1167 1183 1171
rect 1187 1167 1188 1171
rect 1182 1166 1188 1167
rect 438 1163 444 1164
rect 438 1162 439 1163
rect 417 1160 439 1162
rect 438 1159 439 1160
rect 443 1159 444 1163
rect 934 1163 940 1164
rect 934 1162 935 1163
rect 438 1158 444 1159
rect 448 1154 450 1161
rect 520 1160 545 1162
rect 616 1160 641 1162
rect 712 1160 745 1162
rect 905 1160 935 1162
rect 520 1155 522 1160
rect 616 1155 618 1160
rect 712 1155 714 1160
rect 934 1159 935 1160
rect 939 1159 940 1163
rect 934 1158 940 1159
rect 982 1163 988 1164
rect 982 1159 983 1163
rect 987 1159 988 1163
rect 982 1158 988 1159
rect 814 1155 820 1156
rect 366 1153 372 1154
rect 366 1149 367 1153
rect 371 1149 372 1153
rect 437 1152 450 1154
rect 454 1153 460 1154
rect 366 1148 372 1149
rect 454 1149 455 1153
rect 459 1149 460 1153
rect 454 1148 460 1149
rect 550 1153 556 1154
rect 550 1149 551 1153
rect 555 1149 556 1153
rect 550 1148 556 1149
rect 646 1153 652 1154
rect 646 1149 647 1153
rect 651 1149 652 1153
rect 646 1148 652 1149
rect 750 1153 756 1154
rect 750 1149 751 1153
rect 755 1149 756 1153
rect 814 1151 815 1155
rect 819 1151 820 1155
rect 922 1155 928 1156
rect 814 1150 820 1151
rect 854 1153 860 1154
rect 750 1148 756 1149
rect 854 1149 855 1153
rect 859 1149 860 1153
rect 922 1151 923 1155
rect 927 1151 928 1155
rect 922 1150 928 1151
rect 958 1153 964 1154
rect 854 1148 860 1149
rect 958 1149 959 1153
rect 963 1149 964 1153
rect 958 1148 964 1149
rect 1024 1146 1026 1151
rect 1020 1144 1026 1146
rect 934 1139 940 1140
rect 934 1135 935 1139
rect 939 1138 940 1139
rect 1020 1138 1022 1144
rect 939 1136 1022 1138
rect 939 1135 940 1136
rect 934 1134 940 1135
rect 142 1123 148 1124
rect 142 1119 143 1123
rect 147 1119 148 1123
rect 142 1118 148 1119
rect 254 1123 260 1124
rect 254 1119 255 1123
rect 259 1119 260 1123
rect 254 1118 260 1119
rect 414 1123 420 1124
rect 414 1119 415 1123
rect 419 1119 420 1123
rect 414 1118 420 1119
rect 582 1123 588 1124
rect 582 1119 583 1123
rect 587 1119 588 1123
rect 582 1118 588 1119
rect 766 1123 772 1124
rect 766 1119 767 1123
rect 771 1119 772 1123
rect 766 1118 772 1119
rect 830 1123 836 1124
rect 830 1119 831 1123
rect 835 1119 836 1123
rect 830 1118 836 1119
rect 950 1123 956 1124
rect 950 1119 951 1123
rect 955 1119 956 1123
rect 950 1118 956 1119
rect 1014 1119 1020 1120
rect 213 1116 250 1118
rect 325 1116 410 1118
rect 485 1116 578 1118
rect 653 1116 681 1118
rect 193 1112 218 1114
rect 248 1113 250 1116
rect 408 1113 410 1116
rect 576 1113 578 1116
rect 679 1114 681 1116
rect 922 1115 928 1116
rect 679 1112 761 1114
rect 214 1111 220 1112
rect 214 1107 215 1111
rect 219 1107 220 1111
rect 922 1111 923 1115
rect 927 1114 928 1115
rect 1014 1115 1015 1119
rect 1019 1115 1020 1119
rect 1014 1114 1020 1115
rect 927 1112 945 1114
rect 927 1111 928 1112
rect 922 1110 928 1111
rect 214 1106 220 1107
rect 110 1105 116 1106
rect 110 1101 111 1105
rect 115 1101 116 1105
rect 110 1100 116 1101
rect 1182 1105 1188 1106
rect 1182 1101 1183 1105
rect 1187 1101 1188 1105
rect 1182 1100 1188 1101
rect 110 1087 116 1088
rect 110 1083 111 1087
rect 115 1083 116 1087
rect 1182 1087 1188 1088
rect 1182 1083 1183 1087
rect 1187 1083 1188 1087
rect 110 1082 116 1083
rect 146 1082 152 1083
rect 146 1078 147 1082
rect 151 1078 152 1082
rect 146 1077 152 1078
rect 258 1082 264 1083
rect 258 1078 259 1082
rect 263 1078 264 1082
rect 258 1077 264 1078
rect 418 1082 424 1083
rect 418 1078 419 1082
rect 423 1078 424 1082
rect 418 1077 424 1078
rect 586 1082 592 1083
rect 586 1078 587 1082
rect 591 1078 592 1082
rect 586 1077 592 1078
rect 770 1082 776 1083
rect 770 1078 771 1082
rect 775 1078 776 1082
rect 770 1077 776 1078
rect 954 1082 960 1083
rect 1182 1082 1188 1083
rect 954 1078 955 1082
rect 959 1078 960 1082
rect 954 1077 960 1078
rect 154 1026 160 1027
rect 154 1022 155 1026
rect 159 1022 160 1026
rect 110 1021 116 1022
rect 154 1021 160 1022
rect 282 1026 288 1027
rect 282 1022 283 1026
rect 287 1022 288 1026
rect 282 1021 288 1022
rect 426 1026 432 1027
rect 426 1022 427 1026
rect 431 1022 432 1026
rect 426 1021 432 1022
rect 586 1026 592 1027
rect 586 1022 587 1026
rect 591 1022 592 1026
rect 586 1021 592 1022
rect 754 1026 760 1027
rect 754 1022 755 1026
rect 759 1022 760 1026
rect 754 1021 760 1022
rect 938 1026 944 1027
rect 938 1022 939 1026
rect 943 1022 944 1026
rect 938 1021 944 1022
rect 1098 1026 1104 1027
rect 1098 1022 1099 1026
rect 1103 1022 1104 1026
rect 1098 1021 1104 1022
rect 1182 1021 1188 1022
rect 110 1017 111 1021
rect 115 1017 116 1021
rect 110 1016 116 1017
rect 1182 1017 1183 1021
rect 1187 1017 1188 1021
rect 1182 1016 1188 1017
rect 110 1003 116 1004
rect 110 999 111 1003
rect 115 999 116 1003
rect 110 998 116 999
rect 1182 1003 1188 1004
rect 1182 999 1183 1003
rect 1187 999 1188 1003
rect 1182 998 1188 999
rect 239 995 245 996
rect 239 994 240 995
rect 201 992 240 994
rect 239 991 240 992
rect 244 991 245 995
rect 378 995 384 996
rect 378 994 379 995
rect 329 992 379 994
rect 239 990 245 991
rect 378 991 379 992
rect 383 991 384 995
rect 542 995 548 996
rect 542 994 543 995
rect 473 992 543 994
rect 378 990 384 991
rect 542 991 543 992
rect 547 991 548 995
rect 735 995 741 996
rect 735 994 736 995
rect 633 992 736 994
rect 542 990 548 991
rect 735 991 736 992
rect 740 991 741 995
rect 735 990 741 991
rect 762 995 768 996
rect 762 991 763 995
rect 767 991 768 995
rect 1014 995 1020 996
rect 1014 994 1015 995
rect 985 992 1015 994
rect 762 990 768 991
rect 1014 991 1015 992
rect 1019 991 1020 995
rect 1167 995 1173 996
rect 1167 994 1168 995
rect 1145 992 1168 994
rect 1014 990 1020 991
rect 1167 991 1168 992
rect 1172 991 1173 995
rect 1167 990 1173 991
rect 214 987 220 988
rect 150 985 156 986
rect 150 981 151 985
rect 155 981 156 985
rect 214 983 215 987
rect 219 983 220 987
rect 214 982 220 983
rect 278 985 284 986
rect 150 980 156 981
rect 278 981 279 985
rect 283 981 284 985
rect 422 985 428 986
rect 344 982 346 983
rect 278 980 284 981
rect 340 980 346 982
rect 422 981 423 985
rect 427 981 428 985
rect 582 985 588 986
rect 488 982 490 983
rect 422 980 428 981
rect 484 980 490 982
rect 582 981 583 985
rect 587 981 588 985
rect 750 985 756 986
rect 648 982 650 983
rect 582 980 588 981
rect 644 980 650 982
rect 750 981 751 985
rect 755 981 756 985
rect 934 985 940 986
rect 750 980 756 981
rect 239 971 245 972
rect 239 967 240 971
rect 244 970 245 971
rect 340 970 342 980
rect 244 968 342 970
rect 378 971 384 972
rect 244 967 245 968
rect 239 966 245 967
rect 378 967 379 971
rect 383 970 384 971
rect 484 970 486 980
rect 383 968 486 970
rect 542 971 548 972
rect 383 967 384 968
rect 378 966 384 967
rect 542 967 543 971
rect 547 970 548 971
rect 644 970 646 980
rect 547 968 646 970
rect 735 971 741 972
rect 547 967 548 968
rect 542 966 548 967
rect 735 967 736 971
rect 740 970 741 971
rect 816 970 818 983
rect 934 981 935 985
rect 939 981 940 985
rect 1094 985 1100 986
rect 934 980 940 981
rect 990 979 996 980
rect 990 975 991 979
rect 995 978 996 979
rect 1000 978 1002 983
rect 1094 981 1095 985
rect 1099 981 1100 985
rect 1094 980 1100 981
rect 995 976 1002 978
rect 995 975 996 976
rect 990 974 996 975
rect 740 968 818 970
rect 740 967 741 968
rect 735 966 741 967
rect 812 964 958 966
rect 810 963 816 964
rect 810 959 811 963
rect 815 959 816 963
rect 810 958 816 959
rect 956 958 958 964
rect 956 956 962 958
rect 502 955 508 956
rect 502 951 503 955
rect 507 951 508 955
rect 502 950 508 951
rect 590 955 596 956
rect 590 951 591 955
rect 595 951 596 955
rect 590 950 596 951
rect 686 955 692 956
rect 686 951 687 955
rect 691 951 692 955
rect 790 955 796 956
rect 686 950 692 951
rect 762 951 768 952
rect 762 950 763 951
rect 573 948 586 950
rect 661 948 681 950
rect 757 948 763 950
rect 553 944 578 946
rect 584 945 586 948
rect 679 944 681 948
rect 762 947 763 948
rect 767 947 768 951
rect 790 951 791 955
rect 795 951 796 955
rect 894 955 900 956
rect 790 950 796 951
rect 854 951 860 952
rect 762 946 768 947
rect 854 947 855 951
rect 859 947 860 951
rect 894 951 895 955
rect 899 951 900 955
rect 960 953 962 956
rect 1006 955 1012 956
rect 894 950 900 951
rect 1006 951 1007 955
rect 1011 951 1012 955
rect 1006 950 1012 951
rect 1094 955 1100 956
rect 1094 951 1095 955
rect 1099 951 1100 955
rect 1094 950 1100 951
rect 1167 951 1173 952
rect 1167 950 1168 951
rect 1077 948 1090 950
rect 1165 948 1168 950
rect 854 946 860 947
rect 982 947 988 948
rect 982 946 983 947
rect 945 944 983 946
rect 574 943 580 944
rect 574 939 575 943
rect 579 939 580 943
rect 574 938 580 939
rect 810 943 816 944
rect 810 939 811 943
rect 815 939 816 943
rect 982 943 983 944
rect 987 943 988 947
rect 1057 944 1082 946
rect 1088 945 1090 948
rect 1167 947 1168 948
rect 1172 947 1173 951
rect 1167 946 1173 947
rect 982 942 988 943
rect 1078 943 1084 944
rect 810 938 816 939
rect 1078 939 1079 943
rect 1083 939 1084 943
rect 1078 938 1084 939
rect 110 937 116 938
rect 110 933 111 937
rect 115 933 116 937
rect 110 932 116 933
rect 1182 937 1188 938
rect 1182 933 1183 937
rect 1187 933 1188 937
rect 1182 932 1188 933
rect 110 919 116 920
rect 110 915 111 919
rect 115 915 116 919
rect 1182 919 1188 920
rect 1182 915 1183 919
rect 1187 915 1188 919
rect 110 914 116 915
rect 506 914 512 915
rect 506 910 507 914
rect 511 910 512 914
rect 506 909 512 910
rect 594 914 600 915
rect 594 910 595 914
rect 599 910 600 914
rect 594 909 600 910
rect 690 914 696 915
rect 690 910 691 914
rect 695 910 696 914
rect 690 909 696 910
rect 794 914 800 915
rect 794 910 795 914
rect 799 910 800 914
rect 794 909 800 910
rect 898 914 904 915
rect 898 910 899 914
rect 903 910 904 914
rect 898 909 904 910
rect 1010 914 1016 915
rect 1010 910 1011 914
rect 1015 910 1016 914
rect 1010 909 1016 910
rect 1098 914 1104 915
rect 1182 914 1188 915
rect 1098 910 1099 914
rect 1103 910 1104 914
rect 1098 909 1104 910
rect 1078 887 1084 888
rect 1078 883 1079 887
rect 1083 886 1084 887
rect 1158 887 1164 888
rect 1158 886 1159 887
rect 1083 884 1159 886
rect 1083 883 1084 884
rect 1078 882 1084 883
rect 1158 883 1159 884
rect 1163 883 1164 887
rect 1158 882 1164 883
rect 562 866 568 867
rect 562 862 563 866
rect 567 862 568 866
rect 110 861 116 862
rect 562 861 568 862
rect 650 866 656 867
rect 650 862 651 866
rect 655 862 656 866
rect 650 861 656 862
rect 738 866 744 867
rect 738 862 739 866
rect 743 862 744 866
rect 738 861 744 862
rect 826 866 832 867
rect 826 862 827 866
rect 831 862 832 866
rect 826 861 832 862
rect 922 866 928 867
rect 922 862 923 866
rect 927 862 928 866
rect 1010 866 1016 867
rect 922 861 928 862
rect 990 863 996 864
rect 110 857 111 861
rect 115 857 116 861
rect 990 859 991 863
rect 995 862 996 863
rect 999 863 1005 864
rect 999 862 1000 863
rect 995 860 1000 862
rect 995 859 996 860
rect 990 858 996 859
rect 999 859 1000 860
rect 1004 859 1005 863
rect 1010 862 1011 866
rect 1015 862 1016 866
rect 1010 861 1016 862
rect 1098 866 1104 867
rect 1098 862 1099 866
rect 1103 862 1104 866
rect 1098 861 1104 862
rect 1182 861 1188 862
rect 999 858 1005 859
rect 110 856 116 857
rect 1182 857 1183 861
rect 1187 857 1188 861
rect 1182 856 1188 857
rect 110 843 116 844
rect 110 839 111 843
rect 115 839 116 843
rect 110 838 116 839
rect 1182 843 1188 844
rect 1182 839 1183 843
rect 1187 839 1188 843
rect 1182 838 1188 839
rect 630 835 636 836
rect 630 834 631 835
rect 609 832 631 834
rect 630 831 631 832
rect 635 831 636 835
rect 1167 835 1173 836
rect 1167 834 1168 835
rect 630 830 636 831
rect 640 826 642 833
rect 712 832 729 834
rect 800 832 817 834
rect 888 832 913 834
rect 1145 832 1168 834
rect 712 827 714 832
rect 800 827 802 832
rect 888 827 890 832
rect 1167 831 1168 832
rect 1172 831 1173 835
rect 1167 830 1173 831
rect 982 827 988 828
rect 558 825 564 826
rect 558 821 559 825
rect 563 821 564 825
rect 629 824 642 826
rect 646 825 652 826
rect 558 820 564 821
rect 646 821 647 825
rect 651 821 652 825
rect 646 820 652 821
rect 734 825 740 826
rect 734 821 735 825
rect 739 821 740 825
rect 734 820 740 821
rect 822 825 828 826
rect 822 821 823 825
rect 827 821 828 825
rect 822 820 828 821
rect 918 825 924 826
rect 918 821 919 825
rect 923 821 924 825
rect 982 823 983 827
rect 987 823 988 827
rect 1158 827 1164 828
rect 982 822 988 823
rect 1006 825 1012 826
rect 918 820 924 821
rect 1006 821 1007 825
rect 1011 821 1012 825
rect 1094 825 1100 826
rect 1072 822 1074 823
rect 1006 820 1012 821
rect 1068 820 1074 822
rect 1094 821 1095 825
rect 1099 821 1100 825
rect 1158 823 1159 827
rect 1163 823 1164 827
rect 1158 822 1164 823
rect 1094 820 1100 821
rect 998 811 1004 812
rect 998 807 999 811
rect 1003 810 1004 811
rect 1068 810 1070 820
rect 1003 808 1070 810
rect 1003 807 1004 808
rect 998 806 1004 807
rect 390 787 396 788
rect 390 783 391 787
rect 395 783 396 787
rect 390 782 396 783
rect 494 787 500 788
rect 494 783 495 787
rect 499 783 500 787
rect 494 782 500 783
rect 606 787 612 788
rect 606 783 607 787
rect 611 783 612 787
rect 606 782 612 783
rect 726 787 732 788
rect 726 783 727 787
rect 731 783 732 787
rect 726 782 732 783
rect 854 787 860 788
rect 854 783 855 787
rect 859 783 860 787
rect 982 787 988 788
rect 854 782 860 783
rect 918 783 924 784
rect 461 780 490 782
rect 565 780 602 782
rect 677 780 681 782
rect 797 780 850 782
rect 441 776 482 778
rect 488 777 490 780
rect 600 777 602 780
rect 679 778 681 780
rect 679 776 721 778
rect 848 777 850 780
rect 918 779 919 783
rect 923 779 924 783
rect 982 783 983 787
rect 987 783 988 787
rect 1094 787 1100 788
rect 982 782 988 783
rect 1046 783 1052 784
rect 918 778 924 779
rect 1046 779 1047 783
rect 1051 779 1052 783
rect 1094 783 1095 787
rect 1099 783 1100 787
rect 1094 782 1100 783
rect 1167 783 1173 784
rect 1167 782 1168 783
rect 1165 780 1168 782
rect 1046 778 1052 779
rect 1167 779 1168 780
rect 1172 779 1173 783
rect 1167 778 1173 779
rect 478 775 484 776
rect 478 771 479 775
rect 483 771 484 775
rect 478 770 484 771
rect 998 775 1004 776
rect 998 771 999 775
rect 1003 771 1004 775
rect 998 770 1004 771
rect 1118 775 1124 776
rect 1118 771 1119 775
rect 1123 771 1124 775
rect 1118 770 1124 771
rect 110 769 116 770
rect 110 765 111 769
rect 115 765 116 769
rect 110 764 116 765
rect 1182 769 1188 770
rect 1182 765 1183 769
rect 1187 765 1188 769
rect 1182 764 1188 765
rect 110 751 116 752
rect 110 747 111 751
rect 115 747 116 751
rect 1182 751 1188 752
rect 1182 747 1183 751
rect 1187 747 1188 751
rect 110 746 116 747
rect 394 746 400 747
rect 394 742 395 746
rect 399 742 400 746
rect 394 741 400 742
rect 498 746 504 747
rect 498 742 499 746
rect 503 742 504 746
rect 498 741 504 742
rect 610 746 616 747
rect 610 742 611 746
rect 615 742 616 746
rect 610 741 616 742
rect 730 746 736 747
rect 730 742 731 746
rect 735 742 736 746
rect 730 741 736 742
rect 858 746 864 747
rect 858 742 859 746
rect 863 742 864 746
rect 858 741 864 742
rect 986 746 992 747
rect 986 742 987 746
rect 991 742 992 746
rect 986 741 992 742
rect 1098 746 1104 747
rect 1182 746 1188 747
rect 1098 742 1099 746
rect 1103 742 1104 746
rect 1098 741 1104 742
rect 1122 723 1128 724
rect 1122 719 1123 723
rect 1127 722 1128 723
rect 1170 723 1176 724
rect 1170 722 1171 723
rect 1127 720 1171 722
rect 1127 719 1128 720
rect 1122 718 1128 719
rect 1170 719 1171 720
rect 1175 719 1176 723
rect 1170 718 1176 719
rect 210 702 216 703
rect 210 698 211 702
rect 215 698 216 702
rect 110 697 116 698
rect 210 697 216 698
rect 354 702 360 703
rect 354 698 355 702
rect 359 698 360 702
rect 354 697 360 698
rect 522 702 528 703
rect 522 698 523 702
rect 527 698 528 702
rect 522 697 528 698
rect 714 702 720 703
rect 714 698 715 702
rect 719 698 720 702
rect 714 697 720 698
rect 914 702 920 703
rect 914 698 915 702
rect 919 698 920 702
rect 914 697 920 698
rect 1098 702 1104 703
rect 1098 698 1099 702
rect 1103 698 1104 702
rect 1098 697 1104 698
rect 1182 697 1188 698
rect 110 693 111 697
rect 115 693 116 697
rect 110 692 116 693
rect 1182 693 1183 697
rect 1187 693 1188 697
rect 1182 692 1188 693
rect 110 679 116 680
rect 110 675 111 679
rect 115 675 116 679
rect 110 674 116 675
rect 1182 679 1188 680
rect 1182 675 1183 679
rect 1187 675 1188 679
rect 1182 674 1188 675
rect 334 671 340 672
rect 334 670 335 671
rect 257 668 335 670
rect 334 667 335 668
rect 339 667 340 671
rect 1167 671 1173 672
rect 1167 670 1168 671
rect 334 666 340 667
rect 344 662 346 669
rect 416 668 513 670
rect 679 668 705 670
rect 776 668 905 670
rect 1145 668 1168 670
rect 416 663 418 668
rect 679 662 681 668
rect 776 663 778 668
rect 1167 667 1168 668
rect 1172 667 1173 671
rect 1167 666 1173 667
rect 1170 663 1176 664
rect 1170 662 1171 663
rect 206 661 212 662
rect 206 657 207 661
rect 211 657 212 661
rect 277 660 346 662
rect 350 661 356 662
rect 206 656 212 657
rect 350 657 351 661
rect 355 657 356 661
rect 350 656 356 657
rect 518 661 524 662
rect 518 657 519 661
rect 523 657 524 661
rect 589 660 681 662
rect 710 661 716 662
rect 518 656 524 657
rect 710 657 711 661
rect 715 657 716 661
rect 710 656 716 657
rect 910 661 916 662
rect 910 657 911 661
rect 915 657 916 661
rect 1094 661 1100 662
rect 910 656 916 657
rect 478 647 484 648
rect 478 643 479 647
rect 483 646 484 647
rect 976 646 978 659
rect 1094 657 1095 661
rect 1099 657 1100 661
rect 1165 660 1171 662
rect 1170 659 1171 660
rect 1175 659 1176 663
rect 1170 658 1176 659
rect 1094 656 1100 657
rect 483 644 978 646
rect 483 643 484 644
rect 478 642 484 643
rect 1167 639 1173 640
rect 1167 638 1168 639
rect 1160 636 1168 638
rect 142 635 148 636
rect 142 631 143 635
rect 147 631 148 635
rect 142 630 148 631
rect 294 635 300 636
rect 294 631 295 635
rect 299 631 300 635
rect 294 630 300 631
rect 486 635 492 636
rect 486 631 487 635
rect 491 631 492 635
rect 486 630 492 631
rect 686 635 692 636
rect 686 631 687 635
rect 691 631 692 635
rect 686 630 692 631
rect 750 635 756 636
rect 750 631 751 635
rect 755 631 756 635
rect 750 630 756 631
rect 894 635 900 636
rect 894 631 895 635
rect 899 631 900 635
rect 894 630 900 631
rect 958 635 964 636
rect 958 631 959 635
rect 963 631 964 635
rect 958 630 964 631
rect 1094 635 1100 636
rect 1094 631 1095 635
rect 1099 631 1100 635
rect 1160 633 1162 636
rect 1167 635 1168 636
rect 1172 635 1173 639
rect 1167 634 1173 635
rect 1094 630 1100 631
rect 213 628 290 630
rect 365 628 482 630
rect 557 628 681 630
rect 193 624 218 626
rect 288 625 290 628
rect 480 625 482 628
rect 679 624 681 628
rect 1046 627 1052 628
rect 1046 626 1047 627
rect 945 624 1047 626
rect 215 623 221 624
rect 215 619 216 623
rect 220 619 221 623
rect 1046 623 1047 624
rect 1051 623 1052 627
rect 1145 624 1166 626
rect 1046 622 1052 623
rect 1164 622 1166 624
rect 1170 623 1176 624
rect 1170 622 1171 623
rect 1164 620 1171 622
rect 215 618 221 619
rect 1170 619 1171 620
rect 1175 619 1176 623
rect 1170 618 1176 619
rect 110 617 116 618
rect 110 613 111 617
rect 115 613 116 617
rect 110 612 116 613
rect 1182 617 1188 618
rect 1182 613 1183 617
rect 1187 613 1188 617
rect 1182 612 1188 613
rect 110 599 116 600
rect 110 595 111 599
rect 115 595 116 599
rect 1182 599 1188 600
rect 1182 595 1183 599
rect 1187 595 1188 599
rect 110 594 116 595
rect 146 594 152 595
rect 146 590 147 594
rect 151 590 152 594
rect 146 589 152 590
rect 298 594 304 595
rect 298 590 299 594
rect 303 590 304 594
rect 298 589 304 590
rect 490 594 496 595
rect 490 590 491 594
rect 495 590 496 594
rect 490 589 496 590
rect 690 594 696 595
rect 690 590 691 594
rect 695 590 696 594
rect 690 589 696 590
rect 898 594 904 595
rect 898 590 899 594
rect 903 590 904 594
rect 898 589 904 590
rect 1098 594 1104 595
rect 1182 594 1188 595
rect 1098 590 1099 594
rect 1103 590 1104 594
rect 1098 589 1104 590
rect 146 554 152 555
rect 146 550 147 554
rect 151 550 152 554
rect 110 549 116 550
rect 146 549 152 550
rect 282 554 288 555
rect 282 550 283 554
rect 287 550 288 554
rect 282 549 288 550
rect 466 554 472 555
rect 466 550 467 554
rect 471 550 472 554
rect 466 549 472 550
rect 666 554 672 555
rect 666 550 667 554
rect 671 550 672 554
rect 666 549 672 550
rect 882 554 888 555
rect 882 550 883 554
rect 887 550 888 554
rect 882 549 888 550
rect 1098 554 1104 555
rect 1098 550 1099 554
rect 1103 550 1104 554
rect 1098 549 1104 550
rect 1182 549 1188 550
rect 110 545 111 549
rect 115 545 116 549
rect 110 544 116 545
rect 1182 545 1183 549
rect 1187 545 1188 549
rect 1182 544 1188 545
rect 110 531 116 532
rect 110 527 111 531
rect 115 527 116 531
rect 110 526 116 527
rect 1182 531 1188 532
rect 1182 527 1183 531
rect 1187 527 1188 531
rect 1182 526 1188 527
rect 238 523 244 524
rect 238 522 239 523
rect 193 520 239 522
rect 238 519 239 520
rect 243 519 244 523
rect 398 523 404 524
rect 398 522 399 523
rect 329 520 399 522
rect 238 518 244 519
rect 398 519 399 520
rect 403 519 404 523
rect 594 523 600 524
rect 594 522 595 523
rect 513 520 595 522
rect 398 518 404 519
rect 594 519 595 520
rect 599 519 600 523
rect 594 518 600 519
rect 670 523 676 524
rect 670 519 671 523
rect 675 519 676 523
rect 1167 523 1173 524
rect 1167 522 1168 523
rect 670 518 676 519
rect 728 520 873 522
rect 1145 520 1168 522
rect 215 515 221 516
rect 728 515 730 520
rect 1167 519 1168 520
rect 1172 519 1173 523
rect 1167 518 1173 519
rect 1170 515 1176 516
rect 215 514 216 515
rect 142 513 148 514
rect 142 509 143 513
rect 147 509 148 513
rect 213 512 216 514
rect 215 511 216 512
rect 220 511 221 515
rect 1170 514 1171 515
rect 215 510 221 511
rect 278 513 284 514
rect 142 508 148 509
rect 278 509 279 513
rect 283 509 284 513
rect 462 513 468 514
rect 344 510 346 511
rect 278 508 284 509
rect 340 508 346 510
rect 462 509 463 513
rect 467 509 468 513
rect 662 513 668 514
rect 528 510 530 511
rect 462 508 468 509
rect 524 508 530 510
rect 662 509 663 513
rect 667 509 668 513
rect 662 508 668 509
rect 878 513 884 514
rect 878 509 879 513
rect 883 509 884 513
rect 1094 513 1100 514
rect 878 508 884 509
rect 238 499 244 500
rect 238 495 239 499
rect 243 498 244 499
rect 340 498 342 508
rect 243 496 342 498
rect 398 499 404 500
rect 243 495 244 496
rect 238 494 244 495
rect 398 495 399 499
rect 403 498 404 499
rect 524 498 526 508
rect 403 496 526 498
rect 594 499 600 500
rect 403 495 404 496
rect 398 494 404 495
rect 594 495 595 499
rect 599 498 600 499
rect 944 498 946 511
rect 1094 509 1095 513
rect 1099 509 1100 513
rect 1165 512 1171 514
rect 1170 511 1171 512
rect 1175 511 1176 515
rect 1170 510 1176 511
rect 1094 508 1100 509
rect 599 496 946 498
rect 599 495 600 496
rect 594 494 600 495
rect 740 492 902 494
rect 738 491 744 492
rect 738 487 739 491
rect 743 487 744 491
rect 738 486 744 487
rect 900 486 902 492
rect 1167 487 1173 488
rect 1167 486 1168 487
rect 900 484 906 486
rect 1160 484 1168 486
rect 406 483 412 484
rect 406 479 407 483
rect 411 479 412 483
rect 406 478 412 479
rect 502 483 508 484
rect 502 479 503 483
rect 507 479 508 483
rect 502 478 508 479
rect 606 483 612 484
rect 606 479 607 483
rect 611 479 612 483
rect 606 478 612 479
rect 670 483 676 484
rect 670 479 671 483
rect 675 479 676 483
rect 670 478 676 479
rect 718 483 724 484
rect 718 479 719 483
rect 723 479 724 483
rect 838 483 844 484
rect 718 478 724 479
rect 782 479 788 480
rect 477 476 498 478
rect 573 476 602 478
rect 457 472 490 474
rect 496 473 498 476
rect 600 473 602 476
rect 782 475 783 479
rect 787 475 788 479
rect 838 479 839 483
rect 843 479 844 483
rect 904 481 906 484
rect 966 483 972 484
rect 838 478 844 479
rect 966 479 967 483
rect 971 479 972 483
rect 1094 483 1100 484
rect 966 478 972 479
rect 1030 479 1036 480
rect 782 474 788 475
rect 946 475 952 476
rect 946 474 947 475
rect 889 472 947 474
rect 486 471 492 472
rect 486 467 487 471
rect 491 467 492 471
rect 486 466 492 467
rect 738 471 744 472
rect 738 467 739 471
rect 743 467 744 471
rect 946 471 947 472
rect 951 471 952 475
rect 946 470 952 471
rect 958 475 964 476
rect 958 471 959 475
rect 963 471 964 475
rect 1030 475 1031 479
rect 1035 475 1036 479
rect 1094 479 1095 483
rect 1099 479 1100 483
rect 1160 481 1162 484
rect 1167 483 1168 484
rect 1172 483 1173 487
rect 1167 482 1173 483
rect 1094 478 1100 479
rect 1030 474 1036 475
rect 1167 475 1173 476
rect 1167 474 1168 475
rect 1145 472 1168 474
rect 958 470 964 471
rect 1167 471 1168 472
rect 1172 471 1173 475
rect 1167 470 1173 471
rect 738 466 744 467
rect 110 465 116 466
rect 110 461 111 465
rect 115 461 116 465
rect 110 460 116 461
rect 1182 465 1188 466
rect 1182 461 1183 465
rect 1187 461 1188 465
rect 1182 460 1188 461
rect 110 447 116 448
rect 110 443 111 447
rect 115 443 116 447
rect 1182 447 1188 448
rect 1182 443 1183 447
rect 1187 443 1188 447
rect 110 442 116 443
rect 410 442 416 443
rect 410 438 411 442
rect 415 438 416 442
rect 410 437 416 438
rect 506 442 512 443
rect 506 438 507 442
rect 511 438 512 442
rect 506 437 512 438
rect 610 442 616 443
rect 610 438 611 442
rect 615 438 616 442
rect 610 437 616 438
rect 722 442 728 443
rect 722 438 723 442
rect 727 438 728 442
rect 722 437 728 438
rect 842 442 848 443
rect 842 438 843 442
rect 847 438 848 442
rect 842 437 848 438
rect 970 442 976 443
rect 970 438 971 442
rect 975 438 976 442
rect 970 437 976 438
rect 1098 442 1104 443
rect 1182 442 1188 443
rect 1098 438 1099 442
rect 1103 438 1104 442
rect 1098 437 1104 438
rect 978 419 984 420
rect 978 415 979 419
rect 983 418 984 419
rect 1030 419 1036 420
rect 1030 418 1031 419
rect 983 416 1031 418
rect 983 415 984 416
rect 978 414 984 415
rect 1030 415 1031 416
rect 1035 415 1036 419
rect 1030 414 1036 415
rect 586 398 592 399
rect 586 394 587 398
rect 591 394 592 398
rect 110 393 116 394
rect 586 393 592 394
rect 674 398 680 399
rect 674 394 675 398
rect 679 394 680 398
rect 674 393 680 394
rect 770 398 776 399
rect 770 394 771 398
rect 775 394 776 398
rect 770 393 776 394
rect 874 398 880 399
rect 874 394 875 398
rect 879 394 880 398
rect 874 393 880 394
rect 986 398 992 399
rect 986 394 987 398
rect 991 394 992 398
rect 986 393 992 394
rect 1098 398 1104 399
rect 1098 394 1099 398
rect 1103 394 1104 398
rect 1098 393 1104 394
rect 1182 393 1188 394
rect 110 389 111 393
rect 115 389 116 393
rect 110 388 116 389
rect 1182 389 1183 393
rect 1187 389 1188 393
rect 1182 388 1188 389
rect 946 387 952 388
rect 946 383 947 387
rect 951 386 952 387
rect 951 384 1050 386
rect 951 383 952 384
rect 946 382 952 383
rect 1046 383 1052 384
rect 1046 379 1047 383
rect 1051 379 1052 383
rect 1046 378 1052 379
rect 110 375 116 376
rect 110 371 111 375
rect 115 371 116 375
rect 110 370 116 371
rect 1182 375 1188 376
rect 1182 371 1183 375
rect 1187 371 1188 375
rect 1182 370 1188 371
rect 654 367 660 368
rect 654 366 655 367
rect 633 364 655 366
rect 654 363 655 364
rect 659 363 660 367
rect 1166 367 1172 368
rect 1166 366 1167 367
rect 654 362 660 363
rect 664 358 666 365
rect 736 364 761 366
rect 832 364 865 366
rect 936 364 977 366
rect 1145 364 1167 366
rect 736 359 738 364
rect 832 359 834 364
rect 936 359 938 364
rect 1166 363 1167 364
rect 1171 363 1172 367
rect 1166 362 1172 363
rect 1046 359 1052 360
rect 582 357 588 358
rect 582 353 583 357
rect 587 353 588 357
rect 653 356 666 358
rect 670 357 676 358
rect 582 352 588 353
rect 670 353 671 357
rect 675 353 676 357
rect 670 352 676 353
rect 766 357 772 358
rect 766 353 767 357
rect 771 353 772 357
rect 766 352 772 353
rect 870 357 876 358
rect 870 353 871 357
rect 875 353 876 357
rect 870 352 876 353
rect 982 357 988 358
rect 982 353 983 357
rect 987 353 988 357
rect 1046 355 1047 359
rect 1051 355 1052 359
rect 1167 359 1173 360
rect 1167 358 1168 359
rect 1046 354 1052 355
rect 1094 357 1100 358
rect 982 352 988 353
rect 1094 353 1095 357
rect 1099 353 1100 357
rect 1165 356 1168 358
rect 1167 355 1168 356
rect 1172 355 1173 359
rect 1167 354 1173 355
rect 1094 352 1100 353
rect 414 335 420 336
rect 414 331 415 335
rect 419 331 420 335
rect 414 330 420 331
rect 510 335 516 336
rect 510 331 511 335
rect 515 331 516 335
rect 510 330 516 331
rect 614 335 620 336
rect 614 331 615 335
rect 619 331 620 335
rect 614 330 620 331
rect 726 335 732 336
rect 726 331 727 335
rect 731 331 732 335
rect 726 330 732 331
rect 838 335 844 336
rect 838 331 839 335
rect 843 331 844 335
rect 838 330 844 331
rect 902 335 908 336
rect 902 331 903 335
rect 907 331 908 335
rect 902 330 908 331
rect 958 335 964 336
rect 958 331 959 335
rect 963 331 964 335
rect 1086 335 1092 336
rect 958 330 964 331
rect 1026 331 1032 332
rect 485 328 506 330
rect 581 328 610 330
rect 685 328 722 330
rect 797 328 834 330
rect 465 324 498 326
rect 504 325 506 328
rect 608 325 610 328
rect 720 325 722 328
rect 832 325 834 328
rect 1026 327 1027 331
rect 1031 327 1032 331
rect 1086 331 1087 335
rect 1091 331 1092 335
rect 1086 330 1092 331
rect 1166 331 1172 332
rect 1166 330 1167 331
rect 1157 328 1167 330
rect 1026 326 1032 327
rect 1166 327 1167 328
rect 1171 327 1172 331
rect 1166 326 1172 327
rect 1137 324 1162 326
rect 494 323 500 324
rect 494 319 495 323
rect 499 319 500 323
rect 494 318 500 319
rect 974 323 980 324
rect 974 319 975 323
rect 979 319 980 323
rect 974 318 980 319
rect 1158 323 1164 324
rect 1158 319 1159 323
rect 1163 319 1164 323
rect 1158 318 1164 319
rect 110 317 116 318
rect 110 313 111 317
rect 115 313 116 317
rect 110 312 116 313
rect 1182 317 1188 318
rect 1182 313 1183 317
rect 1187 313 1188 317
rect 1182 312 1188 313
rect 110 299 116 300
rect 110 295 111 299
rect 115 295 116 299
rect 1182 299 1188 300
rect 1182 295 1183 299
rect 1187 295 1188 299
rect 110 294 116 295
rect 418 294 424 295
rect 418 290 419 294
rect 423 290 424 294
rect 418 289 424 290
rect 514 294 520 295
rect 514 290 515 294
rect 519 290 520 294
rect 514 289 520 290
rect 618 294 624 295
rect 618 290 619 294
rect 623 290 624 294
rect 618 289 624 290
rect 730 294 736 295
rect 730 290 731 294
rect 735 290 736 294
rect 730 289 736 290
rect 842 294 848 295
rect 842 290 843 294
rect 847 290 848 294
rect 842 289 848 290
rect 962 294 968 295
rect 962 290 963 294
rect 967 290 968 294
rect 962 289 968 290
rect 1090 294 1096 295
rect 1182 294 1188 295
rect 1090 290 1091 294
rect 1095 290 1096 294
rect 1090 289 1096 290
rect 494 271 500 272
rect 494 267 495 271
rect 499 270 500 271
rect 702 271 708 272
rect 702 270 703 271
rect 499 268 703 270
rect 499 267 500 268
rect 494 266 500 267
rect 702 267 703 268
rect 707 267 708 271
rect 702 266 708 267
rect 863 271 869 272
rect 863 267 864 271
rect 868 270 869 271
rect 1026 271 1032 272
rect 1026 270 1027 271
rect 868 268 1027 270
rect 868 267 869 268
rect 863 266 869 267
rect 1026 267 1027 268
rect 1031 267 1032 271
rect 1026 266 1032 267
rect 202 250 208 251
rect 202 246 203 250
rect 207 246 208 250
rect 110 245 116 246
rect 202 245 208 246
rect 306 250 312 251
rect 306 246 307 250
rect 311 246 312 250
rect 306 245 312 246
rect 418 250 424 251
rect 418 246 419 250
rect 423 246 424 250
rect 418 245 424 246
rect 530 250 536 251
rect 530 246 531 250
rect 535 246 536 250
rect 530 245 536 246
rect 642 250 648 251
rect 642 246 643 250
rect 647 246 648 250
rect 642 245 648 246
rect 762 250 768 251
rect 762 246 763 250
rect 767 246 768 250
rect 762 245 768 246
rect 882 250 888 251
rect 882 246 883 250
rect 887 246 888 250
rect 882 245 888 246
rect 1002 250 1008 251
rect 1002 246 1003 250
rect 1007 246 1008 250
rect 1002 245 1008 246
rect 1098 250 1104 251
rect 1098 246 1099 250
rect 1103 246 1104 250
rect 1098 245 1104 246
rect 1182 245 1188 246
rect 110 241 111 245
rect 115 241 116 245
rect 110 240 116 241
rect 1182 241 1183 245
rect 1187 241 1188 245
rect 1182 240 1188 241
rect 110 227 116 228
rect 110 223 111 227
rect 115 223 116 227
rect 110 222 116 223
rect 1182 227 1188 228
rect 1182 223 1183 227
rect 1187 223 1188 227
rect 1182 222 1188 223
rect 287 219 293 220
rect 287 218 288 219
rect 249 216 288 218
rect 287 215 288 216
rect 292 215 293 219
rect 863 219 869 220
rect 863 218 864 219
rect 287 214 293 215
rect 296 210 298 217
rect 368 216 409 218
rect 480 216 521 218
rect 592 216 633 218
rect 809 216 864 218
rect 368 211 370 216
rect 480 211 482 216
rect 592 211 594 216
rect 863 215 864 216
rect 868 215 869 219
rect 863 214 869 215
rect 702 211 708 212
rect 198 209 204 210
rect 198 205 199 209
rect 203 205 204 209
rect 269 208 298 210
rect 302 209 308 210
rect 198 204 204 205
rect 302 205 303 209
rect 307 205 308 209
rect 302 204 308 205
rect 414 209 420 210
rect 414 205 415 209
rect 419 205 420 209
rect 414 204 420 205
rect 526 209 532 210
rect 526 205 527 209
rect 531 205 532 209
rect 526 204 532 205
rect 638 209 644 210
rect 638 205 639 209
rect 643 205 644 209
rect 702 207 703 211
rect 707 207 708 211
rect 872 210 874 217
rect 944 216 993 218
rect 1064 216 1089 218
rect 944 211 946 216
rect 1064 211 1066 216
rect 1158 211 1164 212
rect 702 206 708 207
rect 758 209 764 210
rect 638 204 644 205
rect 758 205 759 209
rect 763 205 764 209
rect 829 208 874 210
rect 878 209 884 210
rect 758 204 764 205
rect 878 205 879 209
rect 883 205 884 209
rect 878 204 884 205
rect 998 209 1004 210
rect 998 205 999 209
rect 1003 205 1004 209
rect 998 204 1004 205
rect 1094 209 1100 210
rect 1094 205 1095 209
rect 1099 205 1100 209
rect 1158 207 1159 211
rect 1163 207 1164 211
rect 1158 206 1164 207
rect 1094 204 1100 205
rect 287 171 293 172
rect 287 167 288 171
rect 292 170 293 171
rect 292 168 826 170
rect 292 167 293 168
rect 287 166 293 167
rect 142 159 148 160
rect 142 155 143 159
rect 147 155 148 159
rect 142 154 148 155
rect 230 159 236 160
rect 230 155 231 159
rect 235 155 236 159
rect 230 154 236 155
rect 318 159 324 160
rect 318 155 319 159
rect 323 155 324 159
rect 318 154 324 155
rect 406 159 412 160
rect 406 155 407 159
rect 411 155 412 159
rect 406 154 412 155
rect 494 159 500 160
rect 494 155 495 159
rect 499 155 500 159
rect 494 154 500 155
rect 582 159 588 160
rect 582 155 583 159
rect 587 155 588 159
rect 582 154 588 155
rect 670 159 676 160
rect 670 155 671 159
rect 675 155 676 159
rect 670 154 676 155
rect 758 159 764 160
rect 758 155 759 159
rect 763 155 764 159
rect 824 157 826 168
rect 758 154 764 155
rect 213 152 226 154
rect 301 152 314 154
rect 389 152 402 154
rect 477 152 490 154
rect 565 152 578 154
rect 653 152 666 154
rect 741 152 754 154
rect 224 149 226 152
rect 312 149 314 152
rect 400 149 402 152
rect 488 149 490 152
rect 576 149 578 152
rect 664 149 666 152
rect 752 149 754 152
rect 110 141 116 142
rect 110 137 111 141
rect 115 137 116 141
rect 110 136 116 137
rect 1182 141 1188 142
rect 1182 137 1183 141
rect 1187 137 1188 141
rect 1182 136 1188 137
rect 110 123 116 124
rect 110 119 111 123
rect 115 119 116 123
rect 1182 123 1188 124
rect 1182 119 1183 123
rect 1187 119 1188 123
rect 110 118 116 119
rect 146 118 152 119
rect 146 114 147 118
rect 151 114 152 118
rect 146 113 152 114
rect 234 118 240 119
rect 234 114 235 118
rect 239 114 240 118
rect 234 113 240 114
rect 322 118 328 119
rect 322 114 323 118
rect 327 114 328 118
rect 322 113 328 114
rect 410 118 416 119
rect 410 114 411 118
rect 415 114 416 118
rect 410 113 416 114
rect 498 118 504 119
rect 498 114 499 118
rect 503 114 504 118
rect 498 113 504 114
rect 586 118 592 119
rect 586 114 587 118
rect 591 114 592 118
rect 586 113 592 114
rect 674 118 680 119
rect 674 114 675 118
rect 679 114 680 118
rect 674 113 680 114
rect 762 118 768 119
rect 1182 118 1188 119
rect 762 114 763 118
rect 767 114 768 118
rect 762 113 768 114
<< m3c >>
rect 663 1271 667 1275
rect 751 1271 755 1275
rect 839 1271 843 1275
rect 927 1271 931 1275
rect 991 1267 995 1271
rect 111 1253 115 1257
rect 1183 1253 1187 1257
rect 111 1235 115 1239
rect 1183 1235 1187 1239
rect 667 1230 671 1234
rect 755 1230 759 1234
rect 843 1230 847 1234
rect 931 1230 935 1234
rect 371 1190 375 1194
rect 459 1190 463 1194
rect 555 1190 559 1194
rect 651 1190 655 1194
rect 755 1190 759 1194
rect 859 1190 863 1194
rect 963 1190 967 1194
rect 111 1185 115 1189
rect 1183 1185 1187 1189
rect 815 1175 819 1179
rect 111 1167 115 1171
rect 1183 1167 1187 1171
rect 439 1159 443 1163
rect 935 1159 939 1163
rect 983 1159 987 1163
rect 367 1149 371 1153
rect 455 1149 459 1153
rect 551 1149 555 1153
rect 647 1149 651 1153
rect 751 1149 755 1153
rect 815 1151 819 1155
rect 855 1149 859 1153
rect 923 1151 927 1155
rect 959 1149 963 1153
rect 935 1135 939 1139
rect 143 1119 147 1123
rect 255 1119 259 1123
rect 415 1119 419 1123
rect 583 1119 587 1123
rect 767 1119 771 1123
rect 831 1119 835 1123
rect 951 1119 955 1123
rect 215 1107 219 1111
rect 923 1111 927 1115
rect 1015 1115 1019 1119
rect 111 1101 115 1105
rect 1183 1101 1187 1105
rect 111 1083 115 1087
rect 1183 1083 1187 1087
rect 147 1078 151 1082
rect 259 1078 263 1082
rect 419 1078 423 1082
rect 587 1078 591 1082
rect 771 1078 775 1082
rect 955 1078 959 1082
rect 155 1022 159 1026
rect 283 1022 287 1026
rect 427 1022 431 1026
rect 587 1022 591 1026
rect 755 1022 759 1026
rect 939 1022 943 1026
rect 1099 1022 1103 1026
rect 111 1017 115 1021
rect 1183 1017 1187 1021
rect 111 999 115 1003
rect 1183 999 1187 1003
rect 379 991 383 995
rect 543 991 547 995
rect 763 991 767 995
rect 1015 991 1019 995
rect 151 981 155 985
rect 215 983 219 987
rect 279 981 283 985
rect 423 981 427 985
rect 583 981 587 985
rect 751 981 755 985
rect 379 967 383 971
rect 543 967 547 971
rect 935 981 939 985
rect 991 975 995 979
rect 1095 981 1099 985
rect 811 959 815 963
rect 503 951 507 955
rect 591 951 595 955
rect 687 951 691 955
rect 763 947 767 951
rect 791 951 795 955
rect 855 947 859 951
rect 895 951 899 955
rect 1007 951 1011 955
rect 1095 951 1099 955
rect 575 939 579 943
rect 811 939 815 943
rect 983 943 987 947
rect 1079 939 1083 943
rect 111 933 115 937
rect 1183 933 1187 937
rect 111 915 115 919
rect 1183 915 1187 919
rect 507 910 511 914
rect 595 910 599 914
rect 691 910 695 914
rect 795 910 799 914
rect 899 910 903 914
rect 1011 910 1015 914
rect 1099 910 1103 914
rect 1079 883 1083 887
rect 1159 883 1163 887
rect 563 862 567 866
rect 651 862 655 866
rect 739 862 743 866
rect 827 862 831 866
rect 923 862 927 866
rect 111 857 115 861
rect 991 859 995 863
rect 1011 862 1015 866
rect 1099 862 1103 866
rect 1183 857 1187 861
rect 111 839 115 843
rect 1183 839 1187 843
rect 631 831 635 835
rect 559 821 563 825
rect 647 821 651 825
rect 735 821 739 825
rect 823 821 827 825
rect 919 821 923 825
rect 983 823 987 827
rect 1007 821 1011 825
rect 1095 821 1099 825
rect 1159 823 1163 827
rect 999 807 1003 811
rect 391 783 395 787
rect 495 783 499 787
rect 607 783 611 787
rect 727 783 731 787
rect 855 783 859 787
rect 919 779 923 783
rect 983 783 987 787
rect 1047 779 1051 783
rect 1095 783 1099 787
rect 479 771 483 775
rect 999 771 1003 775
rect 1119 771 1123 775
rect 111 765 115 769
rect 1183 765 1187 769
rect 111 747 115 751
rect 1183 747 1187 751
rect 395 742 399 746
rect 499 742 503 746
rect 611 742 615 746
rect 731 742 735 746
rect 859 742 863 746
rect 987 742 991 746
rect 1099 742 1103 746
rect 1123 719 1127 723
rect 1171 719 1175 723
rect 211 698 215 702
rect 355 698 359 702
rect 523 698 527 702
rect 715 698 719 702
rect 915 698 919 702
rect 1099 698 1103 702
rect 111 693 115 697
rect 1183 693 1187 697
rect 111 675 115 679
rect 1183 675 1187 679
rect 335 667 339 671
rect 207 657 211 661
rect 351 657 355 661
rect 519 657 523 661
rect 711 657 715 661
rect 911 657 915 661
rect 479 643 483 647
rect 1095 657 1099 661
rect 1171 659 1175 663
rect 143 631 147 635
rect 295 631 299 635
rect 487 631 491 635
rect 687 631 691 635
rect 751 631 755 635
rect 895 631 899 635
rect 959 631 963 635
rect 1095 631 1099 635
rect 1047 623 1051 627
rect 1171 619 1175 623
rect 111 613 115 617
rect 1183 613 1187 617
rect 111 595 115 599
rect 1183 595 1187 599
rect 147 590 151 594
rect 299 590 303 594
rect 491 590 495 594
rect 691 590 695 594
rect 899 590 903 594
rect 1099 590 1103 594
rect 147 550 151 554
rect 283 550 287 554
rect 467 550 471 554
rect 667 550 671 554
rect 883 550 887 554
rect 1099 550 1103 554
rect 111 545 115 549
rect 1183 545 1187 549
rect 111 527 115 531
rect 1183 527 1187 531
rect 239 519 243 523
rect 399 519 403 523
rect 595 519 599 523
rect 671 519 675 523
rect 143 509 147 513
rect 279 509 283 513
rect 463 509 467 513
rect 663 509 667 513
rect 879 509 883 513
rect 239 495 243 499
rect 399 495 403 499
rect 595 495 599 499
rect 1095 509 1099 513
rect 1171 511 1175 515
rect 739 487 743 491
rect 407 479 411 483
rect 503 479 507 483
rect 607 479 611 483
rect 671 479 675 483
rect 719 479 723 483
rect 783 475 787 479
rect 839 479 843 483
rect 967 479 971 483
rect 487 467 491 471
rect 739 467 743 471
rect 947 471 951 475
rect 959 471 963 475
rect 1031 475 1035 479
rect 1095 479 1099 483
rect 111 461 115 465
rect 1183 461 1187 465
rect 111 443 115 447
rect 1183 443 1187 447
rect 411 438 415 442
rect 507 438 511 442
rect 611 438 615 442
rect 723 438 727 442
rect 843 438 847 442
rect 971 438 975 442
rect 1099 438 1103 442
rect 979 415 983 419
rect 1031 415 1035 419
rect 587 394 591 398
rect 675 394 679 398
rect 771 394 775 398
rect 875 394 879 398
rect 987 394 991 398
rect 1099 394 1103 398
rect 111 389 115 393
rect 1183 389 1187 393
rect 947 383 951 387
rect 1047 379 1051 383
rect 111 371 115 375
rect 1183 371 1187 375
rect 655 363 659 367
rect 1167 363 1171 367
rect 583 353 587 357
rect 671 353 675 357
rect 767 353 771 357
rect 871 353 875 357
rect 983 353 987 357
rect 1047 355 1051 359
rect 1095 353 1099 357
rect 415 331 419 335
rect 511 331 515 335
rect 615 331 619 335
rect 727 331 731 335
rect 839 331 843 335
rect 903 331 907 335
rect 959 331 963 335
rect 1027 327 1031 331
rect 1087 331 1091 335
rect 1167 327 1171 331
rect 495 319 499 323
rect 975 319 979 323
rect 1159 319 1163 323
rect 111 313 115 317
rect 1183 313 1187 317
rect 111 295 115 299
rect 1183 295 1187 299
rect 419 290 423 294
rect 515 290 519 294
rect 619 290 623 294
rect 731 290 735 294
rect 843 290 847 294
rect 963 290 967 294
rect 1091 290 1095 294
rect 495 267 499 271
rect 703 267 707 271
rect 1027 267 1031 271
rect 203 246 207 250
rect 307 246 311 250
rect 419 246 423 250
rect 531 246 535 250
rect 643 246 647 250
rect 763 246 767 250
rect 883 246 887 250
rect 1003 246 1007 250
rect 1099 246 1103 250
rect 111 241 115 245
rect 1183 241 1187 245
rect 111 223 115 227
rect 1183 223 1187 227
rect 199 205 203 209
rect 303 205 307 209
rect 415 205 419 209
rect 527 205 531 209
rect 639 205 643 209
rect 703 207 707 211
rect 759 205 763 209
rect 879 205 883 209
rect 999 205 1003 209
rect 1095 205 1099 209
rect 1159 207 1163 211
rect 143 155 147 159
rect 231 155 235 159
rect 319 155 323 159
rect 407 155 411 159
rect 495 155 499 159
rect 583 155 587 159
rect 671 155 675 159
rect 759 155 763 159
rect 111 137 115 141
rect 1183 137 1187 141
rect 111 119 115 123
rect 1183 119 1187 123
rect 147 114 151 118
rect 235 114 239 118
rect 323 114 327 118
rect 411 114 415 118
rect 499 114 503 118
rect 587 114 591 118
rect 675 114 679 118
rect 763 114 767 118
<< m3 >>
rect 111 1286 115 1287
rect 111 1281 115 1282
rect 663 1286 667 1287
rect 663 1281 667 1282
rect 751 1286 755 1287
rect 751 1281 755 1282
rect 839 1286 843 1287
rect 839 1281 843 1282
rect 927 1286 931 1287
rect 927 1281 931 1282
rect 1183 1286 1187 1287
rect 1183 1281 1187 1282
rect 112 1258 114 1281
rect 664 1276 666 1281
rect 752 1276 754 1281
rect 840 1276 842 1281
rect 928 1276 930 1281
rect 662 1275 668 1276
rect 662 1271 663 1275
rect 667 1271 668 1275
rect 662 1270 668 1271
rect 750 1275 756 1276
rect 750 1271 751 1275
rect 755 1271 756 1275
rect 750 1270 756 1271
rect 838 1275 844 1276
rect 838 1271 839 1275
rect 843 1271 844 1275
rect 838 1270 844 1271
rect 926 1275 932 1276
rect 926 1271 927 1275
rect 931 1271 932 1275
rect 926 1270 932 1271
rect 990 1271 996 1272
rect 990 1267 991 1271
rect 995 1267 996 1271
rect 990 1266 996 1267
rect 110 1257 116 1258
rect 110 1253 111 1257
rect 115 1253 116 1257
rect 110 1252 116 1253
rect 110 1239 116 1240
rect 110 1235 111 1239
rect 115 1235 116 1239
rect 110 1234 116 1235
rect 666 1234 672 1235
rect 112 1215 114 1234
rect 666 1230 667 1234
rect 671 1230 672 1234
rect 666 1229 672 1230
rect 754 1234 760 1235
rect 754 1230 755 1234
rect 759 1230 760 1234
rect 754 1229 760 1230
rect 842 1234 848 1235
rect 842 1230 843 1234
rect 847 1230 848 1234
rect 842 1229 848 1230
rect 930 1234 936 1235
rect 930 1230 931 1234
rect 935 1230 936 1234
rect 930 1229 936 1230
rect 668 1215 670 1229
rect 756 1215 758 1229
rect 844 1215 846 1229
rect 932 1215 934 1229
rect 992 1219 994 1266
rect 1184 1258 1186 1281
rect 1182 1257 1188 1258
rect 1182 1253 1183 1257
rect 1187 1253 1188 1257
rect 1182 1252 1188 1253
rect 1182 1239 1188 1240
rect 1182 1235 1183 1239
rect 1187 1235 1188 1239
rect 1182 1234 1188 1235
rect 984 1217 994 1219
rect 111 1214 115 1215
rect 111 1209 115 1210
rect 371 1214 375 1215
rect 371 1209 375 1210
rect 459 1214 463 1215
rect 459 1209 463 1210
rect 555 1214 559 1215
rect 555 1209 559 1210
rect 651 1214 655 1215
rect 651 1209 655 1210
rect 667 1214 671 1215
rect 667 1209 671 1210
rect 755 1214 759 1215
rect 755 1209 759 1210
rect 843 1214 847 1215
rect 843 1209 847 1210
rect 859 1214 863 1215
rect 859 1209 863 1210
rect 931 1214 935 1215
rect 931 1209 935 1210
rect 963 1214 967 1215
rect 963 1209 967 1210
rect 112 1190 114 1209
rect 372 1195 374 1209
rect 460 1195 462 1209
rect 556 1195 558 1209
rect 652 1195 654 1209
rect 756 1195 758 1209
rect 860 1195 862 1209
rect 964 1195 966 1209
rect 370 1194 376 1195
rect 370 1190 371 1194
rect 375 1190 376 1194
rect 110 1189 116 1190
rect 370 1189 376 1190
rect 458 1194 464 1195
rect 458 1190 459 1194
rect 463 1190 464 1194
rect 458 1189 464 1190
rect 554 1194 560 1195
rect 554 1190 555 1194
rect 559 1190 560 1194
rect 554 1189 560 1190
rect 650 1194 656 1195
rect 650 1190 651 1194
rect 655 1190 656 1194
rect 650 1189 656 1190
rect 754 1194 760 1195
rect 754 1190 755 1194
rect 759 1190 760 1194
rect 754 1189 760 1190
rect 858 1194 864 1195
rect 858 1190 859 1194
rect 863 1190 864 1194
rect 858 1189 864 1190
rect 962 1194 968 1195
rect 962 1190 963 1194
rect 967 1190 968 1194
rect 962 1189 968 1190
rect 110 1185 111 1189
rect 115 1185 116 1189
rect 110 1184 116 1185
rect 814 1179 820 1180
rect 814 1175 815 1179
rect 819 1175 820 1179
rect 814 1174 820 1175
rect 110 1171 116 1172
rect 110 1167 111 1171
rect 115 1167 116 1171
rect 110 1166 116 1167
rect 112 1135 114 1166
rect 438 1163 444 1164
rect 438 1159 439 1163
rect 443 1159 444 1163
rect 438 1158 444 1159
rect 366 1153 372 1154
rect 366 1149 367 1153
rect 371 1149 372 1153
rect 366 1148 372 1149
rect 368 1135 370 1148
rect 111 1134 115 1135
rect 111 1129 115 1130
rect 143 1134 147 1135
rect 143 1129 147 1130
rect 255 1134 259 1135
rect 255 1129 259 1130
rect 367 1134 371 1135
rect 367 1129 371 1130
rect 415 1134 419 1135
rect 415 1129 419 1130
rect 112 1106 114 1129
rect 144 1124 146 1129
rect 256 1124 258 1129
rect 416 1124 418 1129
rect 440 1125 442 1158
rect 816 1156 818 1174
rect 984 1164 986 1217
rect 1184 1215 1186 1234
rect 1183 1214 1187 1215
rect 1183 1209 1187 1210
rect 1184 1190 1186 1209
rect 1182 1189 1188 1190
rect 1182 1185 1183 1189
rect 1187 1185 1188 1189
rect 1182 1184 1188 1185
rect 1182 1171 1188 1172
rect 1182 1167 1183 1171
rect 1187 1167 1188 1171
rect 1182 1166 1188 1167
rect 934 1163 940 1164
rect 934 1159 935 1163
rect 939 1159 940 1163
rect 934 1158 940 1159
rect 982 1163 988 1164
rect 982 1159 983 1163
rect 987 1159 988 1163
rect 982 1158 988 1159
rect 814 1155 820 1156
rect 454 1153 460 1154
rect 454 1149 455 1153
rect 459 1149 460 1153
rect 454 1148 460 1149
rect 550 1153 556 1154
rect 550 1149 551 1153
rect 555 1149 556 1153
rect 550 1148 556 1149
rect 646 1153 652 1154
rect 646 1149 647 1153
rect 651 1149 652 1153
rect 646 1148 652 1149
rect 750 1153 756 1154
rect 750 1149 751 1153
rect 755 1149 756 1153
rect 814 1151 815 1155
rect 819 1151 820 1155
rect 922 1155 928 1156
rect 814 1150 820 1151
rect 854 1153 860 1154
rect 750 1148 756 1149
rect 854 1149 855 1153
rect 859 1149 860 1153
rect 922 1151 923 1155
rect 927 1151 928 1155
rect 922 1150 928 1151
rect 854 1148 860 1149
rect 456 1135 458 1148
rect 552 1135 554 1148
rect 648 1135 650 1148
rect 752 1135 754 1148
rect 856 1135 858 1148
rect 455 1134 459 1135
rect 455 1129 459 1130
rect 551 1134 555 1135
rect 551 1129 555 1130
rect 583 1134 587 1135
rect 583 1129 587 1130
rect 647 1134 651 1135
rect 647 1129 651 1130
rect 751 1134 755 1135
rect 751 1129 755 1130
rect 767 1134 771 1135
rect 767 1129 771 1130
rect 855 1134 859 1135
rect 855 1129 859 1130
rect 439 1124 443 1125
rect 584 1124 586 1129
rect 768 1124 770 1129
rect 831 1124 835 1125
rect 142 1123 148 1124
rect 142 1119 143 1123
rect 147 1119 148 1123
rect 142 1118 148 1119
rect 254 1123 260 1124
rect 254 1119 255 1123
rect 259 1119 260 1123
rect 254 1118 260 1119
rect 414 1123 420 1124
rect 414 1119 415 1123
rect 419 1119 420 1123
rect 439 1119 443 1120
rect 582 1123 588 1124
rect 582 1119 583 1123
rect 587 1119 588 1123
rect 414 1118 420 1119
rect 582 1118 588 1119
rect 766 1123 772 1124
rect 766 1119 767 1123
rect 771 1119 772 1123
rect 766 1118 772 1119
rect 830 1119 831 1124
rect 835 1119 836 1124
rect 830 1118 836 1119
rect 924 1116 926 1150
rect 936 1140 938 1158
rect 958 1153 964 1154
rect 958 1149 959 1153
rect 963 1149 964 1153
rect 958 1148 964 1149
rect 934 1139 940 1140
rect 934 1135 935 1139
rect 939 1135 940 1139
rect 960 1135 962 1148
rect 1184 1135 1186 1166
rect 934 1134 940 1135
rect 951 1134 955 1135
rect 951 1129 955 1130
rect 959 1134 963 1135
rect 959 1129 963 1130
rect 1183 1134 1187 1135
rect 1183 1129 1187 1130
rect 952 1124 954 1129
rect 950 1123 956 1124
rect 950 1119 951 1123
rect 955 1119 956 1123
rect 950 1118 956 1119
rect 1014 1119 1020 1120
rect 922 1115 928 1116
rect 214 1111 220 1112
rect 214 1107 215 1111
rect 219 1107 220 1111
rect 922 1111 923 1115
rect 927 1111 928 1115
rect 1014 1115 1015 1119
rect 1019 1115 1020 1119
rect 1014 1114 1020 1115
rect 922 1110 928 1111
rect 214 1106 220 1107
rect 110 1105 116 1106
rect 110 1101 111 1105
rect 115 1101 116 1105
rect 110 1100 116 1101
rect 110 1087 116 1088
rect 110 1083 111 1087
rect 115 1083 116 1087
rect 110 1082 116 1083
rect 146 1082 152 1083
rect 112 1047 114 1082
rect 146 1078 147 1082
rect 151 1078 152 1082
rect 146 1077 152 1078
rect 148 1047 150 1077
rect 111 1046 115 1047
rect 111 1041 115 1042
rect 147 1046 151 1047
rect 147 1041 151 1042
rect 155 1046 159 1047
rect 155 1041 159 1042
rect 112 1022 114 1041
rect 156 1027 158 1041
rect 154 1026 160 1027
rect 154 1022 155 1026
rect 159 1022 160 1026
rect 110 1021 116 1022
rect 154 1021 160 1022
rect 110 1017 111 1021
rect 115 1017 116 1021
rect 110 1016 116 1017
rect 110 1003 116 1004
rect 110 999 111 1003
rect 115 999 116 1003
rect 110 998 116 999
rect 112 967 114 998
rect 216 988 218 1106
rect 258 1082 264 1083
rect 258 1078 259 1082
rect 263 1078 264 1082
rect 258 1077 264 1078
rect 418 1082 424 1083
rect 418 1078 419 1082
rect 423 1078 424 1082
rect 418 1077 424 1078
rect 586 1082 592 1083
rect 586 1078 587 1082
rect 591 1078 592 1082
rect 586 1077 592 1078
rect 770 1082 776 1083
rect 770 1078 771 1082
rect 775 1078 776 1082
rect 770 1077 776 1078
rect 954 1082 960 1083
rect 954 1078 955 1082
rect 959 1078 960 1082
rect 954 1077 960 1078
rect 260 1047 262 1077
rect 420 1047 422 1077
rect 588 1047 590 1077
rect 772 1047 774 1077
rect 956 1047 958 1077
rect 259 1046 263 1047
rect 259 1041 263 1042
rect 283 1046 287 1047
rect 283 1041 287 1042
rect 419 1046 423 1047
rect 419 1041 423 1042
rect 427 1046 431 1047
rect 427 1041 431 1042
rect 587 1046 591 1047
rect 587 1041 591 1042
rect 755 1046 759 1047
rect 755 1041 759 1042
rect 771 1046 775 1047
rect 771 1041 775 1042
rect 939 1046 943 1047
rect 939 1041 943 1042
rect 955 1046 959 1047
rect 955 1041 959 1042
rect 284 1027 286 1041
rect 428 1027 430 1041
rect 588 1027 590 1041
rect 756 1027 758 1041
rect 940 1027 942 1041
rect 282 1026 288 1027
rect 282 1022 283 1026
rect 287 1022 288 1026
rect 282 1021 288 1022
rect 426 1026 432 1027
rect 426 1022 427 1026
rect 431 1022 432 1026
rect 426 1021 432 1022
rect 586 1026 592 1027
rect 586 1022 587 1026
rect 591 1022 592 1026
rect 586 1021 592 1022
rect 754 1026 760 1027
rect 754 1022 755 1026
rect 759 1022 760 1026
rect 754 1021 760 1022
rect 938 1026 944 1027
rect 938 1022 939 1026
rect 943 1022 944 1026
rect 938 1021 944 1022
rect 1016 996 1018 1114
rect 1184 1106 1186 1129
rect 1182 1105 1188 1106
rect 1182 1101 1183 1105
rect 1187 1101 1188 1105
rect 1182 1100 1188 1101
rect 1182 1087 1188 1088
rect 1182 1083 1183 1087
rect 1187 1083 1188 1087
rect 1182 1082 1188 1083
rect 1184 1047 1186 1082
rect 1099 1046 1103 1047
rect 1099 1041 1103 1042
rect 1183 1046 1187 1047
rect 1183 1041 1187 1042
rect 1100 1027 1102 1041
rect 1098 1026 1104 1027
rect 1098 1022 1099 1026
rect 1103 1022 1104 1026
rect 1184 1022 1186 1041
rect 1098 1021 1104 1022
rect 1182 1021 1188 1022
rect 1182 1017 1183 1021
rect 1187 1017 1188 1021
rect 1182 1016 1188 1017
rect 1182 1003 1188 1004
rect 1182 999 1183 1003
rect 1187 999 1188 1003
rect 1182 998 1188 999
rect 378 995 384 996
rect 378 991 379 995
rect 383 991 384 995
rect 378 990 384 991
rect 542 995 548 996
rect 542 991 543 995
rect 547 991 548 995
rect 542 990 548 991
rect 762 995 768 996
rect 762 991 763 995
rect 767 991 768 995
rect 762 990 768 991
rect 1014 995 1020 996
rect 1014 991 1015 995
rect 1019 991 1020 995
rect 1014 990 1020 991
rect 214 987 220 988
rect 150 985 156 986
rect 150 981 151 985
rect 155 981 156 985
rect 214 983 215 987
rect 219 983 220 987
rect 214 982 220 983
rect 278 985 284 986
rect 150 980 156 981
rect 278 981 279 985
rect 283 981 284 985
rect 278 980 284 981
rect 152 967 154 980
rect 280 967 282 980
rect 380 972 382 990
rect 422 985 428 986
rect 422 981 423 985
rect 427 981 428 985
rect 422 980 428 981
rect 378 971 384 972
rect 378 967 379 971
rect 383 967 384 971
rect 424 967 426 980
rect 544 972 546 990
rect 582 985 588 986
rect 582 981 583 985
rect 587 981 588 985
rect 582 980 588 981
rect 750 985 756 986
rect 750 981 751 985
rect 755 981 756 985
rect 750 980 756 981
rect 542 971 548 972
rect 542 967 543 971
rect 547 967 548 971
rect 584 967 586 980
rect 752 967 754 980
rect 111 966 115 967
rect 111 961 115 962
rect 151 966 155 967
rect 151 961 155 962
rect 279 966 283 967
rect 378 966 384 967
rect 423 966 427 967
rect 279 961 283 962
rect 423 961 427 962
rect 503 966 507 967
rect 542 966 548 967
rect 583 966 587 967
rect 503 961 507 962
rect 583 961 587 962
rect 591 966 595 967
rect 591 961 595 962
rect 687 966 691 967
rect 687 961 691 962
rect 751 966 755 967
rect 751 961 755 962
rect 112 938 114 961
rect 504 956 506 961
rect 592 956 594 961
rect 688 956 690 961
rect 502 955 508 956
rect 502 951 503 955
rect 507 951 508 955
rect 502 950 508 951
rect 590 955 596 956
rect 590 951 591 955
rect 595 951 596 955
rect 590 950 596 951
rect 686 955 692 956
rect 686 951 687 955
rect 691 951 692 955
rect 764 952 766 990
rect 934 985 940 986
rect 934 981 935 985
rect 939 981 940 985
rect 934 980 940 981
rect 1094 985 1100 986
rect 1094 981 1095 985
rect 1099 981 1100 985
rect 1094 980 1100 981
rect 936 967 938 980
rect 990 979 996 980
rect 990 975 991 979
rect 995 975 996 979
rect 990 974 996 975
rect 791 966 795 967
rect 895 966 899 967
rect 791 961 795 962
rect 810 963 816 964
rect 792 956 794 961
rect 810 959 811 963
rect 815 959 816 963
rect 895 961 899 962
rect 935 966 939 967
rect 935 961 939 962
rect 810 958 816 959
rect 790 955 796 956
rect 686 950 692 951
rect 762 951 768 952
rect 575 948 579 949
rect 762 947 763 951
rect 767 947 768 951
rect 790 951 791 955
rect 795 951 796 955
rect 790 950 796 951
rect 762 946 768 947
rect 812 944 814 958
rect 896 956 898 961
rect 894 955 900 956
rect 854 951 860 952
rect 854 946 855 951
rect 859 946 860 951
rect 894 951 895 955
rect 899 951 900 955
rect 894 950 900 951
rect 982 947 988 948
rect 574 943 580 944
rect 574 939 575 943
rect 579 939 580 943
rect 574 938 580 939
rect 810 943 816 944
rect 855 943 859 944
rect 982 943 983 947
rect 987 943 988 947
rect 810 939 811 943
rect 815 939 816 943
rect 982 942 988 943
rect 810 938 816 939
rect 110 937 116 938
rect 110 933 111 937
rect 115 933 116 937
rect 110 932 116 933
rect 110 919 116 920
rect 110 915 111 919
rect 115 915 116 919
rect 110 914 116 915
rect 506 914 512 915
rect 112 887 114 914
rect 506 910 507 914
rect 511 910 512 914
rect 506 909 512 910
rect 594 914 600 915
rect 594 910 595 914
rect 599 910 600 914
rect 594 909 600 910
rect 690 914 696 915
rect 690 910 691 914
rect 695 910 696 914
rect 690 909 696 910
rect 794 914 800 915
rect 794 910 795 914
rect 799 910 800 914
rect 794 909 800 910
rect 898 914 904 915
rect 898 910 899 914
rect 903 910 904 914
rect 898 909 904 910
rect 508 887 510 909
rect 596 887 598 909
rect 692 887 694 909
rect 796 887 798 909
rect 900 887 902 909
rect 111 886 115 887
rect 111 881 115 882
rect 507 886 511 887
rect 507 881 511 882
rect 563 886 567 887
rect 563 881 567 882
rect 595 886 599 887
rect 595 881 599 882
rect 651 886 655 887
rect 651 881 655 882
rect 691 886 695 887
rect 691 881 695 882
rect 739 886 743 887
rect 739 881 743 882
rect 795 886 799 887
rect 795 881 799 882
rect 827 886 831 887
rect 827 881 831 882
rect 899 886 903 887
rect 899 881 903 882
rect 923 886 927 887
rect 923 881 927 882
rect 112 862 114 881
rect 564 867 566 881
rect 652 867 654 881
rect 740 867 742 881
rect 828 867 830 881
rect 924 867 926 881
rect 562 866 568 867
rect 562 862 563 866
rect 567 862 568 866
rect 110 861 116 862
rect 562 861 568 862
rect 650 866 656 867
rect 650 862 651 866
rect 655 862 656 866
rect 650 861 656 862
rect 738 866 744 867
rect 738 862 739 866
rect 743 862 744 866
rect 738 861 744 862
rect 826 866 832 867
rect 826 862 827 866
rect 831 862 832 866
rect 826 861 832 862
rect 922 866 928 867
rect 922 862 923 866
rect 927 862 928 866
rect 922 861 928 862
rect 110 857 111 861
rect 115 857 116 861
rect 110 856 116 857
rect 110 843 116 844
rect 110 839 111 843
rect 115 839 116 843
rect 110 838 116 839
rect 112 799 114 838
rect 630 835 636 836
rect 630 831 631 835
rect 635 831 636 835
rect 630 830 636 831
rect 558 825 564 826
rect 558 821 559 825
rect 563 821 564 825
rect 558 820 564 821
rect 560 799 562 820
rect 111 798 115 799
rect 111 793 115 794
rect 391 798 395 799
rect 391 793 395 794
rect 495 798 499 799
rect 495 793 499 794
rect 559 798 563 799
rect 559 793 563 794
rect 607 798 611 799
rect 607 793 611 794
rect 112 770 114 793
rect 392 788 394 793
rect 496 788 498 793
rect 608 788 610 793
rect 390 787 396 788
rect 390 783 391 787
rect 395 783 396 787
rect 390 782 396 783
rect 494 787 500 788
rect 494 783 495 787
rect 499 783 500 787
rect 494 782 500 783
rect 606 787 612 788
rect 606 783 607 787
rect 611 783 612 787
rect 606 782 612 783
rect 478 775 484 776
rect 478 771 479 775
rect 483 771 484 775
rect 632 773 634 830
rect 984 828 986 942
rect 992 864 994 974
rect 1096 967 1098 980
rect 1184 967 1186 998
rect 1007 966 1011 967
rect 1007 961 1011 962
rect 1095 966 1099 967
rect 1095 961 1099 962
rect 1183 966 1187 967
rect 1183 961 1187 962
rect 1008 956 1010 961
rect 1096 956 1098 961
rect 1006 955 1012 956
rect 1006 951 1007 955
rect 1011 951 1012 955
rect 1006 950 1012 951
rect 1094 955 1100 956
rect 1094 951 1095 955
rect 1099 951 1100 955
rect 1094 950 1100 951
rect 1078 943 1084 944
rect 1078 939 1079 943
rect 1083 939 1084 943
rect 1078 938 1084 939
rect 1184 938 1186 961
rect 1010 914 1016 915
rect 1010 910 1011 914
rect 1015 910 1016 914
rect 1010 909 1016 910
rect 1012 887 1014 909
rect 1080 888 1082 938
rect 1182 937 1188 938
rect 1182 933 1183 937
rect 1187 933 1188 937
rect 1182 932 1188 933
rect 1182 919 1188 920
rect 1182 915 1183 919
rect 1187 915 1188 919
rect 1098 914 1104 915
rect 1182 914 1188 915
rect 1098 910 1099 914
rect 1103 910 1104 914
rect 1098 909 1104 910
rect 1078 887 1084 888
rect 1100 887 1102 909
rect 1158 887 1164 888
rect 1184 887 1186 914
rect 1011 886 1015 887
rect 1078 883 1079 887
rect 1083 883 1084 887
rect 1078 882 1084 883
rect 1099 886 1103 887
rect 1158 883 1159 887
rect 1163 883 1164 887
rect 1158 882 1164 883
rect 1183 886 1187 887
rect 1011 881 1015 882
rect 1099 881 1103 882
rect 1012 867 1014 881
rect 1100 867 1102 881
rect 1010 866 1016 867
rect 990 863 996 864
rect 990 859 991 863
rect 995 859 996 863
rect 1010 862 1011 866
rect 1015 862 1016 866
rect 1010 861 1016 862
rect 1098 866 1104 867
rect 1098 862 1099 866
rect 1103 862 1104 866
rect 1098 861 1104 862
rect 990 858 996 859
rect 1160 828 1162 882
rect 1183 881 1187 882
rect 1184 862 1186 881
rect 1182 861 1188 862
rect 1182 857 1183 861
rect 1187 857 1188 861
rect 1182 856 1188 857
rect 1182 843 1188 844
rect 1182 839 1183 843
rect 1187 839 1188 843
rect 1182 838 1188 839
rect 982 827 988 828
rect 646 825 652 826
rect 646 821 647 825
rect 651 821 652 825
rect 646 820 652 821
rect 734 825 740 826
rect 734 821 735 825
rect 739 821 740 825
rect 734 820 740 821
rect 822 825 828 826
rect 822 821 823 825
rect 827 821 828 825
rect 822 820 828 821
rect 918 825 924 826
rect 918 821 919 825
rect 923 821 924 825
rect 982 823 983 827
rect 987 823 988 827
rect 1158 827 1164 828
rect 982 822 988 823
rect 1006 825 1012 826
rect 918 820 924 821
rect 1006 821 1007 825
rect 1011 821 1012 825
rect 1006 820 1012 821
rect 1094 825 1100 826
rect 1094 821 1095 825
rect 1099 821 1100 825
rect 1158 823 1159 827
rect 1163 823 1164 827
rect 1158 822 1164 823
rect 1094 820 1100 821
rect 648 799 650 820
rect 736 799 738 820
rect 824 799 826 820
rect 920 799 922 820
rect 998 811 1004 812
rect 998 807 999 811
rect 1003 807 1004 811
rect 998 806 1004 807
rect 647 798 651 799
rect 647 793 651 794
rect 727 798 731 799
rect 727 793 731 794
rect 735 798 739 799
rect 735 793 739 794
rect 823 798 827 799
rect 823 793 827 794
rect 855 798 859 799
rect 855 793 859 794
rect 919 798 923 799
rect 919 793 923 794
rect 983 798 987 799
rect 983 793 987 794
rect 728 788 730 793
rect 856 788 858 793
rect 984 788 986 793
rect 726 787 732 788
rect 726 783 727 787
rect 731 783 732 787
rect 726 782 732 783
rect 854 787 860 788
rect 854 783 855 787
rect 859 783 860 787
rect 982 787 988 788
rect 854 782 860 783
rect 918 783 924 784
rect 918 779 919 783
rect 923 779 924 783
rect 982 783 983 787
rect 987 783 988 787
rect 982 782 988 783
rect 918 778 924 779
rect 920 773 922 778
rect 1000 776 1002 806
rect 1008 799 1010 820
rect 1096 799 1098 820
rect 1184 799 1186 838
rect 1007 798 1011 799
rect 1007 793 1011 794
rect 1095 798 1099 799
rect 1095 793 1099 794
rect 1183 798 1187 799
rect 1183 793 1187 794
rect 1096 788 1098 793
rect 1094 787 1100 788
rect 1046 783 1052 784
rect 1046 779 1047 783
rect 1051 779 1052 783
rect 1094 783 1095 787
rect 1099 783 1100 787
rect 1094 782 1100 783
rect 1046 778 1052 779
rect 998 775 1004 776
rect 478 770 484 771
rect 631 772 635 773
rect 110 769 116 770
rect 110 765 111 769
rect 115 765 116 769
rect 110 764 116 765
rect 110 751 116 752
rect 110 747 111 751
rect 115 747 116 751
rect 110 746 116 747
rect 394 746 400 747
rect 112 723 114 746
rect 394 742 395 746
rect 399 742 400 746
rect 394 741 400 742
rect 396 723 398 741
rect 111 722 115 723
rect 111 717 115 718
rect 211 722 215 723
rect 211 717 215 718
rect 355 722 359 723
rect 355 717 359 718
rect 395 722 399 723
rect 395 717 399 718
rect 112 698 114 717
rect 212 703 214 717
rect 356 703 358 717
rect 210 702 216 703
rect 210 698 211 702
rect 215 698 216 702
rect 110 697 116 698
rect 210 697 216 698
rect 354 702 360 703
rect 354 698 355 702
rect 359 698 360 702
rect 354 697 360 698
rect 110 693 111 697
rect 115 693 116 697
rect 110 692 116 693
rect 110 679 116 680
rect 110 675 111 679
rect 115 675 116 679
rect 110 674 116 675
rect 112 647 114 674
rect 334 671 340 672
rect 334 667 335 671
rect 339 667 340 671
rect 334 666 340 667
rect 206 661 212 662
rect 206 657 207 661
rect 211 657 212 661
rect 206 656 212 657
rect 208 647 210 656
rect 111 646 115 647
rect 111 641 115 642
rect 143 646 147 647
rect 143 641 147 642
rect 207 646 211 647
rect 207 641 211 642
rect 295 646 299 647
rect 295 641 299 642
rect 112 618 114 641
rect 144 636 146 641
rect 296 636 298 641
rect 336 637 338 666
rect 350 661 356 662
rect 350 657 351 661
rect 355 657 356 661
rect 350 656 356 657
rect 352 647 354 656
rect 480 648 482 770
rect 631 767 635 768
rect 919 772 923 773
rect 998 771 999 775
rect 1003 771 1004 775
rect 998 770 1004 771
rect 919 767 923 768
rect 498 746 504 747
rect 498 742 499 746
rect 503 742 504 746
rect 498 741 504 742
rect 610 746 616 747
rect 610 742 611 746
rect 615 742 616 746
rect 610 741 616 742
rect 730 746 736 747
rect 730 742 731 746
rect 735 742 736 746
rect 730 741 736 742
rect 858 746 864 747
rect 858 742 859 746
rect 863 742 864 746
rect 858 741 864 742
rect 986 746 992 747
rect 986 742 987 746
rect 991 742 992 746
rect 986 741 992 742
rect 500 723 502 741
rect 612 723 614 741
rect 732 723 734 741
rect 860 723 862 741
rect 988 723 990 741
rect 499 722 503 723
rect 499 717 503 718
rect 523 722 527 723
rect 523 717 527 718
rect 611 722 615 723
rect 611 717 615 718
rect 715 722 719 723
rect 715 717 719 718
rect 731 722 735 723
rect 731 717 735 718
rect 859 722 863 723
rect 859 717 863 718
rect 915 722 919 723
rect 915 717 919 718
rect 987 722 991 723
rect 987 717 991 718
rect 524 703 526 717
rect 716 703 718 717
rect 916 703 918 717
rect 522 702 528 703
rect 522 698 523 702
rect 527 698 528 702
rect 522 697 528 698
rect 714 702 720 703
rect 714 698 715 702
rect 719 698 720 702
rect 714 697 720 698
rect 914 702 920 703
rect 914 698 915 702
rect 919 698 920 702
rect 914 697 920 698
rect 518 661 524 662
rect 518 657 519 661
rect 523 657 524 661
rect 518 656 524 657
rect 710 661 716 662
rect 710 657 711 661
rect 715 657 716 661
rect 710 656 716 657
rect 910 661 916 662
rect 910 657 911 661
rect 915 657 916 661
rect 910 656 916 657
rect 478 647 484 648
rect 520 647 522 656
rect 712 647 714 656
rect 912 647 914 656
rect 351 646 355 647
rect 478 643 479 647
rect 483 643 484 647
rect 478 642 484 643
rect 487 646 491 647
rect 351 641 355 642
rect 487 641 491 642
rect 519 646 523 647
rect 519 641 523 642
rect 687 646 691 647
rect 687 641 691 642
rect 711 646 715 647
rect 711 641 715 642
rect 895 646 899 647
rect 895 641 899 642
rect 911 646 915 647
rect 911 641 915 642
rect 335 636 339 637
rect 488 636 490 641
rect 688 636 690 641
rect 751 636 755 637
rect 896 636 898 641
rect 142 635 148 636
rect 142 631 143 635
rect 147 631 148 635
rect 142 630 148 631
rect 294 635 300 636
rect 294 631 295 635
rect 299 631 300 635
rect 335 631 339 632
rect 486 635 492 636
rect 486 631 487 635
rect 491 631 492 635
rect 294 630 300 631
rect 486 630 492 631
rect 686 635 692 636
rect 686 631 687 635
rect 691 631 692 635
rect 686 630 692 631
rect 750 631 751 636
rect 755 631 756 636
rect 750 630 756 631
rect 894 635 900 636
rect 894 631 895 635
rect 899 631 900 635
rect 894 630 900 631
rect 958 635 964 636
rect 958 631 959 635
rect 963 631 964 635
rect 958 630 964 631
rect 110 617 116 618
rect 110 613 111 617
rect 115 613 116 617
rect 110 612 116 613
rect 110 599 116 600
rect 110 595 111 599
rect 115 595 116 599
rect 110 594 116 595
rect 146 594 152 595
rect 112 575 114 594
rect 146 590 147 594
rect 151 590 152 594
rect 146 589 152 590
rect 298 594 304 595
rect 298 590 299 594
rect 303 590 304 594
rect 298 589 304 590
rect 490 594 496 595
rect 490 590 491 594
rect 495 590 496 594
rect 490 589 496 590
rect 690 594 696 595
rect 690 590 691 594
rect 695 590 696 594
rect 690 589 696 590
rect 898 594 904 595
rect 898 590 899 594
rect 903 590 904 594
rect 898 589 904 590
rect 148 575 150 589
rect 300 575 302 589
rect 492 575 494 589
rect 692 575 694 589
rect 900 575 902 589
rect 111 574 115 575
rect 111 569 115 570
rect 147 574 151 575
rect 147 569 151 570
rect 283 574 287 575
rect 283 569 287 570
rect 299 574 303 575
rect 299 569 303 570
rect 467 574 471 575
rect 467 569 471 570
rect 491 574 495 575
rect 491 569 495 570
rect 667 574 671 575
rect 667 569 671 570
rect 691 574 695 575
rect 691 569 695 570
rect 883 574 887 575
rect 883 569 887 570
rect 899 574 903 575
rect 899 569 903 570
rect 112 550 114 569
rect 148 555 150 569
rect 284 555 286 569
rect 468 555 470 569
rect 668 555 670 569
rect 884 555 886 569
rect 146 554 152 555
rect 146 550 147 554
rect 151 550 152 554
rect 110 549 116 550
rect 146 549 152 550
rect 282 554 288 555
rect 282 550 283 554
rect 287 550 288 554
rect 282 549 288 550
rect 466 554 472 555
rect 466 550 467 554
rect 471 550 472 554
rect 466 549 472 550
rect 666 554 672 555
rect 666 550 667 554
rect 671 550 672 554
rect 666 549 672 550
rect 882 554 888 555
rect 882 550 883 554
rect 887 550 888 554
rect 882 549 888 550
rect 110 545 111 549
rect 115 545 116 549
rect 110 544 116 545
rect 110 531 116 532
rect 110 527 111 531
rect 115 527 116 531
rect 110 526 116 527
rect 112 495 114 526
rect 238 523 244 524
rect 238 519 239 523
rect 243 519 244 523
rect 238 518 244 519
rect 398 523 404 524
rect 398 519 399 523
rect 403 519 404 523
rect 398 518 404 519
rect 594 523 600 524
rect 594 519 595 523
rect 599 519 600 523
rect 594 518 600 519
rect 670 523 676 524
rect 670 519 671 523
rect 675 519 676 523
rect 670 518 676 519
rect 142 513 148 514
rect 142 509 143 513
rect 147 509 148 513
rect 142 508 148 509
rect 144 495 146 508
rect 240 500 242 518
rect 278 513 284 514
rect 278 509 279 513
rect 283 509 284 513
rect 278 508 284 509
rect 238 499 244 500
rect 238 495 239 499
rect 243 495 244 499
rect 280 495 282 508
rect 400 500 402 518
rect 462 513 468 514
rect 462 509 463 513
rect 467 509 468 513
rect 462 508 468 509
rect 398 499 404 500
rect 398 495 399 499
rect 403 495 404 499
rect 464 495 466 508
rect 596 500 598 518
rect 662 513 668 514
rect 662 509 663 513
rect 667 509 668 513
rect 662 508 668 509
rect 594 499 600 500
rect 594 495 595 499
rect 599 495 600 499
rect 664 495 666 508
rect 111 494 115 495
rect 111 489 115 490
rect 143 494 147 495
rect 238 494 244 495
rect 279 494 283 495
rect 398 494 404 495
rect 407 494 411 495
rect 143 489 147 490
rect 279 489 283 490
rect 407 489 411 490
rect 463 494 467 495
rect 463 489 467 490
rect 503 494 507 495
rect 594 494 600 495
rect 607 494 611 495
rect 503 489 507 490
rect 607 489 611 490
rect 663 494 667 495
rect 663 489 667 490
rect 112 466 114 489
rect 408 484 410 489
rect 504 484 506 489
rect 608 484 610 489
rect 672 484 674 518
rect 878 513 884 514
rect 878 509 879 513
rect 883 509 884 513
rect 878 508 884 509
rect 880 495 882 508
rect 719 494 723 495
rect 839 494 843 495
rect 719 489 723 490
rect 738 491 744 492
rect 720 484 722 489
rect 738 487 739 491
rect 743 487 744 491
rect 839 489 843 490
rect 879 494 883 495
rect 879 489 883 490
rect 738 486 744 487
rect 406 483 412 484
rect 406 479 407 483
rect 411 479 412 483
rect 406 478 412 479
rect 502 483 508 484
rect 502 479 503 483
rect 507 479 508 483
rect 502 478 508 479
rect 606 483 612 484
rect 606 479 607 483
rect 611 479 612 483
rect 606 478 612 479
rect 670 483 676 484
rect 670 479 671 483
rect 675 479 676 483
rect 670 478 676 479
rect 718 483 724 484
rect 718 479 719 483
rect 723 479 724 483
rect 718 478 724 479
rect 487 476 491 477
rect 740 472 742 486
rect 840 484 842 489
rect 838 483 844 484
rect 782 479 788 480
rect 782 474 783 479
rect 787 474 788 479
rect 838 479 839 483
rect 843 479 844 483
rect 838 478 844 479
rect 960 476 962 630
rect 1048 628 1050 778
rect 1118 775 1124 776
rect 1118 771 1119 775
rect 1123 771 1124 775
rect 1118 770 1124 771
rect 1184 770 1186 793
rect 1098 746 1104 747
rect 1098 742 1099 746
rect 1103 742 1104 746
rect 1098 741 1104 742
rect 1100 723 1102 741
rect 1120 724 1122 770
rect 1182 769 1188 770
rect 1182 765 1183 769
rect 1187 765 1188 769
rect 1182 764 1188 765
rect 1182 751 1188 752
rect 1182 747 1183 751
rect 1187 747 1188 751
rect 1182 746 1188 747
rect 1120 723 1128 724
rect 1099 722 1103 723
rect 1120 721 1123 723
rect 1122 719 1123 721
rect 1127 719 1128 723
rect 1122 718 1128 719
rect 1170 723 1176 724
rect 1184 723 1186 746
rect 1170 719 1171 723
rect 1175 719 1176 723
rect 1170 718 1176 719
rect 1183 722 1187 723
rect 1099 717 1103 718
rect 1100 703 1102 717
rect 1098 702 1104 703
rect 1098 698 1099 702
rect 1103 698 1104 702
rect 1098 697 1104 698
rect 1172 664 1174 718
rect 1183 717 1187 718
rect 1184 698 1186 717
rect 1182 697 1188 698
rect 1182 693 1183 697
rect 1187 693 1188 697
rect 1182 692 1188 693
rect 1182 679 1188 680
rect 1182 675 1183 679
rect 1187 675 1188 679
rect 1182 674 1188 675
rect 1170 663 1176 664
rect 1094 661 1100 662
rect 1094 657 1095 661
rect 1099 657 1100 661
rect 1170 659 1171 663
rect 1175 659 1176 663
rect 1170 658 1176 659
rect 1094 656 1100 657
rect 1096 647 1098 656
rect 1184 647 1186 674
rect 1095 646 1099 647
rect 1095 641 1099 642
rect 1183 646 1187 647
rect 1183 641 1187 642
rect 1096 636 1098 641
rect 1094 635 1100 636
rect 1094 631 1095 635
rect 1099 631 1100 635
rect 1094 630 1100 631
rect 1046 627 1052 628
rect 1046 623 1047 627
rect 1051 623 1052 627
rect 1046 622 1052 623
rect 1170 623 1176 624
rect 1170 619 1171 623
rect 1175 619 1176 623
rect 1170 618 1176 619
rect 1184 618 1186 641
rect 1098 594 1104 595
rect 1098 590 1099 594
rect 1103 590 1104 594
rect 1098 589 1104 590
rect 1100 575 1102 589
rect 1099 574 1103 575
rect 1099 569 1103 570
rect 1100 555 1102 569
rect 1098 554 1104 555
rect 1098 550 1099 554
rect 1103 550 1104 554
rect 1098 549 1104 550
rect 1172 516 1174 618
rect 1182 617 1188 618
rect 1182 613 1183 617
rect 1187 613 1188 617
rect 1182 612 1188 613
rect 1182 599 1188 600
rect 1182 595 1183 599
rect 1187 595 1188 599
rect 1182 594 1188 595
rect 1184 575 1186 594
rect 1183 574 1187 575
rect 1183 569 1187 570
rect 1184 550 1186 569
rect 1182 549 1188 550
rect 1182 545 1183 549
rect 1187 545 1188 549
rect 1182 544 1188 545
rect 1182 531 1188 532
rect 1182 527 1183 531
rect 1187 527 1188 531
rect 1182 526 1188 527
rect 1170 515 1176 516
rect 1094 513 1100 514
rect 1094 509 1095 513
rect 1099 509 1100 513
rect 1170 511 1171 515
rect 1175 511 1176 515
rect 1170 510 1176 511
rect 1094 508 1100 509
rect 1096 495 1098 508
rect 1184 495 1186 526
rect 967 494 971 495
rect 967 489 971 490
rect 1095 494 1099 495
rect 1095 489 1099 490
rect 1183 494 1187 495
rect 1183 489 1187 490
rect 968 484 970 489
rect 1096 484 1098 489
rect 966 483 972 484
rect 966 479 967 483
rect 971 479 972 483
rect 1094 483 1100 484
rect 966 478 972 479
rect 1030 479 1036 480
rect 946 475 952 476
rect 486 471 492 472
rect 486 467 487 471
rect 491 467 492 471
rect 486 466 492 467
rect 738 471 744 472
rect 783 471 787 472
rect 946 471 947 475
rect 951 471 952 475
rect 738 467 739 471
rect 743 467 744 471
rect 946 470 952 471
rect 958 475 964 476
rect 958 471 959 475
rect 963 471 964 475
rect 1030 475 1031 479
rect 1035 475 1036 479
rect 1094 479 1095 483
rect 1099 479 1100 483
rect 1094 478 1100 479
rect 1030 474 1036 475
rect 958 470 964 471
rect 738 466 744 467
rect 110 465 116 466
rect 110 461 111 465
rect 115 461 116 465
rect 110 460 116 461
rect 110 447 116 448
rect 110 443 111 447
rect 115 443 116 447
rect 110 442 116 443
rect 410 442 416 443
rect 112 419 114 442
rect 410 438 411 442
rect 415 438 416 442
rect 410 437 416 438
rect 506 442 512 443
rect 506 438 507 442
rect 511 438 512 442
rect 506 437 512 438
rect 610 442 616 443
rect 610 438 611 442
rect 615 438 616 442
rect 610 437 616 438
rect 722 442 728 443
rect 722 438 723 442
rect 727 438 728 442
rect 722 437 728 438
rect 842 442 848 443
rect 842 438 843 442
rect 847 438 848 442
rect 842 437 848 438
rect 412 419 414 437
rect 508 419 510 437
rect 612 419 614 437
rect 724 419 726 437
rect 844 419 846 437
rect 111 418 115 419
rect 111 413 115 414
rect 411 418 415 419
rect 411 413 415 414
rect 507 418 511 419
rect 507 413 511 414
rect 587 418 591 419
rect 587 413 591 414
rect 611 418 615 419
rect 611 413 615 414
rect 675 418 679 419
rect 675 413 679 414
rect 723 418 727 419
rect 723 413 727 414
rect 771 418 775 419
rect 771 413 775 414
rect 843 418 847 419
rect 843 413 847 414
rect 875 418 879 419
rect 875 413 879 414
rect 112 394 114 413
rect 588 399 590 413
rect 676 399 678 413
rect 772 399 774 413
rect 876 399 878 413
rect 586 398 592 399
rect 586 394 587 398
rect 591 394 592 398
rect 110 393 116 394
rect 586 393 592 394
rect 674 398 680 399
rect 674 394 675 398
rect 679 394 680 398
rect 674 393 680 394
rect 770 398 776 399
rect 770 394 771 398
rect 775 394 776 398
rect 770 393 776 394
rect 874 398 880 399
rect 874 394 875 398
rect 879 394 880 398
rect 874 393 880 394
rect 110 389 111 393
rect 115 389 116 393
rect 110 388 116 389
rect 948 388 950 470
rect 970 442 976 443
rect 970 438 971 442
rect 975 438 976 442
rect 970 437 976 438
rect 972 419 974 437
rect 1032 420 1034 474
rect 1184 466 1186 489
rect 1182 465 1188 466
rect 1182 461 1183 465
rect 1187 461 1188 465
rect 1182 460 1188 461
rect 1182 447 1188 448
rect 1182 443 1183 447
rect 1187 443 1188 447
rect 1098 442 1104 443
rect 1182 442 1188 443
rect 1098 438 1099 442
rect 1103 438 1104 442
rect 1098 437 1104 438
rect 978 419 984 420
rect 1030 419 1036 420
rect 1100 419 1102 437
rect 1184 419 1186 442
rect 971 418 975 419
rect 978 415 979 419
rect 983 415 984 419
rect 978 414 984 415
rect 987 418 991 419
rect 1030 415 1031 419
rect 1035 415 1036 419
rect 1030 414 1036 415
rect 1099 418 1103 419
rect 971 413 975 414
rect 980 411 982 414
rect 987 413 991 414
rect 1099 413 1103 414
rect 1183 418 1187 419
rect 1183 413 1187 414
rect 976 409 982 411
rect 946 387 952 388
rect 946 383 947 387
rect 951 383 952 387
rect 946 382 952 383
rect 110 375 116 376
rect 110 371 111 375
rect 115 371 116 375
rect 110 370 116 371
rect 112 347 114 370
rect 654 367 660 368
rect 654 363 655 367
rect 659 363 660 367
rect 654 362 660 363
rect 582 357 588 358
rect 656 357 658 362
rect 670 357 676 358
rect 582 353 583 357
rect 587 353 588 357
rect 582 352 588 353
rect 655 356 659 357
rect 670 353 671 357
rect 675 353 676 357
rect 670 352 676 353
rect 766 357 772 358
rect 766 353 767 357
rect 771 353 772 357
rect 766 352 772 353
rect 870 357 876 358
rect 870 353 871 357
rect 875 353 876 357
rect 870 352 876 353
rect 903 356 907 357
rect 584 347 586 352
rect 655 351 659 352
rect 672 347 674 352
rect 768 347 770 352
rect 872 347 874 352
rect 903 351 907 352
rect 111 346 115 347
rect 111 341 115 342
rect 415 346 419 347
rect 415 341 419 342
rect 511 346 515 347
rect 511 341 515 342
rect 583 346 587 347
rect 583 341 587 342
rect 615 346 619 347
rect 615 341 619 342
rect 671 346 675 347
rect 671 341 675 342
rect 727 346 731 347
rect 727 341 731 342
rect 767 346 771 347
rect 767 341 771 342
rect 839 346 843 347
rect 839 341 843 342
rect 871 346 875 347
rect 871 341 875 342
rect 112 318 114 341
rect 416 336 418 341
rect 512 336 514 341
rect 616 336 618 341
rect 728 336 730 341
rect 840 336 842 341
rect 904 336 906 351
rect 959 346 963 347
rect 959 341 963 342
rect 960 336 962 341
rect 414 335 420 336
rect 414 331 415 335
rect 419 331 420 335
rect 414 330 420 331
rect 510 335 516 336
rect 510 331 511 335
rect 515 331 516 335
rect 510 330 516 331
rect 614 335 620 336
rect 614 331 615 335
rect 619 331 620 335
rect 614 330 620 331
rect 726 335 732 336
rect 726 331 727 335
rect 731 331 732 335
rect 726 330 732 331
rect 838 335 844 336
rect 838 331 839 335
rect 843 331 844 335
rect 838 330 844 331
rect 902 335 908 336
rect 902 331 903 335
rect 907 331 908 335
rect 902 330 908 331
rect 958 335 964 336
rect 958 331 959 335
rect 963 331 964 335
rect 958 330 964 331
rect 976 324 978 409
rect 988 399 990 413
rect 1100 399 1102 413
rect 986 398 992 399
rect 986 394 987 398
rect 991 394 992 398
rect 986 393 992 394
rect 1098 398 1104 399
rect 1098 394 1099 398
rect 1103 394 1104 398
rect 1184 394 1186 413
rect 1098 393 1104 394
rect 1182 393 1188 394
rect 1182 389 1183 393
rect 1187 389 1188 393
rect 1182 388 1188 389
rect 1046 383 1052 384
rect 1046 379 1047 383
rect 1051 379 1052 383
rect 1046 378 1052 379
rect 1048 360 1050 378
rect 1182 375 1188 376
rect 1182 371 1183 375
rect 1187 371 1188 375
rect 1182 370 1188 371
rect 1166 367 1172 368
rect 1166 363 1167 367
rect 1171 363 1172 367
rect 1166 362 1172 363
rect 1046 359 1052 360
rect 982 357 988 358
rect 982 353 983 357
rect 987 353 988 357
rect 1046 355 1047 359
rect 1051 355 1052 359
rect 1046 354 1052 355
rect 1094 357 1100 358
rect 982 352 988 353
rect 1094 353 1095 357
rect 1099 353 1100 357
rect 1094 352 1100 353
rect 984 347 986 352
rect 1096 347 1098 352
rect 983 346 987 347
rect 983 341 987 342
rect 1087 346 1091 347
rect 1087 341 1091 342
rect 1095 346 1099 347
rect 1095 341 1099 342
rect 1088 336 1090 341
rect 1086 335 1092 336
rect 1026 331 1032 332
rect 1026 327 1027 331
rect 1031 327 1032 331
rect 1086 331 1087 335
rect 1091 331 1092 335
rect 1168 332 1170 362
rect 1184 347 1186 370
rect 1183 346 1187 347
rect 1183 341 1187 342
rect 1086 330 1092 331
rect 1166 331 1172 332
rect 1026 326 1032 327
rect 1166 327 1167 331
rect 1171 327 1172 331
rect 1166 326 1172 327
rect 494 323 500 324
rect 494 319 495 323
rect 499 319 500 323
rect 494 318 500 319
rect 974 323 980 324
rect 974 319 975 323
rect 979 319 980 323
rect 974 318 980 319
rect 110 317 116 318
rect 110 313 111 317
rect 115 313 116 317
rect 110 312 116 313
rect 110 299 116 300
rect 110 295 111 299
rect 115 295 116 299
rect 110 294 116 295
rect 418 294 424 295
rect 112 271 114 294
rect 418 290 419 294
rect 423 290 424 294
rect 418 289 424 290
rect 420 271 422 289
rect 496 272 498 318
rect 514 294 520 295
rect 514 290 515 294
rect 519 290 520 294
rect 514 289 520 290
rect 618 294 624 295
rect 618 290 619 294
rect 623 290 624 294
rect 618 289 624 290
rect 730 294 736 295
rect 730 290 731 294
rect 735 290 736 294
rect 730 289 736 290
rect 842 294 848 295
rect 842 290 843 294
rect 847 290 848 294
rect 842 289 848 290
rect 962 294 968 295
rect 962 290 963 294
rect 967 290 968 294
rect 962 289 968 290
rect 494 271 500 272
rect 516 271 518 289
rect 620 271 622 289
rect 702 271 708 272
rect 732 271 734 289
rect 844 271 846 289
rect 964 271 966 289
rect 1028 272 1030 326
rect 1158 323 1164 324
rect 1158 319 1159 323
rect 1163 319 1164 323
rect 1158 318 1164 319
rect 1184 318 1186 341
rect 1090 294 1096 295
rect 1090 290 1091 294
rect 1095 290 1096 294
rect 1090 289 1096 290
rect 1026 271 1032 272
rect 1092 271 1094 289
rect 111 270 115 271
rect 111 265 115 266
rect 203 270 207 271
rect 203 265 207 266
rect 307 270 311 271
rect 307 265 311 266
rect 419 270 423 271
rect 494 267 495 271
rect 499 267 500 271
rect 494 266 500 267
rect 515 270 519 271
rect 419 265 423 266
rect 515 265 519 266
rect 531 270 535 271
rect 531 265 535 266
rect 619 270 623 271
rect 619 265 623 266
rect 643 270 647 271
rect 702 267 703 271
rect 707 267 708 271
rect 702 266 708 267
rect 731 270 735 271
rect 643 265 647 266
rect 112 246 114 265
rect 204 251 206 265
rect 308 251 310 265
rect 420 251 422 265
rect 532 251 534 265
rect 644 251 646 265
rect 202 250 208 251
rect 202 246 203 250
rect 207 246 208 250
rect 110 245 116 246
rect 202 245 208 246
rect 306 250 312 251
rect 306 246 307 250
rect 311 246 312 250
rect 306 245 312 246
rect 418 250 424 251
rect 418 246 419 250
rect 423 246 424 250
rect 418 245 424 246
rect 530 250 536 251
rect 530 246 531 250
rect 535 246 536 250
rect 530 245 536 246
rect 642 250 648 251
rect 642 246 643 250
rect 647 246 648 250
rect 642 245 648 246
rect 110 241 111 245
rect 115 241 116 245
rect 110 240 116 241
rect 110 227 116 228
rect 110 223 111 227
rect 115 223 116 227
rect 110 222 116 223
rect 112 171 114 222
rect 704 212 706 266
rect 731 265 735 266
rect 763 270 767 271
rect 763 265 767 266
rect 843 270 847 271
rect 843 265 847 266
rect 883 270 887 271
rect 883 265 887 266
rect 963 270 967 271
rect 963 265 967 266
rect 1003 270 1007 271
rect 1026 267 1027 271
rect 1031 267 1032 271
rect 1026 266 1032 267
rect 1091 270 1095 271
rect 1003 265 1007 266
rect 1091 265 1095 266
rect 1099 270 1103 271
rect 1099 265 1103 266
rect 764 251 766 265
rect 884 251 886 265
rect 1004 251 1006 265
rect 1100 251 1102 265
rect 762 250 768 251
rect 762 246 763 250
rect 767 246 768 250
rect 762 245 768 246
rect 882 250 888 251
rect 882 246 883 250
rect 887 246 888 250
rect 882 245 888 246
rect 1002 250 1008 251
rect 1002 246 1003 250
rect 1007 246 1008 250
rect 1002 245 1008 246
rect 1098 250 1104 251
rect 1098 246 1099 250
rect 1103 246 1104 250
rect 1098 245 1104 246
rect 1160 212 1162 318
rect 1182 317 1188 318
rect 1182 313 1183 317
rect 1187 313 1188 317
rect 1182 312 1188 313
rect 1182 299 1188 300
rect 1182 295 1183 299
rect 1187 295 1188 299
rect 1182 294 1188 295
rect 1184 271 1186 294
rect 1183 270 1187 271
rect 1183 265 1187 266
rect 1184 246 1186 265
rect 1182 245 1188 246
rect 1182 241 1183 245
rect 1187 241 1188 245
rect 1182 240 1188 241
rect 1182 227 1188 228
rect 1182 223 1183 227
rect 1187 223 1188 227
rect 1182 222 1188 223
rect 702 211 708 212
rect 198 209 204 210
rect 198 205 199 209
rect 203 205 204 209
rect 198 204 204 205
rect 302 209 308 210
rect 302 205 303 209
rect 307 205 308 209
rect 302 204 308 205
rect 414 209 420 210
rect 414 205 415 209
rect 419 205 420 209
rect 414 204 420 205
rect 526 209 532 210
rect 526 205 527 209
rect 531 205 532 209
rect 526 204 532 205
rect 638 209 644 210
rect 638 205 639 209
rect 643 205 644 209
rect 702 207 703 211
rect 707 207 708 211
rect 1158 211 1164 212
rect 702 206 708 207
rect 758 209 764 210
rect 638 204 644 205
rect 758 205 759 209
rect 763 205 764 209
rect 758 204 764 205
rect 878 209 884 210
rect 878 205 879 209
rect 883 205 884 209
rect 878 204 884 205
rect 998 209 1004 210
rect 998 205 999 209
rect 1003 205 1004 209
rect 998 204 1004 205
rect 1094 209 1100 210
rect 1094 205 1095 209
rect 1099 205 1100 209
rect 1158 207 1159 211
rect 1163 207 1164 211
rect 1158 206 1164 207
rect 1094 204 1100 205
rect 200 171 202 204
rect 304 171 306 204
rect 416 171 418 204
rect 528 171 530 204
rect 640 171 642 204
rect 760 171 762 204
rect 880 171 882 204
rect 1000 171 1002 204
rect 1096 171 1098 204
rect 1184 171 1186 222
rect 111 170 115 171
rect 111 165 115 166
rect 143 170 147 171
rect 143 165 147 166
rect 199 170 203 171
rect 199 165 203 166
rect 231 170 235 171
rect 231 165 235 166
rect 303 170 307 171
rect 303 165 307 166
rect 319 170 323 171
rect 319 165 323 166
rect 407 170 411 171
rect 407 165 411 166
rect 415 170 419 171
rect 415 165 419 166
rect 495 170 499 171
rect 495 165 499 166
rect 527 170 531 171
rect 527 165 531 166
rect 583 170 587 171
rect 583 165 587 166
rect 639 170 643 171
rect 639 165 643 166
rect 671 170 675 171
rect 671 165 675 166
rect 759 170 763 171
rect 759 165 763 166
rect 879 170 883 171
rect 879 165 883 166
rect 999 170 1003 171
rect 999 165 1003 166
rect 1095 170 1099 171
rect 1095 165 1099 166
rect 1183 170 1187 171
rect 1183 165 1187 166
rect 112 142 114 165
rect 144 160 146 165
rect 232 160 234 165
rect 320 160 322 165
rect 408 160 410 165
rect 496 160 498 165
rect 584 160 586 165
rect 672 160 674 165
rect 760 160 762 165
rect 142 159 148 160
rect 142 155 143 159
rect 147 155 148 159
rect 142 154 148 155
rect 230 159 236 160
rect 230 155 231 159
rect 235 155 236 159
rect 230 154 236 155
rect 318 159 324 160
rect 318 155 319 159
rect 323 155 324 159
rect 318 154 324 155
rect 406 159 412 160
rect 406 155 407 159
rect 411 155 412 159
rect 406 154 412 155
rect 494 159 500 160
rect 494 155 495 159
rect 499 155 500 159
rect 494 154 500 155
rect 582 159 588 160
rect 582 155 583 159
rect 587 155 588 159
rect 582 154 588 155
rect 670 159 676 160
rect 670 155 671 159
rect 675 155 676 159
rect 670 154 676 155
rect 758 159 764 160
rect 758 155 759 159
rect 763 155 764 159
rect 758 154 764 155
rect 1184 142 1186 165
rect 110 141 116 142
rect 110 137 111 141
rect 115 137 116 141
rect 110 136 116 137
rect 1182 141 1188 142
rect 1182 137 1183 141
rect 1187 137 1188 141
rect 1182 136 1188 137
rect 110 123 116 124
rect 110 119 111 123
rect 115 119 116 123
rect 1182 123 1188 124
rect 1182 119 1183 123
rect 1187 119 1188 123
rect 110 118 116 119
rect 146 118 152 119
rect 112 99 114 118
rect 146 114 147 118
rect 151 114 152 118
rect 146 113 152 114
rect 234 118 240 119
rect 234 114 235 118
rect 239 114 240 118
rect 234 113 240 114
rect 322 118 328 119
rect 322 114 323 118
rect 327 114 328 118
rect 322 113 328 114
rect 410 118 416 119
rect 410 114 411 118
rect 415 114 416 118
rect 410 113 416 114
rect 498 118 504 119
rect 498 114 499 118
rect 503 114 504 118
rect 498 113 504 114
rect 586 118 592 119
rect 586 114 587 118
rect 591 114 592 118
rect 586 113 592 114
rect 674 118 680 119
rect 674 114 675 118
rect 679 114 680 118
rect 674 113 680 114
rect 762 118 768 119
rect 1182 118 1188 119
rect 762 114 763 118
rect 767 114 768 118
rect 762 113 768 114
rect 148 99 150 113
rect 236 99 238 113
rect 324 99 326 113
rect 412 99 414 113
rect 500 99 502 113
rect 588 99 590 113
rect 676 99 678 113
rect 764 99 766 113
rect 1184 99 1186 118
rect 111 98 115 99
rect 111 93 115 94
rect 147 98 151 99
rect 147 93 151 94
rect 235 98 239 99
rect 235 93 239 94
rect 323 98 327 99
rect 323 93 327 94
rect 411 98 415 99
rect 411 93 415 94
rect 499 98 503 99
rect 499 93 503 94
rect 587 98 591 99
rect 587 93 591 94
rect 675 98 679 99
rect 675 93 679 94
rect 763 98 767 99
rect 763 93 767 94
rect 1183 98 1187 99
rect 1183 93 1187 94
<< m4c >>
rect 111 1282 115 1286
rect 663 1282 667 1286
rect 751 1282 755 1286
rect 839 1282 843 1286
rect 927 1282 931 1286
rect 1183 1282 1187 1286
rect 111 1210 115 1214
rect 371 1210 375 1214
rect 459 1210 463 1214
rect 555 1210 559 1214
rect 651 1210 655 1214
rect 667 1210 671 1214
rect 755 1210 759 1214
rect 843 1210 847 1214
rect 859 1210 863 1214
rect 931 1210 935 1214
rect 963 1210 967 1214
rect 111 1130 115 1134
rect 143 1130 147 1134
rect 255 1130 259 1134
rect 367 1130 371 1134
rect 415 1130 419 1134
rect 1183 1210 1187 1214
rect 455 1130 459 1134
rect 551 1130 555 1134
rect 583 1130 587 1134
rect 647 1130 651 1134
rect 751 1130 755 1134
rect 767 1130 771 1134
rect 855 1130 859 1134
rect 439 1120 443 1124
rect 831 1123 835 1124
rect 831 1120 835 1123
rect 951 1130 955 1134
rect 959 1130 963 1134
rect 1183 1130 1187 1134
rect 111 1042 115 1046
rect 147 1042 151 1046
rect 155 1042 159 1046
rect 259 1042 263 1046
rect 283 1042 287 1046
rect 419 1042 423 1046
rect 427 1042 431 1046
rect 587 1042 591 1046
rect 755 1042 759 1046
rect 771 1042 775 1046
rect 939 1042 943 1046
rect 955 1042 959 1046
rect 1099 1042 1103 1046
rect 1183 1042 1187 1046
rect 111 962 115 966
rect 151 962 155 966
rect 279 962 283 966
rect 423 962 427 966
rect 503 962 507 966
rect 583 962 587 966
rect 591 962 595 966
rect 687 962 691 966
rect 751 962 755 966
rect 791 962 795 966
rect 895 962 899 966
rect 935 962 939 966
rect 575 944 579 948
rect 855 947 859 948
rect 855 944 859 947
rect 111 882 115 886
rect 507 882 511 886
rect 563 882 567 886
rect 595 882 599 886
rect 651 882 655 886
rect 691 882 695 886
rect 739 882 743 886
rect 795 882 799 886
rect 827 882 831 886
rect 899 882 903 886
rect 923 882 927 886
rect 111 794 115 798
rect 391 794 395 798
rect 495 794 499 798
rect 559 794 563 798
rect 607 794 611 798
rect 1007 962 1011 966
rect 1095 962 1099 966
rect 1183 962 1187 966
rect 1011 882 1015 886
rect 1099 882 1103 886
rect 1183 882 1187 886
rect 647 794 651 798
rect 727 794 731 798
rect 735 794 739 798
rect 823 794 827 798
rect 855 794 859 798
rect 919 794 923 798
rect 983 794 987 798
rect 1007 794 1011 798
rect 1095 794 1099 798
rect 1183 794 1187 798
rect 111 718 115 722
rect 211 718 215 722
rect 355 718 359 722
rect 395 718 399 722
rect 111 642 115 646
rect 143 642 147 646
rect 207 642 211 646
rect 295 642 299 646
rect 631 768 635 772
rect 919 768 923 772
rect 499 718 503 722
rect 523 718 527 722
rect 611 718 615 722
rect 715 718 719 722
rect 731 718 735 722
rect 859 718 863 722
rect 915 718 919 722
rect 987 718 991 722
rect 351 642 355 646
rect 487 642 491 646
rect 519 642 523 646
rect 687 642 691 646
rect 711 642 715 646
rect 895 642 899 646
rect 911 642 915 646
rect 335 632 339 636
rect 751 635 755 636
rect 751 632 755 635
rect 111 570 115 574
rect 147 570 151 574
rect 283 570 287 574
rect 299 570 303 574
rect 467 570 471 574
rect 491 570 495 574
rect 667 570 671 574
rect 691 570 695 574
rect 883 570 887 574
rect 899 570 903 574
rect 111 490 115 494
rect 143 490 147 494
rect 279 490 283 494
rect 407 490 411 494
rect 463 490 467 494
rect 503 490 507 494
rect 607 490 611 494
rect 663 490 667 494
rect 719 490 723 494
rect 839 490 843 494
rect 879 490 883 494
rect 487 472 491 476
rect 783 475 787 476
rect 783 472 787 475
rect 1099 718 1103 722
rect 1183 718 1187 722
rect 1095 642 1099 646
rect 1183 642 1187 646
rect 1099 570 1103 574
rect 1183 570 1187 574
rect 967 490 971 494
rect 1095 490 1099 494
rect 1183 490 1187 494
rect 111 414 115 418
rect 411 414 415 418
rect 507 414 511 418
rect 587 414 591 418
rect 611 414 615 418
rect 675 414 679 418
rect 723 414 727 418
rect 771 414 775 418
rect 843 414 847 418
rect 875 414 879 418
rect 971 414 975 418
rect 987 414 991 418
rect 1099 414 1103 418
rect 1183 414 1187 418
rect 655 352 659 356
rect 903 352 907 356
rect 111 342 115 346
rect 415 342 419 346
rect 511 342 515 346
rect 583 342 587 346
rect 615 342 619 346
rect 671 342 675 346
rect 727 342 731 346
rect 767 342 771 346
rect 839 342 843 346
rect 871 342 875 346
rect 959 342 963 346
rect 983 342 987 346
rect 1087 342 1091 346
rect 1095 342 1099 346
rect 1183 342 1187 346
rect 111 266 115 270
rect 203 266 207 270
rect 307 266 311 270
rect 419 266 423 270
rect 515 266 519 270
rect 531 266 535 270
rect 619 266 623 270
rect 643 266 647 270
rect 731 266 735 270
rect 763 266 767 270
rect 843 266 847 270
rect 883 266 887 270
rect 963 266 967 270
rect 1003 266 1007 270
rect 1091 266 1095 270
rect 1099 266 1103 270
rect 1183 266 1187 270
rect 111 166 115 170
rect 143 166 147 170
rect 199 166 203 170
rect 231 166 235 170
rect 303 166 307 170
rect 319 166 323 170
rect 407 166 411 170
rect 415 166 419 170
rect 495 166 499 170
rect 527 166 531 170
rect 583 166 587 170
rect 639 166 643 170
rect 671 166 675 170
rect 759 166 763 170
rect 879 166 883 170
rect 999 166 1003 170
rect 1095 166 1099 170
rect 1183 166 1187 170
rect 111 94 115 98
rect 147 94 151 98
rect 235 94 239 98
rect 323 94 327 98
rect 411 94 415 98
rect 499 94 503 98
rect 587 94 591 98
rect 675 94 679 98
rect 763 94 767 98
rect 1183 94 1187 98
<< m4 >>
rect 96 1281 97 1287
rect 103 1286 1219 1287
rect 103 1282 111 1286
rect 115 1282 663 1286
rect 667 1282 751 1286
rect 755 1282 839 1286
rect 843 1282 927 1286
rect 931 1282 1183 1286
rect 1187 1282 1219 1286
rect 103 1281 1219 1282
rect 1225 1281 1226 1287
rect 84 1209 85 1215
rect 91 1214 1207 1215
rect 91 1210 111 1214
rect 115 1210 371 1214
rect 375 1210 459 1214
rect 463 1210 555 1214
rect 559 1210 651 1214
rect 655 1210 667 1214
rect 671 1210 755 1214
rect 759 1210 843 1214
rect 847 1210 859 1214
rect 863 1210 931 1214
rect 935 1210 963 1214
rect 967 1210 1183 1214
rect 1187 1210 1207 1214
rect 91 1209 1207 1210
rect 1213 1209 1214 1215
rect 96 1129 97 1135
rect 103 1134 1219 1135
rect 103 1130 111 1134
rect 115 1130 143 1134
rect 147 1130 255 1134
rect 259 1130 367 1134
rect 371 1130 415 1134
rect 419 1130 455 1134
rect 459 1130 551 1134
rect 555 1130 583 1134
rect 587 1130 647 1134
rect 651 1130 751 1134
rect 755 1130 767 1134
rect 771 1130 855 1134
rect 859 1130 951 1134
rect 955 1130 959 1134
rect 963 1130 1183 1134
rect 1187 1130 1219 1134
rect 103 1129 1219 1130
rect 1225 1129 1226 1135
rect 438 1124 444 1125
rect 830 1124 836 1125
rect 438 1120 439 1124
rect 443 1120 831 1124
rect 835 1120 836 1124
rect 438 1119 444 1120
rect 830 1119 836 1120
rect 84 1041 85 1047
rect 91 1046 1207 1047
rect 91 1042 111 1046
rect 115 1042 147 1046
rect 151 1042 155 1046
rect 159 1042 259 1046
rect 263 1042 283 1046
rect 287 1042 419 1046
rect 423 1042 427 1046
rect 431 1042 587 1046
rect 591 1042 755 1046
rect 759 1042 771 1046
rect 775 1042 939 1046
rect 943 1042 955 1046
rect 959 1042 1099 1046
rect 1103 1042 1183 1046
rect 1187 1042 1207 1046
rect 91 1041 1207 1042
rect 1213 1041 1214 1047
rect 96 961 97 967
rect 103 966 1219 967
rect 103 962 111 966
rect 115 962 151 966
rect 155 962 279 966
rect 283 962 423 966
rect 427 962 503 966
rect 507 962 583 966
rect 587 962 591 966
rect 595 962 687 966
rect 691 962 751 966
rect 755 962 791 966
rect 795 962 895 966
rect 899 962 935 966
rect 939 962 1007 966
rect 1011 962 1095 966
rect 1099 962 1183 966
rect 1187 962 1219 966
rect 103 961 1219 962
rect 1225 961 1226 967
rect 574 948 580 949
rect 854 948 860 949
rect 574 944 575 948
rect 579 944 855 948
rect 859 944 860 948
rect 574 943 580 944
rect 854 943 860 944
rect 84 881 85 887
rect 91 886 1207 887
rect 91 882 111 886
rect 115 882 507 886
rect 511 882 563 886
rect 567 882 595 886
rect 599 882 651 886
rect 655 882 691 886
rect 695 882 739 886
rect 743 882 795 886
rect 799 882 827 886
rect 831 882 899 886
rect 903 882 923 886
rect 927 882 1011 886
rect 1015 882 1099 886
rect 1103 882 1183 886
rect 1187 882 1207 886
rect 91 881 1207 882
rect 1213 881 1214 887
rect 96 793 97 799
rect 103 798 1219 799
rect 103 794 111 798
rect 115 794 391 798
rect 395 794 495 798
rect 499 794 559 798
rect 563 794 607 798
rect 611 794 647 798
rect 651 794 727 798
rect 731 794 735 798
rect 739 794 823 798
rect 827 794 855 798
rect 859 794 919 798
rect 923 794 983 798
rect 987 794 1007 798
rect 1011 794 1095 798
rect 1099 794 1183 798
rect 1187 794 1219 798
rect 103 793 1219 794
rect 1225 793 1226 799
rect 630 772 636 773
rect 918 772 924 773
rect 630 768 631 772
rect 635 768 919 772
rect 923 768 924 772
rect 630 767 636 768
rect 918 767 924 768
rect 84 717 85 723
rect 91 722 1207 723
rect 91 718 111 722
rect 115 718 211 722
rect 215 718 355 722
rect 359 718 395 722
rect 399 718 499 722
rect 503 718 523 722
rect 527 718 611 722
rect 615 718 715 722
rect 719 718 731 722
rect 735 718 859 722
rect 863 718 915 722
rect 919 718 987 722
rect 991 718 1099 722
rect 1103 718 1183 722
rect 1187 718 1207 722
rect 91 717 1207 718
rect 1213 717 1214 723
rect 96 641 97 647
rect 103 646 1219 647
rect 103 642 111 646
rect 115 642 143 646
rect 147 642 207 646
rect 211 642 295 646
rect 299 642 351 646
rect 355 642 487 646
rect 491 642 519 646
rect 523 642 687 646
rect 691 642 711 646
rect 715 642 895 646
rect 899 642 911 646
rect 915 642 1095 646
rect 1099 642 1183 646
rect 1187 642 1219 646
rect 103 641 1219 642
rect 1225 641 1226 647
rect 334 636 340 637
rect 750 636 756 637
rect 334 632 335 636
rect 339 632 751 636
rect 755 632 756 636
rect 334 631 340 632
rect 750 631 756 632
rect 84 569 85 575
rect 91 574 1207 575
rect 91 570 111 574
rect 115 570 147 574
rect 151 570 283 574
rect 287 570 299 574
rect 303 570 467 574
rect 471 570 491 574
rect 495 570 667 574
rect 671 570 691 574
rect 695 570 883 574
rect 887 570 899 574
rect 903 570 1099 574
rect 1103 570 1183 574
rect 1187 570 1207 574
rect 91 569 1207 570
rect 1213 569 1214 575
rect 96 489 97 495
rect 103 494 1219 495
rect 103 490 111 494
rect 115 490 143 494
rect 147 490 279 494
rect 283 490 407 494
rect 411 490 463 494
rect 467 490 503 494
rect 507 490 607 494
rect 611 490 663 494
rect 667 490 719 494
rect 723 490 839 494
rect 843 490 879 494
rect 883 490 967 494
rect 971 490 1095 494
rect 1099 490 1183 494
rect 1187 490 1219 494
rect 103 489 1219 490
rect 1225 489 1226 495
rect 486 476 492 477
rect 782 476 788 477
rect 486 472 487 476
rect 491 472 783 476
rect 787 472 788 476
rect 486 471 492 472
rect 782 471 788 472
rect 84 413 85 419
rect 91 418 1207 419
rect 91 414 111 418
rect 115 414 411 418
rect 415 414 507 418
rect 511 414 587 418
rect 591 414 611 418
rect 615 414 675 418
rect 679 414 723 418
rect 727 414 771 418
rect 775 414 843 418
rect 847 414 875 418
rect 879 414 971 418
rect 975 414 987 418
rect 991 414 1099 418
rect 1103 414 1183 418
rect 1187 414 1207 418
rect 91 413 1207 414
rect 1213 413 1214 419
rect 654 356 660 357
rect 902 356 908 357
rect 654 352 655 356
rect 659 352 903 356
rect 907 352 908 356
rect 654 351 660 352
rect 902 351 908 352
rect 96 341 97 347
rect 103 346 1219 347
rect 103 342 111 346
rect 115 342 415 346
rect 419 342 511 346
rect 515 342 583 346
rect 587 342 615 346
rect 619 342 671 346
rect 675 342 727 346
rect 731 342 767 346
rect 771 342 839 346
rect 843 342 871 346
rect 875 342 959 346
rect 963 342 983 346
rect 987 342 1087 346
rect 1091 342 1095 346
rect 1099 342 1183 346
rect 1187 342 1219 346
rect 103 341 1219 342
rect 1225 341 1226 347
rect 84 265 85 271
rect 91 270 1207 271
rect 91 266 111 270
rect 115 266 203 270
rect 207 266 307 270
rect 311 266 419 270
rect 423 266 515 270
rect 519 266 531 270
rect 535 266 619 270
rect 623 266 643 270
rect 647 266 731 270
rect 735 266 763 270
rect 767 266 843 270
rect 847 266 883 270
rect 887 266 963 270
rect 967 266 1003 270
rect 1007 266 1091 270
rect 1095 266 1099 270
rect 1103 266 1183 270
rect 1187 266 1207 270
rect 91 265 1207 266
rect 1213 265 1214 271
rect 96 165 97 171
rect 103 170 1219 171
rect 103 166 111 170
rect 115 166 143 170
rect 147 166 199 170
rect 203 166 231 170
rect 235 166 303 170
rect 307 166 319 170
rect 323 166 407 170
rect 411 166 415 170
rect 419 166 495 170
rect 499 166 527 170
rect 531 166 583 170
rect 587 166 639 170
rect 643 166 671 170
rect 675 166 759 170
rect 763 166 879 170
rect 883 166 999 170
rect 1003 166 1095 170
rect 1099 166 1183 170
rect 1187 166 1219 170
rect 103 165 1219 166
rect 1225 165 1226 171
rect 84 93 85 99
rect 91 98 1207 99
rect 91 94 111 98
rect 115 94 147 98
rect 151 94 235 98
rect 239 94 323 98
rect 327 94 411 98
rect 415 94 499 98
rect 503 94 587 98
rect 591 94 675 98
rect 679 94 763 98
rect 767 94 1183 98
rect 1187 94 1207 98
rect 91 93 1207 94
rect 1213 93 1214 99
<< m5c >>
rect 97 1281 103 1287
rect 1219 1281 1225 1287
rect 85 1209 91 1215
rect 1207 1209 1213 1215
rect 97 1129 103 1135
rect 1219 1129 1225 1135
rect 85 1041 91 1047
rect 1207 1041 1213 1047
rect 97 961 103 967
rect 1219 961 1225 967
rect 85 881 91 887
rect 1207 881 1213 887
rect 97 793 103 799
rect 1219 793 1225 799
rect 85 717 91 723
rect 1207 717 1213 723
rect 97 641 103 647
rect 1219 641 1225 647
rect 85 569 91 575
rect 1207 569 1213 575
rect 97 489 103 495
rect 1219 489 1225 495
rect 85 413 91 419
rect 1207 413 1213 419
rect 97 341 103 347
rect 1219 341 1225 347
rect 85 265 91 271
rect 1207 265 1213 271
rect 97 165 103 171
rect 1219 165 1225 171
rect 85 93 91 99
rect 1207 93 1213 99
<< m5 >>
rect 84 1215 92 1296
rect 84 1209 85 1215
rect 91 1209 92 1215
rect 84 1047 92 1209
rect 84 1041 85 1047
rect 91 1041 92 1047
rect 84 887 92 1041
rect 84 881 85 887
rect 91 881 92 887
rect 84 723 92 881
rect 84 717 85 723
rect 91 717 92 723
rect 84 575 92 717
rect 84 569 85 575
rect 91 569 92 575
rect 84 419 92 569
rect 84 413 85 419
rect 91 413 92 419
rect 84 271 92 413
rect 84 265 85 271
rect 91 265 92 271
rect 84 99 92 265
rect 84 93 85 99
rect 91 93 92 99
rect 84 72 92 93
rect 96 1287 104 1296
rect 96 1281 97 1287
rect 103 1281 104 1287
rect 96 1135 104 1281
rect 96 1129 97 1135
rect 103 1129 104 1135
rect 96 967 104 1129
rect 96 961 97 967
rect 103 961 104 967
rect 96 799 104 961
rect 96 793 97 799
rect 103 793 104 799
rect 96 647 104 793
rect 96 641 97 647
rect 103 641 104 647
rect 96 495 104 641
rect 96 489 97 495
rect 103 489 104 495
rect 96 347 104 489
rect 96 341 97 347
rect 103 341 104 347
rect 96 171 104 341
rect 96 165 97 171
rect 103 165 104 171
rect 96 72 104 165
rect 1206 1215 1214 1296
rect 1206 1209 1207 1215
rect 1213 1209 1214 1215
rect 1206 1047 1214 1209
rect 1206 1041 1207 1047
rect 1213 1041 1214 1047
rect 1206 887 1214 1041
rect 1206 881 1207 887
rect 1213 881 1214 887
rect 1206 723 1214 881
rect 1206 717 1207 723
rect 1213 717 1214 723
rect 1206 575 1214 717
rect 1206 569 1207 575
rect 1213 569 1214 575
rect 1206 419 1214 569
rect 1206 413 1207 419
rect 1213 413 1214 419
rect 1206 271 1214 413
rect 1206 265 1207 271
rect 1213 265 1214 271
rect 1206 99 1214 265
rect 1206 93 1207 99
rect 1213 93 1214 99
rect 1206 72 1214 93
rect 1218 1287 1226 1296
rect 1218 1281 1219 1287
rect 1225 1281 1226 1287
rect 1218 1135 1226 1281
rect 1218 1129 1219 1135
rect 1225 1129 1226 1135
rect 1218 967 1226 1129
rect 1218 961 1219 967
rect 1225 961 1226 967
rect 1218 799 1226 961
rect 1218 793 1219 799
rect 1225 793 1226 799
rect 1218 647 1226 793
rect 1218 641 1219 647
rect 1225 641 1226 647
rect 1218 495 1226 641
rect 1218 489 1219 495
rect 1225 489 1226 495
rect 1218 347 1226 489
rect 1218 341 1219 347
rect 1225 341 1226 347
rect 1218 171 1226 341
rect 1218 165 1219 171
rect 1225 165 1226 171
rect 1218 72 1226 165
use _0_0std_0_0cells_0_0LATCH  latch_599_6
timestamp 1730954142
transform 1 0 128 0 1 96
box 7 3 85 69
use welltap_svt  __well_tap__0
timestamp 1730954142
transform 1 0 104 0 1 116
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0LATCH  latch_599_6
timestamp 1730954142
transform 1 0 128 0 1 96
box 7 3 85 69
use welltap_svt  __well_tap__0
timestamp 1730954142
transform 1 0 104 0 1 116
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0LATCH  latch_598_6
timestamp 1730954142
transform 1 0 216 0 1 96
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_598_6
timestamp 1730954142
transform 1 0 216 0 1 96
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_597_6
timestamp 1730954142
transform 1 0 304 0 1 96
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_597_6
timestamp 1730954142
transform 1 0 304 0 1 96
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_596_6
timestamp 1730954142
transform 1 0 392 0 1 96
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_596_6
timestamp 1730954142
transform 1 0 392 0 1 96
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_595_6
timestamp 1730954142
transform 1 0 480 0 1 96
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_595_6
timestamp 1730954142
transform 1 0 480 0 1 96
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_594_6
timestamp 1730954142
transform 1 0 568 0 1 96
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_594_6
timestamp 1730954142
transform 1 0 568 0 1 96
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_593_6
timestamp 1730954142
transform 1 0 656 0 1 96
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_593_6
timestamp 1730954142
transform 1 0 656 0 1 96
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_592_6
timestamp 1730954142
transform 1 0 744 0 1 96
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_592_6
timestamp 1730954142
transform 1 0 744 0 1 96
box 7 3 85 69
use welltap_svt  __well_tap__1
timestamp 1730954142
transform 1 0 1176 0 1 116
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1730954142
transform 1 0 1176 0 1 116
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_591_6
timestamp 1730954142
transform 1 0 184 0 -1 268
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_591_6
timestamp 1730954142
transform 1 0 184 0 -1 268
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_590_6
timestamp 1730954142
transform 1 0 288 0 -1 268
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_590_6
timestamp 1730954142
transform 1 0 288 0 -1 268
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_589_6
timestamp 1730954142
transform 1 0 400 0 -1 268
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_589_6
timestamp 1730954142
transform 1 0 400 0 -1 268
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_588_6
timestamp 1730954142
transform 1 0 512 0 -1 268
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_588_6
timestamp 1730954142
transform 1 0 512 0 -1 268
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_587_6
timestamp 1730954142
transform 1 0 624 0 -1 268
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_587_6
timestamp 1730954142
transform 1 0 624 0 -1 268
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_514_6
timestamp 1730954142
transform 1 0 744 0 -1 268
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_514_6
timestamp 1730954142
transform 1 0 744 0 -1 268
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_513_6
timestamp 1730954142
transform 1 0 864 0 -1 268
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_513_6
timestamp 1730954142
transform 1 0 864 0 -1 268
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_512_6
timestamp 1730954142
transform 1 0 984 0 -1 268
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_512_6
timestamp 1730954142
transform 1 0 984 0 -1 268
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_511_6
timestamp 1730954142
transform 1 0 1080 0 -1 268
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_511_6
timestamp 1730954142
transform 1 0 1080 0 -1 268
box 7 3 85 69
use welltap_svt  __well_tap__2
timestamp 1730954142
transform 1 0 104 0 -1 248
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730954142
transform 1 0 104 0 -1 248
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_586_6
timestamp 1730954142
transform 1 0 400 0 1 272
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_586_6
timestamp 1730954142
transform 1 0 400 0 1 272
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_585_6
timestamp 1730954142
transform 1 0 496 0 1 272
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_585_6
timestamp 1730954142
transform 1 0 496 0 1 272
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_584_6
timestamp 1730954142
transform 1 0 600 0 1 272
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_584_6
timestamp 1730954142
transform 1 0 600 0 1 272
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_583_6
timestamp 1730954142
transform 1 0 712 0 1 272
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_583_6
timestamp 1730954142
transform 1 0 712 0 1 272
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_582_6
timestamp 1730954142
transform 1 0 824 0 1 272
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_582_6
timestamp 1730954142
transform 1 0 824 0 1 272
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_515_6
timestamp 1730954142
transform 1 0 944 0 1 272
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_515_6
timestamp 1730954142
transform 1 0 944 0 1 272
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_510_6
timestamp 1730954142
transform 1 0 1072 0 1 272
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_510_6
timestamp 1730954142
transform 1 0 1072 0 1 272
box 7 3 85 69
use welltap_svt  __well_tap__3
timestamp 1730954142
transform 1 0 1176 0 -1 248
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730954142
transform 1 0 1176 0 -1 248
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730954142
transform 1 0 104 0 1 292
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730954142
transform 1 0 104 0 1 292
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_581_6
timestamp 1730954142
transform 1 0 568 0 -1 416
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_581_6
timestamp 1730954142
transform 1 0 568 0 -1 416
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_580_6
timestamp 1730954142
transform 1 0 656 0 -1 416
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_580_6
timestamp 1730954142
transform 1 0 656 0 -1 416
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_579_6
timestamp 1730954142
transform 1 0 752 0 -1 416
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_579_6
timestamp 1730954142
transform 1 0 752 0 -1 416
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_578_6
timestamp 1730954142
transform 1 0 856 0 -1 416
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_578_6
timestamp 1730954142
transform 1 0 856 0 -1 416
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_577_6
timestamp 1730954142
transform 1 0 968 0 -1 416
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_577_6
timestamp 1730954142
transform 1 0 968 0 -1 416
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_59_6
timestamp 1730954142
transform 1 0 1080 0 -1 416
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_59_6
timestamp 1730954142
transform 1 0 1080 0 -1 416
box 7 3 85 69
use welltap_svt  __well_tap__5
timestamp 1730954142
transform 1 0 1176 0 1 292
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730954142
transform 1 0 1176 0 1 292
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730954142
transform 1 0 104 0 -1 396
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730954142
transform 1 0 104 0 -1 396
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_574_6
timestamp 1730954142
transform 1 0 392 0 1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_574_6
timestamp 1730954142
transform 1 0 392 0 1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_573_6
timestamp 1730954142
transform 1 0 488 0 1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_573_6
timestamp 1730954142
transform 1 0 488 0 1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_572_6
timestamp 1730954142
transform 1 0 592 0 1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_572_6
timestamp 1730954142
transform 1 0 592 0 1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_575_6
timestamp 1730954142
transform 1 0 704 0 1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_575_6
timestamp 1730954142
transform 1 0 704 0 1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_576_6
timestamp 1730954142
transform 1 0 824 0 1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_576_6
timestamp 1730954142
transform 1 0 824 0 1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_516_6
timestamp 1730954142
transform 1 0 952 0 1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_516_6
timestamp 1730954142
transform 1 0 952 0 1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_58_6
timestamp 1730954142
transform 1 0 1080 0 1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_58_6
timestamp 1730954142
transform 1 0 1080 0 1 420
box 7 3 85 69
use welltap_svt  __well_tap__7
timestamp 1730954142
transform 1 0 1176 0 -1 396
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1730954142
transform 1 0 1176 0 -1 396
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730954142
transform 1 0 104 0 1 440
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730954142
transform 1 0 104 0 1 440
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730954142
transform 1 0 1176 0 1 440
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730954142
transform 1 0 1176 0 1 440
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_567_6
timestamp 1730954142
transform 1 0 128 0 -1 572
box 7 3 85 69
use welltap_svt  __well_tap__10
timestamp 1730954142
transform 1 0 104 0 -1 552
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_567_6
timestamp 1730954142
transform 1 0 128 0 -1 572
box 7 3 85 69
use welltap_svt  __well_tap__10
timestamp 1730954142
transform 1 0 104 0 -1 552
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_568_6
timestamp 1730954142
transform 1 0 264 0 -1 572
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_568_6
timestamp 1730954142
transform 1 0 264 0 -1 572
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_569_6
timestamp 1730954142
transform 1 0 448 0 -1 572
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_569_6
timestamp 1730954142
transform 1 0 448 0 -1 572
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_571_6
timestamp 1730954142
transform 1 0 648 0 -1 572
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_571_6
timestamp 1730954142
transform 1 0 648 0 -1 572
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_570_6
timestamp 1730954142
transform 1 0 864 0 -1 572
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_570_6
timestamp 1730954142
transform 1 0 864 0 -1 572
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_57_6
timestamp 1730954142
transform 1 0 1080 0 -1 572
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_57_6
timestamp 1730954142
transform 1 0 1080 0 -1 572
box 7 3 85 69
use welltap_svt  __well_tap__11
timestamp 1730954142
transform 1 0 1176 0 -1 552
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730954142
transform 1 0 1176 0 -1 552
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_566_6
timestamp 1730954142
transform 1 0 128 0 1 572
box 7 3 85 69
use welltap_svt  __well_tap__12
timestamp 1730954142
transform 1 0 104 0 1 592
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_566_6
timestamp 1730954142
transform 1 0 128 0 1 572
box 7 3 85 69
use welltap_svt  __well_tap__12
timestamp 1730954142
transform 1 0 104 0 1 592
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_565_6
timestamp 1730954142
transform 1 0 280 0 1 572
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_565_6
timestamp 1730954142
transform 1 0 280 0 1 572
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_564_6
timestamp 1730954142
transform 1 0 472 0 1 572
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_564_6
timestamp 1730954142
transform 1 0 472 0 1 572
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_563_6
timestamp 1730954142
transform 1 0 672 0 1 572
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_563_6
timestamp 1730954142
transform 1 0 672 0 1 572
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_517_6
timestamp 1730954142
transform 1 0 880 0 1 572
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_517_6
timestamp 1730954142
transform 1 0 880 0 1 572
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_56_6
timestamp 1730954142
transform 1 0 1080 0 1 572
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_56_6
timestamp 1730954142
transform 1 0 1080 0 1 572
box 7 3 85 69
use welltap_svt  __well_tap__13
timestamp 1730954142
transform 1 0 1176 0 1 592
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730954142
transform 1 0 1176 0 1 592
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730954142
transform 1 0 104 0 -1 700
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730954142
transform 1 0 104 0 -1 700
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_562_6
timestamp 1730954142
transform 1 0 192 0 -1 720
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_562_6
timestamp 1730954142
transform 1 0 192 0 -1 720
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_561_6
timestamp 1730954142
transform 1 0 336 0 -1 720
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_561_6
timestamp 1730954142
transform 1 0 336 0 -1 720
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_560_6
timestamp 1730954142
transform 1 0 504 0 -1 720
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_560_6
timestamp 1730954142
transform 1 0 504 0 -1 720
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_559_6
timestamp 1730954142
transform 1 0 696 0 -1 720
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_559_6
timestamp 1730954142
transform 1 0 696 0 -1 720
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_558_6
timestamp 1730954142
transform 1 0 896 0 -1 720
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_558_6
timestamp 1730954142
transform 1 0 896 0 -1 720
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_55_6
timestamp 1730954142
transform 1 0 1080 0 -1 720
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_55_6
timestamp 1730954142
transform 1 0 1080 0 -1 720
box 7 3 85 69
use welltap_svt  __well_tap__15
timestamp 1730954142
transform 1 0 1176 0 -1 700
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1730954142
transform 1 0 1176 0 -1 700
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730954142
transform 1 0 104 0 1 744
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730954142
transform 1 0 104 0 1 744
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_557_6
timestamp 1730954142
transform 1 0 376 0 1 724
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_557_6
timestamp 1730954142
transform 1 0 376 0 1 724
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_556_6
timestamp 1730954142
transform 1 0 480 0 1 724
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_556_6
timestamp 1730954142
transform 1 0 480 0 1 724
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_555_6
timestamp 1730954142
transform 1 0 592 0 1 724
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_555_6
timestamp 1730954142
transform 1 0 592 0 1 724
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_554_6
timestamp 1730954142
transform 1 0 712 0 1 724
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_554_6
timestamp 1730954142
transform 1 0 712 0 1 724
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_553_6
timestamp 1730954142
transform 1 0 840 0 1 724
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_553_6
timestamp 1730954142
transform 1 0 840 0 1 724
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_518_6
timestamp 1730954142
transform 1 0 968 0 1 724
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_518_6
timestamp 1730954142
transform 1 0 968 0 1 724
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_54_6
timestamp 1730954142
transform 1 0 1080 0 1 724
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_54_6
timestamp 1730954142
transform 1 0 1080 0 1 724
box 7 3 85 69
use welltap_svt  __well_tap__17
timestamp 1730954142
transform 1 0 1176 0 1 744
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730954142
transform 1 0 1176 0 1 744
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730954142
transform 1 0 104 0 -1 864
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730954142
transform 1 0 104 0 -1 864
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_552_6
timestamp 1730954142
transform 1 0 544 0 -1 884
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_552_6
timestamp 1730954142
transform 1 0 544 0 -1 884
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_551_6
timestamp 1730954142
transform 1 0 632 0 -1 884
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_551_6
timestamp 1730954142
transform 1 0 632 0 -1 884
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_550_6
timestamp 1730954142
transform 1 0 720 0 -1 884
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_550_6
timestamp 1730954142
transform 1 0 720 0 -1 884
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_549_6
timestamp 1730954142
transform 1 0 808 0 -1 884
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_549_6
timestamp 1730954142
transform 1 0 808 0 -1 884
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_548_6
timestamp 1730954142
transform 1 0 904 0 -1 884
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_548_6
timestamp 1730954142
transform 1 0 904 0 -1 884
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_519_6
timestamp 1730954142
transform 1 0 992 0 -1 884
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_519_6
timestamp 1730954142
transform 1 0 992 0 -1 884
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_53_6
timestamp 1730954142
transform 1 0 1080 0 -1 884
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_53_6
timestamp 1730954142
transform 1 0 1080 0 -1 884
box 7 3 85 69
use welltap_svt  __well_tap__19
timestamp 1730954142
transform 1 0 1176 0 -1 864
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730954142
transform 1 0 1176 0 -1 864
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730954142
transform 1 0 104 0 1 912
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730954142
transform 1 0 104 0 1 912
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_545_6
timestamp 1730954142
transform 1 0 488 0 1 892
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_545_6
timestamp 1730954142
transform 1 0 488 0 1 892
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_544_6
timestamp 1730954142
transform 1 0 576 0 1 892
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_544_6
timestamp 1730954142
transform 1 0 576 0 1 892
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_543_6
timestamp 1730954142
transform 1 0 672 0 1 892
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_543_6
timestamp 1730954142
transform 1 0 672 0 1 892
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_546_6
timestamp 1730954142
transform 1 0 776 0 1 892
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_546_6
timestamp 1730954142
transform 1 0 776 0 1 892
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_547_6
timestamp 1730954142
transform 1 0 880 0 1 892
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_547_6
timestamp 1730954142
transform 1 0 880 0 1 892
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_52_6
timestamp 1730954142
transform 1 0 992 0 1 892
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_52_6
timestamp 1730954142
transform 1 0 992 0 1 892
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_51_6
timestamp 1730954142
transform 1 0 1080 0 1 892
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_51_6
timestamp 1730954142
transform 1 0 1080 0 1 892
box 7 3 85 69
use welltap_svt  __well_tap__21
timestamp 1730954142
transform 1 0 1176 0 1 912
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730954142
transform 1 0 1176 0 1 912
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_538_6
timestamp 1730954142
transform 1 0 136 0 -1 1044
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_538_6
timestamp 1730954142
transform 1 0 136 0 -1 1044
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_539_6
timestamp 1730954142
transform 1 0 264 0 -1 1044
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_539_6
timestamp 1730954142
transform 1 0 264 0 -1 1044
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_540_6
timestamp 1730954142
transform 1 0 408 0 -1 1044
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_540_6
timestamp 1730954142
transform 1 0 408 0 -1 1044
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_541_6
timestamp 1730954142
transform 1 0 568 0 -1 1044
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_541_6
timestamp 1730954142
transform 1 0 568 0 -1 1044
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_542_6
timestamp 1730954142
transform 1 0 736 0 -1 1044
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_542_6
timestamp 1730954142
transform 1 0 736 0 -1 1044
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_520_6
timestamp 1730954142
transform 1 0 920 0 -1 1044
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_520_6
timestamp 1730954142
transform 1 0 920 0 -1 1044
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_50_6
timestamp 1730954142
transform 1 0 1080 0 -1 1044
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_50_6
timestamp 1730954142
transform 1 0 1080 0 -1 1044
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_537_6
timestamp 1730954142
transform 1 0 128 0 1 1060
box 7 3 85 69
use welltap_svt  __well_tap__22
timestamp 1730954142
transform 1 0 104 0 -1 1024
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_537_6
timestamp 1730954142
transform 1 0 128 0 1 1060
box 7 3 85 69
use welltap_svt  __well_tap__22
timestamp 1730954142
transform 1 0 104 0 -1 1024
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_536_6
timestamp 1730954142
transform 1 0 240 0 1 1060
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_536_6
timestamp 1730954142
transform 1 0 240 0 1 1060
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_535_6
timestamp 1730954142
transform 1 0 400 0 1 1060
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_535_6
timestamp 1730954142
transform 1 0 400 0 1 1060
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_534_6
timestamp 1730954142
transform 1 0 568 0 1 1060
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_534_6
timestamp 1730954142
transform 1 0 568 0 1 1060
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_533_6
timestamp 1730954142
transform 1 0 752 0 1 1060
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_533_6
timestamp 1730954142
transform 1 0 752 0 1 1060
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_521_6
timestamp 1730954142
transform 1 0 936 0 1 1060
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_521_6
timestamp 1730954142
transform 1 0 936 0 1 1060
box 7 3 85 69
use welltap_svt  __well_tap__23
timestamp 1730954142
transform 1 0 1176 0 -1 1024
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1730954142
transform 1 0 1176 0 -1 1024
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730954142
transform 1 0 104 0 1 1080
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730954142
transform 1 0 104 0 1 1080
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1730954142
transform 1 0 1176 0 1 1080
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1730954142
transform 1 0 1176 0 1 1080
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730954142
transform 1 0 104 0 -1 1192
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730954142
transform 1 0 104 0 -1 1192
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_532_6
timestamp 1730954142
transform 1 0 352 0 -1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_532_6
timestamp 1730954142
transform 1 0 352 0 -1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_531_6
timestamp 1730954142
transform 1 0 440 0 -1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_531_6
timestamp 1730954142
transform 1 0 440 0 -1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_530_6
timestamp 1730954142
transform 1 0 536 0 -1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_530_6
timestamp 1730954142
transform 1 0 536 0 -1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_529_6
timestamp 1730954142
transform 1 0 632 0 -1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_529_6
timestamp 1730954142
transform 1 0 632 0 -1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_528_6
timestamp 1730954142
transform 1 0 736 0 -1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_528_6
timestamp 1730954142
transform 1 0 736 0 -1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_522_6
timestamp 1730954142
transform 1 0 840 0 -1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_522_6
timestamp 1730954142
transform 1 0 840 0 -1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_523_6
timestamp 1730954142
transform 1 0 944 0 -1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_523_6
timestamp 1730954142
transform 1 0 944 0 -1 1212
box 7 3 85 69
use welltap_svt  __well_tap__27
timestamp 1730954142
transform 1 0 1176 0 -1 1192
box 8 4 12 24
use welltap_svt  __well_tap__27
timestamp 1730954142
transform 1 0 1176 0 -1 1192
box 8 4 12 24
use welltap_svt  __well_tap__28
timestamp 1730954142
transform 1 0 104 0 1 1232
box 8 4 12 24
use welltap_svt  __well_tap__28
timestamp 1730954142
transform 1 0 104 0 1 1232
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_527_6
timestamp 1730954142
transform 1 0 648 0 1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_527_6
timestamp 1730954142
transform 1 0 648 0 1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_526_6
timestamp 1730954142
transform 1 0 736 0 1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_526_6
timestamp 1730954142
transform 1 0 736 0 1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_525_6
timestamp 1730954142
transform 1 0 824 0 1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_525_6
timestamp 1730954142
transform 1 0 824 0 1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_524_6
timestamp 1730954142
transform 1 0 912 0 1 1212
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_524_6
timestamp 1730954142
transform 1 0 912 0 1 1212
box 7 3 85 69
use welltap_svt  __well_tap__29
timestamp 1730954142
transform 1 0 1176 0 1 1232
box 8 4 12 24
use welltap_svt  __well_tap__29
timestamp 1730954142
transform 1 0 1176 0 1 1232
box 8 4 12 24
<< end >>
