magic
tech sky130l
timestamp 1731220469
<< m1 >>
rect 264 5663 268 5699
rect 2352 5487 2356 5527
rect 2560 5487 2564 5527
rect 2920 5487 2924 5527
rect 3112 5487 3116 5527
rect 3464 5487 3468 5527
rect 4384 5483 4388 5523
rect 4552 5483 4556 5523
rect 5016 5483 5020 5523
rect 1488 5363 1492 5403
rect 2648 5255 2652 5295
rect 3184 5255 3188 5295
rect 3520 5255 3524 5295
rect 1104 5215 1108 5251
rect 4480 5223 4484 5263
rect 4944 5223 4948 5263
rect 5128 5223 5132 5263
rect 752 5035 756 5075
rect 888 5035 892 5075
rect 1024 5035 1028 5075
rect 1424 5035 1428 5051
rect 2768 5031 2772 5103
rect 5248 4959 5252 4999
rect 4016 4791 4020 4827
rect 4256 4791 4260 4827
rect 5288 4791 5292 4827
rect 288 4647 292 4683
rect 2168 4599 2172 4635
rect 2576 4563 2580 4635
rect 4296 4563 4300 4599
rect 2344 4519 2348 4559
rect 2568 4519 2572 4559
rect 3400 4519 3404 4559
rect 3536 4519 3540 4559
rect 4648 4331 4652 4367
rect 5224 4331 5228 4367
rect 4040 4255 4044 4295
rect 2672 4123 2676 4159
rect 864 4079 868 4119
rect 2808 4123 2812 4159
rect 1000 4079 1004 4119
rect 4304 3995 4308 4067
rect 4496 3995 4500 4035
rect 4648 3995 4652 4035
rect 4800 3995 4804 4035
rect 4944 3995 4948 4035
rect 5088 3995 5092 4035
rect 5224 3995 5228 4035
rect 5376 3995 5380 4035
rect 2672 3875 2676 3911
rect 720 3803 724 3843
rect 2648 3635 2652 3671
rect 2848 3643 2852 3671
rect 3208 3635 3212 3671
rect 3408 3547 3412 3587
rect 3624 3547 3628 3587
rect 2744 3391 2748 3427
rect 2800 3323 2804 3427
rect 5040 3303 5044 3339
rect 4784 3227 4788 3267
rect 5512 3227 5516 3267
rect 856 3155 860 3191
rect 1784 3155 1788 3191
rect 2632 3127 2636 3163
rect 2992 3127 2996 3163
rect 3464 3039 3468 3079
rect 1304 2895 1308 2931
rect 2996 2835 3004 2839
rect 3000 2795 3004 2835
rect 4136 2835 4140 2871
rect 3992 2751 3996 2791
rect 584 2667 588 2703
rect 824 2667 828 2703
rect 976 2667 980 2703
rect 1520 2667 1524 2703
rect 1352 2591 1356 2631
rect 1672 2591 1676 2631
rect 2688 2555 2692 2595
rect 2960 2555 2964 2595
rect 3096 2555 3100 2595
rect 4080 2527 4084 2567
rect 4576 2527 4580 2567
rect 5072 2527 5076 2567
rect 512 2443 516 2479
rect 728 2443 732 2479
rect 1400 2407 1404 2479
rect 4440 2375 4444 2411
rect 2680 2299 2684 2339
rect 5144 2287 5148 2327
rect 592 2111 596 2151
rect 968 2111 972 2151
rect 1560 2111 1564 2151
rect 1784 2111 1788 2151
rect 3648 2143 3652 2179
rect 4848 2127 4852 2163
rect 800 1959 804 1995
rect 944 1959 948 1995
rect 376 1879 380 1919
rect 3232 1903 3236 1939
rect 3368 1903 3372 1939
rect 4968 1903 4972 1939
rect 5104 1903 5108 1939
rect 768 1723 772 1759
rect 1512 1723 1516 1759
rect 5240 1691 5244 1855
rect 5376 1815 5380 1899
rect 5512 1815 5516 1855
rect 4016 1651 4020 1687
rect 304 1375 308 1459
rect 536 1227 540 1263
rect 544 1227 548 1371
rect 2840 1323 2844 1363
rect 904 1227 908 1263
rect 1328 1139 1332 1179
rect 1648 1139 1652 1179
rect 3120 1151 3124 1187
rect 680 891 684 931
rect 2320 911 2324 947
rect 2328 831 2332 907
rect 2616 831 2620 871
rect 1008 695 1012 763
rect 1320 727 1324 763
rect 3992 659 3996 691
rect 1120 471 1124 539
rect 4432 503 4436 539
rect 5000 503 5004 539
rect 408 267 412 303
rect 808 195 812 303
rect 3624 243 3628 279
rect 5264 263 5268 299
rect 536 151 540 191
<< m2c >>
rect 256 5699 260 5703
rect 264 5699 268 5703
rect 392 5699 396 5703
rect 264 5659 268 5663
rect 2120 5599 2124 5603
rect 2280 5599 2284 5603
rect 2464 5599 2468 5603
rect 2648 5599 2652 5603
rect 2824 5599 2828 5603
rect 2992 5599 2996 5603
rect 3160 5599 3164 5603
rect 3320 5599 3324 5603
rect 3480 5599 3484 5603
rect 3640 5599 3644 5603
rect 3776 5599 3780 5603
rect 4432 5595 4436 5599
rect 4568 5595 4572 5599
rect 4704 5595 4708 5599
rect 4840 5595 4844 5599
rect 4976 5595 4980 5599
rect 5112 5595 5116 5599
rect 256 5583 260 5587
rect 400 5583 404 5587
rect 600 5583 604 5587
rect 824 5583 828 5587
rect 1080 5583 1084 5587
rect 1352 5583 1356 5587
rect 1640 5583 1644 5587
rect 1912 5583 1916 5587
rect 2352 5527 2356 5531
rect 2560 5527 2564 5531
rect 2920 5527 2924 5531
rect 3112 5527 3116 5531
rect 3464 5527 3468 5531
rect 4384 5523 4388 5527
rect 2264 5483 2268 5487
rect 2352 5483 2356 5487
rect 2480 5483 2484 5487
rect 2560 5483 2564 5487
rect 2688 5483 2692 5487
rect 2880 5483 2884 5487
rect 2920 5483 2924 5487
rect 3064 5483 3068 5487
rect 3112 5483 3116 5487
rect 3240 5483 3244 5487
rect 3416 5483 3420 5487
rect 3464 5483 3468 5487
rect 3592 5483 3596 5487
rect 3768 5483 3772 5487
rect 4552 5523 4556 5527
rect 5016 5523 5020 5527
rect 4376 5479 4380 5483
rect 4384 5479 4388 5483
rect 4528 5479 4532 5483
rect 4552 5479 4556 5483
rect 4680 5479 4684 5483
rect 4832 5479 4836 5483
rect 4984 5479 4988 5483
rect 5016 5479 5020 5483
rect 5144 5479 5148 5483
rect 376 5475 380 5479
rect 616 5475 620 5479
rect 864 5475 868 5479
rect 1112 5475 1116 5479
rect 1360 5475 1364 5479
rect 1608 5475 1612 5479
rect 1864 5475 1868 5479
rect 1488 5403 1492 5407
rect 2408 5367 2412 5371
rect 2608 5367 2612 5371
rect 2800 5367 2804 5371
rect 2984 5367 2988 5371
rect 3168 5367 3172 5371
rect 3344 5367 3348 5371
rect 3520 5367 3524 5371
rect 3704 5367 3708 5371
rect 536 5359 540 5363
rect 736 5359 740 5363
rect 944 5359 948 5363
rect 1160 5359 1164 5363
rect 1384 5359 1388 5363
rect 1488 5359 1492 5363
rect 1616 5359 1620 5363
rect 4376 5351 4380 5355
rect 4584 5352 4588 5356
rect 4792 5351 4796 5355
rect 5008 5351 5012 5355
rect 5224 5351 5228 5355
rect 2648 5295 2652 5299
rect 3184 5295 3188 5299
rect 3520 5295 3524 5299
rect 4480 5263 4484 5267
rect 688 5251 692 5255
rect 824 5251 828 5255
rect 960 5251 964 5255
rect 1096 5251 1100 5255
rect 1104 5251 1108 5255
rect 1232 5251 1236 5255
rect 1368 5251 1372 5255
rect 1504 5251 1508 5255
rect 1640 5251 1644 5255
rect 2320 5251 2324 5255
rect 2464 5251 2468 5255
rect 2616 5251 2620 5255
rect 2648 5251 2652 5255
rect 2776 5251 2780 5255
rect 2944 5251 2948 5255
rect 3128 5251 3132 5255
rect 3184 5251 3188 5255
rect 3312 5251 3316 5255
rect 3504 5251 3508 5255
rect 3520 5251 3524 5255
rect 3704 5251 3708 5255
rect 4944 5263 4948 5267
rect 5128 5263 5132 5267
rect 4376 5219 4380 5223
rect 4480 5219 4484 5223
rect 4608 5219 4612 5223
rect 4840 5219 4844 5223
rect 4944 5219 4948 5223
rect 5072 5219 5076 5223
rect 5128 5219 5132 5223
rect 5312 5219 5316 5223
rect 1104 5211 1108 5215
rect 2120 5143 2124 5147
rect 2256 5143 2260 5147
rect 2424 5143 2428 5147
rect 2608 5143 2612 5147
rect 2792 5143 2796 5147
rect 2984 5143 2988 5147
rect 3184 5143 3188 5147
rect 3384 5143 3388 5147
rect 3592 5143 3596 5147
rect 3776 5143 3780 5147
rect 2768 5103 2772 5107
rect 752 5075 756 5079
rect 888 5075 892 5079
rect 1024 5075 1028 5079
rect 1424 5051 1428 5055
rect 472 5031 476 5035
rect 608 5031 612 5035
rect 744 5031 748 5035
rect 752 5031 756 5035
rect 880 5031 884 5035
rect 888 5031 892 5035
rect 1016 5031 1020 5035
rect 1024 5031 1028 5035
rect 1160 5031 1164 5035
rect 1312 5031 1316 5035
rect 1424 5031 1428 5035
rect 1464 5031 1468 5035
rect 1616 5031 1620 5035
rect 1776 5031 1780 5035
rect 1912 5031 1916 5035
rect 3984 5083 3988 5087
rect 4232 5083 4236 5087
rect 4504 5083 4508 5087
rect 4776 5083 4780 5087
rect 5056 5083 5060 5087
rect 5336 5083 5340 5087
rect 3864 5031 3868 5035
rect 2120 5027 2124 5031
rect 2656 5027 2660 5031
rect 2768 5027 2772 5031
rect 3224 5027 3228 5031
rect 3776 5027 3780 5031
rect 5248 4999 5252 5003
rect 3984 4955 3988 4959
rect 4144 4955 4148 4959
rect 4336 4955 4340 4959
rect 4536 4955 4540 4959
rect 4752 4955 4756 4959
rect 4968 4955 4972 4959
rect 5192 4955 5196 4959
rect 5248 4955 5252 4959
rect 5424 4955 5428 4959
rect 256 4923 260 4927
rect 440 4923 444 4927
rect 648 4923 652 4927
rect 848 4923 852 4927
rect 1040 4923 1044 4927
rect 1224 4923 1228 4927
rect 1408 4923 1412 4927
rect 1584 4923 1588 4927
rect 1760 4923 1764 4927
rect 1912 4923 1916 4927
rect 2968 4887 2972 4891
rect 3104 4887 3108 4891
rect 3984 4827 3988 4831
rect 4016 4827 4020 4831
rect 4168 4827 4172 4831
rect 4256 4827 4260 4831
rect 4384 4827 4388 4831
rect 4608 4827 4612 4831
rect 4832 4827 4836 4831
rect 5056 4827 5060 4831
rect 5280 4827 5284 4831
rect 5288 4827 5292 4831
rect 5504 4827 5508 4831
rect 256 4799 260 4803
rect 392 4799 396 4803
rect 528 4799 532 4803
rect 664 4799 668 4803
rect 800 4799 804 4803
rect 4016 4787 4020 4791
rect 4256 4787 4260 4791
rect 5288 4787 5292 4791
rect 2120 4747 2124 4751
rect 2280 4747 2284 4751
rect 2472 4747 2476 4751
rect 2664 4747 2668 4751
rect 2856 4747 2860 4751
rect 3056 4747 3060 4751
rect 3256 4747 3260 4751
rect 4040 4707 4044 4711
rect 4312 4707 4316 4711
rect 4592 4707 4596 4711
rect 4888 4707 4892 4711
rect 5192 4707 5196 4711
rect 5496 4707 5500 4711
rect 256 4683 260 4687
rect 288 4683 292 4687
rect 440 4683 444 4687
rect 664 4683 668 4687
rect 904 4683 908 4687
rect 1152 4683 1156 4687
rect 1408 4683 1412 4687
rect 1672 4683 1676 4687
rect 1912 4683 1916 4687
rect 288 4643 292 4647
rect 2120 4635 2124 4639
rect 2168 4635 2172 4639
rect 2336 4635 2340 4639
rect 2568 4635 2572 4639
rect 2576 4635 2580 4639
rect 2792 4635 2796 4639
rect 3016 4635 3020 4639
rect 3240 4635 3244 4639
rect 3464 4635 3468 4639
rect 2168 4595 2172 4599
rect 4160 4599 4164 4603
rect 4296 4599 4300 4603
rect 4424 4599 4428 4603
rect 4696 4599 4700 4603
rect 4968 4599 4972 4603
rect 5248 4599 5252 4603
rect 5536 4599 5540 4603
rect 2344 4559 2348 4563
rect 296 4551 300 4555
rect 520 4551 524 4555
rect 768 4551 772 4555
rect 1032 4551 1036 4555
rect 1320 4551 1324 4555
rect 1616 4551 1620 4555
rect 1912 4551 1916 4555
rect 2568 4559 2572 4563
rect 2576 4559 2580 4563
rect 3400 4559 3404 4563
rect 3536 4559 3540 4563
rect 4296 4559 4300 4563
rect 2224 4515 2228 4519
rect 2344 4515 2348 4519
rect 2472 4515 2476 4519
rect 2568 4515 2572 4519
rect 2704 4515 2708 4519
rect 2920 4515 2924 4519
rect 3128 4515 3132 4519
rect 3328 4515 3332 4519
rect 3400 4515 3404 4519
rect 3528 4515 3532 4519
rect 3536 4515 3540 4519
rect 3736 4515 3740 4519
rect 4304 4483 4308 4487
rect 4536 4483 4540 4487
rect 4784 4483 4788 4487
rect 5040 4483 5044 4487
rect 5304 4483 5308 4487
rect 5568 4483 5572 4487
rect 544 4439 548 4443
rect 752 4439 756 4443
rect 984 4439 988 4443
rect 1240 4439 1244 4443
rect 1504 4439 1508 4443
rect 1776 4439 1780 4443
rect 2328 4399 2332 4403
rect 2544 4399 2548 4403
rect 2760 4399 2764 4403
rect 2968 4399 2972 4403
rect 3176 4399 3180 4403
rect 3384 4399 3388 4403
rect 3592 4399 3596 4403
rect 3776 4399 3780 4403
rect 4456 4367 4460 4371
rect 4616 4367 4620 4371
rect 4648 4367 4652 4371
rect 4784 4367 4788 4371
rect 4976 4367 4980 4371
rect 5176 4367 5180 4371
rect 5224 4367 5228 4371
rect 5384 4367 5388 4371
rect 5600 4367 5604 4371
rect 4648 4327 4652 4331
rect 5224 4327 5228 4331
rect 792 4319 796 4323
rect 936 4319 940 4323
rect 1088 4319 1092 4323
rect 1248 4319 1252 4323
rect 1416 4319 1420 4323
rect 1592 4319 1596 4323
rect 1776 4319 1780 4323
rect 4040 4295 4044 4299
rect 2432 4275 2436 4279
rect 2584 4275 2588 4279
rect 2752 4275 2756 4279
rect 2936 4275 2940 4279
rect 3136 4275 3140 4279
rect 3352 4275 3356 4279
rect 3576 4275 3580 4279
rect 3776 4275 3780 4279
rect 3984 4251 3988 4255
rect 4040 4251 4044 4255
rect 4168 4251 4172 4255
rect 4376 4251 4380 4255
rect 4600 4251 4604 4255
rect 4840 4251 4844 4255
rect 5096 4251 5100 4255
rect 5360 4251 5364 4255
rect 5624 4251 5628 4255
rect 912 4195 916 4199
rect 1048 4195 1052 4199
rect 1184 4195 1188 4199
rect 1320 4195 1324 4199
rect 1456 4195 1460 4199
rect 1592 4195 1596 4199
rect 1728 4195 1732 4199
rect 1864 4195 1868 4199
rect 2664 4159 2668 4163
rect 2672 4159 2676 4163
rect 2800 4159 2804 4163
rect 2808 4159 2812 4163
rect 2936 4159 2940 4163
rect 3072 4159 3076 4163
rect 864 4119 868 4123
rect 1000 4119 1004 4123
rect 2672 4119 2676 4123
rect 2808 4119 2812 4123
rect 3984 4107 3988 4111
rect 4512 4107 4516 4111
rect 5072 4107 5076 4111
rect 5640 4107 5644 4111
rect 856 4075 860 4079
rect 864 4075 868 4079
rect 992 4075 996 4079
rect 1000 4075 1004 4079
rect 1128 4075 1132 4079
rect 1264 4075 1268 4079
rect 1400 4075 1404 4079
rect 1536 4075 1540 4079
rect 1672 4075 1676 4079
rect 4304 4067 4308 4071
rect 2416 4023 2420 4027
rect 2552 4023 2556 4027
rect 2688 4023 2692 4027
rect 2824 4023 2828 4027
rect 2960 4023 2964 4027
rect 4496 4035 4500 4039
rect 4648 4035 4652 4039
rect 4800 4035 4804 4039
rect 4944 4035 4948 4039
rect 5088 4035 5092 4039
rect 5224 4035 5228 4039
rect 5376 4035 5380 4039
rect 3984 3991 3988 3995
rect 4128 3991 4132 3995
rect 4296 3991 4300 3995
rect 4304 3991 4308 3995
rect 4464 3991 4468 3995
rect 4496 3991 4500 3995
rect 4624 3991 4628 3995
rect 4648 3991 4652 3995
rect 4776 3991 4780 3995
rect 4800 3991 4804 3995
rect 4928 3991 4932 3995
rect 4944 3991 4948 3995
rect 5072 3991 5076 3995
rect 5088 3991 5092 3995
rect 5216 3991 5220 3995
rect 5224 3991 5228 3995
rect 5360 3991 5364 3995
rect 5376 3991 5380 3995
rect 5504 3991 5508 3995
rect 5640 3991 5644 3995
rect 608 3943 612 3947
rect 760 3943 764 3947
rect 920 3943 924 3947
rect 1080 3943 1084 3947
rect 1248 3943 1252 3947
rect 1416 3943 1420 3947
rect 2216 3911 2220 3915
rect 2424 3911 2428 3915
rect 2632 3911 2636 3915
rect 2672 3911 2676 3915
rect 2840 3911 2844 3915
rect 3040 3911 3044 3915
rect 3232 3911 3236 3915
rect 3416 3911 3420 3915
rect 3608 3911 3612 3915
rect 3776 3911 3780 3915
rect 2672 3871 2676 3875
rect 4480 3859 4484 3863
rect 4696 3859 4700 3863
rect 4920 3859 4924 3863
rect 5160 3859 5164 3863
rect 5408 3860 5412 3864
rect 5640 3859 5644 3863
rect 720 3843 724 3847
rect 256 3799 260 3803
rect 432 3799 436 3803
rect 640 3799 644 3803
rect 720 3799 724 3803
rect 848 3799 852 3803
rect 1064 3799 1068 3803
rect 1288 3799 1292 3803
rect 2264 3783 2268 3787
rect 2496 3783 2500 3787
rect 2712 3783 2716 3787
rect 2920 3783 2924 3787
rect 3120 3783 3124 3787
rect 3320 3783 3324 3787
rect 3528 3783 3532 3787
rect 4120 3727 4124 3731
rect 4328 3727 4332 3731
rect 4560 3727 4564 3731
rect 4816 3727 4820 3731
rect 5088 3727 5092 3731
rect 5376 3727 5380 3731
rect 5640 3727 5644 3731
rect 256 3691 260 3695
rect 432 3691 436 3695
rect 624 3691 628 3695
rect 808 3691 812 3695
rect 984 3691 988 3695
rect 1152 3691 1156 3695
rect 1312 3691 1316 3695
rect 1464 3691 1468 3695
rect 1616 3691 1620 3695
rect 1776 3691 1780 3695
rect 1912 3691 1916 3695
rect 2376 3671 2380 3675
rect 2576 3671 2580 3675
rect 2648 3671 2652 3675
rect 2776 3671 2780 3675
rect 2848 3671 2852 3675
rect 2976 3671 2980 3675
rect 3176 3671 3180 3675
rect 3208 3671 3212 3675
rect 3376 3671 3380 3675
rect 2848 3639 2852 3643
rect 2648 3631 2652 3635
rect 3208 3631 3212 3635
rect 4312 3591 4316 3595
rect 4496 3591 4500 3595
rect 4704 3591 4708 3595
rect 4928 3591 4932 3595
rect 5168 3591 5172 3595
rect 5416 3591 5420 3595
rect 5640 3591 5644 3595
rect 3408 3587 3412 3591
rect 272 3563 276 3567
rect 480 3563 484 3567
rect 696 3563 700 3567
rect 928 3563 932 3567
rect 1168 3563 1172 3567
rect 1416 3563 1420 3567
rect 1672 3563 1676 3567
rect 1912 3563 1916 3567
rect 3624 3587 3628 3591
rect 2120 3543 2124 3547
rect 2376 3543 2380 3547
rect 2640 3543 2644 3547
rect 2880 3543 2884 3547
rect 3104 3543 3108 3547
rect 3320 3543 3324 3547
rect 3408 3543 3412 3547
rect 3536 3543 3540 3547
rect 3624 3543 3628 3547
rect 3752 3543 3756 3547
rect 4656 3451 4660 3455
rect 4808 3451 4812 3455
rect 4968 3451 4972 3455
rect 5128 3451 5132 3455
rect 5296 3451 5300 3455
rect 5472 3451 5476 3455
rect 5640 3451 5644 3455
rect 400 3431 404 3435
rect 544 3431 548 3435
rect 696 3431 700 3435
rect 856 3431 860 3435
rect 1032 3431 1036 3435
rect 1208 3431 1212 3435
rect 1392 3431 1396 3435
rect 1584 3431 1588 3435
rect 2120 3427 2124 3431
rect 2288 3427 2292 3431
rect 2496 3427 2500 3431
rect 2712 3427 2716 3431
rect 2744 3427 2748 3431
rect 2744 3387 2748 3391
rect 2800 3427 2804 3431
rect 2928 3427 2932 3431
rect 3144 3427 3148 3431
rect 3360 3427 3364 3431
rect 3576 3427 3580 3431
rect 3776 3427 3780 3431
rect 3984 3339 3988 3343
rect 4248 3339 4252 3343
rect 4520 3339 4524 3343
rect 4768 3339 4772 3343
rect 4992 3339 4996 3343
rect 5040 3339 5044 3343
rect 5208 3339 5212 3343
rect 5424 3339 5428 3343
rect 5640 3339 5644 3343
rect 2800 3319 2804 3323
rect 592 3299 596 3303
rect 792 3299 796 3303
rect 1000 3299 1004 3303
rect 1216 3299 1220 3303
rect 1440 3299 1444 3303
rect 5040 3299 5044 3303
rect 2120 3271 2124 3275
rect 2320 3271 2324 3275
rect 2536 3271 2540 3275
rect 2744 3271 2748 3275
rect 2936 3271 2940 3275
rect 3128 3271 3132 3275
rect 3312 3271 3316 3275
rect 3496 3271 3500 3275
rect 3680 3271 3684 3275
rect 4784 3267 4788 3271
rect 5512 3267 5516 3271
rect 3984 3223 3988 3227
rect 4224 3223 4228 3227
rect 4472 3223 4476 3227
rect 4704 3223 4708 3227
rect 4784 3223 4788 3227
rect 4912 3223 4916 3227
rect 5112 3223 5116 3227
rect 5296 3223 5300 3227
rect 5480 3223 5484 3227
rect 5512 3223 5516 3227
rect 5640 3223 5644 3227
rect 632 3191 636 3195
rect 824 3191 828 3195
rect 856 3191 860 3195
rect 1016 3191 1020 3195
rect 1208 3191 1212 3195
rect 1392 3191 1396 3195
rect 1568 3191 1572 3195
rect 1752 3191 1756 3195
rect 1784 3191 1788 3195
rect 1912 3191 1916 3195
rect 856 3151 860 3155
rect 2560 3163 2564 3167
rect 2632 3163 2636 3167
rect 2760 3163 2764 3167
rect 2960 3163 2964 3167
rect 2992 3163 2996 3167
rect 3152 3163 3156 3167
rect 3336 3163 3340 3167
rect 3528 3163 3532 3167
rect 3720 3163 3724 3167
rect 1784 3151 1788 3155
rect 2632 3123 2636 3127
rect 2992 3123 2996 3127
rect 4000 3099 4004 3103
rect 4232 3099 4236 3103
rect 4456 3099 4460 3103
rect 4680 3099 4684 3103
rect 4904 3099 4908 3103
rect 5128 3099 5132 3103
rect 3464 3079 3468 3083
rect 552 3067 556 3071
rect 688 3067 692 3071
rect 824 3067 828 3071
rect 960 3067 964 3071
rect 1096 3067 1100 3071
rect 1232 3067 1236 3071
rect 1368 3067 1372 3071
rect 1504 3067 1508 3071
rect 1640 3067 1644 3071
rect 1776 3067 1780 3071
rect 1912 3067 1916 3071
rect 2456 3035 2460 3039
rect 2680 3035 2684 3039
rect 2904 3035 2908 3039
rect 3128 3035 3132 3039
rect 3360 3035 3364 3039
rect 3464 3035 3468 3039
rect 3592 3035 3596 3039
rect 4032 2983 4036 2987
rect 4200 2983 4204 2987
rect 4368 2983 4372 2987
rect 4536 2983 4540 2987
rect 4704 2983 4708 2987
rect 4880 2983 4884 2987
rect 296 2931 300 2935
rect 608 2931 612 2935
rect 912 2931 916 2935
rect 1208 2931 1212 2935
rect 1304 2931 1308 2935
rect 1512 2931 1516 2935
rect 1816 2931 1820 2935
rect 2240 2915 2244 2919
rect 2440 2915 2444 2919
rect 2640 2915 2644 2919
rect 2840 2915 2844 2919
rect 3032 2915 3036 2919
rect 3232 2915 3236 2919
rect 3432 2915 3436 2919
rect 1304 2891 1308 2895
rect 3992 2871 3996 2875
rect 4128 2871 4132 2875
rect 4136 2871 4140 2875
rect 4264 2871 4268 2875
rect 4400 2871 4404 2875
rect 4536 2871 4540 2875
rect 4672 2871 4676 2875
rect 2992 2835 2996 2839
rect 256 2815 260 2819
rect 432 2815 436 2819
rect 648 2815 652 2819
rect 888 2815 892 2819
rect 1136 2815 1140 2819
rect 1400 2815 1404 2819
rect 1664 2815 1668 2819
rect 4136 2831 4140 2835
rect 2136 2791 2140 2795
rect 2384 2791 2388 2795
rect 2632 2791 2636 2795
rect 2880 2791 2884 2795
rect 3000 2791 3004 2795
rect 3128 2791 3132 2795
rect 3992 2791 3996 2795
rect 3984 2747 3988 2751
rect 3992 2747 3996 2751
rect 4120 2747 4124 2751
rect 4256 2747 4260 2751
rect 4392 2747 4396 2751
rect 4528 2747 4532 2751
rect 4664 2747 4668 2751
rect 4800 2747 4804 2751
rect 4936 2747 4940 2751
rect 376 2703 380 2707
rect 552 2703 556 2707
rect 584 2703 588 2707
rect 744 2703 748 2707
rect 824 2703 828 2707
rect 952 2703 956 2707
rect 976 2703 980 2707
rect 1176 2703 1180 2707
rect 1408 2703 1412 2707
rect 1520 2703 1524 2707
rect 1648 2703 1652 2707
rect 1896 2703 1900 2707
rect 584 2663 588 2667
rect 824 2663 828 2667
rect 976 2663 980 2667
rect 2120 2679 2124 2683
rect 2344 2679 2348 2683
rect 2600 2679 2604 2683
rect 2856 2679 2860 2683
rect 3112 2679 3116 2683
rect 1520 2663 1524 2667
rect 4056 2639 4060 2643
rect 4352 2639 4356 2643
rect 4640 2639 4644 2643
rect 4920 2639 4924 2643
rect 5208 2639 5212 2643
rect 5496 2639 5500 2643
rect 1352 2631 1356 2635
rect 1672 2631 1676 2635
rect 2688 2595 2692 2599
rect 696 2587 700 2591
rect 856 2587 860 2591
rect 1016 2587 1020 2591
rect 1168 2587 1172 2591
rect 1320 2587 1324 2591
rect 1352 2587 1356 2591
rect 1480 2587 1484 2591
rect 1640 2587 1644 2591
rect 1672 2587 1676 2591
rect 1800 2587 1804 2591
rect 2960 2595 2964 2599
rect 3096 2595 3100 2599
rect 4080 2567 4084 2571
rect 2680 2551 2684 2555
rect 2688 2551 2692 2555
rect 2816 2551 2820 2555
rect 2952 2551 2956 2555
rect 2960 2551 2964 2555
rect 3088 2551 3092 2555
rect 3096 2551 3100 2555
rect 3224 2551 3228 2555
rect 4576 2567 4580 2571
rect 5072 2567 5076 2571
rect 3984 2523 3988 2527
rect 4080 2523 4084 2527
rect 4208 2523 4212 2527
rect 4456 2523 4460 2527
rect 4576 2523 4580 2527
rect 4704 2523 4708 2527
rect 4952 2523 4956 2527
rect 5072 2523 5076 2527
rect 5200 2523 5204 2527
rect 5448 2523 5452 2527
rect 480 2479 484 2483
rect 512 2479 516 2483
rect 696 2479 700 2483
rect 728 2479 732 2483
rect 912 2479 916 2483
rect 1120 2479 1124 2483
rect 1328 2479 1332 2483
rect 1400 2479 1404 2483
rect 1528 2479 1532 2483
rect 1728 2479 1732 2483
rect 1912 2479 1916 2483
rect 512 2439 516 2443
rect 728 2439 732 2443
rect 2120 2419 2124 2423
rect 2320 2419 2324 2423
rect 2544 2419 2548 2423
rect 2776 2419 2780 2423
rect 3024 2419 3028 2423
rect 3280 2419 3284 2423
rect 3536 2419 3540 2423
rect 3776 2419 3780 2423
rect 3984 2411 3988 2415
rect 4184 2411 4188 2415
rect 4424 2411 4428 2415
rect 4440 2411 4444 2415
rect 4680 2411 4684 2415
rect 4944 2411 4948 2415
rect 5216 2411 5220 2415
rect 5496 2411 5500 2415
rect 1400 2403 1404 2407
rect 4440 2371 4444 2375
rect 2000 2367 2004 2371
rect 352 2359 356 2363
rect 648 2359 652 2363
rect 960 2359 964 2363
rect 1280 2359 1284 2363
rect 1608 2359 1612 2363
rect 1912 2359 1916 2363
rect 2680 2339 2684 2343
rect 5144 2327 5148 2331
rect 2120 2295 2124 2299
rect 2280 2295 2284 2299
rect 2472 2295 2476 2299
rect 2664 2295 2668 2299
rect 2680 2295 2684 2299
rect 2856 2295 2860 2299
rect 3048 2295 3052 2299
rect 3240 2295 3244 2299
rect 3424 2295 3428 2299
rect 3608 2295 3612 2299
rect 3776 2295 3780 2299
rect 4568 2283 4572 2287
rect 4736 2283 4740 2287
rect 4912 2284 4916 2288
rect 5088 2283 5092 2287
rect 5144 2283 5148 2287
rect 5272 2283 5276 2287
rect 5464 2283 5468 2287
rect 5640 2283 5644 2287
rect 256 2235 260 2239
rect 464 2235 468 2239
rect 696 2235 700 2239
rect 928 2235 932 2239
rect 1160 2235 1164 2239
rect 2120 2179 2124 2183
rect 2288 2179 2292 2183
rect 2456 2179 2460 2183
rect 2632 2179 2636 2183
rect 2808 2179 2812 2183
rect 2976 2179 2980 2183
rect 3144 2179 3148 2183
rect 3304 2179 3308 2183
rect 3464 2179 3468 2183
rect 3632 2179 3636 2183
rect 3648 2179 3652 2183
rect 3776 2179 3780 2183
rect 592 2151 596 2155
rect 968 2151 972 2155
rect 1560 2151 1564 2155
rect 1784 2151 1788 2155
rect 4640 2163 4644 2167
rect 4816 2163 4820 2167
rect 4848 2163 4852 2167
rect 5008 2163 5012 2167
rect 5216 2163 5220 2167
rect 5432 2163 5436 2167
rect 5640 2163 5644 2167
rect 3648 2139 3652 2143
rect 4848 2123 4852 2127
rect 256 2107 260 2111
rect 472 2107 476 2111
rect 592 2107 596 2111
rect 720 2107 724 2111
rect 960 2107 964 2111
rect 968 2107 972 2111
rect 1200 2107 1204 2111
rect 1440 2107 1444 2111
rect 1560 2107 1564 2111
rect 1688 2107 1692 2111
rect 1784 2107 1788 2111
rect 1912 2107 1916 2111
rect 3232 2047 3236 2051
rect 3368 2047 3372 2051
rect 3504 2047 3508 2051
rect 3640 2047 3644 2051
rect 3776 2047 3780 2051
rect 4760 2047 4764 2051
rect 4896 2047 4900 2051
rect 5032 2047 5036 2051
rect 5168 2047 5172 2051
rect 5304 2047 5308 2051
rect 368 1995 372 1999
rect 504 1995 508 1999
rect 640 1995 644 1999
rect 784 1995 788 1999
rect 800 1995 804 1999
rect 928 1995 932 1999
rect 944 1995 948 1999
rect 1072 1995 1076 1999
rect 1216 1995 1220 1999
rect 1360 1995 1364 1999
rect 1504 1995 1508 1999
rect 1640 1995 1644 1999
rect 1776 1995 1780 1999
rect 1912 1995 1916 1999
rect 800 1955 804 1959
rect 944 1955 948 1959
rect 3224 1939 3228 1943
rect 3232 1939 3236 1943
rect 3360 1939 3364 1943
rect 3368 1939 3372 1943
rect 3496 1939 3500 1943
rect 3632 1939 3636 1943
rect 3768 1939 3772 1943
rect 4960 1939 4964 1943
rect 4968 1939 4972 1943
rect 5096 1939 5100 1943
rect 5104 1939 5108 1943
rect 5232 1939 5236 1943
rect 5368 1939 5372 1943
rect 5504 1939 5508 1943
rect 5640 1939 5644 1943
rect 376 1919 380 1923
rect 3232 1899 3236 1903
rect 3368 1899 3372 1903
rect 4968 1899 4972 1903
rect 5104 1899 5108 1903
rect 5376 1899 5380 1903
rect 312 1875 316 1879
rect 376 1875 380 1879
rect 504 1875 508 1879
rect 712 1875 716 1879
rect 936 1875 940 1879
rect 1176 1875 1180 1879
rect 1424 1875 1428 1879
rect 1680 1875 1684 1879
rect 1912 1875 1916 1879
rect 5240 1855 5244 1859
rect 2120 1811 2124 1815
rect 2352 1811 2356 1815
rect 2592 1811 2596 1815
rect 2816 1811 2820 1815
rect 3032 1811 3036 1815
rect 3232 1811 3236 1815
rect 3424 1811 3428 1815
rect 3608 1811 3612 1815
rect 3776 1811 3780 1815
rect 4800 1811 4804 1815
rect 4944 1811 4948 1815
rect 5088 1811 5092 1815
rect 5232 1811 5236 1815
rect 256 1759 260 1763
rect 472 1759 476 1763
rect 688 1759 692 1763
rect 768 1759 772 1763
rect 896 1759 900 1763
rect 1096 1759 1100 1763
rect 1288 1759 1292 1763
rect 1480 1759 1484 1763
rect 1512 1759 1516 1763
rect 1672 1759 1676 1763
rect 768 1719 772 1723
rect 1512 1719 1516 1723
rect 2120 1695 2124 1699
rect 2256 1695 2260 1699
rect 2408 1695 2412 1699
rect 2568 1695 2572 1699
rect 2736 1695 2740 1699
rect 2904 1695 2908 1699
rect 3072 1695 3076 1699
rect 3248 1695 3252 1699
rect 5512 1855 5516 1859
rect 5368 1811 5372 1815
rect 5376 1811 5380 1815
rect 5504 1811 5508 1815
rect 5512 1811 5516 1815
rect 5640 1811 5644 1815
rect 3984 1687 3988 1691
rect 4016 1687 4020 1691
rect 4176 1687 4180 1691
rect 4400 1687 4404 1691
rect 4632 1687 4636 1691
rect 4872 1687 4876 1691
rect 5120 1687 5124 1691
rect 5240 1687 5244 1691
rect 5376 1687 5380 1691
rect 5632 1687 5636 1691
rect 4016 1647 4020 1651
rect 256 1619 260 1623
rect 520 1619 524 1623
rect 808 1619 812 1623
rect 1104 1619 1108 1623
rect 1400 1619 1404 1623
rect 2216 1571 2220 1575
rect 2352 1571 2356 1575
rect 2488 1571 2492 1575
rect 2624 1571 2628 1575
rect 2760 1571 2764 1575
rect 2896 1571 2900 1575
rect 3032 1571 3036 1575
rect 3168 1571 3172 1575
rect 3304 1571 3308 1575
rect 3984 1571 3988 1575
rect 4120 1571 4124 1575
rect 4280 1571 4284 1575
rect 4480 1571 4484 1575
rect 4712 1571 4716 1575
rect 4976 1571 4980 1575
rect 5256 1571 5260 1575
rect 5544 1571 5548 1575
rect 256 1499 260 1503
rect 472 1499 476 1503
rect 704 1499 708 1503
rect 936 1499 940 1503
rect 1168 1499 1172 1503
rect 1400 1499 1404 1503
rect 3984 1463 3988 1467
rect 4120 1463 4124 1467
rect 4256 1463 4260 1467
rect 4400 1463 4404 1467
rect 4592 1463 4596 1467
rect 4816 1463 4820 1467
rect 5064 1463 5068 1467
rect 5320 1463 5324 1467
rect 5584 1463 5588 1467
rect 304 1459 308 1463
rect 2120 1443 2124 1447
rect 2256 1443 2260 1447
rect 2392 1443 2396 1447
rect 2528 1443 2532 1447
rect 2664 1443 2668 1447
rect 2800 1443 2804 1447
rect 2936 1443 2940 1447
rect 3072 1443 3076 1447
rect 256 1371 260 1375
rect 304 1371 308 1375
rect 536 1371 540 1375
rect 544 1371 548 1375
rect 864 1371 868 1375
rect 1216 1371 1220 1375
rect 1576 1371 1580 1375
rect 1912 1371 1916 1375
rect 2000 1371 2004 1375
rect 256 1263 260 1267
rect 456 1263 460 1267
rect 536 1263 540 1267
rect 536 1223 540 1227
rect 2840 1363 2844 1367
rect 3984 1343 3988 1347
rect 4184 1343 4188 1347
rect 4432 1343 4436 1347
rect 4704 1343 4708 1347
rect 5000 1343 5004 1347
rect 5312 1343 5316 1347
rect 5624 1343 5628 1347
rect 2120 1319 2124 1323
rect 2400 1319 2404 1323
rect 2688 1319 2692 1323
rect 2840 1319 2844 1323
rect 2968 1319 2972 1323
rect 3248 1319 3252 1323
rect 3520 1319 3524 1323
rect 3776 1319 3780 1323
rect 672 1263 676 1267
rect 872 1263 876 1267
rect 904 1263 908 1267
rect 1064 1263 1068 1267
rect 1248 1263 1252 1267
rect 1424 1263 1428 1267
rect 1592 1263 1596 1267
rect 1760 1263 1764 1267
rect 1912 1263 1916 1267
rect 544 1223 548 1227
rect 4712 1227 4716 1231
rect 4888 1227 4892 1231
rect 5072 1227 5076 1231
rect 5264 1227 5268 1231
rect 5464 1227 5468 1231
rect 5640 1227 5644 1231
rect 904 1223 908 1227
rect 2752 1187 2756 1191
rect 2928 1187 2932 1191
rect 3104 1187 3108 1191
rect 3120 1187 3124 1191
rect 3280 1187 3284 1191
rect 3456 1187 3460 1191
rect 3640 1187 3644 1191
rect 1328 1179 1332 1183
rect 1648 1179 1652 1183
rect 3120 1147 3124 1151
rect 256 1135 260 1139
rect 416 1135 420 1139
rect 600 1135 604 1139
rect 784 1135 788 1139
rect 960 1135 964 1139
rect 1128 1135 1132 1139
rect 1296 1135 1300 1139
rect 1328 1135 1332 1139
rect 1456 1135 1460 1139
rect 1616 1135 1620 1139
rect 1648 1135 1652 1139
rect 1776 1135 1780 1139
rect 1912 1135 1916 1139
rect 4960 1107 4964 1111
rect 5096 1107 5100 1111
rect 5232 1107 5236 1111
rect 5368 1107 5372 1111
rect 5504 1107 5508 1111
rect 5640 1107 5644 1111
rect 2120 1055 2124 1059
rect 2296 1055 2300 1059
rect 2488 1055 2492 1059
rect 2672 1055 2676 1059
rect 2848 1055 2852 1059
rect 3016 1055 3020 1059
rect 3184 1055 3188 1059
rect 3344 1055 3348 1059
rect 3512 1055 3516 1059
rect 272 1015 276 1019
rect 528 1015 532 1019
rect 784 1015 788 1019
rect 1048 1015 1052 1019
rect 1312 1015 1316 1019
rect 4904 995 4908 999
rect 5040 995 5044 999
rect 5176 995 5180 999
rect 5312 995 5316 999
rect 5448 995 5452 999
rect 5584 995 5588 999
rect 2120 947 2124 951
rect 2288 947 2292 951
rect 2320 947 2324 951
rect 2472 947 2476 951
rect 2664 947 2668 951
rect 2856 947 2860 951
rect 3040 947 3044 951
rect 3224 947 3228 951
rect 3408 947 3412 951
rect 3592 947 3596 951
rect 3776 947 3780 951
rect 680 931 684 935
rect 2320 907 2324 911
rect 2328 907 2332 911
rect 360 887 364 891
rect 584 887 588 891
rect 680 887 684 891
rect 808 887 812 891
rect 1032 887 1036 891
rect 1256 887 1260 891
rect 1488 887 1492 891
rect 3984 875 3988 879
rect 4120 875 4124 879
rect 4296 875 4300 879
rect 4512 875 4516 879
rect 4768 875 4772 879
rect 5056 875 5060 879
rect 5360 875 5364 879
rect 5640 875 5644 879
rect 2616 871 2620 875
rect 2120 827 2124 831
rect 2304 827 2308 831
rect 2328 827 2332 831
rect 2528 827 2532 831
rect 2616 827 2620 831
rect 2800 827 2804 831
rect 3112 827 3116 831
rect 3448 827 3452 831
rect 3776 827 3780 831
rect 3984 767 3988 771
rect 4120 767 4124 771
rect 4256 767 4260 771
rect 4392 767 4396 771
rect 4528 767 4532 771
rect 4664 767 4668 771
rect 4816 767 4820 771
rect 4992 767 4996 771
rect 5184 767 5188 771
rect 5384 767 5388 771
rect 5584 767 5588 771
rect 272 763 276 767
rect 528 763 532 767
rect 768 763 772 767
rect 1000 763 1004 767
rect 1008 763 1012 767
rect 1224 763 1228 767
rect 1320 763 1324 767
rect 1448 763 1452 767
rect 1672 763 1676 767
rect 1320 723 1324 727
rect 1008 691 1012 695
rect 3992 691 3996 695
rect 3992 655 3996 659
rect 256 647 260 651
rect 440 647 444 651
rect 648 647 652 651
rect 848 647 852 651
rect 1032 647 1036 651
rect 1208 647 1212 651
rect 1384 647 1388 651
rect 1552 647 1556 651
rect 1720 647 1724 651
rect 1896 647 1900 651
rect 3984 647 3988 651
rect 4120 647 4124 651
rect 4256 647 4260 651
rect 4392 647 4396 651
rect 4528 647 4532 651
rect 4664 647 4668 651
rect 4824 647 4828 651
rect 5016 647 5020 651
rect 5224 647 5228 651
rect 5440 647 5444 651
rect 5640 647 5644 651
rect 256 539 260 543
rect 472 539 476 543
rect 696 539 700 543
rect 904 539 908 543
rect 1096 539 1100 543
rect 1120 539 1124 543
rect 1272 539 1276 543
rect 1440 539 1444 543
rect 1608 539 1612 543
rect 1768 539 1772 543
rect 1912 539 1916 543
rect 3984 539 3988 543
rect 4168 539 4172 543
rect 4408 539 4412 543
rect 4432 539 4436 543
rect 4672 539 4676 543
rect 4952 539 4956 543
rect 5000 539 5004 543
rect 5248 539 5252 543
rect 5544 539 5548 543
rect 3232 519 3236 523
rect 3368 519 3372 523
rect 3504 519 3508 523
rect 3640 519 3644 523
rect 3776 519 3780 523
rect 4432 499 4436 503
rect 5000 499 5004 503
rect 1120 467 1124 471
rect 280 423 284 427
rect 608 423 612 427
rect 936 423 940 427
rect 1264 423 1268 427
rect 1600 423 1604 427
rect 1912 423 1916 427
rect 4576 411 4580 415
rect 4768 411 4772 415
rect 4968 411 4972 415
rect 5176 411 5180 415
rect 5392 411 5396 415
rect 5608 411 5612 415
rect 2120 403 2124 407
rect 2328 403 2332 407
rect 2552 403 2556 407
rect 2776 403 2780 407
rect 2984 403 2988 407
rect 3192 403 3196 407
rect 3392 403 3396 407
rect 3592 403 3596 407
rect 3776 403 3780 407
rect 376 303 380 307
rect 408 303 412 307
rect 584 303 588 307
rect 800 303 804 307
rect 808 303 812 307
rect 1016 303 1020 307
rect 1232 303 1236 307
rect 408 263 412 267
rect 4712 299 4716 303
rect 4872 299 4876 303
rect 5048 299 5052 303
rect 5232 299 5236 303
rect 5264 299 5268 303
rect 5424 299 5428 303
rect 5624 299 5628 303
rect 2120 279 2124 283
rect 2256 279 2260 283
rect 2392 279 2396 283
rect 2528 279 2532 283
rect 2664 279 2668 283
rect 2800 279 2804 283
rect 2936 279 2940 283
rect 3072 279 3076 283
rect 3208 279 3212 283
rect 3344 279 3348 283
rect 3480 279 3484 283
rect 3616 279 3620 283
rect 3624 279 3628 283
rect 3752 279 3756 283
rect 5264 259 5268 263
rect 3624 239 3628 243
rect 536 191 540 195
rect 808 191 812 195
rect 256 147 260 151
rect 392 147 396 151
rect 528 147 532 151
rect 536 147 540 151
rect 664 147 668 151
rect 800 147 804 151
rect 936 147 940 151
rect 1072 147 1076 151
rect 1208 147 1212 151
rect 4416 143 4420 147
rect 4552 143 4556 147
rect 4688 143 4692 147
rect 4824 143 4828 147
rect 4960 143 4964 147
rect 5096 143 5100 147
rect 5232 143 5236 147
rect 5368 143 5372 147
rect 5640 143 5644 147
rect 2120 127 2124 131
rect 2256 127 2260 131
rect 2392 127 2396 131
rect 2528 127 2532 131
rect 2664 127 2668 131
rect 2800 127 2804 131
rect 2936 127 2940 131
rect 3072 127 3076 131
rect 3208 127 3212 131
rect 3344 127 3348 131
rect 3480 127 3484 131
rect 3616 127 3620 131
rect 3752 127 3756 131
<< m2 >>
rect 110 5729 116 5730
rect 1934 5729 1940 5730
rect 110 5725 111 5729
rect 115 5725 116 5729
rect 110 5724 116 5725
rect 158 5728 164 5729
rect 158 5724 159 5728
rect 163 5724 164 5728
rect 158 5723 164 5724
rect 294 5728 300 5729
rect 294 5724 295 5728
rect 299 5724 300 5728
rect 1934 5725 1935 5729
rect 1939 5725 1940 5729
rect 1934 5724 1940 5725
rect 294 5723 300 5724
rect 130 5713 136 5714
rect 110 5712 116 5713
rect 110 5708 111 5712
rect 115 5708 116 5712
rect 130 5709 131 5713
rect 135 5709 136 5713
rect 130 5708 136 5709
rect 266 5713 272 5714
rect 266 5709 267 5713
rect 271 5709 272 5713
rect 266 5708 272 5709
rect 1934 5712 1940 5713
rect 1934 5708 1935 5712
rect 1939 5708 1940 5712
rect 110 5707 116 5708
rect 1934 5707 1940 5708
rect 255 5703 261 5704
rect 255 5699 256 5703
rect 260 5702 261 5703
rect 263 5703 269 5704
rect 263 5702 264 5703
rect 260 5700 264 5702
rect 260 5699 261 5700
rect 255 5698 261 5699
rect 263 5699 264 5700
rect 268 5699 269 5703
rect 263 5698 269 5699
rect 378 5703 384 5704
rect 378 5699 379 5703
rect 383 5702 384 5703
rect 391 5703 397 5704
rect 391 5702 392 5703
rect 383 5700 392 5702
rect 383 5699 384 5700
rect 378 5698 384 5699
rect 391 5699 392 5700
rect 396 5699 397 5703
rect 391 5698 397 5699
rect 263 5663 269 5664
rect 263 5659 264 5663
rect 268 5662 269 5663
rect 268 5660 273 5662
rect 268 5659 269 5660
rect 263 5658 269 5659
rect 378 5635 384 5636
rect 378 5634 379 5635
rect 259 5632 379 5634
rect 259 5630 261 5632
rect 378 5631 379 5632
rect 383 5631 384 5635
rect 378 5630 384 5631
rect 1778 5631 1784 5632
rect 1778 5630 1779 5631
rect 229 5628 261 5630
rect 1613 5628 1779 5630
rect 282 5627 288 5628
rect 282 5623 283 5627
rect 287 5623 288 5627
rect 282 5622 288 5623
rect 482 5627 488 5628
rect 482 5623 483 5627
rect 487 5623 488 5627
rect 482 5622 488 5623
rect 706 5627 712 5628
rect 706 5623 707 5627
rect 711 5623 712 5627
rect 706 5622 712 5623
rect 962 5627 968 5628
rect 962 5623 963 5627
rect 967 5623 968 5627
rect 962 5622 968 5623
rect 1234 5627 1240 5628
rect 1234 5623 1235 5627
rect 1239 5623 1240 5627
rect 1778 5627 1779 5628
rect 1783 5627 1784 5631
rect 1974 5629 1980 5630
rect 3798 5629 3804 5630
rect 1778 5626 1784 5627
rect 1794 5627 1800 5628
rect 1234 5622 1240 5623
rect 1794 5623 1795 5627
rect 1799 5623 1800 5627
rect 1974 5625 1975 5629
rect 1979 5625 1980 5629
rect 1974 5624 1980 5625
rect 2022 5628 2028 5629
rect 2022 5624 2023 5628
rect 2027 5624 2028 5628
rect 2022 5623 2028 5624
rect 2182 5628 2188 5629
rect 2182 5624 2183 5628
rect 2187 5624 2188 5628
rect 2182 5623 2188 5624
rect 2366 5628 2372 5629
rect 2366 5624 2367 5628
rect 2371 5624 2372 5628
rect 2366 5623 2372 5624
rect 2550 5628 2556 5629
rect 2550 5624 2551 5628
rect 2555 5624 2556 5628
rect 2550 5623 2556 5624
rect 2726 5628 2732 5629
rect 2726 5624 2727 5628
rect 2731 5624 2732 5628
rect 2726 5623 2732 5624
rect 2894 5628 2900 5629
rect 2894 5624 2895 5628
rect 2899 5624 2900 5628
rect 2894 5623 2900 5624
rect 3062 5628 3068 5629
rect 3062 5624 3063 5628
rect 3067 5624 3068 5628
rect 3062 5623 3068 5624
rect 3222 5628 3228 5629
rect 3222 5624 3223 5628
rect 3227 5624 3228 5628
rect 3222 5623 3228 5624
rect 3382 5628 3388 5629
rect 3382 5624 3383 5628
rect 3387 5624 3388 5628
rect 3382 5623 3388 5624
rect 3542 5628 3548 5629
rect 3542 5624 3543 5628
rect 3547 5624 3548 5628
rect 3542 5623 3548 5624
rect 3678 5628 3684 5629
rect 3678 5624 3679 5628
rect 3683 5624 3684 5628
rect 3798 5625 3799 5629
rect 3803 5625 3804 5629
rect 3798 5624 3804 5625
rect 3838 5625 3844 5626
rect 5662 5625 5668 5626
rect 3678 5623 3684 5624
rect 1794 5622 1800 5623
rect 3838 5621 3839 5625
rect 3843 5621 3844 5625
rect 3838 5620 3844 5621
rect 4334 5624 4340 5625
rect 4334 5620 4335 5624
rect 4339 5620 4340 5624
rect 4334 5619 4340 5620
rect 4470 5624 4476 5625
rect 4470 5620 4471 5624
rect 4475 5620 4476 5624
rect 4470 5619 4476 5620
rect 4606 5624 4612 5625
rect 4606 5620 4607 5624
rect 4611 5620 4612 5624
rect 4606 5619 4612 5620
rect 4742 5624 4748 5625
rect 4742 5620 4743 5624
rect 4747 5620 4748 5624
rect 4742 5619 4748 5620
rect 4878 5624 4884 5625
rect 4878 5620 4879 5624
rect 4883 5620 4884 5624
rect 4878 5619 4884 5620
rect 5014 5624 5020 5625
rect 5014 5620 5015 5624
rect 5019 5620 5020 5624
rect 5662 5621 5663 5625
rect 5667 5621 5668 5625
rect 5662 5620 5668 5621
rect 5014 5619 5020 5620
rect 1994 5613 2000 5614
rect 1974 5612 1980 5613
rect 1974 5608 1975 5612
rect 1979 5608 1980 5612
rect 1994 5609 1995 5613
rect 1999 5609 2000 5613
rect 1994 5608 2000 5609
rect 2154 5613 2160 5614
rect 2154 5609 2155 5613
rect 2159 5609 2160 5613
rect 2154 5608 2160 5609
rect 2338 5613 2344 5614
rect 2338 5609 2339 5613
rect 2343 5609 2344 5613
rect 2338 5608 2344 5609
rect 2522 5613 2528 5614
rect 2522 5609 2523 5613
rect 2527 5609 2528 5613
rect 2522 5608 2528 5609
rect 2698 5613 2704 5614
rect 2698 5609 2699 5613
rect 2703 5609 2704 5613
rect 2698 5608 2704 5609
rect 2866 5613 2872 5614
rect 2866 5609 2867 5613
rect 2871 5609 2872 5613
rect 2866 5608 2872 5609
rect 3034 5613 3040 5614
rect 3034 5609 3035 5613
rect 3039 5609 3040 5613
rect 3034 5608 3040 5609
rect 3194 5613 3200 5614
rect 3194 5609 3195 5613
rect 3199 5609 3200 5613
rect 3194 5608 3200 5609
rect 3354 5613 3360 5614
rect 3354 5609 3355 5613
rect 3359 5609 3360 5613
rect 3354 5608 3360 5609
rect 3514 5613 3520 5614
rect 3514 5609 3515 5613
rect 3519 5609 3520 5613
rect 3514 5608 3520 5609
rect 3650 5613 3656 5614
rect 3650 5609 3651 5613
rect 3655 5609 3656 5613
rect 3650 5608 3656 5609
rect 3798 5612 3804 5613
rect 3798 5608 3799 5612
rect 3803 5608 3804 5612
rect 4306 5609 4312 5610
rect 1974 5607 1980 5608
rect 3798 5607 3804 5608
rect 3838 5608 3844 5609
rect 3838 5604 3839 5608
rect 3843 5604 3844 5608
rect 4306 5605 4307 5609
rect 4311 5605 4312 5609
rect 4306 5604 4312 5605
rect 4442 5609 4448 5610
rect 4442 5605 4443 5609
rect 4447 5605 4448 5609
rect 4442 5604 4448 5605
rect 4578 5609 4584 5610
rect 4578 5605 4579 5609
rect 4583 5605 4584 5609
rect 4578 5604 4584 5605
rect 4714 5609 4720 5610
rect 4714 5605 4715 5609
rect 4719 5605 4720 5609
rect 4714 5604 4720 5605
rect 4850 5609 4856 5610
rect 4850 5605 4851 5609
rect 4855 5605 4856 5609
rect 4850 5604 4856 5605
rect 4986 5609 4992 5610
rect 4986 5605 4987 5609
rect 4991 5605 4992 5609
rect 4986 5604 4992 5605
rect 5662 5608 5668 5609
rect 5662 5604 5663 5608
rect 5667 5604 5668 5608
rect 2119 5603 2125 5604
rect 2119 5599 2120 5603
rect 2124 5602 2125 5603
rect 2142 5603 2148 5604
rect 2142 5602 2143 5603
rect 2124 5600 2143 5602
rect 2124 5599 2125 5600
rect 2119 5598 2125 5599
rect 2142 5599 2143 5600
rect 2147 5599 2148 5603
rect 2142 5598 2148 5599
rect 2279 5603 2288 5604
rect 2279 5599 2280 5603
rect 2287 5599 2288 5603
rect 2279 5598 2288 5599
rect 2463 5603 2472 5604
rect 2463 5599 2464 5603
rect 2471 5599 2472 5603
rect 2463 5598 2472 5599
rect 2646 5603 2653 5604
rect 2646 5599 2647 5603
rect 2652 5599 2653 5603
rect 2646 5598 2653 5599
rect 2823 5603 2832 5604
rect 2823 5599 2824 5603
rect 2831 5599 2832 5603
rect 2823 5598 2832 5599
rect 2991 5603 3000 5604
rect 2991 5599 2992 5603
rect 2999 5599 3000 5603
rect 2991 5598 3000 5599
rect 3159 5603 3165 5604
rect 3159 5599 3160 5603
rect 3164 5602 3165 5603
rect 3182 5603 3188 5604
rect 3182 5602 3183 5603
rect 3164 5600 3183 5602
rect 3164 5599 3165 5600
rect 3159 5598 3165 5599
rect 3182 5599 3183 5600
rect 3187 5599 3188 5603
rect 3182 5598 3188 5599
rect 3319 5603 3325 5604
rect 3319 5599 3320 5603
rect 3324 5602 3325 5603
rect 3342 5603 3348 5604
rect 3342 5602 3343 5603
rect 3324 5600 3343 5602
rect 3324 5599 3325 5600
rect 3319 5598 3325 5599
rect 3342 5599 3343 5600
rect 3347 5599 3348 5603
rect 3342 5598 3348 5599
rect 3479 5603 3485 5604
rect 3479 5599 3480 5603
rect 3484 5602 3485 5603
rect 3502 5603 3508 5604
rect 3502 5602 3503 5603
rect 3484 5600 3503 5602
rect 3484 5599 3485 5600
rect 3479 5598 3485 5599
rect 3502 5599 3503 5600
rect 3507 5599 3508 5603
rect 3502 5598 3508 5599
rect 3639 5603 3648 5604
rect 3639 5599 3640 5603
rect 3647 5599 3648 5603
rect 3639 5598 3648 5599
rect 3738 5603 3744 5604
rect 3738 5599 3739 5603
rect 3743 5602 3744 5603
rect 3775 5603 3781 5604
rect 3838 5603 3844 5604
rect 5662 5603 5668 5604
rect 3775 5602 3776 5603
rect 3743 5600 3776 5602
rect 3743 5599 3744 5600
rect 3738 5598 3744 5599
rect 3775 5599 3776 5600
rect 3780 5599 3781 5603
rect 3775 5598 3781 5599
rect 4431 5599 4440 5600
rect 4431 5595 4432 5599
rect 4439 5595 4440 5599
rect 4431 5594 4440 5595
rect 4567 5599 4576 5600
rect 4567 5595 4568 5599
rect 4575 5595 4576 5599
rect 4567 5594 4576 5595
rect 4703 5599 4712 5600
rect 4703 5595 4704 5599
rect 4711 5595 4712 5599
rect 4703 5594 4712 5595
rect 4839 5599 4848 5600
rect 4839 5595 4840 5599
rect 4847 5595 4848 5599
rect 4839 5594 4848 5595
rect 4975 5599 4984 5600
rect 4975 5595 4976 5599
rect 4983 5595 4984 5599
rect 4975 5594 4984 5595
rect 5110 5599 5117 5600
rect 5110 5595 5111 5599
rect 5116 5595 5117 5599
rect 5110 5594 5117 5595
rect 255 5587 261 5588
rect 255 5583 256 5587
rect 260 5586 261 5587
rect 282 5587 288 5588
rect 282 5586 283 5587
rect 260 5584 283 5586
rect 260 5583 261 5584
rect 255 5582 261 5583
rect 282 5583 283 5584
rect 287 5583 288 5587
rect 282 5582 288 5583
rect 399 5587 405 5588
rect 399 5583 400 5587
rect 404 5586 405 5587
rect 482 5587 488 5588
rect 482 5586 483 5587
rect 404 5584 483 5586
rect 404 5583 405 5584
rect 399 5582 405 5583
rect 482 5583 483 5584
rect 487 5583 488 5587
rect 482 5582 488 5583
rect 599 5587 605 5588
rect 599 5583 600 5587
rect 604 5586 605 5587
rect 706 5587 712 5588
rect 706 5586 707 5587
rect 604 5584 707 5586
rect 604 5583 605 5584
rect 599 5582 605 5583
rect 706 5583 707 5584
rect 711 5583 712 5587
rect 706 5582 712 5583
rect 823 5587 829 5588
rect 823 5583 824 5587
rect 828 5586 829 5587
rect 962 5587 968 5588
rect 962 5586 963 5587
rect 828 5584 963 5586
rect 828 5583 829 5584
rect 823 5582 829 5583
rect 962 5583 963 5584
rect 967 5583 968 5587
rect 962 5582 968 5583
rect 1079 5587 1085 5588
rect 1079 5583 1080 5587
rect 1084 5586 1085 5587
rect 1234 5587 1240 5588
rect 1234 5586 1235 5587
rect 1084 5584 1235 5586
rect 1084 5583 1085 5584
rect 1079 5582 1085 5583
rect 1234 5583 1235 5584
rect 1239 5583 1240 5587
rect 1234 5582 1240 5583
rect 1278 5587 1284 5588
rect 1278 5583 1279 5587
rect 1283 5586 1284 5587
rect 1351 5587 1357 5588
rect 1351 5586 1352 5587
rect 1283 5584 1352 5586
rect 1283 5583 1284 5584
rect 1278 5582 1284 5583
rect 1351 5583 1352 5584
rect 1356 5583 1357 5587
rect 1351 5582 1357 5583
rect 1639 5587 1645 5588
rect 1639 5583 1640 5587
rect 1644 5586 1645 5587
rect 1794 5587 1800 5588
rect 1794 5586 1795 5587
rect 1644 5584 1795 5586
rect 1644 5583 1645 5584
rect 1639 5582 1645 5583
rect 1794 5583 1795 5584
rect 1799 5583 1800 5587
rect 1794 5582 1800 5583
rect 1911 5587 1917 5588
rect 1911 5583 1912 5587
rect 1916 5586 1917 5587
rect 1962 5587 1968 5588
rect 1962 5586 1963 5587
rect 1916 5584 1963 5586
rect 1916 5583 1917 5584
rect 1911 5582 1917 5583
rect 1962 5583 1963 5584
rect 1967 5583 1968 5587
rect 1962 5582 1968 5583
rect 110 5580 116 5581
rect 1934 5580 1940 5581
rect 110 5576 111 5580
rect 115 5576 116 5580
rect 110 5575 116 5576
rect 130 5579 136 5580
rect 130 5575 131 5579
rect 135 5575 136 5579
rect 130 5574 136 5575
rect 274 5579 280 5580
rect 274 5575 275 5579
rect 279 5575 280 5579
rect 274 5574 280 5575
rect 474 5579 480 5580
rect 474 5575 475 5579
rect 479 5575 480 5579
rect 474 5574 480 5575
rect 698 5579 704 5580
rect 698 5575 699 5579
rect 703 5575 704 5579
rect 698 5574 704 5575
rect 954 5579 960 5580
rect 954 5575 955 5579
rect 959 5575 960 5579
rect 954 5574 960 5575
rect 1226 5579 1232 5580
rect 1226 5575 1227 5579
rect 1231 5575 1232 5579
rect 1226 5574 1232 5575
rect 1514 5579 1520 5580
rect 1514 5575 1515 5579
rect 1519 5575 1520 5579
rect 1514 5574 1520 5575
rect 1786 5579 1792 5580
rect 1786 5575 1787 5579
rect 1791 5575 1792 5579
rect 1934 5576 1935 5580
rect 1939 5576 1940 5580
rect 1934 5575 1940 5576
rect 1786 5574 1792 5575
rect 158 5564 164 5565
rect 110 5563 116 5564
rect 110 5559 111 5563
rect 115 5559 116 5563
rect 158 5560 159 5564
rect 163 5560 164 5564
rect 158 5559 164 5560
rect 302 5564 308 5565
rect 302 5560 303 5564
rect 307 5560 308 5564
rect 302 5559 308 5560
rect 502 5564 508 5565
rect 502 5560 503 5564
rect 507 5560 508 5564
rect 502 5559 508 5560
rect 726 5564 732 5565
rect 726 5560 727 5564
rect 731 5560 732 5564
rect 726 5559 732 5560
rect 982 5564 988 5565
rect 982 5560 983 5564
rect 987 5560 988 5564
rect 982 5559 988 5560
rect 1254 5564 1260 5565
rect 1254 5560 1255 5564
rect 1259 5560 1260 5564
rect 1254 5559 1260 5560
rect 1542 5564 1548 5565
rect 1542 5560 1543 5564
rect 1547 5560 1548 5564
rect 1542 5559 1548 5560
rect 1814 5564 1820 5565
rect 1814 5560 1815 5564
rect 1819 5560 1820 5564
rect 1814 5559 1820 5560
rect 1934 5563 1940 5564
rect 1934 5559 1935 5563
rect 1939 5559 1940 5563
rect 110 5558 116 5559
rect 1934 5558 1940 5559
rect 1962 5563 1968 5564
rect 1962 5559 1963 5563
rect 1967 5562 1968 5563
rect 2142 5563 2148 5564
rect 1967 5560 2001 5562
rect 1967 5559 1968 5560
rect 1962 5558 1968 5559
rect 2142 5559 2143 5563
rect 2147 5562 2148 5563
rect 2282 5563 2288 5564
rect 2147 5560 2161 5562
rect 2147 5559 2148 5560
rect 2142 5558 2148 5559
rect 2282 5559 2283 5563
rect 2287 5562 2288 5563
rect 2466 5563 2472 5564
rect 2287 5560 2345 5562
rect 2287 5559 2288 5560
rect 2282 5558 2288 5559
rect 2466 5559 2467 5563
rect 2471 5562 2472 5563
rect 2794 5563 2800 5564
rect 2471 5560 2529 5562
rect 2471 5559 2472 5560
rect 2466 5558 2472 5559
rect 2794 5559 2795 5563
rect 2799 5559 2800 5563
rect 2794 5558 2800 5559
rect 2826 5563 2832 5564
rect 2826 5559 2827 5563
rect 2831 5562 2832 5563
rect 2994 5563 3000 5564
rect 2831 5560 2873 5562
rect 2831 5559 2832 5560
rect 2826 5558 2832 5559
rect 2994 5559 2995 5563
rect 2999 5562 3000 5563
rect 3182 5563 3188 5564
rect 2999 5560 3041 5562
rect 2999 5559 3000 5560
rect 2994 5558 3000 5559
rect 3182 5559 3183 5563
rect 3187 5562 3188 5563
rect 3342 5563 3348 5564
rect 3187 5560 3201 5562
rect 3187 5559 3188 5560
rect 3182 5558 3188 5559
rect 3342 5559 3343 5563
rect 3347 5562 3348 5563
rect 3502 5563 3508 5564
rect 3347 5560 3361 5562
rect 3347 5559 3348 5560
rect 3342 5558 3348 5559
rect 3502 5559 3503 5563
rect 3507 5562 3508 5563
rect 3642 5563 3648 5564
rect 3507 5560 3521 5562
rect 3507 5559 3508 5560
rect 3502 5558 3508 5559
rect 3642 5559 3643 5563
rect 3647 5562 3648 5563
rect 3647 5560 3657 5562
rect 3647 5559 3648 5560
rect 3642 5558 3648 5559
rect 4374 5559 4380 5560
rect 4374 5555 4375 5559
rect 4379 5555 4380 5559
rect 4374 5554 4380 5555
rect 4434 5559 4440 5560
rect 4434 5555 4435 5559
rect 4439 5558 4440 5559
rect 4570 5559 4576 5560
rect 4439 5556 4449 5558
rect 4439 5555 4440 5556
rect 4434 5554 4440 5555
rect 4570 5555 4571 5559
rect 4575 5558 4576 5559
rect 4706 5559 4712 5560
rect 4575 5556 4585 5558
rect 4575 5555 4576 5556
rect 4570 5554 4576 5555
rect 4706 5555 4707 5559
rect 4711 5558 4712 5559
rect 4842 5559 4848 5560
rect 4711 5556 4721 5558
rect 4711 5555 4712 5556
rect 4706 5554 4712 5555
rect 4842 5555 4843 5559
rect 4847 5558 4848 5559
rect 4978 5559 4984 5560
rect 4847 5556 4857 5558
rect 4847 5555 4848 5556
rect 4842 5554 4848 5555
rect 4978 5555 4979 5559
rect 4983 5558 4984 5559
rect 4983 5556 4993 5558
rect 4983 5555 4984 5556
rect 4978 5554 4984 5555
rect 2351 5531 2357 5532
rect 2351 5530 2352 5531
rect 2237 5528 2352 5530
rect 2351 5527 2352 5528
rect 2356 5527 2357 5531
rect 2559 5531 2565 5532
rect 2559 5530 2560 5531
rect 2453 5528 2560 5530
rect 2351 5526 2357 5527
rect 2559 5527 2560 5528
rect 2564 5527 2565 5531
rect 2559 5526 2565 5527
rect 2646 5531 2652 5532
rect 2646 5527 2647 5531
rect 2651 5527 2652 5531
rect 2919 5531 2925 5532
rect 2919 5530 2920 5531
rect 2853 5528 2920 5530
rect 2646 5526 2652 5527
rect 2919 5527 2920 5528
rect 2924 5527 2925 5531
rect 3111 5531 3117 5532
rect 3111 5530 3112 5531
rect 3037 5528 3112 5530
rect 2919 5526 2925 5527
rect 3111 5527 3112 5528
rect 3116 5527 3117 5531
rect 3111 5526 3117 5527
rect 3166 5531 3172 5532
rect 3166 5527 3167 5531
rect 3171 5527 3172 5531
rect 3463 5531 3469 5532
rect 3463 5530 3464 5531
rect 3389 5528 3464 5530
rect 3166 5526 3172 5527
rect 3463 5527 3464 5528
rect 3468 5527 3469 5531
rect 3634 5531 3640 5532
rect 3634 5530 3635 5531
rect 3565 5528 3635 5530
rect 3463 5526 3469 5527
rect 3634 5527 3635 5528
rect 3639 5527 3640 5531
rect 3634 5526 3640 5527
rect 3738 5531 3744 5532
rect 3738 5527 3739 5531
rect 3743 5527 3744 5531
rect 3738 5526 3744 5527
rect 4383 5527 4389 5528
rect 4383 5526 4384 5527
rect 4349 5524 4384 5526
rect 4383 5523 4384 5524
rect 4388 5523 4389 5527
rect 4551 5527 4557 5528
rect 4551 5526 4552 5527
rect 4501 5524 4552 5526
rect 4383 5522 4389 5523
rect 4551 5523 4552 5524
rect 4556 5523 4557 5527
rect 4551 5522 4557 5523
rect 4574 5527 4580 5528
rect 4574 5523 4575 5527
rect 4579 5523 4580 5527
rect 4850 5527 4856 5528
rect 4850 5526 4851 5527
rect 4805 5524 4851 5526
rect 4574 5522 4580 5523
rect 4850 5523 4851 5524
rect 4855 5523 4856 5527
rect 5015 5527 5021 5528
rect 5015 5526 5016 5527
rect 4957 5524 5016 5526
rect 4850 5522 4856 5523
rect 5015 5523 5016 5524
rect 5020 5523 5021 5527
rect 5015 5522 5021 5523
rect 5110 5527 5116 5528
rect 5110 5523 5111 5527
rect 5115 5523 5116 5527
rect 5110 5522 5116 5523
rect 110 5505 116 5506
rect 1934 5505 1940 5506
rect 110 5501 111 5505
rect 115 5501 116 5505
rect 110 5500 116 5501
rect 278 5504 284 5505
rect 278 5500 279 5504
rect 283 5500 284 5504
rect 278 5499 284 5500
rect 518 5504 524 5505
rect 518 5500 519 5504
rect 523 5500 524 5504
rect 518 5499 524 5500
rect 766 5504 772 5505
rect 766 5500 767 5504
rect 771 5500 772 5504
rect 766 5499 772 5500
rect 1014 5504 1020 5505
rect 1014 5500 1015 5504
rect 1019 5500 1020 5504
rect 1014 5499 1020 5500
rect 1262 5504 1268 5505
rect 1262 5500 1263 5504
rect 1267 5500 1268 5504
rect 1262 5499 1268 5500
rect 1510 5504 1516 5505
rect 1510 5500 1511 5504
rect 1515 5500 1516 5504
rect 1510 5499 1516 5500
rect 1766 5504 1772 5505
rect 1766 5500 1767 5504
rect 1771 5500 1772 5504
rect 1934 5501 1935 5505
rect 1939 5501 1940 5505
rect 1934 5500 1940 5501
rect 1766 5499 1772 5500
rect 250 5489 256 5490
rect 110 5488 116 5489
rect 110 5484 111 5488
rect 115 5484 116 5488
rect 250 5485 251 5489
rect 255 5485 256 5489
rect 250 5484 256 5485
rect 490 5489 496 5490
rect 490 5485 491 5489
rect 495 5485 496 5489
rect 490 5484 496 5485
rect 738 5489 744 5490
rect 738 5485 739 5489
rect 743 5485 744 5489
rect 738 5484 744 5485
rect 986 5489 992 5490
rect 986 5485 987 5489
rect 991 5485 992 5489
rect 986 5484 992 5485
rect 1234 5489 1240 5490
rect 1234 5485 1235 5489
rect 1239 5485 1240 5489
rect 1234 5484 1240 5485
rect 1482 5489 1488 5490
rect 1482 5485 1483 5489
rect 1487 5485 1488 5489
rect 1482 5484 1488 5485
rect 1738 5489 1744 5490
rect 1738 5485 1739 5489
rect 1743 5485 1744 5489
rect 1738 5484 1744 5485
rect 1934 5488 1940 5489
rect 1934 5484 1935 5488
rect 1939 5484 1940 5488
rect 110 5483 116 5484
rect 1934 5483 1940 5484
rect 2262 5487 2269 5488
rect 2262 5483 2263 5487
rect 2268 5483 2269 5487
rect 2262 5482 2269 5483
rect 2351 5487 2357 5488
rect 2351 5483 2352 5487
rect 2356 5486 2357 5487
rect 2479 5487 2485 5488
rect 2479 5486 2480 5487
rect 2356 5484 2480 5486
rect 2356 5483 2357 5484
rect 2351 5482 2357 5483
rect 2479 5483 2480 5484
rect 2484 5483 2485 5487
rect 2479 5482 2485 5483
rect 2559 5487 2565 5488
rect 2559 5483 2560 5487
rect 2564 5486 2565 5487
rect 2687 5487 2693 5488
rect 2687 5486 2688 5487
rect 2564 5484 2688 5486
rect 2564 5483 2565 5484
rect 2559 5482 2565 5483
rect 2687 5483 2688 5484
rect 2692 5483 2693 5487
rect 2687 5482 2693 5483
rect 2794 5487 2800 5488
rect 2794 5483 2795 5487
rect 2799 5486 2800 5487
rect 2879 5487 2885 5488
rect 2879 5486 2880 5487
rect 2799 5484 2880 5486
rect 2799 5483 2800 5484
rect 2794 5482 2800 5483
rect 2879 5483 2880 5484
rect 2884 5483 2885 5487
rect 2879 5482 2885 5483
rect 2919 5487 2925 5488
rect 2919 5483 2920 5487
rect 2924 5486 2925 5487
rect 3063 5487 3069 5488
rect 3063 5486 3064 5487
rect 2924 5484 3064 5486
rect 2924 5483 2925 5484
rect 2919 5482 2925 5483
rect 3063 5483 3064 5484
rect 3068 5483 3069 5487
rect 3063 5482 3069 5483
rect 3111 5487 3117 5488
rect 3111 5483 3112 5487
rect 3116 5486 3117 5487
rect 3239 5487 3245 5488
rect 3239 5486 3240 5487
rect 3116 5484 3240 5486
rect 3116 5483 3117 5484
rect 3111 5482 3117 5483
rect 3239 5483 3240 5484
rect 3244 5483 3245 5487
rect 3239 5482 3245 5483
rect 3326 5487 3332 5488
rect 3326 5483 3327 5487
rect 3331 5486 3332 5487
rect 3415 5487 3421 5488
rect 3415 5486 3416 5487
rect 3331 5484 3416 5486
rect 3331 5483 3332 5484
rect 3326 5482 3332 5483
rect 3415 5483 3416 5484
rect 3420 5483 3421 5487
rect 3415 5482 3421 5483
rect 3463 5487 3469 5488
rect 3463 5483 3464 5487
rect 3468 5486 3469 5487
rect 3591 5487 3597 5488
rect 3591 5486 3592 5487
rect 3468 5484 3592 5486
rect 3468 5483 3469 5484
rect 3463 5482 3469 5483
rect 3591 5483 3592 5484
rect 3596 5483 3597 5487
rect 3591 5482 3597 5483
rect 3634 5487 3640 5488
rect 3634 5483 3635 5487
rect 3639 5486 3640 5487
rect 3767 5487 3773 5488
rect 3767 5486 3768 5487
rect 3639 5484 3768 5486
rect 3639 5483 3640 5484
rect 3634 5482 3640 5483
rect 3767 5483 3768 5484
rect 3772 5483 3773 5487
rect 3767 5482 3773 5483
rect 4374 5483 4381 5484
rect 1974 5480 1980 5481
rect 3798 5480 3804 5481
rect 375 5479 384 5480
rect 375 5475 376 5479
rect 383 5475 384 5479
rect 375 5474 384 5475
rect 615 5479 624 5480
rect 615 5475 616 5479
rect 623 5475 624 5479
rect 615 5474 624 5475
rect 863 5479 872 5480
rect 863 5475 864 5479
rect 871 5475 872 5479
rect 1111 5479 1117 5480
rect 1111 5478 1112 5479
rect 863 5474 872 5475
rect 1099 5476 1112 5478
rect 506 5471 512 5472
rect 506 5467 507 5471
rect 511 5470 512 5471
rect 1099 5470 1101 5476
rect 1111 5475 1112 5476
rect 1116 5475 1117 5479
rect 1111 5474 1117 5475
rect 1359 5479 1368 5480
rect 1359 5475 1360 5479
rect 1367 5475 1368 5479
rect 1359 5474 1368 5475
rect 1607 5479 1616 5480
rect 1607 5475 1608 5479
rect 1615 5475 1616 5479
rect 1607 5474 1616 5475
rect 1778 5479 1784 5480
rect 1778 5475 1779 5479
rect 1783 5478 1784 5479
rect 1863 5479 1869 5480
rect 1863 5478 1864 5479
rect 1783 5476 1864 5478
rect 1783 5475 1784 5476
rect 1778 5474 1784 5475
rect 1863 5475 1864 5476
rect 1868 5475 1869 5479
rect 1974 5476 1975 5480
rect 1979 5476 1980 5480
rect 1974 5475 1980 5476
rect 2138 5479 2144 5480
rect 2138 5475 2139 5479
rect 2143 5475 2144 5479
rect 1863 5474 1869 5475
rect 2138 5474 2144 5475
rect 2354 5479 2360 5480
rect 2354 5475 2355 5479
rect 2359 5475 2360 5479
rect 2354 5474 2360 5475
rect 2562 5479 2568 5480
rect 2562 5475 2563 5479
rect 2567 5475 2568 5479
rect 2562 5474 2568 5475
rect 2754 5479 2760 5480
rect 2754 5475 2755 5479
rect 2759 5475 2760 5479
rect 2754 5474 2760 5475
rect 2938 5479 2944 5480
rect 2938 5475 2939 5479
rect 2943 5475 2944 5479
rect 2938 5474 2944 5475
rect 3114 5479 3120 5480
rect 3114 5475 3115 5479
rect 3119 5475 3120 5479
rect 3114 5474 3120 5475
rect 3290 5479 3296 5480
rect 3290 5475 3291 5479
rect 3295 5475 3296 5479
rect 3290 5474 3296 5475
rect 3466 5479 3472 5480
rect 3466 5475 3467 5479
rect 3471 5475 3472 5479
rect 3466 5474 3472 5475
rect 3642 5479 3648 5480
rect 3642 5475 3643 5479
rect 3647 5475 3648 5479
rect 3798 5476 3799 5480
rect 3803 5476 3804 5480
rect 4374 5479 4375 5483
rect 4380 5479 4381 5483
rect 4374 5478 4381 5479
rect 4383 5483 4389 5484
rect 4383 5479 4384 5483
rect 4388 5482 4389 5483
rect 4527 5483 4533 5484
rect 4527 5482 4528 5483
rect 4388 5480 4528 5482
rect 4388 5479 4389 5480
rect 4383 5478 4389 5479
rect 4527 5479 4528 5480
rect 4532 5479 4533 5483
rect 4527 5478 4533 5479
rect 4551 5483 4557 5484
rect 4551 5479 4552 5483
rect 4556 5482 4557 5483
rect 4679 5483 4685 5484
rect 4679 5482 4680 5483
rect 4556 5480 4680 5482
rect 4556 5479 4557 5480
rect 4551 5478 4557 5479
rect 4679 5479 4680 5480
rect 4684 5479 4685 5483
rect 4679 5478 4685 5479
rect 4762 5483 4768 5484
rect 4762 5479 4763 5483
rect 4767 5482 4768 5483
rect 4831 5483 4837 5484
rect 4831 5482 4832 5483
rect 4767 5480 4832 5482
rect 4767 5479 4768 5480
rect 4762 5478 4768 5479
rect 4831 5479 4832 5480
rect 4836 5479 4837 5483
rect 4831 5478 4837 5479
rect 4850 5483 4856 5484
rect 4850 5479 4851 5483
rect 4855 5482 4856 5483
rect 4983 5483 4989 5484
rect 4983 5482 4984 5483
rect 4855 5480 4984 5482
rect 4855 5479 4856 5480
rect 4850 5478 4856 5479
rect 4983 5479 4984 5480
rect 4988 5479 4989 5483
rect 4983 5478 4989 5479
rect 5015 5483 5021 5484
rect 5015 5479 5016 5483
rect 5020 5482 5021 5483
rect 5143 5483 5149 5484
rect 5143 5482 5144 5483
rect 5020 5480 5144 5482
rect 5020 5479 5021 5480
rect 5015 5478 5021 5479
rect 5143 5479 5144 5480
rect 5148 5479 5149 5483
rect 5143 5478 5149 5479
rect 3798 5475 3804 5476
rect 3838 5476 3844 5477
rect 5662 5476 5668 5477
rect 3642 5474 3648 5475
rect 3838 5472 3839 5476
rect 3843 5472 3844 5476
rect 3838 5471 3844 5472
rect 4250 5475 4256 5476
rect 4250 5471 4251 5475
rect 4255 5471 4256 5475
rect 4250 5470 4256 5471
rect 4402 5475 4408 5476
rect 4402 5471 4403 5475
rect 4407 5471 4408 5475
rect 4402 5470 4408 5471
rect 4554 5475 4560 5476
rect 4554 5471 4555 5475
rect 4559 5471 4560 5475
rect 4554 5470 4560 5471
rect 4706 5475 4712 5476
rect 4706 5471 4707 5475
rect 4711 5471 4712 5475
rect 4706 5470 4712 5471
rect 4858 5475 4864 5476
rect 4858 5471 4859 5475
rect 4863 5471 4864 5475
rect 4858 5470 4864 5471
rect 5018 5475 5024 5476
rect 5018 5471 5019 5475
rect 5023 5471 5024 5475
rect 5662 5472 5663 5476
rect 5667 5472 5668 5476
rect 5662 5471 5668 5472
rect 5018 5470 5024 5471
rect 511 5468 1101 5470
rect 511 5467 512 5468
rect 506 5466 512 5467
rect 2166 5464 2172 5465
rect 1974 5463 1980 5464
rect 1974 5459 1975 5463
rect 1979 5459 1980 5463
rect 2166 5460 2167 5464
rect 2171 5460 2172 5464
rect 2166 5459 2172 5460
rect 2382 5464 2388 5465
rect 2382 5460 2383 5464
rect 2387 5460 2388 5464
rect 2382 5459 2388 5460
rect 2590 5464 2596 5465
rect 2590 5460 2591 5464
rect 2595 5460 2596 5464
rect 2590 5459 2596 5460
rect 2782 5464 2788 5465
rect 2782 5460 2783 5464
rect 2787 5460 2788 5464
rect 2782 5459 2788 5460
rect 2966 5464 2972 5465
rect 2966 5460 2967 5464
rect 2971 5460 2972 5464
rect 2966 5459 2972 5460
rect 3142 5464 3148 5465
rect 3142 5460 3143 5464
rect 3147 5460 3148 5464
rect 3142 5459 3148 5460
rect 3318 5464 3324 5465
rect 3318 5460 3319 5464
rect 3323 5460 3324 5464
rect 3318 5459 3324 5460
rect 3494 5464 3500 5465
rect 3494 5460 3495 5464
rect 3499 5460 3500 5464
rect 3494 5459 3500 5460
rect 3670 5464 3676 5465
rect 3670 5460 3671 5464
rect 3675 5460 3676 5464
rect 3670 5459 3676 5460
rect 3798 5463 3804 5464
rect 3798 5459 3799 5463
rect 3803 5459 3804 5463
rect 4278 5460 4284 5461
rect 1974 5458 1980 5459
rect 3798 5458 3804 5459
rect 3838 5459 3844 5460
rect 3838 5455 3839 5459
rect 3843 5455 3844 5459
rect 4278 5456 4279 5460
rect 4283 5456 4284 5460
rect 4278 5455 4284 5456
rect 4430 5460 4436 5461
rect 4430 5456 4431 5460
rect 4435 5456 4436 5460
rect 4430 5455 4436 5456
rect 4582 5460 4588 5461
rect 4582 5456 4583 5460
rect 4587 5456 4588 5460
rect 4582 5455 4588 5456
rect 4734 5460 4740 5461
rect 4734 5456 4735 5460
rect 4739 5456 4740 5460
rect 4734 5455 4740 5456
rect 4886 5460 4892 5461
rect 4886 5456 4887 5460
rect 4891 5456 4892 5460
rect 4886 5455 4892 5456
rect 5046 5460 5052 5461
rect 5046 5456 5047 5460
rect 5051 5456 5052 5460
rect 5046 5455 5052 5456
rect 5662 5459 5668 5460
rect 5662 5455 5663 5459
rect 5667 5455 5668 5459
rect 3838 5454 3844 5455
rect 5662 5454 5668 5455
rect 378 5439 384 5440
rect 348 5430 350 5437
rect 378 5435 379 5439
rect 383 5438 384 5439
rect 618 5439 624 5440
rect 383 5436 497 5438
rect 383 5435 384 5436
rect 378 5434 384 5435
rect 618 5435 619 5439
rect 623 5438 624 5439
rect 866 5439 872 5440
rect 623 5436 745 5438
rect 623 5435 624 5436
rect 618 5434 624 5435
rect 866 5435 867 5439
rect 871 5438 872 5439
rect 1330 5439 1336 5440
rect 871 5436 993 5438
rect 871 5435 872 5436
rect 866 5434 872 5435
rect 1330 5435 1331 5439
rect 1335 5435 1336 5439
rect 1330 5434 1336 5435
rect 1362 5439 1368 5440
rect 1362 5435 1363 5439
rect 1367 5438 1368 5439
rect 1610 5439 1616 5440
rect 1367 5436 1489 5438
rect 1367 5435 1368 5436
rect 1362 5434 1368 5435
rect 1610 5435 1611 5439
rect 1615 5438 1616 5439
rect 1615 5436 1745 5438
rect 1615 5435 1616 5436
rect 1610 5434 1616 5435
rect 1278 5431 1284 5432
rect 1278 5430 1279 5431
rect 348 5428 1279 5430
rect 1278 5427 1279 5428
rect 1283 5427 1284 5431
rect 1278 5426 1284 5427
rect 506 5407 512 5408
rect 506 5403 507 5407
rect 511 5403 512 5407
rect 1487 5407 1493 5408
rect 1487 5406 1488 5407
rect 1357 5404 1488 5406
rect 506 5402 512 5403
rect 618 5403 624 5404
rect 618 5399 619 5403
rect 623 5399 624 5403
rect 618 5398 624 5399
rect 826 5403 832 5404
rect 826 5399 827 5403
rect 831 5399 832 5403
rect 826 5398 832 5399
rect 1042 5403 1048 5404
rect 1042 5399 1043 5403
rect 1047 5399 1048 5403
rect 1487 5403 1488 5404
rect 1492 5403 1493 5407
rect 1487 5402 1493 5403
rect 1586 5403 1592 5404
rect 1042 5398 1048 5399
rect 1586 5399 1587 5403
rect 1591 5399 1592 5403
rect 1586 5398 1592 5399
rect 1974 5397 1980 5398
rect 3798 5397 3804 5398
rect 1974 5393 1975 5397
rect 1979 5393 1980 5397
rect 1974 5392 1980 5393
rect 2310 5396 2316 5397
rect 2310 5392 2311 5396
rect 2315 5392 2316 5396
rect 2310 5391 2316 5392
rect 2510 5396 2516 5397
rect 2510 5392 2511 5396
rect 2515 5392 2516 5396
rect 2510 5391 2516 5392
rect 2702 5396 2708 5397
rect 2702 5392 2703 5396
rect 2707 5392 2708 5396
rect 2702 5391 2708 5392
rect 2886 5396 2892 5397
rect 2886 5392 2887 5396
rect 2891 5392 2892 5396
rect 2886 5391 2892 5392
rect 3070 5396 3076 5397
rect 3070 5392 3071 5396
rect 3075 5392 3076 5396
rect 3070 5391 3076 5392
rect 3246 5396 3252 5397
rect 3246 5392 3247 5396
rect 3251 5392 3252 5396
rect 3246 5391 3252 5392
rect 3422 5396 3428 5397
rect 3422 5392 3423 5396
rect 3427 5392 3428 5396
rect 3422 5391 3428 5392
rect 3606 5396 3612 5397
rect 3606 5392 3607 5396
rect 3611 5392 3612 5396
rect 3798 5393 3799 5397
rect 3803 5393 3804 5397
rect 3798 5392 3804 5393
rect 3606 5391 3612 5392
rect 2282 5381 2288 5382
rect 1974 5380 1980 5381
rect 1974 5376 1975 5380
rect 1979 5376 1980 5380
rect 2282 5377 2283 5381
rect 2287 5377 2288 5381
rect 2282 5376 2288 5377
rect 2482 5381 2488 5382
rect 2482 5377 2483 5381
rect 2487 5377 2488 5381
rect 2482 5376 2488 5377
rect 2674 5381 2680 5382
rect 2674 5377 2675 5381
rect 2679 5377 2680 5381
rect 2674 5376 2680 5377
rect 2858 5381 2864 5382
rect 2858 5377 2859 5381
rect 2863 5377 2864 5381
rect 2858 5376 2864 5377
rect 3042 5381 3048 5382
rect 3042 5377 3043 5381
rect 3047 5377 3048 5381
rect 3042 5376 3048 5377
rect 3218 5381 3224 5382
rect 3218 5377 3219 5381
rect 3223 5377 3224 5381
rect 3218 5376 3224 5377
rect 3394 5381 3400 5382
rect 3394 5377 3395 5381
rect 3399 5377 3400 5381
rect 3394 5376 3400 5377
rect 3578 5381 3584 5382
rect 3838 5381 3844 5382
rect 5662 5381 5668 5382
rect 3578 5377 3579 5381
rect 3583 5377 3584 5381
rect 3578 5376 3584 5377
rect 3798 5380 3804 5381
rect 3798 5376 3799 5380
rect 3803 5376 3804 5380
rect 3838 5377 3839 5381
rect 3843 5377 3844 5381
rect 3838 5376 3844 5377
rect 4278 5380 4284 5381
rect 4278 5376 4279 5380
rect 4283 5376 4284 5380
rect 1974 5375 1980 5376
rect 3798 5375 3804 5376
rect 4278 5375 4284 5376
rect 4486 5380 4492 5381
rect 4486 5376 4487 5380
rect 4491 5376 4492 5380
rect 4486 5375 4492 5376
rect 4694 5380 4700 5381
rect 4694 5376 4695 5380
rect 4699 5376 4700 5380
rect 4694 5375 4700 5376
rect 4910 5380 4916 5381
rect 4910 5376 4911 5380
rect 4915 5376 4916 5380
rect 4910 5375 4916 5376
rect 5126 5380 5132 5381
rect 5126 5376 5127 5380
rect 5131 5376 5132 5380
rect 5662 5377 5663 5381
rect 5667 5377 5668 5381
rect 5662 5376 5668 5377
rect 5126 5375 5132 5376
rect 658 5371 664 5372
rect 658 5367 659 5371
rect 663 5370 664 5371
rect 2407 5371 2413 5372
rect 663 5368 1101 5370
rect 663 5367 664 5368
rect 658 5366 664 5367
rect 535 5363 541 5364
rect 535 5359 536 5363
rect 540 5362 541 5363
rect 618 5363 624 5364
rect 618 5362 619 5363
rect 540 5360 619 5362
rect 540 5359 541 5360
rect 535 5358 541 5359
rect 618 5359 619 5360
rect 623 5359 624 5363
rect 618 5358 624 5359
rect 735 5363 741 5364
rect 735 5359 736 5363
rect 740 5362 741 5363
rect 826 5363 832 5364
rect 826 5362 827 5363
rect 740 5360 827 5362
rect 740 5359 741 5360
rect 735 5358 741 5359
rect 826 5359 827 5360
rect 831 5359 832 5363
rect 826 5358 832 5359
rect 943 5363 949 5364
rect 943 5359 944 5363
rect 948 5362 949 5363
rect 1042 5363 1048 5364
rect 1042 5362 1043 5363
rect 948 5360 1043 5362
rect 948 5359 949 5360
rect 943 5358 949 5359
rect 1042 5359 1043 5360
rect 1047 5359 1048 5363
rect 1099 5362 1101 5368
rect 2407 5367 2408 5371
rect 2412 5370 2413 5371
rect 2442 5371 2448 5372
rect 2442 5370 2443 5371
rect 2412 5368 2443 5370
rect 2412 5367 2413 5368
rect 2407 5366 2413 5367
rect 2442 5367 2443 5368
rect 2447 5367 2448 5371
rect 2442 5366 2448 5367
rect 2607 5371 2616 5372
rect 2607 5367 2608 5371
rect 2615 5367 2616 5371
rect 2607 5366 2616 5367
rect 2799 5371 2805 5372
rect 2799 5367 2800 5371
rect 2804 5370 2805 5371
rect 2810 5371 2816 5372
rect 2810 5370 2811 5371
rect 2804 5368 2811 5370
rect 2804 5367 2805 5368
rect 2799 5366 2805 5367
rect 2810 5367 2811 5368
rect 2815 5367 2816 5371
rect 2810 5366 2816 5367
rect 2983 5371 2992 5372
rect 2983 5367 2984 5371
rect 2991 5367 2992 5371
rect 2983 5366 2992 5367
rect 3166 5371 3173 5372
rect 3166 5367 3167 5371
rect 3172 5367 3173 5371
rect 3166 5366 3173 5367
rect 3343 5371 3352 5372
rect 3343 5367 3344 5371
rect 3351 5367 3352 5371
rect 3343 5366 3352 5367
rect 3519 5371 3528 5372
rect 3519 5367 3520 5371
rect 3527 5367 3528 5371
rect 3519 5366 3528 5367
rect 3674 5371 3680 5372
rect 3674 5367 3675 5371
rect 3679 5370 3680 5371
rect 3703 5371 3709 5372
rect 3703 5370 3704 5371
rect 3679 5368 3704 5370
rect 3679 5367 3680 5368
rect 3674 5366 3680 5367
rect 3703 5367 3704 5368
rect 3708 5367 3709 5371
rect 3703 5366 3709 5367
rect 4250 5365 4256 5366
rect 3838 5364 3844 5365
rect 1159 5363 1165 5364
rect 1159 5362 1160 5363
rect 1099 5360 1160 5362
rect 1042 5358 1048 5359
rect 1159 5359 1160 5360
rect 1164 5359 1165 5363
rect 1159 5358 1165 5359
rect 1330 5363 1336 5364
rect 1330 5359 1331 5363
rect 1335 5362 1336 5363
rect 1383 5363 1389 5364
rect 1383 5362 1384 5363
rect 1335 5360 1384 5362
rect 1335 5359 1336 5360
rect 1330 5358 1336 5359
rect 1383 5359 1384 5360
rect 1388 5359 1389 5363
rect 1383 5358 1389 5359
rect 1487 5363 1493 5364
rect 1487 5359 1488 5363
rect 1492 5362 1493 5363
rect 1615 5363 1621 5364
rect 1615 5362 1616 5363
rect 1492 5360 1616 5362
rect 1492 5359 1493 5360
rect 1487 5358 1493 5359
rect 1615 5359 1616 5360
rect 1620 5359 1621 5363
rect 3838 5360 3839 5364
rect 3843 5360 3844 5364
rect 4250 5361 4251 5365
rect 4255 5361 4256 5365
rect 4250 5360 4256 5361
rect 4458 5365 4464 5366
rect 4458 5361 4459 5365
rect 4463 5361 4464 5365
rect 4458 5360 4464 5361
rect 4666 5365 4672 5366
rect 4666 5361 4667 5365
rect 4671 5361 4672 5365
rect 4666 5360 4672 5361
rect 4882 5365 4888 5366
rect 4882 5361 4883 5365
rect 4887 5361 4888 5365
rect 4882 5360 4888 5361
rect 5098 5365 5104 5366
rect 5098 5361 5099 5365
rect 5103 5361 5104 5365
rect 5098 5360 5104 5361
rect 5662 5364 5668 5365
rect 5662 5360 5663 5364
rect 5667 5360 5668 5364
rect 3838 5359 3844 5360
rect 5662 5359 5668 5360
rect 1615 5358 1621 5359
rect 110 5356 116 5357
rect 1934 5356 1940 5357
rect 4583 5356 4589 5357
rect 110 5352 111 5356
rect 115 5352 116 5356
rect 110 5351 116 5352
rect 410 5355 416 5356
rect 410 5351 411 5355
rect 415 5351 416 5355
rect 410 5350 416 5351
rect 610 5355 616 5356
rect 610 5351 611 5355
rect 615 5351 616 5355
rect 610 5350 616 5351
rect 818 5355 824 5356
rect 818 5351 819 5355
rect 823 5351 824 5355
rect 818 5350 824 5351
rect 1034 5355 1040 5356
rect 1034 5351 1035 5355
rect 1039 5351 1040 5355
rect 1034 5350 1040 5351
rect 1258 5355 1264 5356
rect 1258 5351 1259 5355
rect 1263 5351 1264 5355
rect 1258 5350 1264 5351
rect 1490 5355 1496 5356
rect 1490 5351 1491 5355
rect 1495 5351 1496 5355
rect 1934 5352 1935 5356
rect 1939 5352 1940 5356
rect 1934 5351 1940 5352
rect 4375 5355 4381 5356
rect 4375 5351 4376 5355
rect 4380 5354 4381 5355
rect 4418 5355 4424 5356
rect 4418 5354 4419 5355
rect 4380 5352 4419 5354
rect 4380 5351 4381 5352
rect 1490 5350 1496 5351
rect 4375 5350 4381 5351
rect 4418 5351 4419 5352
rect 4423 5351 4424 5355
rect 4418 5350 4424 5351
rect 4574 5355 4580 5356
rect 4574 5351 4575 5355
rect 4579 5354 4580 5355
rect 4583 5354 4584 5356
rect 4579 5352 4584 5354
rect 4588 5352 4589 5356
rect 4579 5351 4580 5352
rect 4583 5351 4589 5352
rect 4791 5355 4797 5356
rect 4791 5351 4792 5355
rect 4796 5354 4797 5355
rect 4806 5355 4812 5356
rect 4806 5354 4807 5355
rect 4796 5352 4807 5354
rect 4796 5351 4797 5352
rect 4574 5350 4580 5351
rect 4791 5350 4797 5351
rect 4806 5351 4807 5352
rect 4811 5351 4812 5355
rect 4806 5350 4812 5351
rect 5007 5355 5016 5356
rect 5007 5351 5008 5355
rect 5015 5351 5016 5355
rect 5007 5350 5016 5351
rect 5222 5355 5229 5356
rect 5222 5351 5223 5355
rect 5228 5351 5229 5355
rect 5222 5350 5229 5351
rect 438 5340 444 5341
rect 110 5339 116 5340
rect 110 5335 111 5339
rect 115 5335 116 5339
rect 438 5336 439 5340
rect 443 5336 444 5340
rect 438 5335 444 5336
rect 638 5340 644 5341
rect 638 5336 639 5340
rect 643 5336 644 5340
rect 638 5335 644 5336
rect 846 5340 852 5341
rect 846 5336 847 5340
rect 851 5336 852 5340
rect 846 5335 852 5336
rect 1062 5340 1068 5341
rect 1062 5336 1063 5340
rect 1067 5336 1068 5340
rect 1062 5335 1068 5336
rect 1286 5340 1292 5341
rect 1286 5336 1287 5340
rect 1291 5336 1292 5340
rect 1286 5335 1292 5336
rect 1518 5340 1524 5341
rect 1518 5336 1519 5340
rect 1523 5336 1524 5340
rect 1518 5335 1524 5336
rect 1934 5339 1940 5340
rect 1934 5335 1935 5339
rect 1939 5335 1940 5339
rect 110 5334 116 5335
rect 1934 5334 1940 5335
rect 2262 5331 2268 5332
rect 2262 5327 2263 5331
rect 2267 5330 2268 5331
rect 2442 5331 2448 5332
rect 2267 5328 2289 5330
rect 2267 5327 2268 5328
rect 2262 5326 2268 5327
rect 2442 5327 2443 5331
rect 2447 5330 2448 5331
rect 2610 5331 2616 5332
rect 2447 5328 2489 5330
rect 2447 5327 2448 5328
rect 2442 5326 2448 5327
rect 2610 5327 2611 5331
rect 2615 5330 2616 5331
rect 2954 5331 2960 5332
rect 2615 5328 2681 5330
rect 2615 5327 2616 5328
rect 2610 5326 2616 5327
rect 2954 5327 2955 5331
rect 2959 5327 2960 5331
rect 2954 5326 2960 5327
rect 2986 5331 2992 5332
rect 2986 5327 2987 5331
rect 2991 5330 2992 5331
rect 3326 5331 3332 5332
rect 3326 5330 3327 5331
rect 2991 5328 3049 5330
rect 3317 5328 3327 5330
rect 2991 5327 2992 5328
rect 2986 5326 2992 5327
rect 3326 5327 3327 5328
rect 3331 5327 3332 5331
rect 3326 5326 3332 5327
rect 3346 5331 3352 5332
rect 3346 5327 3347 5331
rect 3351 5330 3352 5331
rect 3522 5331 3528 5332
rect 3351 5328 3401 5330
rect 3351 5327 3352 5328
rect 3346 5326 3352 5327
rect 3522 5327 3523 5331
rect 3527 5330 3528 5331
rect 3527 5328 3585 5330
rect 3527 5327 3528 5328
rect 3522 5326 3528 5327
rect 4346 5315 4352 5316
rect 4346 5311 4347 5315
rect 4351 5311 4352 5315
rect 4346 5310 4352 5311
rect 4418 5315 4424 5316
rect 4418 5311 4419 5315
rect 4423 5314 4424 5315
rect 4762 5315 4768 5316
rect 4423 5312 4465 5314
rect 4423 5311 4424 5312
rect 4418 5310 4424 5311
rect 4762 5311 4763 5315
rect 4767 5311 4768 5315
rect 4762 5310 4768 5311
rect 4806 5315 4812 5316
rect 4806 5311 4807 5315
rect 4811 5314 4812 5315
rect 5010 5315 5016 5316
rect 4811 5312 4889 5314
rect 4811 5311 4812 5312
rect 4806 5310 4812 5311
rect 5010 5311 5011 5315
rect 5015 5314 5016 5315
rect 5015 5312 5105 5314
rect 5015 5311 5016 5312
rect 5010 5310 5016 5311
rect 2330 5299 2336 5300
rect 2330 5298 2331 5299
rect 2293 5296 2331 5298
rect 2330 5295 2331 5296
rect 2335 5295 2336 5299
rect 2482 5299 2488 5300
rect 2482 5298 2483 5299
rect 2437 5296 2483 5298
rect 2330 5294 2336 5295
rect 2482 5295 2483 5296
rect 2487 5295 2488 5299
rect 2647 5299 2653 5300
rect 2647 5298 2648 5299
rect 2589 5296 2648 5298
rect 2482 5294 2488 5295
rect 2647 5295 2648 5296
rect 2652 5295 2653 5299
rect 2802 5299 2808 5300
rect 2802 5298 2803 5299
rect 2749 5296 2803 5298
rect 2647 5294 2653 5295
rect 2802 5295 2803 5296
rect 2807 5295 2808 5299
rect 2802 5294 2808 5295
rect 2810 5299 2816 5300
rect 2810 5295 2811 5299
rect 2815 5298 2816 5299
rect 3183 5299 3189 5300
rect 3183 5298 3184 5299
rect 2815 5296 2825 5298
rect 3101 5296 3184 5298
rect 2815 5295 2816 5296
rect 2810 5294 2816 5295
rect 3183 5295 3184 5296
rect 3188 5295 3189 5299
rect 3519 5299 3525 5300
rect 3519 5298 3520 5299
rect 3477 5296 3520 5298
rect 3183 5294 3189 5295
rect 3194 5295 3200 5296
rect 3194 5291 3195 5295
rect 3199 5291 3200 5295
rect 3519 5295 3520 5296
rect 3524 5295 3525 5299
rect 3519 5294 3525 5295
rect 3674 5299 3680 5300
rect 3674 5295 3675 5299
rect 3679 5295 3680 5299
rect 3674 5294 3680 5295
rect 3194 5290 3200 5291
rect 110 5281 116 5282
rect 1934 5281 1940 5282
rect 110 5277 111 5281
rect 115 5277 116 5281
rect 110 5276 116 5277
rect 590 5280 596 5281
rect 590 5276 591 5280
rect 595 5276 596 5280
rect 590 5275 596 5276
rect 726 5280 732 5281
rect 726 5276 727 5280
rect 731 5276 732 5280
rect 726 5275 732 5276
rect 862 5280 868 5281
rect 862 5276 863 5280
rect 867 5276 868 5280
rect 862 5275 868 5276
rect 998 5280 1004 5281
rect 998 5276 999 5280
rect 1003 5276 1004 5280
rect 998 5275 1004 5276
rect 1134 5280 1140 5281
rect 1134 5276 1135 5280
rect 1139 5276 1140 5280
rect 1134 5275 1140 5276
rect 1270 5280 1276 5281
rect 1270 5276 1271 5280
rect 1275 5276 1276 5280
rect 1270 5275 1276 5276
rect 1406 5280 1412 5281
rect 1406 5276 1407 5280
rect 1411 5276 1412 5280
rect 1406 5275 1412 5276
rect 1542 5280 1548 5281
rect 1542 5276 1543 5280
rect 1547 5276 1548 5280
rect 1934 5277 1935 5281
rect 1939 5277 1940 5281
rect 1934 5276 1940 5277
rect 1542 5275 1548 5276
rect 4479 5267 4485 5268
rect 4479 5266 4480 5267
rect 562 5265 568 5266
rect 110 5264 116 5265
rect 110 5260 111 5264
rect 115 5260 116 5264
rect 562 5261 563 5265
rect 567 5261 568 5265
rect 562 5260 568 5261
rect 698 5265 704 5266
rect 698 5261 699 5265
rect 703 5261 704 5265
rect 698 5260 704 5261
rect 834 5265 840 5266
rect 834 5261 835 5265
rect 839 5261 840 5265
rect 834 5260 840 5261
rect 970 5265 976 5266
rect 970 5261 971 5265
rect 975 5261 976 5265
rect 970 5260 976 5261
rect 1106 5265 1112 5266
rect 1106 5261 1107 5265
rect 1111 5261 1112 5265
rect 1106 5260 1112 5261
rect 1242 5265 1248 5266
rect 1242 5261 1243 5265
rect 1247 5261 1248 5265
rect 1242 5260 1248 5261
rect 1378 5265 1384 5266
rect 1378 5261 1379 5265
rect 1383 5261 1384 5265
rect 1378 5260 1384 5261
rect 1514 5265 1520 5266
rect 1514 5261 1515 5265
rect 1519 5261 1520 5265
rect 1514 5260 1520 5261
rect 1934 5264 1940 5265
rect 4349 5264 4480 5266
rect 1934 5260 1935 5264
rect 1939 5260 1940 5264
rect 4479 5263 4480 5264
rect 4484 5263 4485 5267
rect 4479 5262 4485 5263
rect 4502 5267 4508 5268
rect 4502 5263 4503 5267
rect 4507 5263 4508 5267
rect 4943 5267 4949 5268
rect 4943 5266 4944 5267
rect 4813 5264 4944 5266
rect 4502 5262 4508 5263
rect 4943 5263 4944 5264
rect 4948 5263 4949 5267
rect 5127 5267 5133 5268
rect 5127 5266 5128 5267
rect 5045 5264 5128 5266
rect 4943 5262 4949 5263
rect 5127 5263 5128 5264
rect 5132 5263 5133 5267
rect 5127 5262 5133 5263
rect 5222 5267 5228 5268
rect 5222 5263 5223 5267
rect 5227 5263 5228 5267
rect 5222 5262 5228 5263
rect 110 5259 116 5260
rect 1934 5259 1940 5260
rect 687 5255 696 5256
rect 687 5251 688 5255
rect 695 5251 696 5255
rect 687 5250 696 5251
rect 823 5255 832 5256
rect 823 5251 824 5255
rect 831 5251 832 5255
rect 823 5250 832 5251
rect 959 5255 968 5256
rect 959 5251 960 5255
rect 967 5251 968 5255
rect 959 5250 968 5251
rect 1095 5255 1101 5256
rect 1095 5251 1096 5255
rect 1100 5254 1101 5255
rect 1103 5255 1109 5256
rect 1103 5254 1104 5255
rect 1100 5252 1104 5254
rect 1100 5251 1101 5252
rect 1095 5250 1101 5251
rect 1103 5251 1104 5252
rect 1108 5251 1109 5255
rect 1103 5250 1109 5251
rect 1231 5255 1240 5256
rect 1231 5251 1232 5255
rect 1239 5251 1240 5255
rect 1231 5250 1240 5251
rect 1367 5255 1376 5256
rect 1367 5251 1368 5255
rect 1375 5251 1376 5255
rect 1367 5250 1376 5251
rect 1503 5255 1512 5256
rect 1503 5251 1504 5255
rect 1511 5251 1512 5255
rect 1503 5250 1512 5251
rect 1586 5255 1592 5256
rect 1586 5251 1587 5255
rect 1591 5254 1592 5255
rect 1639 5255 1645 5256
rect 1639 5254 1640 5255
rect 1591 5252 1640 5254
rect 1591 5251 1592 5252
rect 1586 5250 1592 5251
rect 1639 5251 1640 5252
rect 1644 5251 1645 5255
rect 1639 5250 1645 5251
rect 2318 5255 2325 5256
rect 2318 5251 2319 5255
rect 2324 5251 2325 5255
rect 2318 5250 2325 5251
rect 2330 5255 2336 5256
rect 2330 5251 2331 5255
rect 2335 5254 2336 5255
rect 2463 5255 2469 5256
rect 2463 5254 2464 5255
rect 2335 5252 2464 5254
rect 2335 5251 2336 5252
rect 2330 5250 2336 5251
rect 2463 5251 2464 5252
rect 2468 5251 2469 5255
rect 2463 5250 2469 5251
rect 2482 5255 2488 5256
rect 2482 5251 2483 5255
rect 2487 5254 2488 5255
rect 2615 5255 2621 5256
rect 2615 5254 2616 5255
rect 2487 5252 2616 5254
rect 2487 5251 2488 5252
rect 2482 5250 2488 5251
rect 2615 5251 2616 5252
rect 2620 5251 2621 5255
rect 2615 5250 2621 5251
rect 2647 5255 2653 5256
rect 2647 5251 2648 5255
rect 2652 5254 2653 5255
rect 2775 5255 2781 5256
rect 2775 5254 2776 5255
rect 2652 5252 2776 5254
rect 2652 5251 2653 5252
rect 2647 5250 2653 5251
rect 2775 5251 2776 5252
rect 2780 5251 2781 5255
rect 2775 5250 2781 5251
rect 2802 5255 2808 5256
rect 2802 5251 2803 5255
rect 2807 5254 2808 5255
rect 2943 5255 2949 5256
rect 2943 5254 2944 5255
rect 2807 5252 2944 5254
rect 2807 5251 2808 5252
rect 2802 5250 2808 5251
rect 2943 5251 2944 5252
rect 2948 5251 2949 5255
rect 2943 5250 2949 5251
rect 2954 5255 2960 5256
rect 2954 5251 2955 5255
rect 2959 5254 2960 5255
rect 3127 5255 3133 5256
rect 3127 5254 3128 5255
rect 2959 5252 3128 5254
rect 2959 5251 2960 5252
rect 2954 5250 2960 5251
rect 3127 5251 3128 5252
rect 3132 5251 3133 5255
rect 3127 5250 3133 5251
rect 3183 5255 3189 5256
rect 3183 5251 3184 5255
rect 3188 5254 3189 5255
rect 3311 5255 3317 5256
rect 3311 5254 3312 5255
rect 3188 5252 3312 5254
rect 3188 5251 3189 5252
rect 3183 5250 3189 5251
rect 3311 5251 3312 5252
rect 3316 5251 3317 5255
rect 3311 5250 3317 5251
rect 3354 5255 3360 5256
rect 3354 5251 3355 5255
rect 3359 5254 3360 5255
rect 3503 5255 3509 5256
rect 3503 5254 3504 5255
rect 3359 5252 3504 5254
rect 3359 5251 3360 5252
rect 3354 5250 3360 5251
rect 3503 5251 3504 5252
rect 3508 5251 3509 5255
rect 3503 5250 3509 5251
rect 3519 5255 3525 5256
rect 3519 5251 3520 5255
rect 3524 5254 3525 5255
rect 3703 5255 3709 5256
rect 3703 5254 3704 5255
rect 3524 5252 3704 5254
rect 3524 5251 3525 5252
rect 3519 5250 3525 5251
rect 3703 5251 3704 5252
rect 3708 5251 3709 5255
rect 3703 5250 3709 5251
rect 1974 5248 1980 5249
rect 3798 5248 3804 5249
rect 1974 5244 1975 5248
rect 1979 5244 1980 5248
rect 1974 5243 1980 5244
rect 2194 5247 2200 5248
rect 2194 5243 2195 5247
rect 2199 5243 2200 5247
rect 2194 5242 2200 5243
rect 2338 5247 2344 5248
rect 2338 5243 2339 5247
rect 2343 5243 2344 5247
rect 2338 5242 2344 5243
rect 2490 5247 2496 5248
rect 2490 5243 2491 5247
rect 2495 5243 2496 5247
rect 2490 5242 2496 5243
rect 2650 5247 2656 5248
rect 2650 5243 2651 5247
rect 2655 5243 2656 5247
rect 2650 5242 2656 5243
rect 2818 5247 2824 5248
rect 2818 5243 2819 5247
rect 2823 5243 2824 5247
rect 2818 5242 2824 5243
rect 3002 5247 3008 5248
rect 3002 5243 3003 5247
rect 3007 5243 3008 5247
rect 3002 5242 3008 5243
rect 3186 5247 3192 5248
rect 3186 5243 3187 5247
rect 3191 5243 3192 5247
rect 3186 5242 3192 5243
rect 3378 5247 3384 5248
rect 3378 5243 3379 5247
rect 3383 5243 3384 5247
rect 3378 5242 3384 5243
rect 3578 5247 3584 5248
rect 3578 5243 3579 5247
rect 3583 5243 3584 5247
rect 3798 5244 3799 5248
rect 3803 5244 3804 5248
rect 3798 5243 3804 5244
rect 3578 5242 3584 5243
rect 2222 5232 2228 5233
rect 1974 5231 1980 5232
rect 1974 5227 1975 5231
rect 1979 5227 1980 5231
rect 2222 5228 2223 5232
rect 2227 5228 2228 5232
rect 2222 5227 2228 5228
rect 2366 5232 2372 5233
rect 2366 5228 2367 5232
rect 2371 5228 2372 5232
rect 2366 5227 2372 5228
rect 2518 5232 2524 5233
rect 2518 5228 2519 5232
rect 2523 5228 2524 5232
rect 2518 5227 2524 5228
rect 2678 5232 2684 5233
rect 2678 5228 2679 5232
rect 2683 5228 2684 5232
rect 2678 5227 2684 5228
rect 2846 5232 2852 5233
rect 2846 5228 2847 5232
rect 2851 5228 2852 5232
rect 2846 5227 2852 5228
rect 3030 5232 3036 5233
rect 3030 5228 3031 5232
rect 3035 5228 3036 5232
rect 3030 5227 3036 5228
rect 3214 5232 3220 5233
rect 3214 5228 3215 5232
rect 3219 5228 3220 5232
rect 3214 5227 3220 5228
rect 3406 5232 3412 5233
rect 3406 5228 3407 5232
rect 3411 5228 3412 5232
rect 3406 5227 3412 5228
rect 3606 5232 3612 5233
rect 3606 5228 3607 5232
rect 3611 5228 3612 5232
rect 3606 5227 3612 5228
rect 3798 5231 3804 5232
rect 3798 5227 3799 5231
rect 3803 5227 3804 5231
rect 1974 5226 1980 5227
rect 3798 5226 3804 5227
rect 4346 5223 4352 5224
rect 4346 5219 4347 5223
rect 4351 5222 4352 5223
rect 4375 5223 4381 5224
rect 4375 5222 4376 5223
rect 4351 5220 4376 5222
rect 4351 5219 4352 5220
rect 4346 5218 4352 5219
rect 4375 5219 4376 5220
rect 4380 5219 4381 5223
rect 4375 5218 4381 5219
rect 4479 5223 4485 5224
rect 4479 5219 4480 5223
rect 4484 5222 4485 5223
rect 4607 5223 4613 5224
rect 4607 5222 4608 5223
rect 4484 5220 4608 5222
rect 4484 5219 4485 5220
rect 4479 5218 4485 5219
rect 4607 5219 4608 5220
rect 4612 5219 4613 5223
rect 4607 5218 4613 5219
rect 4839 5223 4848 5224
rect 4839 5219 4840 5223
rect 4847 5219 4848 5223
rect 4839 5218 4848 5219
rect 4943 5223 4949 5224
rect 4943 5219 4944 5223
rect 4948 5222 4949 5223
rect 5071 5223 5077 5224
rect 5071 5222 5072 5223
rect 4948 5220 5072 5222
rect 4948 5219 4949 5220
rect 4943 5218 4949 5219
rect 5071 5219 5072 5220
rect 5076 5219 5077 5223
rect 5071 5218 5077 5219
rect 5127 5223 5133 5224
rect 5127 5219 5128 5223
rect 5132 5222 5133 5223
rect 5311 5223 5317 5224
rect 5311 5222 5312 5223
rect 5132 5220 5312 5222
rect 5132 5219 5133 5220
rect 5127 5218 5133 5219
rect 5311 5219 5312 5220
rect 5316 5219 5317 5223
rect 5311 5218 5317 5219
rect 3838 5216 3844 5217
rect 5662 5216 5668 5217
rect 658 5215 664 5216
rect 658 5211 659 5215
rect 663 5211 664 5215
rect 658 5210 664 5211
rect 690 5215 696 5216
rect 690 5211 691 5215
rect 695 5214 696 5215
rect 826 5215 832 5216
rect 695 5212 705 5214
rect 695 5211 696 5212
rect 690 5210 696 5211
rect 826 5211 827 5215
rect 831 5214 832 5215
rect 962 5215 968 5216
rect 831 5212 841 5214
rect 831 5211 832 5212
rect 826 5210 832 5211
rect 962 5211 963 5215
rect 967 5214 968 5215
rect 1103 5215 1109 5216
rect 967 5212 977 5214
rect 967 5211 968 5212
rect 962 5210 968 5211
rect 1103 5211 1104 5215
rect 1108 5214 1109 5215
rect 1234 5215 1240 5216
rect 1108 5212 1113 5214
rect 1108 5211 1109 5212
rect 1103 5210 1109 5211
rect 1234 5211 1235 5215
rect 1239 5214 1240 5215
rect 1370 5215 1376 5216
rect 1239 5212 1249 5214
rect 1239 5211 1240 5212
rect 1234 5210 1240 5211
rect 1370 5211 1371 5215
rect 1375 5214 1376 5215
rect 1506 5215 1512 5216
rect 1375 5212 1385 5214
rect 1375 5211 1376 5212
rect 1370 5210 1376 5211
rect 1506 5211 1507 5215
rect 1511 5214 1512 5215
rect 1511 5212 1521 5214
rect 3838 5212 3839 5216
rect 3843 5212 3844 5216
rect 1511 5211 1512 5212
rect 3838 5211 3844 5212
rect 4250 5215 4256 5216
rect 4250 5211 4251 5215
rect 4255 5211 4256 5215
rect 1506 5210 1512 5211
rect 4250 5210 4256 5211
rect 4482 5215 4488 5216
rect 4482 5211 4483 5215
rect 4487 5211 4488 5215
rect 4482 5210 4488 5211
rect 4714 5215 4720 5216
rect 4714 5211 4715 5215
rect 4719 5211 4720 5215
rect 4714 5210 4720 5211
rect 4946 5215 4952 5216
rect 4946 5211 4947 5215
rect 4951 5211 4952 5215
rect 4946 5210 4952 5211
rect 5186 5215 5192 5216
rect 5186 5211 5187 5215
rect 5191 5211 5192 5215
rect 5662 5212 5663 5216
rect 5667 5212 5668 5216
rect 5662 5211 5668 5212
rect 5186 5210 5192 5211
rect 4278 5200 4284 5201
rect 3838 5199 3844 5200
rect 3838 5195 3839 5199
rect 3843 5195 3844 5199
rect 4278 5196 4279 5200
rect 4283 5196 4284 5200
rect 4278 5195 4284 5196
rect 4510 5200 4516 5201
rect 4510 5196 4511 5200
rect 4515 5196 4516 5200
rect 4510 5195 4516 5196
rect 4742 5200 4748 5201
rect 4742 5196 4743 5200
rect 4747 5196 4748 5200
rect 4742 5195 4748 5196
rect 4974 5200 4980 5201
rect 4974 5196 4975 5200
rect 4979 5196 4980 5200
rect 4974 5195 4980 5196
rect 5214 5200 5220 5201
rect 5214 5196 5215 5200
rect 5219 5196 5220 5200
rect 5214 5195 5220 5196
rect 5662 5199 5668 5200
rect 5662 5195 5663 5199
rect 5667 5195 5668 5199
rect 3838 5194 3844 5195
rect 5662 5194 5668 5195
rect 1974 5173 1980 5174
rect 3798 5173 3804 5174
rect 1974 5169 1975 5173
rect 1979 5169 1980 5173
rect 1974 5168 1980 5169
rect 2022 5172 2028 5173
rect 2022 5168 2023 5172
rect 2027 5168 2028 5172
rect 2022 5167 2028 5168
rect 2158 5172 2164 5173
rect 2158 5168 2159 5172
rect 2163 5168 2164 5172
rect 2158 5167 2164 5168
rect 2326 5172 2332 5173
rect 2326 5168 2327 5172
rect 2331 5168 2332 5172
rect 2326 5167 2332 5168
rect 2510 5172 2516 5173
rect 2510 5168 2511 5172
rect 2515 5168 2516 5172
rect 2510 5167 2516 5168
rect 2694 5172 2700 5173
rect 2694 5168 2695 5172
rect 2699 5168 2700 5172
rect 2694 5167 2700 5168
rect 2886 5172 2892 5173
rect 2886 5168 2887 5172
rect 2891 5168 2892 5172
rect 2886 5167 2892 5168
rect 3086 5172 3092 5173
rect 3086 5168 3087 5172
rect 3091 5168 3092 5172
rect 3086 5167 3092 5168
rect 3286 5172 3292 5173
rect 3286 5168 3287 5172
rect 3291 5168 3292 5172
rect 3286 5167 3292 5168
rect 3494 5172 3500 5173
rect 3494 5168 3495 5172
rect 3499 5168 3500 5172
rect 3494 5167 3500 5168
rect 3678 5172 3684 5173
rect 3678 5168 3679 5172
rect 3683 5168 3684 5172
rect 3798 5169 3799 5173
rect 3803 5169 3804 5173
rect 3798 5168 3804 5169
rect 3678 5167 3684 5168
rect 1994 5157 2000 5158
rect 1974 5156 1980 5157
rect 1974 5152 1975 5156
rect 1979 5152 1980 5156
rect 1994 5153 1995 5157
rect 1999 5153 2000 5157
rect 1994 5152 2000 5153
rect 2130 5157 2136 5158
rect 2130 5153 2131 5157
rect 2135 5153 2136 5157
rect 2130 5152 2136 5153
rect 2298 5157 2304 5158
rect 2298 5153 2299 5157
rect 2303 5153 2304 5157
rect 2298 5152 2304 5153
rect 2482 5157 2488 5158
rect 2482 5153 2483 5157
rect 2487 5153 2488 5157
rect 2482 5152 2488 5153
rect 2666 5157 2672 5158
rect 2666 5153 2667 5157
rect 2671 5153 2672 5157
rect 2666 5152 2672 5153
rect 2858 5157 2864 5158
rect 2858 5153 2859 5157
rect 2863 5153 2864 5157
rect 2858 5152 2864 5153
rect 3058 5157 3064 5158
rect 3058 5153 3059 5157
rect 3063 5153 3064 5157
rect 3058 5152 3064 5153
rect 3258 5157 3264 5158
rect 3258 5153 3259 5157
rect 3263 5153 3264 5157
rect 3258 5152 3264 5153
rect 3466 5157 3472 5158
rect 3466 5153 3467 5157
rect 3471 5153 3472 5157
rect 3466 5152 3472 5153
rect 3650 5157 3656 5158
rect 3650 5153 3651 5157
rect 3655 5153 3656 5157
rect 3650 5152 3656 5153
rect 3798 5156 3804 5157
rect 3798 5152 3799 5156
rect 3803 5152 3804 5156
rect 1974 5151 1980 5152
rect 3798 5151 3804 5152
rect 2090 5147 2096 5148
rect 2090 5143 2091 5147
rect 2095 5146 2096 5147
rect 2119 5147 2125 5148
rect 2119 5146 2120 5147
rect 2095 5144 2120 5146
rect 2095 5143 2096 5144
rect 2090 5142 2096 5143
rect 2119 5143 2120 5144
rect 2124 5143 2125 5147
rect 2119 5142 2125 5143
rect 2138 5147 2144 5148
rect 2138 5143 2139 5147
rect 2143 5146 2144 5147
rect 2255 5147 2261 5148
rect 2255 5146 2256 5147
rect 2143 5144 2256 5146
rect 2143 5143 2144 5144
rect 2138 5142 2144 5143
rect 2255 5143 2256 5144
rect 2260 5143 2261 5147
rect 2255 5142 2261 5143
rect 2423 5147 2432 5148
rect 2423 5143 2424 5147
rect 2431 5143 2432 5147
rect 2423 5142 2432 5143
rect 2607 5147 2616 5148
rect 2607 5143 2608 5147
rect 2615 5143 2616 5147
rect 2791 5147 2797 5148
rect 2791 5146 2792 5147
rect 2607 5142 2616 5143
rect 2779 5144 2792 5146
rect 2226 5139 2232 5140
rect 2226 5135 2227 5139
rect 2231 5138 2232 5139
rect 2779 5138 2781 5144
rect 2791 5143 2792 5144
rect 2796 5143 2797 5147
rect 2791 5142 2797 5143
rect 2983 5147 2989 5148
rect 2983 5143 2984 5147
rect 2988 5146 2989 5147
rect 2998 5147 3004 5148
rect 2998 5146 2999 5147
rect 2988 5144 2999 5146
rect 2988 5143 2989 5144
rect 2983 5142 2989 5143
rect 2998 5143 2999 5144
rect 3003 5143 3004 5147
rect 2998 5142 3004 5143
rect 3183 5147 3189 5148
rect 3183 5143 3184 5147
rect 3188 5146 3189 5147
rect 3194 5147 3200 5148
rect 3194 5146 3195 5147
rect 3188 5144 3195 5146
rect 3188 5143 3189 5144
rect 3183 5142 3189 5143
rect 3194 5143 3195 5144
rect 3199 5143 3200 5147
rect 3194 5142 3200 5143
rect 3383 5147 3389 5148
rect 3383 5143 3384 5147
rect 3388 5146 3389 5147
rect 3426 5147 3432 5148
rect 3426 5146 3427 5147
rect 3388 5144 3427 5146
rect 3388 5143 3389 5144
rect 3383 5142 3389 5143
rect 3426 5143 3427 5144
rect 3431 5143 3432 5147
rect 3426 5142 3432 5143
rect 3591 5147 3597 5148
rect 3591 5143 3592 5147
rect 3596 5146 3597 5147
rect 3606 5147 3612 5148
rect 3606 5146 3607 5147
rect 3596 5144 3607 5146
rect 3596 5143 3597 5144
rect 3591 5142 3597 5143
rect 3606 5143 3607 5144
rect 3611 5143 3612 5147
rect 3606 5142 3612 5143
rect 3746 5147 3752 5148
rect 3746 5143 3747 5147
rect 3751 5146 3752 5147
rect 3775 5147 3781 5148
rect 3775 5146 3776 5147
rect 3751 5144 3776 5146
rect 3751 5143 3752 5144
rect 3746 5142 3752 5143
rect 3775 5143 3776 5144
rect 3780 5143 3781 5147
rect 3775 5142 3781 5143
rect 2231 5136 2781 5138
rect 2231 5135 2232 5136
rect 2226 5134 2232 5135
rect 2138 5115 2144 5116
rect 2138 5114 2139 5115
rect 2092 5112 2139 5114
rect 2092 5105 2094 5112
rect 2138 5111 2139 5112
rect 2143 5111 2144 5115
rect 2138 5110 2144 5111
rect 3838 5113 3844 5114
rect 5662 5113 5668 5114
rect 3838 5109 3839 5113
rect 3843 5109 3844 5113
rect 3838 5108 3844 5109
rect 3886 5112 3892 5113
rect 3886 5108 3887 5112
rect 3891 5108 3892 5112
rect 2226 5107 2232 5108
rect 2226 5103 2227 5107
rect 2231 5103 2232 5107
rect 2226 5102 2232 5103
rect 2318 5107 2324 5108
rect 2318 5103 2319 5107
rect 2323 5103 2324 5107
rect 2318 5102 2324 5103
rect 2426 5107 2432 5108
rect 2426 5103 2427 5107
rect 2431 5106 2432 5107
rect 2610 5107 2616 5108
rect 2431 5104 2489 5106
rect 2431 5103 2432 5104
rect 2426 5102 2432 5103
rect 2610 5103 2611 5107
rect 2615 5106 2616 5107
rect 2767 5107 2773 5108
rect 2615 5104 2673 5106
rect 2615 5103 2616 5104
rect 2610 5102 2616 5103
rect 2767 5103 2768 5107
rect 2772 5106 2773 5107
rect 2998 5107 3004 5108
rect 2772 5104 2865 5106
rect 2772 5103 2773 5104
rect 2767 5102 2773 5103
rect 2998 5103 2999 5107
rect 3003 5106 3004 5107
rect 3354 5107 3360 5108
rect 3003 5104 3065 5106
rect 3003 5103 3004 5104
rect 2998 5102 3004 5103
rect 3354 5103 3355 5107
rect 3359 5103 3360 5107
rect 3354 5102 3360 5103
rect 3426 5107 3432 5108
rect 3426 5103 3427 5107
rect 3431 5106 3432 5107
rect 3606 5107 3612 5108
rect 3886 5107 3892 5108
rect 4134 5112 4140 5113
rect 4134 5108 4135 5112
rect 4139 5108 4140 5112
rect 4134 5107 4140 5108
rect 4406 5112 4412 5113
rect 4406 5108 4407 5112
rect 4411 5108 4412 5112
rect 4406 5107 4412 5108
rect 4678 5112 4684 5113
rect 4678 5108 4679 5112
rect 4683 5108 4684 5112
rect 4678 5107 4684 5108
rect 4958 5112 4964 5113
rect 4958 5108 4959 5112
rect 4963 5108 4964 5112
rect 4958 5107 4964 5108
rect 5238 5112 5244 5113
rect 5238 5108 5239 5112
rect 5243 5108 5244 5112
rect 5662 5109 5663 5113
rect 5667 5109 5668 5113
rect 5662 5108 5668 5109
rect 5238 5107 5244 5108
rect 3431 5104 3473 5106
rect 3431 5103 3432 5104
rect 3426 5102 3432 5103
rect 3606 5103 3607 5107
rect 3611 5106 3612 5107
rect 3611 5104 3657 5106
rect 3611 5103 3612 5104
rect 3606 5102 3612 5103
rect 3858 5097 3864 5098
rect 3838 5096 3844 5097
rect 3838 5092 3839 5096
rect 3843 5092 3844 5096
rect 3858 5093 3859 5097
rect 3863 5093 3864 5097
rect 3858 5092 3864 5093
rect 4106 5097 4112 5098
rect 4106 5093 4107 5097
rect 4111 5093 4112 5097
rect 4106 5092 4112 5093
rect 4378 5097 4384 5098
rect 4378 5093 4379 5097
rect 4383 5093 4384 5097
rect 4378 5092 4384 5093
rect 4650 5097 4656 5098
rect 4650 5093 4651 5097
rect 4655 5093 4656 5097
rect 4650 5092 4656 5093
rect 4930 5097 4936 5098
rect 4930 5093 4931 5097
rect 4935 5093 4936 5097
rect 4930 5092 4936 5093
rect 5210 5097 5216 5098
rect 5210 5093 5211 5097
rect 5215 5093 5216 5097
rect 5210 5092 5216 5093
rect 5662 5096 5668 5097
rect 5662 5092 5663 5096
rect 5667 5092 5668 5096
rect 3838 5091 3844 5092
rect 5662 5091 5668 5092
rect 3954 5087 3960 5088
rect 3954 5083 3955 5087
rect 3959 5086 3960 5087
rect 3983 5087 3989 5088
rect 3983 5086 3984 5087
rect 3959 5084 3984 5086
rect 3959 5083 3960 5084
rect 3954 5082 3960 5083
rect 3983 5083 3984 5084
rect 3988 5083 3989 5087
rect 3983 5082 3989 5083
rect 4231 5087 4240 5088
rect 4231 5083 4232 5087
rect 4239 5083 4240 5087
rect 4231 5082 4240 5083
rect 4502 5087 4509 5088
rect 4502 5083 4503 5087
rect 4508 5083 4509 5087
rect 4775 5087 4781 5088
rect 4775 5086 4776 5087
rect 4502 5082 4509 5083
rect 4616 5084 4776 5086
rect 751 5079 757 5080
rect 751 5078 752 5079
rect 717 5076 752 5078
rect 442 5075 448 5076
rect 442 5071 443 5075
rect 447 5071 448 5075
rect 442 5070 448 5071
rect 490 5075 496 5076
rect 490 5071 491 5075
rect 495 5071 496 5075
rect 751 5075 752 5076
rect 756 5075 757 5079
rect 887 5079 893 5080
rect 887 5078 888 5079
rect 853 5076 888 5078
rect 751 5074 757 5075
rect 887 5075 888 5076
rect 892 5075 893 5079
rect 1023 5079 1029 5080
rect 1023 5078 1024 5079
rect 989 5076 1024 5078
rect 887 5074 893 5075
rect 1023 5075 1024 5076
rect 1028 5075 1029 5079
rect 1222 5079 1228 5080
rect 1023 5074 1029 5075
rect 1130 5075 1136 5076
rect 490 5070 496 5071
rect 1130 5071 1131 5075
rect 1135 5071 1136 5075
rect 1222 5075 1223 5079
rect 1227 5075 1228 5079
rect 2118 5079 2124 5080
rect 2118 5078 2119 5079
rect 1885 5076 2119 5078
rect 1222 5074 1228 5075
rect 1346 5075 1352 5076
rect 1130 5070 1136 5071
rect 1346 5071 1347 5075
rect 1351 5071 1352 5075
rect 1346 5070 1352 5071
rect 1586 5075 1592 5076
rect 1586 5071 1587 5075
rect 1591 5071 1592 5075
rect 1586 5070 1592 5071
rect 1658 5075 1664 5076
rect 1658 5071 1659 5075
rect 1663 5071 1664 5075
rect 2118 5075 2119 5076
rect 2123 5075 2124 5079
rect 4202 5079 4208 5080
rect 2118 5074 2124 5075
rect 2954 5075 2960 5076
rect 2954 5074 2955 5075
rect 2629 5072 2955 5074
rect 1658 5070 1664 5071
rect 2090 5071 2096 5072
rect 2090 5067 2091 5071
rect 2095 5067 2096 5071
rect 2954 5071 2955 5072
rect 2959 5071 2960 5075
rect 2954 5070 2960 5071
rect 3018 5075 3024 5076
rect 3018 5071 3019 5075
rect 3023 5074 3024 5075
rect 3746 5075 3752 5076
rect 3023 5072 3105 5074
rect 3023 5071 3024 5072
rect 3018 5070 3024 5071
rect 3746 5071 3747 5075
rect 3751 5071 3752 5075
rect 4202 5075 4203 5079
rect 4207 5078 4208 5079
rect 4616 5078 4618 5084
rect 4775 5083 4776 5084
rect 4780 5083 4781 5087
rect 4775 5082 4781 5083
rect 5055 5087 5064 5088
rect 5055 5083 5056 5087
rect 5063 5083 5064 5087
rect 5055 5082 5064 5083
rect 5334 5087 5341 5088
rect 5334 5083 5335 5087
rect 5340 5083 5341 5087
rect 5334 5082 5341 5083
rect 4207 5076 4618 5078
rect 4207 5075 4208 5076
rect 4202 5074 4208 5075
rect 3746 5070 3752 5071
rect 2090 5066 2096 5067
rect 1130 5055 1136 5056
rect 1130 5051 1131 5055
rect 1135 5054 1136 5055
rect 1423 5055 1429 5056
rect 1423 5054 1424 5055
rect 1135 5052 1424 5054
rect 1135 5051 1136 5052
rect 1130 5050 1136 5051
rect 1423 5051 1424 5052
rect 1428 5051 1429 5055
rect 1423 5050 1429 5051
rect 1586 5055 1592 5056
rect 1586 5051 1587 5055
rect 1591 5054 1592 5055
rect 1910 5055 1916 5056
rect 1910 5054 1911 5055
rect 1591 5052 1911 5054
rect 1591 5051 1592 5052
rect 1586 5050 1592 5051
rect 1910 5051 1911 5052
rect 1915 5051 1916 5055
rect 1910 5050 1916 5051
rect 4202 5047 4208 5048
rect 442 5043 448 5044
rect 442 5039 443 5043
rect 447 5042 448 5043
rect 4202 5043 4203 5047
rect 4207 5043 4208 5047
rect 4202 5042 4208 5043
rect 4234 5047 4240 5048
rect 4234 5043 4235 5047
rect 4239 5046 4240 5047
rect 4746 5047 4752 5048
rect 4239 5044 4385 5046
rect 4239 5043 4240 5044
rect 4234 5042 4240 5043
rect 4746 5043 4747 5047
rect 4751 5043 4752 5047
rect 4746 5042 4752 5043
rect 4842 5047 4848 5048
rect 4842 5043 4843 5047
rect 4847 5046 4848 5047
rect 5058 5047 5064 5048
rect 4847 5044 4937 5046
rect 4847 5043 4848 5044
rect 4842 5042 4848 5043
rect 5058 5043 5059 5047
rect 5063 5046 5064 5047
rect 5063 5044 5217 5046
rect 5063 5043 5064 5044
rect 5058 5042 5064 5043
rect 447 5040 618 5042
rect 447 5039 448 5040
rect 442 5038 448 5039
rect 471 5035 477 5036
rect 471 5031 472 5035
rect 476 5034 477 5035
rect 490 5035 496 5036
rect 490 5034 491 5035
rect 476 5032 491 5034
rect 476 5031 477 5032
rect 471 5030 477 5031
rect 490 5031 491 5032
rect 495 5031 496 5035
rect 490 5030 496 5031
rect 606 5035 613 5036
rect 606 5031 607 5035
rect 612 5031 613 5035
rect 616 5034 618 5040
rect 743 5035 749 5036
rect 743 5034 744 5035
rect 616 5032 744 5034
rect 606 5030 613 5031
rect 743 5031 744 5032
rect 748 5031 749 5035
rect 743 5030 749 5031
rect 751 5035 757 5036
rect 751 5031 752 5035
rect 756 5034 757 5035
rect 879 5035 885 5036
rect 879 5034 880 5035
rect 756 5032 880 5034
rect 756 5031 757 5032
rect 751 5030 757 5031
rect 879 5031 880 5032
rect 884 5031 885 5035
rect 879 5030 885 5031
rect 887 5035 893 5036
rect 887 5031 888 5035
rect 892 5034 893 5035
rect 1015 5035 1021 5036
rect 1015 5034 1016 5035
rect 892 5032 1016 5034
rect 892 5031 893 5032
rect 887 5030 893 5031
rect 1015 5031 1016 5032
rect 1020 5031 1021 5035
rect 1015 5030 1021 5031
rect 1023 5035 1029 5036
rect 1023 5031 1024 5035
rect 1028 5034 1029 5035
rect 1159 5035 1165 5036
rect 1159 5034 1160 5035
rect 1028 5032 1160 5034
rect 1028 5031 1029 5032
rect 1023 5030 1029 5031
rect 1159 5031 1160 5032
rect 1164 5031 1165 5035
rect 1159 5030 1165 5031
rect 1311 5035 1317 5036
rect 1311 5031 1312 5035
rect 1316 5034 1317 5035
rect 1346 5035 1352 5036
rect 1346 5034 1347 5035
rect 1316 5032 1347 5034
rect 1316 5031 1317 5032
rect 1311 5030 1317 5031
rect 1346 5031 1347 5032
rect 1351 5031 1352 5035
rect 1346 5030 1352 5031
rect 1423 5035 1429 5036
rect 1423 5031 1424 5035
rect 1428 5034 1429 5035
rect 1463 5035 1469 5036
rect 1463 5034 1464 5035
rect 1428 5032 1464 5034
rect 1428 5031 1429 5032
rect 1423 5030 1429 5031
rect 1463 5031 1464 5032
rect 1468 5031 1469 5035
rect 1463 5030 1469 5031
rect 1615 5035 1621 5036
rect 1615 5031 1616 5035
rect 1620 5034 1621 5035
rect 1658 5035 1664 5036
rect 1658 5034 1659 5035
rect 1620 5032 1659 5034
rect 1620 5031 1621 5032
rect 1615 5030 1621 5031
rect 1658 5031 1659 5032
rect 1663 5031 1664 5035
rect 1658 5030 1664 5031
rect 1775 5035 1784 5036
rect 1775 5031 1776 5035
rect 1783 5031 1784 5035
rect 1775 5030 1784 5031
rect 1910 5035 1917 5036
rect 1910 5031 1911 5035
rect 1916 5031 1917 5035
rect 3863 5035 3869 5036
rect 3863 5034 3864 5035
rect 3820 5032 3864 5034
rect 1910 5030 1917 5031
rect 2118 5031 2125 5032
rect 110 5028 116 5029
rect 1934 5028 1940 5029
rect 110 5024 111 5028
rect 115 5024 116 5028
rect 110 5023 116 5024
rect 346 5027 352 5028
rect 346 5023 347 5027
rect 351 5023 352 5027
rect 346 5022 352 5023
rect 482 5027 488 5028
rect 482 5023 483 5027
rect 487 5023 488 5027
rect 482 5022 488 5023
rect 618 5027 624 5028
rect 618 5023 619 5027
rect 623 5023 624 5027
rect 618 5022 624 5023
rect 754 5027 760 5028
rect 754 5023 755 5027
rect 759 5023 760 5027
rect 754 5022 760 5023
rect 890 5027 896 5028
rect 890 5023 891 5027
rect 895 5023 896 5027
rect 890 5022 896 5023
rect 1034 5027 1040 5028
rect 1034 5023 1035 5027
rect 1039 5023 1040 5027
rect 1034 5022 1040 5023
rect 1186 5027 1192 5028
rect 1186 5023 1187 5027
rect 1191 5023 1192 5027
rect 1186 5022 1192 5023
rect 1338 5027 1344 5028
rect 1338 5023 1339 5027
rect 1343 5023 1344 5027
rect 1338 5022 1344 5023
rect 1490 5027 1496 5028
rect 1490 5023 1491 5027
rect 1495 5023 1496 5027
rect 1490 5022 1496 5023
rect 1650 5027 1656 5028
rect 1650 5023 1651 5027
rect 1655 5023 1656 5027
rect 1650 5022 1656 5023
rect 1786 5027 1792 5028
rect 1786 5023 1787 5027
rect 1791 5023 1792 5027
rect 1934 5024 1935 5028
rect 1939 5024 1940 5028
rect 2118 5027 2119 5031
rect 2124 5027 2125 5031
rect 2118 5026 2125 5027
rect 2655 5031 2661 5032
rect 2655 5027 2656 5031
rect 2660 5030 2661 5031
rect 2767 5031 2773 5032
rect 2767 5030 2768 5031
rect 2660 5028 2768 5030
rect 2660 5027 2661 5028
rect 2655 5026 2661 5027
rect 2767 5027 2768 5028
rect 2772 5027 2773 5031
rect 2767 5026 2773 5027
rect 2954 5031 2960 5032
rect 2954 5027 2955 5031
rect 2959 5030 2960 5031
rect 3223 5031 3229 5032
rect 3223 5030 3224 5031
rect 2959 5028 3224 5030
rect 2959 5027 2960 5028
rect 2954 5026 2960 5027
rect 3223 5027 3224 5028
rect 3228 5027 3229 5031
rect 3223 5026 3229 5027
rect 3775 5031 3781 5032
rect 3775 5027 3776 5031
rect 3780 5030 3781 5031
rect 3820 5030 3822 5032
rect 3863 5031 3864 5032
rect 3868 5031 3869 5035
rect 3863 5030 3869 5031
rect 3780 5028 3822 5030
rect 3780 5027 3781 5028
rect 3775 5026 3781 5027
rect 1934 5023 1940 5024
rect 1974 5024 1980 5025
rect 3798 5024 3804 5025
rect 1786 5022 1792 5023
rect 1974 5020 1975 5024
rect 1979 5020 1980 5024
rect 1974 5019 1980 5020
rect 1994 5023 2000 5024
rect 1994 5019 1995 5023
rect 1999 5019 2000 5023
rect 1994 5018 2000 5019
rect 2530 5023 2536 5024
rect 2530 5019 2531 5023
rect 2535 5019 2536 5023
rect 2530 5018 2536 5019
rect 3098 5023 3104 5024
rect 3098 5019 3099 5023
rect 3103 5019 3104 5023
rect 3098 5018 3104 5019
rect 3650 5023 3656 5024
rect 3650 5019 3651 5023
rect 3655 5019 3656 5023
rect 3798 5020 3799 5024
rect 3803 5020 3804 5024
rect 3798 5019 3804 5020
rect 3650 5018 3656 5019
rect 374 5012 380 5013
rect 110 5011 116 5012
rect 110 5007 111 5011
rect 115 5007 116 5011
rect 374 5008 375 5012
rect 379 5008 380 5012
rect 374 5007 380 5008
rect 510 5012 516 5013
rect 510 5008 511 5012
rect 515 5008 516 5012
rect 510 5007 516 5008
rect 646 5012 652 5013
rect 646 5008 647 5012
rect 651 5008 652 5012
rect 646 5007 652 5008
rect 782 5012 788 5013
rect 782 5008 783 5012
rect 787 5008 788 5012
rect 782 5007 788 5008
rect 918 5012 924 5013
rect 918 5008 919 5012
rect 923 5008 924 5012
rect 918 5007 924 5008
rect 1062 5012 1068 5013
rect 1062 5008 1063 5012
rect 1067 5008 1068 5012
rect 1062 5007 1068 5008
rect 1214 5012 1220 5013
rect 1214 5008 1215 5012
rect 1219 5008 1220 5012
rect 1214 5007 1220 5008
rect 1366 5012 1372 5013
rect 1366 5008 1367 5012
rect 1371 5008 1372 5012
rect 1366 5007 1372 5008
rect 1518 5012 1524 5013
rect 1518 5008 1519 5012
rect 1523 5008 1524 5012
rect 1518 5007 1524 5008
rect 1678 5012 1684 5013
rect 1678 5008 1679 5012
rect 1683 5008 1684 5012
rect 1678 5007 1684 5008
rect 1814 5012 1820 5013
rect 1814 5008 1815 5012
rect 1819 5008 1820 5012
rect 1814 5007 1820 5008
rect 1934 5011 1940 5012
rect 1934 5007 1935 5011
rect 1939 5007 1940 5011
rect 2022 5008 2028 5009
rect 110 5006 116 5007
rect 1934 5006 1940 5007
rect 1974 5007 1980 5008
rect 1974 5003 1975 5007
rect 1979 5003 1980 5007
rect 2022 5004 2023 5008
rect 2027 5004 2028 5008
rect 2022 5003 2028 5004
rect 2558 5008 2564 5009
rect 2558 5004 2559 5008
rect 2563 5004 2564 5008
rect 2558 5003 2564 5004
rect 3126 5008 3132 5009
rect 3126 5004 3127 5008
rect 3131 5004 3132 5008
rect 3126 5003 3132 5004
rect 3678 5008 3684 5009
rect 3678 5004 3679 5008
rect 3683 5004 3684 5008
rect 3678 5003 3684 5004
rect 3798 5007 3804 5008
rect 3798 5003 3799 5007
rect 3803 5003 3804 5007
rect 4818 5007 4824 5008
rect 4818 5006 4819 5007
rect 4628 5004 4819 5006
rect 1974 5002 1980 5003
rect 3798 5002 3804 5003
rect 3954 5003 3960 5004
rect 3954 4999 3955 5003
rect 3959 4999 3960 5003
rect 4628 5002 4630 5004
rect 4818 5003 4819 5004
rect 4823 5003 4824 5007
rect 4818 5002 4824 5003
rect 5247 5003 5253 5004
rect 5247 5002 5248 5003
rect 4509 5000 4630 5002
rect 5165 5000 5248 5002
rect 3954 4998 3960 4999
rect 4026 4999 4032 5000
rect 4026 4995 4027 4999
rect 4031 4995 4032 4999
rect 4026 4994 4032 4995
rect 4218 4999 4224 5000
rect 4218 4995 4219 4999
rect 4223 4995 4224 4999
rect 4218 4994 4224 4995
rect 4634 4999 4640 5000
rect 4634 4995 4635 4999
rect 4639 4995 4640 4999
rect 4634 4994 4640 4995
rect 4850 4999 4856 5000
rect 4850 4995 4851 4999
rect 4855 4995 4856 4999
rect 5247 4999 5248 5000
rect 5252 4999 5253 5003
rect 5247 4998 5253 4999
rect 5334 5003 5340 5004
rect 5334 4999 5335 5003
rect 5339 4999 5340 5003
rect 5334 4998 5340 4999
rect 4850 4994 4856 4995
rect 3983 4959 3989 4960
rect 3983 4955 3984 4959
rect 3988 4958 3989 4959
rect 4026 4959 4032 4960
rect 4026 4958 4027 4959
rect 3988 4956 4027 4958
rect 3988 4955 3989 4956
rect 3983 4954 3989 4955
rect 4026 4955 4027 4956
rect 4031 4955 4032 4959
rect 4026 4954 4032 4955
rect 4143 4959 4149 4960
rect 4143 4955 4144 4959
rect 4148 4958 4149 4959
rect 4218 4959 4224 4960
rect 4218 4958 4219 4959
rect 4148 4956 4219 4958
rect 4148 4955 4149 4956
rect 4143 4954 4149 4955
rect 4218 4955 4219 4956
rect 4223 4955 4224 4959
rect 4218 4954 4224 4955
rect 4334 4959 4341 4960
rect 4334 4955 4335 4959
rect 4340 4955 4341 4959
rect 4334 4954 4341 4955
rect 4535 4959 4541 4960
rect 4535 4955 4536 4959
rect 4540 4958 4541 4959
rect 4634 4959 4640 4960
rect 4634 4958 4635 4959
rect 4540 4956 4635 4958
rect 4540 4955 4541 4956
rect 4535 4954 4541 4955
rect 4634 4955 4635 4956
rect 4639 4955 4640 4959
rect 4634 4954 4640 4955
rect 4746 4959 4757 4960
rect 4746 4955 4747 4959
rect 4751 4955 4752 4959
rect 4756 4955 4757 4959
rect 4746 4954 4757 4955
rect 4818 4959 4824 4960
rect 4818 4955 4819 4959
rect 4823 4958 4824 4959
rect 4967 4959 4973 4960
rect 4967 4958 4968 4959
rect 4823 4956 4968 4958
rect 4823 4955 4824 4956
rect 4818 4954 4824 4955
rect 4967 4955 4968 4956
rect 4972 4955 4973 4959
rect 4967 4954 4973 4955
rect 5190 4959 5197 4960
rect 5190 4955 5191 4959
rect 5196 4955 5197 4959
rect 5190 4954 5197 4955
rect 5247 4959 5253 4960
rect 5247 4955 5248 4959
rect 5252 4958 5253 4959
rect 5423 4959 5429 4960
rect 5423 4958 5424 4959
rect 5252 4956 5424 4958
rect 5252 4955 5253 4956
rect 5247 4954 5253 4955
rect 5423 4955 5424 4956
rect 5428 4955 5429 4959
rect 5423 4954 5429 4955
rect 110 4953 116 4954
rect 1934 4953 1940 4954
rect 110 4949 111 4953
rect 115 4949 116 4953
rect 110 4948 116 4949
rect 158 4952 164 4953
rect 158 4948 159 4952
rect 163 4948 164 4952
rect 158 4947 164 4948
rect 342 4952 348 4953
rect 342 4948 343 4952
rect 347 4948 348 4952
rect 342 4947 348 4948
rect 550 4952 556 4953
rect 550 4948 551 4952
rect 555 4948 556 4952
rect 550 4947 556 4948
rect 750 4952 756 4953
rect 750 4948 751 4952
rect 755 4948 756 4952
rect 750 4947 756 4948
rect 942 4952 948 4953
rect 942 4948 943 4952
rect 947 4948 948 4952
rect 942 4947 948 4948
rect 1126 4952 1132 4953
rect 1126 4948 1127 4952
rect 1131 4948 1132 4952
rect 1126 4947 1132 4948
rect 1310 4952 1316 4953
rect 1310 4948 1311 4952
rect 1315 4948 1316 4952
rect 1310 4947 1316 4948
rect 1486 4952 1492 4953
rect 1486 4948 1487 4952
rect 1491 4948 1492 4952
rect 1486 4947 1492 4948
rect 1662 4952 1668 4953
rect 1662 4948 1663 4952
rect 1667 4948 1668 4952
rect 1662 4947 1668 4948
rect 1814 4952 1820 4953
rect 1814 4948 1815 4952
rect 1819 4948 1820 4952
rect 1934 4949 1935 4953
rect 1939 4949 1940 4953
rect 1934 4948 1940 4949
rect 3838 4952 3844 4953
rect 5662 4952 5668 4953
rect 3838 4948 3839 4952
rect 3843 4948 3844 4952
rect 1814 4947 1820 4948
rect 3838 4947 3844 4948
rect 3858 4951 3864 4952
rect 3858 4947 3859 4951
rect 3863 4947 3864 4951
rect 3858 4946 3864 4947
rect 4018 4951 4024 4952
rect 4018 4947 4019 4951
rect 4023 4947 4024 4951
rect 4018 4946 4024 4947
rect 4210 4951 4216 4952
rect 4210 4947 4211 4951
rect 4215 4947 4216 4951
rect 4210 4946 4216 4947
rect 4410 4951 4416 4952
rect 4410 4947 4411 4951
rect 4415 4947 4416 4951
rect 4410 4946 4416 4947
rect 4626 4951 4632 4952
rect 4626 4947 4627 4951
rect 4631 4947 4632 4951
rect 4626 4946 4632 4947
rect 4842 4951 4848 4952
rect 4842 4947 4843 4951
rect 4847 4947 4848 4951
rect 4842 4946 4848 4947
rect 5066 4951 5072 4952
rect 5066 4947 5067 4951
rect 5071 4947 5072 4951
rect 5066 4946 5072 4947
rect 5298 4951 5304 4952
rect 5298 4947 5299 4951
rect 5303 4947 5304 4951
rect 5662 4948 5663 4952
rect 5667 4948 5668 4952
rect 5662 4947 5668 4948
rect 5298 4946 5304 4947
rect 130 4937 136 4938
rect 110 4936 116 4937
rect 110 4932 111 4936
rect 115 4932 116 4936
rect 130 4933 131 4937
rect 135 4933 136 4937
rect 130 4932 136 4933
rect 314 4937 320 4938
rect 314 4933 315 4937
rect 319 4933 320 4937
rect 314 4932 320 4933
rect 522 4937 528 4938
rect 522 4933 523 4937
rect 527 4933 528 4937
rect 522 4932 528 4933
rect 722 4937 728 4938
rect 722 4933 723 4937
rect 727 4933 728 4937
rect 722 4932 728 4933
rect 914 4937 920 4938
rect 914 4933 915 4937
rect 919 4933 920 4937
rect 914 4932 920 4933
rect 1098 4937 1104 4938
rect 1098 4933 1099 4937
rect 1103 4933 1104 4937
rect 1098 4932 1104 4933
rect 1282 4937 1288 4938
rect 1282 4933 1283 4937
rect 1287 4933 1288 4937
rect 1282 4932 1288 4933
rect 1458 4937 1464 4938
rect 1458 4933 1459 4937
rect 1463 4933 1464 4937
rect 1458 4932 1464 4933
rect 1634 4937 1640 4938
rect 1634 4933 1635 4937
rect 1639 4933 1640 4937
rect 1634 4932 1640 4933
rect 1786 4937 1792 4938
rect 1786 4933 1787 4937
rect 1791 4933 1792 4937
rect 1786 4932 1792 4933
rect 1934 4936 1940 4937
rect 3886 4936 3892 4937
rect 1934 4932 1935 4936
rect 1939 4932 1940 4936
rect 110 4931 116 4932
rect 1934 4931 1940 4932
rect 3838 4935 3844 4936
rect 3838 4931 3839 4935
rect 3843 4931 3844 4935
rect 3886 4932 3887 4936
rect 3891 4932 3892 4936
rect 3886 4931 3892 4932
rect 4046 4936 4052 4937
rect 4046 4932 4047 4936
rect 4051 4932 4052 4936
rect 4046 4931 4052 4932
rect 4238 4936 4244 4937
rect 4238 4932 4239 4936
rect 4243 4932 4244 4936
rect 4238 4931 4244 4932
rect 4438 4936 4444 4937
rect 4438 4932 4439 4936
rect 4443 4932 4444 4936
rect 4438 4931 4444 4932
rect 4654 4936 4660 4937
rect 4654 4932 4655 4936
rect 4659 4932 4660 4936
rect 4654 4931 4660 4932
rect 4870 4936 4876 4937
rect 4870 4932 4871 4936
rect 4875 4932 4876 4936
rect 4870 4931 4876 4932
rect 5094 4936 5100 4937
rect 5094 4932 5095 4936
rect 5099 4932 5100 4936
rect 5094 4931 5100 4932
rect 5326 4936 5332 4937
rect 5326 4932 5327 4936
rect 5331 4932 5332 4936
rect 5326 4931 5332 4932
rect 5662 4935 5668 4936
rect 5662 4931 5663 4935
rect 5667 4931 5668 4935
rect 3838 4930 3844 4931
rect 5662 4930 5668 4931
rect 226 4927 232 4928
rect 226 4923 227 4927
rect 231 4926 232 4927
rect 255 4927 261 4928
rect 255 4926 256 4927
rect 231 4924 256 4926
rect 231 4923 232 4924
rect 226 4922 232 4923
rect 255 4923 256 4924
rect 260 4923 261 4927
rect 255 4922 261 4923
rect 274 4927 280 4928
rect 274 4923 275 4927
rect 279 4926 280 4927
rect 439 4927 445 4928
rect 439 4926 440 4927
rect 279 4924 440 4926
rect 279 4923 280 4924
rect 274 4922 280 4923
rect 439 4923 440 4924
rect 444 4923 445 4927
rect 439 4922 445 4923
rect 647 4927 653 4928
rect 647 4923 648 4927
rect 652 4926 653 4927
rect 686 4927 692 4928
rect 686 4926 687 4927
rect 652 4924 687 4926
rect 652 4923 653 4924
rect 647 4922 653 4923
rect 686 4923 687 4924
rect 691 4923 692 4927
rect 847 4927 853 4928
rect 847 4926 848 4927
rect 686 4922 692 4923
rect 696 4924 848 4926
rect 410 4919 416 4920
rect 410 4915 411 4919
rect 415 4918 416 4919
rect 696 4918 698 4924
rect 847 4923 848 4924
rect 852 4923 853 4927
rect 847 4922 853 4923
rect 1039 4927 1045 4928
rect 1039 4923 1040 4927
rect 1044 4926 1045 4927
rect 1070 4927 1076 4928
rect 1070 4926 1071 4927
rect 1044 4924 1071 4926
rect 1044 4923 1045 4924
rect 1039 4922 1045 4923
rect 1070 4923 1071 4924
rect 1075 4923 1076 4927
rect 1070 4922 1076 4923
rect 1222 4927 1229 4928
rect 1222 4923 1223 4927
rect 1228 4923 1229 4927
rect 1407 4927 1413 4928
rect 1407 4926 1408 4927
rect 1222 4922 1229 4923
rect 1252 4924 1408 4926
rect 415 4916 698 4918
rect 1010 4919 1016 4920
rect 415 4915 416 4916
rect 410 4914 416 4915
rect 1010 4915 1011 4919
rect 1015 4918 1016 4919
rect 1252 4918 1254 4924
rect 1407 4923 1408 4924
rect 1412 4923 1413 4927
rect 1407 4922 1413 4923
rect 1434 4927 1440 4928
rect 1434 4923 1435 4927
rect 1439 4926 1440 4927
rect 1583 4927 1589 4928
rect 1583 4926 1584 4927
rect 1439 4924 1584 4926
rect 1439 4923 1440 4924
rect 1434 4922 1440 4923
rect 1583 4923 1584 4924
rect 1588 4923 1589 4927
rect 1583 4922 1589 4923
rect 1610 4927 1616 4928
rect 1610 4923 1611 4927
rect 1615 4926 1616 4927
rect 1759 4927 1765 4928
rect 1759 4926 1760 4927
rect 1615 4924 1760 4926
rect 1615 4923 1616 4924
rect 1610 4922 1616 4923
rect 1759 4923 1760 4924
rect 1764 4923 1765 4927
rect 1759 4922 1765 4923
rect 1770 4927 1776 4928
rect 1770 4923 1771 4927
rect 1775 4926 1776 4927
rect 1911 4927 1917 4928
rect 1911 4926 1912 4927
rect 1775 4924 1912 4926
rect 1775 4923 1776 4924
rect 1770 4922 1776 4923
rect 1911 4923 1912 4924
rect 1916 4923 1917 4927
rect 1911 4922 1917 4923
rect 1015 4916 1254 4918
rect 1974 4917 1980 4918
rect 3798 4917 3804 4918
rect 1015 4915 1016 4916
rect 1010 4914 1016 4915
rect 1974 4913 1975 4917
rect 1979 4913 1980 4917
rect 1974 4912 1980 4913
rect 2870 4916 2876 4917
rect 2870 4912 2871 4916
rect 2875 4912 2876 4916
rect 2870 4911 2876 4912
rect 3006 4916 3012 4917
rect 3006 4912 3007 4916
rect 3011 4912 3012 4916
rect 3798 4913 3799 4917
rect 3803 4913 3804 4917
rect 3798 4912 3804 4913
rect 3006 4911 3012 4912
rect 2842 4901 2848 4902
rect 1974 4900 1980 4901
rect 1974 4896 1975 4900
rect 1979 4896 1980 4900
rect 2842 4897 2843 4901
rect 2847 4897 2848 4901
rect 2842 4896 2848 4897
rect 2978 4901 2984 4902
rect 2978 4897 2979 4901
rect 2983 4897 2984 4901
rect 2978 4896 2984 4897
rect 3798 4900 3804 4901
rect 3798 4896 3799 4900
rect 3803 4896 3804 4900
rect 1974 4895 1980 4896
rect 3798 4895 3804 4896
rect 2967 4891 2973 4892
rect 274 4887 280 4888
rect 274 4886 275 4887
rect 229 4884 275 4886
rect 274 4883 275 4884
rect 279 4883 280 4887
rect 274 4882 280 4883
rect 410 4887 416 4888
rect 410 4883 411 4887
rect 415 4883 416 4887
rect 410 4882 416 4883
rect 606 4887 612 4888
rect 606 4883 607 4887
rect 611 4883 612 4887
rect 606 4882 612 4883
rect 686 4887 692 4888
rect 686 4883 687 4887
rect 691 4886 692 4887
rect 1010 4887 1016 4888
rect 691 4884 729 4886
rect 691 4883 692 4884
rect 686 4882 692 4883
rect 1010 4883 1011 4887
rect 1015 4883 1016 4887
rect 1010 4882 1016 4883
rect 1070 4887 1076 4888
rect 1070 4883 1071 4887
rect 1075 4886 1076 4887
rect 1434 4887 1440 4888
rect 1434 4886 1435 4887
rect 1075 4884 1105 4886
rect 1381 4884 1435 4886
rect 1075 4883 1076 4884
rect 1070 4882 1076 4883
rect 1434 4883 1435 4884
rect 1439 4883 1440 4887
rect 1610 4887 1616 4888
rect 1610 4886 1611 4887
rect 1557 4884 1611 4886
rect 1434 4882 1440 4883
rect 1610 4883 1611 4884
rect 1615 4883 1616 4887
rect 1770 4887 1776 4888
rect 1770 4886 1771 4887
rect 1733 4884 1771 4886
rect 1610 4882 1616 4883
rect 1770 4883 1771 4884
rect 1775 4883 1776 4887
rect 1770 4882 1776 4883
rect 1778 4887 1784 4888
rect 1778 4883 1779 4887
rect 1783 4886 1784 4887
rect 2967 4887 2968 4891
rect 2972 4890 2973 4891
rect 3018 4891 3024 4892
rect 3018 4890 3019 4891
rect 2972 4888 3019 4890
rect 2972 4887 2973 4888
rect 2967 4886 2973 4887
rect 3018 4887 3019 4888
rect 3023 4887 3024 4891
rect 3103 4891 3109 4892
rect 3103 4890 3104 4891
rect 3018 4886 3024 4887
rect 3028 4888 3104 4890
rect 1783 4884 1793 4886
rect 1783 4883 1784 4884
rect 1778 4882 1784 4883
rect 2938 4883 2944 4884
rect 2938 4879 2939 4883
rect 2943 4882 2944 4883
rect 3028 4882 3030 4888
rect 3103 4887 3104 4888
rect 3108 4887 3109 4891
rect 3103 4886 3109 4887
rect 2943 4880 3030 4882
rect 2943 4879 2944 4880
rect 2938 4878 2944 4879
rect 3838 4857 3844 4858
rect 5662 4857 5668 4858
rect 3838 4853 3839 4857
rect 3843 4853 3844 4857
rect 3838 4852 3844 4853
rect 3886 4856 3892 4857
rect 3886 4852 3887 4856
rect 3891 4852 3892 4856
rect 2938 4851 2944 4852
rect 226 4847 232 4848
rect 226 4843 227 4847
rect 231 4843 232 4847
rect 2938 4847 2939 4851
rect 2943 4847 2944 4851
rect 3146 4851 3152 4852
rect 3886 4851 3892 4852
rect 4070 4856 4076 4857
rect 4070 4852 4071 4856
rect 4075 4852 4076 4856
rect 4070 4851 4076 4852
rect 4286 4856 4292 4857
rect 4286 4852 4287 4856
rect 4291 4852 4292 4856
rect 4286 4851 4292 4852
rect 4510 4856 4516 4857
rect 4510 4852 4511 4856
rect 4515 4852 4516 4856
rect 4510 4851 4516 4852
rect 4734 4856 4740 4857
rect 4734 4852 4735 4856
rect 4739 4852 4740 4856
rect 4734 4851 4740 4852
rect 4958 4856 4964 4857
rect 4958 4852 4959 4856
rect 4963 4852 4964 4856
rect 4958 4851 4964 4852
rect 5182 4856 5188 4857
rect 5182 4852 5183 4856
rect 5187 4852 5188 4856
rect 5182 4851 5188 4852
rect 5406 4856 5412 4857
rect 5406 4852 5407 4856
rect 5411 4852 5412 4856
rect 5662 4853 5663 4857
rect 5667 4853 5668 4857
rect 5662 4852 5668 4853
rect 5406 4851 5412 4852
rect 3146 4850 3147 4851
rect 3077 4848 3147 4850
rect 2938 4846 2944 4847
rect 3146 4847 3147 4848
rect 3151 4847 3152 4851
rect 3146 4846 3152 4847
rect 226 4842 232 4843
rect 274 4843 280 4844
rect 274 4839 275 4843
rect 279 4839 280 4843
rect 274 4838 280 4839
rect 410 4843 416 4844
rect 410 4839 411 4843
rect 415 4839 416 4843
rect 410 4838 416 4839
rect 546 4843 552 4844
rect 546 4839 547 4843
rect 551 4839 552 4843
rect 546 4838 552 4839
rect 682 4843 688 4844
rect 682 4839 683 4843
rect 687 4839 688 4843
rect 3858 4841 3864 4842
rect 682 4838 688 4839
rect 3838 4840 3844 4841
rect 3838 4836 3839 4840
rect 3843 4836 3844 4840
rect 3858 4837 3859 4841
rect 3863 4837 3864 4841
rect 3858 4836 3864 4837
rect 4042 4841 4048 4842
rect 4042 4837 4043 4841
rect 4047 4837 4048 4841
rect 4042 4836 4048 4837
rect 4258 4841 4264 4842
rect 4258 4837 4259 4841
rect 4263 4837 4264 4841
rect 4258 4836 4264 4837
rect 4482 4841 4488 4842
rect 4482 4837 4483 4841
rect 4487 4837 4488 4841
rect 4482 4836 4488 4837
rect 4706 4841 4712 4842
rect 4706 4837 4707 4841
rect 4711 4837 4712 4841
rect 4706 4836 4712 4837
rect 4930 4841 4936 4842
rect 4930 4837 4931 4841
rect 4935 4837 4936 4841
rect 4930 4836 4936 4837
rect 5154 4841 5160 4842
rect 5154 4837 5155 4841
rect 5159 4837 5160 4841
rect 5154 4836 5160 4837
rect 5378 4841 5384 4842
rect 5378 4837 5379 4841
rect 5383 4837 5384 4841
rect 5378 4836 5384 4837
rect 5662 4840 5668 4841
rect 5662 4836 5663 4840
rect 5667 4836 5668 4840
rect 3838 4835 3844 4836
rect 5662 4835 5668 4836
rect 3982 4831 3989 4832
rect 3982 4827 3983 4831
rect 3988 4827 3989 4831
rect 3982 4826 3989 4827
rect 4015 4831 4021 4832
rect 4015 4827 4016 4831
rect 4020 4830 4021 4831
rect 4167 4831 4173 4832
rect 4167 4830 4168 4831
rect 4020 4828 4168 4830
rect 4020 4827 4021 4828
rect 4015 4826 4021 4827
rect 4167 4827 4168 4828
rect 4172 4827 4173 4831
rect 4167 4826 4173 4827
rect 4255 4831 4261 4832
rect 4255 4827 4256 4831
rect 4260 4830 4261 4831
rect 4383 4831 4389 4832
rect 4383 4830 4384 4831
rect 4260 4828 4384 4830
rect 4260 4827 4261 4828
rect 4255 4826 4261 4827
rect 4383 4827 4384 4828
rect 4388 4827 4389 4831
rect 4383 4826 4389 4827
rect 4607 4831 4616 4832
rect 4607 4827 4608 4831
rect 4615 4827 4616 4831
rect 4607 4826 4616 4827
rect 4831 4831 4837 4832
rect 4831 4827 4832 4831
rect 4836 4830 4837 4831
rect 4850 4831 4856 4832
rect 4850 4830 4851 4831
rect 4836 4828 4851 4830
rect 4836 4827 4837 4828
rect 4831 4826 4837 4827
rect 4850 4827 4851 4828
rect 4855 4827 4856 4831
rect 5055 4831 5061 4832
rect 5055 4830 5056 4831
rect 4850 4826 4856 4827
rect 4884 4828 5056 4830
rect 4578 4823 4584 4824
rect 4578 4819 4579 4823
rect 4583 4822 4584 4823
rect 4884 4822 4886 4828
rect 5055 4827 5056 4828
rect 5060 4827 5061 4831
rect 5055 4826 5061 4827
rect 5279 4831 5285 4832
rect 5279 4827 5280 4831
rect 5284 4830 5285 4831
rect 5287 4831 5293 4832
rect 5287 4830 5288 4831
rect 5284 4828 5288 4830
rect 5284 4827 5285 4828
rect 5279 4826 5285 4827
rect 5287 4827 5288 4828
rect 5292 4827 5293 4831
rect 5287 4826 5293 4827
rect 5466 4831 5472 4832
rect 5466 4827 5467 4831
rect 5471 4830 5472 4831
rect 5503 4831 5509 4832
rect 5503 4830 5504 4831
rect 5471 4828 5504 4830
rect 5471 4827 5472 4828
rect 5466 4826 5472 4827
rect 5503 4827 5504 4828
rect 5508 4827 5509 4831
rect 5503 4826 5509 4827
rect 4583 4820 4886 4822
rect 4583 4819 4584 4820
rect 4578 4818 4584 4819
rect 255 4803 261 4804
rect 255 4799 256 4803
rect 260 4802 261 4803
rect 274 4803 280 4804
rect 274 4802 275 4803
rect 260 4800 275 4802
rect 260 4799 261 4800
rect 255 4798 261 4799
rect 274 4799 275 4800
rect 279 4799 280 4803
rect 274 4798 280 4799
rect 391 4803 397 4804
rect 391 4799 392 4803
rect 396 4802 397 4803
rect 410 4803 416 4804
rect 410 4802 411 4803
rect 396 4800 411 4802
rect 396 4799 397 4800
rect 391 4798 397 4799
rect 410 4799 411 4800
rect 415 4799 416 4803
rect 410 4798 416 4799
rect 527 4803 533 4804
rect 527 4799 528 4803
rect 532 4802 533 4803
rect 546 4803 552 4804
rect 546 4802 547 4803
rect 532 4800 547 4802
rect 532 4799 533 4800
rect 527 4798 533 4799
rect 546 4799 547 4800
rect 551 4799 552 4803
rect 546 4798 552 4799
rect 663 4803 669 4804
rect 663 4799 664 4803
rect 668 4802 669 4803
rect 682 4803 688 4804
rect 682 4802 683 4803
rect 668 4800 683 4802
rect 668 4799 669 4800
rect 663 4798 669 4799
rect 682 4799 683 4800
rect 687 4799 688 4803
rect 682 4798 688 4799
rect 690 4803 696 4804
rect 690 4799 691 4803
rect 695 4802 696 4803
rect 799 4803 805 4804
rect 799 4802 800 4803
rect 695 4800 800 4802
rect 695 4799 696 4800
rect 690 4798 696 4799
rect 799 4799 800 4800
rect 804 4799 805 4803
rect 799 4798 805 4799
rect 110 4796 116 4797
rect 1934 4796 1940 4797
rect 110 4792 111 4796
rect 115 4792 116 4796
rect 110 4791 116 4792
rect 130 4795 136 4796
rect 130 4791 131 4795
rect 135 4791 136 4795
rect 130 4790 136 4791
rect 266 4795 272 4796
rect 266 4791 267 4795
rect 271 4791 272 4795
rect 266 4790 272 4791
rect 402 4795 408 4796
rect 402 4791 403 4795
rect 407 4791 408 4795
rect 402 4790 408 4791
rect 538 4795 544 4796
rect 538 4791 539 4795
rect 543 4791 544 4795
rect 538 4790 544 4791
rect 674 4795 680 4796
rect 674 4791 675 4795
rect 679 4791 680 4795
rect 1934 4792 1935 4796
rect 1939 4792 1940 4796
rect 1934 4791 1940 4792
rect 1966 4795 1972 4796
rect 1966 4791 1967 4795
rect 1971 4794 1972 4795
rect 2790 4795 2796 4796
rect 1971 4792 2001 4794
rect 1971 4791 1972 4792
rect 674 4790 680 4791
rect 1966 4790 1972 4791
rect 2162 4791 2168 4792
rect 2162 4787 2163 4791
rect 2167 4787 2168 4791
rect 2162 4786 2168 4787
rect 2354 4791 2360 4792
rect 2354 4787 2355 4791
rect 2359 4787 2360 4791
rect 2354 4786 2360 4787
rect 2546 4791 2552 4792
rect 2546 4787 2547 4791
rect 2551 4787 2552 4791
rect 2790 4791 2791 4795
rect 2795 4791 2796 4795
rect 2790 4790 2796 4791
rect 2938 4791 2944 4792
rect 2546 4786 2552 4787
rect 2938 4787 2939 4791
rect 2943 4787 2944 4791
rect 2938 4786 2944 4787
rect 3138 4791 3144 4792
rect 3138 4787 3139 4791
rect 3143 4787 3144 4791
rect 4015 4791 4021 4792
rect 4015 4790 4016 4791
rect 3957 4788 4016 4790
rect 3138 4786 3144 4787
rect 4015 4787 4016 4788
rect 4020 4787 4021 4791
rect 4255 4791 4261 4792
rect 4255 4790 4256 4791
rect 4141 4788 4256 4790
rect 4015 4786 4021 4787
rect 4255 4787 4256 4788
rect 4260 4787 4261 4791
rect 4255 4786 4261 4787
rect 4334 4791 4340 4792
rect 4334 4787 4335 4791
rect 4339 4787 4340 4791
rect 4334 4786 4340 4787
rect 4578 4791 4584 4792
rect 4578 4787 4579 4791
rect 4583 4787 4584 4791
rect 4578 4786 4584 4787
rect 4610 4791 4616 4792
rect 4610 4787 4611 4791
rect 4615 4790 4616 4791
rect 5082 4791 5088 4792
rect 5082 4790 5083 4791
rect 4615 4788 4713 4790
rect 5029 4788 5083 4790
rect 4615 4787 4616 4788
rect 4610 4786 4616 4787
rect 5082 4787 5083 4788
rect 5087 4787 5088 4791
rect 5082 4786 5088 4787
rect 5190 4791 5196 4792
rect 5190 4787 5191 4791
rect 5195 4787 5196 4791
rect 5190 4786 5196 4787
rect 5287 4791 5293 4792
rect 5287 4787 5288 4791
rect 5292 4790 5293 4791
rect 5292 4788 5385 4790
rect 5292 4787 5293 4788
rect 5287 4786 5293 4787
rect 158 4780 164 4781
rect 110 4779 116 4780
rect 110 4775 111 4779
rect 115 4775 116 4779
rect 158 4776 159 4780
rect 163 4776 164 4780
rect 158 4775 164 4776
rect 294 4780 300 4781
rect 294 4776 295 4780
rect 299 4776 300 4780
rect 294 4775 300 4776
rect 430 4780 436 4781
rect 430 4776 431 4780
rect 435 4776 436 4780
rect 430 4775 436 4776
rect 566 4780 572 4781
rect 566 4776 567 4780
rect 571 4776 572 4780
rect 566 4775 572 4776
rect 702 4780 708 4781
rect 702 4776 703 4780
rect 707 4776 708 4780
rect 702 4775 708 4776
rect 1934 4779 1940 4780
rect 1934 4775 1935 4779
rect 1939 4775 1940 4779
rect 110 4774 116 4775
rect 1934 4774 1940 4775
rect 3982 4755 3988 4756
rect 2119 4751 2125 4752
rect 2119 4747 2120 4751
rect 2124 4750 2125 4751
rect 2162 4751 2168 4752
rect 2162 4750 2163 4751
rect 2124 4748 2163 4750
rect 2124 4747 2125 4748
rect 2119 4746 2125 4747
rect 2162 4747 2163 4748
rect 2167 4747 2168 4751
rect 2162 4746 2168 4747
rect 2279 4751 2285 4752
rect 2279 4747 2280 4751
rect 2284 4750 2285 4751
rect 2354 4751 2360 4752
rect 2354 4750 2355 4751
rect 2284 4748 2355 4750
rect 2284 4747 2285 4748
rect 2279 4746 2285 4747
rect 2354 4747 2355 4748
rect 2359 4747 2360 4751
rect 2354 4746 2360 4747
rect 2471 4751 2477 4752
rect 2471 4747 2472 4751
rect 2476 4750 2477 4751
rect 2546 4751 2552 4752
rect 2546 4750 2547 4751
rect 2476 4748 2547 4750
rect 2476 4747 2477 4748
rect 2471 4746 2477 4747
rect 2546 4747 2547 4748
rect 2551 4747 2552 4751
rect 2546 4746 2552 4747
rect 2658 4751 2669 4752
rect 2658 4747 2659 4751
rect 2663 4747 2664 4751
rect 2668 4747 2669 4751
rect 2658 4746 2669 4747
rect 2855 4751 2861 4752
rect 2855 4747 2856 4751
rect 2860 4750 2861 4751
rect 2938 4751 2944 4752
rect 2938 4750 2939 4751
rect 2860 4748 2939 4750
rect 2860 4747 2861 4748
rect 2855 4746 2861 4747
rect 2938 4747 2939 4748
rect 2943 4747 2944 4751
rect 2938 4746 2944 4747
rect 3055 4751 3061 4752
rect 3055 4747 3056 4751
rect 3060 4750 3061 4751
rect 3138 4751 3144 4752
rect 3138 4750 3139 4751
rect 3060 4748 3139 4750
rect 3060 4747 3061 4748
rect 3055 4746 3061 4747
rect 3138 4747 3139 4748
rect 3143 4747 3144 4751
rect 3138 4746 3144 4747
rect 3146 4751 3152 4752
rect 3146 4747 3147 4751
rect 3151 4750 3152 4751
rect 3255 4751 3261 4752
rect 3255 4750 3256 4751
rect 3151 4748 3256 4750
rect 3151 4747 3152 4748
rect 3146 4746 3152 4747
rect 3255 4747 3256 4748
rect 3260 4747 3261 4751
rect 3982 4751 3983 4755
rect 3987 4751 3988 4755
rect 5466 4755 5472 4756
rect 3982 4750 3988 4751
rect 4194 4751 4200 4752
rect 3255 4746 3261 4747
rect 4194 4747 4195 4751
rect 4199 4747 4200 4751
rect 4194 4746 4200 4747
rect 4474 4751 4480 4752
rect 4474 4747 4475 4751
rect 4479 4747 4480 4751
rect 4474 4746 4480 4747
rect 4858 4751 4864 4752
rect 4858 4747 4859 4751
rect 4863 4747 4864 4751
rect 4858 4746 4864 4747
rect 5074 4751 5080 4752
rect 5074 4747 5075 4751
rect 5079 4747 5080 4751
rect 5466 4751 5467 4755
rect 5471 4751 5472 4755
rect 5466 4750 5472 4751
rect 5074 4746 5080 4747
rect 1974 4744 1980 4745
rect 3798 4744 3804 4745
rect 226 4743 232 4744
rect 226 4739 227 4743
rect 231 4742 232 4743
rect 690 4743 696 4744
rect 690 4742 691 4743
rect 231 4740 691 4742
rect 231 4739 232 4740
rect 226 4738 232 4739
rect 690 4739 691 4740
rect 695 4739 696 4743
rect 1974 4740 1975 4744
rect 1979 4740 1980 4744
rect 1974 4739 1980 4740
rect 1994 4743 2000 4744
rect 1994 4739 1995 4743
rect 1999 4739 2000 4743
rect 690 4738 696 4739
rect 1994 4738 2000 4739
rect 2154 4743 2160 4744
rect 2154 4739 2155 4743
rect 2159 4739 2160 4743
rect 2154 4738 2160 4739
rect 2346 4743 2352 4744
rect 2346 4739 2347 4743
rect 2351 4739 2352 4743
rect 2346 4738 2352 4739
rect 2538 4743 2544 4744
rect 2538 4739 2539 4743
rect 2543 4739 2544 4743
rect 2538 4738 2544 4739
rect 2730 4743 2736 4744
rect 2730 4739 2731 4743
rect 2735 4739 2736 4743
rect 2730 4738 2736 4739
rect 2930 4743 2936 4744
rect 2930 4739 2931 4743
rect 2935 4739 2936 4743
rect 2930 4738 2936 4739
rect 3130 4743 3136 4744
rect 3130 4739 3131 4743
rect 3135 4739 3136 4743
rect 3798 4740 3799 4744
rect 3803 4740 3804 4744
rect 3798 4739 3804 4740
rect 3130 4738 3136 4739
rect 2022 4728 2028 4729
rect 1974 4727 1980 4728
rect 1974 4723 1975 4727
rect 1979 4723 1980 4727
rect 2022 4724 2023 4728
rect 2027 4724 2028 4728
rect 2022 4723 2028 4724
rect 2182 4728 2188 4729
rect 2182 4724 2183 4728
rect 2187 4724 2188 4728
rect 2182 4723 2188 4724
rect 2374 4728 2380 4729
rect 2374 4724 2375 4728
rect 2379 4724 2380 4728
rect 2374 4723 2380 4724
rect 2566 4728 2572 4729
rect 2566 4724 2567 4728
rect 2571 4724 2572 4728
rect 2566 4723 2572 4724
rect 2758 4728 2764 4729
rect 2758 4724 2759 4728
rect 2763 4724 2764 4728
rect 2758 4723 2764 4724
rect 2958 4728 2964 4729
rect 2958 4724 2959 4728
rect 2963 4724 2964 4728
rect 2958 4723 2964 4724
rect 3158 4728 3164 4729
rect 3158 4724 3159 4728
rect 3163 4724 3164 4728
rect 3158 4723 3164 4724
rect 3798 4727 3804 4728
rect 3798 4723 3799 4727
rect 3803 4723 3804 4727
rect 1974 4722 1980 4723
rect 3798 4722 3804 4723
rect 110 4713 116 4714
rect 1934 4713 1940 4714
rect 110 4709 111 4713
rect 115 4709 116 4713
rect 110 4708 116 4709
rect 158 4712 164 4713
rect 158 4708 159 4712
rect 163 4708 164 4712
rect 158 4707 164 4708
rect 342 4712 348 4713
rect 342 4708 343 4712
rect 347 4708 348 4712
rect 342 4707 348 4708
rect 566 4712 572 4713
rect 566 4708 567 4712
rect 571 4708 572 4712
rect 566 4707 572 4708
rect 806 4712 812 4713
rect 806 4708 807 4712
rect 811 4708 812 4712
rect 806 4707 812 4708
rect 1054 4712 1060 4713
rect 1054 4708 1055 4712
rect 1059 4708 1060 4712
rect 1054 4707 1060 4708
rect 1310 4712 1316 4713
rect 1310 4708 1311 4712
rect 1315 4708 1316 4712
rect 1310 4707 1316 4708
rect 1574 4712 1580 4713
rect 1574 4708 1575 4712
rect 1579 4708 1580 4712
rect 1574 4707 1580 4708
rect 1814 4712 1820 4713
rect 1814 4708 1815 4712
rect 1819 4708 1820 4712
rect 1934 4709 1935 4713
rect 1939 4709 1940 4713
rect 1934 4708 1940 4709
rect 4039 4711 4045 4712
rect 1814 4707 1820 4708
rect 4039 4707 4040 4711
rect 4044 4710 4045 4711
rect 4194 4711 4200 4712
rect 4194 4710 4195 4711
rect 4044 4708 4195 4710
rect 4044 4707 4045 4708
rect 4039 4706 4045 4707
rect 4194 4707 4195 4708
rect 4199 4707 4200 4711
rect 4194 4706 4200 4707
rect 4311 4711 4317 4712
rect 4311 4707 4312 4711
rect 4316 4710 4317 4711
rect 4474 4711 4480 4712
rect 4474 4710 4475 4711
rect 4316 4708 4475 4710
rect 4316 4707 4317 4708
rect 4311 4706 4317 4707
rect 4474 4707 4475 4708
rect 4479 4707 4480 4711
rect 4474 4706 4480 4707
rect 4590 4711 4597 4712
rect 4590 4707 4591 4711
rect 4596 4707 4597 4711
rect 4590 4706 4597 4707
rect 4887 4711 4893 4712
rect 4887 4707 4888 4711
rect 4892 4710 4893 4711
rect 5074 4711 5080 4712
rect 5074 4710 5075 4711
rect 4892 4708 5075 4710
rect 4892 4707 4893 4708
rect 4887 4706 4893 4707
rect 5074 4707 5075 4708
rect 5079 4707 5080 4711
rect 5074 4706 5080 4707
rect 5082 4711 5088 4712
rect 5082 4707 5083 4711
rect 5087 4710 5088 4711
rect 5191 4711 5197 4712
rect 5191 4710 5192 4711
rect 5087 4708 5192 4710
rect 5087 4707 5088 4708
rect 5082 4706 5088 4707
rect 5191 4707 5192 4708
rect 5196 4707 5197 4711
rect 5191 4706 5197 4707
rect 5494 4711 5501 4712
rect 5494 4707 5495 4711
rect 5500 4707 5501 4711
rect 5494 4706 5501 4707
rect 3838 4704 3844 4705
rect 5662 4704 5668 4705
rect 3838 4700 3839 4704
rect 3843 4700 3844 4704
rect 3838 4699 3844 4700
rect 3914 4703 3920 4704
rect 3914 4699 3915 4703
rect 3919 4699 3920 4703
rect 3914 4698 3920 4699
rect 4186 4703 4192 4704
rect 4186 4699 4187 4703
rect 4191 4699 4192 4703
rect 4186 4698 4192 4699
rect 4466 4703 4472 4704
rect 4466 4699 4467 4703
rect 4471 4699 4472 4703
rect 4466 4698 4472 4699
rect 4762 4703 4768 4704
rect 4762 4699 4763 4703
rect 4767 4699 4768 4703
rect 4762 4698 4768 4699
rect 5066 4703 5072 4704
rect 5066 4699 5067 4703
rect 5071 4699 5072 4703
rect 5066 4698 5072 4699
rect 5370 4703 5376 4704
rect 5370 4699 5371 4703
rect 5375 4699 5376 4703
rect 5662 4700 5663 4704
rect 5667 4700 5668 4704
rect 5662 4699 5668 4700
rect 5370 4698 5376 4699
rect 130 4697 136 4698
rect 110 4696 116 4697
rect 110 4692 111 4696
rect 115 4692 116 4696
rect 130 4693 131 4697
rect 135 4693 136 4697
rect 130 4692 136 4693
rect 314 4697 320 4698
rect 314 4693 315 4697
rect 319 4693 320 4697
rect 314 4692 320 4693
rect 538 4697 544 4698
rect 538 4693 539 4697
rect 543 4693 544 4697
rect 538 4692 544 4693
rect 778 4697 784 4698
rect 778 4693 779 4697
rect 783 4693 784 4697
rect 778 4692 784 4693
rect 1026 4697 1032 4698
rect 1026 4693 1027 4697
rect 1031 4693 1032 4697
rect 1026 4692 1032 4693
rect 1282 4697 1288 4698
rect 1282 4693 1283 4697
rect 1287 4693 1288 4697
rect 1282 4692 1288 4693
rect 1546 4697 1552 4698
rect 1546 4693 1547 4697
rect 1551 4693 1552 4697
rect 1546 4692 1552 4693
rect 1786 4697 1792 4698
rect 1786 4693 1787 4697
rect 1791 4693 1792 4697
rect 1786 4692 1792 4693
rect 1934 4696 1940 4697
rect 1934 4692 1935 4696
rect 1939 4692 1940 4696
rect 110 4691 116 4692
rect 1934 4691 1940 4692
rect 3942 4688 3948 4689
rect 255 4687 261 4688
rect 255 4683 256 4687
rect 260 4686 261 4687
rect 287 4687 293 4688
rect 287 4686 288 4687
rect 260 4684 288 4686
rect 260 4683 261 4684
rect 255 4682 261 4683
rect 287 4683 288 4684
rect 292 4683 293 4687
rect 287 4682 293 4683
rect 439 4687 448 4688
rect 439 4683 440 4687
rect 447 4683 448 4687
rect 439 4682 448 4683
rect 663 4687 672 4688
rect 663 4683 664 4687
rect 671 4683 672 4687
rect 663 4682 672 4683
rect 903 4687 912 4688
rect 903 4683 904 4687
rect 911 4683 912 4687
rect 903 4682 912 4683
rect 1010 4687 1016 4688
rect 1010 4683 1011 4687
rect 1015 4686 1016 4687
rect 1151 4687 1157 4688
rect 1151 4686 1152 4687
rect 1015 4684 1152 4686
rect 1015 4683 1016 4684
rect 1010 4682 1016 4683
rect 1151 4683 1152 4684
rect 1156 4683 1157 4687
rect 1151 4682 1157 4683
rect 1407 4687 1416 4688
rect 1407 4683 1408 4687
rect 1415 4683 1416 4687
rect 1407 4682 1416 4683
rect 1671 4687 1680 4688
rect 1671 4683 1672 4687
rect 1679 4683 1680 4687
rect 1671 4682 1680 4683
rect 1911 4687 1917 4688
rect 1911 4683 1912 4687
rect 1916 4686 1917 4687
rect 1966 4687 1972 4688
rect 1966 4686 1967 4687
rect 1916 4684 1967 4686
rect 1916 4683 1917 4684
rect 1911 4682 1917 4683
rect 1966 4683 1967 4684
rect 1971 4683 1972 4687
rect 1966 4682 1972 4683
rect 3838 4687 3844 4688
rect 3838 4683 3839 4687
rect 3843 4683 3844 4687
rect 3942 4684 3943 4688
rect 3947 4684 3948 4688
rect 3942 4683 3948 4684
rect 4214 4688 4220 4689
rect 4214 4684 4215 4688
rect 4219 4684 4220 4688
rect 4214 4683 4220 4684
rect 4494 4688 4500 4689
rect 4494 4684 4495 4688
rect 4499 4684 4500 4688
rect 4494 4683 4500 4684
rect 4790 4688 4796 4689
rect 4790 4684 4791 4688
rect 4795 4684 4796 4688
rect 4790 4683 4796 4684
rect 5094 4688 5100 4689
rect 5094 4684 5095 4688
rect 5099 4684 5100 4688
rect 5094 4683 5100 4684
rect 5398 4688 5404 4689
rect 5398 4684 5399 4688
rect 5403 4684 5404 4688
rect 5398 4683 5404 4684
rect 5662 4687 5668 4688
rect 5662 4683 5663 4687
rect 5667 4683 5668 4687
rect 3838 4682 3844 4683
rect 5662 4682 5668 4683
rect 1974 4665 1980 4666
rect 3798 4665 3804 4666
rect 1974 4661 1975 4665
rect 1979 4661 1980 4665
rect 1974 4660 1980 4661
rect 2022 4664 2028 4665
rect 2022 4660 2023 4664
rect 2027 4660 2028 4664
rect 2022 4659 2028 4660
rect 2238 4664 2244 4665
rect 2238 4660 2239 4664
rect 2243 4660 2244 4664
rect 2238 4659 2244 4660
rect 2470 4664 2476 4665
rect 2470 4660 2471 4664
rect 2475 4660 2476 4664
rect 2470 4659 2476 4660
rect 2694 4664 2700 4665
rect 2694 4660 2695 4664
rect 2699 4660 2700 4664
rect 2694 4659 2700 4660
rect 2918 4664 2924 4665
rect 2918 4660 2919 4664
rect 2923 4660 2924 4664
rect 2918 4659 2924 4660
rect 3142 4664 3148 4665
rect 3142 4660 3143 4664
rect 3147 4660 3148 4664
rect 3142 4659 3148 4660
rect 3366 4664 3372 4665
rect 3366 4660 3367 4664
rect 3371 4660 3372 4664
rect 3798 4661 3799 4665
rect 3803 4661 3804 4665
rect 3798 4660 3804 4661
rect 3366 4659 3372 4660
rect 1994 4649 2000 4650
rect 1974 4648 1980 4649
rect 226 4647 232 4648
rect 226 4643 227 4647
rect 231 4643 232 4647
rect 226 4642 232 4643
rect 287 4647 293 4648
rect 287 4643 288 4647
rect 292 4646 293 4647
rect 442 4647 448 4648
rect 292 4644 321 4646
rect 292 4643 293 4644
rect 287 4642 293 4643
rect 442 4643 443 4647
rect 447 4646 448 4647
rect 666 4647 672 4648
rect 447 4644 545 4646
rect 447 4643 448 4644
rect 442 4642 448 4643
rect 666 4643 667 4647
rect 671 4646 672 4647
rect 906 4647 912 4648
rect 671 4644 785 4646
rect 671 4643 672 4644
rect 666 4642 672 4643
rect 906 4643 907 4647
rect 911 4646 912 4647
rect 1410 4647 1416 4648
rect 911 4644 1033 4646
rect 911 4643 912 4644
rect 906 4642 912 4643
rect 1380 4638 1382 4645
rect 1410 4643 1411 4647
rect 1415 4646 1416 4647
rect 1674 4647 1680 4648
rect 1415 4644 1553 4646
rect 1415 4643 1416 4644
rect 1410 4642 1416 4643
rect 1674 4643 1675 4647
rect 1679 4646 1680 4647
rect 1679 4644 1793 4646
rect 1974 4644 1975 4648
rect 1979 4644 1980 4648
rect 1994 4645 1995 4649
rect 1999 4645 2000 4649
rect 1994 4644 2000 4645
rect 2210 4649 2216 4650
rect 2210 4645 2211 4649
rect 2215 4645 2216 4649
rect 2210 4644 2216 4645
rect 2442 4649 2448 4650
rect 2442 4645 2443 4649
rect 2447 4645 2448 4649
rect 2442 4644 2448 4645
rect 2666 4649 2672 4650
rect 2666 4645 2667 4649
rect 2671 4645 2672 4649
rect 2666 4644 2672 4645
rect 2890 4649 2896 4650
rect 2890 4645 2891 4649
rect 2895 4645 2896 4649
rect 2890 4644 2896 4645
rect 3114 4649 3120 4650
rect 3114 4645 3115 4649
rect 3119 4645 3120 4649
rect 3114 4644 3120 4645
rect 3338 4649 3344 4650
rect 3338 4645 3339 4649
rect 3343 4645 3344 4649
rect 3338 4644 3344 4645
rect 3798 4648 3804 4649
rect 3798 4644 3799 4648
rect 3803 4644 3804 4648
rect 1679 4643 1680 4644
rect 1974 4643 1980 4644
rect 3798 4643 3804 4644
rect 1674 4642 1680 4643
rect 1518 4639 1524 4640
rect 1518 4638 1519 4639
rect 1380 4636 1519 4638
rect 1518 4635 1519 4636
rect 1523 4635 1524 4639
rect 1518 4634 1524 4635
rect 2119 4639 2125 4640
rect 2119 4635 2120 4639
rect 2124 4638 2125 4639
rect 2167 4639 2173 4640
rect 2167 4638 2168 4639
rect 2124 4636 2168 4638
rect 2124 4635 2125 4636
rect 2119 4634 2125 4635
rect 2167 4635 2168 4636
rect 2172 4635 2173 4639
rect 2167 4634 2173 4635
rect 2335 4639 2344 4640
rect 2335 4635 2336 4639
rect 2343 4635 2344 4639
rect 2335 4634 2344 4635
rect 2567 4639 2573 4640
rect 2567 4635 2568 4639
rect 2572 4638 2573 4639
rect 2575 4639 2581 4640
rect 2575 4638 2576 4639
rect 2572 4636 2576 4638
rect 2572 4635 2573 4636
rect 2567 4634 2573 4635
rect 2575 4635 2576 4636
rect 2580 4635 2581 4639
rect 2575 4634 2581 4635
rect 2790 4639 2797 4640
rect 2790 4635 2791 4639
rect 2796 4635 2797 4639
rect 2790 4634 2797 4635
rect 2882 4639 2888 4640
rect 2882 4635 2883 4639
rect 2887 4638 2888 4639
rect 3015 4639 3021 4640
rect 3015 4638 3016 4639
rect 2887 4636 3016 4638
rect 2887 4635 2888 4636
rect 2882 4634 2888 4635
rect 3015 4635 3016 4636
rect 3020 4635 3021 4639
rect 3015 4634 3021 4635
rect 3239 4639 3248 4640
rect 3239 4635 3240 4639
rect 3247 4635 3248 4639
rect 3463 4639 3469 4640
rect 3463 4638 3464 4639
rect 3239 4634 3248 4635
rect 3252 4636 3464 4638
rect 2986 4631 2992 4632
rect 2986 4627 2987 4631
rect 2991 4630 2992 4631
rect 3252 4630 3254 4636
rect 3463 4635 3464 4636
rect 3468 4635 3469 4639
rect 3463 4634 3469 4635
rect 2991 4628 3254 4630
rect 3838 4629 3844 4630
rect 5662 4629 5668 4630
rect 2991 4627 2992 4628
rect 2986 4626 2992 4627
rect 3838 4625 3839 4629
rect 3843 4625 3844 4629
rect 3838 4624 3844 4625
rect 4062 4628 4068 4629
rect 4062 4624 4063 4628
rect 4067 4624 4068 4628
rect 4062 4623 4068 4624
rect 4326 4628 4332 4629
rect 4326 4624 4327 4628
rect 4331 4624 4332 4628
rect 4326 4623 4332 4624
rect 4598 4628 4604 4629
rect 4598 4624 4599 4628
rect 4603 4624 4604 4628
rect 4598 4623 4604 4624
rect 4870 4628 4876 4629
rect 4870 4624 4871 4628
rect 4875 4624 4876 4628
rect 4870 4623 4876 4624
rect 5150 4628 5156 4629
rect 5150 4624 5151 4628
rect 5155 4624 5156 4628
rect 5150 4623 5156 4624
rect 5438 4628 5444 4629
rect 5438 4624 5439 4628
rect 5443 4624 5444 4628
rect 5662 4625 5663 4629
rect 5667 4625 5668 4629
rect 5662 4624 5668 4625
rect 5438 4623 5444 4624
rect 4034 4613 4040 4614
rect 3838 4612 3844 4613
rect 3838 4608 3839 4612
rect 3843 4608 3844 4612
rect 4034 4609 4035 4613
rect 4039 4609 4040 4613
rect 4034 4608 4040 4609
rect 4298 4613 4304 4614
rect 4298 4609 4299 4613
rect 4303 4609 4304 4613
rect 4298 4608 4304 4609
rect 4570 4613 4576 4614
rect 4570 4609 4571 4613
rect 4575 4609 4576 4613
rect 4570 4608 4576 4609
rect 4842 4613 4848 4614
rect 4842 4609 4843 4613
rect 4847 4609 4848 4613
rect 4842 4608 4848 4609
rect 5122 4613 5128 4614
rect 5122 4609 5123 4613
rect 5127 4609 5128 4613
rect 5122 4608 5128 4609
rect 5410 4613 5416 4614
rect 5410 4609 5411 4613
rect 5415 4609 5416 4613
rect 5410 4608 5416 4609
rect 5662 4612 5668 4613
rect 5662 4608 5663 4612
rect 5667 4608 5668 4612
rect 3838 4607 3844 4608
rect 5662 4607 5668 4608
rect 1010 4603 1016 4604
rect 1010 4602 1011 4603
rect 396 4600 1011 4602
rect 396 4598 398 4600
rect 1010 4599 1011 4600
rect 1015 4599 1016 4603
rect 1906 4603 1912 4604
rect 1906 4602 1907 4603
rect 1010 4598 1016 4599
rect 1784 4600 1907 4602
rect 1784 4598 1786 4600
rect 1906 4599 1907 4600
rect 1911 4599 1912 4603
rect 4159 4603 4165 4604
rect 1906 4598 1912 4599
rect 2167 4599 2173 4600
rect 269 4596 398 4598
rect 1589 4596 1786 4598
rect 402 4595 408 4596
rect 402 4591 403 4595
rect 407 4591 408 4595
rect 402 4590 408 4591
rect 650 4595 656 4596
rect 650 4591 651 4595
rect 655 4591 656 4595
rect 650 4590 656 4591
rect 914 4595 920 4596
rect 914 4591 915 4595
rect 919 4591 920 4595
rect 914 4590 920 4591
rect 1202 4595 1208 4596
rect 1202 4591 1203 4595
rect 1207 4591 1208 4595
rect 1202 4590 1208 4591
rect 1794 4595 1800 4596
rect 1794 4591 1795 4595
rect 1799 4591 1800 4595
rect 1794 4590 1800 4591
rect 2092 4590 2094 4597
rect 2167 4595 2168 4599
rect 2172 4598 2173 4599
rect 2338 4599 2344 4600
rect 2172 4596 2217 4598
rect 2172 4595 2173 4596
rect 2167 4594 2173 4595
rect 2338 4595 2339 4599
rect 2343 4598 2344 4599
rect 2882 4599 2888 4600
rect 2882 4598 2883 4599
rect 2343 4596 2449 4598
rect 2765 4596 2883 4598
rect 2343 4595 2344 4596
rect 2338 4594 2344 4595
rect 2882 4595 2883 4596
rect 2887 4595 2888 4599
rect 2882 4594 2888 4595
rect 2986 4599 2992 4600
rect 2986 4595 2987 4599
rect 2991 4595 2992 4599
rect 2986 4594 2992 4595
rect 3126 4599 3132 4600
rect 3126 4595 3127 4599
rect 3131 4595 3132 4599
rect 3126 4594 3132 4595
rect 3242 4599 3248 4600
rect 3242 4595 3243 4599
rect 3247 4598 3248 4599
rect 4159 4599 4160 4603
rect 4164 4602 4165 4603
rect 4170 4603 4176 4604
rect 4170 4602 4171 4603
rect 4164 4600 4171 4602
rect 4164 4599 4165 4600
rect 4159 4598 4165 4599
rect 4170 4599 4171 4600
rect 4175 4599 4176 4603
rect 4170 4598 4176 4599
rect 4295 4603 4301 4604
rect 4295 4599 4296 4603
rect 4300 4602 4301 4603
rect 4423 4603 4429 4604
rect 4423 4602 4424 4603
rect 4300 4600 4424 4602
rect 4300 4599 4301 4600
rect 4295 4598 4301 4599
rect 4423 4599 4424 4600
rect 4428 4599 4429 4603
rect 4423 4598 4429 4599
rect 4542 4603 4548 4604
rect 4542 4599 4543 4603
rect 4547 4602 4548 4603
rect 4695 4603 4701 4604
rect 4695 4602 4696 4603
rect 4547 4600 4696 4602
rect 4547 4599 4548 4600
rect 4542 4598 4548 4599
rect 4695 4599 4696 4600
rect 4700 4599 4701 4603
rect 4695 4598 4701 4599
rect 4858 4603 4864 4604
rect 4858 4599 4859 4603
rect 4863 4602 4864 4603
rect 4967 4603 4973 4604
rect 4967 4602 4968 4603
rect 4863 4600 4968 4602
rect 4863 4599 4864 4600
rect 4858 4598 4864 4599
rect 4967 4599 4968 4600
rect 4972 4599 4973 4603
rect 4967 4598 4973 4599
rect 5066 4603 5072 4604
rect 5066 4599 5067 4603
rect 5071 4602 5072 4603
rect 5247 4603 5253 4604
rect 5247 4602 5248 4603
rect 5071 4600 5248 4602
rect 5071 4599 5072 4600
rect 5066 4598 5072 4599
rect 5247 4599 5248 4600
rect 5252 4599 5253 4603
rect 5247 4598 5253 4599
rect 5534 4603 5541 4604
rect 5534 4599 5535 4603
rect 5540 4599 5541 4603
rect 5534 4598 5541 4599
rect 3247 4596 3345 4598
rect 3247 4595 3248 4596
rect 3242 4594 3248 4595
rect 2658 4591 2664 4592
rect 2658 4590 2659 4591
rect 2092 4588 2659 4590
rect 2658 4587 2659 4588
rect 2663 4587 2664 4591
rect 2658 4586 2664 4587
rect 2343 4563 2349 4564
rect 2343 4562 2344 4563
rect 2197 4560 2344 4562
rect 2343 4559 2344 4560
rect 2348 4559 2349 4563
rect 2567 4563 2573 4564
rect 2567 4562 2568 4563
rect 2445 4560 2568 4562
rect 2343 4558 2349 4559
rect 2567 4559 2568 4560
rect 2572 4559 2573 4563
rect 2567 4558 2573 4559
rect 2575 4563 2581 4564
rect 2575 4559 2576 4563
rect 2580 4562 2581 4563
rect 3399 4563 3405 4564
rect 3399 4562 3400 4563
rect 2580 4560 2585 4562
rect 3301 4560 3400 4562
rect 2580 4559 2581 4560
rect 2575 4558 2581 4559
rect 2890 4559 2896 4560
rect 295 4555 301 4556
rect 295 4551 296 4555
rect 300 4554 301 4555
rect 402 4555 408 4556
rect 402 4554 403 4555
rect 300 4552 403 4554
rect 300 4551 301 4552
rect 295 4550 301 4551
rect 402 4551 403 4552
rect 407 4551 408 4555
rect 402 4550 408 4551
rect 519 4555 525 4556
rect 519 4551 520 4555
rect 524 4554 525 4555
rect 650 4555 656 4556
rect 650 4554 651 4555
rect 524 4552 651 4554
rect 524 4551 525 4552
rect 519 4550 525 4551
rect 650 4551 651 4552
rect 655 4551 656 4555
rect 650 4550 656 4551
rect 767 4555 773 4556
rect 767 4551 768 4555
rect 772 4554 773 4555
rect 914 4555 920 4556
rect 914 4554 915 4555
rect 772 4552 915 4554
rect 772 4551 773 4552
rect 767 4550 773 4551
rect 914 4551 915 4552
rect 919 4551 920 4555
rect 914 4550 920 4551
rect 1031 4555 1037 4556
rect 1031 4551 1032 4555
rect 1036 4554 1037 4555
rect 1202 4555 1208 4556
rect 1202 4554 1203 4555
rect 1036 4552 1203 4554
rect 1036 4551 1037 4552
rect 1031 4550 1037 4551
rect 1202 4551 1203 4552
rect 1207 4551 1208 4555
rect 1202 4550 1208 4551
rect 1230 4555 1236 4556
rect 1230 4551 1231 4555
rect 1235 4554 1236 4555
rect 1319 4555 1325 4556
rect 1319 4554 1320 4555
rect 1235 4552 1320 4554
rect 1235 4551 1236 4552
rect 1230 4550 1236 4551
rect 1319 4551 1320 4552
rect 1324 4551 1325 4555
rect 1319 4550 1325 4551
rect 1518 4555 1524 4556
rect 1518 4551 1519 4555
rect 1523 4554 1524 4555
rect 1615 4555 1621 4556
rect 1615 4554 1616 4555
rect 1523 4552 1616 4554
rect 1523 4551 1524 4552
rect 1518 4550 1524 4551
rect 1615 4551 1616 4552
rect 1620 4551 1621 4555
rect 1615 4550 1621 4551
rect 1906 4555 1917 4556
rect 1906 4551 1907 4555
rect 1911 4551 1912 4555
rect 1916 4551 1917 4555
rect 2890 4555 2891 4559
rect 2895 4555 2896 4559
rect 2890 4554 2896 4555
rect 3010 4559 3016 4560
rect 3010 4555 3011 4559
rect 3015 4555 3016 4559
rect 3399 4559 3400 4560
rect 3404 4559 3405 4563
rect 3535 4563 3541 4564
rect 3535 4562 3536 4563
rect 3501 4560 3536 4562
rect 3399 4558 3405 4559
rect 3535 4559 3536 4560
rect 3540 4559 3541 4563
rect 4295 4563 4301 4564
rect 4295 4562 4296 4563
rect 4133 4560 4296 4562
rect 3535 4558 3541 4559
rect 3706 4559 3712 4560
rect 3010 4554 3016 4555
rect 3706 4555 3707 4559
rect 3711 4555 3712 4559
rect 4295 4559 4296 4560
rect 4300 4559 4301 4563
rect 4542 4563 4548 4564
rect 4542 4562 4543 4563
rect 4397 4560 4543 4562
rect 4295 4558 4301 4559
rect 4542 4559 4543 4560
rect 4547 4559 4548 4563
rect 4542 4558 4548 4559
rect 4590 4563 4596 4564
rect 4590 4559 4591 4563
rect 4595 4559 4596 4563
rect 5066 4563 5072 4564
rect 5066 4562 5067 4563
rect 4941 4560 5067 4562
rect 4590 4558 4596 4559
rect 5066 4559 5067 4560
rect 5071 4559 5072 4563
rect 5066 4558 5072 4559
rect 5218 4563 5224 4564
rect 5218 4559 5219 4563
rect 5223 4559 5224 4563
rect 5218 4558 5224 4559
rect 5494 4563 5500 4564
rect 5494 4559 5495 4563
rect 5499 4559 5500 4563
rect 5494 4558 5500 4559
rect 3706 4554 3712 4555
rect 1906 4550 1917 4551
rect 110 4548 116 4549
rect 1934 4548 1940 4549
rect 110 4544 111 4548
rect 115 4544 116 4548
rect 110 4543 116 4544
rect 170 4547 176 4548
rect 170 4543 171 4547
rect 175 4543 176 4547
rect 170 4542 176 4543
rect 394 4547 400 4548
rect 394 4543 395 4547
rect 399 4543 400 4547
rect 394 4542 400 4543
rect 642 4547 648 4548
rect 642 4543 643 4547
rect 647 4543 648 4547
rect 642 4542 648 4543
rect 906 4547 912 4548
rect 906 4543 907 4547
rect 911 4543 912 4547
rect 906 4542 912 4543
rect 1194 4547 1200 4548
rect 1194 4543 1195 4547
rect 1199 4543 1200 4547
rect 1194 4542 1200 4543
rect 1490 4547 1496 4548
rect 1490 4543 1491 4547
rect 1495 4543 1496 4547
rect 1490 4542 1496 4543
rect 1786 4547 1792 4548
rect 1786 4543 1787 4547
rect 1791 4543 1792 4547
rect 1934 4544 1935 4548
rect 1939 4544 1940 4548
rect 1934 4543 1940 4544
rect 1786 4542 1792 4543
rect 198 4532 204 4533
rect 110 4531 116 4532
rect 110 4527 111 4531
rect 115 4527 116 4531
rect 198 4528 199 4532
rect 203 4528 204 4532
rect 198 4527 204 4528
rect 422 4532 428 4533
rect 422 4528 423 4532
rect 427 4528 428 4532
rect 422 4527 428 4528
rect 670 4532 676 4533
rect 670 4528 671 4532
rect 675 4528 676 4532
rect 670 4527 676 4528
rect 934 4532 940 4533
rect 934 4528 935 4532
rect 939 4528 940 4532
rect 934 4527 940 4528
rect 1222 4532 1228 4533
rect 1222 4528 1223 4532
rect 1227 4528 1228 4532
rect 1222 4527 1228 4528
rect 1518 4532 1524 4533
rect 1518 4528 1519 4532
rect 1523 4528 1524 4532
rect 1518 4527 1524 4528
rect 1814 4532 1820 4533
rect 1814 4528 1815 4532
rect 1819 4528 1820 4532
rect 1814 4527 1820 4528
rect 1934 4531 1940 4532
rect 1934 4527 1935 4531
rect 1939 4527 1940 4531
rect 4170 4531 4176 4532
rect 110 4526 116 4527
rect 1934 4526 1940 4527
rect 2890 4527 2896 4528
rect 2890 4523 2891 4527
rect 2895 4526 2896 4527
rect 4170 4527 4171 4531
rect 4175 4530 4176 4531
rect 4974 4531 4980 4532
rect 4175 4528 4185 4530
rect 4175 4527 4176 4528
rect 4170 4526 4176 4527
rect 4418 4527 4424 4528
rect 2895 4524 3138 4526
rect 2895 4523 2896 4524
rect 2890 4522 2896 4523
rect 2222 4519 2229 4520
rect 2222 4515 2223 4519
rect 2228 4515 2229 4519
rect 2222 4514 2229 4515
rect 2343 4519 2349 4520
rect 2343 4515 2344 4519
rect 2348 4518 2349 4519
rect 2471 4519 2477 4520
rect 2471 4518 2472 4519
rect 2348 4516 2472 4518
rect 2348 4515 2349 4516
rect 2343 4514 2349 4515
rect 2471 4515 2472 4516
rect 2476 4515 2477 4519
rect 2471 4514 2477 4515
rect 2567 4519 2573 4520
rect 2567 4515 2568 4519
rect 2572 4518 2573 4519
rect 2703 4519 2709 4520
rect 2703 4518 2704 4519
rect 2572 4516 2704 4518
rect 2572 4515 2573 4516
rect 2567 4514 2573 4515
rect 2703 4515 2704 4516
rect 2708 4515 2709 4519
rect 2703 4514 2709 4515
rect 2919 4519 2925 4520
rect 2919 4515 2920 4519
rect 2924 4518 2925 4519
rect 3010 4519 3016 4520
rect 3010 4518 3011 4519
rect 2924 4516 3011 4518
rect 2924 4515 2925 4516
rect 2919 4514 2925 4515
rect 3010 4515 3011 4516
rect 3015 4515 3016 4519
rect 3010 4514 3016 4515
rect 3126 4519 3133 4520
rect 3126 4515 3127 4519
rect 3132 4515 3133 4519
rect 3136 4518 3138 4524
rect 4418 4523 4419 4527
rect 4423 4523 4424 4527
rect 4418 4522 4424 4523
rect 4666 4527 4672 4528
rect 4666 4523 4667 4527
rect 4671 4523 4672 4527
rect 4974 4527 4975 4531
rect 4979 4527 4980 4531
rect 5534 4531 5540 4532
rect 4974 4526 4980 4527
rect 5186 4527 5192 4528
rect 4666 4522 4672 4523
rect 5186 4523 5187 4527
rect 5191 4523 5192 4527
rect 5534 4527 5535 4531
rect 5539 4527 5540 4531
rect 5534 4526 5540 4527
rect 5186 4522 5192 4523
rect 3327 4519 3333 4520
rect 3327 4518 3328 4519
rect 3136 4516 3328 4518
rect 3126 4514 3133 4515
rect 3327 4515 3328 4516
rect 3332 4515 3333 4519
rect 3327 4514 3333 4515
rect 3399 4519 3405 4520
rect 3399 4515 3400 4519
rect 3404 4518 3405 4519
rect 3527 4519 3533 4520
rect 3527 4518 3528 4519
rect 3404 4516 3528 4518
rect 3404 4515 3405 4516
rect 3399 4514 3405 4515
rect 3527 4515 3528 4516
rect 3532 4515 3533 4519
rect 3527 4514 3533 4515
rect 3535 4519 3541 4520
rect 3535 4515 3536 4519
rect 3540 4518 3541 4519
rect 3735 4519 3741 4520
rect 3735 4518 3736 4519
rect 3540 4516 3736 4518
rect 3540 4515 3541 4516
rect 3535 4514 3541 4515
rect 3735 4515 3736 4516
rect 3740 4515 3741 4519
rect 3735 4514 3741 4515
rect 1974 4512 1980 4513
rect 3798 4512 3804 4513
rect 1974 4508 1975 4512
rect 1979 4508 1980 4512
rect 1974 4507 1980 4508
rect 2098 4511 2104 4512
rect 2098 4507 2099 4511
rect 2103 4507 2104 4511
rect 2098 4506 2104 4507
rect 2346 4511 2352 4512
rect 2346 4507 2347 4511
rect 2351 4507 2352 4511
rect 2346 4506 2352 4507
rect 2578 4511 2584 4512
rect 2578 4507 2579 4511
rect 2583 4507 2584 4511
rect 2578 4506 2584 4507
rect 2794 4511 2800 4512
rect 2794 4507 2795 4511
rect 2799 4507 2800 4511
rect 2794 4506 2800 4507
rect 3002 4511 3008 4512
rect 3002 4507 3003 4511
rect 3007 4507 3008 4511
rect 3002 4506 3008 4507
rect 3202 4511 3208 4512
rect 3202 4507 3203 4511
rect 3207 4507 3208 4511
rect 3202 4506 3208 4507
rect 3402 4511 3408 4512
rect 3402 4507 3403 4511
rect 3407 4507 3408 4511
rect 3402 4506 3408 4507
rect 3610 4511 3616 4512
rect 3610 4507 3611 4511
rect 3615 4507 3616 4511
rect 3798 4508 3799 4512
rect 3803 4508 3804 4512
rect 3798 4507 3804 4508
rect 3610 4506 3616 4507
rect 2126 4496 2132 4497
rect 1974 4495 1980 4496
rect 1974 4491 1975 4495
rect 1979 4491 1980 4495
rect 2126 4492 2127 4496
rect 2131 4492 2132 4496
rect 2126 4491 2132 4492
rect 2374 4496 2380 4497
rect 2374 4492 2375 4496
rect 2379 4492 2380 4496
rect 2374 4491 2380 4492
rect 2606 4496 2612 4497
rect 2606 4492 2607 4496
rect 2611 4492 2612 4496
rect 2606 4491 2612 4492
rect 2822 4496 2828 4497
rect 2822 4492 2823 4496
rect 2827 4492 2828 4496
rect 2822 4491 2828 4492
rect 3030 4496 3036 4497
rect 3030 4492 3031 4496
rect 3035 4492 3036 4496
rect 3030 4491 3036 4492
rect 3230 4496 3236 4497
rect 3230 4492 3231 4496
rect 3235 4492 3236 4496
rect 3230 4491 3236 4492
rect 3430 4496 3436 4497
rect 3430 4492 3431 4496
rect 3435 4492 3436 4496
rect 3430 4491 3436 4492
rect 3638 4496 3644 4497
rect 3638 4492 3639 4496
rect 3643 4492 3644 4496
rect 3638 4491 3644 4492
rect 3798 4495 3804 4496
rect 3798 4491 3799 4495
rect 3803 4491 3804 4495
rect 1974 4490 1980 4491
rect 3798 4490 3804 4491
rect 4303 4487 4309 4488
rect 4303 4483 4304 4487
rect 4308 4486 4309 4487
rect 4418 4487 4424 4488
rect 4418 4486 4419 4487
rect 4308 4484 4419 4486
rect 4308 4483 4309 4484
rect 4303 4482 4309 4483
rect 4418 4483 4419 4484
rect 4423 4483 4424 4487
rect 4418 4482 4424 4483
rect 4535 4487 4541 4488
rect 4535 4483 4536 4487
rect 4540 4486 4541 4487
rect 4666 4487 4672 4488
rect 4666 4486 4667 4487
rect 4540 4484 4667 4486
rect 4540 4483 4541 4484
rect 4535 4482 4541 4483
rect 4666 4483 4667 4484
rect 4671 4483 4672 4487
rect 4666 4482 4672 4483
rect 4754 4487 4760 4488
rect 4754 4483 4755 4487
rect 4759 4486 4760 4487
rect 4783 4487 4789 4488
rect 4783 4486 4784 4487
rect 4759 4484 4784 4486
rect 4759 4483 4760 4484
rect 4754 4482 4760 4483
rect 4783 4483 4784 4484
rect 4788 4483 4789 4487
rect 4783 4482 4789 4483
rect 5039 4487 5045 4488
rect 5039 4483 5040 4487
rect 5044 4486 5045 4487
rect 5186 4487 5192 4488
rect 5186 4486 5187 4487
rect 5044 4484 5187 4486
rect 5044 4483 5045 4484
rect 5039 4482 5045 4483
rect 5186 4483 5187 4484
rect 5191 4483 5192 4487
rect 5186 4482 5192 4483
rect 5218 4487 5224 4488
rect 5218 4483 5219 4487
rect 5223 4486 5224 4487
rect 5303 4487 5309 4488
rect 5303 4486 5304 4487
rect 5223 4484 5304 4486
rect 5223 4483 5224 4484
rect 5218 4482 5224 4483
rect 5303 4483 5304 4484
rect 5308 4483 5309 4487
rect 5303 4482 5309 4483
rect 5566 4487 5573 4488
rect 5566 4483 5567 4487
rect 5572 4483 5573 4487
rect 5566 4482 5573 4483
rect 3838 4480 3844 4481
rect 5662 4480 5668 4481
rect 3838 4476 3839 4480
rect 3843 4476 3844 4480
rect 3838 4475 3844 4476
rect 4178 4479 4184 4480
rect 4178 4475 4179 4479
rect 4183 4475 4184 4479
rect 4178 4474 4184 4475
rect 4410 4479 4416 4480
rect 4410 4475 4411 4479
rect 4415 4475 4416 4479
rect 4410 4474 4416 4475
rect 4658 4479 4664 4480
rect 4658 4475 4659 4479
rect 4663 4475 4664 4479
rect 4658 4474 4664 4475
rect 4914 4479 4920 4480
rect 4914 4475 4915 4479
rect 4919 4475 4920 4479
rect 4914 4474 4920 4475
rect 5178 4479 5184 4480
rect 5178 4475 5179 4479
rect 5183 4475 5184 4479
rect 5178 4474 5184 4475
rect 5442 4479 5448 4480
rect 5442 4475 5443 4479
rect 5447 4475 5448 4479
rect 5662 4476 5663 4480
rect 5667 4476 5668 4480
rect 5662 4475 5668 4476
rect 5442 4474 5448 4475
rect 110 4469 116 4470
rect 1934 4469 1940 4470
rect 110 4465 111 4469
rect 115 4465 116 4469
rect 110 4464 116 4465
rect 446 4468 452 4469
rect 446 4464 447 4468
rect 451 4464 452 4468
rect 446 4463 452 4464
rect 654 4468 660 4469
rect 654 4464 655 4468
rect 659 4464 660 4468
rect 654 4463 660 4464
rect 886 4468 892 4469
rect 886 4464 887 4468
rect 891 4464 892 4468
rect 886 4463 892 4464
rect 1142 4468 1148 4469
rect 1142 4464 1143 4468
rect 1147 4464 1148 4468
rect 1142 4463 1148 4464
rect 1406 4468 1412 4469
rect 1406 4464 1407 4468
rect 1411 4464 1412 4468
rect 1406 4463 1412 4464
rect 1678 4468 1684 4469
rect 1678 4464 1679 4468
rect 1683 4464 1684 4468
rect 1934 4465 1935 4469
rect 1939 4465 1940 4469
rect 1934 4464 1940 4465
rect 4206 4464 4212 4465
rect 1678 4463 1684 4464
rect 3838 4463 3844 4464
rect 3838 4459 3839 4463
rect 3843 4459 3844 4463
rect 4206 4460 4207 4464
rect 4211 4460 4212 4464
rect 4206 4459 4212 4460
rect 4438 4464 4444 4465
rect 4438 4460 4439 4464
rect 4443 4460 4444 4464
rect 4438 4459 4444 4460
rect 4686 4464 4692 4465
rect 4686 4460 4687 4464
rect 4691 4460 4692 4464
rect 4686 4459 4692 4460
rect 4942 4464 4948 4465
rect 4942 4460 4943 4464
rect 4947 4460 4948 4464
rect 4942 4459 4948 4460
rect 5206 4464 5212 4465
rect 5206 4460 5207 4464
rect 5211 4460 5212 4464
rect 5206 4459 5212 4460
rect 5470 4464 5476 4465
rect 5470 4460 5471 4464
rect 5475 4460 5476 4464
rect 5470 4459 5476 4460
rect 5662 4463 5668 4464
rect 5662 4459 5663 4463
rect 5667 4459 5668 4463
rect 3838 4458 3844 4459
rect 5662 4458 5668 4459
rect 418 4453 424 4454
rect 110 4452 116 4453
rect 110 4448 111 4452
rect 115 4448 116 4452
rect 418 4449 419 4453
rect 423 4449 424 4453
rect 418 4448 424 4449
rect 626 4453 632 4454
rect 626 4449 627 4453
rect 631 4449 632 4453
rect 626 4448 632 4449
rect 858 4453 864 4454
rect 858 4449 859 4453
rect 863 4449 864 4453
rect 858 4448 864 4449
rect 1114 4453 1120 4454
rect 1114 4449 1115 4453
rect 1119 4449 1120 4453
rect 1114 4448 1120 4449
rect 1378 4453 1384 4454
rect 1378 4449 1379 4453
rect 1383 4449 1384 4453
rect 1378 4448 1384 4449
rect 1650 4453 1656 4454
rect 1650 4449 1651 4453
rect 1655 4449 1656 4453
rect 1650 4448 1656 4449
rect 1934 4452 1940 4453
rect 1934 4448 1935 4452
rect 1939 4448 1940 4452
rect 110 4447 116 4448
rect 1934 4447 1940 4448
rect 543 4443 549 4444
rect 543 4439 544 4443
rect 548 4442 549 4443
rect 586 4443 592 4444
rect 586 4442 587 4443
rect 548 4440 587 4442
rect 548 4439 549 4440
rect 543 4438 549 4439
rect 586 4439 587 4440
rect 591 4439 592 4443
rect 586 4438 592 4439
rect 751 4443 760 4444
rect 751 4439 752 4443
rect 759 4439 760 4443
rect 751 4438 760 4439
rect 983 4443 989 4444
rect 983 4439 984 4443
rect 988 4442 989 4443
rect 1078 4443 1084 4444
rect 1078 4442 1079 4443
rect 988 4440 1079 4442
rect 988 4439 989 4440
rect 983 4438 989 4439
rect 1078 4439 1079 4440
rect 1083 4439 1084 4443
rect 1078 4438 1084 4439
rect 1239 4443 1248 4444
rect 1239 4439 1240 4443
rect 1247 4439 1248 4443
rect 1239 4438 1248 4439
rect 1274 4443 1280 4444
rect 1274 4439 1275 4443
rect 1279 4442 1280 4443
rect 1503 4443 1509 4444
rect 1503 4442 1504 4443
rect 1279 4440 1504 4442
rect 1279 4439 1280 4440
rect 1274 4438 1280 4439
rect 1503 4439 1504 4440
rect 1508 4439 1509 4443
rect 1503 4438 1509 4439
rect 1775 4443 1781 4444
rect 1775 4439 1776 4443
rect 1780 4442 1781 4443
rect 1794 4443 1800 4444
rect 1794 4442 1795 4443
rect 1780 4440 1795 4442
rect 1780 4439 1781 4440
rect 1775 4438 1781 4439
rect 1794 4439 1795 4440
rect 1799 4439 1800 4443
rect 1794 4438 1800 4439
rect 514 4435 520 4436
rect 514 4431 515 4435
rect 519 4434 520 4435
rect 1230 4435 1236 4436
rect 1230 4434 1231 4435
rect 519 4432 1231 4434
rect 519 4431 520 4432
rect 514 4430 520 4431
rect 1230 4431 1231 4432
rect 1235 4431 1236 4435
rect 1230 4430 1236 4431
rect 1974 4429 1980 4430
rect 3798 4429 3804 4430
rect 1974 4425 1975 4429
rect 1979 4425 1980 4429
rect 1974 4424 1980 4425
rect 2230 4428 2236 4429
rect 2230 4424 2231 4428
rect 2235 4424 2236 4428
rect 2230 4423 2236 4424
rect 2446 4428 2452 4429
rect 2446 4424 2447 4428
rect 2451 4424 2452 4428
rect 2446 4423 2452 4424
rect 2662 4428 2668 4429
rect 2662 4424 2663 4428
rect 2667 4424 2668 4428
rect 2662 4423 2668 4424
rect 2870 4428 2876 4429
rect 2870 4424 2871 4428
rect 2875 4424 2876 4428
rect 2870 4423 2876 4424
rect 3078 4428 3084 4429
rect 3078 4424 3079 4428
rect 3083 4424 3084 4428
rect 3078 4423 3084 4424
rect 3286 4428 3292 4429
rect 3286 4424 3287 4428
rect 3291 4424 3292 4428
rect 3286 4423 3292 4424
rect 3494 4428 3500 4429
rect 3494 4424 3495 4428
rect 3499 4424 3500 4428
rect 3494 4423 3500 4424
rect 3678 4428 3684 4429
rect 3678 4424 3679 4428
rect 3683 4424 3684 4428
rect 3798 4425 3799 4429
rect 3803 4425 3804 4429
rect 3798 4424 3804 4425
rect 3678 4423 3684 4424
rect 2202 4413 2208 4414
rect 1974 4412 1980 4413
rect 1974 4408 1975 4412
rect 1979 4408 1980 4412
rect 2202 4409 2203 4413
rect 2207 4409 2208 4413
rect 2202 4408 2208 4409
rect 2418 4413 2424 4414
rect 2418 4409 2419 4413
rect 2423 4409 2424 4413
rect 2418 4408 2424 4409
rect 2634 4413 2640 4414
rect 2634 4409 2635 4413
rect 2639 4409 2640 4413
rect 2634 4408 2640 4409
rect 2842 4413 2848 4414
rect 2842 4409 2843 4413
rect 2847 4409 2848 4413
rect 2842 4408 2848 4409
rect 3050 4413 3056 4414
rect 3050 4409 3051 4413
rect 3055 4409 3056 4413
rect 3050 4408 3056 4409
rect 3258 4413 3264 4414
rect 3258 4409 3259 4413
rect 3263 4409 3264 4413
rect 3258 4408 3264 4409
rect 3466 4413 3472 4414
rect 3466 4409 3467 4413
rect 3471 4409 3472 4413
rect 3466 4408 3472 4409
rect 3650 4413 3656 4414
rect 3650 4409 3651 4413
rect 3655 4409 3656 4413
rect 3650 4408 3656 4409
rect 3798 4412 3804 4413
rect 3798 4408 3799 4412
rect 3803 4408 3804 4412
rect 1974 4407 1980 4408
rect 3798 4407 3804 4408
rect 514 4403 520 4404
rect 514 4399 515 4403
rect 519 4399 520 4403
rect 514 4398 520 4399
rect 586 4403 592 4404
rect 586 4399 587 4403
rect 591 4402 592 4403
rect 754 4403 760 4404
rect 591 4400 633 4402
rect 591 4399 592 4400
rect 586 4398 592 4399
rect 754 4399 755 4403
rect 759 4402 760 4403
rect 1078 4403 1084 4404
rect 759 4400 865 4402
rect 759 4399 760 4400
rect 754 4398 760 4399
rect 1078 4399 1079 4403
rect 1083 4402 1084 4403
rect 1242 4403 1248 4404
rect 1083 4400 1121 4402
rect 1083 4399 1084 4400
rect 1078 4398 1084 4399
rect 1242 4399 1243 4403
rect 1247 4402 1248 4403
rect 1746 4403 1752 4404
rect 1247 4400 1385 4402
rect 1247 4399 1248 4400
rect 1242 4398 1248 4399
rect 1746 4399 1747 4403
rect 1751 4399 1752 4403
rect 1746 4398 1752 4399
rect 2327 4403 2336 4404
rect 2327 4399 2328 4403
rect 2335 4399 2336 4403
rect 2327 4398 2336 4399
rect 2543 4403 2552 4404
rect 2543 4399 2544 4403
rect 2551 4399 2552 4403
rect 2543 4398 2552 4399
rect 2759 4403 2765 4404
rect 2759 4399 2760 4403
rect 2764 4402 2765 4403
rect 2786 4403 2792 4404
rect 2786 4402 2787 4403
rect 2764 4400 2787 4402
rect 2764 4399 2765 4400
rect 2759 4398 2765 4399
rect 2786 4399 2787 4400
rect 2791 4399 2792 4403
rect 2786 4398 2792 4399
rect 2914 4403 2920 4404
rect 2914 4399 2915 4403
rect 2919 4402 2920 4403
rect 2967 4403 2973 4404
rect 2967 4402 2968 4403
rect 2919 4400 2968 4402
rect 2919 4399 2920 4400
rect 2914 4398 2920 4399
rect 2967 4399 2968 4400
rect 2972 4399 2973 4403
rect 2967 4398 2973 4399
rect 3175 4403 3181 4404
rect 3175 4399 3176 4403
rect 3180 4402 3181 4403
rect 3190 4403 3196 4404
rect 3190 4402 3191 4403
rect 3180 4400 3191 4402
rect 3180 4399 3181 4400
rect 3175 4398 3181 4399
rect 3190 4399 3191 4400
rect 3195 4399 3196 4403
rect 3190 4398 3196 4399
rect 3383 4403 3389 4404
rect 3383 4399 3384 4403
rect 3388 4402 3389 4403
rect 3430 4403 3436 4404
rect 3430 4402 3431 4403
rect 3388 4400 3431 4402
rect 3388 4399 3389 4400
rect 3383 4398 3389 4399
rect 3430 4399 3431 4400
rect 3435 4399 3436 4403
rect 3430 4398 3436 4399
rect 3591 4403 3597 4404
rect 3591 4399 3592 4403
rect 3596 4402 3597 4403
rect 3606 4403 3612 4404
rect 3606 4402 3607 4403
rect 3596 4400 3607 4402
rect 3596 4399 3597 4400
rect 3591 4398 3597 4399
rect 3606 4399 3607 4400
rect 3611 4399 3612 4403
rect 3606 4398 3612 4399
rect 3706 4403 3712 4404
rect 3706 4399 3707 4403
rect 3711 4402 3712 4403
rect 3775 4403 3781 4404
rect 3775 4402 3776 4403
rect 3711 4400 3776 4402
rect 3711 4399 3712 4400
rect 3706 4398 3712 4399
rect 3775 4399 3776 4400
rect 3780 4399 3781 4403
rect 3775 4398 3781 4399
rect 3838 4397 3844 4398
rect 5662 4397 5668 4398
rect 3838 4393 3839 4397
rect 3843 4393 3844 4397
rect 3838 4392 3844 4393
rect 4358 4396 4364 4397
rect 4358 4392 4359 4396
rect 4363 4392 4364 4396
rect 4358 4391 4364 4392
rect 4518 4396 4524 4397
rect 4518 4392 4519 4396
rect 4523 4392 4524 4396
rect 4518 4391 4524 4392
rect 4686 4396 4692 4397
rect 4686 4392 4687 4396
rect 4691 4392 4692 4396
rect 4686 4391 4692 4392
rect 4878 4396 4884 4397
rect 4878 4392 4879 4396
rect 4883 4392 4884 4396
rect 4878 4391 4884 4392
rect 5078 4396 5084 4397
rect 5078 4392 5079 4396
rect 5083 4392 5084 4396
rect 5078 4391 5084 4392
rect 5286 4396 5292 4397
rect 5286 4392 5287 4396
rect 5291 4392 5292 4396
rect 5286 4391 5292 4392
rect 5502 4396 5508 4397
rect 5502 4392 5503 4396
rect 5507 4392 5508 4396
rect 5662 4393 5663 4397
rect 5667 4393 5668 4397
rect 5662 4392 5668 4393
rect 5502 4391 5508 4392
rect 4330 4381 4336 4382
rect 3838 4380 3844 4381
rect 3838 4376 3839 4380
rect 3843 4376 3844 4380
rect 4330 4377 4331 4381
rect 4335 4377 4336 4381
rect 4330 4376 4336 4377
rect 4490 4381 4496 4382
rect 4490 4377 4491 4381
rect 4495 4377 4496 4381
rect 4490 4376 4496 4377
rect 4658 4381 4664 4382
rect 4658 4377 4659 4381
rect 4663 4377 4664 4381
rect 4658 4376 4664 4377
rect 4850 4381 4856 4382
rect 4850 4377 4851 4381
rect 4855 4377 4856 4381
rect 4850 4376 4856 4377
rect 5050 4381 5056 4382
rect 5050 4377 5051 4381
rect 5055 4377 5056 4381
rect 5050 4376 5056 4377
rect 5258 4381 5264 4382
rect 5258 4377 5259 4381
rect 5263 4377 5264 4381
rect 5258 4376 5264 4377
rect 5474 4381 5480 4382
rect 5474 4377 5475 4381
rect 5479 4377 5480 4381
rect 5474 4376 5480 4377
rect 5662 4380 5668 4381
rect 5662 4376 5663 4380
rect 5667 4376 5668 4380
rect 3838 4375 3844 4376
rect 5662 4375 5668 4376
rect 1274 4371 1280 4372
rect 1274 4370 1275 4371
rect 812 4368 1275 4370
rect 812 4366 814 4368
rect 1274 4367 1275 4368
rect 1279 4367 1280 4371
rect 1274 4366 1280 4367
rect 4346 4371 4352 4372
rect 4346 4367 4347 4371
rect 4351 4370 4352 4371
rect 4455 4371 4461 4372
rect 4455 4370 4456 4371
rect 4351 4368 4456 4370
rect 4351 4367 4352 4368
rect 4346 4366 4352 4367
rect 4455 4367 4456 4368
rect 4460 4367 4461 4371
rect 4455 4366 4461 4367
rect 4482 4371 4488 4372
rect 4482 4367 4483 4371
rect 4487 4370 4488 4371
rect 4615 4371 4621 4372
rect 4615 4370 4616 4371
rect 4487 4368 4616 4370
rect 4487 4367 4488 4368
rect 4482 4366 4488 4367
rect 4615 4367 4616 4368
rect 4620 4367 4621 4371
rect 4615 4366 4621 4367
rect 4647 4371 4653 4372
rect 4647 4367 4648 4371
rect 4652 4370 4653 4371
rect 4783 4371 4789 4372
rect 4783 4370 4784 4371
rect 4652 4368 4784 4370
rect 4652 4367 4653 4368
rect 4647 4366 4653 4367
rect 4783 4367 4784 4368
rect 4788 4367 4789 4371
rect 4783 4366 4789 4367
rect 4974 4371 4981 4372
rect 4974 4367 4975 4371
rect 4980 4367 4981 4371
rect 4974 4366 4981 4367
rect 5010 4371 5016 4372
rect 5010 4367 5011 4371
rect 5015 4370 5016 4371
rect 5175 4371 5181 4372
rect 5175 4370 5176 4371
rect 5015 4368 5176 4370
rect 5015 4367 5016 4368
rect 5010 4366 5016 4367
rect 5175 4367 5176 4368
rect 5180 4367 5181 4371
rect 5175 4366 5181 4367
rect 5223 4371 5229 4372
rect 5223 4367 5224 4371
rect 5228 4370 5229 4371
rect 5383 4371 5389 4372
rect 5383 4370 5384 4371
rect 5228 4368 5384 4370
rect 5228 4367 5229 4368
rect 5223 4366 5229 4367
rect 5383 4367 5384 4368
rect 5388 4367 5389 4371
rect 5383 4366 5389 4367
rect 5594 4371 5605 4372
rect 5594 4367 5595 4371
rect 5599 4367 5600 4371
rect 5604 4367 5605 4371
rect 5594 4366 5605 4367
rect 765 4364 814 4366
rect 818 4363 824 4364
rect 818 4359 819 4363
rect 823 4359 824 4363
rect 818 4358 824 4359
rect 970 4363 976 4364
rect 970 4359 971 4363
rect 975 4359 976 4363
rect 970 4358 976 4359
rect 1130 4363 1136 4364
rect 1130 4359 1131 4363
rect 1135 4359 1136 4363
rect 1130 4358 1136 4359
rect 1298 4363 1304 4364
rect 1298 4359 1299 4363
rect 1303 4359 1304 4363
rect 1298 4358 1304 4359
rect 1562 4363 1568 4364
rect 1562 4359 1563 4363
rect 1567 4359 1568 4363
rect 1562 4358 1568 4359
rect 1658 4363 1664 4364
rect 1658 4359 1659 4363
rect 1663 4359 1664 4363
rect 1658 4358 1664 4359
rect 2222 4363 2228 4364
rect 2222 4359 2223 4363
rect 2227 4359 2228 4363
rect 2222 4358 2228 4359
rect 2330 4363 2336 4364
rect 2330 4359 2331 4363
rect 2335 4362 2336 4363
rect 2546 4363 2552 4364
rect 2335 4360 2425 4362
rect 2335 4359 2336 4360
rect 2330 4358 2336 4359
rect 2546 4359 2547 4363
rect 2551 4362 2552 4363
rect 2786 4363 2792 4364
rect 2551 4360 2641 4362
rect 2551 4359 2552 4360
rect 2546 4358 2552 4359
rect 2786 4359 2787 4363
rect 2791 4362 2792 4363
rect 3190 4363 3196 4364
rect 2791 4360 2849 4362
rect 2791 4359 2792 4360
rect 2786 4358 2792 4359
rect 3148 4354 3150 4361
rect 3190 4359 3191 4363
rect 3195 4362 3196 4363
rect 3430 4363 3436 4364
rect 3195 4360 3265 4362
rect 3195 4359 3196 4360
rect 3190 4358 3196 4359
rect 3430 4359 3431 4363
rect 3435 4362 3436 4363
rect 3606 4363 3612 4364
rect 3435 4360 3473 4362
rect 3435 4359 3436 4360
rect 3430 4358 3436 4359
rect 3606 4359 3607 4363
rect 3611 4362 3612 4363
rect 3611 4360 3657 4362
rect 3611 4359 3612 4360
rect 3606 4358 3612 4359
rect 3438 4355 3444 4356
rect 3438 4354 3439 4355
rect 3148 4352 3439 4354
rect 3438 4351 3439 4352
rect 3443 4351 3444 4355
rect 3438 4350 3444 4351
rect 4482 4331 4488 4332
rect 4482 4330 4483 4331
rect 4429 4328 4483 4330
rect 2914 4327 2920 4328
rect 2914 4326 2915 4327
rect 2460 4324 2915 4326
rect 791 4323 797 4324
rect 791 4319 792 4323
rect 796 4322 797 4323
rect 818 4323 824 4324
rect 818 4322 819 4323
rect 796 4320 819 4322
rect 796 4319 797 4320
rect 791 4318 797 4319
rect 818 4319 819 4320
rect 823 4319 824 4323
rect 818 4318 824 4319
rect 935 4323 941 4324
rect 935 4319 936 4323
rect 940 4322 941 4323
rect 970 4323 976 4324
rect 970 4322 971 4323
rect 940 4320 971 4322
rect 940 4319 941 4320
rect 935 4318 941 4319
rect 970 4319 971 4320
rect 975 4319 976 4323
rect 970 4318 976 4319
rect 1087 4323 1093 4324
rect 1087 4319 1088 4323
rect 1092 4322 1093 4323
rect 1130 4323 1136 4324
rect 1130 4322 1131 4323
rect 1092 4320 1131 4322
rect 1092 4319 1093 4320
rect 1087 4318 1093 4319
rect 1130 4319 1131 4320
rect 1135 4319 1136 4323
rect 1130 4318 1136 4319
rect 1247 4323 1253 4324
rect 1247 4319 1248 4323
rect 1252 4322 1253 4323
rect 1298 4323 1304 4324
rect 1298 4322 1299 4323
rect 1252 4320 1299 4322
rect 1252 4319 1253 4320
rect 1247 4318 1253 4319
rect 1298 4319 1299 4320
rect 1303 4319 1304 4323
rect 1298 4318 1304 4319
rect 1306 4323 1312 4324
rect 1306 4319 1307 4323
rect 1311 4322 1312 4323
rect 1415 4323 1421 4324
rect 1415 4322 1416 4323
rect 1311 4320 1416 4322
rect 1311 4319 1312 4320
rect 1306 4318 1312 4319
rect 1415 4319 1416 4320
rect 1420 4319 1421 4323
rect 1415 4318 1421 4319
rect 1591 4323 1597 4324
rect 1591 4319 1592 4323
rect 1596 4322 1597 4323
rect 1658 4323 1664 4324
rect 1658 4322 1659 4323
rect 1596 4320 1659 4322
rect 1596 4319 1597 4320
rect 1591 4318 1597 4319
rect 1658 4319 1659 4320
rect 1663 4319 1664 4323
rect 1658 4318 1664 4319
rect 1746 4323 1752 4324
rect 1746 4319 1747 4323
rect 1751 4322 1752 4323
rect 1775 4323 1781 4324
rect 1775 4322 1776 4323
rect 1751 4320 1776 4322
rect 1751 4319 1752 4320
rect 1746 4318 1752 4319
rect 1775 4319 1776 4320
rect 1780 4319 1781 4323
rect 2460 4322 2462 4324
rect 2914 4323 2915 4324
rect 2919 4323 2920 4327
rect 4482 4327 4483 4328
rect 4487 4327 4488 4331
rect 4647 4331 4653 4332
rect 4647 4330 4648 4331
rect 4589 4328 4648 4330
rect 4482 4326 4488 4327
rect 4647 4327 4648 4328
rect 4652 4327 4653 4331
rect 4647 4326 4653 4327
rect 4754 4331 4760 4332
rect 4754 4327 4755 4331
rect 4759 4327 4760 4331
rect 5010 4331 5016 4332
rect 5010 4330 5011 4331
rect 4949 4328 5011 4330
rect 4754 4326 4760 4327
rect 5010 4327 5011 4328
rect 5015 4327 5016 4331
rect 5223 4331 5229 4332
rect 5223 4330 5224 4331
rect 5149 4328 5224 4330
rect 5010 4326 5016 4327
rect 5223 4327 5224 4328
rect 5228 4327 5229 4331
rect 5223 4326 5229 4327
rect 5354 4331 5360 4332
rect 5354 4327 5355 4331
rect 5359 4327 5360 4331
rect 5354 4326 5360 4327
rect 5566 4331 5572 4332
rect 5566 4327 5567 4331
rect 5571 4327 5572 4331
rect 5566 4326 5572 4327
rect 2914 4322 2920 4323
rect 3642 4323 3648 4324
rect 3642 4322 3643 4323
rect 2405 4320 2462 4322
rect 3549 4320 3643 4322
rect 1775 4318 1781 4319
rect 2466 4319 2472 4320
rect 110 4316 116 4317
rect 1934 4316 1940 4317
rect 110 4312 111 4316
rect 115 4312 116 4316
rect 110 4311 116 4312
rect 666 4315 672 4316
rect 666 4311 667 4315
rect 671 4311 672 4315
rect 666 4310 672 4311
rect 810 4315 816 4316
rect 810 4311 811 4315
rect 815 4311 816 4315
rect 810 4310 816 4311
rect 962 4315 968 4316
rect 962 4311 963 4315
rect 967 4311 968 4315
rect 962 4310 968 4311
rect 1122 4315 1128 4316
rect 1122 4311 1123 4315
rect 1127 4311 1128 4315
rect 1122 4310 1128 4311
rect 1290 4315 1296 4316
rect 1290 4311 1291 4315
rect 1295 4311 1296 4315
rect 1290 4310 1296 4311
rect 1466 4315 1472 4316
rect 1466 4311 1467 4315
rect 1471 4311 1472 4315
rect 1466 4310 1472 4311
rect 1650 4315 1656 4316
rect 1650 4311 1651 4315
rect 1655 4311 1656 4315
rect 1934 4312 1935 4316
rect 1939 4312 1940 4316
rect 2466 4315 2467 4319
rect 2471 4315 2472 4319
rect 2466 4314 2472 4315
rect 2634 4319 2640 4320
rect 2634 4315 2635 4319
rect 2639 4315 2640 4319
rect 2634 4314 2640 4315
rect 2818 4319 2824 4320
rect 2818 4315 2819 4319
rect 2823 4315 2824 4319
rect 2818 4314 2824 4315
rect 3018 4319 3024 4320
rect 3018 4315 3019 4319
rect 3023 4315 3024 4319
rect 3018 4314 3024 4315
rect 3234 4319 3240 4320
rect 3234 4315 3235 4319
rect 3239 4315 3240 4319
rect 3642 4319 3643 4320
rect 3647 4319 3648 4323
rect 3982 4323 3988 4324
rect 3982 4322 3983 4323
rect 3749 4320 3983 4322
rect 3642 4318 3648 4319
rect 3982 4319 3983 4320
rect 3987 4319 3988 4323
rect 3982 4318 3988 4319
rect 3234 4314 3240 4315
rect 1934 4311 1940 4312
rect 1650 4310 1656 4311
rect 694 4300 700 4301
rect 110 4299 116 4300
rect 110 4295 111 4299
rect 115 4295 116 4299
rect 694 4296 695 4300
rect 699 4296 700 4300
rect 694 4295 700 4296
rect 838 4300 844 4301
rect 838 4296 839 4300
rect 843 4296 844 4300
rect 838 4295 844 4296
rect 990 4300 996 4301
rect 990 4296 991 4300
rect 995 4296 996 4300
rect 990 4295 996 4296
rect 1150 4300 1156 4301
rect 1150 4296 1151 4300
rect 1155 4296 1156 4300
rect 1150 4295 1156 4296
rect 1318 4300 1324 4301
rect 1318 4296 1319 4300
rect 1323 4296 1324 4300
rect 1318 4295 1324 4296
rect 1494 4300 1500 4301
rect 1494 4296 1495 4300
rect 1499 4296 1500 4300
rect 1494 4295 1500 4296
rect 1678 4300 1684 4301
rect 1678 4296 1679 4300
rect 1683 4296 1684 4300
rect 1678 4295 1684 4296
rect 1934 4299 1940 4300
rect 1934 4295 1935 4299
rect 1939 4295 1940 4299
rect 4039 4299 4045 4300
rect 4039 4298 4040 4299
rect 3957 4296 4040 4298
rect 110 4294 116 4295
rect 1934 4294 1940 4295
rect 4039 4295 4040 4296
rect 4044 4295 4045 4299
rect 4346 4299 4352 4300
rect 4039 4294 4045 4295
rect 4050 4295 4056 4296
rect 4050 4291 4051 4295
rect 4055 4291 4056 4295
rect 4346 4295 4347 4299
rect 4351 4295 4352 4299
rect 5594 4299 5600 4300
rect 4346 4294 4352 4295
rect 4482 4295 4488 4296
rect 4050 4290 4056 4291
rect 4482 4291 4483 4295
rect 4487 4291 4488 4295
rect 4482 4290 4488 4291
rect 4722 4295 4728 4296
rect 4722 4291 4723 4295
rect 4727 4291 4728 4295
rect 4722 4290 4728 4291
rect 4978 4295 4984 4296
rect 4978 4291 4979 4295
rect 4983 4291 4984 4295
rect 4978 4290 4984 4291
rect 5242 4295 5248 4296
rect 5242 4291 5243 4295
rect 5247 4291 5248 4295
rect 5594 4295 5595 4299
rect 5599 4295 5600 4299
rect 5594 4294 5600 4295
rect 5242 4290 5248 4291
rect 2431 4279 2437 4280
rect 2431 4275 2432 4279
rect 2436 4278 2437 4279
rect 2466 4279 2472 4280
rect 2466 4278 2467 4279
rect 2436 4276 2467 4278
rect 2436 4275 2437 4276
rect 2431 4274 2437 4275
rect 2466 4275 2467 4276
rect 2471 4275 2472 4279
rect 2466 4274 2472 4275
rect 2583 4279 2589 4280
rect 2583 4275 2584 4279
rect 2588 4278 2589 4279
rect 2634 4279 2640 4280
rect 2634 4278 2635 4279
rect 2588 4276 2635 4278
rect 2588 4275 2589 4276
rect 2583 4274 2589 4275
rect 2634 4275 2635 4276
rect 2639 4275 2640 4279
rect 2634 4274 2640 4275
rect 2751 4279 2757 4280
rect 2751 4275 2752 4279
rect 2756 4278 2757 4279
rect 2818 4279 2824 4280
rect 2818 4278 2819 4279
rect 2756 4276 2819 4278
rect 2756 4275 2757 4276
rect 2751 4274 2757 4275
rect 2818 4275 2819 4276
rect 2823 4275 2824 4279
rect 2818 4274 2824 4275
rect 2935 4279 2941 4280
rect 2935 4275 2936 4279
rect 2940 4278 2941 4279
rect 3018 4279 3024 4280
rect 3018 4278 3019 4279
rect 2940 4276 3019 4278
rect 2940 4275 2941 4276
rect 2935 4274 2941 4275
rect 3018 4275 3019 4276
rect 3023 4275 3024 4279
rect 3018 4274 3024 4275
rect 3135 4279 3141 4280
rect 3135 4275 3136 4279
rect 3140 4278 3141 4279
rect 3234 4279 3240 4280
rect 3234 4278 3235 4279
rect 3140 4276 3235 4278
rect 3140 4275 3141 4276
rect 3135 4274 3141 4275
rect 3234 4275 3235 4276
rect 3239 4275 3240 4279
rect 3234 4274 3240 4275
rect 3350 4279 3357 4280
rect 3350 4275 3351 4279
rect 3356 4275 3357 4279
rect 3350 4274 3357 4275
rect 3438 4279 3444 4280
rect 3438 4275 3439 4279
rect 3443 4278 3444 4279
rect 3575 4279 3581 4280
rect 3575 4278 3576 4279
rect 3443 4276 3576 4278
rect 3443 4275 3444 4276
rect 3438 4274 3444 4275
rect 3575 4275 3576 4276
rect 3580 4275 3581 4279
rect 3575 4274 3581 4275
rect 3642 4279 3648 4280
rect 3642 4275 3643 4279
rect 3647 4278 3648 4279
rect 3775 4279 3781 4280
rect 3775 4278 3776 4279
rect 3647 4276 3776 4278
rect 3647 4275 3648 4276
rect 3642 4274 3648 4275
rect 3775 4275 3776 4276
rect 3780 4275 3781 4279
rect 3775 4274 3781 4275
rect 1974 4272 1980 4273
rect 3798 4272 3804 4273
rect 1974 4268 1975 4272
rect 1979 4268 1980 4272
rect 1974 4267 1980 4268
rect 2306 4271 2312 4272
rect 2306 4267 2307 4271
rect 2311 4267 2312 4271
rect 2306 4266 2312 4267
rect 2458 4271 2464 4272
rect 2458 4267 2459 4271
rect 2463 4267 2464 4271
rect 2458 4266 2464 4267
rect 2626 4271 2632 4272
rect 2626 4267 2627 4271
rect 2631 4267 2632 4271
rect 2626 4266 2632 4267
rect 2810 4271 2816 4272
rect 2810 4267 2811 4271
rect 2815 4267 2816 4271
rect 2810 4266 2816 4267
rect 3010 4271 3016 4272
rect 3010 4267 3011 4271
rect 3015 4267 3016 4271
rect 3010 4266 3016 4267
rect 3226 4271 3232 4272
rect 3226 4267 3227 4271
rect 3231 4267 3232 4271
rect 3226 4266 3232 4267
rect 3450 4271 3456 4272
rect 3450 4267 3451 4271
rect 3455 4267 3456 4271
rect 3450 4266 3456 4267
rect 3650 4271 3656 4272
rect 3650 4267 3651 4271
rect 3655 4267 3656 4271
rect 3798 4268 3799 4272
rect 3803 4268 3804 4272
rect 3798 4267 3804 4268
rect 3650 4266 3656 4267
rect 2334 4256 2340 4257
rect 1974 4255 1980 4256
rect 1974 4251 1975 4255
rect 1979 4251 1980 4255
rect 2334 4252 2335 4256
rect 2339 4252 2340 4256
rect 2334 4251 2340 4252
rect 2486 4256 2492 4257
rect 2486 4252 2487 4256
rect 2491 4252 2492 4256
rect 2486 4251 2492 4252
rect 2654 4256 2660 4257
rect 2654 4252 2655 4256
rect 2659 4252 2660 4256
rect 2654 4251 2660 4252
rect 2838 4256 2844 4257
rect 2838 4252 2839 4256
rect 2843 4252 2844 4256
rect 2838 4251 2844 4252
rect 3038 4256 3044 4257
rect 3038 4252 3039 4256
rect 3043 4252 3044 4256
rect 3038 4251 3044 4252
rect 3254 4256 3260 4257
rect 3254 4252 3255 4256
rect 3259 4252 3260 4256
rect 3254 4251 3260 4252
rect 3478 4256 3484 4257
rect 3478 4252 3479 4256
rect 3483 4252 3484 4256
rect 3478 4251 3484 4252
rect 3678 4256 3684 4257
rect 3678 4252 3679 4256
rect 3683 4252 3684 4256
rect 3678 4251 3684 4252
rect 3798 4255 3804 4256
rect 3798 4251 3799 4255
rect 3803 4251 3804 4255
rect 1974 4250 1980 4251
rect 3798 4250 3804 4251
rect 3982 4255 3989 4256
rect 3982 4251 3983 4255
rect 3988 4251 3989 4255
rect 3982 4250 3989 4251
rect 4039 4255 4045 4256
rect 4039 4251 4040 4255
rect 4044 4254 4045 4255
rect 4167 4255 4173 4256
rect 4167 4254 4168 4255
rect 4044 4252 4168 4254
rect 4044 4251 4045 4252
rect 4039 4250 4045 4251
rect 4167 4251 4168 4252
rect 4172 4251 4173 4255
rect 4167 4250 4173 4251
rect 4375 4255 4381 4256
rect 4375 4251 4376 4255
rect 4380 4254 4381 4255
rect 4482 4255 4488 4256
rect 4482 4254 4483 4255
rect 4380 4252 4483 4254
rect 4380 4251 4381 4252
rect 4375 4250 4381 4251
rect 4482 4251 4483 4252
rect 4487 4251 4488 4255
rect 4482 4250 4488 4251
rect 4599 4255 4605 4256
rect 4599 4251 4600 4255
rect 4604 4254 4605 4255
rect 4722 4255 4728 4256
rect 4722 4254 4723 4255
rect 4604 4252 4723 4254
rect 4604 4251 4605 4252
rect 4599 4250 4605 4251
rect 4722 4251 4723 4252
rect 4727 4251 4728 4255
rect 4722 4250 4728 4251
rect 4839 4255 4845 4256
rect 4839 4251 4840 4255
rect 4844 4254 4845 4255
rect 4978 4255 4984 4256
rect 4978 4254 4979 4255
rect 4844 4252 4979 4254
rect 4844 4251 4845 4252
rect 4839 4250 4845 4251
rect 4978 4251 4979 4252
rect 4983 4251 4984 4255
rect 4978 4250 4984 4251
rect 5095 4255 5101 4256
rect 5095 4251 5096 4255
rect 5100 4254 5101 4255
rect 5242 4255 5248 4256
rect 5242 4254 5243 4255
rect 5100 4252 5243 4254
rect 5100 4251 5101 4252
rect 5095 4250 5101 4251
rect 5242 4251 5243 4252
rect 5247 4251 5248 4255
rect 5242 4250 5248 4251
rect 5354 4255 5365 4256
rect 5354 4251 5355 4255
rect 5359 4251 5360 4255
rect 5364 4251 5365 4255
rect 5354 4250 5365 4251
rect 5610 4255 5616 4256
rect 5610 4251 5611 4255
rect 5615 4254 5616 4255
rect 5623 4255 5629 4256
rect 5623 4254 5624 4255
rect 5615 4252 5624 4254
rect 5615 4251 5616 4252
rect 5610 4250 5616 4251
rect 5623 4251 5624 4252
rect 5628 4251 5629 4255
rect 5623 4250 5629 4251
rect 3838 4248 3844 4249
rect 5662 4248 5668 4249
rect 3838 4244 3839 4248
rect 3843 4244 3844 4248
rect 3838 4243 3844 4244
rect 3858 4247 3864 4248
rect 3858 4243 3859 4247
rect 3863 4243 3864 4247
rect 3858 4242 3864 4243
rect 4042 4247 4048 4248
rect 4042 4243 4043 4247
rect 4047 4243 4048 4247
rect 4042 4242 4048 4243
rect 4250 4247 4256 4248
rect 4250 4243 4251 4247
rect 4255 4243 4256 4247
rect 4250 4242 4256 4243
rect 4474 4247 4480 4248
rect 4474 4243 4475 4247
rect 4479 4243 4480 4247
rect 4474 4242 4480 4243
rect 4714 4247 4720 4248
rect 4714 4243 4715 4247
rect 4719 4243 4720 4247
rect 4714 4242 4720 4243
rect 4970 4247 4976 4248
rect 4970 4243 4971 4247
rect 4975 4243 4976 4247
rect 4970 4242 4976 4243
rect 5234 4247 5240 4248
rect 5234 4243 5235 4247
rect 5239 4243 5240 4247
rect 5234 4242 5240 4243
rect 5498 4247 5504 4248
rect 5498 4243 5499 4247
rect 5503 4243 5504 4247
rect 5662 4244 5663 4248
rect 5667 4244 5668 4248
rect 5662 4243 5668 4244
rect 5498 4242 5504 4243
rect 3886 4232 3892 4233
rect 3838 4231 3844 4232
rect 3838 4227 3839 4231
rect 3843 4227 3844 4231
rect 3886 4228 3887 4232
rect 3891 4228 3892 4232
rect 3886 4227 3892 4228
rect 4070 4232 4076 4233
rect 4070 4228 4071 4232
rect 4075 4228 4076 4232
rect 4070 4227 4076 4228
rect 4278 4232 4284 4233
rect 4278 4228 4279 4232
rect 4283 4228 4284 4232
rect 4278 4227 4284 4228
rect 4502 4232 4508 4233
rect 4502 4228 4503 4232
rect 4507 4228 4508 4232
rect 4502 4227 4508 4228
rect 4742 4232 4748 4233
rect 4742 4228 4743 4232
rect 4747 4228 4748 4232
rect 4742 4227 4748 4228
rect 4998 4232 5004 4233
rect 4998 4228 4999 4232
rect 5003 4228 5004 4232
rect 4998 4227 5004 4228
rect 5262 4232 5268 4233
rect 5262 4228 5263 4232
rect 5267 4228 5268 4232
rect 5262 4227 5268 4228
rect 5526 4232 5532 4233
rect 5526 4228 5527 4232
rect 5531 4228 5532 4232
rect 5526 4227 5532 4228
rect 5662 4231 5668 4232
rect 5662 4227 5663 4231
rect 5667 4227 5668 4231
rect 3838 4226 3844 4227
rect 5662 4226 5668 4227
rect 110 4225 116 4226
rect 1934 4225 1940 4226
rect 110 4221 111 4225
rect 115 4221 116 4225
rect 110 4220 116 4221
rect 814 4224 820 4225
rect 814 4220 815 4224
rect 819 4220 820 4224
rect 814 4219 820 4220
rect 950 4224 956 4225
rect 950 4220 951 4224
rect 955 4220 956 4224
rect 950 4219 956 4220
rect 1086 4224 1092 4225
rect 1086 4220 1087 4224
rect 1091 4220 1092 4224
rect 1086 4219 1092 4220
rect 1222 4224 1228 4225
rect 1222 4220 1223 4224
rect 1227 4220 1228 4224
rect 1222 4219 1228 4220
rect 1358 4224 1364 4225
rect 1358 4220 1359 4224
rect 1363 4220 1364 4224
rect 1358 4219 1364 4220
rect 1494 4224 1500 4225
rect 1494 4220 1495 4224
rect 1499 4220 1500 4224
rect 1494 4219 1500 4220
rect 1630 4224 1636 4225
rect 1630 4220 1631 4224
rect 1635 4220 1636 4224
rect 1630 4219 1636 4220
rect 1766 4224 1772 4225
rect 1766 4220 1767 4224
rect 1771 4220 1772 4224
rect 1934 4221 1935 4225
rect 1939 4221 1940 4225
rect 1934 4220 1940 4221
rect 1766 4219 1772 4220
rect 786 4209 792 4210
rect 110 4208 116 4209
rect 110 4204 111 4208
rect 115 4204 116 4208
rect 786 4205 787 4209
rect 791 4205 792 4209
rect 786 4204 792 4205
rect 922 4209 928 4210
rect 922 4205 923 4209
rect 927 4205 928 4209
rect 922 4204 928 4205
rect 1058 4209 1064 4210
rect 1058 4205 1059 4209
rect 1063 4205 1064 4209
rect 1058 4204 1064 4205
rect 1194 4209 1200 4210
rect 1194 4205 1195 4209
rect 1199 4205 1200 4209
rect 1194 4204 1200 4205
rect 1330 4209 1336 4210
rect 1330 4205 1331 4209
rect 1335 4205 1336 4209
rect 1330 4204 1336 4205
rect 1466 4209 1472 4210
rect 1466 4205 1467 4209
rect 1471 4205 1472 4209
rect 1466 4204 1472 4205
rect 1602 4209 1608 4210
rect 1602 4205 1603 4209
rect 1607 4205 1608 4209
rect 1602 4204 1608 4205
rect 1738 4209 1744 4210
rect 1738 4205 1739 4209
rect 1743 4205 1744 4209
rect 1738 4204 1744 4205
rect 1934 4208 1940 4209
rect 1934 4204 1935 4208
rect 1939 4204 1940 4208
rect 110 4203 116 4204
rect 1934 4203 1940 4204
rect 911 4199 920 4200
rect 911 4195 912 4199
rect 919 4195 920 4199
rect 911 4194 920 4195
rect 1047 4199 1056 4200
rect 1047 4195 1048 4199
rect 1055 4195 1056 4199
rect 1047 4194 1056 4195
rect 1183 4199 1192 4200
rect 1183 4195 1184 4199
rect 1191 4195 1192 4199
rect 1183 4194 1192 4195
rect 1319 4199 1328 4200
rect 1319 4195 1320 4199
rect 1327 4195 1328 4199
rect 1319 4194 1328 4195
rect 1378 4199 1384 4200
rect 1378 4195 1379 4199
rect 1383 4198 1384 4199
rect 1455 4199 1461 4200
rect 1455 4198 1456 4199
rect 1383 4196 1456 4198
rect 1383 4195 1384 4196
rect 1378 4194 1384 4195
rect 1455 4195 1456 4196
rect 1460 4195 1461 4199
rect 1455 4194 1461 4195
rect 1562 4199 1568 4200
rect 1562 4195 1563 4199
rect 1567 4198 1568 4199
rect 1591 4199 1597 4200
rect 1591 4198 1592 4199
rect 1567 4196 1592 4198
rect 1567 4195 1568 4196
rect 1562 4194 1568 4195
rect 1591 4195 1592 4196
rect 1596 4195 1597 4199
rect 1591 4194 1597 4195
rect 1727 4199 1736 4200
rect 1727 4195 1728 4199
rect 1735 4195 1736 4199
rect 1863 4199 1869 4200
rect 1863 4198 1864 4199
rect 1727 4194 1736 4195
rect 1740 4196 1864 4198
rect 1562 4191 1568 4192
rect 1562 4187 1563 4191
rect 1567 4190 1568 4191
rect 1740 4190 1742 4196
rect 1863 4195 1864 4196
rect 1868 4195 1869 4199
rect 1863 4194 1869 4195
rect 1567 4188 1742 4190
rect 1974 4189 1980 4190
rect 3798 4189 3804 4190
rect 1567 4187 1568 4188
rect 1562 4186 1568 4187
rect 1974 4185 1975 4189
rect 1979 4185 1980 4189
rect 1974 4184 1980 4185
rect 2566 4188 2572 4189
rect 2566 4184 2567 4188
rect 2571 4184 2572 4188
rect 2566 4183 2572 4184
rect 2702 4188 2708 4189
rect 2702 4184 2703 4188
rect 2707 4184 2708 4188
rect 2702 4183 2708 4184
rect 2838 4188 2844 4189
rect 2838 4184 2839 4188
rect 2843 4184 2844 4188
rect 2838 4183 2844 4184
rect 2974 4188 2980 4189
rect 2974 4184 2975 4188
rect 2979 4184 2980 4188
rect 3798 4185 3799 4189
rect 3803 4185 3804 4189
rect 3798 4184 3804 4185
rect 2974 4183 2980 4184
rect 2538 4173 2544 4174
rect 1974 4172 1980 4173
rect 1974 4168 1975 4172
rect 1979 4168 1980 4172
rect 2538 4169 2539 4173
rect 2543 4169 2544 4173
rect 2538 4168 2544 4169
rect 2674 4173 2680 4174
rect 2674 4169 2675 4173
rect 2679 4169 2680 4173
rect 2674 4168 2680 4169
rect 2810 4173 2816 4174
rect 2810 4169 2811 4173
rect 2815 4169 2816 4173
rect 2810 4168 2816 4169
rect 2946 4173 2952 4174
rect 2946 4169 2947 4173
rect 2951 4169 2952 4173
rect 2946 4168 2952 4169
rect 3798 4172 3804 4173
rect 3798 4168 3799 4172
rect 3803 4168 3804 4172
rect 1974 4167 1980 4168
rect 3798 4167 3804 4168
rect 2658 4163 2669 4164
rect 914 4159 920 4160
rect 884 4150 886 4157
rect 914 4155 915 4159
rect 919 4158 920 4159
rect 1050 4159 1056 4160
rect 919 4156 929 4158
rect 919 4155 920 4156
rect 914 4154 920 4155
rect 1050 4155 1051 4159
rect 1055 4158 1056 4159
rect 1186 4159 1192 4160
rect 1055 4156 1065 4158
rect 1055 4155 1056 4156
rect 1050 4154 1056 4155
rect 1186 4155 1187 4159
rect 1191 4158 1192 4159
rect 1322 4159 1328 4160
rect 1191 4156 1201 4158
rect 1191 4155 1192 4156
rect 1186 4154 1192 4155
rect 1322 4155 1323 4159
rect 1327 4158 1328 4159
rect 1562 4159 1568 4160
rect 1327 4156 1337 4158
rect 1327 4155 1328 4156
rect 1322 4154 1328 4155
rect 1562 4155 1563 4159
rect 1567 4155 1568 4159
rect 1562 4154 1568 4155
rect 1670 4159 1676 4160
rect 1670 4155 1671 4159
rect 1675 4155 1676 4159
rect 1670 4154 1676 4155
rect 1730 4159 1736 4160
rect 1730 4155 1731 4159
rect 1735 4158 1736 4159
rect 2658 4159 2659 4163
rect 2663 4159 2664 4163
rect 2668 4159 2669 4163
rect 2658 4158 2669 4159
rect 2671 4163 2677 4164
rect 2671 4159 2672 4163
rect 2676 4162 2677 4163
rect 2799 4163 2805 4164
rect 2799 4162 2800 4163
rect 2676 4160 2800 4162
rect 2676 4159 2677 4160
rect 2671 4158 2677 4159
rect 2799 4159 2800 4160
rect 2804 4159 2805 4163
rect 2799 4158 2805 4159
rect 2807 4163 2813 4164
rect 2807 4159 2808 4163
rect 2812 4162 2813 4163
rect 2935 4163 2941 4164
rect 2935 4162 2936 4163
rect 2812 4160 2936 4162
rect 2812 4159 2813 4160
rect 2807 4158 2813 4159
rect 2935 4159 2936 4160
rect 2940 4159 2941 4163
rect 2935 4158 2941 4159
rect 2954 4163 2960 4164
rect 2954 4159 2955 4163
rect 2959 4162 2960 4163
rect 3071 4163 3077 4164
rect 3071 4162 3072 4163
rect 2959 4160 3072 4162
rect 2959 4159 2960 4160
rect 2954 4158 2960 4159
rect 3071 4159 3072 4160
rect 3076 4159 3077 4163
rect 3071 4158 3077 4159
rect 1735 4156 1745 4158
rect 1735 4155 1736 4156
rect 1730 4154 1736 4155
rect 1306 4151 1312 4152
rect 1306 4150 1307 4151
rect 884 4148 1307 4150
rect 1306 4147 1307 4148
rect 1311 4147 1312 4151
rect 1306 4146 1312 4147
rect 3838 4137 3844 4138
rect 5662 4137 5668 4138
rect 3838 4133 3839 4137
rect 3843 4133 3844 4137
rect 3838 4132 3844 4133
rect 3886 4136 3892 4137
rect 3886 4132 3887 4136
rect 3891 4132 3892 4136
rect 2954 4131 2960 4132
rect 3886 4131 3892 4132
rect 4414 4136 4420 4137
rect 4414 4132 4415 4136
rect 4419 4132 4420 4136
rect 4414 4131 4420 4132
rect 4974 4136 4980 4137
rect 4974 4132 4975 4136
rect 4979 4132 4980 4136
rect 4974 4131 4980 4132
rect 5542 4136 5548 4137
rect 5542 4132 5543 4136
rect 5547 4132 5548 4136
rect 5662 4133 5663 4137
rect 5667 4133 5668 4137
rect 5662 4132 5668 4133
rect 5542 4131 5548 4132
rect 2954 4130 2955 4131
rect 2908 4128 2955 4130
rect 1378 4127 1384 4128
rect 1378 4126 1379 4127
rect 1276 4124 1379 4126
rect 863 4123 869 4124
rect 863 4122 864 4123
rect 829 4120 864 4122
rect 863 4119 864 4120
rect 868 4119 869 4123
rect 999 4123 1005 4124
rect 999 4122 1000 4123
rect 965 4120 1000 4122
rect 863 4118 869 4119
rect 999 4119 1000 4120
rect 1004 4119 1005 4123
rect 1276 4122 1278 4124
rect 1378 4123 1379 4124
rect 1383 4123 1384 4127
rect 1378 4122 1384 4123
rect 2671 4123 2677 4124
rect 2671 4122 2672 4123
rect 1237 4120 1278 4122
rect 2637 4120 2672 4122
rect 999 4118 1005 4119
rect 1098 4119 1104 4120
rect 1098 4115 1099 4119
rect 1103 4115 1104 4119
rect 1098 4114 1104 4115
rect 1370 4119 1376 4120
rect 1370 4115 1371 4119
rect 1375 4115 1376 4119
rect 1370 4114 1376 4115
rect 1418 4119 1424 4120
rect 1418 4115 1419 4119
rect 1423 4115 1424 4119
rect 1418 4114 1424 4115
rect 1554 4119 1560 4120
rect 1554 4115 1555 4119
rect 1559 4115 1560 4119
rect 2671 4119 2672 4120
rect 2676 4119 2677 4123
rect 2807 4123 2813 4124
rect 2807 4122 2808 4123
rect 2773 4120 2808 4122
rect 2671 4118 2677 4119
rect 2807 4119 2808 4120
rect 2812 4119 2813 4123
rect 2908 4121 2910 4128
rect 2954 4127 2955 4128
rect 2959 4127 2960 4131
rect 2954 4126 2960 4127
rect 3350 4123 3356 4124
rect 3350 4122 3351 4123
rect 3045 4120 3351 4122
rect 2807 4118 2813 4119
rect 3350 4119 3351 4120
rect 3355 4119 3356 4123
rect 3858 4121 3864 4122
rect 3350 4118 3356 4119
rect 3838 4120 3844 4121
rect 3838 4116 3839 4120
rect 3843 4116 3844 4120
rect 3858 4117 3859 4121
rect 3863 4117 3864 4121
rect 3858 4116 3864 4117
rect 4386 4121 4392 4122
rect 4386 4117 4387 4121
rect 4391 4117 4392 4121
rect 4386 4116 4392 4117
rect 4946 4121 4952 4122
rect 4946 4117 4947 4121
rect 4951 4117 4952 4121
rect 4946 4116 4952 4117
rect 5514 4121 5520 4122
rect 5514 4117 5515 4121
rect 5519 4117 5520 4121
rect 5514 4116 5520 4117
rect 5662 4120 5668 4121
rect 5662 4116 5663 4120
rect 5667 4116 5668 4120
rect 3838 4115 3844 4116
rect 5662 4115 5668 4116
rect 1554 4114 1560 4115
rect 3983 4111 3989 4112
rect 3983 4107 3984 4111
rect 3988 4110 3989 4111
rect 4050 4111 4056 4112
rect 4050 4110 4051 4111
rect 3988 4108 4051 4110
rect 3988 4107 3989 4108
rect 3983 4106 3989 4107
rect 4050 4107 4051 4108
rect 4055 4107 4056 4111
rect 4050 4106 4056 4107
rect 4511 4111 4517 4112
rect 4511 4107 4512 4111
rect 4516 4110 4517 4111
rect 4878 4111 4884 4112
rect 4878 4110 4879 4111
rect 4516 4108 4879 4110
rect 4516 4107 4517 4108
rect 4511 4106 4517 4107
rect 4878 4107 4879 4108
rect 4883 4107 4884 4111
rect 5071 4111 5077 4112
rect 5071 4110 5072 4111
rect 4878 4106 4884 4107
rect 4888 4108 5072 4110
rect 3954 4103 3960 4104
rect 3954 4099 3955 4103
rect 3959 4102 3960 4103
rect 4888 4102 4890 4108
rect 5071 4107 5072 4108
rect 5076 4107 5077 4111
rect 5071 4106 5077 4107
rect 5618 4111 5624 4112
rect 5618 4107 5619 4111
rect 5623 4110 5624 4111
rect 5639 4111 5645 4112
rect 5639 4110 5640 4111
rect 5623 4108 5640 4110
rect 5623 4107 5624 4108
rect 5618 4106 5624 4107
rect 5639 4107 5640 4108
rect 5644 4107 5645 4111
rect 5639 4106 5645 4107
rect 3959 4100 4890 4102
rect 3959 4099 3960 4100
rect 3954 4098 3960 4099
rect 1098 4087 1104 4088
rect 1098 4083 1099 4087
rect 1103 4086 1104 4087
rect 1103 4084 1186 4086
rect 1103 4083 1104 4084
rect 1098 4082 1104 4083
rect 854 4079 861 4080
rect 854 4075 855 4079
rect 860 4075 861 4079
rect 854 4074 861 4075
rect 863 4079 869 4080
rect 863 4075 864 4079
rect 868 4078 869 4079
rect 991 4079 997 4080
rect 991 4078 992 4079
rect 868 4076 992 4078
rect 868 4075 869 4076
rect 863 4074 869 4075
rect 991 4075 992 4076
rect 996 4075 997 4079
rect 991 4074 997 4075
rect 999 4079 1005 4080
rect 999 4075 1000 4079
rect 1004 4078 1005 4079
rect 1127 4079 1133 4080
rect 1127 4078 1128 4079
rect 1004 4076 1128 4078
rect 1004 4075 1005 4076
rect 999 4074 1005 4075
rect 1127 4075 1128 4076
rect 1132 4075 1133 4079
rect 1184 4078 1186 4084
rect 1263 4079 1269 4080
rect 1263 4078 1264 4079
rect 1184 4076 1264 4078
rect 1127 4074 1133 4075
rect 1263 4075 1264 4076
rect 1268 4075 1269 4079
rect 1263 4074 1269 4075
rect 1399 4079 1405 4080
rect 1399 4075 1400 4079
rect 1404 4078 1405 4079
rect 1418 4079 1424 4080
rect 1418 4078 1419 4079
rect 1404 4076 1419 4078
rect 1404 4075 1405 4076
rect 1399 4074 1405 4075
rect 1418 4075 1419 4076
rect 1423 4075 1424 4079
rect 1418 4074 1424 4075
rect 1535 4079 1541 4080
rect 1535 4075 1536 4079
rect 1540 4078 1541 4079
rect 1554 4079 1560 4080
rect 1554 4078 1555 4079
rect 1540 4076 1555 4078
rect 1540 4075 1541 4076
rect 1535 4074 1541 4075
rect 1554 4075 1555 4076
rect 1559 4075 1560 4079
rect 1554 4074 1560 4075
rect 1670 4079 1677 4080
rect 1670 4075 1671 4079
rect 1676 4075 1677 4079
rect 1670 4074 1677 4075
rect 110 4072 116 4073
rect 1934 4072 1940 4073
rect 110 4068 111 4072
rect 115 4068 116 4072
rect 110 4067 116 4068
rect 730 4071 736 4072
rect 730 4067 731 4071
rect 735 4067 736 4071
rect 730 4066 736 4067
rect 866 4071 872 4072
rect 866 4067 867 4071
rect 871 4067 872 4071
rect 866 4066 872 4067
rect 1002 4071 1008 4072
rect 1002 4067 1003 4071
rect 1007 4067 1008 4071
rect 1002 4066 1008 4067
rect 1138 4071 1144 4072
rect 1138 4067 1139 4071
rect 1143 4067 1144 4071
rect 1138 4066 1144 4067
rect 1274 4071 1280 4072
rect 1274 4067 1275 4071
rect 1279 4067 1280 4071
rect 1274 4066 1280 4067
rect 1410 4071 1416 4072
rect 1410 4067 1411 4071
rect 1415 4067 1416 4071
rect 1410 4066 1416 4067
rect 1546 4071 1552 4072
rect 1546 4067 1547 4071
rect 1551 4067 1552 4071
rect 1934 4068 1935 4072
rect 1939 4068 1940 4072
rect 2658 4071 2664 4072
rect 1934 4067 1940 4068
rect 2386 4067 2392 4068
rect 1546 4066 1552 4067
rect 2386 4063 2387 4067
rect 2391 4063 2392 4067
rect 2386 4062 2392 4063
rect 2434 4067 2440 4068
rect 2434 4063 2435 4067
rect 2439 4063 2440 4067
rect 2658 4067 2659 4071
rect 2663 4067 2664 4071
rect 3954 4071 3960 4072
rect 2658 4066 2664 4067
rect 2706 4067 2712 4068
rect 2434 4062 2440 4063
rect 2706 4063 2707 4067
rect 2711 4063 2712 4067
rect 2706 4062 2712 4063
rect 2842 4067 2848 4068
rect 2842 4063 2843 4067
rect 2847 4063 2848 4067
rect 3954 4067 3955 4071
rect 3959 4067 3960 4071
rect 3954 4066 3960 4067
rect 4303 4071 4309 4072
rect 4303 4067 4304 4071
rect 4308 4070 4309 4071
rect 4878 4071 4884 4072
rect 4308 4068 4393 4070
rect 4308 4067 4309 4068
rect 4303 4066 4309 4067
rect 4878 4067 4879 4071
rect 4883 4070 4884 4071
rect 5610 4071 5616 4072
rect 4883 4068 4953 4070
rect 4883 4067 4884 4068
rect 4878 4066 4884 4067
rect 5610 4067 5611 4071
rect 5615 4067 5616 4071
rect 5610 4066 5616 4067
rect 2842 4062 2848 4063
rect 758 4056 764 4057
rect 110 4055 116 4056
rect 110 4051 111 4055
rect 115 4051 116 4055
rect 758 4052 759 4056
rect 763 4052 764 4056
rect 758 4051 764 4052
rect 894 4056 900 4057
rect 894 4052 895 4056
rect 899 4052 900 4056
rect 894 4051 900 4052
rect 1030 4056 1036 4057
rect 1030 4052 1031 4056
rect 1035 4052 1036 4056
rect 1030 4051 1036 4052
rect 1166 4056 1172 4057
rect 1166 4052 1167 4056
rect 1171 4052 1172 4056
rect 1166 4051 1172 4052
rect 1302 4056 1308 4057
rect 1302 4052 1303 4056
rect 1307 4052 1308 4056
rect 1302 4051 1308 4052
rect 1438 4056 1444 4057
rect 1438 4052 1439 4056
rect 1443 4052 1444 4056
rect 1438 4051 1444 4052
rect 1574 4056 1580 4057
rect 1574 4052 1575 4056
rect 1579 4052 1580 4056
rect 1574 4051 1580 4052
rect 1934 4055 1940 4056
rect 1934 4051 1935 4055
rect 1939 4051 1940 4055
rect 110 4050 116 4051
rect 1934 4050 1940 4051
rect 4495 4039 4501 4040
rect 4495 4038 4496 4039
rect 4437 4036 4496 4038
rect 3866 4035 3872 4036
rect 3866 4031 3867 4035
rect 3871 4031 3872 4035
rect 3866 4030 3872 4031
rect 4010 4035 4016 4036
rect 4010 4031 4011 4035
rect 4015 4031 4016 4035
rect 4010 4030 4016 4031
rect 4178 4035 4184 4036
rect 4178 4031 4179 4035
rect 4183 4031 4184 4035
rect 4495 4035 4496 4036
rect 4500 4035 4501 4039
rect 4647 4039 4653 4040
rect 4647 4038 4648 4039
rect 4597 4036 4648 4038
rect 4495 4034 4501 4035
rect 4647 4035 4648 4036
rect 4652 4035 4653 4039
rect 4799 4039 4805 4040
rect 4799 4038 4800 4039
rect 4749 4036 4800 4038
rect 4647 4034 4653 4035
rect 4799 4035 4800 4036
rect 4804 4035 4805 4039
rect 4943 4039 4949 4040
rect 4943 4038 4944 4039
rect 4901 4036 4944 4038
rect 4799 4034 4805 4035
rect 4943 4035 4944 4036
rect 4948 4035 4949 4039
rect 5087 4039 5093 4040
rect 5087 4038 5088 4039
rect 5045 4036 5088 4038
rect 4943 4034 4949 4035
rect 5087 4035 5088 4036
rect 5092 4035 5093 4039
rect 5223 4039 5229 4040
rect 5223 4038 5224 4039
rect 5189 4036 5224 4038
rect 5087 4034 5093 4035
rect 5223 4035 5224 4036
rect 5228 4035 5229 4039
rect 5375 4039 5381 4040
rect 5375 4038 5376 4039
rect 5333 4036 5376 4038
rect 5223 4034 5229 4035
rect 5375 4035 5376 4036
rect 5380 4035 5381 4039
rect 5375 4034 5381 4035
rect 5398 4039 5404 4040
rect 5398 4035 5399 4039
rect 5403 4035 5404 4039
rect 5618 4039 5624 4040
rect 5618 4038 5619 4039
rect 5613 4036 5619 4038
rect 5398 4034 5404 4035
rect 5618 4035 5619 4036
rect 5623 4035 5624 4039
rect 5618 4034 5624 4035
rect 4178 4030 4184 4031
rect 2415 4027 2421 4028
rect 2415 4023 2416 4027
rect 2420 4026 2421 4027
rect 2434 4027 2440 4028
rect 2434 4026 2435 4027
rect 2420 4024 2435 4026
rect 2420 4023 2421 4024
rect 2415 4022 2421 4023
rect 2434 4023 2435 4024
rect 2439 4023 2440 4027
rect 2434 4022 2440 4023
rect 2550 4027 2557 4028
rect 2550 4023 2551 4027
rect 2556 4023 2557 4027
rect 2550 4022 2557 4023
rect 2687 4027 2693 4028
rect 2687 4023 2688 4027
rect 2692 4026 2693 4027
rect 2706 4027 2712 4028
rect 2706 4026 2707 4027
rect 2692 4024 2707 4026
rect 2692 4023 2693 4024
rect 2687 4022 2693 4023
rect 2706 4023 2707 4024
rect 2711 4023 2712 4027
rect 2706 4022 2712 4023
rect 2823 4027 2829 4028
rect 2823 4023 2824 4027
rect 2828 4026 2829 4027
rect 2842 4027 2848 4028
rect 2842 4026 2843 4027
rect 2828 4024 2843 4026
rect 2828 4023 2829 4024
rect 2823 4022 2829 4023
rect 2842 4023 2843 4024
rect 2847 4023 2848 4027
rect 2842 4022 2848 4023
rect 2958 4027 2965 4028
rect 2958 4023 2959 4027
rect 2964 4023 2965 4027
rect 2958 4022 2965 4023
rect 1974 4020 1980 4021
rect 3798 4020 3804 4021
rect 1974 4016 1975 4020
rect 1979 4016 1980 4020
rect 1974 4015 1980 4016
rect 2290 4019 2296 4020
rect 2290 4015 2291 4019
rect 2295 4015 2296 4019
rect 2290 4014 2296 4015
rect 2426 4019 2432 4020
rect 2426 4015 2427 4019
rect 2431 4015 2432 4019
rect 2426 4014 2432 4015
rect 2562 4019 2568 4020
rect 2562 4015 2563 4019
rect 2567 4015 2568 4019
rect 2562 4014 2568 4015
rect 2698 4019 2704 4020
rect 2698 4015 2699 4019
rect 2703 4015 2704 4019
rect 2698 4014 2704 4015
rect 2834 4019 2840 4020
rect 2834 4015 2835 4019
rect 2839 4015 2840 4019
rect 3798 4016 3799 4020
rect 3803 4016 3804 4020
rect 3798 4015 3804 4016
rect 2834 4014 2840 4015
rect 2318 4004 2324 4005
rect 1974 4003 1980 4004
rect 1974 3999 1975 4003
rect 1979 3999 1980 4003
rect 2318 4000 2319 4004
rect 2323 4000 2324 4004
rect 2318 3999 2324 4000
rect 2454 4004 2460 4005
rect 2454 4000 2455 4004
rect 2459 4000 2460 4004
rect 2454 3999 2460 4000
rect 2590 4004 2596 4005
rect 2590 4000 2591 4004
rect 2595 4000 2596 4004
rect 2590 3999 2596 4000
rect 2726 4004 2732 4005
rect 2726 4000 2727 4004
rect 2731 4000 2732 4004
rect 2726 3999 2732 4000
rect 2862 4004 2868 4005
rect 2862 4000 2863 4004
rect 2867 4000 2868 4004
rect 2862 3999 2868 4000
rect 3798 4003 3804 4004
rect 3798 3999 3799 4003
rect 3803 3999 3804 4003
rect 1974 3998 1980 3999
rect 3798 3998 3804 3999
rect 3983 3995 3989 3996
rect 3983 3991 3984 3995
rect 3988 3994 3989 3995
rect 4010 3995 4016 3996
rect 4010 3994 4011 3995
rect 3988 3992 4011 3994
rect 3988 3991 3989 3992
rect 3983 3990 3989 3991
rect 4010 3991 4011 3992
rect 4015 3991 4016 3995
rect 4010 3990 4016 3991
rect 4127 3995 4133 3996
rect 4127 3991 4128 3995
rect 4132 3994 4133 3995
rect 4178 3995 4184 3996
rect 4178 3994 4179 3995
rect 4132 3992 4179 3994
rect 4132 3991 4133 3992
rect 4127 3990 4133 3991
rect 4178 3991 4179 3992
rect 4183 3991 4184 3995
rect 4178 3990 4184 3991
rect 4295 3995 4301 3996
rect 4295 3991 4296 3995
rect 4300 3994 4301 3995
rect 4303 3995 4309 3996
rect 4303 3994 4304 3995
rect 4300 3992 4304 3994
rect 4300 3991 4301 3992
rect 4295 3990 4301 3991
rect 4303 3991 4304 3992
rect 4308 3991 4309 3995
rect 4303 3990 4309 3991
rect 4450 3995 4456 3996
rect 4450 3991 4451 3995
rect 4455 3994 4456 3995
rect 4463 3995 4469 3996
rect 4463 3994 4464 3995
rect 4455 3992 4464 3994
rect 4455 3991 4456 3992
rect 4450 3990 4456 3991
rect 4463 3991 4464 3992
rect 4468 3991 4469 3995
rect 4463 3990 4469 3991
rect 4495 3995 4501 3996
rect 4495 3991 4496 3995
rect 4500 3994 4501 3995
rect 4623 3995 4629 3996
rect 4623 3994 4624 3995
rect 4500 3992 4624 3994
rect 4500 3991 4501 3992
rect 4495 3990 4501 3991
rect 4623 3991 4624 3992
rect 4628 3991 4629 3995
rect 4623 3990 4629 3991
rect 4647 3995 4653 3996
rect 4647 3991 4648 3995
rect 4652 3994 4653 3995
rect 4775 3995 4781 3996
rect 4775 3994 4776 3995
rect 4652 3992 4776 3994
rect 4652 3991 4653 3992
rect 4647 3990 4653 3991
rect 4775 3991 4776 3992
rect 4780 3991 4781 3995
rect 4775 3990 4781 3991
rect 4799 3995 4805 3996
rect 4799 3991 4800 3995
rect 4804 3994 4805 3995
rect 4927 3995 4933 3996
rect 4927 3994 4928 3995
rect 4804 3992 4928 3994
rect 4804 3991 4805 3992
rect 4799 3990 4805 3991
rect 4927 3991 4928 3992
rect 4932 3991 4933 3995
rect 4927 3990 4933 3991
rect 4943 3995 4949 3996
rect 4943 3991 4944 3995
rect 4948 3994 4949 3995
rect 5071 3995 5077 3996
rect 5071 3994 5072 3995
rect 4948 3992 5072 3994
rect 4948 3991 4949 3992
rect 4943 3990 4949 3991
rect 5071 3991 5072 3992
rect 5076 3991 5077 3995
rect 5071 3990 5077 3991
rect 5087 3995 5093 3996
rect 5087 3991 5088 3995
rect 5092 3994 5093 3995
rect 5215 3995 5221 3996
rect 5215 3994 5216 3995
rect 5092 3992 5216 3994
rect 5092 3991 5093 3992
rect 5087 3990 5093 3991
rect 5215 3991 5216 3992
rect 5220 3991 5221 3995
rect 5215 3990 5221 3991
rect 5223 3995 5229 3996
rect 5223 3991 5224 3995
rect 5228 3994 5229 3995
rect 5359 3995 5365 3996
rect 5359 3994 5360 3995
rect 5228 3992 5360 3994
rect 5228 3991 5229 3992
rect 5223 3990 5229 3991
rect 5359 3991 5360 3992
rect 5364 3991 5365 3995
rect 5359 3990 5365 3991
rect 5375 3995 5381 3996
rect 5375 3991 5376 3995
rect 5380 3994 5381 3995
rect 5503 3995 5509 3996
rect 5503 3994 5504 3995
rect 5380 3992 5504 3994
rect 5380 3991 5381 3992
rect 5375 3990 5381 3991
rect 5503 3991 5504 3992
rect 5508 3991 5509 3995
rect 5503 3990 5509 3991
rect 5634 3995 5645 3996
rect 5634 3991 5635 3995
rect 5639 3991 5640 3995
rect 5644 3991 5645 3995
rect 5634 3990 5645 3991
rect 3838 3988 3844 3989
rect 5662 3988 5668 3989
rect 3838 3984 3839 3988
rect 3843 3984 3844 3988
rect 3838 3983 3844 3984
rect 3858 3987 3864 3988
rect 3858 3983 3859 3987
rect 3863 3983 3864 3987
rect 3858 3982 3864 3983
rect 4002 3987 4008 3988
rect 4002 3983 4003 3987
rect 4007 3983 4008 3987
rect 4002 3982 4008 3983
rect 4170 3987 4176 3988
rect 4170 3983 4171 3987
rect 4175 3983 4176 3987
rect 4170 3982 4176 3983
rect 4338 3987 4344 3988
rect 4338 3983 4339 3987
rect 4343 3983 4344 3987
rect 4338 3982 4344 3983
rect 4498 3987 4504 3988
rect 4498 3983 4499 3987
rect 4503 3983 4504 3987
rect 4498 3982 4504 3983
rect 4650 3987 4656 3988
rect 4650 3983 4651 3987
rect 4655 3983 4656 3987
rect 4650 3982 4656 3983
rect 4802 3987 4808 3988
rect 4802 3983 4803 3987
rect 4807 3983 4808 3987
rect 4802 3982 4808 3983
rect 4946 3987 4952 3988
rect 4946 3983 4947 3987
rect 4951 3983 4952 3987
rect 4946 3982 4952 3983
rect 5090 3987 5096 3988
rect 5090 3983 5091 3987
rect 5095 3983 5096 3987
rect 5090 3982 5096 3983
rect 5234 3987 5240 3988
rect 5234 3983 5235 3987
rect 5239 3983 5240 3987
rect 5234 3982 5240 3983
rect 5378 3987 5384 3988
rect 5378 3983 5379 3987
rect 5383 3983 5384 3987
rect 5378 3982 5384 3983
rect 5514 3987 5520 3988
rect 5514 3983 5515 3987
rect 5519 3983 5520 3987
rect 5662 3984 5663 3988
rect 5667 3984 5668 3988
rect 5662 3983 5668 3984
rect 5514 3982 5520 3983
rect 110 3973 116 3974
rect 1934 3973 1940 3974
rect 110 3969 111 3973
rect 115 3969 116 3973
rect 110 3968 116 3969
rect 510 3972 516 3973
rect 510 3968 511 3972
rect 515 3968 516 3972
rect 510 3967 516 3968
rect 662 3972 668 3973
rect 662 3968 663 3972
rect 667 3968 668 3972
rect 662 3967 668 3968
rect 822 3972 828 3973
rect 822 3968 823 3972
rect 827 3968 828 3972
rect 822 3967 828 3968
rect 982 3972 988 3973
rect 982 3968 983 3972
rect 987 3968 988 3972
rect 982 3967 988 3968
rect 1150 3972 1156 3973
rect 1150 3968 1151 3972
rect 1155 3968 1156 3972
rect 1150 3967 1156 3968
rect 1318 3972 1324 3973
rect 1318 3968 1319 3972
rect 1323 3968 1324 3972
rect 1934 3969 1935 3973
rect 1939 3969 1940 3973
rect 3886 3972 3892 3973
rect 1934 3968 1940 3969
rect 3838 3971 3844 3972
rect 1318 3967 1324 3968
rect 3838 3967 3839 3971
rect 3843 3967 3844 3971
rect 3886 3968 3887 3972
rect 3891 3968 3892 3972
rect 3886 3967 3892 3968
rect 4030 3972 4036 3973
rect 4030 3968 4031 3972
rect 4035 3968 4036 3972
rect 4030 3967 4036 3968
rect 4198 3972 4204 3973
rect 4198 3968 4199 3972
rect 4203 3968 4204 3972
rect 4198 3967 4204 3968
rect 4366 3972 4372 3973
rect 4366 3968 4367 3972
rect 4371 3968 4372 3972
rect 4366 3967 4372 3968
rect 4526 3972 4532 3973
rect 4526 3968 4527 3972
rect 4531 3968 4532 3972
rect 4526 3967 4532 3968
rect 4678 3972 4684 3973
rect 4678 3968 4679 3972
rect 4683 3968 4684 3972
rect 4678 3967 4684 3968
rect 4830 3972 4836 3973
rect 4830 3968 4831 3972
rect 4835 3968 4836 3972
rect 4830 3967 4836 3968
rect 4974 3972 4980 3973
rect 4974 3968 4975 3972
rect 4979 3968 4980 3972
rect 4974 3967 4980 3968
rect 5118 3972 5124 3973
rect 5118 3968 5119 3972
rect 5123 3968 5124 3972
rect 5118 3967 5124 3968
rect 5262 3972 5268 3973
rect 5262 3968 5263 3972
rect 5267 3968 5268 3972
rect 5262 3967 5268 3968
rect 5406 3972 5412 3973
rect 5406 3968 5407 3972
rect 5411 3968 5412 3972
rect 5406 3967 5412 3968
rect 5542 3972 5548 3973
rect 5542 3968 5543 3972
rect 5547 3968 5548 3972
rect 5542 3967 5548 3968
rect 5662 3971 5668 3972
rect 5662 3967 5663 3971
rect 5667 3967 5668 3971
rect 3838 3966 3844 3967
rect 5662 3966 5668 3967
rect 482 3957 488 3958
rect 110 3956 116 3957
rect 110 3952 111 3956
rect 115 3952 116 3956
rect 482 3953 483 3957
rect 487 3953 488 3957
rect 482 3952 488 3953
rect 634 3957 640 3958
rect 634 3953 635 3957
rect 639 3953 640 3957
rect 634 3952 640 3953
rect 794 3957 800 3958
rect 794 3953 795 3957
rect 799 3953 800 3957
rect 794 3952 800 3953
rect 954 3957 960 3958
rect 954 3953 955 3957
rect 959 3953 960 3957
rect 954 3952 960 3953
rect 1122 3957 1128 3958
rect 1122 3953 1123 3957
rect 1127 3953 1128 3957
rect 1122 3952 1128 3953
rect 1290 3957 1296 3958
rect 1290 3953 1291 3957
rect 1295 3953 1296 3957
rect 1290 3952 1296 3953
rect 1934 3956 1940 3957
rect 1934 3952 1935 3956
rect 1939 3952 1940 3956
rect 110 3951 116 3952
rect 1934 3951 1940 3952
rect 607 3947 616 3948
rect 607 3943 608 3947
rect 615 3943 616 3947
rect 607 3942 616 3943
rect 758 3947 765 3948
rect 758 3943 759 3947
rect 764 3943 765 3947
rect 758 3942 765 3943
rect 919 3947 925 3948
rect 919 3943 920 3947
rect 924 3946 925 3947
rect 942 3947 948 3948
rect 942 3946 943 3947
rect 924 3944 943 3946
rect 924 3943 925 3944
rect 919 3942 925 3943
rect 942 3943 943 3944
rect 947 3943 948 3947
rect 1079 3947 1085 3948
rect 1079 3946 1080 3947
rect 942 3942 948 3943
rect 952 3944 1080 3946
rect 578 3939 584 3940
rect 578 3935 579 3939
rect 583 3938 584 3939
rect 952 3938 954 3944
rect 1079 3943 1080 3944
rect 1084 3943 1085 3947
rect 1079 3942 1085 3943
rect 1247 3947 1256 3948
rect 1247 3943 1248 3947
rect 1255 3943 1256 3947
rect 1247 3942 1256 3943
rect 1370 3947 1376 3948
rect 1370 3943 1371 3947
rect 1375 3946 1376 3947
rect 1415 3947 1421 3948
rect 1415 3946 1416 3947
rect 1375 3944 1416 3946
rect 1375 3943 1376 3944
rect 1370 3942 1376 3943
rect 1415 3943 1416 3944
rect 1420 3943 1421 3947
rect 1415 3942 1421 3943
rect 583 3936 954 3938
rect 1974 3941 1980 3942
rect 3798 3941 3804 3942
rect 1974 3937 1975 3941
rect 1979 3937 1980 3941
rect 1974 3936 1980 3937
rect 2118 3940 2124 3941
rect 2118 3936 2119 3940
rect 2123 3936 2124 3940
rect 583 3935 584 3936
rect 2118 3935 2124 3936
rect 2326 3940 2332 3941
rect 2326 3936 2327 3940
rect 2331 3936 2332 3940
rect 2326 3935 2332 3936
rect 2534 3940 2540 3941
rect 2534 3936 2535 3940
rect 2539 3936 2540 3940
rect 2534 3935 2540 3936
rect 2742 3940 2748 3941
rect 2742 3936 2743 3940
rect 2747 3936 2748 3940
rect 2742 3935 2748 3936
rect 2942 3940 2948 3941
rect 2942 3936 2943 3940
rect 2947 3936 2948 3940
rect 2942 3935 2948 3936
rect 3134 3940 3140 3941
rect 3134 3936 3135 3940
rect 3139 3936 3140 3940
rect 3134 3935 3140 3936
rect 3318 3940 3324 3941
rect 3318 3936 3319 3940
rect 3323 3936 3324 3940
rect 3318 3935 3324 3936
rect 3510 3940 3516 3941
rect 3510 3936 3511 3940
rect 3515 3936 3516 3940
rect 3510 3935 3516 3936
rect 3678 3940 3684 3941
rect 3678 3936 3679 3940
rect 3683 3936 3684 3940
rect 3798 3937 3799 3941
rect 3803 3937 3804 3941
rect 3798 3936 3804 3937
rect 3678 3935 3684 3936
rect 578 3934 584 3935
rect 2090 3925 2096 3926
rect 1974 3924 1980 3925
rect 1974 3920 1975 3924
rect 1979 3920 1980 3924
rect 2090 3921 2091 3925
rect 2095 3921 2096 3925
rect 2090 3920 2096 3921
rect 2298 3925 2304 3926
rect 2298 3921 2299 3925
rect 2303 3921 2304 3925
rect 2298 3920 2304 3921
rect 2506 3925 2512 3926
rect 2506 3921 2507 3925
rect 2511 3921 2512 3925
rect 2506 3920 2512 3921
rect 2714 3925 2720 3926
rect 2714 3921 2715 3925
rect 2719 3921 2720 3925
rect 2714 3920 2720 3921
rect 2914 3925 2920 3926
rect 2914 3921 2915 3925
rect 2919 3921 2920 3925
rect 2914 3920 2920 3921
rect 3106 3925 3112 3926
rect 3106 3921 3107 3925
rect 3111 3921 3112 3925
rect 3106 3920 3112 3921
rect 3290 3925 3296 3926
rect 3290 3921 3291 3925
rect 3295 3921 3296 3925
rect 3290 3920 3296 3921
rect 3482 3925 3488 3926
rect 3482 3921 3483 3925
rect 3487 3921 3488 3925
rect 3482 3920 3488 3921
rect 3650 3925 3656 3926
rect 3650 3921 3651 3925
rect 3655 3921 3656 3925
rect 3650 3920 3656 3921
rect 3798 3924 3804 3925
rect 3798 3920 3799 3924
rect 3803 3920 3804 3924
rect 1974 3919 1980 3920
rect 3798 3919 3804 3920
rect 2214 3915 2221 3916
rect 2214 3911 2215 3915
rect 2220 3911 2221 3915
rect 2214 3910 2221 3911
rect 2290 3915 2296 3916
rect 2290 3911 2291 3915
rect 2295 3914 2296 3915
rect 2423 3915 2429 3916
rect 2423 3914 2424 3915
rect 2295 3912 2424 3914
rect 2295 3911 2296 3912
rect 2290 3910 2296 3911
rect 2423 3911 2424 3912
rect 2428 3911 2429 3915
rect 2423 3910 2429 3911
rect 2631 3915 2637 3916
rect 2631 3911 2632 3915
rect 2636 3914 2637 3915
rect 2671 3915 2677 3916
rect 2671 3914 2672 3915
rect 2636 3912 2672 3914
rect 2636 3911 2637 3912
rect 2631 3910 2637 3911
rect 2671 3911 2672 3912
rect 2676 3911 2677 3915
rect 2839 3915 2845 3916
rect 2839 3914 2840 3915
rect 2671 3910 2677 3911
rect 2779 3912 2840 3914
rect 578 3907 584 3908
rect 578 3903 579 3907
rect 583 3903 584 3907
rect 578 3902 584 3903
rect 610 3907 616 3908
rect 610 3903 611 3907
rect 615 3906 616 3907
rect 854 3907 860 3908
rect 615 3904 641 3906
rect 615 3903 616 3904
rect 610 3902 616 3903
rect 854 3903 855 3907
rect 859 3903 860 3907
rect 854 3902 860 3903
rect 942 3907 948 3908
rect 942 3903 943 3907
rect 947 3906 948 3907
rect 1218 3907 1224 3908
rect 947 3904 961 3906
rect 947 3903 948 3904
rect 942 3902 948 3903
rect 1218 3903 1219 3907
rect 1223 3903 1224 3907
rect 1218 3902 1224 3903
rect 1250 3907 1256 3908
rect 1250 3903 1251 3907
rect 1255 3906 1256 3907
rect 2394 3907 2400 3908
rect 1255 3904 1297 3906
rect 1255 3903 1256 3904
rect 1250 3902 1256 3903
rect 2394 3903 2395 3907
rect 2399 3906 2400 3907
rect 2779 3906 2781 3912
rect 2839 3911 2840 3912
rect 2844 3911 2845 3915
rect 2839 3910 2845 3911
rect 3039 3915 3048 3916
rect 3039 3911 3040 3915
rect 3047 3911 3048 3915
rect 3039 3910 3048 3911
rect 3231 3915 3240 3916
rect 3231 3911 3232 3915
rect 3239 3911 3240 3915
rect 3231 3910 3240 3911
rect 3415 3915 3424 3916
rect 3415 3911 3416 3915
rect 3423 3911 3424 3915
rect 3415 3910 3424 3911
rect 3607 3915 3616 3916
rect 3607 3911 3608 3915
rect 3615 3911 3616 3915
rect 3607 3910 3616 3911
rect 3775 3915 3781 3916
rect 3775 3911 3776 3915
rect 3780 3914 3781 3915
rect 3866 3915 3872 3916
rect 3866 3914 3867 3915
rect 3780 3912 3867 3914
rect 3780 3911 3781 3912
rect 3775 3910 3781 3911
rect 3866 3911 3867 3912
rect 3871 3911 3872 3915
rect 3866 3910 3872 3911
rect 2399 3904 2781 3906
rect 2399 3903 2400 3904
rect 2394 3902 2400 3903
rect 3838 3889 3844 3890
rect 5662 3889 5668 3890
rect 3838 3885 3839 3889
rect 3843 3885 3844 3889
rect 3838 3884 3844 3885
rect 4382 3888 4388 3889
rect 4382 3884 4383 3888
rect 4387 3884 4388 3888
rect 4382 3883 4388 3884
rect 4598 3888 4604 3889
rect 4598 3884 4599 3888
rect 4603 3884 4604 3888
rect 4598 3883 4604 3884
rect 4822 3888 4828 3889
rect 4822 3884 4823 3888
rect 4827 3884 4828 3888
rect 4822 3883 4828 3884
rect 5062 3888 5068 3889
rect 5062 3884 5063 3888
rect 5067 3884 5068 3888
rect 5062 3883 5068 3884
rect 5310 3888 5316 3889
rect 5310 3884 5311 3888
rect 5315 3884 5316 3888
rect 5310 3883 5316 3884
rect 5542 3888 5548 3889
rect 5542 3884 5543 3888
rect 5547 3884 5548 3888
rect 5662 3885 5663 3889
rect 5667 3885 5668 3889
rect 5662 3884 5668 3885
rect 5542 3883 5548 3884
rect 2290 3875 2296 3876
rect 2290 3874 2291 3875
rect 2189 3872 2291 3874
rect 2290 3871 2291 3872
rect 2295 3871 2296 3875
rect 2290 3870 2296 3871
rect 2394 3875 2400 3876
rect 2394 3871 2395 3875
rect 2399 3871 2400 3875
rect 2394 3870 2400 3871
rect 2550 3875 2556 3876
rect 2550 3871 2551 3875
rect 2555 3871 2556 3875
rect 2550 3870 2556 3871
rect 2671 3875 2677 3876
rect 2671 3871 2672 3875
rect 2676 3874 2677 3875
rect 3010 3875 3016 3876
rect 2676 3872 2721 3874
rect 2676 3871 2677 3872
rect 2671 3870 2677 3871
rect 3010 3871 3011 3875
rect 3015 3871 3016 3875
rect 3010 3870 3016 3871
rect 3042 3875 3048 3876
rect 3042 3871 3043 3875
rect 3047 3874 3048 3875
rect 3234 3875 3240 3876
rect 3047 3872 3113 3874
rect 3047 3871 3048 3872
rect 3042 3870 3048 3871
rect 3234 3871 3235 3875
rect 3239 3874 3240 3875
rect 3418 3875 3424 3876
rect 3239 3872 3297 3874
rect 3239 3871 3240 3872
rect 3234 3870 3240 3871
rect 3418 3871 3419 3875
rect 3423 3874 3424 3875
rect 3610 3875 3616 3876
rect 3423 3872 3489 3874
rect 3423 3871 3424 3872
rect 3418 3870 3424 3871
rect 3610 3871 3611 3875
rect 3615 3874 3616 3875
rect 3615 3872 3657 3874
rect 4354 3873 4360 3874
rect 3838 3872 3844 3873
rect 3615 3871 3616 3872
rect 3610 3870 3616 3871
rect 3838 3868 3839 3872
rect 3843 3868 3844 3872
rect 4354 3869 4355 3873
rect 4359 3869 4360 3873
rect 4354 3868 4360 3869
rect 4570 3873 4576 3874
rect 4570 3869 4571 3873
rect 4575 3869 4576 3873
rect 4570 3868 4576 3869
rect 4794 3873 4800 3874
rect 4794 3869 4795 3873
rect 4799 3869 4800 3873
rect 4794 3868 4800 3869
rect 5034 3873 5040 3874
rect 5034 3869 5035 3873
rect 5039 3869 5040 3873
rect 5034 3868 5040 3869
rect 5282 3873 5288 3874
rect 5282 3869 5283 3873
rect 5287 3869 5288 3873
rect 5282 3868 5288 3869
rect 5514 3873 5520 3874
rect 5514 3869 5515 3873
rect 5519 3869 5520 3873
rect 5514 3868 5520 3869
rect 5662 3872 5668 3873
rect 5662 3868 5663 3872
rect 5667 3868 5668 3872
rect 3838 3867 3844 3868
rect 5662 3867 5668 3868
rect 5407 3864 5413 3865
rect 4479 3863 4488 3864
rect 4479 3859 4480 3863
rect 4487 3859 4488 3863
rect 4479 3858 4488 3859
rect 4695 3863 4704 3864
rect 4695 3859 4696 3863
rect 4703 3859 4704 3863
rect 4695 3858 4704 3859
rect 4919 3863 4928 3864
rect 4919 3859 4920 3863
rect 4927 3859 4928 3863
rect 4919 3858 4928 3859
rect 5058 3863 5064 3864
rect 5058 3859 5059 3863
rect 5063 3862 5064 3863
rect 5159 3863 5165 3864
rect 5159 3862 5160 3863
rect 5063 3860 5160 3862
rect 5063 3859 5064 3860
rect 5058 3858 5064 3859
rect 5159 3859 5160 3860
rect 5164 3859 5165 3863
rect 5159 3858 5165 3859
rect 5398 3863 5404 3864
rect 5398 3859 5399 3863
rect 5403 3862 5404 3863
rect 5407 3862 5408 3864
rect 5403 3860 5408 3862
rect 5412 3860 5413 3864
rect 5403 3859 5404 3860
rect 5407 3859 5413 3860
rect 5610 3863 5616 3864
rect 5610 3859 5611 3863
rect 5615 3862 5616 3863
rect 5639 3863 5645 3864
rect 5639 3862 5640 3863
rect 5615 3860 5640 3862
rect 5615 3859 5616 3860
rect 5398 3858 5404 3859
rect 5610 3858 5616 3859
rect 5639 3859 5640 3860
rect 5644 3859 5645 3863
rect 5639 3858 5645 3859
rect 626 3855 632 3856
rect 626 3854 627 3855
rect 259 3852 627 3854
rect 259 3846 261 3852
rect 626 3851 627 3852
rect 631 3851 632 3855
rect 626 3850 632 3851
rect 719 3847 725 3848
rect 719 3846 720 3847
rect 229 3844 261 3846
rect 613 3844 720 3846
rect 314 3843 320 3844
rect 314 3839 315 3843
rect 319 3839 320 3843
rect 719 3843 720 3844
rect 724 3843 725 3847
rect 719 3842 725 3843
rect 758 3847 764 3848
rect 758 3843 759 3847
rect 763 3843 764 3847
rect 1150 3847 1156 3848
rect 1150 3846 1151 3847
rect 1037 3844 1151 3846
rect 758 3842 764 3843
rect 1150 3843 1151 3844
rect 1155 3843 1156 3847
rect 1150 3842 1156 3843
rect 1170 3843 1176 3844
rect 314 3838 320 3839
rect 1170 3839 1171 3843
rect 1175 3839 1176 3843
rect 1170 3838 1176 3839
rect 2214 3831 2220 3832
rect 2214 3827 2215 3831
rect 2219 3827 2220 3831
rect 2214 3826 2220 3827
rect 2378 3827 2384 3828
rect 2378 3823 2379 3827
rect 2383 3823 2384 3827
rect 2378 3822 2384 3823
rect 2594 3827 2600 3828
rect 2594 3823 2595 3827
rect 2599 3823 2600 3827
rect 2594 3822 2600 3823
rect 2802 3827 2808 3828
rect 2802 3823 2803 3827
rect 2807 3823 2808 3827
rect 2802 3822 2808 3823
rect 3002 3827 3008 3828
rect 3002 3823 3003 3827
rect 3007 3823 3008 3827
rect 3002 3822 3008 3823
rect 3202 3827 3208 3828
rect 3202 3823 3203 3827
rect 3207 3823 3208 3827
rect 3202 3822 3208 3823
rect 3410 3827 3416 3828
rect 3410 3823 3411 3827
rect 3415 3823 3416 3827
rect 3410 3822 3416 3823
rect 4450 3823 4456 3824
rect 4450 3819 4451 3823
rect 4455 3819 4456 3823
rect 4450 3818 4456 3819
rect 4482 3823 4488 3824
rect 4482 3819 4483 3823
rect 4487 3822 4488 3823
rect 4698 3823 4704 3824
rect 4487 3820 4577 3822
rect 4487 3819 4488 3820
rect 4482 3818 4488 3819
rect 4698 3819 4699 3823
rect 4703 3822 4704 3823
rect 4922 3823 4928 3824
rect 4703 3820 4801 3822
rect 4703 3819 4704 3820
rect 4698 3818 4704 3819
rect 4922 3819 4923 3823
rect 4927 3822 4928 3823
rect 5374 3823 5380 3824
rect 4927 3820 5041 3822
rect 4927 3819 4928 3820
rect 4922 3818 4928 3819
rect 5374 3819 5375 3823
rect 5379 3819 5380 3823
rect 5634 3823 5640 3824
rect 5634 3822 5635 3823
rect 5613 3820 5635 3822
rect 5374 3818 5380 3819
rect 5634 3819 5635 3820
rect 5639 3819 5640 3823
rect 5634 3818 5640 3819
rect 255 3803 261 3804
rect 255 3799 256 3803
rect 260 3802 261 3803
rect 314 3803 320 3804
rect 314 3802 315 3803
rect 260 3800 315 3802
rect 260 3799 261 3800
rect 255 3798 261 3799
rect 314 3799 315 3800
rect 319 3799 320 3803
rect 314 3798 320 3799
rect 402 3803 408 3804
rect 402 3799 403 3803
rect 407 3802 408 3803
rect 431 3803 437 3804
rect 431 3802 432 3803
rect 407 3800 432 3802
rect 407 3799 408 3800
rect 402 3798 408 3799
rect 431 3799 432 3800
rect 436 3799 437 3803
rect 431 3798 437 3799
rect 626 3803 632 3804
rect 626 3799 627 3803
rect 631 3802 632 3803
rect 639 3803 645 3804
rect 639 3802 640 3803
rect 631 3800 640 3802
rect 631 3799 632 3800
rect 626 3798 632 3799
rect 639 3799 640 3800
rect 644 3799 645 3803
rect 639 3798 645 3799
rect 719 3803 725 3804
rect 719 3799 720 3803
rect 724 3802 725 3803
rect 847 3803 853 3804
rect 847 3802 848 3803
rect 724 3800 848 3802
rect 724 3799 725 3800
rect 719 3798 725 3799
rect 847 3799 848 3800
rect 852 3799 853 3803
rect 847 3798 853 3799
rect 1063 3803 1069 3804
rect 1063 3799 1064 3803
rect 1068 3802 1069 3803
rect 1170 3803 1176 3804
rect 1170 3802 1171 3803
rect 1068 3800 1171 3802
rect 1068 3799 1069 3800
rect 1063 3798 1069 3799
rect 1170 3799 1171 3800
rect 1175 3799 1176 3803
rect 1170 3798 1176 3799
rect 1218 3803 1224 3804
rect 1218 3799 1219 3803
rect 1223 3802 1224 3803
rect 1287 3803 1293 3804
rect 1287 3802 1288 3803
rect 1223 3800 1288 3802
rect 1223 3799 1224 3800
rect 1218 3798 1224 3799
rect 1287 3799 1288 3800
rect 1292 3799 1293 3803
rect 1287 3798 1293 3799
rect 110 3796 116 3797
rect 1934 3796 1940 3797
rect 110 3792 111 3796
rect 115 3792 116 3796
rect 110 3791 116 3792
rect 130 3795 136 3796
rect 130 3791 131 3795
rect 135 3791 136 3795
rect 130 3790 136 3791
rect 306 3795 312 3796
rect 306 3791 307 3795
rect 311 3791 312 3795
rect 306 3790 312 3791
rect 514 3795 520 3796
rect 514 3791 515 3795
rect 519 3791 520 3795
rect 514 3790 520 3791
rect 722 3795 728 3796
rect 722 3791 723 3795
rect 727 3791 728 3795
rect 722 3790 728 3791
rect 938 3795 944 3796
rect 938 3791 939 3795
rect 943 3791 944 3795
rect 938 3790 944 3791
rect 1162 3795 1168 3796
rect 1162 3791 1163 3795
rect 1167 3791 1168 3795
rect 1934 3792 1935 3796
rect 1939 3792 1940 3796
rect 1934 3791 1940 3792
rect 1162 3790 1168 3791
rect 2263 3787 2269 3788
rect 2263 3783 2264 3787
rect 2268 3786 2269 3787
rect 2378 3787 2384 3788
rect 2378 3786 2379 3787
rect 2268 3784 2379 3786
rect 2268 3783 2269 3784
rect 2263 3782 2269 3783
rect 2378 3783 2379 3784
rect 2383 3783 2384 3787
rect 2378 3782 2384 3783
rect 2390 3787 2396 3788
rect 2390 3783 2391 3787
rect 2395 3786 2396 3787
rect 2495 3787 2501 3788
rect 2495 3786 2496 3787
rect 2395 3784 2496 3786
rect 2395 3783 2396 3784
rect 2390 3782 2396 3783
rect 2495 3783 2496 3784
rect 2500 3783 2501 3787
rect 2495 3782 2501 3783
rect 2711 3787 2717 3788
rect 2711 3783 2712 3787
rect 2716 3786 2717 3787
rect 2802 3787 2808 3788
rect 2802 3786 2803 3787
rect 2716 3784 2803 3786
rect 2716 3783 2717 3784
rect 2711 3782 2717 3783
rect 2802 3783 2803 3784
rect 2807 3783 2808 3787
rect 2802 3782 2808 3783
rect 2919 3787 2925 3788
rect 2919 3783 2920 3787
rect 2924 3786 2925 3787
rect 3002 3787 3008 3788
rect 3002 3786 3003 3787
rect 2924 3784 3003 3786
rect 2924 3783 2925 3784
rect 2919 3782 2925 3783
rect 3002 3783 3003 3784
rect 3007 3783 3008 3787
rect 3002 3782 3008 3783
rect 3119 3787 3125 3788
rect 3119 3783 3120 3787
rect 3124 3786 3125 3787
rect 3202 3787 3208 3788
rect 3202 3786 3203 3787
rect 3124 3784 3203 3786
rect 3124 3783 3125 3784
rect 3119 3782 3125 3783
rect 3202 3783 3203 3784
rect 3207 3783 3208 3787
rect 3202 3782 3208 3783
rect 3319 3787 3325 3788
rect 3319 3783 3320 3787
rect 3324 3786 3325 3787
rect 3410 3787 3416 3788
rect 3410 3786 3411 3787
rect 3324 3784 3411 3786
rect 3324 3783 3325 3784
rect 3319 3782 3325 3783
rect 3410 3783 3411 3784
rect 3415 3783 3416 3787
rect 3410 3782 3416 3783
rect 3418 3787 3424 3788
rect 3418 3783 3419 3787
rect 3423 3786 3424 3787
rect 3527 3787 3533 3788
rect 3527 3786 3528 3787
rect 3423 3784 3528 3786
rect 3423 3783 3424 3784
rect 3418 3782 3424 3783
rect 3527 3783 3528 3784
rect 3532 3783 3533 3787
rect 3527 3782 3533 3783
rect 158 3780 164 3781
rect 110 3779 116 3780
rect 110 3775 111 3779
rect 115 3775 116 3779
rect 158 3776 159 3780
rect 163 3776 164 3780
rect 158 3775 164 3776
rect 334 3780 340 3781
rect 334 3776 335 3780
rect 339 3776 340 3780
rect 334 3775 340 3776
rect 542 3780 548 3781
rect 542 3776 543 3780
rect 547 3776 548 3780
rect 542 3775 548 3776
rect 750 3780 756 3781
rect 750 3776 751 3780
rect 755 3776 756 3780
rect 750 3775 756 3776
rect 966 3780 972 3781
rect 966 3776 967 3780
rect 971 3776 972 3780
rect 966 3775 972 3776
rect 1190 3780 1196 3781
rect 1974 3780 1980 3781
rect 3798 3780 3804 3781
rect 1190 3776 1191 3780
rect 1195 3776 1196 3780
rect 1190 3775 1196 3776
rect 1934 3779 1940 3780
rect 1934 3775 1935 3779
rect 1939 3775 1940 3779
rect 1974 3776 1975 3780
rect 1979 3776 1980 3780
rect 1974 3775 1980 3776
rect 2138 3779 2144 3780
rect 2138 3775 2139 3779
rect 2143 3775 2144 3779
rect 110 3774 116 3775
rect 1934 3774 1940 3775
rect 2138 3774 2144 3775
rect 2370 3779 2376 3780
rect 2370 3775 2371 3779
rect 2375 3775 2376 3779
rect 2370 3774 2376 3775
rect 2586 3779 2592 3780
rect 2586 3775 2587 3779
rect 2591 3775 2592 3779
rect 2586 3774 2592 3775
rect 2794 3779 2800 3780
rect 2794 3775 2795 3779
rect 2799 3775 2800 3779
rect 2794 3774 2800 3775
rect 2994 3779 3000 3780
rect 2994 3775 2995 3779
rect 2999 3775 3000 3779
rect 2994 3774 3000 3775
rect 3194 3779 3200 3780
rect 3194 3775 3195 3779
rect 3199 3775 3200 3779
rect 3194 3774 3200 3775
rect 3402 3779 3408 3780
rect 3402 3775 3403 3779
rect 3407 3775 3408 3779
rect 3798 3776 3799 3780
rect 3803 3776 3804 3780
rect 3798 3775 3804 3776
rect 5058 3775 5064 3776
rect 3402 3774 3408 3775
rect 4090 3771 4096 3772
rect 4090 3767 4091 3771
rect 4095 3767 4096 3771
rect 4090 3766 4096 3767
rect 4210 3771 4216 3772
rect 4210 3767 4211 3771
rect 4215 3767 4216 3771
rect 4210 3766 4216 3767
rect 4442 3771 4448 3772
rect 4442 3767 4443 3771
rect 4447 3767 4448 3771
rect 4442 3766 4448 3767
rect 4698 3771 4704 3772
rect 4698 3767 4699 3771
rect 4703 3767 4704 3771
rect 5058 3771 5059 3775
rect 5063 3771 5064 3775
rect 5610 3775 5616 3776
rect 5058 3770 5064 3771
rect 5346 3771 5352 3772
rect 4698 3766 4704 3767
rect 5346 3767 5347 3771
rect 5351 3767 5352 3771
rect 5610 3771 5611 3775
rect 5615 3771 5616 3775
rect 5610 3770 5616 3771
rect 5346 3766 5352 3767
rect 2166 3764 2172 3765
rect 1974 3763 1980 3764
rect 1974 3759 1975 3763
rect 1979 3759 1980 3763
rect 2166 3760 2167 3764
rect 2171 3760 2172 3764
rect 2166 3759 2172 3760
rect 2398 3764 2404 3765
rect 2398 3760 2399 3764
rect 2403 3760 2404 3764
rect 2398 3759 2404 3760
rect 2614 3764 2620 3765
rect 2614 3760 2615 3764
rect 2619 3760 2620 3764
rect 2614 3759 2620 3760
rect 2822 3764 2828 3765
rect 2822 3760 2823 3764
rect 2827 3760 2828 3764
rect 2822 3759 2828 3760
rect 3022 3764 3028 3765
rect 3022 3760 3023 3764
rect 3027 3760 3028 3764
rect 3022 3759 3028 3760
rect 3222 3764 3228 3765
rect 3222 3760 3223 3764
rect 3227 3760 3228 3764
rect 3222 3759 3228 3760
rect 3430 3764 3436 3765
rect 3430 3760 3431 3764
rect 3435 3760 3436 3764
rect 3430 3759 3436 3760
rect 3798 3763 3804 3764
rect 3798 3759 3799 3763
rect 3803 3759 3804 3763
rect 1974 3758 1980 3759
rect 3798 3758 3804 3759
rect 4119 3731 4125 3732
rect 4119 3727 4120 3731
rect 4124 3730 4125 3731
rect 4210 3731 4216 3732
rect 4210 3730 4211 3731
rect 4124 3728 4211 3730
rect 4124 3727 4125 3728
rect 4119 3726 4125 3727
rect 4210 3727 4211 3728
rect 4215 3727 4216 3731
rect 4210 3726 4216 3727
rect 4327 3731 4333 3732
rect 4327 3727 4328 3731
rect 4332 3730 4333 3731
rect 4442 3731 4448 3732
rect 4442 3730 4443 3731
rect 4332 3728 4443 3730
rect 4332 3727 4333 3728
rect 4327 3726 4333 3727
rect 4442 3727 4443 3728
rect 4447 3727 4448 3731
rect 4442 3726 4448 3727
rect 4559 3731 4565 3732
rect 4559 3727 4560 3731
rect 4564 3730 4565 3731
rect 4698 3731 4704 3732
rect 4698 3730 4699 3731
rect 4564 3728 4699 3730
rect 4564 3727 4565 3728
rect 4559 3726 4565 3727
rect 4698 3727 4699 3728
rect 4703 3727 4704 3731
rect 4698 3726 4704 3727
rect 4814 3731 4821 3732
rect 4814 3727 4815 3731
rect 4820 3727 4821 3731
rect 4814 3726 4821 3727
rect 4938 3731 4944 3732
rect 4938 3727 4939 3731
rect 4943 3730 4944 3731
rect 5087 3731 5093 3732
rect 5087 3730 5088 3731
rect 4943 3728 5088 3730
rect 4943 3727 4944 3728
rect 4938 3726 4944 3727
rect 5087 3727 5088 3728
rect 5092 3727 5093 3731
rect 5087 3726 5093 3727
rect 5374 3731 5381 3732
rect 5374 3727 5375 3731
rect 5380 3727 5381 3731
rect 5374 3726 5381 3727
rect 5626 3731 5632 3732
rect 5626 3727 5627 3731
rect 5631 3730 5632 3731
rect 5639 3731 5645 3732
rect 5639 3730 5640 3731
rect 5631 3728 5640 3730
rect 5631 3727 5632 3728
rect 5626 3726 5632 3727
rect 5639 3727 5640 3728
rect 5644 3727 5645 3731
rect 5639 3726 5645 3727
rect 3838 3724 3844 3725
rect 5662 3724 5668 3725
rect 110 3721 116 3722
rect 1934 3721 1940 3722
rect 110 3717 111 3721
rect 115 3717 116 3721
rect 110 3716 116 3717
rect 158 3720 164 3721
rect 158 3716 159 3720
rect 163 3716 164 3720
rect 158 3715 164 3716
rect 334 3720 340 3721
rect 334 3716 335 3720
rect 339 3716 340 3720
rect 334 3715 340 3716
rect 526 3720 532 3721
rect 526 3716 527 3720
rect 531 3716 532 3720
rect 526 3715 532 3716
rect 710 3720 716 3721
rect 710 3716 711 3720
rect 715 3716 716 3720
rect 710 3715 716 3716
rect 886 3720 892 3721
rect 886 3716 887 3720
rect 891 3716 892 3720
rect 886 3715 892 3716
rect 1054 3720 1060 3721
rect 1054 3716 1055 3720
rect 1059 3716 1060 3720
rect 1054 3715 1060 3716
rect 1214 3720 1220 3721
rect 1214 3716 1215 3720
rect 1219 3716 1220 3720
rect 1214 3715 1220 3716
rect 1366 3720 1372 3721
rect 1366 3716 1367 3720
rect 1371 3716 1372 3720
rect 1366 3715 1372 3716
rect 1518 3720 1524 3721
rect 1518 3716 1519 3720
rect 1523 3716 1524 3720
rect 1518 3715 1524 3716
rect 1678 3720 1684 3721
rect 1678 3716 1679 3720
rect 1683 3716 1684 3720
rect 1678 3715 1684 3716
rect 1814 3720 1820 3721
rect 1814 3716 1815 3720
rect 1819 3716 1820 3720
rect 1934 3717 1935 3721
rect 1939 3717 1940 3721
rect 3838 3720 3839 3724
rect 3843 3720 3844 3724
rect 3838 3719 3844 3720
rect 3994 3723 4000 3724
rect 3994 3719 3995 3723
rect 3999 3719 4000 3723
rect 3994 3718 4000 3719
rect 4202 3723 4208 3724
rect 4202 3719 4203 3723
rect 4207 3719 4208 3723
rect 4202 3718 4208 3719
rect 4434 3723 4440 3724
rect 4434 3719 4435 3723
rect 4439 3719 4440 3723
rect 4434 3718 4440 3719
rect 4690 3723 4696 3724
rect 4690 3719 4691 3723
rect 4695 3719 4696 3723
rect 4690 3718 4696 3719
rect 4962 3723 4968 3724
rect 4962 3719 4963 3723
rect 4967 3719 4968 3723
rect 4962 3718 4968 3719
rect 5250 3723 5256 3724
rect 5250 3719 5251 3723
rect 5255 3719 5256 3723
rect 5250 3718 5256 3719
rect 5514 3723 5520 3724
rect 5514 3719 5515 3723
rect 5519 3719 5520 3723
rect 5662 3720 5663 3724
rect 5667 3720 5668 3724
rect 5662 3719 5668 3720
rect 5514 3718 5520 3719
rect 1934 3716 1940 3717
rect 1814 3715 1820 3716
rect 4022 3708 4028 3709
rect 3838 3707 3844 3708
rect 130 3705 136 3706
rect 110 3704 116 3705
rect 110 3700 111 3704
rect 115 3700 116 3704
rect 130 3701 131 3705
rect 135 3701 136 3705
rect 130 3700 136 3701
rect 306 3705 312 3706
rect 306 3701 307 3705
rect 311 3701 312 3705
rect 306 3700 312 3701
rect 498 3705 504 3706
rect 498 3701 499 3705
rect 503 3701 504 3705
rect 498 3700 504 3701
rect 682 3705 688 3706
rect 682 3701 683 3705
rect 687 3701 688 3705
rect 682 3700 688 3701
rect 858 3705 864 3706
rect 858 3701 859 3705
rect 863 3701 864 3705
rect 858 3700 864 3701
rect 1026 3705 1032 3706
rect 1026 3701 1027 3705
rect 1031 3701 1032 3705
rect 1026 3700 1032 3701
rect 1186 3705 1192 3706
rect 1186 3701 1187 3705
rect 1191 3701 1192 3705
rect 1186 3700 1192 3701
rect 1338 3705 1344 3706
rect 1338 3701 1339 3705
rect 1343 3701 1344 3705
rect 1338 3700 1344 3701
rect 1490 3705 1496 3706
rect 1490 3701 1491 3705
rect 1495 3701 1496 3705
rect 1490 3700 1496 3701
rect 1650 3705 1656 3706
rect 1650 3701 1651 3705
rect 1655 3701 1656 3705
rect 1650 3700 1656 3701
rect 1786 3705 1792 3706
rect 1786 3701 1787 3705
rect 1791 3701 1792 3705
rect 1786 3700 1792 3701
rect 1934 3704 1940 3705
rect 1934 3700 1935 3704
rect 1939 3700 1940 3704
rect 3838 3703 3839 3707
rect 3843 3703 3844 3707
rect 4022 3704 4023 3708
rect 4027 3704 4028 3708
rect 4022 3703 4028 3704
rect 4230 3708 4236 3709
rect 4230 3704 4231 3708
rect 4235 3704 4236 3708
rect 4230 3703 4236 3704
rect 4462 3708 4468 3709
rect 4462 3704 4463 3708
rect 4467 3704 4468 3708
rect 4462 3703 4468 3704
rect 4718 3708 4724 3709
rect 4718 3704 4719 3708
rect 4723 3704 4724 3708
rect 4718 3703 4724 3704
rect 4990 3708 4996 3709
rect 4990 3704 4991 3708
rect 4995 3704 4996 3708
rect 4990 3703 4996 3704
rect 5278 3708 5284 3709
rect 5278 3704 5279 3708
rect 5283 3704 5284 3708
rect 5278 3703 5284 3704
rect 5542 3708 5548 3709
rect 5542 3704 5543 3708
rect 5547 3704 5548 3708
rect 5542 3703 5548 3704
rect 5662 3707 5668 3708
rect 5662 3703 5663 3707
rect 5667 3703 5668 3707
rect 3838 3702 3844 3703
rect 5662 3702 5668 3703
rect 110 3699 116 3700
rect 1934 3699 1940 3700
rect 1974 3701 1980 3702
rect 3798 3701 3804 3702
rect 1974 3697 1975 3701
rect 1979 3697 1980 3701
rect 1974 3696 1980 3697
rect 2278 3700 2284 3701
rect 2278 3696 2279 3700
rect 2283 3696 2284 3700
rect 242 3695 248 3696
rect 242 3691 243 3695
rect 247 3694 248 3695
rect 255 3695 261 3696
rect 255 3694 256 3695
rect 247 3692 256 3694
rect 247 3691 248 3692
rect 242 3690 248 3691
rect 255 3691 256 3692
rect 260 3691 261 3695
rect 255 3690 261 3691
rect 431 3695 440 3696
rect 431 3691 432 3695
rect 439 3691 440 3695
rect 623 3695 629 3696
rect 623 3694 624 3695
rect 431 3690 440 3691
rect 444 3692 624 3694
rect 226 3687 232 3688
rect 226 3683 227 3687
rect 231 3686 232 3687
rect 444 3686 446 3692
rect 623 3691 624 3692
rect 628 3691 629 3695
rect 623 3690 629 3691
rect 807 3695 816 3696
rect 807 3691 808 3695
rect 815 3691 816 3695
rect 807 3690 816 3691
rect 983 3695 989 3696
rect 983 3691 984 3695
rect 988 3694 989 3695
rect 1130 3695 1136 3696
rect 1130 3694 1131 3695
rect 988 3692 1131 3694
rect 988 3691 989 3692
rect 983 3690 989 3691
rect 1130 3691 1131 3692
rect 1135 3691 1136 3695
rect 1130 3690 1136 3691
rect 1150 3695 1157 3696
rect 1150 3691 1151 3695
rect 1156 3691 1157 3695
rect 1150 3690 1157 3691
rect 1311 3695 1320 3696
rect 1311 3691 1312 3695
rect 1319 3691 1320 3695
rect 1311 3690 1320 3691
rect 1463 3695 1472 3696
rect 1463 3691 1464 3695
rect 1471 3691 1472 3695
rect 1463 3690 1472 3691
rect 1615 3695 1621 3696
rect 1615 3691 1616 3695
rect 1620 3694 1621 3695
rect 1638 3695 1644 3696
rect 1638 3694 1639 3695
rect 1620 3692 1639 3694
rect 1620 3691 1621 3692
rect 1615 3690 1621 3691
rect 1638 3691 1639 3692
rect 1643 3691 1644 3695
rect 1638 3690 1644 3691
rect 1775 3695 1784 3696
rect 1775 3691 1776 3695
rect 1783 3691 1784 3695
rect 1775 3690 1784 3691
rect 1882 3695 1888 3696
rect 1882 3691 1883 3695
rect 1887 3694 1888 3695
rect 1911 3695 1917 3696
rect 2278 3695 2284 3696
rect 2478 3700 2484 3701
rect 2478 3696 2479 3700
rect 2483 3696 2484 3700
rect 2478 3695 2484 3696
rect 2678 3700 2684 3701
rect 2678 3696 2679 3700
rect 2683 3696 2684 3700
rect 2678 3695 2684 3696
rect 2878 3700 2884 3701
rect 2878 3696 2879 3700
rect 2883 3696 2884 3700
rect 2878 3695 2884 3696
rect 3078 3700 3084 3701
rect 3078 3696 3079 3700
rect 3083 3696 3084 3700
rect 3078 3695 3084 3696
rect 3278 3700 3284 3701
rect 3278 3696 3279 3700
rect 3283 3696 3284 3700
rect 3798 3697 3799 3701
rect 3803 3697 3804 3701
rect 3798 3696 3804 3697
rect 3278 3695 3284 3696
rect 1911 3694 1912 3695
rect 1887 3692 1912 3694
rect 1887 3691 1888 3692
rect 1882 3690 1888 3691
rect 1911 3691 1912 3692
rect 1916 3691 1917 3695
rect 1911 3690 1917 3691
rect 231 3684 446 3686
rect 2250 3685 2256 3686
rect 1974 3684 1980 3685
rect 231 3683 232 3684
rect 226 3682 232 3683
rect 1974 3680 1975 3684
rect 1979 3680 1980 3684
rect 2250 3681 2251 3685
rect 2255 3681 2256 3685
rect 2250 3680 2256 3681
rect 2450 3685 2456 3686
rect 2450 3681 2451 3685
rect 2455 3681 2456 3685
rect 2450 3680 2456 3681
rect 2650 3685 2656 3686
rect 2650 3681 2651 3685
rect 2655 3681 2656 3685
rect 2650 3680 2656 3681
rect 2850 3685 2856 3686
rect 2850 3681 2851 3685
rect 2855 3681 2856 3685
rect 2850 3680 2856 3681
rect 3050 3685 3056 3686
rect 3050 3681 3051 3685
rect 3055 3681 3056 3685
rect 3050 3680 3056 3681
rect 3250 3685 3256 3686
rect 3250 3681 3251 3685
rect 3255 3681 3256 3685
rect 3250 3680 3256 3681
rect 3798 3684 3804 3685
rect 3798 3680 3799 3684
rect 3803 3680 3804 3684
rect 1974 3679 1980 3680
rect 3798 3679 3804 3680
rect 2346 3675 2352 3676
rect 2346 3671 2347 3675
rect 2351 3674 2352 3675
rect 2375 3675 2381 3676
rect 2375 3674 2376 3675
rect 2351 3672 2376 3674
rect 2351 3671 2352 3672
rect 2346 3670 2352 3671
rect 2375 3671 2376 3672
rect 2380 3671 2381 3675
rect 2375 3670 2381 3671
rect 2575 3675 2581 3676
rect 2575 3671 2576 3675
rect 2580 3674 2581 3675
rect 2594 3675 2600 3676
rect 2594 3674 2595 3675
rect 2580 3672 2595 3674
rect 2580 3671 2581 3672
rect 2575 3670 2581 3671
rect 2594 3671 2595 3672
rect 2599 3671 2600 3675
rect 2594 3670 2600 3671
rect 2647 3675 2653 3676
rect 2647 3671 2648 3675
rect 2652 3674 2653 3675
rect 2775 3675 2781 3676
rect 2775 3674 2776 3675
rect 2652 3672 2776 3674
rect 2652 3671 2653 3672
rect 2647 3670 2653 3671
rect 2775 3671 2776 3672
rect 2780 3671 2781 3675
rect 2775 3670 2781 3671
rect 2847 3675 2853 3676
rect 2847 3671 2848 3675
rect 2852 3674 2853 3675
rect 2975 3675 2981 3676
rect 2975 3674 2976 3675
rect 2852 3672 2976 3674
rect 2852 3671 2853 3672
rect 2847 3670 2853 3671
rect 2975 3671 2976 3672
rect 2980 3671 2981 3675
rect 2975 3670 2981 3671
rect 3175 3675 3181 3676
rect 3175 3671 3176 3675
rect 3180 3674 3181 3675
rect 3207 3675 3213 3676
rect 3207 3674 3208 3675
rect 3180 3672 3208 3674
rect 3180 3671 3181 3672
rect 3175 3670 3181 3671
rect 3207 3671 3208 3672
rect 3212 3671 3213 3675
rect 3375 3675 3381 3676
rect 3375 3674 3376 3675
rect 3207 3670 3213 3671
rect 3256 3672 3376 3674
rect 2946 3667 2952 3668
rect 2946 3663 2947 3667
rect 2951 3666 2952 3667
rect 3256 3666 3258 3672
rect 3375 3671 3376 3672
rect 3380 3671 3381 3675
rect 3375 3670 3381 3671
rect 2951 3664 3258 3666
rect 2951 3663 2952 3664
rect 2946 3662 2952 3663
rect 226 3655 232 3656
rect 226 3651 227 3655
rect 231 3651 232 3655
rect 226 3650 232 3651
rect 402 3655 408 3656
rect 402 3651 403 3655
rect 407 3651 408 3655
rect 402 3650 408 3651
rect 434 3655 440 3656
rect 434 3651 435 3655
rect 439 3654 440 3655
rect 810 3655 816 3656
rect 439 3652 505 3654
rect 439 3651 440 3652
rect 434 3650 440 3651
rect 780 3646 782 3653
rect 810 3651 811 3655
rect 815 3654 816 3655
rect 1122 3655 1128 3656
rect 815 3652 865 3654
rect 815 3651 816 3652
rect 810 3650 816 3651
rect 1122 3651 1123 3655
rect 1127 3651 1128 3655
rect 1122 3650 1128 3651
rect 1130 3655 1136 3656
rect 1130 3651 1131 3655
rect 1135 3654 1136 3655
rect 1314 3655 1320 3656
rect 1135 3652 1193 3654
rect 1135 3651 1136 3652
rect 1130 3650 1136 3651
rect 1314 3651 1315 3655
rect 1319 3654 1320 3655
rect 1466 3655 1472 3656
rect 1319 3652 1345 3654
rect 1319 3651 1320 3652
rect 1314 3650 1320 3651
rect 1466 3651 1467 3655
rect 1471 3654 1472 3655
rect 1638 3655 1644 3656
rect 1471 3652 1497 3654
rect 1471 3651 1472 3652
rect 1466 3650 1472 3651
rect 1638 3651 1639 3655
rect 1643 3654 1644 3655
rect 1778 3655 1784 3656
rect 1643 3652 1657 3654
rect 1643 3651 1644 3652
rect 1638 3650 1644 3651
rect 1778 3651 1779 3655
rect 1783 3654 1784 3655
rect 1783 3652 1793 3654
rect 1783 3651 1784 3652
rect 1778 3650 1784 3651
rect 1414 3647 1420 3648
rect 1414 3646 1415 3647
rect 780 3644 1415 3646
rect 1414 3643 1415 3644
rect 1419 3643 1420 3647
rect 1414 3642 1420 3643
rect 2847 3643 2853 3644
rect 2847 3642 2848 3643
rect 2779 3640 2848 3642
rect 2390 3635 2396 3636
rect 2390 3634 2391 3635
rect 2349 3632 2391 3634
rect 2390 3631 2391 3632
rect 2395 3631 2396 3635
rect 2647 3635 2653 3636
rect 2647 3634 2648 3635
rect 2549 3632 2648 3634
rect 2390 3630 2396 3631
rect 2647 3631 2648 3632
rect 2652 3631 2653 3635
rect 2779 3634 2781 3640
rect 2847 3639 2848 3640
rect 2852 3639 2853 3643
rect 2847 3638 2853 3639
rect 2749 3632 2781 3634
rect 2946 3635 2952 3636
rect 2647 3630 2653 3631
rect 2946 3631 2947 3635
rect 2951 3631 2952 3635
rect 2946 3630 2952 3631
rect 3102 3635 3108 3636
rect 3102 3631 3103 3635
rect 3107 3631 3108 3635
rect 3102 3630 3108 3631
rect 3207 3635 3213 3636
rect 3207 3631 3208 3635
rect 3212 3634 3213 3635
rect 3212 3632 3257 3634
rect 3212 3631 3213 3632
rect 3207 3630 3213 3631
rect 3838 3621 3844 3622
rect 5662 3621 5668 3622
rect 1670 3619 1676 3620
rect 1670 3618 1671 3619
rect 1480 3616 1671 3618
rect 242 3611 248 3612
rect 242 3607 243 3611
rect 247 3607 248 3611
rect 1480 3610 1482 3616
rect 1670 3615 1671 3616
rect 1675 3615 1676 3619
rect 3838 3617 3839 3621
rect 3843 3617 3844 3621
rect 3838 3616 3844 3617
rect 4214 3620 4220 3621
rect 4214 3616 4215 3620
rect 4219 3616 4220 3620
rect 4214 3615 4220 3616
rect 4398 3620 4404 3621
rect 4398 3616 4399 3620
rect 4403 3616 4404 3620
rect 4398 3615 4404 3616
rect 4606 3620 4612 3621
rect 4606 3616 4607 3620
rect 4611 3616 4612 3620
rect 4606 3615 4612 3616
rect 4830 3620 4836 3621
rect 4830 3616 4831 3620
rect 4835 3616 4836 3620
rect 4830 3615 4836 3616
rect 5070 3620 5076 3621
rect 5070 3616 5071 3620
rect 5075 3616 5076 3620
rect 5070 3615 5076 3616
rect 5318 3620 5324 3621
rect 5318 3616 5319 3620
rect 5323 3616 5324 3620
rect 5318 3615 5324 3616
rect 5542 3620 5548 3621
rect 5542 3616 5543 3620
rect 5547 3616 5548 3620
rect 5662 3617 5663 3621
rect 5667 3617 5668 3621
rect 5662 3616 5668 3617
rect 5542 3615 5548 3616
rect 1670 3614 1676 3615
rect 1389 3608 1482 3610
rect 1582 3611 1588 3612
rect 242 3606 248 3607
rect 362 3607 368 3608
rect 362 3603 363 3607
rect 367 3603 368 3607
rect 362 3602 368 3603
rect 578 3607 584 3608
rect 578 3603 579 3607
rect 583 3603 584 3607
rect 578 3602 584 3603
rect 810 3607 816 3608
rect 810 3603 811 3607
rect 815 3603 816 3607
rect 810 3602 816 3603
rect 1138 3607 1144 3608
rect 1138 3603 1139 3607
rect 1143 3603 1144 3607
rect 1582 3607 1583 3611
rect 1587 3607 1588 3611
rect 1582 3606 1588 3607
rect 1882 3611 1888 3612
rect 1882 3607 1883 3611
rect 1887 3607 1888 3611
rect 1882 3606 1888 3607
rect 4186 3605 4192 3606
rect 1138 3602 1144 3603
rect 3838 3604 3844 3605
rect 3838 3600 3839 3604
rect 3843 3600 3844 3604
rect 4186 3601 4187 3605
rect 4191 3601 4192 3605
rect 4186 3600 4192 3601
rect 4370 3605 4376 3606
rect 4370 3601 4371 3605
rect 4375 3601 4376 3605
rect 4370 3600 4376 3601
rect 4578 3605 4584 3606
rect 4578 3601 4579 3605
rect 4583 3601 4584 3605
rect 4578 3600 4584 3601
rect 4802 3605 4808 3606
rect 4802 3601 4803 3605
rect 4807 3601 4808 3605
rect 4802 3600 4808 3601
rect 5042 3605 5048 3606
rect 5042 3601 5043 3605
rect 5047 3601 5048 3605
rect 5042 3600 5048 3601
rect 5290 3605 5296 3606
rect 5290 3601 5291 3605
rect 5295 3601 5296 3605
rect 5290 3600 5296 3601
rect 5514 3605 5520 3606
rect 5514 3601 5515 3605
rect 5519 3601 5520 3605
rect 5514 3600 5520 3601
rect 5662 3604 5668 3605
rect 5662 3600 5663 3604
rect 5667 3600 5668 3604
rect 3838 3599 3844 3600
rect 5662 3599 5668 3600
rect 4311 3595 4317 3596
rect 1922 3591 1928 3592
rect 1922 3587 1923 3591
rect 1927 3590 1928 3591
rect 2346 3591 2352 3592
rect 1927 3588 2001 3590
rect 1927 3587 1928 3588
rect 1922 3586 1928 3587
rect 2346 3587 2347 3591
rect 2351 3587 2352 3591
rect 3407 3591 3413 3592
rect 3407 3590 3408 3591
rect 3293 3588 3408 3590
rect 2346 3586 2352 3587
rect 2522 3587 2528 3588
rect 2522 3583 2523 3587
rect 2527 3583 2528 3587
rect 2522 3582 2528 3583
rect 2850 3587 2856 3588
rect 2850 3583 2851 3587
rect 2855 3583 2856 3587
rect 2850 3582 2856 3583
rect 2986 3587 2992 3588
rect 2986 3583 2987 3587
rect 2991 3583 2992 3587
rect 3407 3587 3408 3588
rect 3412 3587 3413 3591
rect 3623 3591 3629 3592
rect 3623 3590 3624 3591
rect 3509 3588 3624 3590
rect 3407 3586 3413 3587
rect 3623 3587 3624 3588
rect 3628 3587 3629 3591
rect 4311 3591 4312 3595
rect 4316 3594 4317 3595
rect 4326 3595 4332 3596
rect 4326 3594 4327 3595
rect 4316 3592 4327 3594
rect 4316 3591 4317 3592
rect 4311 3590 4317 3591
rect 4326 3591 4327 3592
rect 4331 3591 4332 3595
rect 4326 3590 4332 3591
rect 4495 3595 4501 3596
rect 4495 3591 4496 3595
rect 4500 3594 4501 3595
rect 4538 3595 4544 3596
rect 4538 3594 4539 3595
rect 4500 3592 4539 3594
rect 4500 3591 4501 3592
rect 4495 3590 4501 3591
rect 4538 3591 4539 3592
rect 4543 3591 4544 3595
rect 4538 3590 4544 3591
rect 4703 3595 4712 3596
rect 4703 3591 4704 3595
rect 4711 3591 4712 3595
rect 4703 3590 4712 3591
rect 4927 3595 4936 3596
rect 4927 3591 4928 3595
rect 4935 3591 4936 3595
rect 5167 3595 5173 3596
rect 5167 3594 5168 3595
rect 4927 3590 4936 3591
rect 4940 3592 5168 3594
rect 3623 3586 3629 3587
rect 3634 3587 3640 3588
rect 2986 3582 2992 3583
rect 3634 3583 3635 3587
rect 3639 3583 3640 3587
rect 3634 3582 3640 3583
rect 4626 3587 4632 3588
rect 4626 3583 4627 3587
rect 4631 3586 4632 3587
rect 4940 3586 4942 3592
rect 5167 3591 5168 3592
rect 5172 3591 5173 3595
rect 5167 3590 5173 3591
rect 5346 3595 5352 3596
rect 5346 3591 5347 3595
rect 5351 3594 5352 3595
rect 5415 3595 5421 3596
rect 5415 3594 5416 3595
rect 5351 3592 5416 3594
rect 5351 3591 5352 3592
rect 5346 3590 5352 3591
rect 5415 3591 5416 3592
rect 5420 3591 5421 3595
rect 5415 3590 5421 3591
rect 5610 3595 5616 3596
rect 5610 3591 5611 3595
rect 5615 3594 5616 3595
rect 5639 3595 5645 3596
rect 5639 3594 5640 3595
rect 5615 3592 5640 3594
rect 5615 3591 5616 3592
rect 5610 3590 5616 3591
rect 5639 3591 5640 3592
rect 5644 3591 5645 3595
rect 5639 3590 5645 3591
rect 4631 3584 4942 3586
rect 4631 3583 4632 3584
rect 4626 3582 4632 3583
rect 271 3567 277 3568
rect 271 3563 272 3567
rect 276 3566 277 3567
rect 362 3567 368 3568
rect 362 3566 363 3567
rect 276 3564 363 3566
rect 276 3563 277 3564
rect 271 3562 277 3563
rect 362 3563 363 3564
rect 367 3563 368 3567
rect 362 3562 368 3563
rect 479 3567 485 3568
rect 479 3563 480 3567
rect 484 3566 485 3567
rect 578 3567 584 3568
rect 578 3566 579 3567
rect 484 3564 579 3566
rect 484 3563 485 3564
rect 479 3562 485 3563
rect 578 3563 579 3564
rect 583 3563 584 3567
rect 578 3562 584 3563
rect 695 3567 701 3568
rect 695 3563 696 3567
rect 700 3566 701 3567
rect 810 3567 816 3568
rect 810 3566 811 3567
rect 700 3564 811 3566
rect 700 3563 701 3564
rect 695 3562 701 3563
rect 810 3563 811 3564
rect 815 3563 816 3567
rect 810 3562 816 3563
rect 926 3567 933 3568
rect 926 3563 927 3567
rect 932 3563 933 3567
rect 926 3562 933 3563
rect 1122 3567 1128 3568
rect 1122 3563 1123 3567
rect 1127 3566 1128 3567
rect 1167 3567 1173 3568
rect 1167 3566 1168 3567
rect 1127 3564 1168 3566
rect 1127 3563 1128 3564
rect 1122 3562 1128 3563
rect 1167 3563 1168 3564
rect 1172 3563 1173 3567
rect 1167 3562 1173 3563
rect 1414 3567 1421 3568
rect 1414 3563 1415 3567
rect 1420 3563 1421 3567
rect 1414 3562 1421 3563
rect 1670 3567 1677 3568
rect 1670 3563 1671 3567
rect 1676 3563 1677 3567
rect 1670 3562 1677 3563
rect 1911 3567 1917 3568
rect 1911 3563 1912 3567
rect 1916 3566 1917 3567
rect 1922 3567 1928 3568
rect 1922 3566 1923 3567
rect 1916 3564 1923 3566
rect 1916 3563 1917 3564
rect 1911 3562 1917 3563
rect 1922 3563 1923 3564
rect 1927 3563 1928 3567
rect 1922 3562 1928 3563
rect 110 3560 116 3561
rect 1934 3560 1940 3561
rect 110 3556 111 3560
rect 115 3556 116 3560
rect 110 3555 116 3556
rect 146 3559 152 3560
rect 146 3555 147 3559
rect 151 3555 152 3559
rect 146 3554 152 3555
rect 354 3559 360 3560
rect 354 3555 355 3559
rect 359 3555 360 3559
rect 354 3554 360 3555
rect 570 3559 576 3560
rect 570 3555 571 3559
rect 575 3555 576 3559
rect 570 3554 576 3555
rect 802 3559 808 3560
rect 802 3555 803 3559
rect 807 3555 808 3559
rect 802 3554 808 3555
rect 1042 3559 1048 3560
rect 1042 3555 1043 3559
rect 1047 3555 1048 3559
rect 1042 3554 1048 3555
rect 1290 3559 1296 3560
rect 1290 3555 1291 3559
rect 1295 3555 1296 3559
rect 1290 3554 1296 3555
rect 1546 3559 1552 3560
rect 1546 3555 1547 3559
rect 1551 3555 1552 3559
rect 1546 3554 1552 3555
rect 1786 3559 1792 3560
rect 1786 3555 1787 3559
rect 1791 3555 1792 3559
rect 1934 3556 1935 3560
rect 1939 3556 1940 3560
rect 1934 3555 1940 3556
rect 2850 3555 2856 3556
rect 1786 3554 1792 3555
rect 2850 3551 2851 3555
rect 2855 3554 2856 3555
rect 4326 3555 4332 3556
rect 2855 3552 3206 3554
rect 2855 3551 2856 3552
rect 2850 3550 2856 3551
rect 2090 3547 2096 3548
rect 174 3544 180 3545
rect 110 3543 116 3544
rect 110 3539 111 3543
rect 115 3539 116 3543
rect 174 3540 175 3544
rect 179 3540 180 3544
rect 174 3539 180 3540
rect 382 3544 388 3545
rect 382 3540 383 3544
rect 387 3540 388 3544
rect 382 3539 388 3540
rect 598 3544 604 3545
rect 598 3540 599 3544
rect 603 3540 604 3544
rect 598 3539 604 3540
rect 830 3544 836 3545
rect 830 3540 831 3544
rect 835 3540 836 3544
rect 830 3539 836 3540
rect 1070 3544 1076 3545
rect 1070 3540 1071 3544
rect 1075 3540 1076 3544
rect 1070 3539 1076 3540
rect 1318 3544 1324 3545
rect 1318 3540 1319 3544
rect 1323 3540 1324 3544
rect 1318 3539 1324 3540
rect 1574 3544 1580 3545
rect 1574 3540 1575 3544
rect 1579 3540 1580 3544
rect 1574 3539 1580 3540
rect 1814 3544 1820 3545
rect 1814 3540 1815 3544
rect 1819 3540 1820 3544
rect 1814 3539 1820 3540
rect 1934 3543 1940 3544
rect 1934 3539 1935 3543
rect 1939 3539 1940 3543
rect 2090 3543 2091 3547
rect 2095 3546 2096 3547
rect 2119 3547 2125 3548
rect 2119 3546 2120 3547
rect 2095 3544 2120 3546
rect 2095 3543 2096 3544
rect 2090 3542 2096 3543
rect 2119 3543 2120 3544
rect 2124 3543 2125 3547
rect 2119 3542 2125 3543
rect 2375 3547 2381 3548
rect 2375 3543 2376 3547
rect 2380 3546 2381 3547
rect 2522 3547 2528 3548
rect 2522 3546 2523 3547
rect 2380 3544 2523 3546
rect 2380 3543 2381 3544
rect 2375 3542 2381 3543
rect 2522 3543 2523 3544
rect 2527 3543 2528 3547
rect 2522 3542 2528 3543
rect 2638 3547 2645 3548
rect 2638 3543 2639 3547
rect 2644 3543 2645 3547
rect 2638 3542 2645 3543
rect 2879 3547 2885 3548
rect 2879 3543 2880 3547
rect 2884 3546 2885 3547
rect 2986 3547 2992 3548
rect 2986 3546 2987 3547
rect 2884 3544 2987 3546
rect 2884 3543 2885 3544
rect 2879 3542 2885 3543
rect 2986 3543 2987 3544
rect 2991 3543 2992 3547
rect 2986 3542 2992 3543
rect 3102 3547 3109 3548
rect 3102 3543 3103 3547
rect 3108 3543 3109 3547
rect 3204 3546 3206 3552
rect 3319 3547 3325 3548
rect 3319 3546 3320 3547
rect 3204 3544 3320 3546
rect 3102 3542 3109 3543
rect 3319 3543 3320 3544
rect 3324 3543 3325 3547
rect 3319 3542 3325 3543
rect 3407 3547 3413 3548
rect 3407 3543 3408 3547
rect 3412 3546 3413 3547
rect 3535 3547 3541 3548
rect 3535 3546 3536 3547
rect 3412 3544 3536 3546
rect 3412 3543 3413 3544
rect 3407 3542 3413 3543
rect 3535 3543 3536 3544
rect 3540 3543 3541 3547
rect 3535 3542 3541 3543
rect 3623 3547 3629 3548
rect 3623 3543 3624 3547
rect 3628 3546 3629 3547
rect 3751 3547 3757 3548
rect 3751 3546 3752 3547
rect 3628 3544 3752 3546
rect 3628 3543 3629 3544
rect 3623 3542 3629 3543
rect 3751 3543 3752 3544
rect 3756 3543 3757 3547
rect 4284 3546 4286 3553
rect 4326 3551 4327 3555
rect 4331 3554 4332 3555
rect 4538 3555 4544 3556
rect 4331 3552 4377 3554
rect 4331 3551 4332 3552
rect 4326 3550 4332 3551
rect 4538 3551 4539 3555
rect 4543 3554 4544 3555
rect 4706 3555 4712 3556
rect 4543 3552 4585 3554
rect 4543 3551 4544 3552
rect 4538 3550 4544 3551
rect 4706 3551 4707 3555
rect 4711 3554 4712 3555
rect 4930 3555 4936 3556
rect 4711 3552 4809 3554
rect 4711 3551 4712 3552
rect 4706 3550 4712 3551
rect 4930 3551 4931 3555
rect 4935 3554 4936 3555
rect 5386 3555 5392 3556
rect 4935 3552 5049 3554
rect 4935 3551 4936 3552
rect 4930 3550 4936 3551
rect 5386 3551 5387 3555
rect 5391 3551 5392 3555
rect 5626 3555 5632 3556
rect 5626 3554 5627 3555
rect 5613 3552 5627 3554
rect 5386 3550 5392 3551
rect 5626 3551 5627 3552
rect 5631 3551 5632 3555
rect 5626 3550 5632 3551
rect 4814 3547 4820 3548
rect 4814 3546 4815 3547
rect 4284 3544 4815 3546
rect 3751 3542 3757 3543
rect 4814 3543 4815 3544
rect 4819 3543 4820 3547
rect 4814 3542 4820 3543
rect 110 3538 116 3539
rect 1934 3538 1940 3539
rect 1974 3540 1980 3541
rect 3798 3540 3804 3541
rect 1974 3536 1975 3540
rect 1979 3536 1980 3540
rect 1974 3535 1980 3536
rect 1994 3539 2000 3540
rect 1994 3535 1995 3539
rect 1999 3535 2000 3539
rect 1994 3534 2000 3535
rect 2250 3539 2256 3540
rect 2250 3535 2251 3539
rect 2255 3535 2256 3539
rect 2250 3534 2256 3535
rect 2514 3539 2520 3540
rect 2514 3535 2515 3539
rect 2519 3535 2520 3539
rect 2514 3534 2520 3535
rect 2754 3539 2760 3540
rect 2754 3535 2755 3539
rect 2759 3535 2760 3539
rect 2754 3534 2760 3535
rect 2978 3539 2984 3540
rect 2978 3535 2979 3539
rect 2983 3535 2984 3539
rect 2978 3534 2984 3535
rect 3194 3539 3200 3540
rect 3194 3535 3195 3539
rect 3199 3535 3200 3539
rect 3194 3534 3200 3535
rect 3410 3539 3416 3540
rect 3410 3535 3411 3539
rect 3415 3535 3416 3539
rect 3410 3534 3416 3535
rect 3626 3539 3632 3540
rect 3626 3535 3627 3539
rect 3631 3535 3632 3539
rect 3798 3536 3799 3540
rect 3803 3536 3804 3540
rect 3798 3535 3804 3536
rect 3626 3534 3632 3535
rect 2022 3524 2028 3525
rect 1974 3523 1980 3524
rect 1974 3519 1975 3523
rect 1979 3519 1980 3523
rect 2022 3520 2023 3524
rect 2027 3520 2028 3524
rect 2022 3519 2028 3520
rect 2278 3524 2284 3525
rect 2278 3520 2279 3524
rect 2283 3520 2284 3524
rect 2278 3519 2284 3520
rect 2542 3524 2548 3525
rect 2542 3520 2543 3524
rect 2547 3520 2548 3524
rect 2542 3519 2548 3520
rect 2782 3524 2788 3525
rect 2782 3520 2783 3524
rect 2787 3520 2788 3524
rect 2782 3519 2788 3520
rect 3006 3524 3012 3525
rect 3006 3520 3007 3524
rect 3011 3520 3012 3524
rect 3006 3519 3012 3520
rect 3222 3524 3228 3525
rect 3222 3520 3223 3524
rect 3227 3520 3228 3524
rect 3222 3519 3228 3520
rect 3438 3524 3444 3525
rect 3438 3520 3439 3524
rect 3443 3520 3444 3524
rect 3438 3519 3444 3520
rect 3654 3524 3660 3525
rect 3654 3520 3655 3524
rect 3659 3520 3660 3524
rect 3654 3519 3660 3520
rect 3798 3523 3804 3524
rect 3798 3519 3799 3523
rect 3803 3519 3804 3523
rect 1974 3518 1980 3519
rect 3798 3518 3804 3519
rect 4626 3499 4632 3500
rect 4626 3495 4627 3499
rect 4631 3495 4632 3499
rect 5318 3499 5324 3500
rect 4626 3494 4632 3495
rect 4690 3495 4696 3496
rect 4690 3491 4691 3495
rect 4695 3491 4696 3495
rect 4690 3490 4696 3491
rect 4850 3495 4856 3496
rect 4850 3491 4851 3495
rect 4855 3491 4856 3495
rect 4850 3490 4856 3491
rect 5010 3495 5016 3496
rect 5010 3491 5011 3495
rect 5015 3491 5016 3495
rect 5010 3490 5016 3491
rect 5178 3495 5184 3496
rect 5178 3491 5179 3495
rect 5183 3491 5184 3495
rect 5318 3495 5319 3499
rect 5323 3498 5324 3499
rect 5610 3499 5616 3500
rect 5323 3496 5353 3498
rect 5323 3495 5324 3496
rect 5318 3494 5324 3495
rect 5610 3495 5611 3499
rect 5615 3495 5616 3499
rect 5610 3494 5616 3495
rect 5178 3490 5184 3491
rect 110 3461 116 3462
rect 1934 3461 1940 3462
rect 110 3457 111 3461
rect 115 3457 116 3461
rect 110 3456 116 3457
rect 302 3460 308 3461
rect 302 3456 303 3460
rect 307 3456 308 3460
rect 302 3455 308 3456
rect 446 3460 452 3461
rect 446 3456 447 3460
rect 451 3456 452 3460
rect 446 3455 452 3456
rect 598 3460 604 3461
rect 598 3456 599 3460
rect 603 3456 604 3460
rect 598 3455 604 3456
rect 758 3460 764 3461
rect 758 3456 759 3460
rect 763 3456 764 3460
rect 758 3455 764 3456
rect 934 3460 940 3461
rect 934 3456 935 3460
rect 939 3456 940 3460
rect 934 3455 940 3456
rect 1110 3460 1116 3461
rect 1110 3456 1111 3460
rect 1115 3456 1116 3460
rect 1110 3455 1116 3456
rect 1294 3460 1300 3461
rect 1294 3456 1295 3460
rect 1299 3456 1300 3460
rect 1294 3455 1300 3456
rect 1486 3460 1492 3461
rect 1486 3456 1487 3460
rect 1491 3456 1492 3460
rect 1934 3457 1935 3461
rect 1939 3457 1940 3461
rect 1934 3456 1940 3457
rect 1974 3457 1980 3458
rect 3798 3457 3804 3458
rect 1486 3455 1492 3456
rect 1974 3453 1975 3457
rect 1979 3453 1980 3457
rect 1974 3452 1980 3453
rect 2022 3456 2028 3457
rect 2022 3452 2023 3456
rect 2027 3452 2028 3456
rect 2022 3451 2028 3452
rect 2190 3456 2196 3457
rect 2190 3452 2191 3456
rect 2195 3452 2196 3456
rect 2190 3451 2196 3452
rect 2398 3456 2404 3457
rect 2398 3452 2399 3456
rect 2403 3452 2404 3456
rect 2398 3451 2404 3452
rect 2614 3456 2620 3457
rect 2614 3452 2615 3456
rect 2619 3452 2620 3456
rect 2614 3451 2620 3452
rect 2830 3456 2836 3457
rect 2830 3452 2831 3456
rect 2835 3452 2836 3456
rect 2830 3451 2836 3452
rect 3046 3456 3052 3457
rect 3046 3452 3047 3456
rect 3051 3452 3052 3456
rect 3046 3451 3052 3452
rect 3262 3456 3268 3457
rect 3262 3452 3263 3456
rect 3267 3452 3268 3456
rect 3262 3451 3268 3452
rect 3478 3456 3484 3457
rect 3478 3452 3479 3456
rect 3483 3452 3484 3456
rect 3478 3451 3484 3452
rect 3678 3456 3684 3457
rect 3678 3452 3679 3456
rect 3683 3452 3684 3456
rect 3798 3453 3799 3457
rect 3803 3453 3804 3457
rect 3798 3452 3804 3453
rect 4655 3455 4661 3456
rect 3678 3451 3684 3452
rect 4655 3451 4656 3455
rect 4660 3454 4661 3455
rect 4690 3455 4696 3456
rect 4690 3454 4691 3455
rect 4660 3452 4691 3454
rect 4660 3451 4661 3452
rect 4655 3450 4661 3451
rect 4690 3451 4691 3452
rect 4695 3451 4696 3455
rect 4690 3450 4696 3451
rect 4807 3455 4813 3456
rect 4807 3451 4808 3455
rect 4812 3454 4813 3455
rect 4850 3455 4856 3456
rect 4850 3454 4851 3455
rect 4812 3452 4851 3454
rect 4812 3451 4813 3452
rect 4807 3450 4813 3451
rect 4850 3451 4851 3452
rect 4855 3451 4856 3455
rect 4850 3450 4856 3451
rect 4967 3455 4973 3456
rect 4967 3451 4968 3455
rect 4972 3454 4973 3455
rect 5010 3455 5016 3456
rect 5010 3454 5011 3455
rect 4972 3452 5011 3454
rect 4972 3451 4973 3452
rect 4967 3450 4973 3451
rect 5010 3451 5011 3452
rect 5015 3451 5016 3455
rect 5010 3450 5016 3451
rect 5127 3455 5133 3456
rect 5127 3451 5128 3455
rect 5132 3454 5133 3455
rect 5178 3455 5184 3456
rect 5178 3454 5179 3455
rect 5132 3452 5179 3454
rect 5132 3451 5133 3452
rect 5127 3450 5133 3451
rect 5178 3451 5179 3452
rect 5183 3451 5184 3455
rect 5178 3450 5184 3451
rect 5238 3455 5244 3456
rect 5238 3451 5239 3455
rect 5243 3454 5244 3455
rect 5295 3455 5301 3456
rect 5295 3454 5296 3455
rect 5243 3452 5296 3454
rect 5243 3451 5244 3452
rect 5238 3450 5244 3451
rect 5295 3451 5296 3452
rect 5300 3451 5301 3455
rect 5295 3450 5301 3451
rect 5386 3455 5392 3456
rect 5386 3451 5387 3455
rect 5391 3454 5392 3455
rect 5471 3455 5477 3456
rect 5471 3454 5472 3455
rect 5391 3452 5472 3454
rect 5391 3451 5392 3452
rect 5386 3450 5392 3451
rect 5471 3451 5472 3452
rect 5476 3451 5477 3455
rect 5471 3450 5477 3451
rect 5638 3455 5645 3456
rect 5638 3451 5639 3455
rect 5644 3451 5645 3455
rect 5638 3450 5645 3451
rect 3838 3448 3844 3449
rect 5662 3448 5668 3449
rect 274 3445 280 3446
rect 110 3444 116 3445
rect 110 3440 111 3444
rect 115 3440 116 3444
rect 274 3441 275 3445
rect 279 3441 280 3445
rect 274 3440 280 3441
rect 418 3445 424 3446
rect 418 3441 419 3445
rect 423 3441 424 3445
rect 418 3440 424 3441
rect 570 3445 576 3446
rect 570 3441 571 3445
rect 575 3441 576 3445
rect 570 3440 576 3441
rect 730 3445 736 3446
rect 730 3441 731 3445
rect 735 3441 736 3445
rect 730 3440 736 3441
rect 906 3445 912 3446
rect 906 3441 907 3445
rect 911 3441 912 3445
rect 906 3440 912 3441
rect 1082 3445 1088 3446
rect 1082 3441 1083 3445
rect 1087 3441 1088 3445
rect 1082 3440 1088 3441
rect 1266 3445 1272 3446
rect 1266 3441 1267 3445
rect 1271 3441 1272 3445
rect 1266 3440 1272 3441
rect 1458 3445 1464 3446
rect 1458 3441 1459 3445
rect 1463 3441 1464 3445
rect 1458 3440 1464 3441
rect 1934 3444 1940 3445
rect 1934 3440 1935 3444
rect 1939 3440 1940 3444
rect 3838 3444 3839 3448
rect 3843 3444 3844 3448
rect 3838 3443 3844 3444
rect 4530 3447 4536 3448
rect 4530 3443 4531 3447
rect 4535 3443 4536 3447
rect 4530 3442 4536 3443
rect 4682 3447 4688 3448
rect 4682 3443 4683 3447
rect 4687 3443 4688 3447
rect 4682 3442 4688 3443
rect 4842 3447 4848 3448
rect 4842 3443 4843 3447
rect 4847 3443 4848 3447
rect 4842 3442 4848 3443
rect 5002 3447 5008 3448
rect 5002 3443 5003 3447
rect 5007 3443 5008 3447
rect 5002 3442 5008 3443
rect 5170 3447 5176 3448
rect 5170 3443 5171 3447
rect 5175 3443 5176 3447
rect 5170 3442 5176 3443
rect 5346 3447 5352 3448
rect 5346 3443 5347 3447
rect 5351 3443 5352 3447
rect 5346 3442 5352 3443
rect 5514 3447 5520 3448
rect 5514 3443 5515 3447
rect 5519 3443 5520 3447
rect 5662 3444 5663 3448
rect 5667 3444 5668 3448
rect 5662 3443 5668 3444
rect 5514 3442 5520 3443
rect 1994 3441 2000 3442
rect 110 3439 116 3440
rect 1934 3439 1940 3440
rect 1974 3440 1980 3441
rect 1974 3436 1975 3440
rect 1979 3436 1980 3440
rect 1994 3437 1995 3441
rect 1999 3437 2000 3441
rect 1994 3436 2000 3437
rect 2162 3441 2168 3442
rect 2162 3437 2163 3441
rect 2167 3437 2168 3441
rect 2162 3436 2168 3437
rect 2370 3441 2376 3442
rect 2370 3437 2371 3441
rect 2375 3437 2376 3441
rect 2370 3436 2376 3437
rect 2586 3441 2592 3442
rect 2586 3437 2587 3441
rect 2591 3437 2592 3441
rect 2586 3436 2592 3437
rect 2802 3441 2808 3442
rect 2802 3437 2803 3441
rect 2807 3437 2808 3441
rect 2802 3436 2808 3437
rect 3018 3441 3024 3442
rect 3018 3437 3019 3441
rect 3023 3437 3024 3441
rect 3018 3436 3024 3437
rect 3234 3441 3240 3442
rect 3234 3437 3235 3441
rect 3239 3437 3240 3441
rect 3234 3436 3240 3437
rect 3450 3441 3456 3442
rect 3450 3437 3451 3441
rect 3455 3437 3456 3441
rect 3450 3436 3456 3437
rect 3650 3441 3656 3442
rect 3650 3437 3651 3441
rect 3655 3437 3656 3441
rect 3650 3436 3656 3437
rect 3798 3440 3804 3441
rect 3798 3436 3799 3440
rect 3803 3436 3804 3440
rect 399 3435 408 3436
rect 399 3431 400 3435
rect 407 3431 408 3435
rect 399 3430 408 3431
rect 543 3435 552 3436
rect 543 3431 544 3435
rect 551 3431 552 3435
rect 543 3430 552 3431
rect 695 3435 701 3436
rect 695 3431 696 3435
rect 700 3434 701 3435
rect 718 3435 724 3436
rect 718 3434 719 3435
rect 700 3432 719 3434
rect 700 3431 701 3432
rect 695 3430 701 3431
rect 718 3431 719 3432
rect 723 3431 724 3435
rect 718 3430 724 3431
rect 762 3435 768 3436
rect 762 3431 763 3435
rect 767 3434 768 3435
rect 855 3435 861 3436
rect 855 3434 856 3435
rect 767 3432 856 3434
rect 767 3431 768 3432
rect 762 3430 768 3431
rect 855 3431 856 3432
rect 860 3431 861 3435
rect 855 3430 861 3431
rect 1031 3435 1040 3436
rect 1031 3431 1032 3435
rect 1039 3431 1040 3435
rect 1031 3430 1040 3431
rect 1138 3435 1144 3436
rect 1138 3431 1139 3435
rect 1143 3434 1144 3435
rect 1207 3435 1213 3436
rect 1207 3434 1208 3435
rect 1143 3432 1208 3434
rect 1143 3431 1144 3432
rect 1138 3430 1144 3431
rect 1207 3431 1208 3432
rect 1212 3431 1213 3435
rect 1207 3430 1213 3431
rect 1391 3435 1400 3436
rect 1391 3431 1392 3435
rect 1399 3431 1400 3435
rect 1391 3430 1400 3431
rect 1582 3435 1589 3436
rect 1974 3435 1980 3436
rect 3798 3435 3804 3436
rect 1582 3431 1583 3435
rect 1588 3431 1589 3435
rect 4558 3432 4564 3433
rect 1582 3430 1589 3431
rect 2119 3431 2128 3432
rect 2119 3427 2120 3431
rect 2127 3427 2128 3431
rect 2119 3426 2128 3427
rect 2287 3431 2293 3432
rect 2287 3427 2288 3431
rect 2292 3430 2293 3431
rect 2334 3431 2340 3432
rect 2334 3430 2335 3431
rect 2292 3428 2335 3430
rect 2292 3427 2293 3428
rect 2287 3426 2293 3427
rect 2334 3427 2335 3428
rect 2339 3427 2340 3431
rect 2334 3426 2340 3427
rect 2346 3431 2352 3432
rect 2346 3427 2347 3431
rect 2351 3430 2352 3431
rect 2495 3431 2501 3432
rect 2495 3430 2496 3431
rect 2351 3428 2496 3430
rect 2351 3427 2352 3428
rect 2346 3426 2352 3427
rect 2495 3427 2496 3428
rect 2500 3427 2501 3431
rect 2495 3426 2501 3427
rect 2711 3431 2717 3432
rect 2711 3427 2712 3431
rect 2716 3430 2717 3431
rect 2743 3431 2749 3432
rect 2743 3430 2744 3431
rect 2716 3428 2744 3430
rect 2716 3427 2717 3428
rect 2711 3426 2717 3427
rect 2743 3427 2744 3428
rect 2748 3427 2749 3431
rect 2743 3426 2749 3427
rect 2799 3431 2805 3432
rect 2799 3427 2800 3431
rect 2804 3430 2805 3431
rect 2927 3431 2933 3432
rect 2927 3430 2928 3431
rect 2804 3428 2928 3430
rect 2804 3427 2805 3428
rect 2799 3426 2805 3427
rect 2927 3427 2928 3428
rect 2932 3427 2933 3431
rect 2927 3426 2933 3427
rect 3143 3431 3152 3432
rect 3143 3427 3144 3431
rect 3151 3427 3152 3431
rect 3143 3426 3152 3427
rect 3359 3431 3368 3432
rect 3359 3427 3360 3431
rect 3367 3427 3368 3431
rect 3359 3426 3368 3427
rect 3575 3431 3581 3432
rect 3575 3427 3576 3431
rect 3580 3430 3581 3431
rect 3634 3431 3640 3432
rect 3634 3430 3635 3431
rect 3580 3428 3635 3430
rect 3580 3427 3581 3428
rect 3575 3426 3581 3427
rect 3634 3427 3635 3428
rect 3639 3427 3640 3431
rect 3634 3426 3640 3427
rect 3690 3431 3696 3432
rect 3690 3427 3691 3431
rect 3695 3430 3696 3431
rect 3775 3431 3781 3432
rect 3775 3430 3776 3431
rect 3695 3428 3776 3430
rect 3695 3427 3696 3428
rect 3690 3426 3696 3427
rect 3775 3427 3776 3428
rect 3780 3427 3781 3431
rect 3775 3426 3781 3427
rect 3838 3431 3844 3432
rect 3838 3427 3839 3431
rect 3843 3427 3844 3431
rect 4558 3428 4559 3432
rect 4563 3428 4564 3432
rect 4558 3427 4564 3428
rect 4710 3432 4716 3433
rect 4710 3428 4711 3432
rect 4715 3428 4716 3432
rect 4710 3427 4716 3428
rect 4870 3432 4876 3433
rect 4870 3428 4871 3432
rect 4875 3428 4876 3432
rect 4870 3427 4876 3428
rect 5030 3432 5036 3433
rect 5030 3428 5031 3432
rect 5035 3428 5036 3432
rect 5030 3427 5036 3428
rect 5198 3432 5204 3433
rect 5198 3428 5199 3432
rect 5203 3428 5204 3432
rect 5198 3427 5204 3428
rect 5374 3432 5380 3433
rect 5374 3428 5375 3432
rect 5379 3428 5380 3432
rect 5374 3427 5380 3428
rect 5542 3432 5548 3433
rect 5542 3428 5543 3432
rect 5547 3428 5548 3432
rect 5542 3427 5548 3428
rect 5662 3431 5668 3432
rect 5662 3427 5663 3431
rect 5667 3427 5668 3431
rect 3838 3426 3844 3427
rect 5662 3426 5668 3427
rect 402 3395 408 3396
rect 372 3386 374 3393
rect 402 3391 403 3395
rect 407 3394 408 3395
rect 546 3395 552 3396
rect 407 3392 425 3394
rect 407 3391 408 3392
rect 402 3390 408 3391
rect 546 3391 547 3395
rect 551 3394 552 3395
rect 718 3395 724 3396
rect 551 3392 577 3394
rect 551 3391 552 3392
rect 546 3390 552 3391
rect 718 3391 719 3395
rect 723 3394 724 3395
rect 834 3395 840 3396
rect 723 3392 737 3394
rect 723 3391 724 3392
rect 718 3390 724 3391
rect 834 3391 835 3395
rect 839 3394 840 3395
rect 1034 3395 1040 3396
rect 839 3392 913 3394
rect 839 3391 840 3392
rect 834 3390 840 3391
rect 1034 3391 1035 3395
rect 1039 3394 1040 3395
rect 1362 3395 1368 3396
rect 1039 3392 1089 3394
rect 1039 3391 1040 3392
rect 1034 3390 1040 3391
rect 1362 3391 1363 3395
rect 1367 3391 1368 3395
rect 1362 3390 1368 3391
rect 1394 3395 1400 3396
rect 1394 3391 1395 3395
rect 1399 3394 1400 3395
rect 1399 3392 1465 3394
rect 1399 3391 1400 3392
rect 1394 3390 1400 3391
rect 2090 3391 2096 3392
rect 926 3387 932 3388
rect 926 3386 927 3387
rect 372 3384 927 3386
rect 926 3383 927 3384
rect 931 3383 932 3387
rect 2090 3387 2091 3391
rect 2095 3387 2096 3391
rect 2090 3386 2096 3387
rect 2122 3391 2128 3392
rect 2122 3387 2123 3391
rect 2127 3390 2128 3391
rect 2334 3391 2340 3392
rect 2127 3388 2169 3390
rect 2127 3387 2128 3388
rect 2122 3386 2128 3387
rect 2334 3387 2335 3391
rect 2339 3390 2340 3391
rect 2638 3391 2644 3392
rect 2339 3388 2377 3390
rect 2339 3387 2340 3388
rect 2334 3386 2340 3387
rect 2638 3387 2639 3391
rect 2643 3387 2644 3391
rect 2638 3386 2644 3387
rect 2743 3391 2749 3392
rect 2743 3387 2744 3391
rect 2748 3390 2749 3391
rect 3146 3391 3152 3392
rect 2748 3388 2809 3390
rect 2748 3387 2749 3388
rect 2743 3386 2749 3387
rect 926 3382 932 3383
rect 3116 3374 3118 3389
rect 3146 3387 3147 3391
rect 3151 3390 3152 3391
rect 3362 3391 3368 3392
rect 3151 3388 3241 3390
rect 3151 3387 3152 3388
rect 3146 3386 3152 3387
rect 3362 3387 3363 3391
rect 3367 3390 3368 3391
rect 3746 3391 3752 3392
rect 3367 3388 3457 3390
rect 3367 3387 3368 3388
rect 3362 3386 3368 3387
rect 3746 3387 3747 3391
rect 3751 3387 3752 3391
rect 3746 3386 3752 3387
rect 3690 3375 3696 3376
rect 3690 3374 3691 3375
rect 3116 3372 3691 3374
rect 3690 3371 3691 3372
rect 3695 3371 3696 3375
rect 3690 3370 3696 3371
rect 3838 3369 3844 3370
rect 5662 3369 5668 3370
rect 3838 3365 3839 3369
rect 3843 3365 3844 3369
rect 3838 3364 3844 3365
rect 3886 3368 3892 3369
rect 3886 3364 3887 3368
rect 3891 3364 3892 3368
rect 3886 3363 3892 3364
rect 4150 3368 4156 3369
rect 4150 3364 4151 3368
rect 4155 3364 4156 3368
rect 4150 3363 4156 3364
rect 4422 3368 4428 3369
rect 4422 3364 4423 3368
rect 4427 3364 4428 3368
rect 4422 3363 4428 3364
rect 4670 3368 4676 3369
rect 4670 3364 4671 3368
rect 4675 3364 4676 3368
rect 4670 3363 4676 3364
rect 4894 3368 4900 3369
rect 4894 3364 4895 3368
rect 4899 3364 4900 3368
rect 4894 3363 4900 3364
rect 5110 3368 5116 3369
rect 5110 3364 5111 3368
rect 5115 3364 5116 3368
rect 5110 3363 5116 3364
rect 5326 3368 5332 3369
rect 5326 3364 5327 3368
rect 5331 3364 5332 3368
rect 5326 3363 5332 3364
rect 5542 3368 5548 3369
rect 5542 3364 5543 3368
rect 5547 3364 5548 3368
rect 5662 3365 5663 3369
rect 5667 3365 5668 3369
rect 5662 3364 5668 3365
rect 5542 3363 5548 3364
rect 3858 3353 3864 3354
rect 3838 3352 3844 3353
rect 3838 3348 3839 3352
rect 3843 3348 3844 3352
rect 3858 3349 3859 3353
rect 3863 3349 3864 3353
rect 3858 3348 3864 3349
rect 4122 3353 4128 3354
rect 4122 3349 4123 3353
rect 4127 3349 4128 3353
rect 4122 3348 4128 3349
rect 4394 3353 4400 3354
rect 4394 3349 4395 3353
rect 4399 3349 4400 3353
rect 4394 3348 4400 3349
rect 4642 3353 4648 3354
rect 4642 3349 4643 3353
rect 4647 3349 4648 3353
rect 4642 3348 4648 3349
rect 4866 3353 4872 3354
rect 4866 3349 4867 3353
rect 4871 3349 4872 3353
rect 4866 3348 4872 3349
rect 5082 3353 5088 3354
rect 5082 3349 5083 3353
rect 5087 3349 5088 3353
rect 5082 3348 5088 3349
rect 5298 3353 5304 3354
rect 5298 3349 5299 3353
rect 5303 3349 5304 3353
rect 5298 3348 5304 3349
rect 5514 3353 5520 3354
rect 5514 3349 5515 3353
rect 5519 3349 5520 3353
rect 5514 3348 5520 3349
rect 5662 3352 5668 3353
rect 5662 3348 5663 3352
rect 5667 3348 5668 3352
rect 762 3347 768 3348
rect 562 3343 568 3344
rect 562 3339 563 3343
rect 567 3339 568 3343
rect 762 3343 763 3347
rect 767 3343 768 3347
rect 1390 3347 1396 3348
rect 3838 3347 3844 3348
rect 5662 3347 5668 3348
rect 762 3342 768 3343
rect 882 3343 888 3344
rect 562 3338 568 3339
rect 882 3339 883 3343
rect 887 3339 888 3343
rect 882 3338 888 3339
rect 1098 3343 1104 3344
rect 1098 3339 1099 3343
rect 1103 3339 1104 3343
rect 1390 3343 1391 3347
rect 1395 3343 1396 3347
rect 1390 3342 1396 3343
rect 3746 3343 3752 3344
rect 1098 3338 1104 3339
rect 3746 3339 3747 3343
rect 3751 3342 3752 3343
rect 3983 3343 3989 3344
rect 3983 3342 3984 3343
rect 3751 3340 3984 3342
rect 3751 3339 3752 3340
rect 3746 3338 3752 3339
rect 3983 3339 3984 3340
rect 3988 3339 3989 3343
rect 3983 3338 3989 3339
rect 4130 3343 4136 3344
rect 4130 3339 4131 3343
rect 4135 3342 4136 3343
rect 4247 3343 4253 3344
rect 4247 3342 4248 3343
rect 4135 3340 4248 3342
rect 4135 3339 4136 3340
rect 4130 3338 4136 3339
rect 4247 3339 4248 3340
rect 4252 3339 4253 3343
rect 4247 3338 4253 3339
rect 4519 3343 4528 3344
rect 4519 3339 4520 3343
rect 4527 3339 4528 3343
rect 4519 3338 4528 3339
rect 4767 3343 4776 3344
rect 4767 3339 4768 3343
rect 4775 3339 4776 3343
rect 4767 3338 4776 3339
rect 4991 3343 4997 3344
rect 4991 3339 4992 3343
rect 4996 3342 4997 3343
rect 5039 3343 5045 3344
rect 5039 3342 5040 3343
rect 4996 3340 5040 3342
rect 4996 3339 4997 3340
rect 4991 3338 4997 3339
rect 5039 3339 5040 3340
rect 5044 3339 5045 3343
rect 5039 3338 5045 3339
rect 5207 3343 5213 3344
rect 5207 3339 5208 3343
rect 5212 3342 5213 3343
rect 5254 3343 5260 3344
rect 5254 3342 5255 3343
rect 5212 3340 5255 3342
rect 5212 3339 5213 3340
rect 5207 3338 5213 3339
rect 5254 3339 5255 3340
rect 5259 3339 5260 3343
rect 5423 3343 5429 3344
rect 5423 3342 5424 3343
rect 5254 3338 5260 3339
rect 5299 3340 5424 3342
rect 5142 3335 5148 3336
rect 5142 3331 5143 3335
rect 5147 3334 5148 3335
rect 5299 3334 5301 3340
rect 5423 3339 5424 3340
rect 5428 3339 5429 3343
rect 5423 3338 5429 3339
rect 5610 3343 5616 3344
rect 5610 3339 5611 3343
rect 5615 3342 5616 3343
rect 5639 3343 5645 3344
rect 5639 3342 5640 3343
rect 5615 3340 5640 3342
rect 5615 3339 5616 3340
rect 5610 3338 5616 3339
rect 5639 3339 5640 3340
rect 5644 3339 5645 3343
rect 5639 3338 5645 3339
rect 5147 3332 5301 3334
rect 5147 3331 5148 3332
rect 5142 3330 5148 3331
rect 2799 3323 2805 3324
rect 2799 3322 2800 3323
rect 2620 3320 2800 3322
rect 2186 3319 2192 3320
rect 2186 3318 2187 3319
rect 2093 3316 2187 3318
rect 2186 3315 2187 3316
rect 2191 3315 2192 3319
rect 2346 3319 2352 3320
rect 2346 3318 2347 3319
rect 2293 3316 2347 3318
rect 2186 3314 2192 3315
rect 2346 3315 2347 3316
rect 2351 3315 2352 3319
rect 2620 3318 2622 3320
rect 2799 3319 2800 3320
rect 2804 3319 2805 3323
rect 2799 3318 2805 3319
rect 2509 3316 2622 3318
rect 2346 3314 2352 3315
rect 2626 3315 2632 3316
rect 834 3311 840 3312
rect 834 3310 835 3311
rect 752 3308 835 3310
rect 591 3303 597 3304
rect 591 3299 592 3303
rect 596 3302 597 3303
rect 752 3302 754 3308
rect 834 3307 835 3308
rect 839 3307 840 3311
rect 2626 3311 2627 3315
rect 2631 3311 2632 3315
rect 2626 3310 2632 3311
rect 2906 3315 2912 3316
rect 2906 3311 2907 3315
rect 2911 3311 2912 3315
rect 2906 3310 2912 3311
rect 3010 3315 3016 3316
rect 3010 3311 3011 3315
rect 3015 3311 3016 3315
rect 3010 3310 3016 3311
rect 3194 3315 3200 3316
rect 3194 3311 3195 3315
rect 3199 3311 3200 3315
rect 3194 3310 3200 3311
rect 3378 3315 3384 3316
rect 3378 3311 3379 3315
rect 3383 3311 3384 3315
rect 3378 3310 3384 3311
rect 3562 3315 3568 3316
rect 3562 3311 3563 3315
rect 3567 3311 3568 3315
rect 3562 3310 3568 3311
rect 4130 3311 4136 3312
rect 4130 3310 4131 3311
rect 834 3306 840 3307
rect 3956 3308 4131 3310
rect 596 3300 754 3302
rect 791 3303 797 3304
rect 596 3299 597 3300
rect 591 3298 597 3299
rect 791 3299 792 3303
rect 796 3302 797 3303
rect 882 3303 888 3304
rect 882 3302 883 3303
rect 796 3300 883 3302
rect 796 3299 797 3300
rect 791 3298 797 3299
rect 882 3299 883 3300
rect 887 3299 888 3303
rect 882 3298 888 3299
rect 999 3303 1005 3304
rect 999 3299 1000 3303
rect 1004 3302 1005 3303
rect 1098 3303 1104 3304
rect 1098 3302 1099 3303
rect 1004 3300 1099 3302
rect 1004 3299 1005 3300
rect 999 3298 1005 3299
rect 1098 3299 1099 3300
rect 1103 3299 1104 3303
rect 1098 3298 1104 3299
rect 1154 3303 1160 3304
rect 1154 3299 1155 3303
rect 1159 3302 1160 3303
rect 1215 3303 1221 3304
rect 1215 3302 1216 3303
rect 1159 3300 1216 3302
rect 1159 3299 1160 3300
rect 1154 3298 1160 3299
rect 1215 3299 1216 3300
rect 1220 3299 1221 3303
rect 1215 3298 1221 3299
rect 1362 3303 1368 3304
rect 1362 3299 1363 3303
rect 1367 3302 1368 3303
rect 1439 3303 1445 3304
rect 1439 3302 1440 3303
rect 1367 3300 1440 3302
rect 1367 3299 1368 3300
rect 1362 3298 1368 3299
rect 1439 3299 1440 3300
rect 1444 3299 1445 3303
rect 3956 3301 3958 3308
rect 4130 3307 4131 3308
rect 4135 3307 4136 3311
rect 4130 3306 4136 3307
rect 3986 3303 3992 3304
rect 1439 3298 1445 3299
rect 3986 3299 3987 3303
rect 3991 3302 3992 3303
rect 4522 3303 4528 3304
rect 3991 3300 4129 3302
rect 3991 3299 3992 3300
rect 3986 3298 3992 3299
rect 110 3296 116 3297
rect 1934 3296 1940 3297
rect 110 3292 111 3296
rect 115 3292 116 3296
rect 110 3291 116 3292
rect 466 3295 472 3296
rect 466 3291 467 3295
rect 471 3291 472 3295
rect 466 3290 472 3291
rect 666 3295 672 3296
rect 666 3291 667 3295
rect 671 3291 672 3295
rect 666 3290 672 3291
rect 874 3295 880 3296
rect 874 3291 875 3295
rect 879 3291 880 3295
rect 874 3290 880 3291
rect 1090 3295 1096 3296
rect 1090 3291 1091 3295
rect 1095 3291 1096 3295
rect 1090 3290 1096 3291
rect 1314 3295 1320 3296
rect 1314 3291 1315 3295
rect 1319 3291 1320 3295
rect 1934 3292 1935 3296
rect 1939 3292 1940 3296
rect 4492 3294 4494 3301
rect 4522 3299 4523 3303
rect 4527 3302 4528 3303
rect 4770 3303 4776 3304
rect 4527 3300 4649 3302
rect 4527 3299 4528 3300
rect 4522 3298 4528 3299
rect 4770 3299 4771 3303
rect 4775 3302 4776 3303
rect 5039 3303 5045 3304
rect 4775 3300 4873 3302
rect 4775 3299 4776 3300
rect 4770 3298 4776 3299
rect 5039 3299 5040 3303
rect 5044 3302 5045 3303
rect 5254 3303 5260 3304
rect 5044 3300 5089 3302
rect 5044 3299 5045 3300
rect 5039 3298 5045 3299
rect 5254 3299 5255 3303
rect 5259 3302 5260 3303
rect 5638 3303 5644 3304
rect 5638 3302 5639 3303
rect 5259 3300 5305 3302
rect 5613 3300 5639 3302
rect 5259 3299 5260 3300
rect 5254 3298 5260 3299
rect 5638 3299 5639 3300
rect 5643 3299 5644 3303
rect 5638 3298 5644 3299
rect 5238 3295 5244 3296
rect 5238 3294 5239 3295
rect 4492 3292 5239 3294
rect 1934 3291 1940 3292
rect 5238 3291 5239 3292
rect 5243 3291 5244 3295
rect 1314 3290 1320 3291
rect 5238 3290 5244 3291
rect 494 3280 500 3281
rect 110 3279 116 3280
rect 110 3275 111 3279
rect 115 3275 116 3279
rect 494 3276 495 3280
rect 499 3276 500 3280
rect 494 3275 500 3276
rect 694 3280 700 3281
rect 694 3276 695 3280
rect 699 3276 700 3280
rect 694 3275 700 3276
rect 902 3280 908 3281
rect 902 3276 903 3280
rect 907 3276 908 3280
rect 902 3275 908 3276
rect 1118 3280 1124 3281
rect 1118 3276 1119 3280
rect 1123 3276 1124 3280
rect 1118 3275 1124 3276
rect 1342 3280 1348 3281
rect 1342 3276 1343 3280
rect 1347 3276 1348 3280
rect 1342 3275 1348 3276
rect 1934 3279 1940 3280
rect 1934 3275 1935 3279
rect 1939 3275 1940 3279
rect 110 3274 116 3275
rect 1934 3274 1940 3275
rect 1950 3275 1956 3276
rect 1950 3271 1951 3275
rect 1955 3274 1956 3275
rect 2119 3275 2125 3276
rect 2119 3274 2120 3275
rect 1955 3272 2120 3274
rect 1955 3271 1956 3272
rect 1950 3270 1956 3271
rect 2119 3271 2120 3272
rect 2124 3271 2125 3275
rect 2119 3270 2125 3271
rect 2186 3275 2192 3276
rect 2186 3271 2187 3275
rect 2191 3274 2192 3275
rect 2319 3275 2325 3276
rect 2319 3274 2320 3275
rect 2191 3272 2320 3274
rect 2191 3271 2192 3272
rect 2186 3270 2192 3271
rect 2319 3271 2320 3272
rect 2324 3271 2325 3275
rect 2319 3270 2325 3271
rect 2535 3275 2541 3276
rect 2535 3271 2536 3275
rect 2540 3274 2541 3275
rect 2626 3275 2632 3276
rect 2626 3274 2627 3275
rect 2540 3272 2627 3274
rect 2540 3271 2541 3272
rect 2535 3270 2541 3271
rect 2626 3271 2627 3272
rect 2631 3271 2632 3275
rect 2626 3270 2632 3271
rect 2730 3275 2736 3276
rect 2730 3271 2731 3275
rect 2735 3274 2736 3275
rect 2743 3275 2749 3276
rect 2743 3274 2744 3275
rect 2735 3272 2744 3274
rect 2735 3271 2736 3272
rect 2730 3270 2736 3271
rect 2743 3271 2744 3272
rect 2748 3271 2749 3275
rect 2743 3270 2749 3271
rect 2935 3275 2941 3276
rect 2935 3271 2936 3275
rect 2940 3274 2941 3275
rect 3010 3275 3016 3276
rect 3010 3274 3011 3275
rect 2940 3272 3011 3274
rect 2940 3271 2941 3272
rect 2935 3270 2941 3271
rect 3010 3271 3011 3272
rect 3015 3271 3016 3275
rect 3010 3270 3016 3271
rect 3127 3275 3133 3276
rect 3127 3271 3128 3275
rect 3132 3274 3133 3275
rect 3194 3275 3200 3276
rect 3194 3274 3195 3275
rect 3132 3272 3195 3274
rect 3132 3271 3133 3272
rect 3127 3270 3133 3271
rect 3194 3271 3195 3272
rect 3199 3271 3200 3275
rect 3194 3270 3200 3271
rect 3311 3275 3317 3276
rect 3311 3271 3312 3275
rect 3316 3274 3317 3275
rect 3378 3275 3384 3276
rect 3378 3274 3379 3275
rect 3316 3272 3379 3274
rect 3316 3271 3317 3272
rect 3311 3270 3317 3271
rect 3378 3271 3379 3272
rect 3383 3271 3384 3275
rect 3378 3270 3384 3271
rect 3495 3275 3501 3276
rect 3495 3271 3496 3275
rect 3500 3274 3501 3275
rect 3562 3275 3568 3276
rect 3562 3274 3563 3275
rect 3500 3272 3563 3274
rect 3500 3271 3501 3272
rect 3495 3270 3501 3271
rect 3562 3271 3563 3272
rect 3567 3271 3568 3275
rect 3562 3270 3568 3271
rect 3678 3275 3685 3276
rect 3678 3271 3679 3275
rect 3684 3271 3685 3275
rect 3678 3270 3685 3271
rect 4783 3271 4789 3272
rect 4783 3270 4784 3271
rect 1974 3268 1980 3269
rect 3798 3268 3804 3269
rect 4677 3268 4784 3270
rect 1974 3264 1975 3268
rect 1979 3264 1980 3268
rect 1974 3263 1980 3264
rect 1994 3267 2000 3268
rect 1994 3263 1995 3267
rect 1999 3263 2000 3267
rect 1994 3262 2000 3263
rect 2194 3267 2200 3268
rect 2194 3263 2195 3267
rect 2199 3263 2200 3267
rect 2194 3262 2200 3263
rect 2410 3267 2416 3268
rect 2410 3263 2411 3267
rect 2415 3263 2416 3267
rect 2410 3262 2416 3263
rect 2618 3267 2624 3268
rect 2618 3263 2619 3267
rect 2623 3263 2624 3267
rect 2618 3262 2624 3263
rect 2810 3267 2816 3268
rect 2810 3263 2811 3267
rect 2815 3263 2816 3267
rect 2810 3262 2816 3263
rect 3002 3267 3008 3268
rect 3002 3263 3003 3267
rect 3007 3263 3008 3267
rect 3002 3262 3008 3263
rect 3186 3267 3192 3268
rect 3186 3263 3187 3267
rect 3191 3263 3192 3267
rect 3186 3262 3192 3263
rect 3370 3267 3376 3268
rect 3370 3263 3371 3267
rect 3375 3263 3376 3267
rect 3370 3262 3376 3263
rect 3554 3267 3560 3268
rect 3554 3263 3555 3267
rect 3559 3263 3560 3267
rect 3798 3264 3799 3268
rect 3803 3264 3804 3268
rect 3798 3263 3804 3264
rect 3954 3267 3960 3268
rect 3954 3263 3955 3267
rect 3959 3263 3960 3267
rect 3554 3262 3560 3263
rect 3954 3262 3960 3263
rect 4194 3267 4200 3268
rect 4194 3263 4195 3267
rect 4199 3263 4200 3267
rect 4194 3262 4200 3263
rect 4354 3267 4360 3268
rect 4354 3263 4355 3267
rect 4359 3263 4360 3267
rect 4783 3267 4784 3268
rect 4788 3267 4789 3271
rect 4978 3271 4984 3272
rect 4978 3270 4979 3271
rect 4885 3268 4979 3270
rect 4783 3266 4789 3267
rect 4978 3267 4979 3268
rect 4983 3267 4984 3271
rect 5142 3271 5148 3272
rect 5142 3270 5143 3271
rect 5085 3268 5143 3270
rect 4978 3266 4984 3267
rect 5142 3267 5143 3268
rect 5147 3267 5148 3271
rect 5346 3271 5352 3272
rect 5346 3270 5347 3271
rect 5269 3268 5347 3270
rect 5142 3266 5148 3267
rect 5346 3267 5347 3268
rect 5351 3267 5352 3271
rect 5511 3271 5517 3272
rect 5511 3270 5512 3271
rect 5453 3268 5512 3270
rect 5346 3266 5352 3267
rect 5511 3267 5512 3268
rect 5516 3267 5517 3271
rect 5511 3266 5517 3267
rect 5610 3271 5616 3272
rect 5610 3267 5611 3271
rect 5615 3267 5616 3271
rect 5610 3266 5616 3267
rect 4354 3262 4360 3263
rect 2022 3252 2028 3253
rect 1974 3251 1980 3252
rect 1974 3247 1975 3251
rect 1979 3247 1980 3251
rect 2022 3248 2023 3252
rect 2027 3248 2028 3252
rect 2022 3247 2028 3248
rect 2222 3252 2228 3253
rect 2222 3248 2223 3252
rect 2227 3248 2228 3252
rect 2222 3247 2228 3248
rect 2438 3252 2444 3253
rect 2438 3248 2439 3252
rect 2443 3248 2444 3252
rect 2438 3247 2444 3248
rect 2646 3252 2652 3253
rect 2646 3248 2647 3252
rect 2651 3248 2652 3252
rect 2646 3247 2652 3248
rect 2838 3252 2844 3253
rect 2838 3248 2839 3252
rect 2843 3248 2844 3252
rect 2838 3247 2844 3248
rect 3030 3252 3036 3253
rect 3030 3248 3031 3252
rect 3035 3248 3036 3252
rect 3030 3247 3036 3248
rect 3214 3252 3220 3253
rect 3214 3248 3215 3252
rect 3219 3248 3220 3252
rect 3214 3247 3220 3248
rect 3398 3252 3404 3253
rect 3398 3248 3399 3252
rect 3403 3248 3404 3252
rect 3398 3247 3404 3248
rect 3582 3252 3588 3253
rect 3582 3248 3583 3252
rect 3587 3248 3588 3252
rect 3582 3247 3588 3248
rect 3798 3251 3804 3252
rect 3798 3247 3799 3251
rect 3803 3247 3804 3251
rect 1974 3246 1980 3247
rect 3798 3246 3804 3247
rect 4194 3235 4200 3236
rect 4194 3231 4195 3235
rect 4199 3234 4200 3235
rect 4199 3232 4586 3234
rect 4199 3231 4200 3232
rect 4194 3230 4200 3231
rect 3983 3227 3992 3228
rect 3983 3223 3984 3227
rect 3991 3223 3992 3227
rect 3983 3222 3992 3223
rect 4223 3227 4229 3228
rect 4223 3223 4224 3227
rect 4228 3226 4229 3227
rect 4354 3227 4360 3228
rect 4354 3226 4355 3227
rect 4228 3224 4355 3226
rect 4228 3223 4229 3224
rect 4223 3222 4229 3223
rect 4354 3223 4355 3224
rect 4359 3223 4360 3227
rect 4354 3222 4360 3223
rect 4471 3227 4480 3228
rect 4471 3223 4472 3227
rect 4479 3223 4480 3227
rect 4584 3226 4586 3232
rect 4703 3227 4709 3228
rect 4703 3226 4704 3227
rect 4584 3224 4704 3226
rect 4471 3222 4480 3223
rect 4703 3223 4704 3224
rect 4708 3223 4709 3227
rect 4703 3222 4709 3223
rect 4783 3227 4789 3228
rect 4783 3223 4784 3227
rect 4788 3226 4789 3227
rect 4911 3227 4917 3228
rect 4911 3226 4912 3227
rect 4788 3224 4912 3226
rect 4788 3223 4789 3224
rect 4783 3222 4789 3223
rect 4911 3223 4912 3224
rect 4916 3223 4917 3227
rect 4911 3222 4917 3223
rect 4978 3227 4984 3228
rect 4978 3223 4979 3227
rect 4983 3226 4984 3227
rect 5111 3227 5117 3228
rect 5111 3226 5112 3227
rect 4983 3224 5112 3226
rect 4983 3223 4984 3224
rect 4978 3222 4984 3223
rect 5111 3223 5112 3224
rect 5116 3223 5117 3227
rect 5111 3222 5117 3223
rect 5295 3227 5301 3228
rect 5295 3223 5296 3227
rect 5300 3226 5301 3227
rect 5318 3227 5324 3228
rect 5318 3226 5319 3227
rect 5300 3224 5319 3226
rect 5300 3223 5301 3224
rect 5295 3222 5301 3223
rect 5318 3223 5319 3224
rect 5323 3223 5324 3227
rect 5318 3222 5324 3223
rect 5346 3227 5352 3228
rect 5346 3223 5347 3227
rect 5351 3226 5352 3227
rect 5479 3227 5485 3228
rect 5479 3226 5480 3227
rect 5351 3224 5480 3226
rect 5351 3223 5352 3224
rect 5346 3222 5352 3223
rect 5479 3223 5480 3224
rect 5484 3223 5485 3227
rect 5479 3222 5485 3223
rect 5511 3227 5517 3228
rect 5511 3223 5512 3227
rect 5516 3226 5517 3227
rect 5639 3227 5645 3228
rect 5639 3226 5640 3227
rect 5516 3224 5640 3226
rect 5516 3223 5517 3224
rect 5511 3222 5517 3223
rect 5639 3223 5640 3224
rect 5644 3223 5645 3227
rect 5639 3222 5645 3223
rect 110 3221 116 3222
rect 1934 3221 1940 3222
rect 110 3217 111 3221
rect 115 3217 116 3221
rect 110 3216 116 3217
rect 534 3220 540 3221
rect 534 3216 535 3220
rect 539 3216 540 3220
rect 534 3215 540 3216
rect 726 3220 732 3221
rect 726 3216 727 3220
rect 731 3216 732 3220
rect 726 3215 732 3216
rect 918 3220 924 3221
rect 918 3216 919 3220
rect 923 3216 924 3220
rect 918 3215 924 3216
rect 1110 3220 1116 3221
rect 1110 3216 1111 3220
rect 1115 3216 1116 3220
rect 1110 3215 1116 3216
rect 1294 3220 1300 3221
rect 1294 3216 1295 3220
rect 1299 3216 1300 3220
rect 1294 3215 1300 3216
rect 1470 3220 1476 3221
rect 1470 3216 1471 3220
rect 1475 3216 1476 3220
rect 1470 3215 1476 3216
rect 1654 3220 1660 3221
rect 1654 3216 1655 3220
rect 1659 3216 1660 3220
rect 1654 3215 1660 3216
rect 1814 3220 1820 3221
rect 1814 3216 1815 3220
rect 1819 3216 1820 3220
rect 1934 3217 1935 3221
rect 1939 3217 1940 3221
rect 1934 3216 1940 3217
rect 3838 3220 3844 3221
rect 5662 3220 5668 3221
rect 3838 3216 3839 3220
rect 3843 3216 3844 3220
rect 1814 3215 1820 3216
rect 3838 3215 3844 3216
rect 3858 3219 3864 3220
rect 3858 3215 3859 3219
rect 3863 3215 3864 3219
rect 3858 3214 3864 3215
rect 4098 3219 4104 3220
rect 4098 3215 4099 3219
rect 4103 3215 4104 3219
rect 4098 3214 4104 3215
rect 4346 3219 4352 3220
rect 4346 3215 4347 3219
rect 4351 3215 4352 3219
rect 4346 3214 4352 3215
rect 4578 3219 4584 3220
rect 4578 3215 4579 3219
rect 4583 3215 4584 3219
rect 4578 3214 4584 3215
rect 4786 3219 4792 3220
rect 4786 3215 4787 3219
rect 4791 3215 4792 3219
rect 4786 3214 4792 3215
rect 4986 3219 4992 3220
rect 4986 3215 4987 3219
rect 4991 3215 4992 3219
rect 4986 3214 4992 3215
rect 5170 3219 5176 3220
rect 5170 3215 5171 3219
rect 5175 3215 5176 3219
rect 5170 3214 5176 3215
rect 5354 3219 5360 3220
rect 5354 3215 5355 3219
rect 5359 3215 5360 3219
rect 5354 3214 5360 3215
rect 5514 3219 5520 3220
rect 5514 3215 5515 3219
rect 5519 3215 5520 3219
rect 5662 3216 5663 3220
rect 5667 3216 5668 3220
rect 5662 3215 5668 3216
rect 5514 3214 5520 3215
rect 506 3205 512 3206
rect 110 3204 116 3205
rect 110 3200 111 3204
rect 115 3200 116 3204
rect 506 3201 507 3205
rect 511 3201 512 3205
rect 506 3200 512 3201
rect 698 3205 704 3206
rect 698 3201 699 3205
rect 703 3201 704 3205
rect 698 3200 704 3201
rect 890 3205 896 3206
rect 890 3201 891 3205
rect 895 3201 896 3205
rect 890 3200 896 3201
rect 1082 3205 1088 3206
rect 1082 3201 1083 3205
rect 1087 3201 1088 3205
rect 1082 3200 1088 3201
rect 1266 3205 1272 3206
rect 1266 3201 1267 3205
rect 1271 3201 1272 3205
rect 1266 3200 1272 3201
rect 1442 3205 1448 3206
rect 1442 3201 1443 3205
rect 1447 3201 1448 3205
rect 1442 3200 1448 3201
rect 1626 3205 1632 3206
rect 1626 3201 1627 3205
rect 1631 3201 1632 3205
rect 1626 3200 1632 3201
rect 1786 3205 1792 3206
rect 1786 3201 1787 3205
rect 1791 3201 1792 3205
rect 1786 3200 1792 3201
rect 1934 3204 1940 3205
rect 3886 3204 3892 3205
rect 1934 3200 1935 3204
rect 1939 3200 1940 3204
rect 110 3199 116 3200
rect 1934 3199 1940 3200
rect 3838 3203 3844 3204
rect 3838 3199 3839 3203
rect 3843 3199 3844 3203
rect 3886 3200 3887 3204
rect 3891 3200 3892 3204
rect 3886 3199 3892 3200
rect 4126 3204 4132 3205
rect 4126 3200 4127 3204
rect 4131 3200 4132 3204
rect 4126 3199 4132 3200
rect 4374 3204 4380 3205
rect 4374 3200 4375 3204
rect 4379 3200 4380 3204
rect 4374 3199 4380 3200
rect 4606 3204 4612 3205
rect 4606 3200 4607 3204
rect 4611 3200 4612 3204
rect 4606 3199 4612 3200
rect 4814 3204 4820 3205
rect 4814 3200 4815 3204
rect 4819 3200 4820 3204
rect 4814 3199 4820 3200
rect 5014 3204 5020 3205
rect 5014 3200 5015 3204
rect 5019 3200 5020 3204
rect 5014 3199 5020 3200
rect 5198 3204 5204 3205
rect 5198 3200 5199 3204
rect 5203 3200 5204 3204
rect 5198 3199 5204 3200
rect 5382 3204 5388 3205
rect 5382 3200 5383 3204
rect 5387 3200 5388 3204
rect 5382 3199 5388 3200
rect 5542 3204 5548 3205
rect 5542 3200 5543 3204
rect 5547 3200 5548 3204
rect 5542 3199 5548 3200
rect 5662 3203 5668 3204
rect 5662 3199 5663 3203
rect 5667 3199 5668 3203
rect 3838 3198 3844 3199
rect 5662 3198 5668 3199
rect 562 3195 568 3196
rect 562 3191 563 3195
rect 567 3194 568 3195
rect 631 3195 637 3196
rect 631 3194 632 3195
rect 567 3192 632 3194
rect 567 3191 568 3192
rect 562 3190 568 3191
rect 631 3191 632 3192
rect 636 3191 637 3195
rect 631 3190 637 3191
rect 658 3195 664 3196
rect 658 3191 659 3195
rect 663 3194 664 3195
rect 823 3195 829 3196
rect 823 3194 824 3195
rect 663 3192 824 3194
rect 663 3191 664 3192
rect 658 3190 664 3191
rect 823 3191 824 3192
rect 828 3191 829 3195
rect 823 3190 829 3191
rect 855 3195 861 3196
rect 855 3191 856 3195
rect 860 3194 861 3195
rect 1015 3195 1021 3196
rect 1015 3194 1016 3195
rect 860 3192 1016 3194
rect 860 3191 861 3192
rect 855 3190 861 3191
rect 1015 3191 1016 3192
rect 1020 3191 1021 3195
rect 1015 3190 1021 3191
rect 1207 3195 1216 3196
rect 1207 3191 1208 3195
rect 1215 3191 1216 3195
rect 1207 3190 1216 3191
rect 1390 3195 1397 3196
rect 1390 3191 1391 3195
rect 1396 3191 1397 3195
rect 1390 3190 1397 3191
rect 1566 3195 1573 3196
rect 1566 3191 1567 3195
rect 1572 3191 1573 3195
rect 1566 3190 1573 3191
rect 1594 3195 1600 3196
rect 1594 3191 1595 3195
rect 1599 3194 1600 3195
rect 1751 3195 1757 3196
rect 1751 3194 1752 3195
rect 1599 3192 1752 3194
rect 1599 3191 1600 3192
rect 1594 3190 1600 3191
rect 1751 3191 1752 3192
rect 1756 3191 1757 3195
rect 1751 3190 1757 3191
rect 1783 3195 1789 3196
rect 1783 3191 1784 3195
rect 1788 3194 1789 3195
rect 1911 3195 1917 3196
rect 1911 3194 1912 3195
rect 1788 3192 1912 3194
rect 1788 3191 1789 3192
rect 1783 3190 1789 3191
rect 1911 3191 1912 3192
rect 1916 3191 1917 3195
rect 1911 3190 1917 3191
rect 1974 3193 1980 3194
rect 3798 3193 3804 3194
rect 1974 3189 1975 3193
rect 1979 3189 1980 3193
rect 1974 3188 1980 3189
rect 2462 3192 2468 3193
rect 2462 3188 2463 3192
rect 2467 3188 2468 3192
rect 2462 3187 2468 3188
rect 2662 3192 2668 3193
rect 2662 3188 2663 3192
rect 2667 3188 2668 3192
rect 2662 3187 2668 3188
rect 2862 3192 2868 3193
rect 2862 3188 2863 3192
rect 2867 3188 2868 3192
rect 2862 3187 2868 3188
rect 3054 3192 3060 3193
rect 3054 3188 3055 3192
rect 3059 3188 3060 3192
rect 3054 3187 3060 3188
rect 3238 3192 3244 3193
rect 3238 3188 3239 3192
rect 3243 3188 3244 3192
rect 3238 3187 3244 3188
rect 3430 3192 3436 3193
rect 3430 3188 3431 3192
rect 3435 3188 3436 3192
rect 3430 3187 3436 3188
rect 3622 3192 3628 3193
rect 3622 3188 3623 3192
rect 3627 3188 3628 3192
rect 3798 3189 3799 3193
rect 3803 3189 3804 3193
rect 3798 3188 3804 3189
rect 3622 3187 3628 3188
rect 2434 3177 2440 3178
rect 1974 3176 1980 3177
rect 1974 3172 1975 3176
rect 1979 3172 1980 3176
rect 2434 3173 2435 3177
rect 2439 3173 2440 3177
rect 2434 3172 2440 3173
rect 2634 3177 2640 3178
rect 2634 3173 2635 3177
rect 2639 3173 2640 3177
rect 2634 3172 2640 3173
rect 2834 3177 2840 3178
rect 2834 3173 2835 3177
rect 2839 3173 2840 3177
rect 2834 3172 2840 3173
rect 3026 3177 3032 3178
rect 3026 3173 3027 3177
rect 3031 3173 3032 3177
rect 3026 3172 3032 3173
rect 3210 3177 3216 3178
rect 3210 3173 3211 3177
rect 3215 3173 3216 3177
rect 3210 3172 3216 3173
rect 3402 3177 3408 3178
rect 3402 3173 3403 3177
rect 3407 3173 3408 3177
rect 3402 3172 3408 3173
rect 3594 3177 3600 3178
rect 3594 3173 3595 3177
rect 3599 3173 3600 3177
rect 3594 3172 3600 3173
rect 3798 3176 3804 3177
rect 3798 3172 3799 3176
rect 3803 3172 3804 3176
rect 1974 3171 1980 3172
rect 3798 3171 3804 3172
rect 2426 3167 2432 3168
rect 2426 3163 2427 3167
rect 2431 3166 2432 3167
rect 2559 3167 2565 3168
rect 2559 3166 2560 3167
rect 2431 3164 2560 3166
rect 2431 3163 2432 3164
rect 2426 3162 2432 3163
rect 2559 3163 2560 3164
rect 2564 3163 2565 3167
rect 2559 3162 2565 3163
rect 2631 3167 2637 3168
rect 2631 3163 2632 3167
rect 2636 3166 2637 3167
rect 2759 3167 2765 3168
rect 2759 3166 2760 3167
rect 2636 3164 2760 3166
rect 2636 3163 2637 3164
rect 2631 3162 2637 3163
rect 2759 3163 2760 3164
rect 2764 3163 2765 3167
rect 2759 3162 2765 3163
rect 2906 3167 2912 3168
rect 2906 3163 2907 3167
rect 2911 3166 2912 3167
rect 2959 3167 2965 3168
rect 2959 3166 2960 3167
rect 2911 3164 2960 3166
rect 2911 3163 2912 3164
rect 2906 3162 2912 3163
rect 2959 3163 2960 3164
rect 2964 3163 2965 3167
rect 2959 3162 2965 3163
rect 2991 3167 2997 3168
rect 2991 3163 2992 3167
rect 2996 3166 2997 3167
rect 3151 3167 3157 3168
rect 3151 3166 3152 3167
rect 2996 3164 3152 3166
rect 2996 3163 2997 3164
rect 2991 3162 2997 3163
rect 3151 3163 3152 3164
rect 3156 3163 3157 3167
rect 3151 3162 3157 3163
rect 3335 3167 3344 3168
rect 3335 3163 3336 3167
rect 3343 3163 3344 3167
rect 3335 3162 3344 3163
rect 3526 3167 3533 3168
rect 3526 3163 3527 3167
rect 3532 3163 3533 3167
rect 3719 3167 3725 3168
rect 3719 3166 3720 3167
rect 3526 3162 3533 3163
rect 3619 3164 3720 3166
rect 3306 3159 3312 3160
rect 550 3155 556 3156
rect 550 3151 551 3155
rect 555 3151 556 3155
rect 855 3155 861 3156
rect 855 3154 856 3155
rect 797 3152 856 3154
rect 550 3150 556 3151
rect 855 3151 856 3152
rect 860 3151 861 3155
rect 1210 3155 1216 3156
rect 855 3150 861 3151
rect 988 3146 990 3153
rect 1154 3147 1160 3148
rect 1154 3146 1155 3147
rect 988 3144 1155 3146
rect 1154 3143 1155 3144
rect 1159 3143 1160 3147
rect 1180 3146 1182 3153
rect 1210 3151 1211 3155
rect 1215 3154 1216 3155
rect 1594 3155 1600 3156
rect 1594 3154 1595 3155
rect 1215 3152 1273 3154
rect 1541 3152 1595 3154
rect 1215 3151 1216 3152
rect 1210 3150 1216 3151
rect 1594 3151 1595 3152
rect 1599 3151 1600 3155
rect 1783 3155 1789 3156
rect 1783 3154 1784 3155
rect 1725 3152 1784 3154
rect 1594 3150 1600 3151
rect 1783 3151 1784 3152
rect 1788 3151 1789 3155
rect 1950 3155 1956 3156
rect 1950 3154 1951 3155
rect 1885 3152 1951 3154
rect 1783 3150 1789 3151
rect 1950 3151 1951 3152
rect 1955 3151 1956 3155
rect 3306 3155 3307 3159
rect 3311 3158 3312 3159
rect 3619 3158 3621 3164
rect 3719 3163 3720 3164
rect 3724 3163 3725 3167
rect 3719 3162 3725 3163
rect 3311 3156 3621 3158
rect 3311 3155 3312 3156
rect 3306 3154 3312 3155
rect 1950 3150 1956 3151
rect 1398 3147 1404 3148
rect 1398 3146 1399 3147
rect 1180 3144 1399 3146
rect 1154 3142 1160 3143
rect 1398 3143 1399 3144
rect 1403 3143 1404 3147
rect 1398 3142 1404 3143
rect 3838 3129 3844 3130
rect 5662 3129 5668 3130
rect 2631 3127 2637 3128
rect 2631 3126 2632 3127
rect 2533 3124 2632 3126
rect 2631 3123 2632 3124
rect 2636 3123 2637 3127
rect 2631 3122 2637 3123
rect 2730 3127 2736 3128
rect 2730 3123 2731 3127
rect 2735 3123 2736 3127
rect 2991 3127 2997 3128
rect 2991 3126 2992 3127
rect 2933 3124 2992 3126
rect 2730 3122 2736 3123
rect 2991 3123 2992 3124
rect 2996 3123 2997 3127
rect 2991 3122 2997 3123
rect 3122 3127 3128 3128
rect 3122 3123 3123 3127
rect 3127 3123 3128 3127
rect 3122 3122 3128 3123
rect 3306 3127 3312 3128
rect 3306 3123 3307 3127
rect 3311 3123 3312 3127
rect 3306 3122 3312 3123
rect 3338 3127 3344 3128
rect 3338 3123 3339 3127
rect 3343 3126 3344 3127
rect 3678 3127 3684 3128
rect 3343 3124 3409 3126
rect 3343 3123 3344 3124
rect 3338 3122 3344 3123
rect 3678 3123 3679 3127
rect 3683 3123 3684 3127
rect 3838 3125 3839 3129
rect 3843 3125 3844 3129
rect 3838 3124 3844 3125
rect 3902 3128 3908 3129
rect 3902 3124 3903 3128
rect 3907 3124 3908 3128
rect 3902 3123 3908 3124
rect 4134 3128 4140 3129
rect 4134 3124 4135 3128
rect 4139 3124 4140 3128
rect 4134 3123 4140 3124
rect 4358 3128 4364 3129
rect 4358 3124 4359 3128
rect 4363 3124 4364 3128
rect 4358 3123 4364 3124
rect 4582 3128 4588 3129
rect 4582 3124 4583 3128
rect 4587 3124 4588 3128
rect 4582 3123 4588 3124
rect 4806 3128 4812 3129
rect 4806 3124 4807 3128
rect 4811 3124 4812 3128
rect 4806 3123 4812 3124
rect 5030 3128 5036 3129
rect 5030 3124 5031 3128
rect 5035 3124 5036 3128
rect 5662 3125 5663 3129
rect 5667 3125 5668 3129
rect 5662 3124 5668 3125
rect 5030 3123 5036 3124
rect 3678 3122 3684 3123
rect 658 3115 664 3116
rect 434 3111 440 3112
rect 434 3107 435 3111
rect 439 3107 440 3111
rect 658 3111 659 3115
rect 663 3111 664 3115
rect 1566 3115 1572 3116
rect 658 3110 664 3111
rect 706 3111 712 3112
rect 434 3106 440 3107
rect 706 3107 707 3111
rect 711 3107 712 3111
rect 706 3106 712 3107
rect 842 3111 848 3112
rect 842 3107 843 3111
rect 847 3107 848 3111
rect 842 3106 848 3107
rect 978 3111 984 3112
rect 978 3107 979 3111
rect 983 3107 984 3111
rect 978 3106 984 3107
rect 1114 3111 1120 3112
rect 1114 3107 1115 3111
rect 1119 3107 1120 3111
rect 1114 3106 1120 3107
rect 1250 3111 1256 3112
rect 1250 3107 1251 3111
rect 1255 3107 1256 3111
rect 1250 3106 1256 3107
rect 1386 3111 1392 3112
rect 1386 3107 1387 3111
rect 1391 3107 1392 3111
rect 1566 3111 1567 3115
rect 1571 3111 1572 3115
rect 3874 3113 3880 3114
rect 3838 3112 3844 3113
rect 1566 3110 1572 3111
rect 1658 3111 1664 3112
rect 1386 3106 1392 3107
rect 1658 3107 1659 3111
rect 1663 3107 1664 3111
rect 1658 3106 1664 3107
rect 1794 3111 1800 3112
rect 1794 3107 1795 3111
rect 1799 3107 1800 3111
rect 3838 3108 3839 3112
rect 3843 3108 3844 3112
rect 3874 3109 3875 3113
rect 3879 3109 3880 3113
rect 3874 3108 3880 3109
rect 4106 3113 4112 3114
rect 4106 3109 4107 3113
rect 4111 3109 4112 3113
rect 4106 3108 4112 3109
rect 4330 3113 4336 3114
rect 4330 3109 4331 3113
rect 4335 3109 4336 3113
rect 4330 3108 4336 3109
rect 4554 3113 4560 3114
rect 4554 3109 4555 3113
rect 4559 3109 4560 3113
rect 4554 3108 4560 3109
rect 4778 3113 4784 3114
rect 4778 3109 4779 3113
rect 4783 3109 4784 3113
rect 4778 3108 4784 3109
rect 5002 3113 5008 3114
rect 5002 3109 5003 3113
rect 5007 3109 5008 3113
rect 5002 3108 5008 3109
rect 5662 3112 5668 3113
rect 5662 3108 5663 3112
rect 5667 3108 5668 3112
rect 3838 3107 3844 3108
rect 5662 3107 5668 3108
rect 1794 3106 1800 3107
rect 3954 3103 3960 3104
rect 3954 3099 3955 3103
rect 3959 3102 3960 3103
rect 3999 3103 4005 3104
rect 3999 3102 4000 3103
rect 3959 3100 4000 3102
rect 3959 3099 3960 3100
rect 3954 3098 3960 3099
rect 3999 3099 4000 3100
rect 4004 3099 4005 3103
rect 3999 3098 4005 3099
rect 4231 3103 4240 3104
rect 4231 3099 4232 3103
rect 4239 3099 4240 3103
rect 4231 3098 4240 3099
rect 4454 3103 4461 3104
rect 4454 3099 4455 3103
rect 4460 3099 4461 3103
rect 4454 3098 4461 3099
rect 4679 3103 4688 3104
rect 4679 3099 4680 3103
rect 4687 3099 4688 3103
rect 4679 3098 4688 3099
rect 4903 3103 4912 3104
rect 4903 3099 4904 3103
rect 4911 3099 4912 3103
rect 5127 3103 5133 3104
rect 5127 3102 5128 3103
rect 4903 3098 4912 3099
rect 4916 3100 5128 3102
rect 4202 3095 4208 3096
rect 4202 3091 4203 3095
rect 4207 3094 4208 3095
rect 4916 3094 4918 3100
rect 5127 3099 5128 3100
rect 5132 3099 5133 3103
rect 5127 3098 5133 3099
rect 4207 3092 4918 3094
rect 4207 3091 4208 3092
rect 4202 3090 4208 3091
rect 2426 3083 2432 3084
rect 2426 3079 2427 3083
rect 2431 3079 2432 3083
rect 2838 3083 2844 3084
rect 2426 3078 2432 3079
rect 2562 3079 2568 3080
rect 2562 3075 2563 3079
rect 2567 3075 2568 3079
rect 2838 3079 2839 3083
rect 2843 3079 2844 3083
rect 3463 3083 3469 3084
rect 3463 3082 3464 3083
rect 3333 3080 3464 3082
rect 2838 3078 2844 3079
rect 3010 3079 3016 3080
rect 2562 3074 2568 3075
rect 3010 3075 3011 3079
rect 3015 3075 3016 3079
rect 3463 3079 3464 3080
rect 3468 3079 3469 3083
rect 3463 3078 3469 3079
rect 3526 3083 3532 3084
rect 3526 3079 3527 3083
rect 3531 3079 3532 3083
rect 3526 3078 3532 3079
rect 3010 3074 3016 3075
rect 550 3071 557 3072
rect 550 3067 551 3071
rect 556 3067 557 3071
rect 550 3066 557 3067
rect 687 3071 693 3072
rect 687 3067 688 3071
rect 692 3070 693 3071
rect 706 3071 712 3072
rect 706 3070 707 3071
rect 692 3068 707 3070
rect 692 3067 693 3068
rect 687 3066 693 3067
rect 706 3067 707 3068
rect 711 3067 712 3071
rect 706 3066 712 3067
rect 823 3071 829 3072
rect 823 3067 824 3071
rect 828 3070 829 3071
rect 842 3071 848 3072
rect 842 3070 843 3071
rect 828 3068 843 3070
rect 828 3067 829 3068
rect 823 3066 829 3067
rect 842 3067 843 3068
rect 847 3067 848 3071
rect 842 3066 848 3067
rect 959 3071 965 3072
rect 959 3067 960 3071
rect 964 3070 965 3071
rect 978 3071 984 3072
rect 978 3070 979 3071
rect 964 3068 979 3070
rect 964 3067 965 3068
rect 959 3066 965 3067
rect 978 3067 979 3068
rect 983 3067 984 3071
rect 978 3066 984 3067
rect 1095 3071 1101 3072
rect 1095 3067 1096 3071
rect 1100 3070 1101 3071
rect 1114 3071 1120 3072
rect 1114 3070 1115 3071
rect 1100 3068 1115 3070
rect 1100 3067 1101 3068
rect 1095 3066 1101 3067
rect 1114 3067 1115 3068
rect 1119 3067 1120 3071
rect 1114 3066 1120 3067
rect 1231 3071 1237 3072
rect 1231 3067 1232 3071
rect 1236 3070 1237 3071
rect 1250 3071 1256 3072
rect 1250 3070 1251 3071
rect 1236 3068 1251 3070
rect 1236 3067 1237 3068
rect 1231 3066 1237 3067
rect 1250 3067 1251 3068
rect 1255 3067 1256 3071
rect 1250 3066 1256 3067
rect 1367 3071 1373 3072
rect 1367 3067 1368 3071
rect 1372 3070 1373 3071
rect 1386 3071 1392 3072
rect 1386 3070 1387 3071
rect 1372 3068 1387 3070
rect 1372 3067 1373 3068
rect 1367 3066 1373 3067
rect 1386 3067 1387 3068
rect 1391 3067 1392 3071
rect 1386 3066 1392 3067
rect 1398 3071 1404 3072
rect 1398 3067 1399 3071
rect 1403 3070 1404 3071
rect 1503 3071 1509 3072
rect 1503 3070 1504 3071
rect 1403 3068 1504 3070
rect 1403 3067 1404 3068
rect 1398 3066 1404 3067
rect 1503 3067 1504 3068
rect 1508 3067 1509 3071
rect 1503 3066 1509 3067
rect 1639 3071 1645 3072
rect 1639 3067 1640 3071
rect 1644 3070 1645 3071
rect 1658 3071 1664 3072
rect 1658 3070 1659 3071
rect 1644 3068 1659 3070
rect 1644 3067 1645 3068
rect 1639 3066 1645 3067
rect 1658 3067 1659 3068
rect 1663 3067 1664 3071
rect 1658 3066 1664 3067
rect 1775 3071 1781 3072
rect 1775 3067 1776 3071
rect 1780 3070 1781 3071
rect 1794 3071 1800 3072
rect 1794 3070 1795 3071
rect 1780 3068 1795 3070
rect 1780 3067 1781 3068
rect 1775 3066 1781 3067
rect 1794 3067 1795 3068
rect 1799 3067 1800 3071
rect 1794 3066 1800 3067
rect 1906 3071 1917 3072
rect 1906 3067 1907 3071
rect 1911 3067 1912 3071
rect 1916 3067 1917 3071
rect 1906 3066 1917 3067
rect 110 3064 116 3065
rect 1934 3064 1940 3065
rect 110 3060 111 3064
rect 115 3060 116 3064
rect 110 3059 116 3060
rect 426 3063 432 3064
rect 426 3059 427 3063
rect 431 3059 432 3063
rect 426 3058 432 3059
rect 562 3063 568 3064
rect 562 3059 563 3063
rect 567 3059 568 3063
rect 562 3058 568 3059
rect 698 3063 704 3064
rect 698 3059 699 3063
rect 703 3059 704 3063
rect 698 3058 704 3059
rect 834 3063 840 3064
rect 834 3059 835 3063
rect 839 3059 840 3063
rect 834 3058 840 3059
rect 970 3063 976 3064
rect 970 3059 971 3063
rect 975 3059 976 3063
rect 970 3058 976 3059
rect 1106 3063 1112 3064
rect 1106 3059 1107 3063
rect 1111 3059 1112 3063
rect 1106 3058 1112 3059
rect 1242 3063 1248 3064
rect 1242 3059 1243 3063
rect 1247 3059 1248 3063
rect 1242 3058 1248 3059
rect 1378 3063 1384 3064
rect 1378 3059 1379 3063
rect 1383 3059 1384 3063
rect 1378 3058 1384 3059
rect 1514 3063 1520 3064
rect 1514 3059 1515 3063
rect 1519 3059 1520 3063
rect 1514 3058 1520 3059
rect 1650 3063 1656 3064
rect 1650 3059 1651 3063
rect 1655 3059 1656 3063
rect 1650 3058 1656 3059
rect 1786 3063 1792 3064
rect 1786 3059 1787 3063
rect 1791 3059 1792 3063
rect 1934 3060 1935 3064
rect 1939 3060 1940 3064
rect 1934 3059 1940 3060
rect 3970 3063 3976 3064
rect 3970 3059 3971 3063
rect 3975 3059 3976 3063
rect 1786 3058 1792 3059
rect 3970 3058 3976 3059
rect 4202 3063 4208 3064
rect 4202 3059 4203 3063
rect 4207 3059 4208 3063
rect 4202 3058 4208 3059
rect 4234 3063 4240 3064
rect 4234 3059 4235 3063
rect 4239 3062 4240 3063
rect 4474 3063 4480 3064
rect 4239 3060 4337 3062
rect 4239 3059 4240 3060
rect 4234 3058 4240 3059
rect 4474 3059 4475 3063
rect 4479 3062 4480 3063
rect 4682 3063 4688 3064
rect 4479 3060 4561 3062
rect 4479 3059 4480 3060
rect 4474 3058 4480 3059
rect 4682 3059 4683 3063
rect 4687 3062 4688 3063
rect 4906 3063 4912 3064
rect 4687 3060 4785 3062
rect 4687 3059 4688 3060
rect 4682 3058 4688 3059
rect 4906 3059 4907 3063
rect 4911 3062 4912 3063
rect 4911 3060 5009 3062
rect 4911 3059 4912 3060
rect 4906 3058 4912 3059
rect 454 3048 460 3049
rect 110 3047 116 3048
rect 110 3043 111 3047
rect 115 3043 116 3047
rect 454 3044 455 3048
rect 459 3044 460 3048
rect 454 3043 460 3044
rect 590 3048 596 3049
rect 590 3044 591 3048
rect 595 3044 596 3048
rect 590 3043 596 3044
rect 726 3048 732 3049
rect 726 3044 727 3048
rect 731 3044 732 3048
rect 726 3043 732 3044
rect 862 3048 868 3049
rect 862 3044 863 3048
rect 867 3044 868 3048
rect 862 3043 868 3044
rect 998 3048 1004 3049
rect 998 3044 999 3048
rect 1003 3044 1004 3048
rect 998 3043 1004 3044
rect 1134 3048 1140 3049
rect 1134 3044 1135 3048
rect 1139 3044 1140 3048
rect 1134 3043 1140 3044
rect 1270 3048 1276 3049
rect 1270 3044 1271 3048
rect 1275 3044 1276 3048
rect 1270 3043 1276 3044
rect 1406 3048 1412 3049
rect 1406 3044 1407 3048
rect 1411 3044 1412 3048
rect 1406 3043 1412 3044
rect 1542 3048 1548 3049
rect 1542 3044 1543 3048
rect 1547 3044 1548 3048
rect 1542 3043 1548 3044
rect 1678 3048 1684 3049
rect 1678 3044 1679 3048
rect 1683 3044 1684 3048
rect 1678 3043 1684 3044
rect 1814 3048 1820 3049
rect 1814 3044 1815 3048
rect 1819 3044 1820 3048
rect 1814 3043 1820 3044
rect 1934 3047 1940 3048
rect 1934 3043 1935 3047
rect 1939 3043 1940 3047
rect 110 3042 116 3043
rect 1934 3042 1940 3043
rect 2455 3039 2461 3040
rect 2455 3035 2456 3039
rect 2460 3038 2461 3039
rect 2562 3039 2568 3040
rect 2562 3038 2563 3039
rect 2460 3036 2563 3038
rect 2460 3035 2461 3036
rect 2455 3034 2461 3035
rect 2562 3035 2563 3036
rect 2567 3035 2568 3039
rect 2562 3034 2568 3035
rect 2610 3039 2616 3040
rect 2610 3035 2611 3039
rect 2615 3038 2616 3039
rect 2679 3039 2685 3040
rect 2679 3038 2680 3039
rect 2615 3036 2680 3038
rect 2615 3035 2616 3036
rect 2610 3034 2616 3035
rect 2679 3035 2680 3036
rect 2684 3035 2685 3039
rect 2679 3034 2685 3035
rect 2903 3039 2909 3040
rect 2903 3035 2904 3039
rect 2908 3038 2909 3039
rect 3010 3039 3016 3040
rect 3010 3038 3011 3039
rect 2908 3036 3011 3038
rect 2908 3035 2909 3036
rect 2903 3034 2909 3035
rect 3010 3035 3011 3036
rect 3015 3035 3016 3039
rect 3010 3034 3016 3035
rect 3122 3039 3133 3040
rect 3122 3035 3123 3039
rect 3127 3035 3128 3039
rect 3132 3035 3133 3039
rect 3122 3034 3133 3035
rect 3358 3039 3365 3040
rect 3358 3035 3359 3039
rect 3364 3035 3365 3039
rect 3358 3034 3365 3035
rect 3463 3039 3469 3040
rect 3463 3035 3464 3039
rect 3468 3038 3469 3039
rect 3591 3039 3597 3040
rect 3591 3038 3592 3039
rect 3468 3036 3592 3038
rect 3468 3035 3469 3036
rect 3463 3034 3469 3035
rect 3591 3035 3592 3036
rect 3596 3035 3597 3039
rect 4878 3039 4884 3040
rect 4878 3038 4879 3039
rect 3591 3034 3597 3035
rect 4244 3036 4879 3038
rect 1974 3032 1980 3033
rect 3798 3032 3804 3033
rect 1974 3028 1975 3032
rect 1979 3028 1980 3032
rect 1974 3027 1980 3028
rect 2330 3031 2336 3032
rect 2330 3027 2331 3031
rect 2335 3027 2336 3031
rect 2330 3026 2336 3027
rect 2554 3031 2560 3032
rect 2554 3027 2555 3031
rect 2559 3027 2560 3031
rect 2554 3026 2560 3027
rect 2778 3031 2784 3032
rect 2778 3027 2779 3031
rect 2783 3027 2784 3031
rect 2778 3026 2784 3027
rect 3002 3031 3008 3032
rect 3002 3027 3003 3031
rect 3007 3027 3008 3031
rect 3002 3026 3008 3027
rect 3234 3031 3240 3032
rect 3234 3027 3235 3031
rect 3239 3027 3240 3031
rect 3234 3026 3240 3027
rect 3466 3031 3472 3032
rect 3466 3027 3467 3031
rect 3471 3027 3472 3031
rect 3798 3028 3799 3032
rect 3803 3028 3804 3032
rect 3798 3027 3804 3028
rect 3990 3031 3996 3032
rect 3990 3027 3991 3031
rect 3995 3027 3996 3031
rect 4244 3030 4246 3036
rect 4878 3035 4879 3036
rect 4883 3035 4884 3039
rect 4878 3034 4884 3035
rect 4173 3028 4246 3030
rect 4454 3031 4460 3032
rect 3466 3026 3472 3027
rect 3990 3026 3996 3027
rect 4250 3027 4256 3028
rect 4250 3023 4251 3027
rect 4255 3023 4256 3027
rect 4454 3027 4455 3031
rect 4459 3027 4460 3031
rect 4454 3026 4460 3027
rect 4586 3027 4592 3028
rect 4250 3022 4256 3023
rect 4586 3023 4587 3027
rect 4591 3023 4592 3027
rect 4586 3022 4592 3023
rect 4762 3027 4768 3028
rect 4762 3023 4763 3027
rect 4767 3023 4768 3027
rect 4762 3022 4768 3023
rect 2358 3016 2364 3017
rect 1974 3015 1980 3016
rect 1974 3011 1975 3015
rect 1979 3011 1980 3015
rect 2358 3012 2359 3016
rect 2363 3012 2364 3016
rect 2358 3011 2364 3012
rect 2582 3016 2588 3017
rect 2582 3012 2583 3016
rect 2587 3012 2588 3016
rect 2582 3011 2588 3012
rect 2806 3016 2812 3017
rect 2806 3012 2807 3016
rect 2811 3012 2812 3016
rect 2806 3011 2812 3012
rect 3030 3016 3036 3017
rect 3030 3012 3031 3016
rect 3035 3012 3036 3016
rect 3030 3011 3036 3012
rect 3262 3016 3268 3017
rect 3262 3012 3263 3016
rect 3267 3012 3268 3016
rect 3262 3011 3268 3012
rect 3494 3016 3500 3017
rect 3494 3012 3495 3016
rect 3499 3012 3500 3016
rect 3494 3011 3500 3012
rect 3798 3015 3804 3016
rect 3798 3011 3799 3015
rect 3803 3011 3804 3015
rect 1974 3010 1980 3011
rect 3798 3010 3804 3011
rect 3970 2987 3976 2988
rect 3970 2983 3971 2987
rect 3975 2986 3976 2987
rect 4031 2987 4037 2988
rect 4031 2986 4032 2987
rect 3975 2984 4032 2986
rect 3975 2983 3976 2984
rect 3970 2982 3976 2983
rect 4031 2983 4032 2984
rect 4036 2983 4037 2987
rect 4031 2982 4037 2983
rect 4199 2987 4205 2988
rect 4199 2983 4200 2987
rect 4204 2986 4205 2987
rect 4250 2987 4256 2988
rect 4250 2986 4251 2987
rect 4204 2984 4251 2986
rect 4204 2983 4205 2984
rect 4199 2982 4205 2983
rect 4250 2983 4251 2984
rect 4255 2983 4256 2987
rect 4250 2982 4256 2983
rect 4366 2987 4373 2988
rect 4366 2983 4367 2987
rect 4372 2983 4373 2987
rect 4366 2982 4373 2983
rect 4535 2987 4541 2988
rect 4535 2983 4536 2987
rect 4540 2986 4541 2987
rect 4586 2987 4592 2988
rect 4586 2986 4587 2987
rect 4540 2984 4587 2986
rect 4540 2983 4541 2984
rect 4535 2982 4541 2983
rect 4586 2983 4587 2984
rect 4591 2983 4592 2987
rect 4586 2982 4592 2983
rect 4703 2987 4709 2988
rect 4703 2983 4704 2987
rect 4708 2986 4709 2987
rect 4762 2987 4768 2988
rect 4762 2986 4763 2987
rect 4708 2984 4763 2986
rect 4708 2983 4709 2984
rect 4703 2982 4709 2983
rect 4762 2983 4763 2984
rect 4767 2983 4768 2987
rect 4762 2982 4768 2983
rect 4878 2987 4885 2988
rect 4878 2983 4879 2987
rect 4884 2983 4885 2987
rect 4878 2982 4885 2983
rect 3838 2980 3844 2981
rect 5662 2980 5668 2981
rect 3838 2976 3839 2980
rect 3843 2976 3844 2980
rect 3838 2975 3844 2976
rect 3906 2979 3912 2980
rect 3906 2975 3907 2979
rect 3911 2975 3912 2979
rect 3906 2974 3912 2975
rect 4074 2979 4080 2980
rect 4074 2975 4075 2979
rect 4079 2975 4080 2979
rect 4074 2974 4080 2975
rect 4242 2979 4248 2980
rect 4242 2975 4243 2979
rect 4247 2975 4248 2979
rect 4242 2974 4248 2975
rect 4410 2979 4416 2980
rect 4410 2975 4411 2979
rect 4415 2975 4416 2979
rect 4410 2974 4416 2975
rect 4578 2979 4584 2980
rect 4578 2975 4579 2979
rect 4583 2975 4584 2979
rect 4578 2974 4584 2975
rect 4754 2979 4760 2980
rect 4754 2975 4755 2979
rect 4759 2975 4760 2979
rect 5662 2976 5663 2980
rect 5667 2976 5668 2980
rect 5662 2975 5668 2976
rect 4754 2974 4760 2975
rect 3934 2964 3940 2965
rect 3838 2963 3844 2964
rect 110 2961 116 2962
rect 1934 2961 1940 2962
rect 110 2957 111 2961
rect 115 2957 116 2961
rect 110 2956 116 2957
rect 198 2960 204 2961
rect 198 2956 199 2960
rect 203 2956 204 2960
rect 198 2955 204 2956
rect 510 2960 516 2961
rect 510 2956 511 2960
rect 515 2956 516 2960
rect 510 2955 516 2956
rect 814 2960 820 2961
rect 814 2956 815 2960
rect 819 2956 820 2960
rect 814 2955 820 2956
rect 1110 2960 1116 2961
rect 1110 2956 1111 2960
rect 1115 2956 1116 2960
rect 1110 2955 1116 2956
rect 1414 2960 1420 2961
rect 1414 2956 1415 2960
rect 1419 2956 1420 2960
rect 1414 2955 1420 2956
rect 1718 2960 1724 2961
rect 1718 2956 1719 2960
rect 1723 2956 1724 2960
rect 1934 2957 1935 2961
rect 1939 2957 1940 2961
rect 3838 2959 3839 2963
rect 3843 2959 3844 2963
rect 3934 2960 3935 2964
rect 3939 2960 3940 2964
rect 3934 2959 3940 2960
rect 4102 2964 4108 2965
rect 4102 2960 4103 2964
rect 4107 2960 4108 2964
rect 4102 2959 4108 2960
rect 4270 2964 4276 2965
rect 4270 2960 4271 2964
rect 4275 2960 4276 2964
rect 4270 2959 4276 2960
rect 4438 2964 4444 2965
rect 4438 2960 4439 2964
rect 4443 2960 4444 2964
rect 4438 2959 4444 2960
rect 4606 2964 4612 2965
rect 4606 2960 4607 2964
rect 4611 2960 4612 2964
rect 4606 2959 4612 2960
rect 4782 2964 4788 2965
rect 4782 2960 4783 2964
rect 4787 2960 4788 2964
rect 4782 2959 4788 2960
rect 5662 2963 5668 2964
rect 5662 2959 5663 2963
rect 5667 2959 5668 2963
rect 3838 2958 3844 2959
rect 5662 2958 5668 2959
rect 1934 2956 1940 2957
rect 1718 2955 1724 2956
rect 170 2945 176 2946
rect 110 2944 116 2945
rect 110 2940 111 2944
rect 115 2940 116 2944
rect 170 2941 171 2945
rect 175 2941 176 2945
rect 170 2940 176 2941
rect 482 2945 488 2946
rect 482 2941 483 2945
rect 487 2941 488 2945
rect 482 2940 488 2941
rect 786 2945 792 2946
rect 786 2941 787 2945
rect 791 2941 792 2945
rect 786 2940 792 2941
rect 1082 2945 1088 2946
rect 1082 2941 1083 2945
rect 1087 2941 1088 2945
rect 1082 2940 1088 2941
rect 1386 2945 1392 2946
rect 1386 2941 1387 2945
rect 1391 2941 1392 2945
rect 1386 2940 1392 2941
rect 1690 2945 1696 2946
rect 1974 2945 1980 2946
rect 3798 2945 3804 2946
rect 1690 2941 1691 2945
rect 1695 2941 1696 2945
rect 1690 2940 1696 2941
rect 1934 2944 1940 2945
rect 1934 2940 1935 2944
rect 1939 2940 1940 2944
rect 1974 2941 1975 2945
rect 1979 2941 1980 2945
rect 1974 2940 1980 2941
rect 2142 2944 2148 2945
rect 2142 2940 2143 2944
rect 2147 2940 2148 2944
rect 110 2939 116 2940
rect 1934 2939 1940 2940
rect 2142 2939 2148 2940
rect 2342 2944 2348 2945
rect 2342 2940 2343 2944
rect 2347 2940 2348 2944
rect 2342 2939 2348 2940
rect 2542 2944 2548 2945
rect 2542 2940 2543 2944
rect 2547 2940 2548 2944
rect 2542 2939 2548 2940
rect 2742 2944 2748 2945
rect 2742 2940 2743 2944
rect 2747 2940 2748 2944
rect 2742 2939 2748 2940
rect 2934 2944 2940 2945
rect 2934 2940 2935 2944
rect 2939 2940 2940 2944
rect 2934 2939 2940 2940
rect 3134 2944 3140 2945
rect 3134 2940 3135 2944
rect 3139 2940 3140 2944
rect 3134 2939 3140 2940
rect 3334 2944 3340 2945
rect 3334 2940 3335 2944
rect 3339 2940 3340 2944
rect 3798 2941 3799 2945
rect 3803 2941 3804 2945
rect 3798 2940 3804 2941
rect 3334 2939 3340 2940
rect 295 2935 301 2936
rect 295 2931 296 2935
rect 300 2934 301 2935
rect 434 2935 440 2936
rect 434 2934 435 2935
rect 300 2932 435 2934
rect 300 2931 301 2932
rect 295 2930 301 2931
rect 434 2931 435 2932
rect 439 2931 440 2935
rect 434 2930 440 2931
rect 442 2935 448 2936
rect 442 2931 443 2935
rect 447 2934 448 2935
rect 607 2935 613 2936
rect 607 2934 608 2935
rect 447 2932 608 2934
rect 447 2931 448 2932
rect 442 2930 448 2931
rect 607 2931 608 2932
rect 612 2931 613 2935
rect 607 2930 613 2931
rect 722 2935 728 2936
rect 722 2931 723 2935
rect 727 2934 728 2935
rect 911 2935 917 2936
rect 911 2934 912 2935
rect 727 2932 912 2934
rect 727 2931 728 2932
rect 722 2930 728 2931
rect 911 2931 912 2932
rect 916 2931 917 2935
rect 911 2930 917 2931
rect 1207 2935 1216 2936
rect 1207 2931 1208 2935
rect 1215 2931 1216 2935
rect 1207 2930 1216 2931
rect 1303 2935 1309 2936
rect 1303 2931 1304 2935
rect 1308 2934 1309 2935
rect 1511 2935 1517 2936
rect 1511 2934 1512 2935
rect 1308 2932 1512 2934
rect 1308 2931 1309 2932
rect 1303 2930 1309 2931
rect 1511 2931 1512 2932
rect 1516 2931 1517 2935
rect 1511 2930 1517 2931
rect 1670 2935 1676 2936
rect 1670 2931 1671 2935
rect 1675 2934 1676 2935
rect 1815 2935 1821 2936
rect 1815 2934 1816 2935
rect 1675 2932 1816 2934
rect 1675 2931 1676 2932
rect 1670 2930 1676 2931
rect 1815 2931 1816 2932
rect 1820 2931 1821 2935
rect 1815 2930 1821 2931
rect 2114 2929 2120 2930
rect 1974 2928 1980 2929
rect 1974 2924 1975 2928
rect 1979 2924 1980 2928
rect 2114 2925 2115 2929
rect 2119 2925 2120 2929
rect 2114 2924 2120 2925
rect 2314 2929 2320 2930
rect 2314 2925 2315 2929
rect 2319 2925 2320 2929
rect 2314 2924 2320 2925
rect 2514 2929 2520 2930
rect 2514 2925 2515 2929
rect 2519 2925 2520 2929
rect 2514 2924 2520 2925
rect 2714 2929 2720 2930
rect 2714 2925 2715 2929
rect 2719 2925 2720 2929
rect 2714 2924 2720 2925
rect 2906 2929 2912 2930
rect 2906 2925 2907 2929
rect 2911 2925 2912 2929
rect 2906 2924 2912 2925
rect 3106 2929 3112 2930
rect 3106 2925 3107 2929
rect 3111 2925 3112 2929
rect 3106 2924 3112 2925
rect 3306 2929 3312 2930
rect 3306 2925 3307 2929
rect 3311 2925 3312 2929
rect 3306 2924 3312 2925
rect 3798 2928 3804 2929
rect 3798 2924 3799 2928
rect 3803 2924 3804 2928
rect 1974 2923 1980 2924
rect 3798 2923 3804 2924
rect 2239 2919 2245 2920
rect 2239 2915 2240 2919
rect 2244 2918 2245 2919
rect 2250 2919 2256 2920
rect 2250 2918 2251 2919
rect 2244 2916 2251 2918
rect 2244 2915 2245 2916
rect 2239 2914 2245 2915
rect 2250 2915 2251 2916
rect 2255 2915 2256 2919
rect 2250 2914 2256 2915
rect 2274 2919 2280 2920
rect 2274 2915 2275 2919
rect 2279 2918 2280 2919
rect 2439 2919 2445 2920
rect 2439 2918 2440 2919
rect 2279 2916 2440 2918
rect 2279 2915 2280 2916
rect 2274 2914 2280 2915
rect 2439 2915 2440 2916
rect 2444 2915 2445 2919
rect 2439 2914 2445 2915
rect 2474 2919 2480 2920
rect 2474 2915 2475 2919
rect 2479 2918 2480 2919
rect 2639 2919 2645 2920
rect 2639 2918 2640 2919
rect 2479 2916 2640 2918
rect 2479 2915 2480 2916
rect 2474 2914 2480 2915
rect 2639 2915 2640 2916
rect 2644 2915 2645 2919
rect 2639 2914 2645 2915
rect 2838 2919 2845 2920
rect 2838 2915 2839 2919
rect 2844 2915 2845 2919
rect 2838 2914 2845 2915
rect 3030 2919 3037 2920
rect 3030 2915 3031 2919
rect 3036 2915 3037 2919
rect 3030 2914 3037 2915
rect 3066 2919 3072 2920
rect 3066 2915 3067 2919
rect 3071 2918 3072 2919
rect 3231 2919 3237 2920
rect 3231 2918 3232 2919
rect 3071 2916 3232 2918
rect 3071 2915 3072 2916
rect 3066 2914 3072 2915
rect 3231 2915 3232 2916
rect 3236 2915 3237 2919
rect 3231 2914 3237 2915
rect 3266 2919 3272 2920
rect 3266 2915 3267 2919
rect 3271 2918 3272 2919
rect 3431 2919 3437 2920
rect 3431 2918 3432 2919
rect 3271 2916 3432 2918
rect 3271 2915 3272 2916
rect 3266 2914 3272 2915
rect 3431 2915 3432 2916
rect 3436 2915 3437 2919
rect 3431 2914 3437 2915
rect 3838 2901 3844 2902
rect 5662 2901 5668 2902
rect 3838 2897 3839 2901
rect 3843 2897 3844 2901
rect 3838 2896 3844 2897
rect 3894 2900 3900 2901
rect 3894 2896 3895 2900
rect 3899 2896 3900 2900
rect 442 2895 448 2896
rect 442 2894 443 2895
rect 269 2892 443 2894
rect 442 2891 443 2892
rect 447 2891 448 2895
rect 722 2895 728 2896
rect 722 2894 723 2895
rect 581 2892 723 2894
rect 442 2890 448 2891
rect 722 2891 723 2892
rect 727 2891 728 2895
rect 1026 2895 1032 2896
rect 1026 2894 1027 2895
rect 885 2892 1027 2894
rect 722 2890 728 2891
rect 1026 2891 1027 2892
rect 1031 2891 1032 2895
rect 1303 2895 1309 2896
rect 1303 2894 1304 2895
rect 1181 2892 1304 2894
rect 1026 2890 1032 2891
rect 1303 2891 1304 2892
rect 1308 2891 1309 2895
rect 1670 2895 1676 2896
rect 1670 2894 1671 2895
rect 1485 2892 1671 2894
rect 1303 2890 1309 2891
rect 1670 2891 1671 2892
rect 1675 2891 1676 2895
rect 1906 2895 1912 2896
rect 3894 2895 3900 2896
rect 4030 2900 4036 2901
rect 4030 2896 4031 2900
rect 4035 2896 4036 2900
rect 4030 2895 4036 2896
rect 4166 2900 4172 2901
rect 4166 2896 4167 2900
rect 4171 2896 4172 2900
rect 4166 2895 4172 2896
rect 4302 2900 4308 2901
rect 4302 2896 4303 2900
rect 4307 2896 4308 2900
rect 4302 2895 4308 2896
rect 4438 2900 4444 2901
rect 4438 2896 4439 2900
rect 4443 2896 4444 2900
rect 4438 2895 4444 2896
rect 4574 2900 4580 2901
rect 4574 2896 4575 2900
rect 4579 2896 4580 2900
rect 5662 2897 5663 2901
rect 5667 2897 5668 2901
rect 5662 2896 5668 2897
rect 4574 2895 4580 2896
rect 1906 2894 1907 2895
rect 1789 2892 1907 2894
rect 1670 2890 1676 2891
rect 1906 2891 1907 2892
rect 1911 2891 1912 2895
rect 1906 2890 1912 2891
rect 3866 2885 3872 2886
rect 3838 2884 3844 2885
rect 3838 2880 3839 2884
rect 3843 2880 3844 2884
rect 3866 2881 3867 2885
rect 3871 2881 3872 2885
rect 3866 2880 3872 2881
rect 4002 2885 4008 2886
rect 4002 2881 4003 2885
rect 4007 2881 4008 2885
rect 4002 2880 4008 2881
rect 4138 2885 4144 2886
rect 4138 2881 4139 2885
rect 4143 2881 4144 2885
rect 4138 2880 4144 2881
rect 4274 2885 4280 2886
rect 4274 2881 4275 2885
rect 4279 2881 4280 2885
rect 4274 2880 4280 2881
rect 4410 2885 4416 2886
rect 4410 2881 4411 2885
rect 4415 2881 4416 2885
rect 4410 2880 4416 2881
rect 4546 2885 4552 2886
rect 4546 2881 4547 2885
rect 4551 2881 4552 2885
rect 4546 2880 4552 2881
rect 5662 2884 5668 2885
rect 5662 2880 5663 2884
rect 5667 2880 5668 2884
rect 2274 2879 2280 2880
rect 2274 2878 2275 2879
rect 2213 2876 2275 2878
rect 2274 2875 2275 2876
rect 2279 2875 2280 2879
rect 2474 2879 2480 2880
rect 2474 2878 2475 2879
rect 2413 2876 2475 2878
rect 2274 2874 2280 2875
rect 2474 2875 2475 2876
rect 2479 2875 2480 2879
rect 2474 2874 2480 2875
rect 2610 2879 2616 2880
rect 2610 2875 2611 2879
rect 2615 2875 2616 2879
rect 2610 2874 2616 2875
rect 2634 2879 2640 2880
rect 2634 2875 2635 2879
rect 2639 2878 2640 2879
rect 3066 2879 3072 2880
rect 3066 2878 3067 2879
rect 2639 2876 2721 2878
rect 3005 2876 3067 2878
rect 2639 2875 2640 2876
rect 2634 2874 2640 2875
rect 3066 2875 3067 2876
rect 3071 2875 3072 2879
rect 3266 2879 3272 2880
rect 3266 2878 3267 2879
rect 3205 2876 3267 2878
rect 3066 2874 3072 2875
rect 3266 2875 3267 2876
rect 3271 2875 3272 2879
rect 3266 2874 3272 2875
rect 3358 2879 3364 2880
rect 3838 2879 3844 2880
rect 5662 2879 5668 2880
rect 3358 2875 3359 2879
rect 3363 2875 3364 2879
rect 3358 2874 3364 2875
rect 3990 2875 3997 2876
rect 3990 2871 3991 2875
rect 3996 2871 3997 2875
rect 3990 2870 3997 2871
rect 4122 2875 4133 2876
rect 4122 2871 4123 2875
rect 4127 2871 4128 2875
rect 4132 2871 4133 2875
rect 4122 2870 4133 2871
rect 4135 2875 4141 2876
rect 4135 2871 4136 2875
rect 4140 2874 4141 2875
rect 4263 2875 4269 2876
rect 4263 2874 4264 2875
rect 4140 2872 4264 2874
rect 4140 2871 4141 2872
rect 4135 2870 4141 2871
rect 4263 2871 4264 2872
rect 4268 2871 4269 2875
rect 4263 2870 4269 2871
rect 4399 2875 4408 2876
rect 4399 2871 4400 2875
rect 4407 2871 4408 2875
rect 4399 2870 4408 2871
rect 4535 2875 4544 2876
rect 4535 2871 4536 2875
rect 4543 2871 4544 2875
rect 4671 2875 4677 2876
rect 4671 2874 4672 2875
rect 4535 2870 4544 2871
rect 4564 2872 4672 2874
rect 4234 2867 4240 2868
rect 298 2863 304 2864
rect 298 2862 299 2863
rect 229 2860 299 2862
rect 298 2859 299 2860
rect 303 2859 304 2863
rect 1210 2863 1216 2864
rect 298 2858 304 2859
rect 314 2859 320 2860
rect 314 2855 315 2859
rect 319 2855 320 2859
rect 314 2854 320 2855
rect 530 2859 536 2860
rect 530 2855 531 2859
rect 535 2855 536 2859
rect 530 2854 536 2855
rect 770 2859 776 2860
rect 770 2855 771 2859
rect 775 2855 776 2859
rect 770 2854 776 2855
rect 1018 2859 1024 2860
rect 1018 2855 1019 2859
rect 1023 2855 1024 2859
rect 1210 2859 1211 2863
rect 1215 2862 1216 2863
rect 4234 2863 4235 2867
rect 4239 2866 4240 2867
rect 4564 2866 4566 2872
rect 4671 2871 4672 2872
rect 4676 2871 4677 2875
rect 4671 2870 4677 2871
rect 4239 2864 4566 2866
rect 4239 2863 4240 2864
rect 4234 2862 4240 2863
rect 1215 2860 1281 2862
rect 1215 2859 1216 2860
rect 1210 2858 1216 2859
rect 1546 2859 1552 2860
rect 1018 2854 1024 2855
rect 1546 2855 1547 2859
rect 1551 2855 1552 2859
rect 1546 2854 1552 2855
rect 2154 2839 2160 2840
rect 2154 2838 2155 2839
rect 2109 2836 2155 2838
rect 2154 2835 2155 2836
rect 2159 2835 2160 2839
rect 2154 2834 2160 2835
rect 2250 2839 2256 2840
rect 2250 2835 2251 2839
rect 2255 2838 2256 2839
rect 2991 2839 2997 2840
rect 2991 2838 2992 2839
rect 2255 2836 2265 2838
rect 2853 2836 2992 2838
rect 2255 2835 2256 2836
rect 2250 2834 2256 2835
rect 2514 2835 2520 2836
rect 2514 2831 2515 2835
rect 2519 2831 2520 2835
rect 2991 2835 2992 2836
rect 2996 2835 2997 2839
rect 2991 2834 2997 2835
rect 3030 2839 3036 2840
rect 3030 2835 3031 2839
rect 3035 2835 3036 2839
rect 3030 2834 3036 2835
rect 3962 2835 3968 2836
rect 2514 2830 2520 2831
rect 3962 2831 3963 2835
rect 3967 2831 3968 2835
rect 4135 2835 4141 2836
rect 4135 2834 4136 2835
rect 4101 2832 4136 2834
rect 3962 2830 3968 2831
rect 4135 2831 4136 2832
rect 4140 2831 4141 2835
rect 4135 2830 4141 2831
rect 4234 2835 4240 2836
rect 4234 2831 4235 2835
rect 4239 2831 4240 2835
rect 4234 2830 4240 2831
rect 4366 2835 4372 2836
rect 4366 2831 4367 2835
rect 4371 2831 4372 2835
rect 4366 2830 4372 2831
rect 4402 2835 4408 2836
rect 4402 2831 4403 2835
rect 4407 2834 4408 2835
rect 4538 2835 4544 2836
rect 4407 2832 4417 2834
rect 4407 2831 4408 2832
rect 4402 2830 4408 2831
rect 4538 2831 4539 2835
rect 4543 2834 4544 2835
rect 4543 2832 4553 2834
rect 4543 2831 4544 2832
rect 4538 2830 4544 2831
rect 255 2819 261 2820
rect 255 2815 256 2819
rect 260 2818 261 2819
rect 314 2819 320 2820
rect 314 2818 315 2819
rect 260 2816 315 2818
rect 260 2815 261 2816
rect 255 2814 261 2815
rect 314 2815 315 2816
rect 319 2815 320 2819
rect 314 2814 320 2815
rect 431 2819 437 2820
rect 431 2815 432 2819
rect 436 2818 437 2819
rect 530 2819 536 2820
rect 530 2818 531 2819
rect 436 2816 531 2818
rect 436 2815 437 2816
rect 431 2814 437 2815
rect 530 2815 531 2816
rect 535 2815 536 2819
rect 530 2814 536 2815
rect 647 2819 653 2820
rect 647 2815 648 2819
rect 652 2818 653 2819
rect 770 2819 776 2820
rect 770 2818 771 2819
rect 652 2816 771 2818
rect 652 2815 653 2816
rect 647 2814 653 2815
rect 770 2815 771 2816
rect 775 2815 776 2819
rect 770 2814 776 2815
rect 887 2819 893 2820
rect 887 2815 888 2819
rect 892 2818 893 2819
rect 1018 2819 1024 2820
rect 1018 2818 1019 2819
rect 892 2816 1019 2818
rect 892 2815 893 2816
rect 887 2814 893 2815
rect 1018 2815 1019 2816
rect 1023 2815 1024 2819
rect 1018 2814 1024 2815
rect 1026 2819 1032 2820
rect 1026 2815 1027 2819
rect 1031 2818 1032 2819
rect 1135 2819 1141 2820
rect 1135 2818 1136 2819
rect 1031 2816 1136 2818
rect 1031 2815 1032 2816
rect 1026 2814 1032 2815
rect 1135 2815 1136 2816
rect 1140 2815 1141 2819
rect 1135 2814 1141 2815
rect 1399 2819 1405 2820
rect 1399 2815 1400 2819
rect 1404 2818 1405 2819
rect 1546 2819 1552 2820
rect 1546 2818 1547 2819
rect 1404 2816 1547 2818
rect 1404 2815 1405 2816
rect 1399 2814 1405 2815
rect 1546 2815 1547 2816
rect 1551 2815 1552 2819
rect 1546 2814 1552 2815
rect 1618 2819 1624 2820
rect 1618 2815 1619 2819
rect 1623 2818 1624 2819
rect 1663 2819 1669 2820
rect 1663 2818 1664 2819
rect 1623 2816 1664 2818
rect 1623 2815 1624 2816
rect 1618 2814 1624 2815
rect 1663 2815 1664 2816
rect 1668 2815 1669 2819
rect 1663 2814 1669 2815
rect 110 2812 116 2813
rect 1934 2812 1940 2813
rect 110 2808 111 2812
rect 115 2808 116 2812
rect 110 2807 116 2808
rect 130 2811 136 2812
rect 130 2807 131 2811
rect 135 2807 136 2811
rect 130 2806 136 2807
rect 306 2811 312 2812
rect 306 2807 307 2811
rect 311 2807 312 2811
rect 306 2806 312 2807
rect 522 2811 528 2812
rect 522 2807 523 2811
rect 527 2807 528 2811
rect 522 2806 528 2807
rect 762 2811 768 2812
rect 762 2807 763 2811
rect 767 2807 768 2811
rect 762 2806 768 2807
rect 1010 2811 1016 2812
rect 1010 2807 1011 2811
rect 1015 2807 1016 2811
rect 1010 2806 1016 2807
rect 1274 2811 1280 2812
rect 1274 2807 1275 2811
rect 1279 2807 1280 2811
rect 1274 2806 1280 2807
rect 1538 2811 1544 2812
rect 1538 2807 1539 2811
rect 1543 2807 1544 2811
rect 1934 2808 1935 2812
rect 1939 2808 1940 2812
rect 1934 2807 1940 2808
rect 1538 2806 1544 2807
rect 158 2796 164 2797
rect 110 2795 116 2796
rect 110 2791 111 2795
rect 115 2791 116 2795
rect 158 2792 159 2796
rect 163 2792 164 2796
rect 158 2791 164 2792
rect 334 2796 340 2797
rect 334 2792 335 2796
rect 339 2792 340 2796
rect 334 2791 340 2792
rect 550 2796 556 2797
rect 550 2792 551 2796
rect 555 2792 556 2796
rect 550 2791 556 2792
rect 790 2796 796 2797
rect 790 2792 791 2796
rect 795 2792 796 2796
rect 790 2791 796 2792
rect 1038 2796 1044 2797
rect 1038 2792 1039 2796
rect 1043 2792 1044 2796
rect 1038 2791 1044 2792
rect 1302 2796 1308 2797
rect 1302 2792 1303 2796
rect 1307 2792 1308 2796
rect 1302 2791 1308 2792
rect 1566 2796 1572 2797
rect 1566 2792 1567 2796
rect 1571 2792 1572 2796
rect 1566 2791 1572 2792
rect 1934 2795 1940 2796
rect 1934 2791 1935 2795
rect 1939 2791 1940 2795
rect 110 2790 116 2791
rect 1934 2790 1940 2791
rect 2090 2795 2096 2796
rect 2090 2791 2091 2795
rect 2095 2794 2096 2795
rect 2135 2795 2141 2796
rect 2135 2794 2136 2795
rect 2095 2792 2136 2794
rect 2095 2791 2096 2792
rect 2090 2790 2096 2791
rect 2135 2791 2136 2792
rect 2140 2791 2141 2795
rect 2135 2790 2141 2791
rect 2154 2795 2160 2796
rect 2154 2791 2155 2795
rect 2159 2794 2160 2795
rect 2383 2795 2389 2796
rect 2383 2794 2384 2795
rect 2159 2792 2384 2794
rect 2159 2791 2160 2792
rect 2154 2790 2160 2791
rect 2383 2791 2384 2792
rect 2388 2791 2389 2795
rect 2383 2790 2389 2791
rect 2631 2795 2640 2796
rect 2631 2791 2632 2795
rect 2639 2791 2640 2795
rect 2631 2790 2640 2791
rect 2806 2795 2812 2796
rect 2806 2791 2807 2795
rect 2811 2794 2812 2795
rect 2879 2795 2885 2796
rect 2879 2794 2880 2795
rect 2811 2792 2880 2794
rect 2811 2791 2812 2792
rect 2806 2790 2812 2791
rect 2879 2791 2880 2792
rect 2884 2791 2885 2795
rect 2879 2790 2885 2791
rect 2999 2795 3005 2796
rect 2999 2791 3000 2795
rect 3004 2794 3005 2795
rect 3127 2795 3133 2796
rect 3127 2794 3128 2795
rect 3004 2792 3128 2794
rect 3004 2791 3005 2792
rect 2999 2790 3005 2791
rect 3127 2791 3128 2792
rect 3132 2791 3133 2795
rect 3991 2795 3997 2796
rect 3991 2794 3992 2795
rect 3957 2792 3992 2794
rect 3127 2790 3133 2791
rect 3991 2791 3992 2792
rect 3996 2791 3997 2795
rect 3991 2790 3997 2791
rect 4054 2795 4060 2796
rect 4054 2791 4055 2795
rect 4059 2791 4060 2795
rect 4054 2790 4060 2791
rect 4122 2795 4128 2796
rect 4122 2791 4123 2795
rect 4127 2794 4128 2795
rect 4127 2792 4137 2794
rect 4127 2791 4128 2792
rect 4122 2790 4128 2791
rect 4274 2791 4280 2792
rect 1974 2788 1980 2789
rect 3798 2788 3804 2789
rect 1974 2784 1975 2788
rect 1979 2784 1980 2788
rect 1974 2783 1980 2784
rect 2010 2787 2016 2788
rect 2010 2783 2011 2787
rect 2015 2783 2016 2787
rect 2010 2782 2016 2783
rect 2258 2787 2264 2788
rect 2258 2783 2259 2787
rect 2263 2783 2264 2787
rect 2258 2782 2264 2783
rect 2506 2787 2512 2788
rect 2506 2783 2507 2787
rect 2511 2783 2512 2787
rect 2506 2782 2512 2783
rect 2754 2787 2760 2788
rect 2754 2783 2755 2787
rect 2759 2783 2760 2787
rect 2754 2782 2760 2783
rect 3002 2787 3008 2788
rect 3002 2783 3003 2787
rect 3007 2783 3008 2787
rect 3798 2784 3799 2788
rect 3803 2784 3804 2788
rect 4274 2787 4275 2791
rect 4279 2787 4280 2791
rect 4274 2786 4280 2787
rect 4410 2791 4416 2792
rect 4410 2787 4411 2791
rect 4415 2787 4416 2791
rect 4410 2786 4416 2787
rect 4546 2791 4552 2792
rect 4546 2787 4547 2791
rect 4551 2787 4552 2791
rect 4546 2786 4552 2787
rect 4682 2791 4688 2792
rect 4682 2787 4683 2791
rect 4687 2787 4688 2791
rect 4682 2786 4688 2787
rect 4818 2791 4824 2792
rect 4818 2787 4819 2791
rect 4823 2787 4824 2791
rect 4818 2786 4824 2787
rect 3798 2783 3804 2784
rect 3002 2782 3008 2783
rect 2038 2772 2044 2773
rect 1974 2771 1980 2772
rect 1974 2767 1975 2771
rect 1979 2767 1980 2771
rect 2038 2768 2039 2772
rect 2043 2768 2044 2772
rect 2038 2767 2044 2768
rect 2286 2772 2292 2773
rect 2286 2768 2287 2772
rect 2291 2768 2292 2772
rect 2286 2767 2292 2768
rect 2534 2772 2540 2773
rect 2534 2768 2535 2772
rect 2539 2768 2540 2772
rect 2534 2767 2540 2768
rect 2782 2772 2788 2773
rect 2782 2768 2783 2772
rect 2787 2768 2788 2772
rect 2782 2767 2788 2768
rect 3030 2772 3036 2773
rect 3030 2768 3031 2772
rect 3035 2768 3036 2772
rect 3030 2767 3036 2768
rect 3798 2771 3804 2772
rect 3798 2767 3799 2771
rect 3803 2767 3804 2771
rect 1974 2766 1980 2767
rect 3798 2766 3804 2767
rect 3962 2751 3968 2752
rect 3962 2747 3963 2751
rect 3967 2750 3968 2751
rect 3983 2751 3989 2752
rect 3983 2750 3984 2751
rect 3967 2748 3984 2750
rect 3967 2747 3968 2748
rect 3962 2746 3968 2747
rect 3983 2747 3984 2748
rect 3988 2747 3989 2751
rect 3983 2746 3989 2747
rect 3991 2751 3997 2752
rect 3991 2747 3992 2751
rect 3996 2750 3997 2751
rect 4119 2751 4125 2752
rect 4119 2750 4120 2751
rect 3996 2748 4120 2750
rect 3996 2747 3997 2748
rect 3991 2746 3997 2747
rect 4119 2747 4120 2748
rect 4124 2747 4125 2751
rect 4119 2746 4125 2747
rect 4255 2751 4261 2752
rect 4255 2747 4256 2751
rect 4260 2750 4261 2751
rect 4274 2751 4280 2752
rect 4274 2750 4275 2751
rect 4260 2748 4275 2750
rect 4260 2747 4261 2748
rect 4255 2746 4261 2747
rect 4274 2747 4275 2748
rect 4279 2747 4280 2751
rect 4274 2746 4280 2747
rect 4391 2751 4397 2752
rect 4391 2747 4392 2751
rect 4396 2750 4397 2751
rect 4410 2751 4416 2752
rect 4410 2750 4411 2751
rect 4396 2748 4411 2750
rect 4396 2747 4397 2748
rect 4391 2746 4397 2747
rect 4410 2747 4411 2748
rect 4415 2747 4416 2751
rect 4410 2746 4416 2747
rect 4527 2751 4533 2752
rect 4527 2747 4528 2751
rect 4532 2750 4533 2751
rect 4546 2751 4552 2752
rect 4546 2750 4547 2751
rect 4532 2748 4547 2750
rect 4532 2747 4533 2748
rect 4527 2746 4533 2747
rect 4546 2747 4547 2748
rect 4551 2747 4552 2751
rect 4546 2746 4552 2747
rect 4663 2751 4669 2752
rect 4663 2747 4664 2751
rect 4668 2750 4669 2751
rect 4682 2751 4688 2752
rect 4682 2750 4683 2751
rect 4668 2748 4683 2750
rect 4668 2747 4669 2748
rect 4663 2746 4669 2747
rect 4682 2747 4683 2748
rect 4687 2747 4688 2751
rect 4682 2746 4688 2747
rect 4799 2751 4805 2752
rect 4799 2747 4800 2751
rect 4804 2750 4805 2751
rect 4818 2751 4824 2752
rect 4818 2750 4819 2751
rect 4804 2748 4819 2750
rect 4804 2747 4805 2748
rect 4799 2746 4805 2747
rect 4818 2747 4819 2748
rect 4823 2747 4824 2751
rect 4818 2746 4824 2747
rect 4830 2751 4836 2752
rect 4830 2747 4831 2751
rect 4835 2750 4836 2751
rect 4935 2751 4941 2752
rect 4935 2750 4936 2751
rect 4835 2748 4936 2750
rect 4835 2747 4836 2748
rect 4830 2746 4836 2747
rect 4935 2747 4936 2748
rect 4940 2747 4941 2751
rect 4935 2746 4941 2747
rect 3838 2744 3844 2745
rect 5662 2744 5668 2745
rect 3838 2740 3839 2744
rect 3843 2740 3844 2744
rect 3838 2739 3844 2740
rect 3858 2743 3864 2744
rect 3858 2739 3859 2743
rect 3863 2739 3864 2743
rect 3858 2738 3864 2739
rect 3994 2743 4000 2744
rect 3994 2739 3995 2743
rect 3999 2739 4000 2743
rect 3994 2738 4000 2739
rect 4130 2743 4136 2744
rect 4130 2739 4131 2743
rect 4135 2739 4136 2743
rect 4130 2738 4136 2739
rect 4266 2743 4272 2744
rect 4266 2739 4267 2743
rect 4271 2739 4272 2743
rect 4266 2738 4272 2739
rect 4402 2743 4408 2744
rect 4402 2739 4403 2743
rect 4407 2739 4408 2743
rect 4402 2738 4408 2739
rect 4538 2743 4544 2744
rect 4538 2739 4539 2743
rect 4543 2739 4544 2743
rect 4538 2738 4544 2739
rect 4674 2743 4680 2744
rect 4674 2739 4675 2743
rect 4679 2739 4680 2743
rect 4674 2738 4680 2739
rect 4810 2743 4816 2744
rect 4810 2739 4811 2743
rect 4815 2739 4816 2743
rect 5662 2740 5663 2744
rect 5667 2740 5668 2744
rect 5662 2739 5668 2740
rect 4810 2738 4816 2739
rect 110 2733 116 2734
rect 1934 2733 1940 2734
rect 110 2729 111 2733
rect 115 2729 116 2733
rect 110 2728 116 2729
rect 278 2732 284 2733
rect 278 2728 279 2732
rect 283 2728 284 2732
rect 278 2727 284 2728
rect 454 2732 460 2733
rect 454 2728 455 2732
rect 459 2728 460 2732
rect 454 2727 460 2728
rect 646 2732 652 2733
rect 646 2728 647 2732
rect 651 2728 652 2732
rect 646 2727 652 2728
rect 854 2732 860 2733
rect 854 2728 855 2732
rect 859 2728 860 2732
rect 854 2727 860 2728
rect 1078 2732 1084 2733
rect 1078 2728 1079 2732
rect 1083 2728 1084 2732
rect 1078 2727 1084 2728
rect 1310 2732 1316 2733
rect 1310 2728 1311 2732
rect 1315 2728 1316 2732
rect 1310 2727 1316 2728
rect 1550 2732 1556 2733
rect 1550 2728 1551 2732
rect 1555 2728 1556 2732
rect 1550 2727 1556 2728
rect 1798 2732 1804 2733
rect 1798 2728 1799 2732
rect 1803 2728 1804 2732
rect 1934 2729 1935 2733
rect 1939 2729 1940 2733
rect 1934 2728 1940 2729
rect 3886 2728 3892 2729
rect 1798 2727 1804 2728
rect 3838 2727 3844 2728
rect 3838 2723 3839 2727
rect 3843 2723 3844 2727
rect 3886 2724 3887 2728
rect 3891 2724 3892 2728
rect 3886 2723 3892 2724
rect 4022 2728 4028 2729
rect 4022 2724 4023 2728
rect 4027 2724 4028 2728
rect 4022 2723 4028 2724
rect 4158 2728 4164 2729
rect 4158 2724 4159 2728
rect 4163 2724 4164 2728
rect 4158 2723 4164 2724
rect 4294 2728 4300 2729
rect 4294 2724 4295 2728
rect 4299 2724 4300 2728
rect 4294 2723 4300 2724
rect 4430 2728 4436 2729
rect 4430 2724 4431 2728
rect 4435 2724 4436 2728
rect 4430 2723 4436 2724
rect 4566 2728 4572 2729
rect 4566 2724 4567 2728
rect 4571 2724 4572 2728
rect 4566 2723 4572 2724
rect 4702 2728 4708 2729
rect 4702 2724 4703 2728
rect 4707 2724 4708 2728
rect 4702 2723 4708 2724
rect 4838 2728 4844 2729
rect 4838 2724 4839 2728
rect 4843 2724 4844 2728
rect 4838 2723 4844 2724
rect 5662 2727 5668 2728
rect 5662 2723 5663 2727
rect 5667 2723 5668 2727
rect 3838 2722 3844 2723
rect 5662 2722 5668 2723
rect 250 2717 256 2718
rect 110 2716 116 2717
rect 110 2712 111 2716
rect 115 2712 116 2716
rect 250 2713 251 2717
rect 255 2713 256 2717
rect 250 2712 256 2713
rect 426 2717 432 2718
rect 426 2713 427 2717
rect 431 2713 432 2717
rect 426 2712 432 2713
rect 618 2717 624 2718
rect 618 2713 619 2717
rect 623 2713 624 2717
rect 618 2712 624 2713
rect 826 2717 832 2718
rect 826 2713 827 2717
rect 831 2713 832 2717
rect 826 2712 832 2713
rect 1050 2717 1056 2718
rect 1050 2713 1051 2717
rect 1055 2713 1056 2717
rect 1050 2712 1056 2713
rect 1282 2717 1288 2718
rect 1282 2713 1283 2717
rect 1287 2713 1288 2717
rect 1282 2712 1288 2713
rect 1522 2717 1528 2718
rect 1522 2713 1523 2717
rect 1527 2713 1528 2717
rect 1522 2712 1528 2713
rect 1770 2717 1776 2718
rect 1770 2713 1771 2717
rect 1775 2713 1776 2717
rect 1770 2712 1776 2713
rect 1934 2716 1940 2717
rect 1934 2712 1935 2716
rect 1939 2712 1940 2716
rect 110 2711 116 2712
rect 1934 2711 1940 2712
rect 1974 2709 1980 2710
rect 3798 2709 3804 2710
rect 298 2707 304 2708
rect 298 2703 299 2707
rect 303 2706 304 2707
rect 375 2707 381 2708
rect 375 2706 376 2707
rect 303 2704 376 2706
rect 303 2703 304 2704
rect 298 2702 304 2703
rect 375 2703 376 2704
rect 380 2703 381 2707
rect 375 2702 381 2703
rect 406 2707 412 2708
rect 406 2703 407 2707
rect 411 2706 412 2707
rect 551 2707 557 2708
rect 551 2706 552 2707
rect 411 2704 552 2706
rect 411 2703 412 2704
rect 406 2702 412 2703
rect 551 2703 552 2704
rect 556 2703 557 2707
rect 551 2702 557 2703
rect 583 2707 589 2708
rect 583 2703 584 2707
rect 588 2706 589 2707
rect 743 2707 749 2708
rect 743 2706 744 2707
rect 588 2704 744 2706
rect 588 2703 589 2704
rect 583 2702 589 2703
rect 743 2703 744 2704
rect 748 2703 749 2707
rect 743 2702 749 2703
rect 823 2707 829 2708
rect 823 2703 824 2707
rect 828 2706 829 2707
rect 951 2707 957 2708
rect 951 2706 952 2707
rect 828 2704 952 2706
rect 828 2703 829 2704
rect 823 2702 829 2703
rect 951 2703 952 2704
rect 956 2703 957 2707
rect 951 2702 957 2703
rect 975 2707 981 2708
rect 975 2703 976 2707
rect 980 2706 981 2707
rect 1175 2707 1181 2708
rect 1175 2706 1176 2707
rect 980 2704 1176 2706
rect 980 2703 981 2704
rect 975 2702 981 2703
rect 1175 2703 1176 2704
rect 1180 2703 1181 2707
rect 1175 2702 1181 2703
rect 1406 2707 1413 2708
rect 1406 2703 1407 2707
rect 1412 2703 1413 2707
rect 1406 2702 1413 2703
rect 1519 2707 1525 2708
rect 1519 2703 1520 2707
rect 1524 2706 1525 2707
rect 1647 2707 1653 2708
rect 1647 2706 1648 2707
rect 1524 2704 1648 2706
rect 1524 2703 1525 2704
rect 1519 2702 1525 2703
rect 1647 2703 1648 2704
rect 1652 2703 1653 2707
rect 1647 2702 1653 2703
rect 1786 2707 1792 2708
rect 1786 2703 1787 2707
rect 1791 2706 1792 2707
rect 1895 2707 1901 2708
rect 1895 2706 1896 2707
rect 1791 2704 1896 2706
rect 1791 2703 1792 2704
rect 1786 2702 1792 2703
rect 1895 2703 1896 2704
rect 1900 2703 1901 2707
rect 1974 2705 1975 2709
rect 1979 2705 1980 2709
rect 1974 2704 1980 2705
rect 2022 2708 2028 2709
rect 2022 2704 2023 2708
rect 2027 2704 2028 2708
rect 2022 2703 2028 2704
rect 2246 2708 2252 2709
rect 2246 2704 2247 2708
rect 2251 2704 2252 2708
rect 2246 2703 2252 2704
rect 2502 2708 2508 2709
rect 2502 2704 2503 2708
rect 2507 2704 2508 2708
rect 2502 2703 2508 2704
rect 2758 2708 2764 2709
rect 2758 2704 2759 2708
rect 2763 2704 2764 2708
rect 2758 2703 2764 2704
rect 3014 2708 3020 2709
rect 3014 2704 3015 2708
rect 3019 2704 3020 2708
rect 3798 2705 3799 2709
rect 3803 2705 3804 2709
rect 3798 2704 3804 2705
rect 3014 2703 3020 2704
rect 1895 2702 1901 2703
rect 1994 2693 2000 2694
rect 1974 2692 1980 2693
rect 1974 2688 1975 2692
rect 1979 2688 1980 2692
rect 1994 2689 1995 2693
rect 1999 2689 2000 2693
rect 1994 2688 2000 2689
rect 2218 2693 2224 2694
rect 2218 2689 2219 2693
rect 2223 2689 2224 2693
rect 2218 2688 2224 2689
rect 2474 2693 2480 2694
rect 2474 2689 2475 2693
rect 2479 2689 2480 2693
rect 2474 2688 2480 2689
rect 2730 2693 2736 2694
rect 2730 2689 2731 2693
rect 2735 2689 2736 2693
rect 2730 2688 2736 2689
rect 2986 2693 2992 2694
rect 2986 2689 2987 2693
rect 2991 2689 2992 2693
rect 2986 2688 2992 2689
rect 3798 2692 3804 2693
rect 3798 2688 3799 2692
rect 3803 2688 3804 2692
rect 1974 2687 1980 2688
rect 3798 2687 3804 2688
rect 2119 2683 2125 2684
rect 2119 2682 2120 2683
rect 1939 2680 2120 2682
rect 406 2667 412 2668
rect 406 2666 407 2667
rect 349 2664 407 2666
rect 406 2663 407 2664
rect 411 2663 412 2667
rect 583 2667 589 2668
rect 583 2666 584 2667
rect 525 2664 584 2666
rect 406 2662 412 2663
rect 583 2663 584 2664
rect 588 2663 589 2667
rect 823 2667 829 2668
rect 823 2666 824 2667
rect 717 2664 824 2666
rect 583 2662 589 2663
rect 823 2663 824 2664
rect 828 2663 829 2667
rect 975 2667 981 2668
rect 975 2666 976 2667
rect 925 2664 976 2666
rect 823 2662 829 2663
rect 975 2663 976 2664
rect 980 2663 981 2667
rect 975 2662 981 2663
rect 1018 2667 1024 2668
rect 1018 2663 1019 2667
rect 1023 2666 1024 2667
rect 1519 2667 1525 2668
rect 1519 2666 1520 2667
rect 1023 2664 1057 2666
rect 1381 2664 1520 2666
rect 1023 2663 1024 2664
rect 1018 2662 1024 2663
rect 1519 2663 1520 2664
rect 1524 2663 1525 2667
rect 1519 2662 1525 2663
rect 1618 2667 1624 2668
rect 1618 2663 1619 2667
rect 1623 2663 1624 2667
rect 1939 2666 1941 2680
rect 2119 2679 2120 2680
rect 2124 2679 2125 2683
rect 2119 2678 2125 2679
rect 2343 2683 2349 2684
rect 2343 2679 2344 2683
rect 2348 2682 2349 2683
rect 2514 2683 2520 2684
rect 2514 2682 2515 2683
rect 2348 2680 2515 2682
rect 2348 2679 2349 2680
rect 2343 2678 2349 2679
rect 2514 2679 2515 2680
rect 2519 2679 2520 2683
rect 2514 2678 2520 2679
rect 2599 2683 2608 2684
rect 2599 2679 2600 2683
rect 2607 2679 2608 2683
rect 2599 2678 2608 2679
rect 2855 2683 2864 2684
rect 2855 2679 2856 2683
rect 2863 2679 2864 2683
rect 2855 2678 2864 2679
rect 3110 2683 3117 2684
rect 3110 2679 3111 2683
rect 3116 2679 3117 2683
rect 3110 2678 3117 2679
rect 1869 2664 1941 2666
rect 3838 2669 3844 2670
rect 5662 2669 5668 2670
rect 3838 2665 3839 2669
rect 3843 2665 3844 2669
rect 3838 2664 3844 2665
rect 3958 2668 3964 2669
rect 3958 2664 3959 2668
rect 3963 2664 3964 2668
rect 3958 2663 3964 2664
rect 4254 2668 4260 2669
rect 4254 2664 4255 2668
rect 4259 2664 4260 2668
rect 4254 2663 4260 2664
rect 4542 2668 4548 2669
rect 4542 2664 4543 2668
rect 4547 2664 4548 2668
rect 4542 2663 4548 2664
rect 4822 2668 4828 2669
rect 4822 2664 4823 2668
rect 4827 2664 4828 2668
rect 4822 2663 4828 2664
rect 5110 2668 5116 2669
rect 5110 2664 5111 2668
rect 5115 2664 5116 2668
rect 5110 2663 5116 2664
rect 5398 2668 5404 2669
rect 5398 2664 5399 2668
rect 5403 2664 5404 2668
rect 5662 2665 5663 2669
rect 5667 2665 5668 2669
rect 5662 2664 5668 2665
rect 5398 2663 5404 2664
rect 1618 2662 1624 2663
rect 3930 2653 3936 2654
rect 3838 2652 3844 2653
rect 3838 2648 3839 2652
rect 3843 2648 3844 2652
rect 3930 2649 3931 2653
rect 3935 2649 3936 2653
rect 3930 2648 3936 2649
rect 4226 2653 4232 2654
rect 4226 2649 4227 2653
rect 4231 2649 4232 2653
rect 4226 2648 4232 2649
rect 4514 2653 4520 2654
rect 4514 2649 4515 2653
rect 4519 2649 4520 2653
rect 4514 2648 4520 2649
rect 4794 2653 4800 2654
rect 4794 2649 4795 2653
rect 4799 2649 4800 2653
rect 4794 2648 4800 2649
rect 5082 2653 5088 2654
rect 5082 2649 5083 2653
rect 5087 2649 5088 2653
rect 5082 2648 5088 2649
rect 5370 2653 5376 2654
rect 5370 2649 5371 2653
rect 5375 2649 5376 2653
rect 5370 2648 5376 2649
rect 5662 2652 5668 2653
rect 5662 2648 5663 2652
rect 5667 2648 5668 2652
rect 3838 2647 3844 2648
rect 5662 2647 5668 2648
rect 2090 2643 2096 2644
rect 882 2639 888 2640
rect 882 2638 883 2639
rect 732 2636 883 2638
rect 732 2634 734 2636
rect 882 2635 883 2636
rect 887 2635 888 2639
rect 2090 2639 2091 2643
rect 2095 2639 2096 2643
rect 2602 2643 2608 2644
rect 2090 2638 2096 2639
rect 882 2634 888 2635
rect 1186 2635 1192 2636
rect 1186 2634 1187 2635
rect 669 2632 734 2634
rect 1141 2632 1187 2634
rect 738 2631 744 2632
rect 738 2627 739 2631
rect 743 2627 744 2631
rect 738 2626 744 2627
rect 898 2631 904 2632
rect 898 2627 899 2631
rect 903 2627 904 2631
rect 1186 2631 1187 2632
rect 1191 2631 1192 2635
rect 1351 2635 1357 2636
rect 1351 2634 1352 2635
rect 1293 2632 1352 2634
rect 1186 2630 1192 2631
rect 1351 2631 1352 2632
rect 1356 2631 1357 2635
rect 1351 2630 1357 2631
rect 1406 2635 1412 2636
rect 1406 2631 1407 2635
rect 1411 2631 1412 2635
rect 1671 2635 1677 2636
rect 1671 2634 1672 2635
rect 1613 2632 1672 2634
rect 1406 2630 1412 2631
rect 1671 2631 1672 2632
rect 1676 2631 1677 2635
rect 1786 2635 1792 2636
rect 1786 2634 1787 2635
rect 1773 2632 1787 2634
rect 1671 2630 1677 2631
rect 1786 2631 1787 2632
rect 1791 2631 1792 2635
rect 2316 2634 2318 2641
rect 2538 2635 2544 2636
rect 2538 2634 2539 2635
rect 2316 2632 2539 2634
rect 1786 2630 1792 2631
rect 2538 2631 2539 2632
rect 2543 2631 2544 2635
rect 2572 2634 2574 2641
rect 2602 2639 2603 2643
rect 2607 2642 2608 2643
rect 2858 2643 2864 2644
rect 2607 2640 2737 2642
rect 2607 2639 2608 2640
rect 2602 2638 2608 2639
rect 2858 2639 2859 2643
rect 2863 2642 2864 2643
rect 4054 2643 4061 2644
rect 2863 2640 2993 2642
rect 2863 2639 2864 2640
rect 2858 2638 2864 2639
rect 4054 2639 4055 2643
rect 4060 2639 4061 2643
rect 4054 2638 4061 2639
rect 4351 2643 4357 2644
rect 4351 2639 4352 2643
rect 4356 2642 4357 2643
rect 4442 2643 4448 2644
rect 4442 2642 4443 2643
rect 4356 2640 4443 2642
rect 4356 2639 4357 2640
rect 4351 2638 4357 2639
rect 4442 2639 4443 2640
rect 4447 2639 4448 2643
rect 4442 2638 4448 2639
rect 4638 2643 4645 2644
rect 4638 2639 4639 2643
rect 4644 2639 4645 2643
rect 4638 2638 4645 2639
rect 4919 2643 4925 2644
rect 4919 2639 4920 2643
rect 4924 2642 4925 2643
rect 4974 2643 4980 2644
rect 4974 2642 4975 2643
rect 4924 2640 4975 2642
rect 4924 2639 4925 2640
rect 4919 2638 4925 2639
rect 4974 2639 4975 2640
rect 4979 2639 4980 2643
rect 4974 2638 4980 2639
rect 5207 2643 5213 2644
rect 5207 2639 5208 2643
rect 5212 2642 5213 2643
rect 5266 2643 5272 2644
rect 5266 2642 5267 2643
rect 5212 2640 5267 2642
rect 5212 2639 5213 2640
rect 5207 2638 5213 2639
rect 5266 2639 5267 2640
rect 5271 2639 5272 2643
rect 5266 2638 5272 2639
rect 5418 2643 5424 2644
rect 5418 2639 5419 2643
rect 5423 2642 5424 2643
rect 5495 2643 5501 2644
rect 5495 2642 5496 2643
rect 5423 2640 5496 2642
rect 5423 2639 5424 2640
rect 5418 2638 5424 2639
rect 5495 2639 5496 2640
rect 5500 2639 5501 2643
rect 5495 2638 5501 2639
rect 2806 2635 2812 2636
rect 2806 2634 2807 2635
rect 2572 2632 2807 2634
rect 2538 2630 2544 2631
rect 2806 2631 2807 2632
rect 2811 2631 2812 2635
rect 2806 2630 2812 2631
rect 898 2626 904 2627
rect 4322 2627 4328 2628
rect 4322 2623 4323 2627
rect 4327 2626 4328 2627
rect 4830 2627 4836 2628
rect 4830 2626 4831 2627
rect 4327 2624 4831 2626
rect 4327 2623 4328 2624
rect 4322 2622 4328 2623
rect 4830 2623 4831 2624
rect 4835 2623 4836 2627
rect 4830 2622 4836 2623
rect 3982 2603 3988 2604
rect 2687 2599 2693 2600
rect 2687 2598 2688 2599
rect 2653 2596 2688 2598
rect 2687 2595 2688 2596
rect 2692 2595 2693 2599
rect 2687 2594 2693 2595
rect 2774 2599 2780 2600
rect 2774 2595 2775 2599
rect 2779 2595 2780 2599
rect 2959 2599 2965 2600
rect 2959 2598 2960 2599
rect 2925 2596 2960 2598
rect 2774 2594 2780 2595
rect 2959 2595 2960 2596
rect 2964 2595 2965 2599
rect 3095 2599 3101 2600
rect 3095 2598 3096 2599
rect 3061 2596 3096 2598
rect 2959 2594 2965 2595
rect 3095 2595 3096 2596
rect 3100 2595 3101 2599
rect 3095 2594 3101 2595
rect 3110 2599 3116 2600
rect 3110 2595 3111 2599
rect 3115 2595 3116 2599
rect 3982 2599 3983 2603
rect 3987 2599 3988 2603
rect 3982 2598 3988 2599
rect 4322 2603 4328 2604
rect 4322 2599 4323 2603
rect 4327 2599 4328 2603
rect 4322 2598 4328 2599
rect 4442 2603 4448 2604
rect 4442 2599 4443 2603
rect 4447 2602 4448 2603
rect 4890 2603 4896 2604
rect 4447 2600 4521 2602
rect 4447 2599 4448 2600
rect 4442 2598 4448 2599
rect 4890 2599 4891 2603
rect 4895 2599 4896 2603
rect 4890 2598 4896 2599
rect 4974 2603 4980 2604
rect 4974 2599 4975 2603
rect 4979 2602 4980 2603
rect 5266 2603 5272 2604
rect 4979 2600 5089 2602
rect 4979 2599 4980 2600
rect 4974 2598 4980 2599
rect 5266 2599 5267 2603
rect 5271 2602 5272 2603
rect 5271 2600 5377 2602
rect 5271 2599 5272 2600
rect 5266 2598 5272 2599
rect 3110 2594 3116 2595
rect 695 2591 701 2592
rect 695 2587 696 2591
rect 700 2590 701 2591
rect 738 2591 744 2592
rect 738 2590 739 2591
rect 700 2588 739 2590
rect 700 2587 701 2588
rect 695 2586 701 2587
rect 738 2587 739 2588
rect 743 2587 744 2591
rect 738 2586 744 2587
rect 855 2591 861 2592
rect 855 2587 856 2591
rect 860 2590 861 2591
rect 898 2591 904 2592
rect 898 2590 899 2591
rect 860 2588 899 2590
rect 860 2587 861 2588
rect 855 2586 861 2587
rect 898 2587 899 2588
rect 903 2587 904 2591
rect 898 2586 904 2587
rect 1015 2591 1024 2592
rect 1015 2587 1016 2591
rect 1023 2587 1024 2591
rect 1015 2586 1024 2587
rect 1090 2591 1096 2592
rect 1090 2587 1091 2591
rect 1095 2590 1096 2591
rect 1167 2591 1173 2592
rect 1167 2590 1168 2591
rect 1095 2588 1168 2590
rect 1095 2587 1096 2588
rect 1090 2586 1096 2587
rect 1167 2587 1168 2588
rect 1172 2587 1173 2591
rect 1167 2586 1173 2587
rect 1186 2591 1192 2592
rect 1186 2587 1187 2591
rect 1191 2590 1192 2591
rect 1319 2591 1325 2592
rect 1319 2590 1320 2591
rect 1191 2588 1320 2590
rect 1191 2587 1192 2588
rect 1186 2586 1192 2587
rect 1319 2587 1320 2588
rect 1324 2587 1325 2591
rect 1319 2586 1325 2587
rect 1351 2591 1357 2592
rect 1351 2587 1352 2591
rect 1356 2590 1357 2591
rect 1479 2591 1485 2592
rect 1479 2590 1480 2591
rect 1356 2588 1480 2590
rect 1356 2587 1357 2588
rect 1351 2586 1357 2587
rect 1479 2587 1480 2588
rect 1484 2587 1485 2591
rect 1479 2586 1485 2587
rect 1498 2591 1504 2592
rect 1498 2587 1499 2591
rect 1503 2590 1504 2591
rect 1639 2591 1645 2592
rect 1639 2590 1640 2591
rect 1503 2588 1640 2590
rect 1503 2587 1504 2588
rect 1498 2586 1504 2587
rect 1639 2587 1640 2588
rect 1644 2587 1645 2591
rect 1639 2586 1645 2587
rect 1671 2591 1677 2592
rect 1671 2587 1672 2591
rect 1676 2590 1677 2591
rect 1799 2591 1805 2592
rect 1799 2590 1800 2591
rect 1676 2588 1800 2590
rect 1676 2587 1677 2588
rect 1671 2586 1677 2587
rect 1799 2587 1800 2588
rect 1804 2587 1805 2591
rect 1799 2586 1805 2587
rect 110 2584 116 2585
rect 1934 2584 1940 2585
rect 110 2580 111 2584
rect 115 2580 116 2584
rect 110 2579 116 2580
rect 570 2583 576 2584
rect 570 2579 571 2583
rect 575 2579 576 2583
rect 570 2578 576 2579
rect 730 2583 736 2584
rect 730 2579 731 2583
rect 735 2579 736 2583
rect 730 2578 736 2579
rect 890 2583 896 2584
rect 890 2579 891 2583
rect 895 2579 896 2583
rect 890 2578 896 2579
rect 1042 2583 1048 2584
rect 1042 2579 1043 2583
rect 1047 2579 1048 2583
rect 1042 2578 1048 2579
rect 1194 2583 1200 2584
rect 1194 2579 1195 2583
rect 1199 2579 1200 2583
rect 1194 2578 1200 2579
rect 1354 2583 1360 2584
rect 1354 2579 1355 2583
rect 1359 2579 1360 2583
rect 1354 2578 1360 2579
rect 1514 2583 1520 2584
rect 1514 2579 1515 2583
rect 1519 2579 1520 2583
rect 1514 2578 1520 2579
rect 1674 2583 1680 2584
rect 1674 2579 1675 2583
rect 1679 2579 1680 2583
rect 1934 2580 1935 2584
rect 1939 2580 1940 2584
rect 1934 2579 1940 2580
rect 1674 2578 1680 2579
rect 4079 2571 4085 2572
rect 4079 2570 4080 2571
rect 598 2568 604 2569
rect 110 2567 116 2568
rect 110 2563 111 2567
rect 115 2563 116 2567
rect 598 2564 599 2568
rect 603 2564 604 2568
rect 598 2563 604 2564
rect 758 2568 764 2569
rect 758 2564 759 2568
rect 763 2564 764 2568
rect 758 2563 764 2564
rect 918 2568 924 2569
rect 918 2564 919 2568
rect 923 2564 924 2568
rect 918 2563 924 2564
rect 1070 2568 1076 2569
rect 1070 2564 1071 2568
rect 1075 2564 1076 2568
rect 1070 2563 1076 2564
rect 1222 2568 1228 2569
rect 1222 2564 1223 2568
rect 1227 2564 1228 2568
rect 1222 2563 1228 2564
rect 1382 2568 1388 2569
rect 1382 2564 1383 2568
rect 1387 2564 1388 2568
rect 1382 2563 1388 2564
rect 1542 2568 1548 2569
rect 1542 2564 1543 2568
rect 1547 2564 1548 2568
rect 1542 2563 1548 2564
rect 1702 2568 1708 2569
rect 3957 2568 4080 2570
rect 1702 2564 1703 2568
rect 1707 2564 1708 2568
rect 1702 2563 1708 2564
rect 1934 2567 1940 2568
rect 1934 2563 1935 2567
rect 1939 2563 1940 2567
rect 4079 2567 4080 2568
rect 4084 2567 4085 2571
rect 4575 2571 4581 2572
rect 4575 2570 4576 2571
rect 4429 2568 4576 2570
rect 4079 2566 4085 2567
rect 4178 2567 4184 2568
rect 110 2562 116 2563
rect 1934 2562 1940 2563
rect 4178 2563 4179 2567
rect 4183 2563 4184 2567
rect 4575 2567 4576 2568
rect 4580 2567 4581 2571
rect 4575 2566 4581 2567
rect 4638 2571 4644 2572
rect 4638 2567 4639 2571
rect 4643 2567 4644 2571
rect 5071 2571 5077 2572
rect 5071 2570 5072 2571
rect 4925 2568 5072 2570
rect 4638 2566 4644 2567
rect 5071 2567 5072 2568
rect 5076 2567 5077 2571
rect 5418 2571 5424 2572
rect 5071 2566 5077 2567
rect 5170 2567 5176 2568
rect 4178 2562 4184 2563
rect 5170 2563 5171 2567
rect 5175 2563 5176 2567
rect 5418 2567 5419 2571
rect 5423 2567 5424 2571
rect 5418 2566 5424 2567
rect 5170 2562 5176 2563
rect 2538 2555 2544 2556
rect 2538 2551 2539 2555
rect 2543 2554 2544 2555
rect 2679 2555 2685 2556
rect 2679 2554 2680 2555
rect 2543 2552 2680 2554
rect 2543 2551 2544 2552
rect 2538 2550 2544 2551
rect 2679 2551 2680 2552
rect 2684 2551 2685 2555
rect 2679 2550 2685 2551
rect 2687 2555 2693 2556
rect 2687 2551 2688 2555
rect 2692 2554 2693 2555
rect 2815 2555 2821 2556
rect 2815 2554 2816 2555
rect 2692 2552 2816 2554
rect 2692 2551 2693 2552
rect 2687 2550 2693 2551
rect 2815 2551 2816 2552
rect 2820 2551 2821 2555
rect 2815 2550 2821 2551
rect 2950 2555 2957 2556
rect 2950 2551 2951 2555
rect 2956 2551 2957 2555
rect 2950 2550 2957 2551
rect 2959 2555 2965 2556
rect 2959 2551 2960 2555
rect 2964 2554 2965 2555
rect 3087 2555 3093 2556
rect 3087 2554 3088 2555
rect 2964 2552 3088 2554
rect 2964 2551 2965 2552
rect 2959 2550 2965 2551
rect 3087 2551 3088 2552
rect 3092 2551 3093 2555
rect 3087 2550 3093 2551
rect 3095 2555 3101 2556
rect 3095 2551 3096 2555
rect 3100 2554 3101 2555
rect 3223 2555 3229 2556
rect 3223 2554 3224 2555
rect 3100 2552 3224 2554
rect 3100 2551 3101 2552
rect 3095 2550 3101 2551
rect 3223 2551 3224 2552
rect 3228 2551 3229 2555
rect 3223 2550 3229 2551
rect 1974 2548 1980 2549
rect 3798 2548 3804 2549
rect 1974 2544 1975 2548
rect 1979 2544 1980 2548
rect 1974 2543 1980 2544
rect 2554 2547 2560 2548
rect 2554 2543 2555 2547
rect 2559 2543 2560 2547
rect 2554 2542 2560 2543
rect 2690 2547 2696 2548
rect 2690 2543 2691 2547
rect 2695 2543 2696 2547
rect 2690 2542 2696 2543
rect 2826 2547 2832 2548
rect 2826 2543 2827 2547
rect 2831 2543 2832 2547
rect 2826 2542 2832 2543
rect 2962 2547 2968 2548
rect 2962 2543 2963 2547
rect 2967 2543 2968 2547
rect 2962 2542 2968 2543
rect 3098 2547 3104 2548
rect 3098 2543 3099 2547
rect 3103 2543 3104 2547
rect 3798 2544 3799 2548
rect 3803 2544 3804 2548
rect 3798 2543 3804 2544
rect 3098 2542 3104 2543
rect 2582 2532 2588 2533
rect 1974 2531 1980 2532
rect 1974 2527 1975 2531
rect 1979 2527 1980 2531
rect 2582 2528 2583 2532
rect 2587 2528 2588 2532
rect 2582 2527 2588 2528
rect 2718 2532 2724 2533
rect 2718 2528 2719 2532
rect 2723 2528 2724 2532
rect 2718 2527 2724 2528
rect 2854 2532 2860 2533
rect 2854 2528 2855 2532
rect 2859 2528 2860 2532
rect 2854 2527 2860 2528
rect 2990 2532 2996 2533
rect 2990 2528 2991 2532
rect 2995 2528 2996 2532
rect 2990 2527 2996 2528
rect 3126 2532 3132 2533
rect 3126 2528 3127 2532
rect 3131 2528 3132 2532
rect 3126 2527 3132 2528
rect 3798 2531 3804 2532
rect 3798 2527 3799 2531
rect 3803 2527 3804 2531
rect 1974 2526 1980 2527
rect 3798 2526 3804 2527
rect 3982 2527 3989 2528
rect 3982 2523 3983 2527
rect 3988 2523 3989 2527
rect 3982 2522 3989 2523
rect 4079 2527 4085 2528
rect 4079 2523 4080 2527
rect 4084 2526 4085 2527
rect 4207 2527 4213 2528
rect 4207 2526 4208 2527
rect 4084 2524 4208 2526
rect 4084 2523 4085 2524
rect 4079 2522 4085 2523
rect 4207 2523 4208 2524
rect 4212 2523 4213 2527
rect 4207 2522 4213 2523
rect 4394 2527 4400 2528
rect 4394 2523 4395 2527
rect 4399 2526 4400 2527
rect 4455 2527 4461 2528
rect 4455 2526 4456 2527
rect 4399 2524 4456 2526
rect 4399 2523 4400 2524
rect 4394 2522 4400 2523
rect 4455 2523 4456 2524
rect 4460 2523 4461 2527
rect 4455 2522 4461 2523
rect 4575 2527 4581 2528
rect 4575 2523 4576 2527
rect 4580 2526 4581 2527
rect 4703 2527 4709 2528
rect 4703 2526 4704 2527
rect 4580 2524 4704 2526
rect 4580 2523 4581 2524
rect 4575 2522 4581 2523
rect 4703 2523 4704 2524
rect 4708 2523 4709 2527
rect 4703 2522 4709 2523
rect 4890 2527 4896 2528
rect 4890 2523 4891 2527
rect 4895 2526 4896 2527
rect 4951 2527 4957 2528
rect 4951 2526 4952 2527
rect 4895 2524 4952 2526
rect 4895 2523 4896 2524
rect 4890 2522 4896 2523
rect 4951 2523 4952 2524
rect 4956 2523 4957 2527
rect 4951 2522 4957 2523
rect 5071 2527 5077 2528
rect 5071 2523 5072 2527
rect 5076 2526 5077 2527
rect 5199 2527 5205 2528
rect 5199 2526 5200 2527
rect 5076 2524 5200 2526
rect 5076 2523 5077 2524
rect 5071 2522 5077 2523
rect 5199 2523 5200 2524
rect 5204 2523 5205 2527
rect 5199 2522 5205 2523
rect 5446 2527 5453 2528
rect 5446 2523 5447 2527
rect 5452 2523 5453 2527
rect 5446 2522 5453 2523
rect 3838 2520 3844 2521
rect 5662 2520 5668 2521
rect 3838 2516 3839 2520
rect 3843 2516 3844 2520
rect 3838 2515 3844 2516
rect 3858 2519 3864 2520
rect 3858 2515 3859 2519
rect 3863 2515 3864 2519
rect 3858 2514 3864 2515
rect 4082 2519 4088 2520
rect 4082 2515 4083 2519
rect 4087 2515 4088 2519
rect 4082 2514 4088 2515
rect 4330 2519 4336 2520
rect 4330 2515 4331 2519
rect 4335 2515 4336 2519
rect 4330 2514 4336 2515
rect 4578 2519 4584 2520
rect 4578 2515 4579 2519
rect 4583 2515 4584 2519
rect 4578 2514 4584 2515
rect 4826 2519 4832 2520
rect 4826 2515 4827 2519
rect 4831 2515 4832 2519
rect 4826 2514 4832 2515
rect 5074 2519 5080 2520
rect 5074 2515 5075 2519
rect 5079 2515 5080 2519
rect 5074 2514 5080 2515
rect 5322 2519 5328 2520
rect 5322 2515 5323 2519
rect 5327 2515 5328 2519
rect 5662 2516 5663 2520
rect 5667 2516 5668 2520
rect 5662 2515 5668 2516
rect 5322 2514 5328 2515
rect 110 2509 116 2510
rect 1934 2509 1940 2510
rect 110 2505 111 2509
rect 115 2505 116 2509
rect 110 2504 116 2505
rect 382 2508 388 2509
rect 382 2504 383 2508
rect 387 2504 388 2508
rect 382 2503 388 2504
rect 598 2508 604 2509
rect 598 2504 599 2508
rect 603 2504 604 2508
rect 598 2503 604 2504
rect 814 2508 820 2509
rect 814 2504 815 2508
rect 819 2504 820 2508
rect 814 2503 820 2504
rect 1022 2508 1028 2509
rect 1022 2504 1023 2508
rect 1027 2504 1028 2508
rect 1022 2503 1028 2504
rect 1230 2508 1236 2509
rect 1230 2504 1231 2508
rect 1235 2504 1236 2508
rect 1230 2503 1236 2504
rect 1430 2508 1436 2509
rect 1430 2504 1431 2508
rect 1435 2504 1436 2508
rect 1430 2503 1436 2504
rect 1630 2508 1636 2509
rect 1630 2504 1631 2508
rect 1635 2504 1636 2508
rect 1630 2503 1636 2504
rect 1814 2508 1820 2509
rect 1814 2504 1815 2508
rect 1819 2504 1820 2508
rect 1934 2505 1935 2509
rect 1939 2505 1940 2509
rect 1934 2504 1940 2505
rect 3886 2504 3892 2505
rect 1814 2503 1820 2504
rect 3838 2503 3844 2504
rect 3838 2499 3839 2503
rect 3843 2499 3844 2503
rect 3886 2500 3887 2504
rect 3891 2500 3892 2504
rect 3886 2499 3892 2500
rect 4110 2504 4116 2505
rect 4110 2500 4111 2504
rect 4115 2500 4116 2504
rect 4110 2499 4116 2500
rect 4358 2504 4364 2505
rect 4358 2500 4359 2504
rect 4363 2500 4364 2504
rect 4358 2499 4364 2500
rect 4606 2504 4612 2505
rect 4606 2500 4607 2504
rect 4611 2500 4612 2504
rect 4606 2499 4612 2500
rect 4854 2504 4860 2505
rect 4854 2500 4855 2504
rect 4859 2500 4860 2504
rect 4854 2499 4860 2500
rect 5102 2504 5108 2505
rect 5102 2500 5103 2504
rect 5107 2500 5108 2504
rect 5102 2499 5108 2500
rect 5350 2504 5356 2505
rect 5350 2500 5351 2504
rect 5355 2500 5356 2504
rect 5350 2499 5356 2500
rect 5662 2503 5668 2504
rect 5662 2499 5663 2503
rect 5667 2499 5668 2503
rect 3838 2498 3844 2499
rect 5662 2498 5668 2499
rect 354 2493 360 2494
rect 110 2492 116 2493
rect 110 2488 111 2492
rect 115 2488 116 2492
rect 354 2489 355 2493
rect 359 2489 360 2493
rect 354 2488 360 2489
rect 570 2493 576 2494
rect 570 2489 571 2493
rect 575 2489 576 2493
rect 570 2488 576 2489
rect 786 2493 792 2494
rect 786 2489 787 2493
rect 791 2489 792 2493
rect 786 2488 792 2489
rect 994 2493 1000 2494
rect 994 2489 995 2493
rect 999 2489 1000 2493
rect 994 2488 1000 2489
rect 1202 2493 1208 2494
rect 1202 2489 1203 2493
rect 1207 2489 1208 2493
rect 1202 2488 1208 2489
rect 1402 2493 1408 2494
rect 1402 2489 1403 2493
rect 1407 2489 1408 2493
rect 1402 2488 1408 2489
rect 1602 2493 1608 2494
rect 1602 2489 1603 2493
rect 1607 2489 1608 2493
rect 1602 2488 1608 2489
rect 1786 2493 1792 2494
rect 1786 2489 1787 2493
rect 1791 2489 1792 2493
rect 1786 2488 1792 2489
rect 1934 2492 1940 2493
rect 1934 2488 1935 2492
rect 1939 2488 1940 2492
rect 110 2487 116 2488
rect 1934 2487 1940 2488
rect 479 2483 485 2484
rect 479 2479 480 2483
rect 484 2482 485 2483
rect 511 2483 517 2484
rect 511 2482 512 2483
rect 484 2480 512 2482
rect 484 2479 485 2480
rect 479 2478 485 2479
rect 511 2479 512 2480
rect 516 2479 517 2483
rect 511 2478 517 2479
rect 695 2483 701 2484
rect 695 2479 696 2483
rect 700 2482 701 2483
rect 727 2483 733 2484
rect 727 2482 728 2483
rect 700 2480 728 2482
rect 700 2479 701 2480
rect 695 2478 701 2479
rect 727 2479 728 2480
rect 732 2479 733 2483
rect 727 2478 733 2479
rect 882 2483 888 2484
rect 882 2479 883 2483
rect 887 2482 888 2483
rect 911 2483 917 2484
rect 911 2482 912 2483
rect 887 2480 912 2482
rect 887 2479 888 2480
rect 882 2478 888 2479
rect 911 2479 912 2480
rect 916 2479 917 2483
rect 911 2478 917 2479
rect 1119 2483 1125 2484
rect 1119 2479 1120 2483
rect 1124 2482 1125 2483
rect 1166 2483 1172 2484
rect 1166 2482 1167 2483
rect 1124 2480 1167 2482
rect 1124 2479 1125 2480
rect 1119 2478 1125 2479
rect 1166 2479 1167 2480
rect 1171 2479 1172 2483
rect 1166 2478 1172 2479
rect 1327 2483 1333 2484
rect 1327 2479 1328 2483
rect 1332 2482 1333 2483
rect 1399 2483 1405 2484
rect 1399 2482 1400 2483
rect 1332 2480 1400 2482
rect 1332 2479 1333 2480
rect 1327 2478 1333 2479
rect 1399 2479 1400 2480
rect 1404 2479 1405 2483
rect 1399 2478 1405 2479
rect 1527 2483 1533 2484
rect 1527 2479 1528 2483
rect 1532 2482 1533 2483
rect 1562 2483 1568 2484
rect 1562 2482 1563 2483
rect 1532 2480 1563 2482
rect 1532 2479 1533 2480
rect 1527 2478 1533 2479
rect 1562 2479 1563 2480
rect 1567 2479 1568 2483
rect 1562 2478 1568 2479
rect 1727 2483 1736 2484
rect 1727 2479 1728 2483
rect 1735 2479 1736 2483
rect 1727 2478 1736 2479
rect 1882 2483 1888 2484
rect 1882 2479 1883 2483
rect 1887 2482 1888 2483
rect 1911 2483 1917 2484
rect 1911 2482 1912 2483
rect 1887 2480 1912 2482
rect 1887 2479 1888 2480
rect 1882 2478 1888 2479
rect 1911 2479 1912 2480
rect 1916 2479 1917 2483
rect 1911 2478 1917 2479
rect 1974 2449 1980 2450
rect 3798 2449 3804 2450
rect 1974 2445 1975 2449
rect 1979 2445 1980 2449
rect 1974 2444 1980 2445
rect 2022 2448 2028 2449
rect 2022 2444 2023 2448
rect 2027 2444 2028 2448
rect 362 2443 368 2444
rect 362 2439 363 2443
rect 367 2439 368 2443
rect 362 2438 368 2439
rect 511 2443 517 2444
rect 511 2439 512 2443
rect 516 2442 517 2443
rect 727 2443 733 2444
rect 516 2440 577 2442
rect 516 2439 517 2440
rect 511 2438 517 2439
rect 727 2439 728 2443
rect 732 2442 733 2443
rect 1090 2443 1096 2444
rect 732 2440 793 2442
rect 732 2439 733 2440
rect 727 2438 733 2439
rect 1090 2439 1091 2443
rect 1095 2439 1096 2443
rect 1090 2438 1096 2439
rect 1166 2443 1172 2444
rect 1166 2439 1167 2443
rect 1171 2442 1172 2443
rect 1498 2443 1504 2444
rect 1171 2440 1209 2442
rect 1171 2439 1172 2440
rect 1166 2438 1172 2439
rect 1498 2439 1499 2443
rect 1503 2439 1504 2443
rect 1498 2438 1504 2439
rect 1562 2443 1568 2444
rect 1562 2439 1563 2443
rect 1567 2442 1568 2443
rect 1730 2443 1736 2444
rect 2022 2443 2028 2444
rect 2222 2448 2228 2449
rect 2222 2444 2223 2448
rect 2227 2444 2228 2448
rect 2222 2443 2228 2444
rect 2446 2448 2452 2449
rect 2446 2444 2447 2448
rect 2451 2444 2452 2448
rect 2446 2443 2452 2444
rect 2678 2448 2684 2449
rect 2678 2444 2679 2448
rect 2683 2444 2684 2448
rect 2678 2443 2684 2444
rect 2926 2448 2932 2449
rect 2926 2444 2927 2448
rect 2931 2444 2932 2448
rect 2926 2443 2932 2444
rect 3182 2448 3188 2449
rect 3182 2444 3183 2448
rect 3187 2444 3188 2448
rect 3182 2443 3188 2444
rect 3438 2448 3444 2449
rect 3438 2444 3439 2448
rect 3443 2444 3444 2448
rect 3438 2443 3444 2444
rect 3678 2448 3684 2449
rect 3678 2444 3679 2448
rect 3683 2444 3684 2448
rect 3798 2445 3799 2449
rect 3803 2445 3804 2449
rect 3798 2444 3804 2445
rect 3678 2443 3684 2444
rect 1567 2440 1609 2442
rect 1567 2439 1568 2440
rect 1562 2438 1568 2439
rect 1730 2439 1731 2443
rect 1735 2442 1736 2443
rect 1735 2440 1793 2442
rect 3838 2441 3844 2442
rect 5662 2441 5668 2442
rect 1735 2439 1736 2440
rect 1730 2438 1736 2439
rect 3838 2437 3839 2441
rect 3843 2437 3844 2441
rect 3838 2436 3844 2437
rect 3886 2440 3892 2441
rect 3886 2436 3887 2440
rect 3891 2436 3892 2440
rect 3886 2435 3892 2436
rect 4086 2440 4092 2441
rect 4086 2436 4087 2440
rect 4091 2436 4092 2440
rect 4086 2435 4092 2436
rect 4326 2440 4332 2441
rect 4326 2436 4327 2440
rect 4331 2436 4332 2440
rect 4326 2435 4332 2436
rect 4582 2440 4588 2441
rect 4582 2436 4583 2440
rect 4587 2436 4588 2440
rect 4582 2435 4588 2436
rect 4846 2440 4852 2441
rect 4846 2436 4847 2440
rect 4851 2436 4852 2440
rect 4846 2435 4852 2436
rect 5118 2440 5124 2441
rect 5118 2436 5119 2440
rect 5123 2436 5124 2440
rect 5118 2435 5124 2436
rect 5398 2440 5404 2441
rect 5398 2436 5399 2440
rect 5403 2436 5404 2440
rect 5662 2437 5663 2441
rect 5667 2437 5668 2441
rect 5662 2436 5668 2437
rect 5398 2435 5404 2436
rect 1994 2433 2000 2434
rect 1974 2432 1980 2433
rect 1974 2428 1975 2432
rect 1979 2428 1980 2432
rect 1994 2429 1995 2433
rect 1999 2429 2000 2433
rect 1994 2428 2000 2429
rect 2194 2433 2200 2434
rect 2194 2429 2195 2433
rect 2199 2429 2200 2433
rect 2194 2428 2200 2429
rect 2418 2433 2424 2434
rect 2418 2429 2419 2433
rect 2423 2429 2424 2433
rect 2418 2428 2424 2429
rect 2650 2433 2656 2434
rect 2650 2429 2651 2433
rect 2655 2429 2656 2433
rect 2650 2428 2656 2429
rect 2898 2433 2904 2434
rect 2898 2429 2899 2433
rect 2903 2429 2904 2433
rect 2898 2428 2904 2429
rect 3154 2433 3160 2434
rect 3154 2429 3155 2433
rect 3159 2429 3160 2433
rect 3154 2428 3160 2429
rect 3410 2433 3416 2434
rect 3410 2429 3411 2433
rect 3415 2429 3416 2433
rect 3410 2428 3416 2429
rect 3650 2433 3656 2434
rect 3650 2429 3651 2433
rect 3655 2429 3656 2433
rect 3650 2428 3656 2429
rect 3798 2432 3804 2433
rect 3798 2428 3799 2432
rect 3803 2428 3804 2432
rect 1974 2427 1980 2428
rect 3798 2427 3804 2428
rect 3858 2425 3864 2426
rect 3838 2424 3844 2425
rect 2090 2423 2096 2424
rect 2090 2419 2091 2423
rect 2095 2422 2096 2423
rect 2119 2423 2125 2424
rect 2119 2422 2120 2423
rect 2095 2420 2120 2422
rect 2095 2419 2096 2420
rect 2090 2418 2096 2419
rect 2119 2419 2120 2420
rect 2124 2419 2125 2423
rect 2119 2418 2125 2419
rect 2319 2423 2328 2424
rect 2319 2419 2320 2423
rect 2327 2419 2328 2423
rect 2319 2418 2328 2419
rect 2543 2423 2552 2424
rect 2543 2419 2544 2423
rect 2551 2419 2552 2423
rect 2543 2418 2552 2419
rect 2774 2423 2781 2424
rect 2774 2419 2775 2423
rect 2780 2419 2781 2423
rect 2774 2418 2781 2419
rect 3023 2423 3032 2424
rect 3023 2419 3024 2423
rect 3031 2419 3032 2423
rect 3023 2418 3032 2419
rect 3279 2423 3288 2424
rect 3279 2419 3280 2423
rect 3287 2419 3288 2423
rect 3279 2418 3288 2419
rect 3534 2423 3541 2424
rect 3534 2419 3535 2423
rect 3540 2419 3541 2423
rect 3534 2418 3541 2419
rect 3775 2423 3781 2424
rect 3775 2419 3776 2423
rect 3780 2422 3781 2423
rect 3822 2423 3828 2424
rect 3822 2422 3823 2423
rect 3780 2420 3823 2422
rect 3780 2419 3781 2420
rect 3775 2418 3781 2419
rect 3822 2419 3823 2420
rect 3827 2419 3828 2423
rect 3838 2420 3839 2424
rect 3843 2420 3844 2424
rect 3858 2421 3859 2425
rect 3863 2421 3864 2425
rect 3858 2420 3864 2421
rect 4058 2425 4064 2426
rect 4058 2421 4059 2425
rect 4063 2421 4064 2425
rect 4058 2420 4064 2421
rect 4298 2425 4304 2426
rect 4298 2421 4299 2425
rect 4303 2421 4304 2425
rect 4298 2420 4304 2421
rect 4554 2425 4560 2426
rect 4554 2421 4555 2425
rect 4559 2421 4560 2425
rect 4554 2420 4560 2421
rect 4818 2425 4824 2426
rect 4818 2421 4819 2425
rect 4823 2421 4824 2425
rect 4818 2420 4824 2421
rect 5090 2425 5096 2426
rect 5090 2421 5091 2425
rect 5095 2421 5096 2425
rect 5090 2420 5096 2421
rect 5370 2425 5376 2426
rect 5370 2421 5371 2425
rect 5375 2421 5376 2425
rect 5370 2420 5376 2421
rect 5662 2424 5668 2425
rect 5662 2420 5663 2424
rect 5667 2420 5668 2424
rect 3838 2419 3844 2420
rect 5662 2419 5668 2420
rect 3822 2418 3828 2419
rect 1278 2415 1284 2416
rect 1278 2414 1279 2415
rect 1099 2412 1279 2414
rect 454 2407 460 2408
rect 454 2406 455 2407
rect 325 2404 455 2406
rect 454 2403 455 2404
rect 459 2403 460 2407
rect 1099 2406 1101 2412
rect 1278 2411 1279 2412
rect 1283 2411 1284 2415
rect 1594 2415 1600 2416
rect 1594 2414 1595 2415
rect 1278 2410 1284 2411
rect 1384 2412 1595 2414
rect 1384 2406 1386 2412
rect 1594 2411 1595 2412
rect 1599 2411 1600 2415
rect 1594 2410 1600 2411
rect 3983 2415 3989 2416
rect 3983 2411 3984 2415
rect 3988 2414 3989 2415
rect 4022 2415 4028 2416
rect 4022 2414 4023 2415
rect 3988 2412 4023 2414
rect 3988 2411 3989 2412
rect 3983 2410 3989 2411
rect 4022 2411 4023 2412
rect 4027 2411 4028 2415
rect 4022 2410 4028 2411
rect 4178 2415 4189 2416
rect 4178 2411 4179 2415
rect 4183 2411 4184 2415
rect 4188 2411 4189 2415
rect 4178 2410 4189 2411
rect 4423 2415 4429 2416
rect 4423 2411 4424 2415
rect 4428 2414 4429 2415
rect 4439 2415 4445 2416
rect 4439 2414 4440 2415
rect 4428 2412 4440 2414
rect 4428 2411 4429 2412
rect 4423 2410 4429 2411
rect 4439 2411 4440 2412
rect 4444 2411 4445 2415
rect 4439 2410 4445 2411
rect 4679 2415 4688 2416
rect 4679 2411 4680 2415
rect 4687 2411 4688 2415
rect 4679 2410 4688 2411
rect 4890 2415 4896 2416
rect 4890 2411 4891 2415
rect 4895 2414 4896 2415
rect 4943 2415 4949 2416
rect 4943 2414 4944 2415
rect 4895 2412 4944 2414
rect 4895 2411 4896 2412
rect 4890 2410 4896 2411
rect 4943 2411 4944 2412
rect 4948 2411 4949 2415
rect 4943 2410 4949 2411
rect 5170 2415 5176 2416
rect 5170 2411 5171 2415
rect 5175 2414 5176 2415
rect 5215 2415 5221 2416
rect 5215 2414 5216 2415
rect 5175 2412 5216 2414
rect 5175 2411 5176 2412
rect 5170 2410 5176 2411
rect 5215 2411 5216 2412
rect 5220 2411 5221 2415
rect 5215 2410 5221 2411
rect 5434 2415 5440 2416
rect 5434 2411 5435 2415
rect 5439 2414 5440 2415
rect 5495 2415 5501 2416
rect 5495 2414 5496 2415
rect 5439 2412 5496 2414
rect 5439 2411 5440 2412
rect 5434 2410 5440 2411
rect 5495 2411 5496 2412
rect 5500 2411 5501 2415
rect 5495 2410 5501 2411
rect 933 2404 1101 2406
rect 1253 2404 1386 2406
rect 1399 2407 1405 2408
rect 454 2402 460 2403
rect 618 2403 624 2404
rect 618 2399 619 2403
rect 623 2399 624 2403
rect 1399 2403 1400 2407
rect 1404 2406 1405 2407
rect 1882 2407 1888 2408
rect 1404 2404 1489 2406
rect 1404 2403 1405 2404
rect 1399 2402 1405 2403
rect 1882 2403 1883 2407
rect 1887 2403 1888 2407
rect 1882 2402 1888 2403
rect 618 2398 624 2399
rect 2322 2383 2328 2384
rect 2292 2374 2294 2381
rect 2322 2379 2323 2383
rect 2327 2382 2328 2383
rect 2546 2383 2552 2384
rect 2327 2380 2425 2382
rect 2327 2379 2328 2380
rect 2322 2378 2328 2379
rect 2546 2379 2547 2383
rect 2551 2382 2552 2383
rect 2950 2383 2956 2384
rect 2551 2380 2657 2382
rect 2551 2379 2552 2380
rect 2546 2378 2552 2379
rect 2950 2379 2951 2383
rect 2955 2379 2956 2383
rect 2950 2378 2956 2379
rect 3026 2383 3032 2384
rect 3026 2379 3027 2383
rect 3031 2382 3032 2383
rect 3282 2383 3288 2384
rect 3031 2380 3161 2382
rect 3031 2379 3032 2380
rect 3026 2378 3032 2379
rect 3282 2379 3283 2383
rect 3287 2382 3288 2383
rect 3746 2383 3752 2384
rect 3287 2380 3417 2382
rect 3287 2379 3288 2380
rect 3282 2378 3288 2379
rect 3746 2379 3747 2383
rect 3751 2379 3752 2383
rect 3746 2378 3752 2379
rect 2546 2375 2552 2376
rect 2546 2374 2547 2375
rect 2292 2372 2547 2374
rect 1999 2371 2005 2372
rect 1999 2370 2000 2371
rect 1939 2368 2000 2370
rect 351 2363 357 2364
rect 351 2359 352 2363
rect 356 2362 357 2363
rect 362 2363 368 2364
rect 362 2362 363 2363
rect 356 2360 363 2362
rect 356 2359 357 2360
rect 351 2358 357 2359
rect 362 2359 363 2360
rect 367 2359 368 2363
rect 362 2358 368 2359
rect 454 2363 460 2364
rect 454 2359 455 2363
rect 459 2362 460 2363
rect 647 2363 653 2364
rect 647 2362 648 2363
rect 459 2360 648 2362
rect 459 2359 460 2360
rect 454 2358 460 2359
rect 647 2359 648 2360
rect 652 2359 653 2363
rect 647 2358 653 2359
rect 898 2363 904 2364
rect 898 2359 899 2363
rect 903 2362 904 2363
rect 959 2363 965 2364
rect 959 2362 960 2363
rect 903 2360 960 2362
rect 903 2359 904 2360
rect 898 2358 904 2359
rect 959 2359 960 2360
rect 964 2359 965 2363
rect 959 2358 965 2359
rect 1278 2363 1285 2364
rect 1278 2359 1279 2363
rect 1284 2359 1285 2363
rect 1278 2358 1285 2359
rect 1594 2363 1600 2364
rect 1594 2359 1595 2363
rect 1599 2362 1600 2363
rect 1607 2363 1613 2364
rect 1607 2362 1608 2363
rect 1599 2360 1608 2362
rect 1599 2359 1600 2360
rect 1594 2358 1600 2359
rect 1607 2359 1608 2360
rect 1612 2359 1613 2363
rect 1607 2358 1613 2359
rect 1911 2363 1917 2364
rect 1911 2359 1912 2363
rect 1916 2362 1917 2363
rect 1939 2362 1941 2368
rect 1999 2367 2000 2368
rect 2004 2367 2005 2371
rect 2546 2371 2547 2372
rect 2551 2371 2552 2375
rect 2546 2370 2552 2371
rect 3822 2375 3828 2376
rect 3822 2371 3823 2375
rect 3827 2374 3828 2375
rect 4022 2375 4028 2376
rect 3827 2372 3865 2374
rect 3827 2371 3828 2372
rect 3822 2370 3828 2371
rect 4022 2371 4023 2375
rect 4027 2374 4028 2375
rect 4394 2375 4400 2376
rect 4027 2372 4065 2374
rect 4027 2371 4028 2372
rect 4022 2370 4028 2371
rect 4394 2371 4395 2375
rect 4399 2371 4400 2375
rect 4394 2370 4400 2371
rect 4439 2375 4445 2376
rect 4439 2371 4440 2375
rect 4444 2374 4445 2375
rect 4682 2375 4688 2376
rect 4444 2372 4561 2374
rect 4444 2371 4445 2372
rect 4439 2370 4445 2371
rect 4682 2371 4683 2375
rect 4687 2374 4688 2375
rect 5098 2375 5104 2376
rect 4687 2372 4825 2374
rect 4687 2371 4688 2372
rect 4682 2370 4688 2371
rect 5098 2371 5099 2375
rect 5103 2371 5104 2375
rect 5098 2370 5104 2371
rect 5446 2375 5452 2376
rect 5446 2371 5447 2375
rect 5451 2371 5452 2375
rect 5446 2370 5452 2371
rect 1999 2366 2005 2367
rect 1916 2360 1941 2362
rect 1916 2359 1917 2360
rect 1911 2358 1917 2359
rect 110 2356 116 2357
rect 1934 2356 1940 2357
rect 110 2352 111 2356
rect 115 2352 116 2356
rect 110 2351 116 2352
rect 226 2355 232 2356
rect 226 2351 227 2355
rect 231 2351 232 2355
rect 226 2350 232 2351
rect 522 2355 528 2356
rect 522 2351 523 2355
rect 527 2351 528 2355
rect 522 2350 528 2351
rect 834 2355 840 2356
rect 834 2351 835 2355
rect 839 2351 840 2355
rect 834 2350 840 2351
rect 1154 2355 1160 2356
rect 1154 2351 1155 2355
rect 1159 2351 1160 2355
rect 1154 2350 1160 2351
rect 1482 2355 1488 2356
rect 1482 2351 1483 2355
rect 1487 2351 1488 2355
rect 1482 2350 1488 2351
rect 1786 2355 1792 2356
rect 1786 2351 1787 2355
rect 1791 2351 1792 2355
rect 1934 2352 1935 2356
rect 1939 2352 1940 2356
rect 1934 2351 1940 2352
rect 1786 2350 1792 2351
rect 2090 2343 2096 2344
rect 254 2340 260 2341
rect 110 2339 116 2340
rect 110 2335 111 2339
rect 115 2335 116 2339
rect 254 2336 255 2340
rect 259 2336 260 2340
rect 254 2335 260 2336
rect 550 2340 556 2341
rect 550 2336 551 2340
rect 555 2336 556 2340
rect 550 2335 556 2336
rect 862 2340 868 2341
rect 862 2336 863 2340
rect 867 2336 868 2340
rect 862 2335 868 2336
rect 1182 2340 1188 2341
rect 1182 2336 1183 2340
rect 1187 2336 1188 2340
rect 1182 2335 1188 2336
rect 1510 2340 1516 2341
rect 1510 2336 1511 2340
rect 1515 2336 1516 2340
rect 1510 2335 1516 2336
rect 1814 2340 1820 2341
rect 1814 2336 1815 2340
rect 1819 2336 1820 2340
rect 1814 2335 1820 2336
rect 1934 2339 1940 2340
rect 1934 2335 1935 2339
rect 1939 2335 1940 2339
rect 2090 2339 2091 2343
rect 2095 2339 2096 2343
rect 2679 2343 2685 2344
rect 2679 2342 2680 2343
rect 2637 2340 2680 2342
rect 2090 2338 2096 2339
rect 2162 2339 2168 2340
rect 110 2334 116 2335
rect 1934 2334 1940 2335
rect 2162 2335 2163 2339
rect 2167 2335 2168 2339
rect 2162 2334 2168 2335
rect 2354 2339 2360 2340
rect 2354 2335 2355 2339
rect 2359 2335 2360 2339
rect 2679 2339 2680 2340
rect 2684 2339 2685 2343
rect 2679 2338 2685 2339
rect 2806 2343 2812 2344
rect 2806 2339 2807 2343
rect 2811 2339 2812 2343
rect 3534 2343 3540 2344
rect 2806 2338 2812 2339
rect 3018 2339 3024 2340
rect 2354 2334 2360 2335
rect 3018 2335 3019 2339
rect 3023 2335 3024 2339
rect 3018 2334 3024 2335
rect 3122 2339 3128 2340
rect 3122 2335 3123 2339
rect 3127 2335 3128 2339
rect 3122 2334 3128 2335
rect 3394 2339 3400 2340
rect 3394 2335 3395 2339
rect 3399 2335 3400 2339
rect 3534 2339 3535 2343
rect 3539 2339 3540 2343
rect 3534 2338 3540 2339
rect 3658 2339 3664 2340
rect 3394 2334 3400 2335
rect 3658 2335 3659 2339
rect 3663 2335 3664 2339
rect 3658 2334 3664 2335
rect 4890 2335 4896 2336
rect 4890 2334 4891 2335
rect 4612 2332 4891 2334
rect 4612 2330 4614 2332
rect 4890 2331 4891 2332
rect 4895 2331 4896 2335
rect 4890 2330 4896 2331
rect 5143 2331 5149 2332
rect 5143 2330 5144 2331
rect 4541 2328 4614 2330
rect 5061 2328 5144 2330
rect 4618 2327 4624 2328
rect 4618 2323 4619 2327
rect 4623 2323 4624 2327
rect 4618 2322 4624 2323
rect 4794 2327 4800 2328
rect 4794 2323 4795 2327
rect 4799 2323 4800 2327
rect 5143 2327 5144 2328
rect 5148 2327 5149 2331
rect 5326 2331 5332 2332
rect 5326 2330 5327 2331
rect 5245 2328 5327 2330
rect 5143 2326 5149 2327
rect 5326 2327 5327 2328
rect 5331 2327 5332 2331
rect 5326 2326 5332 2327
rect 5434 2331 5440 2332
rect 5434 2327 5435 2331
rect 5439 2327 5440 2331
rect 5434 2326 5440 2327
rect 5522 2327 5528 2328
rect 4794 2322 4800 2323
rect 5522 2323 5523 2327
rect 5527 2323 5528 2327
rect 5522 2322 5528 2323
rect 3018 2307 3024 2308
rect 3018 2303 3019 2307
rect 3023 2306 3024 2307
rect 3023 2304 3250 2306
rect 3023 2303 3024 2304
rect 3018 2302 3024 2303
rect 2119 2299 2125 2300
rect 2119 2295 2120 2299
rect 2124 2298 2125 2299
rect 2162 2299 2168 2300
rect 2162 2298 2163 2299
rect 2124 2296 2163 2298
rect 2124 2295 2125 2296
rect 2119 2294 2125 2295
rect 2162 2295 2163 2296
rect 2167 2295 2168 2299
rect 2162 2294 2168 2295
rect 2279 2299 2285 2300
rect 2279 2295 2280 2299
rect 2284 2298 2285 2299
rect 2354 2299 2360 2300
rect 2354 2298 2355 2299
rect 2284 2296 2355 2298
rect 2284 2295 2285 2296
rect 2279 2294 2285 2295
rect 2354 2295 2355 2296
rect 2359 2295 2360 2299
rect 2354 2294 2360 2295
rect 2470 2299 2477 2300
rect 2470 2295 2471 2299
rect 2476 2295 2477 2299
rect 2470 2294 2477 2295
rect 2546 2299 2552 2300
rect 2546 2295 2547 2299
rect 2551 2298 2552 2299
rect 2663 2299 2669 2300
rect 2663 2298 2664 2299
rect 2551 2296 2664 2298
rect 2551 2295 2552 2296
rect 2546 2294 2552 2295
rect 2663 2295 2664 2296
rect 2668 2295 2669 2299
rect 2663 2294 2669 2295
rect 2679 2299 2685 2300
rect 2679 2295 2680 2299
rect 2684 2298 2685 2299
rect 2855 2299 2861 2300
rect 2855 2298 2856 2299
rect 2684 2296 2856 2298
rect 2684 2295 2685 2296
rect 2679 2294 2685 2295
rect 2855 2295 2856 2296
rect 2860 2295 2861 2299
rect 2855 2294 2861 2295
rect 3047 2299 3053 2300
rect 3047 2295 3048 2299
rect 3052 2298 3053 2299
rect 3122 2299 3128 2300
rect 3122 2298 3123 2299
rect 3052 2296 3123 2298
rect 3052 2295 3053 2296
rect 3047 2294 3053 2295
rect 3122 2295 3123 2296
rect 3127 2295 3128 2299
rect 3122 2294 3128 2295
rect 3238 2299 3245 2300
rect 3238 2295 3239 2299
rect 3244 2295 3245 2299
rect 3248 2298 3250 2304
rect 3423 2299 3429 2300
rect 3423 2298 3424 2299
rect 3248 2296 3424 2298
rect 3238 2294 3245 2295
rect 3423 2295 3424 2296
rect 3428 2295 3429 2299
rect 3423 2294 3429 2295
rect 3607 2299 3613 2300
rect 3607 2295 3608 2299
rect 3612 2298 3613 2299
rect 3658 2299 3664 2300
rect 3658 2298 3659 2299
rect 3612 2296 3659 2298
rect 3612 2295 3613 2296
rect 3607 2294 3613 2295
rect 3658 2295 3659 2296
rect 3663 2295 3664 2299
rect 3658 2294 3664 2295
rect 3746 2299 3752 2300
rect 3746 2295 3747 2299
rect 3751 2298 3752 2299
rect 3775 2299 3781 2300
rect 3775 2298 3776 2299
rect 3751 2296 3776 2298
rect 3751 2295 3752 2296
rect 3746 2294 3752 2295
rect 3775 2295 3776 2296
rect 3780 2295 3781 2299
rect 3775 2294 3781 2295
rect 1974 2292 1980 2293
rect 3798 2292 3804 2293
rect 1974 2288 1975 2292
rect 1979 2288 1980 2292
rect 1974 2287 1980 2288
rect 1994 2291 2000 2292
rect 1994 2287 1995 2291
rect 1999 2287 2000 2291
rect 1994 2286 2000 2287
rect 2154 2291 2160 2292
rect 2154 2287 2155 2291
rect 2159 2287 2160 2291
rect 2154 2286 2160 2287
rect 2346 2291 2352 2292
rect 2346 2287 2347 2291
rect 2351 2287 2352 2291
rect 2346 2286 2352 2287
rect 2538 2291 2544 2292
rect 2538 2287 2539 2291
rect 2543 2287 2544 2291
rect 2538 2286 2544 2287
rect 2730 2291 2736 2292
rect 2730 2287 2731 2291
rect 2735 2287 2736 2291
rect 2730 2286 2736 2287
rect 2922 2291 2928 2292
rect 2922 2287 2923 2291
rect 2927 2287 2928 2291
rect 2922 2286 2928 2287
rect 3114 2291 3120 2292
rect 3114 2287 3115 2291
rect 3119 2287 3120 2291
rect 3114 2286 3120 2287
rect 3298 2291 3304 2292
rect 3298 2287 3299 2291
rect 3303 2287 3304 2291
rect 3298 2286 3304 2287
rect 3482 2291 3488 2292
rect 3482 2287 3483 2291
rect 3487 2287 3488 2291
rect 3482 2286 3488 2287
rect 3650 2291 3656 2292
rect 3650 2287 3651 2291
rect 3655 2287 3656 2291
rect 3798 2288 3799 2292
rect 3803 2288 3804 2292
rect 4911 2288 4917 2289
rect 3798 2287 3804 2288
rect 4567 2287 4573 2288
rect 3650 2286 3656 2287
rect 4567 2283 4568 2287
rect 4572 2286 4573 2287
rect 4618 2287 4624 2288
rect 4618 2286 4619 2287
rect 4572 2284 4619 2286
rect 4572 2283 4573 2284
rect 4567 2282 4573 2283
rect 4618 2283 4619 2284
rect 4623 2283 4624 2287
rect 4618 2282 4624 2283
rect 4735 2287 4741 2288
rect 4735 2283 4736 2287
rect 4740 2286 4741 2287
rect 4794 2287 4800 2288
rect 4794 2286 4795 2287
rect 4740 2284 4795 2286
rect 4740 2283 4741 2284
rect 4735 2282 4741 2283
rect 4794 2283 4795 2284
rect 4799 2283 4800 2287
rect 4794 2282 4800 2283
rect 4902 2287 4908 2288
rect 4902 2283 4903 2287
rect 4907 2286 4908 2287
rect 4911 2286 4912 2288
rect 4907 2284 4912 2286
rect 4916 2284 4917 2288
rect 4907 2283 4908 2284
rect 4911 2283 4917 2284
rect 5087 2287 5093 2288
rect 5087 2283 5088 2287
rect 5092 2286 5093 2287
rect 5098 2287 5104 2288
rect 5098 2286 5099 2287
rect 5092 2284 5099 2286
rect 5092 2283 5093 2284
rect 4902 2282 4908 2283
rect 5087 2282 5093 2283
rect 5098 2283 5099 2284
rect 5103 2283 5104 2287
rect 5098 2282 5104 2283
rect 5143 2287 5149 2288
rect 5143 2283 5144 2287
rect 5148 2286 5149 2287
rect 5271 2287 5277 2288
rect 5271 2286 5272 2287
rect 5148 2284 5272 2286
rect 5148 2283 5149 2284
rect 5143 2282 5149 2283
rect 5271 2283 5272 2284
rect 5276 2283 5277 2287
rect 5271 2282 5277 2283
rect 5463 2287 5469 2288
rect 5463 2283 5464 2287
rect 5468 2286 5469 2287
rect 5522 2287 5528 2288
rect 5522 2286 5523 2287
rect 5468 2284 5523 2286
rect 5468 2283 5469 2284
rect 5463 2282 5469 2283
rect 5522 2283 5523 2284
rect 5527 2283 5528 2287
rect 5522 2282 5528 2283
rect 5610 2287 5616 2288
rect 5610 2283 5611 2287
rect 5615 2286 5616 2287
rect 5639 2287 5645 2288
rect 5639 2286 5640 2287
rect 5615 2284 5640 2286
rect 5615 2283 5616 2284
rect 5610 2282 5616 2283
rect 5639 2283 5640 2284
rect 5644 2283 5645 2287
rect 5639 2282 5645 2283
rect 3838 2280 3844 2281
rect 5662 2280 5668 2281
rect 2022 2276 2028 2277
rect 1974 2275 1980 2276
rect 1974 2271 1975 2275
rect 1979 2271 1980 2275
rect 2022 2272 2023 2276
rect 2027 2272 2028 2276
rect 2022 2271 2028 2272
rect 2182 2276 2188 2277
rect 2182 2272 2183 2276
rect 2187 2272 2188 2276
rect 2182 2271 2188 2272
rect 2374 2276 2380 2277
rect 2374 2272 2375 2276
rect 2379 2272 2380 2276
rect 2374 2271 2380 2272
rect 2566 2276 2572 2277
rect 2566 2272 2567 2276
rect 2571 2272 2572 2276
rect 2566 2271 2572 2272
rect 2758 2276 2764 2277
rect 2758 2272 2759 2276
rect 2763 2272 2764 2276
rect 2758 2271 2764 2272
rect 2950 2276 2956 2277
rect 2950 2272 2951 2276
rect 2955 2272 2956 2276
rect 2950 2271 2956 2272
rect 3142 2276 3148 2277
rect 3142 2272 3143 2276
rect 3147 2272 3148 2276
rect 3142 2271 3148 2272
rect 3326 2276 3332 2277
rect 3326 2272 3327 2276
rect 3331 2272 3332 2276
rect 3326 2271 3332 2272
rect 3510 2276 3516 2277
rect 3510 2272 3511 2276
rect 3515 2272 3516 2276
rect 3510 2271 3516 2272
rect 3678 2276 3684 2277
rect 3838 2276 3839 2280
rect 3843 2276 3844 2280
rect 3678 2272 3679 2276
rect 3683 2272 3684 2276
rect 3678 2271 3684 2272
rect 3798 2275 3804 2276
rect 3838 2275 3844 2276
rect 4442 2279 4448 2280
rect 4442 2275 4443 2279
rect 4447 2275 4448 2279
rect 3798 2271 3799 2275
rect 3803 2271 3804 2275
rect 4442 2274 4448 2275
rect 4610 2279 4616 2280
rect 4610 2275 4611 2279
rect 4615 2275 4616 2279
rect 4610 2274 4616 2275
rect 4786 2279 4792 2280
rect 4786 2275 4787 2279
rect 4791 2275 4792 2279
rect 4786 2274 4792 2275
rect 4962 2279 4968 2280
rect 4962 2275 4963 2279
rect 4967 2275 4968 2279
rect 4962 2274 4968 2275
rect 5146 2279 5152 2280
rect 5146 2275 5147 2279
rect 5151 2275 5152 2279
rect 5146 2274 5152 2275
rect 5338 2279 5344 2280
rect 5338 2275 5339 2279
rect 5343 2275 5344 2279
rect 5338 2274 5344 2275
rect 5514 2279 5520 2280
rect 5514 2275 5515 2279
rect 5519 2275 5520 2279
rect 5662 2276 5663 2280
rect 5667 2276 5668 2280
rect 5662 2275 5668 2276
rect 5514 2274 5520 2275
rect 1974 2270 1980 2271
rect 3798 2270 3804 2271
rect 110 2265 116 2266
rect 1934 2265 1940 2266
rect 110 2261 111 2265
rect 115 2261 116 2265
rect 110 2260 116 2261
rect 158 2264 164 2265
rect 158 2260 159 2264
rect 163 2260 164 2264
rect 158 2259 164 2260
rect 366 2264 372 2265
rect 366 2260 367 2264
rect 371 2260 372 2264
rect 366 2259 372 2260
rect 598 2264 604 2265
rect 598 2260 599 2264
rect 603 2260 604 2264
rect 598 2259 604 2260
rect 830 2264 836 2265
rect 830 2260 831 2264
rect 835 2260 836 2264
rect 830 2259 836 2260
rect 1062 2264 1068 2265
rect 1062 2260 1063 2264
rect 1067 2260 1068 2264
rect 1934 2261 1935 2265
rect 1939 2261 1940 2265
rect 4470 2264 4476 2265
rect 1934 2260 1940 2261
rect 3838 2263 3844 2264
rect 1062 2259 1068 2260
rect 3838 2259 3839 2263
rect 3843 2259 3844 2263
rect 4470 2260 4471 2264
rect 4475 2260 4476 2264
rect 4470 2259 4476 2260
rect 4638 2264 4644 2265
rect 4638 2260 4639 2264
rect 4643 2260 4644 2264
rect 4638 2259 4644 2260
rect 4814 2264 4820 2265
rect 4814 2260 4815 2264
rect 4819 2260 4820 2264
rect 4814 2259 4820 2260
rect 4990 2264 4996 2265
rect 4990 2260 4991 2264
rect 4995 2260 4996 2264
rect 4990 2259 4996 2260
rect 5174 2264 5180 2265
rect 5174 2260 5175 2264
rect 5179 2260 5180 2264
rect 5174 2259 5180 2260
rect 5366 2264 5372 2265
rect 5366 2260 5367 2264
rect 5371 2260 5372 2264
rect 5366 2259 5372 2260
rect 5542 2264 5548 2265
rect 5542 2260 5543 2264
rect 5547 2260 5548 2264
rect 5542 2259 5548 2260
rect 5662 2263 5668 2264
rect 5662 2259 5663 2263
rect 5667 2259 5668 2263
rect 3838 2258 3844 2259
rect 5662 2258 5668 2259
rect 130 2249 136 2250
rect 110 2248 116 2249
rect 110 2244 111 2248
rect 115 2244 116 2248
rect 130 2245 131 2249
rect 135 2245 136 2249
rect 130 2244 136 2245
rect 338 2249 344 2250
rect 338 2245 339 2249
rect 343 2245 344 2249
rect 338 2244 344 2245
rect 570 2249 576 2250
rect 570 2245 571 2249
rect 575 2245 576 2249
rect 570 2244 576 2245
rect 802 2249 808 2250
rect 802 2245 803 2249
rect 807 2245 808 2249
rect 802 2244 808 2245
rect 1034 2249 1040 2250
rect 1034 2245 1035 2249
rect 1039 2245 1040 2249
rect 1034 2244 1040 2245
rect 1934 2248 1940 2249
rect 1934 2244 1935 2248
rect 1939 2244 1940 2248
rect 110 2243 116 2244
rect 1934 2243 1940 2244
rect 255 2239 261 2240
rect 255 2235 256 2239
rect 260 2238 261 2239
rect 278 2239 284 2240
rect 278 2238 279 2239
rect 260 2236 279 2238
rect 260 2235 261 2236
rect 255 2234 261 2235
rect 278 2235 279 2236
rect 283 2235 284 2239
rect 278 2234 284 2235
rect 463 2239 472 2240
rect 463 2235 464 2239
rect 471 2235 472 2239
rect 463 2234 472 2235
rect 618 2239 624 2240
rect 618 2235 619 2239
rect 623 2238 624 2239
rect 695 2239 701 2240
rect 695 2238 696 2239
rect 623 2236 696 2238
rect 623 2235 624 2236
rect 618 2234 624 2235
rect 695 2235 696 2236
rect 700 2235 701 2239
rect 695 2234 701 2235
rect 927 2239 936 2240
rect 927 2235 928 2239
rect 935 2235 936 2239
rect 927 2234 936 2235
rect 1158 2239 1165 2240
rect 1158 2235 1159 2239
rect 1164 2235 1165 2239
rect 1158 2234 1165 2235
rect 1974 2209 1980 2210
rect 3798 2209 3804 2210
rect 1974 2205 1975 2209
rect 1979 2205 1980 2209
rect 1974 2204 1980 2205
rect 2022 2208 2028 2209
rect 2022 2204 2023 2208
rect 2027 2204 2028 2208
rect 2022 2203 2028 2204
rect 2190 2208 2196 2209
rect 2190 2204 2191 2208
rect 2195 2204 2196 2208
rect 2190 2203 2196 2204
rect 2358 2208 2364 2209
rect 2358 2204 2359 2208
rect 2363 2204 2364 2208
rect 2358 2203 2364 2204
rect 2534 2208 2540 2209
rect 2534 2204 2535 2208
rect 2539 2204 2540 2208
rect 2534 2203 2540 2204
rect 2710 2208 2716 2209
rect 2710 2204 2711 2208
rect 2715 2204 2716 2208
rect 2710 2203 2716 2204
rect 2878 2208 2884 2209
rect 2878 2204 2879 2208
rect 2883 2204 2884 2208
rect 2878 2203 2884 2204
rect 3046 2208 3052 2209
rect 3046 2204 3047 2208
rect 3051 2204 3052 2208
rect 3046 2203 3052 2204
rect 3206 2208 3212 2209
rect 3206 2204 3207 2208
rect 3211 2204 3212 2208
rect 3206 2203 3212 2204
rect 3366 2208 3372 2209
rect 3366 2204 3367 2208
rect 3371 2204 3372 2208
rect 3366 2203 3372 2204
rect 3534 2208 3540 2209
rect 3534 2204 3535 2208
rect 3539 2204 3540 2208
rect 3534 2203 3540 2204
rect 3678 2208 3684 2209
rect 3678 2204 3679 2208
rect 3683 2204 3684 2208
rect 3798 2205 3799 2209
rect 3803 2205 3804 2209
rect 3798 2204 3804 2205
rect 3678 2203 3684 2204
rect 226 2199 232 2200
rect 226 2195 227 2199
rect 231 2195 232 2199
rect 226 2194 232 2195
rect 278 2199 284 2200
rect 278 2195 279 2199
rect 283 2198 284 2199
rect 466 2199 472 2200
rect 283 2196 345 2198
rect 283 2195 284 2196
rect 278 2194 284 2195
rect 466 2195 467 2199
rect 471 2198 472 2199
rect 898 2199 904 2200
rect 471 2196 577 2198
rect 471 2195 472 2196
rect 466 2194 472 2195
rect 898 2195 899 2199
rect 903 2195 904 2199
rect 898 2194 904 2195
rect 930 2199 936 2200
rect 930 2195 931 2199
rect 935 2198 936 2199
rect 935 2196 1041 2198
rect 935 2195 936 2196
rect 930 2194 936 2195
rect 1994 2193 2000 2194
rect 1974 2192 1980 2193
rect 1974 2188 1975 2192
rect 1979 2188 1980 2192
rect 1994 2189 1995 2193
rect 1999 2189 2000 2193
rect 1994 2188 2000 2189
rect 2162 2193 2168 2194
rect 2162 2189 2163 2193
rect 2167 2189 2168 2193
rect 2162 2188 2168 2189
rect 2330 2193 2336 2194
rect 2330 2189 2331 2193
rect 2335 2189 2336 2193
rect 2330 2188 2336 2189
rect 2506 2193 2512 2194
rect 2506 2189 2507 2193
rect 2511 2189 2512 2193
rect 2506 2188 2512 2189
rect 2682 2193 2688 2194
rect 2682 2189 2683 2193
rect 2687 2189 2688 2193
rect 2682 2188 2688 2189
rect 2850 2193 2856 2194
rect 2850 2189 2851 2193
rect 2855 2189 2856 2193
rect 2850 2188 2856 2189
rect 3018 2193 3024 2194
rect 3018 2189 3019 2193
rect 3023 2189 3024 2193
rect 3018 2188 3024 2189
rect 3178 2193 3184 2194
rect 3178 2189 3179 2193
rect 3183 2189 3184 2193
rect 3178 2188 3184 2189
rect 3338 2193 3344 2194
rect 3338 2189 3339 2193
rect 3343 2189 3344 2193
rect 3338 2188 3344 2189
rect 3506 2193 3512 2194
rect 3506 2189 3507 2193
rect 3511 2189 3512 2193
rect 3506 2188 3512 2189
rect 3650 2193 3656 2194
rect 3838 2193 3844 2194
rect 5662 2193 5668 2194
rect 3650 2189 3651 2193
rect 3655 2189 3656 2193
rect 3650 2188 3656 2189
rect 3798 2192 3804 2193
rect 3798 2188 3799 2192
rect 3803 2188 3804 2192
rect 3838 2189 3839 2193
rect 3843 2189 3844 2193
rect 3838 2188 3844 2189
rect 4542 2192 4548 2193
rect 4542 2188 4543 2192
rect 4547 2188 4548 2192
rect 1974 2187 1980 2188
rect 3798 2187 3804 2188
rect 4542 2187 4548 2188
rect 4718 2192 4724 2193
rect 4718 2188 4719 2192
rect 4723 2188 4724 2192
rect 4718 2187 4724 2188
rect 4910 2192 4916 2193
rect 4910 2188 4911 2192
rect 4915 2188 4916 2192
rect 4910 2187 4916 2188
rect 5118 2192 5124 2193
rect 5118 2188 5119 2192
rect 5123 2188 5124 2192
rect 5118 2187 5124 2188
rect 5334 2192 5340 2193
rect 5334 2188 5335 2192
rect 5339 2188 5340 2192
rect 5334 2187 5340 2188
rect 5542 2192 5548 2193
rect 5542 2188 5543 2192
rect 5547 2188 5548 2192
rect 5662 2189 5663 2193
rect 5667 2189 5668 2193
rect 5662 2188 5668 2189
rect 5542 2187 5548 2188
rect 2119 2183 2128 2184
rect 2119 2179 2120 2183
rect 2127 2179 2128 2183
rect 2119 2178 2128 2179
rect 2287 2183 2296 2184
rect 2287 2179 2288 2183
rect 2295 2179 2296 2183
rect 2287 2178 2296 2179
rect 2455 2183 2464 2184
rect 2455 2179 2456 2183
rect 2463 2179 2464 2183
rect 2455 2178 2464 2179
rect 2631 2183 2640 2184
rect 2631 2179 2632 2183
rect 2639 2179 2640 2183
rect 2631 2178 2640 2179
rect 2806 2183 2813 2184
rect 2806 2179 2807 2183
rect 2812 2179 2813 2183
rect 2806 2178 2813 2179
rect 2975 2183 2984 2184
rect 2975 2179 2976 2183
rect 2983 2179 2984 2183
rect 2975 2178 2984 2179
rect 3142 2183 3149 2184
rect 3142 2179 3143 2183
rect 3148 2179 3149 2183
rect 3303 2183 3309 2184
rect 3303 2182 3304 2183
rect 3142 2178 3149 2179
rect 3152 2180 3304 2182
rect 2946 2175 2952 2176
rect 2946 2171 2947 2175
rect 2951 2174 2952 2175
rect 3152 2174 3154 2180
rect 3303 2179 3304 2180
rect 3308 2179 3309 2183
rect 3303 2178 3309 2179
rect 3394 2183 3400 2184
rect 3394 2179 3395 2183
rect 3399 2182 3400 2183
rect 3463 2183 3469 2184
rect 3463 2182 3464 2183
rect 3399 2180 3464 2182
rect 3399 2179 3400 2180
rect 3394 2178 3400 2179
rect 3463 2179 3464 2180
rect 3468 2179 3469 2183
rect 3463 2178 3469 2179
rect 3478 2183 3484 2184
rect 3478 2179 3479 2183
rect 3483 2182 3484 2183
rect 3631 2183 3637 2184
rect 3631 2182 3632 2183
rect 3483 2180 3632 2182
rect 3483 2179 3484 2180
rect 3478 2178 3484 2179
rect 3631 2179 3632 2180
rect 3636 2179 3637 2183
rect 3631 2178 3637 2179
rect 3647 2183 3653 2184
rect 3647 2179 3648 2183
rect 3652 2182 3653 2183
rect 3775 2183 3781 2184
rect 3775 2182 3776 2183
rect 3652 2180 3776 2182
rect 3652 2179 3653 2180
rect 3647 2178 3653 2179
rect 3775 2179 3776 2180
rect 3780 2179 3781 2183
rect 3775 2178 3781 2179
rect 4514 2177 4520 2178
rect 2951 2172 3154 2174
rect 3838 2176 3844 2177
rect 3838 2172 3839 2176
rect 3843 2172 3844 2176
rect 4514 2173 4515 2177
rect 4519 2173 4520 2177
rect 4514 2172 4520 2173
rect 4690 2177 4696 2178
rect 4690 2173 4691 2177
rect 4695 2173 4696 2177
rect 4690 2172 4696 2173
rect 4882 2177 4888 2178
rect 4882 2173 4883 2177
rect 4887 2173 4888 2177
rect 4882 2172 4888 2173
rect 5090 2177 5096 2178
rect 5090 2173 5091 2177
rect 5095 2173 5096 2177
rect 5090 2172 5096 2173
rect 5306 2177 5312 2178
rect 5306 2173 5307 2177
rect 5311 2173 5312 2177
rect 5306 2172 5312 2173
rect 5514 2177 5520 2178
rect 5514 2173 5515 2177
rect 5519 2173 5520 2177
rect 5514 2172 5520 2173
rect 5662 2176 5668 2177
rect 5662 2172 5663 2176
rect 5667 2172 5668 2176
rect 2951 2171 2952 2172
rect 3838 2171 3844 2172
rect 5662 2171 5668 2172
rect 2946 2170 2952 2171
rect 4639 2167 4648 2168
rect 4639 2163 4640 2167
rect 4647 2163 4648 2167
rect 4639 2162 4648 2163
rect 4670 2167 4676 2168
rect 4670 2163 4671 2167
rect 4675 2166 4676 2167
rect 4815 2167 4821 2168
rect 4815 2166 4816 2167
rect 4675 2164 4816 2166
rect 4675 2163 4676 2164
rect 4670 2162 4676 2163
rect 4815 2163 4816 2164
rect 4820 2163 4821 2167
rect 4815 2162 4821 2163
rect 4847 2167 4853 2168
rect 4847 2163 4848 2167
rect 4852 2166 4853 2167
rect 5007 2167 5013 2168
rect 5007 2166 5008 2167
rect 4852 2164 5008 2166
rect 4852 2163 4853 2164
rect 4847 2162 4853 2163
rect 5007 2163 5008 2164
rect 5012 2163 5013 2167
rect 5007 2162 5013 2163
rect 5215 2167 5221 2168
rect 5215 2163 5216 2167
rect 5220 2166 5221 2167
rect 5278 2167 5284 2168
rect 5278 2166 5279 2167
rect 5220 2164 5279 2166
rect 5220 2163 5221 2164
rect 5215 2162 5221 2163
rect 5278 2163 5279 2164
rect 5283 2163 5284 2167
rect 5278 2162 5284 2163
rect 5326 2167 5332 2168
rect 5326 2163 5327 2167
rect 5331 2166 5332 2167
rect 5431 2167 5437 2168
rect 5431 2166 5432 2167
rect 5331 2164 5432 2166
rect 5331 2163 5332 2164
rect 5326 2162 5332 2163
rect 5431 2163 5432 2164
rect 5436 2163 5437 2167
rect 5431 2162 5437 2163
rect 5638 2167 5645 2168
rect 5638 2163 5639 2167
rect 5644 2163 5645 2167
rect 5638 2162 5645 2163
rect 338 2155 344 2156
rect 338 2154 339 2155
rect 229 2152 339 2154
rect 338 2151 339 2152
rect 343 2151 344 2155
rect 591 2155 597 2156
rect 591 2154 592 2155
rect 445 2152 592 2154
rect 338 2150 344 2151
rect 591 2151 592 2152
rect 596 2151 597 2155
rect 591 2150 597 2151
rect 638 2155 644 2156
rect 638 2151 639 2155
rect 643 2151 644 2155
rect 967 2155 973 2156
rect 967 2154 968 2155
rect 933 2152 968 2154
rect 638 2150 644 2151
rect 967 2151 968 2152
rect 972 2151 973 2155
rect 967 2150 973 2151
rect 1158 2155 1164 2156
rect 1158 2151 1159 2155
rect 1163 2151 1164 2155
rect 1559 2155 1565 2156
rect 1559 2154 1560 2155
rect 1413 2152 1560 2154
rect 1158 2150 1164 2151
rect 1559 2151 1560 2152
rect 1564 2151 1565 2155
rect 1783 2155 1789 2156
rect 1783 2154 1784 2155
rect 1661 2152 1784 2154
rect 1559 2150 1565 2151
rect 1783 2151 1784 2152
rect 1788 2151 1789 2155
rect 1783 2150 1789 2151
rect 1794 2151 1800 2152
rect 1794 2147 1795 2151
rect 1799 2147 1800 2151
rect 1794 2146 1800 2147
rect 2122 2143 2128 2144
rect 2092 2134 2094 2141
rect 2122 2139 2123 2143
rect 2127 2142 2128 2143
rect 2290 2143 2296 2144
rect 2127 2140 2169 2142
rect 2127 2139 2128 2140
rect 2122 2138 2128 2139
rect 2290 2139 2291 2143
rect 2295 2142 2296 2143
rect 2458 2143 2464 2144
rect 2295 2140 2337 2142
rect 2295 2139 2296 2140
rect 2290 2138 2296 2139
rect 2458 2139 2459 2143
rect 2463 2142 2464 2143
rect 2634 2143 2640 2144
rect 2463 2140 2513 2142
rect 2463 2139 2464 2140
rect 2458 2138 2464 2139
rect 2634 2139 2635 2143
rect 2639 2142 2640 2143
rect 2946 2143 2952 2144
rect 2639 2140 2689 2142
rect 2639 2139 2640 2140
rect 2634 2138 2640 2139
rect 2946 2139 2947 2143
rect 2951 2139 2952 2143
rect 2946 2138 2952 2139
rect 2978 2143 2984 2144
rect 2978 2139 2979 2143
rect 2983 2142 2984 2143
rect 3238 2143 3244 2144
rect 2983 2140 3025 2142
rect 2983 2139 2984 2140
rect 2978 2138 2984 2139
rect 3238 2139 3239 2143
rect 3243 2139 3244 2143
rect 3478 2143 3484 2144
rect 3478 2142 3479 2143
rect 3437 2140 3479 2142
rect 3238 2138 3244 2139
rect 3478 2139 3479 2140
rect 3483 2139 3484 2143
rect 3647 2143 3653 2144
rect 3647 2142 3648 2143
rect 3605 2140 3648 2142
rect 3478 2138 3484 2139
rect 3647 2139 3648 2140
rect 3652 2139 3653 2143
rect 3647 2138 3653 2139
rect 3746 2143 3752 2144
rect 3746 2139 3747 2143
rect 3751 2139 3752 2143
rect 3746 2138 3752 2139
rect 2470 2135 2476 2136
rect 2470 2134 2471 2135
rect 2092 2132 2471 2134
rect 2470 2131 2471 2132
rect 2475 2131 2476 2135
rect 2470 2130 2476 2131
rect 4670 2127 4676 2128
rect 4670 2126 4671 2127
rect 4613 2124 4671 2126
rect 4670 2123 4671 2124
rect 4675 2123 4676 2127
rect 4847 2127 4853 2128
rect 4847 2126 4848 2127
rect 4789 2124 4848 2126
rect 4670 2122 4676 2123
rect 4847 2123 4848 2124
rect 4852 2123 4853 2127
rect 4847 2122 4853 2123
rect 4902 2127 4908 2128
rect 4902 2123 4903 2127
rect 4907 2123 4908 2127
rect 4902 2122 4908 2123
rect 5166 2127 5172 2128
rect 5166 2123 5167 2127
rect 5171 2123 5172 2127
rect 5166 2122 5172 2123
rect 5278 2127 5284 2128
rect 5278 2123 5279 2127
rect 5283 2126 5284 2127
rect 5610 2127 5616 2128
rect 5283 2124 5313 2126
rect 5283 2123 5284 2124
rect 5278 2122 5284 2123
rect 5610 2123 5611 2127
rect 5615 2123 5616 2127
rect 5610 2122 5616 2123
rect 226 2111 232 2112
rect 226 2107 227 2111
rect 231 2110 232 2111
rect 255 2111 261 2112
rect 255 2110 256 2111
rect 231 2108 256 2110
rect 231 2107 232 2108
rect 226 2106 232 2107
rect 255 2107 256 2108
rect 260 2107 261 2111
rect 255 2106 261 2107
rect 338 2111 344 2112
rect 338 2107 339 2111
rect 343 2110 344 2111
rect 471 2111 477 2112
rect 471 2110 472 2111
rect 343 2108 472 2110
rect 343 2107 344 2108
rect 338 2106 344 2107
rect 471 2107 472 2108
rect 476 2107 477 2111
rect 471 2106 477 2107
rect 591 2111 597 2112
rect 591 2107 592 2111
rect 596 2110 597 2111
rect 719 2111 725 2112
rect 719 2110 720 2111
rect 596 2108 720 2110
rect 596 2107 597 2108
rect 591 2106 597 2107
rect 719 2107 720 2108
rect 724 2107 725 2111
rect 719 2106 725 2107
rect 958 2111 965 2112
rect 958 2107 959 2111
rect 964 2107 965 2111
rect 958 2106 965 2107
rect 967 2111 973 2112
rect 967 2107 968 2111
rect 972 2110 973 2111
rect 1199 2111 1205 2112
rect 1199 2110 1200 2111
rect 972 2108 1200 2110
rect 972 2107 973 2108
rect 967 2106 973 2107
rect 1199 2107 1200 2108
rect 1204 2107 1205 2111
rect 1199 2106 1205 2107
rect 1438 2111 1445 2112
rect 1438 2107 1439 2111
rect 1444 2107 1445 2111
rect 1438 2106 1445 2107
rect 1559 2111 1565 2112
rect 1559 2107 1560 2111
rect 1564 2110 1565 2111
rect 1687 2111 1693 2112
rect 1687 2110 1688 2111
rect 1564 2108 1688 2110
rect 1564 2107 1565 2108
rect 1559 2106 1565 2107
rect 1687 2107 1688 2108
rect 1692 2107 1693 2111
rect 1687 2106 1693 2107
rect 1783 2111 1789 2112
rect 1783 2107 1784 2111
rect 1788 2110 1789 2111
rect 1911 2111 1917 2112
rect 1911 2110 1912 2111
rect 1788 2108 1912 2110
rect 1788 2107 1789 2108
rect 1783 2106 1789 2107
rect 1911 2107 1912 2108
rect 1916 2107 1917 2111
rect 1911 2106 1917 2107
rect 110 2104 116 2105
rect 1934 2104 1940 2105
rect 110 2100 111 2104
rect 115 2100 116 2104
rect 110 2099 116 2100
rect 130 2103 136 2104
rect 130 2099 131 2103
rect 135 2099 136 2103
rect 130 2098 136 2099
rect 346 2103 352 2104
rect 346 2099 347 2103
rect 351 2099 352 2103
rect 346 2098 352 2099
rect 594 2103 600 2104
rect 594 2099 595 2103
rect 599 2099 600 2103
rect 594 2098 600 2099
rect 834 2103 840 2104
rect 834 2099 835 2103
rect 839 2099 840 2103
rect 834 2098 840 2099
rect 1074 2103 1080 2104
rect 1074 2099 1075 2103
rect 1079 2099 1080 2103
rect 1074 2098 1080 2099
rect 1314 2103 1320 2104
rect 1314 2099 1315 2103
rect 1319 2099 1320 2103
rect 1314 2098 1320 2099
rect 1562 2103 1568 2104
rect 1562 2099 1563 2103
rect 1567 2099 1568 2103
rect 1562 2098 1568 2099
rect 1786 2103 1792 2104
rect 1786 2099 1787 2103
rect 1791 2099 1792 2103
rect 1934 2100 1935 2104
rect 1939 2100 1940 2104
rect 1934 2099 1940 2100
rect 3766 2099 3772 2100
rect 1786 2098 1792 2099
rect 3766 2098 3767 2099
rect 3619 2096 3767 2098
rect 3142 2095 3148 2096
rect 3142 2091 3143 2095
rect 3147 2091 3148 2095
rect 3619 2094 3621 2096
rect 3766 2095 3767 2096
rect 3771 2095 3772 2099
rect 3766 2094 3772 2095
rect 4642 2095 4648 2096
rect 3613 2092 3621 2094
rect 3142 2090 3148 2091
rect 3250 2091 3256 2092
rect 158 2088 164 2089
rect 110 2087 116 2088
rect 110 2083 111 2087
rect 115 2083 116 2087
rect 158 2084 159 2088
rect 163 2084 164 2088
rect 158 2083 164 2084
rect 374 2088 380 2089
rect 374 2084 375 2088
rect 379 2084 380 2088
rect 374 2083 380 2084
rect 622 2088 628 2089
rect 622 2084 623 2088
rect 627 2084 628 2088
rect 622 2083 628 2084
rect 862 2088 868 2089
rect 862 2084 863 2088
rect 867 2084 868 2088
rect 862 2083 868 2084
rect 1102 2088 1108 2089
rect 1102 2084 1103 2088
rect 1107 2084 1108 2088
rect 1102 2083 1108 2084
rect 1342 2088 1348 2089
rect 1342 2084 1343 2088
rect 1347 2084 1348 2088
rect 1342 2083 1348 2084
rect 1590 2088 1596 2089
rect 1590 2084 1591 2088
rect 1595 2084 1596 2088
rect 1590 2083 1596 2084
rect 1814 2088 1820 2089
rect 1814 2084 1815 2088
rect 1819 2084 1820 2088
rect 1814 2083 1820 2084
rect 1934 2087 1940 2088
rect 1934 2083 1935 2087
rect 1939 2083 1940 2087
rect 3250 2087 3251 2091
rect 3255 2087 3256 2091
rect 3250 2086 3256 2087
rect 3386 2091 3392 2092
rect 3386 2087 3387 2091
rect 3391 2087 3392 2091
rect 3386 2086 3392 2087
rect 3658 2091 3664 2092
rect 3658 2087 3659 2091
rect 3663 2087 3664 2091
rect 4642 2091 4643 2095
rect 4647 2091 4648 2095
rect 5366 2095 5372 2096
rect 5366 2094 5367 2095
rect 5277 2092 5367 2094
rect 4642 2090 4648 2091
rect 4778 2091 4784 2092
rect 3658 2086 3664 2087
rect 4778 2087 4779 2091
rect 4783 2087 4784 2091
rect 4778 2086 4784 2087
rect 4914 2091 4920 2092
rect 4914 2087 4915 2091
rect 4919 2087 4920 2091
rect 4914 2086 4920 2087
rect 5050 2091 5056 2092
rect 5050 2087 5051 2091
rect 5055 2087 5056 2091
rect 5366 2091 5367 2092
rect 5371 2091 5372 2095
rect 5366 2090 5372 2091
rect 5050 2086 5056 2087
rect 110 2082 116 2083
rect 1934 2082 1940 2083
rect 3231 2051 3237 2052
rect 3231 2047 3232 2051
rect 3236 2050 3237 2051
rect 3250 2051 3256 2052
rect 3250 2050 3251 2051
rect 3236 2048 3251 2050
rect 3236 2047 3237 2048
rect 3231 2046 3237 2047
rect 3250 2047 3251 2048
rect 3255 2047 3256 2051
rect 3250 2046 3256 2047
rect 3367 2051 3373 2052
rect 3367 2047 3368 2051
rect 3372 2050 3373 2051
rect 3386 2051 3392 2052
rect 3386 2050 3387 2051
rect 3372 2048 3387 2050
rect 3372 2047 3373 2048
rect 3367 2046 3373 2047
rect 3386 2047 3387 2048
rect 3391 2047 3392 2051
rect 3386 2046 3392 2047
rect 3466 2051 3472 2052
rect 3466 2047 3467 2051
rect 3471 2050 3472 2051
rect 3503 2051 3509 2052
rect 3503 2050 3504 2051
rect 3471 2048 3504 2050
rect 3471 2047 3472 2048
rect 3466 2046 3472 2047
rect 3503 2047 3504 2048
rect 3508 2047 3509 2051
rect 3503 2046 3509 2047
rect 3639 2051 3645 2052
rect 3639 2047 3640 2051
rect 3644 2050 3645 2051
rect 3658 2051 3664 2052
rect 3658 2050 3659 2051
rect 3644 2048 3659 2050
rect 3644 2047 3645 2048
rect 3639 2046 3645 2047
rect 3658 2047 3659 2048
rect 3663 2047 3664 2051
rect 3658 2046 3664 2047
rect 3746 2051 3752 2052
rect 3746 2047 3747 2051
rect 3751 2050 3752 2051
rect 3775 2051 3781 2052
rect 3775 2050 3776 2051
rect 3751 2048 3776 2050
rect 3751 2047 3752 2048
rect 3746 2046 3752 2047
rect 3775 2047 3776 2048
rect 3780 2047 3781 2051
rect 3775 2046 3781 2047
rect 4759 2051 4765 2052
rect 4759 2047 4760 2051
rect 4764 2050 4765 2051
rect 4778 2051 4784 2052
rect 4778 2050 4779 2051
rect 4764 2048 4779 2050
rect 4764 2047 4765 2048
rect 4759 2046 4765 2047
rect 4778 2047 4779 2048
rect 4783 2047 4784 2051
rect 4778 2046 4784 2047
rect 4895 2051 4901 2052
rect 4895 2047 4896 2051
rect 4900 2050 4901 2051
rect 4914 2051 4920 2052
rect 4914 2050 4915 2051
rect 4900 2048 4915 2050
rect 4900 2047 4901 2048
rect 4895 2046 4901 2047
rect 4914 2047 4915 2048
rect 4919 2047 4920 2051
rect 4914 2046 4920 2047
rect 5031 2051 5037 2052
rect 5031 2047 5032 2051
rect 5036 2050 5037 2051
rect 5050 2051 5056 2052
rect 5050 2050 5051 2051
rect 5036 2048 5051 2050
rect 5036 2047 5037 2048
rect 5031 2046 5037 2047
rect 5050 2047 5051 2048
rect 5055 2047 5056 2051
rect 5050 2046 5056 2047
rect 5166 2051 5173 2052
rect 5166 2047 5167 2051
rect 5172 2047 5173 2051
rect 5166 2046 5173 2047
rect 5218 2051 5224 2052
rect 5218 2047 5219 2051
rect 5223 2050 5224 2051
rect 5303 2051 5309 2052
rect 5303 2050 5304 2051
rect 5223 2048 5304 2050
rect 5223 2047 5224 2048
rect 5218 2046 5224 2047
rect 5303 2047 5304 2048
rect 5308 2047 5309 2051
rect 5303 2046 5309 2047
rect 1974 2044 1980 2045
rect 3798 2044 3804 2045
rect 1974 2040 1975 2044
rect 1979 2040 1980 2044
rect 1974 2039 1980 2040
rect 3106 2043 3112 2044
rect 3106 2039 3107 2043
rect 3111 2039 3112 2043
rect 3106 2038 3112 2039
rect 3242 2043 3248 2044
rect 3242 2039 3243 2043
rect 3247 2039 3248 2043
rect 3242 2038 3248 2039
rect 3378 2043 3384 2044
rect 3378 2039 3379 2043
rect 3383 2039 3384 2043
rect 3378 2038 3384 2039
rect 3514 2043 3520 2044
rect 3514 2039 3515 2043
rect 3519 2039 3520 2043
rect 3514 2038 3520 2039
rect 3650 2043 3656 2044
rect 3650 2039 3651 2043
rect 3655 2039 3656 2043
rect 3798 2040 3799 2044
rect 3803 2040 3804 2044
rect 3798 2039 3804 2040
rect 3838 2044 3844 2045
rect 5662 2044 5668 2045
rect 3838 2040 3839 2044
rect 3843 2040 3844 2044
rect 3838 2039 3844 2040
rect 4634 2043 4640 2044
rect 4634 2039 4635 2043
rect 4639 2039 4640 2043
rect 3650 2038 3656 2039
rect 4634 2038 4640 2039
rect 4770 2043 4776 2044
rect 4770 2039 4771 2043
rect 4775 2039 4776 2043
rect 4770 2038 4776 2039
rect 4906 2043 4912 2044
rect 4906 2039 4907 2043
rect 4911 2039 4912 2043
rect 4906 2038 4912 2039
rect 5042 2043 5048 2044
rect 5042 2039 5043 2043
rect 5047 2039 5048 2043
rect 5042 2038 5048 2039
rect 5178 2043 5184 2044
rect 5178 2039 5179 2043
rect 5183 2039 5184 2043
rect 5662 2040 5663 2044
rect 5667 2040 5668 2044
rect 5662 2039 5668 2040
rect 5178 2038 5184 2039
rect 3134 2028 3140 2029
rect 1974 2027 1980 2028
rect 110 2025 116 2026
rect 1934 2025 1940 2026
rect 110 2021 111 2025
rect 115 2021 116 2025
rect 110 2020 116 2021
rect 270 2024 276 2025
rect 270 2020 271 2024
rect 275 2020 276 2024
rect 270 2019 276 2020
rect 406 2024 412 2025
rect 406 2020 407 2024
rect 411 2020 412 2024
rect 406 2019 412 2020
rect 542 2024 548 2025
rect 542 2020 543 2024
rect 547 2020 548 2024
rect 542 2019 548 2020
rect 686 2024 692 2025
rect 686 2020 687 2024
rect 691 2020 692 2024
rect 686 2019 692 2020
rect 830 2024 836 2025
rect 830 2020 831 2024
rect 835 2020 836 2024
rect 830 2019 836 2020
rect 974 2024 980 2025
rect 974 2020 975 2024
rect 979 2020 980 2024
rect 974 2019 980 2020
rect 1118 2024 1124 2025
rect 1118 2020 1119 2024
rect 1123 2020 1124 2024
rect 1118 2019 1124 2020
rect 1262 2024 1268 2025
rect 1262 2020 1263 2024
rect 1267 2020 1268 2024
rect 1262 2019 1268 2020
rect 1406 2024 1412 2025
rect 1406 2020 1407 2024
rect 1411 2020 1412 2024
rect 1406 2019 1412 2020
rect 1542 2024 1548 2025
rect 1542 2020 1543 2024
rect 1547 2020 1548 2024
rect 1542 2019 1548 2020
rect 1678 2024 1684 2025
rect 1678 2020 1679 2024
rect 1683 2020 1684 2024
rect 1678 2019 1684 2020
rect 1814 2024 1820 2025
rect 1814 2020 1815 2024
rect 1819 2020 1820 2024
rect 1934 2021 1935 2025
rect 1939 2021 1940 2025
rect 1974 2023 1975 2027
rect 1979 2023 1980 2027
rect 3134 2024 3135 2028
rect 3139 2024 3140 2028
rect 3134 2023 3140 2024
rect 3270 2028 3276 2029
rect 3270 2024 3271 2028
rect 3275 2024 3276 2028
rect 3270 2023 3276 2024
rect 3406 2028 3412 2029
rect 3406 2024 3407 2028
rect 3411 2024 3412 2028
rect 3406 2023 3412 2024
rect 3542 2028 3548 2029
rect 3542 2024 3543 2028
rect 3547 2024 3548 2028
rect 3542 2023 3548 2024
rect 3678 2028 3684 2029
rect 4662 2028 4668 2029
rect 3678 2024 3679 2028
rect 3683 2024 3684 2028
rect 3678 2023 3684 2024
rect 3798 2027 3804 2028
rect 3798 2023 3799 2027
rect 3803 2023 3804 2027
rect 1974 2022 1980 2023
rect 3798 2022 3804 2023
rect 3838 2027 3844 2028
rect 3838 2023 3839 2027
rect 3843 2023 3844 2027
rect 4662 2024 4663 2028
rect 4667 2024 4668 2028
rect 4662 2023 4668 2024
rect 4798 2028 4804 2029
rect 4798 2024 4799 2028
rect 4803 2024 4804 2028
rect 4798 2023 4804 2024
rect 4934 2028 4940 2029
rect 4934 2024 4935 2028
rect 4939 2024 4940 2028
rect 4934 2023 4940 2024
rect 5070 2028 5076 2029
rect 5070 2024 5071 2028
rect 5075 2024 5076 2028
rect 5070 2023 5076 2024
rect 5206 2028 5212 2029
rect 5206 2024 5207 2028
rect 5211 2024 5212 2028
rect 5206 2023 5212 2024
rect 5662 2027 5668 2028
rect 5662 2023 5663 2027
rect 5667 2023 5668 2027
rect 3838 2022 3844 2023
rect 5662 2022 5668 2023
rect 1934 2020 1940 2021
rect 1814 2019 1820 2020
rect 242 2009 248 2010
rect 110 2008 116 2009
rect 110 2004 111 2008
rect 115 2004 116 2008
rect 242 2005 243 2009
rect 247 2005 248 2009
rect 242 2004 248 2005
rect 378 2009 384 2010
rect 378 2005 379 2009
rect 383 2005 384 2009
rect 378 2004 384 2005
rect 514 2009 520 2010
rect 514 2005 515 2009
rect 519 2005 520 2009
rect 514 2004 520 2005
rect 658 2009 664 2010
rect 658 2005 659 2009
rect 663 2005 664 2009
rect 658 2004 664 2005
rect 802 2009 808 2010
rect 802 2005 803 2009
rect 807 2005 808 2009
rect 802 2004 808 2005
rect 946 2009 952 2010
rect 946 2005 947 2009
rect 951 2005 952 2009
rect 946 2004 952 2005
rect 1090 2009 1096 2010
rect 1090 2005 1091 2009
rect 1095 2005 1096 2009
rect 1090 2004 1096 2005
rect 1234 2009 1240 2010
rect 1234 2005 1235 2009
rect 1239 2005 1240 2009
rect 1234 2004 1240 2005
rect 1378 2009 1384 2010
rect 1378 2005 1379 2009
rect 1383 2005 1384 2009
rect 1378 2004 1384 2005
rect 1514 2009 1520 2010
rect 1514 2005 1515 2009
rect 1519 2005 1520 2009
rect 1514 2004 1520 2005
rect 1650 2009 1656 2010
rect 1650 2005 1651 2009
rect 1655 2005 1656 2009
rect 1650 2004 1656 2005
rect 1786 2009 1792 2010
rect 1786 2005 1787 2009
rect 1791 2005 1792 2009
rect 1786 2004 1792 2005
rect 1934 2008 1940 2009
rect 1934 2004 1935 2008
rect 1939 2004 1940 2008
rect 110 2003 116 2004
rect 1934 2003 1940 2004
rect 367 1999 376 2000
rect 367 1995 368 1999
rect 375 1995 376 1999
rect 367 1994 376 1995
rect 503 1999 512 2000
rect 503 1995 504 1999
rect 511 1995 512 1999
rect 503 1994 512 1995
rect 638 1999 645 2000
rect 638 1995 639 1999
rect 644 1995 645 1999
rect 638 1994 645 1995
rect 682 1999 688 2000
rect 682 1995 683 1999
rect 687 1998 688 1999
rect 783 1999 789 2000
rect 783 1998 784 1999
rect 687 1996 784 1998
rect 687 1995 688 1996
rect 682 1994 688 1995
rect 783 1995 784 1996
rect 788 1995 789 1999
rect 783 1994 789 1995
rect 799 1999 805 2000
rect 799 1995 800 1999
rect 804 1998 805 1999
rect 927 1999 933 2000
rect 927 1998 928 1999
rect 804 1996 928 1998
rect 804 1995 805 1996
rect 799 1994 805 1995
rect 927 1995 928 1996
rect 932 1995 933 1999
rect 927 1994 933 1995
rect 943 1999 949 2000
rect 943 1995 944 1999
rect 948 1998 949 1999
rect 1071 1999 1077 2000
rect 1071 1998 1072 1999
rect 948 1996 1072 1998
rect 948 1995 949 1996
rect 943 1994 949 1995
rect 1071 1995 1072 1996
rect 1076 1995 1077 1999
rect 1071 1994 1077 1995
rect 1215 1999 1224 2000
rect 1215 1995 1216 1999
rect 1223 1995 1224 1999
rect 1215 1994 1224 1995
rect 1358 1999 1365 2000
rect 1358 1995 1359 1999
rect 1364 1995 1365 1999
rect 1358 1994 1365 1995
rect 1503 1999 1512 2000
rect 1503 1995 1504 1999
rect 1511 1995 1512 1999
rect 1639 1999 1645 2000
rect 1639 1998 1640 1999
rect 1503 1994 1512 1995
rect 1548 1996 1640 1998
rect 1186 1991 1192 1992
rect 1186 1987 1187 1991
rect 1191 1990 1192 1991
rect 1548 1990 1550 1996
rect 1639 1995 1640 1996
rect 1644 1995 1645 1999
rect 1639 1994 1645 1995
rect 1775 1999 1781 2000
rect 1775 1995 1776 1999
rect 1780 1998 1781 1999
rect 1794 1999 1800 2000
rect 1794 1998 1795 1999
rect 1780 1996 1795 1998
rect 1780 1995 1781 1996
rect 1775 1994 1781 1995
rect 1794 1995 1795 1996
rect 1799 1995 1800 1999
rect 1794 1994 1800 1995
rect 1911 1999 1917 2000
rect 1911 1995 1912 1999
rect 1916 1995 1917 1999
rect 1911 1994 1917 1995
rect 1191 1988 1550 1990
rect 1746 1991 1752 1992
rect 1191 1987 1192 1988
rect 1186 1986 1192 1987
rect 1746 1987 1747 1991
rect 1751 1990 1752 1991
rect 1913 1990 1915 1994
rect 1751 1988 1915 1990
rect 1751 1987 1752 1988
rect 1746 1986 1752 1987
rect 1974 1969 1980 1970
rect 3798 1969 3804 1970
rect 1974 1965 1975 1969
rect 1979 1965 1980 1969
rect 1974 1964 1980 1965
rect 3126 1968 3132 1969
rect 3126 1964 3127 1968
rect 3131 1964 3132 1968
rect 3126 1963 3132 1964
rect 3262 1968 3268 1969
rect 3262 1964 3263 1968
rect 3267 1964 3268 1968
rect 3262 1963 3268 1964
rect 3398 1968 3404 1969
rect 3398 1964 3399 1968
rect 3403 1964 3404 1968
rect 3398 1963 3404 1964
rect 3534 1968 3540 1969
rect 3534 1964 3535 1968
rect 3539 1964 3540 1968
rect 3534 1963 3540 1964
rect 3670 1968 3676 1969
rect 3670 1964 3671 1968
rect 3675 1964 3676 1968
rect 3798 1965 3799 1969
rect 3803 1965 3804 1969
rect 3798 1964 3804 1965
rect 3838 1969 3844 1970
rect 5662 1969 5668 1970
rect 3838 1965 3839 1969
rect 3843 1965 3844 1969
rect 3838 1964 3844 1965
rect 4862 1968 4868 1969
rect 4862 1964 4863 1968
rect 4867 1964 4868 1968
rect 3670 1963 3676 1964
rect 4862 1963 4868 1964
rect 4998 1968 5004 1969
rect 4998 1964 4999 1968
rect 5003 1964 5004 1968
rect 4998 1963 5004 1964
rect 5134 1968 5140 1969
rect 5134 1964 5135 1968
rect 5139 1964 5140 1968
rect 5134 1963 5140 1964
rect 5270 1968 5276 1969
rect 5270 1964 5271 1968
rect 5275 1964 5276 1968
rect 5270 1963 5276 1964
rect 5406 1968 5412 1969
rect 5406 1964 5407 1968
rect 5411 1964 5412 1968
rect 5406 1963 5412 1964
rect 5542 1968 5548 1969
rect 5542 1964 5543 1968
rect 5547 1964 5548 1968
rect 5662 1965 5663 1969
rect 5667 1965 5668 1969
rect 5662 1964 5668 1965
rect 5542 1963 5548 1964
rect 310 1959 316 1960
rect 310 1955 311 1959
rect 315 1955 316 1959
rect 310 1954 316 1955
rect 370 1959 376 1960
rect 370 1955 371 1959
rect 375 1958 376 1959
rect 506 1959 512 1960
rect 375 1956 385 1958
rect 375 1955 376 1956
rect 370 1954 376 1955
rect 506 1955 507 1959
rect 511 1958 512 1959
rect 799 1959 805 1960
rect 799 1958 800 1959
rect 511 1956 521 1958
rect 757 1956 800 1958
rect 511 1955 512 1956
rect 506 1954 512 1955
rect 799 1955 800 1956
rect 804 1955 805 1959
rect 943 1959 949 1960
rect 943 1958 944 1959
rect 901 1956 944 1958
rect 799 1954 805 1955
rect 943 1955 944 1956
rect 948 1955 949 1959
rect 943 1954 949 1955
rect 958 1959 964 1960
rect 958 1955 959 1959
rect 963 1955 964 1959
rect 958 1954 964 1955
rect 1186 1959 1192 1960
rect 1186 1955 1187 1959
rect 1191 1955 1192 1959
rect 1186 1954 1192 1955
rect 1218 1959 1224 1960
rect 1218 1955 1219 1959
rect 1223 1958 1224 1959
rect 1438 1959 1444 1960
rect 1223 1956 1241 1958
rect 1223 1955 1224 1956
rect 1218 1954 1224 1955
rect 1438 1955 1439 1959
rect 1443 1955 1444 1959
rect 1438 1954 1444 1955
rect 1506 1959 1512 1960
rect 1506 1955 1507 1959
rect 1511 1958 1512 1959
rect 1746 1959 1752 1960
rect 1511 1956 1521 1958
rect 1511 1955 1512 1956
rect 1506 1954 1512 1955
rect 1746 1955 1747 1959
rect 1751 1955 1752 1959
rect 1746 1954 1752 1955
rect 1882 1959 1888 1960
rect 1882 1955 1883 1959
rect 1887 1955 1888 1959
rect 1882 1954 1888 1955
rect 3098 1953 3104 1954
rect 1974 1952 1980 1953
rect 1974 1948 1975 1952
rect 1979 1948 1980 1952
rect 3098 1949 3099 1953
rect 3103 1949 3104 1953
rect 3098 1948 3104 1949
rect 3234 1953 3240 1954
rect 3234 1949 3235 1953
rect 3239 1949 3240 1953
rect 3234 1948 3240 1949
rect 3370 1953 3376 1954
rect 3370 1949 3371 1953
rect 3375 1949 3376 1953
rect 3370 1948 3376 1949
rect 3506 1953 3512 1954
rect 3506 1949 3507 1953
rect 3511 1949 3512 1953
rect 3506 1948 3512 1949
rect 3642 1953 3648 1954
rect 4834 1953 4840 1954
rect 3642 1949 3643 1953
rect 3647 1949 3648 1953
rect 3642 1948 3648 1949
rect 3798 1952 3804 1953
rect 3798 1948 3799 1952
rect 3803 1948 3804 1952
rect 1974 1947 1980 1948
rect 3798 1947 3804 1948
rect 3838 1952 3844 1953
rect 3838 1948 3839 1952
rect 3843 1948 3844 1952
rect 4834 1949 4835 1953
rect 4839 1949 4840 1953
rect 4834 1948 4840 1949
rect 4970 1953 4976 1954
rect 4970 1949 4971 1953
rect 4975 1949 4976 1953
rect 4970 1948 4976 1949
rect 5106 1953 5112 1954
rect 5106 1949 5107 1953
rect 5111 1949 5112 1953
rect 5106 1948 5112 1949
rect 5242 1953 5248 1954
rect 5242 1949 5243 1953
rect 5247 1949 5248 1953
rect 5242 1948 5248 1949
rect 5378 1953 5384 1954
rect 5378 1949 5379 1953
rect 5383 1949 5384 1953
rect 5378 1948 5384 1949
rect 5514 1953 5520 1954
rect 5514 1949 5515 1953
rect 5519 1949 5520 1953
rect 5514 1948 5520 1949
rect 5662 1952 5668 1953
rect 5662 1948 5663 1952
rect 5667 1948 5668 1952
rect 3838 1947 3844 1948
rect 5662 1947 5668 1948
rect 3202 1943 3208 1944
rect 3202 1939 3203 1943
rect 3207 1942 3208 1943
rect 3223 1943 3229 1944
rect 3223 1942 3224 1943
rect 3207 1940 3224 1942
rect 3207 1939 3208 1940
rect 3202 1938 3208 1939
rect 3223 1939 3224 1940
rect 3228 1939 3229 1943
rect 3223 1938 3229 1939
rect 3231 1943 3237 1944
rect 3231 1939 3232 1943
rect 3236 1942 3237 1943
rect 3359 1943 3365 1944
rect 3359 1942 3360 1943
rect 3236 1940 3360 1942
rect 3236 1939 3237 1940
rect 3231 1938 3237 1939
rect 3359 1939 3360 1940
rect 3364 1939 3365 1943
rect 3359 1938 3365 1939
rect 3367 1943 3373 1944
rect 3367 1939 3368 1943
rect 3372 1942 3373 1943
rect 3495 1943 3501 1944
rect 3495 1942 3496 1943
rect 3372 1940 3496 1942
rect 3372 1939 3373 1940
rect 3367 1938 3373 1939
rect 3495 1939 3496 1940
rect 3500 1939 3501 1943
rect 3495 1938 3501 1939
rect 3631 1943 3640 1944
rect 3631 1939 3632 1943
rect 3639 1939 3640 1943
rect 3631 1938 3640 1939
rect 3766 1943 3773 1944
rect 3766 1939 3767 1943
rect 3772 1939 3773 1943
rect 3766 1938 3773 1939
rect 4770 1943 4776 1944
rect 4770 1939 4771 1943
rect 4775 1942 4776 1943
rect 4959 1943 4965 1944
rect 4959 1942 4960 1943
rect 4775 1940 4960 1942
rect 4775 1939 4776 1940
rect 4770 1938 4776 1939
rect 4959 1939 4960 1940
rect 4964 1939 4965 1943
rect 4959 1938 4965 1939
rect 4967 1943 4973 1944
rect 4967 1939 4968 1943
rect 4972 1942 4973 1943
rect 5095 1943 5101 1944
rect 5095 1942 5096 1943
rect 4972 1940 5096 1942
rect 4972 1939 4973 1940
rect 4967 1938 4973 1939
rect 5095 1939 5096 1940
rect 5100 1939 5101 1943
rect 5095 1938 5101 1939
rect 5103 1943 5109 1944
rect 5103 1939 5104 1943
rect 5108 1942 5109 1943
rect 5231 1943 5237 1944
rect 5231 1942 5232 1943
rect 5108 1940 5232 1942
rect 5108 1939 5109 1940
rect 5103 1938 5109 1939
rect 5231 1939 5232 1940
rect 5236 1939 5237 1943
rect 5231 1938 5237 1939
rect 5366 1943 5373 1944
rect 5366 1939 5367 1943
rect 5372 1939 5373 1943
rect 5366 1938 5373 1939
rect 5386 1943 5392 1944
rect 5386 1939 5387 1943
rect 5391 1942 5392 1943
rect 5503 1943 5509 1944
rect 5503 1942 5504 1943
rect 5391 1940 5504 1942
rect 5391 1939 5392 1940
rect 5386 1938 5392 1939
rect 5503 1939 5504 1940
rect 5508 1939 5509 1943
rect 5503 1938 5509 1939
rect 5610 1943 5616 1944
rect 5610 1939 5611 1943
rect 5615 1942 5616 1943
rect 5639 1943 5645 1944
rect 5639 1942 5640 1943
rect 5615 1940 5640 1942
rect 5615 1939 5616 1940
rect 5610 1938 5616 1939
rect 5639 1939 5640 1940
rect 5644 1939 5645 1943
rect 5639 1938 5645 1939
rect 375 1923 381 1924
rect 375 1922 376 1923
rect 285 1920 376 1922
rect 375 1919 376 1920
rect 380 1919 381 1923
rect 682 1923 688 1924
rect 375 1918 381 1919
rect 474 1919 480 1920
rect 474 1915 475 1919
rect 479 1915 480 1919
rect 682 1919 683 1923
rect 687 1919 688 1923
rect 1358 1923 1364 1924
rect 682 1918 688 1919
rect 818 1919 824 1920
rect 474 1914 480 1915
rect 818 1915 819 1919
rect 823 1915 824 1919
rect 818 1914 824 1915
rect 1058 1919 1064 1920
rect 1058 1915 1059 1919
rect 1063 1915 1064 1919
rect 1358 1919 1359 1923
rect 1363 1919 1364 1923
rect 2118 1923 2124 1924
rect 2118 1922 2119 1923
rect 1885 1920 2119 1922
rect 1358 1918 1364 1919
rect 1562 1919 1568 1920
rect 1058 1914 1064 1915
rect 1562 1915 1563 1919
rect 1567 1915 1568 1919
rect 2118 1919 2119 1920
rect 2123 1919 2124 1923
rect 2118 1918 2124 1919
rect 1562 1914 1568 1915
rect 5386 1911 5392 1912
rect 5386 1910 5387 1911
rect 5340 1908 5387 1910
rect 3231 1903 3237 1904
rect 3231 1902 3232 1903
rect 3197 1900 3232 1902
rect 3231 1899 3232 1900
rect 3236 1899 3237 1903
rect 3367 1903 3373 1904
rect 3367 1902 3368 1903
rect 3333 1900 3368 1902
rect 3231 1898 3237 1899
rect 3367 1899 3368 1900
rect 3372 1899 3373 1903
rect 3367 1898 3373 1899
rect 3466 1903 3472 1904
rect 3466 1899 3467 1903
rect 3471 1899 3472 1903
rect 3466 1898 3472 1899
rect 3602 1903 3608 1904
rect 3602 1899 3603 1903
rect 3607 1899 3608 1903
rect 3602 1898 3608 1899
rect 3634 1903 3640 1904
rect 3634 1899 3635 1903
rect 3639 1902 3640 1903
rect 4967 1903 4973 1904
rect 4967 1902 4968 1903
rect 3639 1900 3649 1902
rect 4933 1900 4968 1902
rect 3639 1899 3640 1900
rect 3634 1898 3640 1899
rect 4967 1899 4968 1900
rect 4972 1899 4973 1903
rect 5103 1903 5109 1904
rect 5103 1902 5104 1903
rect 5069 1900 5104 1902
rect 4967 1898 4973 1899
rect 5103 1899 5104 1900
rect 5108 1899 5109 1903
rect 5218 1903 5224 1904
rect 5218 1902 5219 1903
rect 5205 1900 5219 1902
rect 5103 1898 5109 1899
rect 5218 1899 5219 1900
rect 5223 1899 5224 1903
rect 5340 1901 5342 1908
rect 5386 1907 5387 1908
rect 5391 1907 5392 1911
rect 5386 1906 5392 1907
rect 5375 1903 5381 1904
rect 5218 1898 5224 1899
rect 5375 1899 5376 1903
rect 5380 1902 5381 1903
rect 5638 1903 5644 1904
rect 5638 1902 5639 1903
rect 5380 1900 5385 1902
rect 5613 1900 5639 1902
rect 5380 1899 5381 1900
rect 5375 1898 5381 1899
rect 5638 1899 5639 1900
rect 5643 1899 5644 1903
rect 5638 1898 5644 1899
rect 310 1879 317 1880
rect 310 1875 311 1879
rect 316 1875 317 1879
rect 310 1874 317 1875
rect 375 1879 381 1880
rect 375 1875 376 1879
rect 380 1878 381 1879
rect 503 1879 509 1880
rect 503 1878 504 1879
rect 380 1876 504 1878
rect 380 1875 381 1876
rect 375 1874 381 1875
rect 503 1875 504 1876
rect 508 1875 509 1879
rect 503 1874 509 1875
rect 711 1879 717 1880
rect 711 1875 712 1879
rect 716 1878 717 1879
rect 818 1879 824 1880
rect 818 1878 819 1879
rect 716 1876 819 1878
rect 716 1875 717 1876
rect 711 1874 717 1875
rect 818 1875 819 1876
rect 823 1875 824 1879
rect 818 1874 824 1875
rect 935 1879 941 1880
rect 935 1875 936 1879
rect 940 1878 941 1879
rect 1058 1879 1064 1880
rect 1058 1878 1059 1879
rect 940 1876 1059 1878
rect 940 1875 941 1876
rect 935 1874 941 1875
rect 1058 1875 1059 1876
rect 1063 1875 1064 1879
rect 1058 1874 1064 1875
rect 1134 1879 1140 1880
rect 1134 1875 1135 1879
rect 1139 1878 1140 1879
rect 1175 1879 1181 1880
rect 1175 1878 1176 1879
rect 1139 1876 1176 1878
rect 1139 1875 1140 1876
rect 1134 1874 1140 1875
rect 1175 1875 1176 1876
rect 1180 1875 1181 1879
rect 1175 1874 1181 1875
rect 1423 1879 1429 1880
rect 1423 1875 1424 1879
rect 1428 1878 1429 1879
rect 1562 1879 1568 1880
rect 1562 1878 1563 1879
rect 1428 1876 1563 1878
rect 1428 1875 1429 1876
rect 1423 1874 1429 1875
rect 1562 1875 1563 1876
rect 1567 1875 1568 1879
rect 1562 1874 1568 1875
rect 1642 1879 1648 1880
rect 1642 1875 1643 1879
rect 1647 1878 1648 1879
rect 1679 1879 1685 1880
rect 1679 1878 1680 1879
rect 1647 1876 1680 1878
rect 1647 1875 1648 1876
rect 1642 1874 1648 1875
rect 1679 1875 1680 1876
rect 1684 1875 1685 1879
rect 1679 1874 1685 1875
rect 1882 1879 1888 1880
rect 1882 1875 1883 1879
rect 1887 1878 1888 1879
rect 1911 1879 1917 1880
rect 1911 1878 1912 1879
rect 1887 1876 1912 1878
rect 1887 1875 1888 1876
rect 1882 1874 1888 1875
rect 1911 1875 1912 1876
rect 1916 1875 1917 1879
rect 1911 1874 1917 1875
rect 110 1872 116 1873
rect 1934 1872 1940 1873
rect 110 1868 111 1872
rect 115 1868 116 1872
rect 110 1867 116 1868
rect 186 1871 192 1872
rect 186 1867 187 1871
rect 191 1867 192 1871
rect 186 1866 192 1867
rect 378 1871 384 1872
rect 378 1867 379 1871
rect 383 1867 384 1871
rect 378 1866 384 1867
rect 586 1871 592 1872
rect 586 1867 587 1871
rect 591 1867 592 1871
rect 586 1866 592 1867
rect 810 1871 816 1872
rect 810 1867 811 1871
rect 815 1867 816 1871
rect 810 1866 816 1867
rect 1050 1871 1056 1872
rect 1050 1867 1051 1871
rect 1055 1867 1056 1871
rect 1050 1866 1056 1867
rect 1298 1871 1304 1872
rect 1298 1867 1299 1871
rect 1303 1867 1304 1871
rect 1298 1866 1304 1867
rect 1554 1871 1560 1872
rect 1554 1867 1555 1871
rect 1559 1867 1560 1871
rect 1554 1866 1560 1867
rect 1786 1871 1792 1872
rect 1786 1867 1787 1871
rect 1791 1867 1792 1871
rect 1934 1868 1935 1872
rect 1939 1868 1940 1872
rect 1934 1867 1940 1868
rect 1786 1866 1792 1867
rect 2218 1859 2224 1860
rect 2218 1858 2219 1859
rect 214 1856 220 1857
rect 110 1855 116 1856
rect 110 1851 111 1855
rect 115 1851 116 1855
rect 214 1852 215 1856
rect 219 1852 220 1856
rect 214 1851 220 1852
rect 406 1856 412 1857
rect 406 1852 407 1856
rect 411 1852 412 1856
rect 406 1851 412 1852
rect 614 1856 620 1857
rect 614 1852 615 1856
rect 619 1852 620 1856
rect 614 1851 620 1852
rect 838 1856 844 1857
rect 838 1852 839 1856
rect 843 1852 844 1856
rect 838 1851 844 1852
rect 1078 1856 1084 1857
rect 1078 1852 1079 1856
rect 1083 1852 1084 1856
rect 1078 1851 1084 1852
rect 1326 1856 1332 1857
rect 1326 1852 1327 1856
rect 1331 1852 1332 1856
rect 1326 1851 1332 1852
rect 1582 1856 1588 1857
rect 1582 1852 1583 1856
rect 1587 1852 1588 1856
rect 1582 1851 1588 1852
rect 1814 1856 1820 1857
rect 2093 1856 2219 1858
rect 1814 1852 1815 1856
rect 1819 1852 1820 1856
rect 1814 1851 1820 1852
rect 1934 1855 1940 1856
rect 1934 1851 1935 1855
rect 1939 1851 1940 1855
rect 2218 1855 2219 1856
rect 2223 1855 2224 1859
rect 2402 1859 2408 1860
rect 2402 1858 2403 1859
rect 2325 1856 2403 1858
rect 2218 1854 2224 1855
rect 2402 1855 2403 1856
rect 2407 1855 2408 1859
rect 2402 1854 2408 1855
rect 2410 1859 2416 1860
rect 2410 1855 2411 1859
rect 2415 1858 2416 1859
rect 3202 1859 3208 1860
rect 2415 1856 2473 1858
rect 2415 1855 2416 1856
rect 2410 1854 2416 1855
rect 2786 1855 2792 1856
rect 110 1850 116 1851
rect 1934 1850 1940 1851
rect 2786 1851 2787 1855
rect 2791 1851 2792 1855
rect 2786 1850 2792 1851
rect 2914 1855 2920 1856
rect 2914 1851 2915 1855
rect 2919 1851 2920 1855
rect 3202 1855 3203 1859
rect 3207 1855 3208 1859
rect 3982 1859 3988 1860
rect 3982 1858 3983 1859
rect 3749 1856 3983 1858
rect 3202 1854 3208 1855
rect 3394 1855 3400 1856
rect 2914 1850 2920 1851
rect 3394 1851 3395 1855
rect 3399 1851 3400 1855
rect 3394 1850 3400 1851
rect 3490 1855 3496 1856
rect 3490 1851 3491 1855
rect 3495 1851 3496 1855
rect 3982 1855 3983 1856
rect 3987 1855 3988 1859
rect 3982 1854 3988 1855
rect 4770 1859 4776 1860
rect 4770 1855 4771 1859
rect 4775 1855 4776 1859
rect 5239 1859 5245 1860
rect 5239 1858 5240 1859
rect 5205 1856 5240 1858
rect 4770 1854 4776 1855
rect 4826 1855 4832 1856
rect 3490 1850 3496 1851
rect 4826 1851 4827 1855
rect 4831 1851 4832 1855
rect 4826 1850 4832 1851
rect 4970 1855 4976 1856
rect 4970 1851 4971 1855
rect 4975 1851 4976 1855
rect 5239 1855 5240 1856
rect 5244 1855 5245 1859
rect 5511 1859 5517 1860
rect 5511 1858 5512 1859
rect 5477 1856 5512 1858
rect 5239 1854 5245 1855
rect 5250 1855 5256 1856
rect 4970 1850 4976 1851
rect 5250 1851 5251 1855
rect 5255 1851 5256 1855
rect 5511 1855 5512 1856
rect 5516 1855 5517 1859
rect 5511 1854 5517 1855
rect 5610 1859 5616 1860
rect 5610 1855 5611 1859
rect 5615 1855 5616 1859
rect 5610 1854 5616 1855
rect 5250 1850 5256 1851
rect 2786 1823 2792 1824
rect 2786 1819 2787 1823
rect 2791 1822 2792 1823
rect 3394 1823 3400 1824
rect 2791 1820 3042 1822
rect 2791 1819 2792 1820
rect 2786 1818 2792 1819
rect 2118 1815 2125 1816
rect 2118 1811 2119 1815
rect 2124 1811 2125 1815
rect 2118 1810 2125 1811
rect 2218 1815 2224 1816
rect 2218 1811 2219 1815
rect 2223 1814 2224 1815
rect 2351 1815 2357 1816
rect 2351 1814 2352 1815
rect 2223 1812 2352 1814
rect 2223 1811 2224 1812
rect 2218 1810 2224 1811
rect 2351 1811 2352 1812
rect 2356 1811 2357 1815
rect 2351 1810 2357 1811
rect 2402 1815 2408 1816
rect 2402 1811 2403 1815
rect 2407 1814 2408 1815
rect 2591 1815 2597 1816
rect 2591 1814 2592 1815
rect 2407 1812 2592 1814
rect 2407 1811 2408 1812
rect 2402 1810 2408 1811
rect 2591 1811 2592 1812
rect 2596 1811 2597 1815
rect 2591 1810 2597 1811
rect 2815 1815 2821 1816
rect 2815 1811 2816 1815
rect 2820 1814 2821 1815
rect 2914 1815 2920 1816
rect 2914 1814 2915 1815
rect 2820 1812 2915 1814
rect 2820 1811 2821 1812
rect 2815 1810 2821 1811
rect 2914 1811 2915 1812
rect 2919 1811 2920 1815
rect 2914 1810 2920 1811
rect 3030 1815 3037 1816
rect 3030 1811 3031 1815
rect 3036 1811 3037 1815
rect 3040 1814 3042 1820
rect 3394 1819 3395 1823
rect 3399 1822 3400 1823
rect 3399 1820 3621 1822
rect 3399 1819 3400 1820
rect 3394 1818 3400 1819
rect 3231 1815 3237 1816
rect 3231 1814 3232 1815
rect 3040 1812 3232 1814
rect 3030 1810 3037 1811
rect 3231 1811 3232 1812
rect 3236 1811 3237 1815
rect 3231 1810 3237 1811
rect 3423 1815 3429 1816
rect 3423 1811 3424 1815
rect 3428 1814 3429 1815
rect 3490 1815 3496 1816
rect 3490 1814 3491 1815
rect 3428 1812 3491 1814
rect 3428 1811 3429 1812
rect 3423 1810 3429 1811
rect 3490 1811 3491 1812
rect 3495 1811 3496 1815
rect 3490 1810 3496 1811
rect 3602 1815 3613 1816
rect 3602 1811 3603 1815
rect 3607 1811 3608 1815
rect 3612 1811 3613 1815
rect 3619 1814 3621 1820
rect 3775 1815 3781 1816
rect 3775 1814 3776 1815
rect 3619 1812 3776 1814
rect 3602 1810 3613 1811
rect 3775 1811 3776 1812
rect 3780 1811 3781 1815
rect 3775 1810 3781 1811
rect 4799 1815 4805 1816
rect 4799 1811 4800 1815
rect 4804 1814 4805 1815
rect 4826 1815 4832 1816
rect 4826 1814 4827 1815
rect 4804 1812 4827 1814
rect 4804 1811 4805 1812
rect 4799 1810 4805 1811
rect 4826 1811 4827 1812
rect 4831 1811 4832 1815
rect 4826 1810 4832 1811
rect 4943 1815 4949 1816
rect 4943 1811 4944 1815
rect 4948 1814 4949 1815
rect 4970 1815 4976 1816
rect 4970 1814 4971 1815
rect 4948 1812 4971 1814
rect 4948 1811 4949 1812
rect 4943 1810 4949 1811
rect 4970 1811 4971 1812
rect 4975 1811 4976 1815
rect 4970 1810 4976 1811
rect 5086 1815 5093 1816
rect 5086 1811 5087 1815
rect 5092 1811 5093 1815
rect 5086 1810 5093 1811
rect 5231 1815 5237 1816
rect 5231 1811 5232 1815
rect 5236 1814 5237 1815
rect 5250 1815 5256 1816
rect 5250 1814 5251 1815
rect 5236 1812 5251 1814
rect 5236 1811 5237 1812
rect 5231 1810 5237 1811
rect 5250 1811 5251 1812
rect 5255 1811 5256 1815
rect 5250 1810 5256 1811
rect 5367 1815 5373 1816
rect 5367 1811 5368 1815
rect 5372 1814 5373 1815
rect 5375 1815 5381 1816
rect 5375 1814 5376 1815
rect 5372 1812 5376 1814
rect 5372 1811 5373 1812
rect 5367 1810 5373 1811
rect 5375 1811 5376 1812
rect 5380 1811 5381 1815
rect 5375 1810 5381 1811
rect 5498 1815 5509 1816
rect 5498 1811 5499 1815
rect 5503 1811 5504 1815
rect 5508 1811 5509 1815
rect 5498 1810 5509 1811
rect 5511 1815 5517 1816
rect 5511 1811 5512 1815
rect 5516 1814 5517 1815
rect 5639 1815 5645 1816
rect 5639 1814 5640 1815
rect 5516 1812 5640 1814
rect 5516 1811 5517 1812
rect 5511 1810 5517 1811
rect 5639 1811 5640 1812
rect 5644 1811 5645 1815
rect 5639 1810 5645 1811
rect 1974 1808 1980 1809
rect 3798 1808 3804 1809
rect 1974 1804 1975 1808
rect 1979 1804 1980 1808
rect 1974 1803 1980 1804
rect 1994 1807 2000 1808
rect 1994 1803 1995 1807
rect 1999 1803 2000 1807
rect 1994 1802 2000 1803
rect 2226 1807 2232 1808
rect 2226 1803 2227 1807
rect 2231 1803 2232 1807
rect 2226 1802 2232 1803
rect 2466 1807 2472 1808
rect 2466 1803 2467 1807
rect 2471 1803 2472 1807
rect 2466 1802 2472 1803
rect 2690 1807 2696 1808
rect 2690 1803 2691 1807
rect 2695 1803 2696 1807
rect 2690 1802 2696 1803
rect 2906 1807 2912 1808
rect 2906 1803 2907 1807
rect 2911 1803 2912 1807
rect 2906 1802 2912 1803
rect 3106 1807 3112 1808
rect 3106 1803 3107 1807
rect 3111 1803 3112 1807
rect 3106 1802 3112 1803
rect 3298 1807 3304 1808
rect 3298 1803 3299 1807
rect 3303 1803 3304 1807
rect 3298 1802 3304 1803
rect 3482 1807 3488 1808
rect 3482 1803 3483 1807
rect 3487 1803 3488 1807
rect 3482 1802 3488 1803
rect 3650 1807 3656 1808
rect 3650 1803 3651 1807
rect 3655 1803 3656 1807
rect 3798 1804 3799 1808
rect 3803 1804 3804 1808
rect 3798 1803 3804 1804
rect 3838 1808 3844 1809
rect 5662 1808 5668 1809
rect 3838 1804 3839 1808
rect 3843 1804 3844 1808
rect 3838 1803 3844 1804
rect 4674 1807 4680 1808
rect 4674 1803 4675 1807
rect 4679 1803 4680 1807
rect 3650 1802 3656 1803
rect 4674 1802 4680 1803
rect 4818 1807 4824 1808
rect 4818 1803 4819 1807
rect 4823 1803 4824 1807
rect 4818 1802 4824 1803
rect 4962 1807 4968 1808
rect 4962 1803 4963 1807
rect 4967 1803 4968 1807
rect 4962 1802 4968 1803
rect 5106 1807 5112 1808
rect 5106 1803 5107 1807
rect 5111 1803 5112 1807
rect 5106 1802 5112 1803
rect 5242 1807 5248 1808
rect 5242 1803 5243 1807
rect 5247 1803 5248 1807
rect 5242 1802 5248 1803
rect 5378 1807 5384 1808
rect 5378 1803 5379 1807
rect 5383 1803 5384 1807
rect 5378 1802 5384 1803
rect 5514 1807 5520 1808
rect 5514 1803 5515 1807
rect 5519 1803 5520 1807
rect 5662 1804 5663 1808
rect 5667 1804 5668 1808
rect 5662 1803 5668 1804
rect 5514 1802 5520 1803
rect 2022 1792 2028 1793
rect 1974 1791 1980 1792
rect 110 1789 116 1790
rect 1934 1789 1940 1790
rect 110 1785 111 1789
rect 115 1785 116 1789
rect 110 1784 116 1785
rect 158 1788 164 1789
rect 158 1784 159 1788
rect 163 1784 164 1788
rect 158 1783 164 1784
rect 374 1788 380 1789
rect 374 1784 375 1788
rect 379 1784 380 1788
rect 374 1783 380 1784
rect 590 1788 596 1789
rect 590 1784 591 1788
rect 595 1784 596 1788
rect 590 1783 596 1784
rect 798 1788 804 1789
rect 798 1784 799 1788
rect 803 1784 804 1788
rect 798 1783 804 1784
rect 998 1788 1004 1789
rect 998 1784 999 1788
rect 1003 1784 1004 1788
rect 998 1783 1004 1784
rect 1190 1788 1196 1789
rect 1190 1784 1191 1788
rect 1195 1784 1196 1788
rect 1190 1783 1196 1784
rect 1382 1788 1388 1789
rect 1382 1784 1383 1788
rect 1387 1784 1388 1788
rect 1382 1783 1388 1784
rect 1574 1788 1580 1789
rect 1574 1784 1575 1788
rect 1579 1784 1580 1788
rect 1934 1785 1935 1789
rect 1939 1785 1940 1789
rect 1974 1787 1975 1791
rect 1979 1787 1980 1791
rect 2022 1788 2023 1792
rect 2027 1788 2028 1792
rect 2022 1787 2028 1788
rect 2254 1792 2260 1793
rect 2254 1788 2255 1792
rect 2259 1788 2260 1792
rect 2254 1787 2260 1788
rect 2494 1792 2500 1793
rect 2494 1788 2495 1792
rect 2499 1788 2500 1792
rect 2494 1787 2500 1788
rect 2718 1792 2724 1793
rect 2718 1788 2719 1792
rect 2723 1788 2724 1792
rect 2718 1787 2724 1788
rect 2934 1792 2940 1793
rect 2934 1788 2935 1792
rect 2939 1788 2940 1792
rect 2934 1787 2940 1788
rect 3134 1792 3140 1793
rect 3134 1788 3135 1792
rect 3139 1788 3140 1792
rect 3134 1787 3140 1788
rect 3326 1792 3332 1793
rect 3326 1788 3327 1792
rect 3331 1788 3332 1792
rect 3326 1787 3332 1788
rect 3510 1792 3516 1793
rect 3510 1788 3511 1792
rect 3515 1788 3516 1792
rect 3510 1787 3516 1788
rect 3678 1792 3684 1793
rect 4702 1792 4708 1793
rect 3678 1788 3679 1792
rect 3683 1788 3684 1792
rect 3678 1787 3684 1788
rect 3798 1791 3804 1792
rect 3798 1787 3799 1791
rect 3803 1787 3804 1791
rect 1974 1786 1980 1787
rect 3798 1786 3804 1787
rect 3838 1791 3844 1792
rect 3838 1787 3839 1791
rect 3843 1787 3844 1791
rect 4702 1788 4703 1792
rect 4707 1788 4708 1792
rect 4702 1787 4708 1788
rect 4846 1792 4852 1793
rect 4846 1788 4847 1792
rect 4851 1788 4852 1792
rect 4846 1787 4852 1788
rect 4990 1792 4996 1793
rect 4990 1788 4991 1792
rect 4995 1788 4996 1792
rect 4990 1787 4996 1788
rect 5134 1792 5140 1793
rect 5134 1788 5135 1792
rect 5139 1788 5140 1792
rect 5134 1787 5140 1788
rect 5270 1792 5276 1793
rect 5270 1788 5271 1792
rect 5275 1788 5276 1792
rect 5270 1787 5276 1788
rect 5406 1792 5412 1793
rect 5406 1788 5407 1792
rect 5411 1788 5412 1792
rect 5406 1787 5412 1788
rect 5542 1792 5548 1793
rect 5542 1788 5543 1792
rect 5547 1788 5548 1792
rect 5542 1787 5548 1788
rect 5662 1791 5668 1792
rect 5662 1787 5663 1791
rect 5667 1787 5668 1791
rect 3838 1786 3844 1787
rect 5662 1786 5668 1787
rect 1934 1784 1940 1785
rect 1574 1783 1580 1784
rect 130 1773 136 1774
rect 110 1772 116 1773
rect 110 1768 111 1772
rect 115 1768 116 1772
rect 130 1769 131 1773
rect 135 1769 136 1773
rect 130 1768 136 1769
rect 346 1773 352 1774
rect 346 1769 347 1773
rect 351 1769 352 1773
rect 346 1768 352 1769
rect 562 1773 568 1774
rect 562 1769 563 1773
rect 567 1769 568 1773
rect 562 1768 568 1769
rect 770 1773 776 1774
rect 770 1769 771 1773
rect 775 1769 776 1773
rect 770 1768 776 1769
rect 970 1773 976 1774
rect 970 1769 971 1773
rect 975 1769 976 1773
rect 970 1768 976 1769
rect 1162 1773 1168 1774
rect 1162 1769 1163 1773
rect 1167 1769 1168 1773
rect 1162 1768 1168 1769
rect 1354 1773 1360 1774
rect 1354 1769 1355 1773
rect 1359 1769 1360 1773
rect 1354 1768 1360 1769
rect 1546 1773 1552 1774
rect 1546 1769 1547 1773
rect 1551 1769 1552 1773
rect 1546 1768 1552 1769
rect 1934 1772 1940 1773
rect 1934 1768 1935 1772
rect 1939 1768 1940 1772
rect 110 1767 116 1768
rect 1934 1767 1940 1768
rect 255 1763 261 1764
rect 255 1759 256 1763
rect 260 1762 261 1763
rect 290 1763 296 1764
rect 290 1762 291 1763
rect 260 1760 291 1762
rect 260 1759 261 1760
rect 255 1758 261 1759
rect 290 1759 291 1760
rect 295 1759 296 1763
rect 290 1758 296 1759
rect 471 1763 480 1764
rect 471 1759 472 1763
rect 479 1759 480 1763
rect 471 1758 480 1759
rect 490 1763 496 1764
rect 490 1759 491 1763
rect 495 1762 496 1763
rect 687 1763 693 1764
rect 687 1762 688 1763
rect 495 1760 688 1762
rect 495 1759 496 1760
rect 490 1758 496 1759
rect 687 1759 688 1760
rect 692 1759 693 1763
rect 687 1758 693 1759
rect 767 1763 773 1764
rect 767 1759 768 1763
rect 772 1762 773 1763
rect 895 1763 901 1764
rect 895 1762 896 1763
rect 772 1760 896 1762
rect 772 1759 773 1760
rect 767 1758 773 1759
rect 895 1759 896 1760
rect 900 1759 901 1763
rect 895 1758 901 1759
rect 1095 1763 1101 1764
rect 1095 1759 1096 1763
rect 1100 1762 1101 1763
rect 1106 1763 1112 1764
rect 1106 1762 1107 1763
rect 1100 1760 1107 1762
rect 1100 1759 1101 1760
rect 1095 1758 1101 1759
rect 1106 1759 1107 1760
rect 1111 1759 1112 1763
rect 1106 1758 1112 1759
rect 1286 1763 1293 1764
rect 1286 1759 1287 1763
rect 1292 1759 1293 1763
rect 1479 1763 1485 1764
rect 1479 1762 1480 1763
rect 1286 1758 1293 1759
rect 1296 1760 1480 1762
rect 1066 1755 1072 1756
rect 1066 1751 1067 1755
rect 1071 1754 1072 1755
rect 1296 1754 1298 1760
rect 1479 1759 1480 1760
rect 1484 1759 1485 1763
rect 1479 1758 1485 1759
rect 1511 1763 1517 1764
rect 1511 1759 1512 1763
rect 1516 1762 1517 1763
rect 1671 1763 1677 1764
rect 1671 1762 1672 1763
rect 1516 1760 1672 1762
rect 1516 1759 1517 1760
rect 1511 1758 1517 1759
rect 1671 1759 1672 1760
rect 1676 1759 1677 1763
rect 1671 1758 1677 1759
rect 1071 1752 1298 1754
rect 1071 1751 1072 1752
rect 1066 1750 1072 1751
rect 1974 1725 1980 1726
rect 3798 1725 3804 1726
rect 226 1723 232 1724
rect 226 1719 227 1723
rect 231 1719 232 1723
rect 226 1718 232 1719
rect 290 1723 296 1724
rect 290 1719 291 1723
rect 295 1722 296 1723
rect 767 1723 773 1724
rect 767 1722 768 1723
rect 295 1720 353 1722
rect 661 1720 768 1722
rect 295 1719 296 1720
rect 290 1718 296 1719
rect 767 1719 768 1720
rect 772 1719 773 1723
rect 1066 1723 1072 1724
rect 767 1718 773 1719
rect 868 1714 870 1721
rect 1066 1719 1067 1723
rect 1071 1719 1072 1723
rect 1066 1718 1072 1719
rect 1106 1723 1112 1724
rect 1106 1719 1107 1723
rect 1111 1722 1112 1723
rect 1511 1723 1517 1724
rect 1511 1722 1512 1723
rect 1111 1720 1169 1722
rect 1453 1720 1512 1722
rect 1111 1719 1112 1720
rect 1106 1718 1112 1719
rect 1511 1719 1512 1720
rect 1516 1719 1517 1723
rect 1511 1718 1517 1719
rect 1642 1723 1648 1724
rect 1642 1719 1643 1723
rect 1647 1719 1648 1723
rect 1974 1721 1975 1725
rect 1979 1721 1980 1725
rect 1974 1720 1980 1721
rect 2022 1724 2028 1725
rect 2022 1720 2023 1724
rect 2027 1720 2028 1724
rect 2022 1719 2028 1720
rect 2158 1724 2164 1725
rect 2158 1720 2159 1724
rect 2163 1720 2164 1724
rect 2158 1719 2164 1720
rect 2310 1724 2316 1725
rect 2310 1720 2311 1724
rect 2315 1720 2316 1724
rect 2310 1719 2316 1720
rect 2470 1724 2476 1725
rect 2470 1720 2471 1724
rect 2475 1720 2476 1724
rect 2470 1719 2476 1720
rect 2638 1724 2644 1725
rect 2638 1720 2639 1724
rect 2643 1720 2644 1724
rect 2638 1719 2644 1720
rect 2806 1724 2812 1725
rect 2806 1720 2807 1724
rect 2811 1720 2812 1724
rect 2806 1719 2812 1720
rect 2974 1724 2980 1725
rect 2974 1720 2975 1724
rect 2979 1720 2980 1724
rect 2974 1719 2980 1720
rect 3150 1724 3156 1725
rect 3150 1720 3151 1724
rect 3155 1720 3156 1724
rect 3798 1721 3799 1725
rect 3803 1721 3804 1725
rect 3798 1720 3804 1721
rect 3150 1719 3156 1720
rect 1642 1718 1648 1719
rect 3838 1717 3844 1718
rect 5662 1717 5668 1718
rect 1134 1715 1140 1716
rect 1134 1714 1135 1715
rect 868 1712 1135 1714
rect 1134 1711 1135 1712
rect 1139 1711 1140 1715
rect 3838 1713 3839 1717
rect 3843 1713 3844 1717
rect 3838 1712 3844 1713
rect 3886 1716 3892 1717
rect 3886 1712 3887 1716
rect 3891 1712 3892 1716
rect 3886 1711 3892 1712
rect 4078 1716 4084 1717
rect 4078 1712 4079 1716
rect 4083 1712 4084 1716
rect 4078 1711 4084 1712
rect 4302 1716 4308 1717
rect 4302 1712 4303 1716
rect 4307 1712 4308 1716
rect 4302 1711 4308 1712
rect 4534 1716 4540 1717
rect 4534 1712 4535 1716
rect 4539 1712 4540 1716
rect 4534 1711 4540 1712
rect 4774 1716 4780 1717
rect 4774 1712 4775 1716
rect 4779 1712 4780 1716
rect 4774 1711 4780 1712
rect 5022 1716 5028 1717
rect 5022 1712 5023 1716
rect 5027 1712 5028 1716
rect 5022 1711 5028 1712
rect 5278 1716 5284 1717
rect 5278 1712 5279 1716
rect 5283 1712 5284 1716
rect 5278 1711 5284 1712
rect 5534 1716 5540 1717
rect 5534 1712 5535 1716
rect 5539 1712 5540 1716
rect 5662 1713 5663 1717
rect 5667 1713 5668 1717
rect 5662 1712 5668 1713
rect 5534 1711 5540 1712
rect 1134 1710 1140 1711
rect 1994 1709 2000 1710
rect 1974 1708 1980 1709
rect 1974 1704 1975 1708
rect 1979 1704 1980 1708
rect 1994 1705 1995 1709
rect 1999 1705 2000 1709
rect 1994 1704 2000 1705
rect 2130 1709 2136 1710
rect 2130 1705 2131 1709
rect 2135 1705 2136 1709
rect 2130 1704 2136 1705
rect 2282 1709 2288 1710
rect 2282 1705 2283 1709
rect 2287 1705 2288 1709
rect 2282 1704 2288 1705
rect 2442 1709 2448 1710
rect 2442 1705 2443 1709
rect 2447 1705 2448 1709
rect 2442 1704 2448 1705
rect 2610 1709 2616 1710
rect 2610 1705 2611 1709
rect 2615 1705 2616 1709
rect 2610 1704 2616 1705
rect 2778 1709 2784 1710
rect 2778 1705 2779 1709
rect 2783 1705 2784 1709
rect 2778 1704 2784 1705
rect 2946 1709 2952 1710
rect 2946 1705 2947 1709
rect 2951 1705 2952 1709
rect 2946 1704 2952 1705
rect 3122 1709 3128 1710
rect 3122 1705 3123 1709
rect 3127 1705 3128 1709
rect 3122 1704 3128 1705
rect 3798 1708 3804 1709
rect 3798 1704 3799 1708
rect 3803 1704 3804 1708
rect 1974 1703 1980 1704
rect 3798 1703 3804 1704
rect 3858 1701 3864 1702
rect 3838 1700 3844 1701
rect 2119 1699 2128 1700
rect 2119 1695 2120 1699
rect 2127 1695 2128 1699
rect 2119 1694 2128 1695
rect 2255 1699 2264 1700
rect 2255 1695 2256 1699
rect 2263 1695 2264 1699
rect 2255 1694 2264 1695
rect 2407 1699 2416 1700
rect 2407 1695 2408 1699
rect 2415 1695 2416 1699
rect 2567 1699 2573 1700
rect 2567 1698 2568 1699
rect 2407 1694 2416 1695
rect 2420 1696 2568 1698
rect 2090 1691 2096 1692
rect 2090 1687 2091 1691
rect 2095 1690 2096 1691
rect 2420 1690 2422 1696
rect 2567 1695 2568 1696
rect 2572 1695 2573 1699
rect 2567 1694 2573 1695
rect 2602 1699 2608 1700
rect 2602 1695 2603 1699
rect 2607 1698 2608 1699
rect 2735 1699 2741 1700
rect 2735 1698 2736 1699
rect 2607 1696 2736 1698
rect 2607 1695 2608 1696
rect 2602 1694 2608 1695
rect 2735 1695 2736 1696
rect 2740 1695 2741 1699
rect 2735 1694 2741 1695
rect 2903 1699 2909 1700
rect 2903 1695 2904 1699
rect 2908 1698 2909 1699
rect 2914 1699 2920 1700
rect 2914 1698 2915 1699
rect 2908 1696 2915 1698
rect 2908 1695 2909 1696
rect 2903 1694 2909 1695
rect 2914 1695 2915 1696
rect 2919 1695 2920 1699
rect 2914 1694 2920 1695
rect 3071 1699 3080 1700
rect 3071 1695 3072 1699
rect 3079 1695 3080 1699
rect 3247 1699 3253 1700
rect 3247 1698 3248 1699
rect 3071 1694 3080 1695
rect 3084 1696 3248 1698
rect 2095 1688 2422 1690
rect 2874 1691 2880 1692
rect 2095 1687 2096 1688
rect 2090 1686 2096 1687
rect 2874 1687 2875 1691
rect 2879 1690 2880 1691
rect 3084 1690 3086 1696
rect 3247 1695 3248 1696
rect 3252 1695 3253 1699
rect 3838 1696 3839 1700
rect 3843 1696 3844 1700
rect 3858 1697 3859 1701
rect 3863 1697 3864 1701
rect 3858 1696 3864 1697
rect 4050 1701 4056 1702
rect 4050 1697 4051 1701
rect 4055 1697 4056 1701
rect 4050 1696 4056 1697
rect 4274 1701 4280 1702
rect 4274 1697 4275 1701
rect 4279 1697 4280 1701
rect 4274 1696 4280 1697
rect 4506 1701 4512 1702
rect 4506 1697 4507 1701
rect 4511 1697 4512 1701
rect 4506 1696 4512 1697
rect 4746 1701 4752 1702
rect 4746 1697 4747 1701
rect 4751 1697 4752 1701
rect 4746 1696 4752 1697
rect 4994 1701 5000 1702
rect 4994 1697 4995 1701
rect 4999 1697 5000 1701
rect 4994 1696 5000 1697
rect 5250 1701 5256 1702
rect 5250 1697 5251 1701
rect 5255 1697 5256 1701
rect 5250 1696 5256 1697
rect 5506 1701 5512 1702
rect 5506 1697 5507 1701
rect 5511 1697 5512 1701
rect 5506 1696 5512 1697
rect 5662 1700 5668 1701
rect 5662 1696 5663 1700
rect 5667 1696 5668 1700
rect 3838 1695 3844 1696
rect 5662 1695 5668 1696
rect 3247 1694 3253 1695
rect 2879 1688 3086 1690
rect 3982 1691 3989 1692
rect 2879 1687 2880 1688
rect 2874 1686 2880 1687
rect 3982 1687 3983 1691
rect 3988 1687 3989 1691
rect 3982 1686 3989 1687
rect 4015 1691 4021 1692
rect 4015 1687 4016 1691
rect 4020 1690 4021 1691
rect 4175 1691 4181 1692
rect 4175 1690 4176 1691
rect 4020 1688 4176 1690
rect 4020 1687 4021 1688
rect 4015 1686 4021 1687
rect 4175 1687 4176 1688
rect 4180 1687 4181 1691
rect 4175 1686 4181 1687
rect 4399 1691 4405 1692
rect 4399 1687 4400 1691
rect 4404 1690 4405 1691
rect 4434 1691 4440 1692
rect 4434 1690 4435 1691
rect 4404 1688 4435 1690
rect 4404 1687 4405 1688
rect 4399 1686 4405 1687
rect 4434 1687 4435 1688
rect 4439 1687 4440 1691
rect 4434 1686 4440 1687
rect 4631 1691 4640 1692
rect 4631 1687 4632 1691
rect 4639 1687 4640 1691
rect 4631 1686 4640 1687
rect 4870 1691 4877 1692
rect 4870 1687 4871 1691
rect 4876 1687 4877 1691
rect 5119 1691 5125 1692
rect 5119 1690 5120 1691
rect 4870 1686 4877 1687
rect 4880 1688 5120 1690
rect 4370 1683 4376 1684
rect 4370 1679 4371 1683
rect 4375 1682 4376 1683
rect 4880 1682 4882 1688
rect 5119 1687 5120 1688
rect 5124 1687 5125 1691
rect 5119 1686 5125 1687
rect 5239 1691 5245 1692
rect 5239 1687 5240 1691
rect 5244 1690 5245 1691
rect 5375 1691 5381 1692
rect 5375 1690 5376 1691
rect 5244 1688 5376 1690
rect 5244 1687 5245 1688
rect 5239 1686 5245 1687
rect 5375 1687 5376 1688
rect 5380 1687 5381 1691
rect 5375 1686 5381 1687
rect 5554 1691 5560 1692
rect 5554 1687 5555 1691
rect 5559 1690 5560 1691
rect 5631 1691 5637 1692
rect 5631 1690 5632 1691
rect 5559 1688 5632 1690
rect 5559 1687 5560 1688
rect 5554 1686 5560 1687
rect 5631 1687 5632 1688
rect 5636 1687 5637 1691
rect 5631 1686 5637 1687
rect 4375 1680 4882 1682
rect 4375 1679 4376 1680
rect 4370 1678 4376 1679
rect 238 1667 244 1668
rect 238 1666 239 1667
rect 229 1664 239 1666
rect 238 1663 239 1664
rect 243 1663 244 1667
rect 238 1662 244 1663
rect 490 1667 496 1668
rect 490 1663 491 1667
rect 495 1663 496 1667
rect 1286 1667 1292 1668
rect 490 1662 496 1663
rect 690 1663 696 1664
rect 690 1659 691 1663
rect 695 1659 696 1663
rect 690 1658 696 1659
rect 1074 1663 1080 1664
rect 1074 1659 1075 1663
rect 1079 1659 1080 1663
rect 1286 1663 1287 1667
rect 1291 1663 1292 1667
rect 1286 1662 1292 1663
rect 1074 1658 1080 1659
rect 2090 1659 2096 1660
rect 2090 1655 2091 1659
rect 2095 1655 2096 1659
rect 2090 1654 2096 1655
rect 2122 1659 2128 1660
rect 2122 1655 2123 1659
rect 2127 1658 2128 1659
rect 2258 1659 2264 1660
rect 2127 1656 2137 1658
rect 2127 1655 2128 1656
rect 2122 1654 2128 1655
rect 2258 1655 2259 1659
rect 2263 1658 2264 1659
rect 2602 1659 2608 1660
rect 2602 1658 2603 1659
rect 2263 1656 2289 1658
rect 2541 1656 2603 1658
rect 2263 1655 2264 1656
rect 2258 1654 2264 1655
rect 2602 1655 2603 1656
rect 2607 1655 2608 1659
rect 2602 1654 2608 1655
rect 2706 1659 2712 1660
rect 2706 1655 2707 1659
rect 2711 1655 2712 1659
rect 2706 1654 2712 1655
rect 2874 1659 2880 1660
rect 2874 1655 2875 1659
rect 2879 1655 2880 1659
rect 2874 1654 2880 1655
rect 3030 1659 3036 1660
rect 3030 1655 3031 1659
rect 3035 1655 3036 1659
rect 3030 1654 3036 1655
rect 3074 1659 3080 1660
rect 3074 1655 3075 1659
rect 3079 1658 3080 1659
rect 3079 1656 3129 1658
rect 3079 1655 3080 1656
rect 3074 1654 3080 1655
rect 4015 1651 4021 1652
rect 4015 1650 4016 1651
rect 3957 1648 4016 1650
rect 4015 1647 4016 1648
rect 4020 1647 4021 1651
rect 4015 1646 4021 1647
rect 4146 1651 4152 1652
rect 4146 1647 4147 1651
rect 4151 1647 4152 1651
rect 4146 1646 4152 1647
rect 4370 1651 4376 1652
rect 4370 1647 4371 1651
rect 4375 1647 4376 1651
rect 4370 1646 4376 1647
rect 4434 1651 4440 1652
rect 4434 1647 4435 1651
rect 4439 1650 4440 1651
rect 4634 1651 4640 1652
rect 4439 1648 4513 1650
rect 4439 1647 4440 1648
rect 4434 1646 4440 1647
rect 4634 1647 4635 1651
rect 4639 1650 4640 1651
rect 5086 1651 5092 1652
rect 4639 1648 4753 1650
rect 4639 1647 4640 1648
rect 4634 1646 4640 1647
rect 5086 1647 5087 1651
rect 5091 1647 5092 1651
rect 5086 1646 5092 1647
rect 5346 1651 5352 1652
rect 5346 1647 5347 1651
rect 5351 1647 5352 1651
rect 5346 1646 5352 1647
rect 5498 1651 5504 1652
rect 5498 1647 5499 1651
rect 5503 1650 5504 1651
rect 5503 1648 5513 1650
rect 5503 1647 5504 1648
rect 5498 1646 5504 1647
rect 1074 1635 1080 1636
rect 1074 1631 1075 1635
rect 1079 1634 1080 1635
rect 1079 1632 1282 1634
rect 1079 1631 1080 1632
rect 1074 1630 1080 1631
rect 226 1623 232 1624
rect 226 1619 227 1623
rect 231 1622 232 1623
rect 255 1623 261 1624
rect 255 1622 256 1623
rect 231 1620 256 1622
rect 231 1619 232 1620
rect 226 1618 232 1619
rect 255 1619 256 1620
rect 260 1619 261 1623
rect 255 1618 261 1619
rect 519 1623 525 1624
rect 519 1619 520 1623
rect 524 1622 525 1623
rect 690 1623 696 1624
rect 690 1622 691 1623
rect 524 1620 691 1622
rect 524 1619 525 1620
rect 519 1618 525 1619
rect 690 1619 691 1620
rect 695 1619 696 1623
rect 690 1618 696 1619
rect 807 1623 813 1624
rect 807 1619 808 1623
rect 812 1622 813 1623
rect 986 1623 992 1624
rect 986 1622 987 1623
rect 812 1620 987 1622
rect 812 1619 813 1620
rect 807 1618 813 1619
rect 986 1619 987 1620
rect 991 1619 992 1623
rect 986 1618 992 1619
rect 994 1623 1000 1624
rect 994 1619 995 1623
rect 999 1622 1000 1623
rect 1103 1623 1109 1624
rect 1103 1622 1104 1623
rect 999 1620 1104 1622
rect 999 1619 1000 1620
rect 994 1618 1000 1619
rect 1103 1619 1104 1620
rect 1108 1619 1109 1623
rect 1280 1622 1282 1632
rect 1399 1623 1405 1624
rect 1399 1622 1400 1623
rect 1280 1620 1400 1622
rect 1103 1618 1109 1619
rect 1399 1619 1400 1620
rect 1404 1619 1405 1623
rect 1399 1618 1405 1619
rect 2914 1619 2920 1620
rect 110 1616 116 1617
rect 1934 1616 1940 1617
rect 110 1612 111 1616
rect 115 1612 116 1616
rect 110 1611 116 1612
rect 130 1615 136 1616
rect 130 1611 131 1615
rect 135 1611 136 1615
rect 130 1610 136 1611
rect 394 1615 400 1616
rect 394 1611 395 1615
rect 399 1611 400 1615
rect 394 1610 400 1611
rect 682 1615 688 1616
rect 682 1611 683 1615
rect 687 1611 688 1615
rect 682 1610 688 1611
rect 978 1615 984 1616
rect 978 1611 979 1615
rect 983 1611 984 1615
rect 978 1610 984 1611
rect 1274 1615 1280 1616
rect 1274 1611 1275 1615
rect 1279 1611 1280 1615
rect 1934 1612 1935 1616
rect 1939 1612 1940 1616
rect 1934 1611 1940 1612
rect 2186 1615 2192 1616
rect 2186 1611 2187 1615
rect 2191 1611 2192 1615
rect 1274 1610 1280 1611
rect 2186 1610 2192 1611
rect 2234 1615 2240 1616
rect 2234 1611 2235 1615
rect 2239 1611 2240 1615
rect 2234 1610 2240 1611
rect 2370 1615 2376 1616
rect 2370 1611 2371 1615
rect 2375 1611 2376 1615
rect 2370 1610 2376 1611
rect 2506 1615 2512 1616
rect 2506 1611 2507 1615
rect 2511 1611 2512 1615
rect 2506 1610 2512 1611
rect 2642 1615 2648 1616
rect 2642 1611 2643 1615
rect 2647 1611 2648 1615
rect 2642 1610 2648 1611
rect 2778 1615 2784 1616
rect 2778 1611 2779 1615
rect 2783 1611 2784 1615
rect 2914 1615 2915 1619
rect 2919 1615 2920 1619
rect 4398 1619 4404 1620
rect 2914 1614 2920 1615
rect 3050 1615 3056 1616
rect 2778 1610 2784 1611
rect 3050 1611 3051 1615
rect 3055 1611 3056 1615
rect 3050 1610 3056 1611
rect 3186 1615 3192 1616
rect 3186 1611 3187 1615
rect 3191 1611 3192 1615
rect 3186 1610 3192 1611
rect 3954 1615 3960 1616
rect 3954 1611 3955 1615
rect 3959 1611 3960 1615
rect 3954 1610 3960 1611
rect 4002 1615 4008 1616
rect 4002 1611 4003 1615
rect 4007 1611 4008 1615
rect 4002 1610 4008 1611
rect 4250 1615 4256 1616
rect 4250 1611 4251 1615
rect 4255 1611 4256 1615
rect 4398 1615 4399 1619
rect 4403 1615 4404 1619
rect 4870 1619 4876 1620
rect 4398 1614 4404 1615
rect 4682 1615 4688 1616
rect 4250 1610 4256 1611
rect 4682 1611 4683 1615
rect 4687 1611 4688 1615
rect 4870 1615 4871 1619
rect 4875 1615 4876 1619
rect 5466 1619 5472 1620
rect 4870 1614 4876 1615
rect 5138 1615 5144 1616
rect 4682 1610 4688 1611
rect 5138 1611 5139 1615
rect 5143 1611 5144 1615
rect 5466 1615 5467 1619
rect 5471 1615 5472 1619
rect 5466 1614 5472 1615
rect 5138 1610 5144 1611
rect 158 1600 164 1601
rect 110 1599 116 1600
rect 110 1595 111 1599
rect 115 1595 116 1599
rect 158 1596 159 1600
rect 163 1596 164 1600
rect 158 1595 164 1596
rect 422 1600 428 1601
rect 422 1596 423 1600
rect 427 1596 428 1600
rect 422 1595 428 1596
rect 710 1600 716 1601
rect 710 1596 711 1600
rect 715 1596 716 1600
rect 710 1595 716 1596
rect 1006 1600 1012 1601
rect 1006 1596 1007 1600
rect 1011 1596 1012 1600
rect 1006 1595 1012 1596
rect 1302 1600 1308 1601
rect 1302 1596 1303 1600
rect 1307 1596 1308 1600
rect 1302 1595 1308 1596
rect 1934 1599 1940 1600
rect 1934 1595 1935 1599
rect 1939 1595 1940 1599
rect 110 1594 116 1595
rect 1934 1594 1940 1595
rect 2706 1583 2712 1584
rect 2706 1579 2707 1583
rect 2711 1582 2712 1583
rect 3954 1583 3960 1584
rect 2711 1580 2842 1582
rect 2711 1579 2712 1580
rect 2706 1578 2712 1579
rect 2215 1575 2221 1576
rect 2215 1571 2216 1575
rect 2220 1574 2221 1575
rect 2234 1575 2240 1576
rect 2234 1574 2235 1575
rect 2220 1572 2235 1574
rect 2220 1571 2221 1572
rect 2215 1570 2221 1571
rect 2234 1571 2235 1572
rect 2239 1571 2240 1575
rect 2234 1570 2240 1571
rect 2351 1575 2357 1576
rect 2351 1571 2352 1575
rect 2356 1574 2357 1575
rect 2370 1575 2376 1576
rect 2370 1574 2371 1575
rect 2356 1572 2371 1574
rect 2356 1571 2357 1572
rect 2351 1570 2357 1571
rect 2370 1571 2371 1572
rect 2375 1571 2376 1575
rect 2370 1570 2376 1571
rect 2487 1575 2493 1576
rect 2487 1571 2488 1575
rect 2492 1574 2493 1575
rect 2506 1575 2512 1576
rect 2506 1574 2507 1575
rect 2492 1572 2507 1574
rect 2492 1571 2493 1572
rect 2487 1570 2493 1571
rect 2506 1571 2507 1572
rect 2511 1571 2512 1575
rect 2506 1570 2512 1571
rect 2623 1575 2629 1576
rect 2623 1571 2624 1575
rect 2628 1574 2629 1575
rect 2642 1575 2648 1576
rect 2642 1574 2643 1575
rect 2628 1572 2643 1574
rect 2628 1571 2629 1572
rect 2623 1570 2629 1571
rect 2642 1571 2643 1572
rect 2647 1571 2648 1575
rect 2642 1570 2648 1571
rect 2759 1575 2765 1576
rect 2759 1571 2760 1575
rect 2764 1574 2765 1575
rect 2778 1575 2784 1576
rect 2778 1574 2779 1575
rect 2764 1572 2779 1574
rect 2764 1571 2765 1572
rect 2759 1570 2765 1571
rect 2778 1571 2779 1572
rect 2783 1571 2784 1575
rect 2840 1574 2842 1580
rect 3954 1579 3955 1583
rect 3959 1582 3960 1583
rect 4682 1583 4688 1584
rect 3959 1580 4590 1582
rect 3959 1579 3960 1580
rect 3954 1578 3960 1579
rect 2895 1575 2901 1576
rect 2895 1574 2896 1575
rect 2840 1572 2896 1574
rect 2778 1570 2784 1571
rect 2895 1571 2896 1572
rect 2900 1571 2901 1575
rect 2895 1570 2901 1571
rect 3031 1575 3037 1576
rect 3031 1571 3032 1575
rect 3036 1574 3037 1575
rect 3050 1575 3056 1576
rect 3050 1574 3051 1575
rect 3036 1572 3051 1574
rect 3036 1571 3037 1572
rect 3031 1570 3037 1571
rect 3050 1571 3051 1572
rect 3055 1571 3056 1575
rect 3050 1570 3056 1571
rect 3167 1575 3173 1576
rect 3167 1571 3168 1575
rect 3172 1574 3173 1575
rect 3186 1575 3192 1576
rect 3186 1574 3187 1575
rect 3172 1572 3187 1574
rect 3172 1571 3173 1572
rect 3167 1570 3173 1571
rect 3186 1571 3187 1572
rect 3191 1571 3192 1575
rect 3186 1570 3192 1571
rect 3298 1575 3309 1576
rect 3298 1571 3299 1575
rect 3303 1571 3304 1575
rect 3308 1571 3309 1575
rect 3298 1570 3309 1571
rect 3983 1575 3989 1576
rect 3983 1571 3984 1575
rect 3988 1574 3989 1575
rect 4002 1575 4008 1576
rect 4002 1574 4003 1575
rect 3988 1572 4003 1574
rect 3988 1571 3989 1572
rect 3983 1570 3989 1571
rect 4002 1571 4003 1572
rect 4007 1571 4008 1575
rect 4002 1570 4008 1571
rect 4119 1575 4128 1576
rect 4119 1571 4120 1575
rect 4127 1571 4128 1575
rect 4119 1570 4128 1571
rect 4146 1575 4152 1576
rect 4146 1571 4147 1575
rect 4151 1574 4152 1575
rect 4279 1575 4285 1576
rect 4279 1574 4280 1575
rect 4151 1572 4280 1574
rect 4151 1571 4152 1572
rect 4146 1570 4152 1571
rect 4279 1571 4280 1572
rect 4284 1571 4285 1575
rect 4279 1570 4285 1571
rect 4478 1575 4485 1576
rect 4478 1571 4479 1575
rect 4484 1571 4485 1575
rect 4588 1574 4590 1580
rect 4682 1579 4683 1583
rect 4687 1582 4688 1583
rect 4687 1580 5150 1582
rect 4687 1579 4688 1580
rect 4682 1578 4688 1579
rect 4711 1575 4717 1576
rect 4711 1574 4712 1575
rect 4588 1572 4712 1574
rect 4478 1570 4485 1571
rect 4711 1571 4712 1572
rect 4716 1571 4717 1575
rect 4711 1570 4717 1571
rect 4975 1575 4981 1576
rect 4975 1571 4976 1575
rect 4980 1574 4981 1575
rect 5138 1575 5144 1576
rect 5138 1574 5139 1575
rect 4980 1572 5139 1574
rect 4980 1571 4981 1572
rect 4975 1570 4981 1571
rect 5138 1571 5139 1572
rect 5143 1571 5144 1575
rect 5148 1574 5150 1580
rect 5255 1575 5261 1576
rect 5255 1574 5256 1575
rect 5148 1572 5256 1574
rect 5138 1570 5144 1571
rect 5255 1571 5256 1572
rect 5260 1571 5261 1575
rect 5255 1570 5261 1571
rect 5346 1575 5352 1576
rect 5346 1571 5347 1575
rect 5351 1574 5352 1575
rect 5543 1575 5549 1576
rect 5543 1574 5544 1575
rect 5351 1572 5544 1574
rect 5351 1571 5352 1572
rect 5346 1570 5352 1571
rect 5543 1571 5544 1572
rect 5548 1571 5549 1575
rect 5543 1570 5549 1571
rect 1974 1568 1980 1569
rect 3798 1568 3804 1569
rect 1974 1564 1975 1568
rect 1979 1564 1980 1568
rect 1974 1563 1980 1564
rect 2090 1567 2096 1568
rect 2090 1563 2091 1567
rect 2095 1563 2096 1567
rect 2090 1562 2096 1563
rect 2226 1567 2232 1568
rect 2226 1563 2227 1567
rect 2231 1563 2232 1567
rect 2226 1562 2232 1563
rect 2362 1567 2368 1568
rect 2362 1563 2363 1567
rect 2367 1563 2368 1567
rect 2362 1562 2368 1563
rect 2498 1567 2504 1568
rect 2498 1563 2499 1567
rect 2503 1563 2504 1567
rect 2498 1562 2504 1563
rect 2634 1567 2640 1568
rect 2634 1563 2635 1567
rect 2639 1563 2640 1567
rect 2634 1562 2640 1563
rect 2770 1567 2776 1568
rect 2770 1563 2771 1567
rect 2775 1563 2776 1567
rect 2770 1562 2776 1563
rect 2906 1567 2912 1568
rect 2906 1563 2907 1567
rect 2911 1563 2912 1567
rect 2906 1562 2912 1563
rect 3042 1567 3048 1568
rect 3042 1563 3043 1567
rect 3047 1563 3048 1567
rect 3042 1562 3048 1563
rect 3178 1567 3184 1568
rect 3178 1563 3179 1567
rect 3183 1563 3184 1567
rect 3798 1564 3799 1568
rect 3803 1564 3804 1568
rect 3798 1563 3804 1564
rect 3838 1568 3844 1569
rect 5662 1568 5668 1569
rect 3838 1564 3839 1568
rect 3843 1564 3844 1568
rect 3838 1563 3844 1564
rect 3858 1567 3864 1568
rect 3858 1563 3859 1567
rect 3863 1563 3864 1567
rect 3178 1562 3184 1563
rect 3858 1562 3864 1563
rect 3994 1567 4000 1568
rect 3994 1563 3995 1567
rect 3999 1563 4000 1567
rect 3994 1562 4000 1563
rect 4154 1567 4160 1568
rect 4154 1563 4155 1567
rect 4159 1563 4160 1567
rect 4154 1562 4160 1563
rect 4354 1567 4360 1568
rect 4354 1563 4355 1567
rect 4359 1563 4360 1567
rect 4354 1562 4360 1563
rect 4586 1567 4592 1568
rect 4586 1563 4587 1567
rect 4591 1563 4592 1567
rect 4586 1562 4592 1563
rect 4850 1567 4856 1568
rect 4850 1563 4851 1567
rect 4855 1563 4856 1567
rect 4850 1562 4856 1563
rect 5130 1567 5136 1568
rect 5130 1563 5131 1567
rect 5135 1563 5136 1567
rect 5130 1562 5136 1563
rect 5418 1567 5424 1568
rect 5418 1563 5419 1567
rect 5423 1563 5424 1567
rect 5662 1564 5663 1568
rect 5667 1564 5668 1568
rect 5662 1563 5668 1564
rect 5418 1562 5424 1563
rect 2118 1552 2124 1553
rect 1974 1551 1980 1552
rect 1974 1547 1975 1551
rect 1979 1547 1980 1551
rect 2118 1548 2119 1552
rect 2123 1548 2124 1552
rect 2118 1547 2124 1548
rect 2254 1552 2260 1553
rect 2254 1548 2255 1552
rect 2259 1548 2260 1552
rect 2254 1547 2260 1548
rect 2390 1552 2396 1553
rect 2390 1548 2391 1552
rect 2395 1548 2396 1552
rect 2390 1547 2396 1548
rect 2526 1552 2532 1553
rect 2526 1548 2527 1552
rect 2531 1548 2532 1552
rect 2526 1547 2532 1548
rect 2662 1552 2668 1553
rect 2662 1548 2663 1552
rect 2667 1548 2668 1552
rect 2662 1547 2668 1548
rect 2798 1552 2804 1553
rect 2798 1548 2799 1552
rect 2803 1548 2804 1552
rect 2798 1547 2804 1548
rect 2934 1552 2940 1553
rect 2934 1548 2935 1552
rect 2939 1548 2940 1552
rect 2934 1547 2940 1548
rect 3070 1552 3076 1553
rect 3070 1548 3071 1552
rect 3075 1548 3076 1552
rect 3070 1547 3076 1548
rect 3206 1552 3212 1553
rect 3886 1552 3892 1553
rect 3206 1548 3207 1552
rect 3211 1548 3212 1552
rect 3206 1547 3212 1548
rect 3798 1551 3804 1552
rect 3798 1547 3799 1551
rect 3803 1547 3804 1551
rect 1974 1546 1980 1547
rect 3798 1546 3804 1547
rect 3838 1551 3844 1552
rect 3838 1547 3839 1551
rect 3843 1547 3844 1551
rect 3886 1548 3887 1552
rect 3891 1548 3892 1552
rect 3886 1547 3892 1548
rect 4022 1552 4028 1553
rect 4022 1548 4023 1552
rect 4027 1548 4028 1552
rect 4022 1547 4028 1548
rect 4182 1552 4188 1553
rect 4182 1548 4183 1552
rect 4187 1548 4188 1552
rect 4182 1547 4188 1548
rect 4382 1552 4388 1553
rect 4382 1548 4383 1552
rect 4387 1548 4388 1552
rect 4382 1547 4388 1548
rect 4614 1552 4620 1553
rect 4614 1548 4615 1552
rect 4619 1548 4620 1552
rect 4614 1547 4620 1548
rect 4878 1552 4884 1553
rect 4878 1548 4879 1552
rect 4883 1548 4884 1552
rect 4878 1547 4884 1548
rect 5158 1552 5164 1553
rect 5158 1548 5159 1552
rect 5163 1548 5164 1552
rect 5158 1547 5164 1548
rect 5446 1552 5452 1553
rect 5446 1548 5447 1552
rect 5451 1548 5452 1552
rect 5446 1547 5452 1548
rect 5662 1551 5668 1552
rect 5662 1547 5663 1551
rect 5667 1547 5668 1551
rect 3838 1546 3844 1547
rect 5662 1546 5668 1547
rect 110 1529 116 1530
rect 1934 1529 1940 1530
rect 110 1525 111 1529
rect 115 1525 116 1529
rect 110 1524 116 1525
rect 158 1528 164 1529
rect 158 1524 159 1528
rect 163 1524 164 1528
rect 158 1523 164 1524
rect 374 1528 380 1529
rect 374 1524 375 1528
rect 379 1524 380 1528
rect 374 1523 380 1524
rect 606 1528 612 1529
rect 606 1524 607 1528
rect 611 1524 612 1528
rect 606 1523 612 1524
rect 838 1528 844 1529
rect 838 1524 839 1528
rect 843 1524 844 1528
rect 838 1523 844 1524
rect 1070 1528 1076 1529
rect 1070 1524 1071 1528
rect 1075 1524 1076 1528
rect 1070 1523 1076 1524
rect 1302 1528 1308 1529
rect 1302 1524 1303 1528
rect 1307 1524 1308 1528
rect 1934 1525 1935 1529
rect 1939 1525 1940 1529
rect 1934 1524 1940 1525
rect 1302 1523 1308 1524
rect 130 1513 136 1514
rect 110 1512 116 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 130 1509 131 1513
rect 135 1509 136 1513
rect 130 1508 136 1509
rect 346 1513 352 1514
rect 346 1509 347 1513
rect 351 1509 352 1513
rect 346 1508 352 1509
rect 578 1513 584 1514
rect 578 1509 579 1513
rect 583 1509 584 1513
rect 578 1508 584 1509
rect 810 1513 816 1514
rect 810 1509 811 1513
rect 815 1509 816 1513
rect 810 1508 816 1509
rect 1042 1513 1048 1514
rect 1042 1509 1043 1513
rect 1047 1509 1048 1513
rect 1042 1508 1048 1509
rect 1274 1513 1280 1514
rect 1274 1509 1275 1513
rect 1279 1509 1280 1513
rect 1274 1508 1280 1509
rect 1934 1512 1940 1513
rect 1934 1508 1935 1512
rect 1939 1508 1940 1512
rect 110 1507 116 1508
rect 1934 1507 1940 1508
rect 2186 1511 2192 1512
rect 2186 1507 2187 1511
rect 2191 1510 2192 1511
rect 2654 1511 2660 1512
rect 2654 1510 2655 1511
rect 2191 1508 2655 1510
rect 2191 1507 2192 1508
rect 2186 1506 2192 1507
rect 2654 1507 2655 1508
rect 2659 1507 2660 1511
rect 2654 1506 2660 1507
rect 4122 1507 4128 1508
rect 238 1503 244 1504
rect 238 1499 239 1503
rect 243 1502 244 1503
rect 255 1503 261 1504
rect 255 1502 256 1503
rect 243 1500 256 1502
rect 243 1499 244 1500
rect 238 1498 244 1499
rect 255 1499 256 1500
rect 260 1499 261 1503
rect 255 1498 261 1499
rect 354 1503 360 1504
rect 354 1499 355 1503
rect 359 1502 360 1503
rect 471 1503 477 1504
rect 471 1502 472 1503
rect 359 1500 472 1502
rect 359 1499 360 1500
rect 354 1498 360 1499
rect 471 1499 472 1500
rect 476 1499 477 1503
rect 471 1498 477 1499
rect 703 1503 709 1504
rect 703 1499 704 1503
rect 708 1502 709 1503
rect 718 1503 724 1504
rect 718 1502 719 1503
rect 708 1500 719 1502
rect 708 1499 709 1500
rect 703 1498 709 1499
rect 718 1499 719 1500
rect 723 1499 724 1503
rect 718 1498 724 1499
rect 802 1503 808 1504
rect 802 1499 803 1503
rect 807 1502 808 1503
rect 935 1503 941 1504
rect 935 1502 936 1503
rect 807 1500 936 1502
rect 807 1499 808 1500
rect 802 1498 808 1499
rect 935 1499 936 1500
rect 940 1499 941 1503
rect 935 1498 941 1499
rect 1167 1503 1176 1504
rect 1167 1499 1168 1503
rect 1175 1499 1176 1503
rect 1167 1498 1176 1499
rect 1399 1503 1408 1504
rect 1399 1499 1400 1503
rect 1407 1499 1408 1503
rect 4122 1503 4123 1507
rect 4127 1506 4128 1507
rect 4258 1507 4264 1508
rect 4258 1506 4259 1507
rect 4127 1504 4259 1506
rect 4127 1503 4128 1504
rect 4122 1502 4128 1503
rect 4258 1503 4259 1504
rect 4263 1503 4264 1507
rect 4258 1502 4264 1503
rect 1399 1498 1408 1499
rect 3838 1493 3844 1494
rect 5662 1493 5668 1494
rect 3838 1489 3839 1493
rect 3843 1489 3844 1493
rect 3838 1488 3844 1489
rect 3886 1492 3892 1493
rect 3886 1488 3887 1492
rect 3891 1488 3892 1492
rect 3886 1487 3892 1488
rect 4022 1492 4028 1493
rect 4022 1488 4023 1492
rect 4027 1488 4028 1492
rect 4022 1487 4028 1488
rect 4158 1492 4164 1493
rect 4158 1488 4159 1492
rect 4163 1488 4164 1492
rect 4158 1487 4164 1488
rect 4302 1492 4308 1493
rect 4302 1488 4303 1492
rect 4307 1488 4308 1492
rect 4302 1487 4308 1488
rect 4494 1492 4500 1493
rect 4494 1488 4495 1492
rect 4499 1488 4500 1492
rect 4494 1487 4500 1488
rect 4718 1492 4724 1493
rect 4718 1488 4719 1492
rect 4723 1488 4724 1492
rect 4718 1487 4724 1488
rect 4966 1492 4972 1493
rect 4966 1488 4967 1492
rect 4971 1488 4972 1492
rect 4966 1487 4972 1488
rect 5222 1492 5228 1493
rect 5222 1488 5223 1492
rect 5227 1488 5228 1492
rect 5222 1487 5228 1488
rect 5486 1492 5492 1493
rect 5486 1488 5487 1492
rect 5491 1488 5492 1492
rect 5662 1489 5663 1493
rect 5667 1489 5668 1493
rect 5662 1488 5668 1489
rect 5486 1487 5492 1488
rect 3858 1477 3864 1478
rect 3838 1476 3844 1477
rect 1974 1473 1980 1474
rect 3798 1473 3804 1474
rect 354 1471 360 1472
rect 354 1470 355 1471
rect 228 1468 355 1470
rect 228 1461 230 1468
rect 354 1467 355 1468
rect 359 1467 360 1471
rect 994 1471 1000 1472
rect 994 1470 995 1471
rect 354 1466 360 1467
rect 908 1468 995 1470
rect 303 1463 309 1464
rect 303 1459 304 1463
rect 308 1462 309 1463
rect 802 1463 808 1464
rect 802 1462 803 1463
rect 308 1460 353 1462
rect 677 1460 803 1462
rect 308 1459 309 1460
rect 303 1458 309 1459
rect 802 1459 803 1460
rect 807 1459 808 1463
rect 908 1461 910 1468
rect 994 1467 995 1468
rect 999 1467 1000 1471
rect 1974 1469 1975 1473
rect 1979 1469 1980 1473
rect 1974 1468 1980 1469
rect 2022 1472 2028 1473
rect 2022 1468 2023 1472
rect 2027 1468 2028 1472
rect 2022 1467 2028 1468
rect 2158 1472 2164 1473
rect 2158 1468 2159 1472
rect 2163 1468 2164 1472
rect 2158 1467 2164 1468
rect 2294 1472 2300 1473
rect 2294 1468 2295 1472
rect 2299 1468 2300 1472
rect 2294 1467 2300 1468
rect 2430 1472 2436 1473
rect 2430 1468 2431 1472
rect 2435 1468 2436 1472
rect 2430 1467 2436 1468
rect 2566 1472 2572 1473
rect 2566 1468 2567 1472
rect 2571 1468 2572 1472
rect 2566 1467 2572 1468
rect 2702 1472 2708 1473
rect 2702 1468 2703 1472
rect 2707 1468 2708 1472
rect 2702 1467 2708 1468
rect 2838 1472 2844 1473
rect 2838 1468 2839 1472
rect 2843 1468 2844 1472
rect 2838 1467 2844 1468
rect 2974 1472 2980 1473
rect 2974 1468 2975 1472
rect 2979 1468 2980 1472
rect 3798 1469 3799 1473
rect 3803 1469 3804 1473
rect 3838 1472 3839 1476
rect 3843 1472 3844 1476
rect 3858 1473 3859 1477
rect 3863 1473 3864 1477
rect 3858 1472 3864 1473
rect 3994 1477 4000 1478
rect 3994 1473 3995 1477
rect 3999 1473 4000 1477
rect 3994 1472 4000 1473
rect 4130 1477 4136 1478
rect 4130 1473 4131 1477
rect 4135 1473 4136 1477
rect 4130 1472 4136 1473
rect 4274 1477 4280 1478
rect 4274 1473 4275 1477
rect 4279 1473 4280 1477
rect 4274 1472 4280 1473
rect 4466 1477 4472 1478
rect 4466 1473 4467 1477
rect 4471 1473 4472 1477
rect 4466 1472 4472 1473
rect 4690 1477 4696 1478
rect 4690 1473 4691 1477
rect 4695 1473 4696 1477
rect 4690 1472 4696 1473
rect 4938 1477 4944 1478
rect 4938 1473 4939 1477
rect 4943 1473 4944 1477
rect 4938 1472 4944 1473
rect 5194 1477 5200 1478
rect 5194 1473 5195 1477
rect 5199 1473 5200 1477
rect 5194 1472 5200 1473
rect 5458 1477 5464 1478
rect 5458 1473 5459 1477
rect 5463 1473 5464 1477
rect 5458 1472 5464 1473
rect 5662 1476 5668 1477
rect 5662 1472 5663 1476
rect 5667 1472 5668 1476
rect 3838 1471 3844 1472
rect 5662 1471 5668 1472
rect 3798 1468 3804 1469
rect 2974 1467 2980 1468
rect 3983 1467 3992 1468
rect 994 1466 1000 1467
rect 986 1463 992 1464
rect 802 1458 808 1459
rect 986 1459 987 1463
rect 991 1462 992 1463
rect 1170 1463 1176 1464
rect 991 1460 1049 1462
rect 991 1459 992 1460
rect 986 1458 992 1459
rect 1170 1459 1171 1463
rect 1175 1462 1176 1463
rect 3983 1463 3984 1467
rect 3991 1463 3992 1467
rect 3983 1462 3992 1463
rect 4119 1467 4128 1468
rect 4119 1463 4120 1467
rect 4127 1463 4128 1467
rect 4119 1462 4128 1463
rect 4250 1467 4261 1468
rect 4250 1463 4251 1467
rect 4255 1463 4256 1467
rect 4260 1463 4261 1467
rect 4250 1462 4261 1463
rect 4398 1467 4405 1468
rect 4398 1463 4399 1467
rect 4404 1463 4405 1467
rect 4398 1462 4405 1463
rect 4591 1467 4600 1468
rect 4591 1463 4592 1467
rect 4599 1463 4600 1467
rect 4591 1462 4600 1463
rect 4815 1467 4824 1468
rect 4815 1463 4816 1467
rect 4823 1463 4824 1467
rect 4815 1462 4824 1463
rect 5063 1467 5072 1468
rect 5063 1463 5064 1467
rect 5071 1463 5072 1467
rect 5319 1467 5325 1468
rect 5319 1466 5320 1467
rect 5063 1462 5072 1463
rect 5299 1464 5320 1466
rect 1175 1460 1281 1462
rect 1175 1459 1176 1460
rect 1170 1458 1176 1459
rect 4154 1459 4160 1460
rect 1994 1457 2000 1458
rect 1974 1456 1980 1457
rect 1974 1452 1975 1456
rect 1979 1452 1980 1456
rect 1994 1453 1995 1457
rect 1999 1453 2000 1457
rect 1994 1452 2000 1453
rect 2130 1457 2136 1458
rect 2130 1453 2131 1457
rect 2135 1453 2136 1457
rect 2130 1452 2136 1453
rect 2266 1457 2272 1458
rect 2266 1453 2267 1457
rect 2271 1453 2272 1457
rect 2266 1452 2272 1453
rect 2402 1457 2408 1458
rect 2402 1453 2403 1457
rect 2407 1453 2408 1457
rect 2402 1452 2408 1453
rect 2538 1457 2544 1458
rect 2538 1453 2539 1457
rect 2543 1453 2544 1457
rect 2538 1452 2544 1453
rect 2674 1457 2680 1458
rect 2674 1453 2675 1457
rect 2679 1453 2680 1457
rect 2674 1452 2680 1453
rect 2810 1457 2816 1458
rect 2810 1453 2811 1457
rect 2815 1453 2816 1457
rect 2810 1452 2816 1453
rect 2946 1457 2952 1458
rect 2946 1453 2947 1457
rect 2951 1453 2952 1457
rect 2946 1452 2952 1453
rect 3798 1456 3804 1457
rect 3798 1452 3799 1456
rect 3803 1452 3804 1456
rect 4154 1455 4155 1459
rect 4159 1458 4160 1459
rect 5299 1458 5301 1464
rect 5319 1463 5320 1464
rect 5324 1463 5325 1467
rect 5319 1462 5325 1463
rect 5582 1467 5589 1468
rect 5582 1463 5583 1467
rect 5588 1463 5589 1467
rect 5582 1462 5589 1463
rect 4159 1456 5301 1458
rect 4159 1455 4160 1456
rect 4154 1454 4160 1455
rect 1974 1451 1980 1452
rect 3798 1451 3804 1452
rect 2119 1447 2128 1448
rect 2119 1443 2120 1447
rect 2127 1443 2128 1447
rect 2119 1442 2128 1443
rect 2255 1447 2264 1448
rect 2255 1443 2256 1447
rect 2263 1443 2264 1447
rect 2255 1442 2264 1443
rect 2391 1447 2400 1448
rect 2391 1443 2392 1447
rect 2399 1443 2400 1447
rect 2391 1442 2400 1443
rect 2527 1447 2536 1448
rect 2527 1443 2528 1447
rect 2535 1443 2536 1447
rect 2527 1442 2536 1443
rect 2654 1447 2660 1448
rect 2654 1443 2655 1447
rect 2659 1446 2660 1447
rect 2663 1447 2669 1448
rect 2663 1446 2664 1447
rect 2659 1444 2664 1446
rect 2659 1443 2660 1444
rect 2654 1442 2660 1443
rect 2663 1443 2664 1444
rect 2668 1443 2669 1447
rect 2663 1442 2669 1443
rect 2799 1447 2808 1448
rect 2799 1443 2800 1447
rect 2807 1443 2808 1447
rect 2799 1442 2808 1443
rect 2934 1447 2941 1448
rect 2934 1443 2935 1447
rect 2940 1443 2941 1447
rect 3071 1447 3077 1448
rect 3071 1446 3072 1447
rect 2934 1442 2941 1443
rect 2944 1444 3072 1446
rect 2770 1439 2776 1440
rect 2770 1435 2771 1439
rect 2775 1438 2776 1439
rect 2944 1438 2946 1444
rect 3071 1443 3072 1444
rect 3076 1443 3077 1447
rect 3071 1442 3077 1443
rect 2775 1436 2946 1438
rect 2775 1435 2776 1436
rect 2770 1434 2776 1435
rect 3954 1427 3960 1428
rect 3954 1423 3955 1427
rect 3959 1423 3960 1427
rect 3954 1422 3960 1423
rect 3986 1427 3992 1428
rect 3986 1423 3987 1427
rect 3991 1426 3992 1427
rect 4122 1427 4128 1428
rect 3991 1424 4001 1426
rect 3991 1423 3992 1424
rect 3986 1422 3992 1423
rect 4122 1423 4123 1427
rect 4127 1426 4128 1427
rect 4258 1427 4264 1428
rect 4127 1424 4137 1426
rect 4127 1423 4128 1424
rect 4122 1422 4128 1423
rect 4258 1423 4259 1427
rect 4263 1426 4264 1427
rect 4478 1427 4484 1428
rect 4263 1424 4281 1426
rect 4263 1423 4264 1424
rect 4258 1422 4264 1423
rect 4478 1423 4479 1427
rect 4483 1423 4484 1427
rect 4478 1422 4484 1423
rect 4594 1427 4600 1428
rect 4594 1423 4595 1427
rect 4599 1426 4600 1427
rect 4818 1427 4824 1428
rect 4599 1424 4697 1426
rect 4599 1423 4600 1424
rect 4594 1422 4600 1423
rect 4818 1423 4819 1427
rect 4823 1426 4824 1427
rect 5066 1427 5072 1428
rect 4823 1424 4945 1426
rect 4823 1423 4824 1424
rect 4818 1422 4824 1423
rect 5066 1423 5067 1427
rect 5071 1426 5072 1427
rect 5554 1427 5560 1428
rect 5071 1424 5201 1426
rect 5071 1423 5072 1424
rect 5066 1422 5072 1423
rect 5554 1423 5555 1427
rect 5559 1423 5560 1427
rect 5554 1422 5560 1423
rect 718 1419 724 1420
rect 226 1415 232 1416
rect 226 1411 227 1415
rect 231 1411 232 1415
rect 226 1410 232 1411
rect 506 1415 512 1416
rect 506 1411 507 1415
rect 511 1411 512 1415
rect 718 1415 719 1419
rect 723 1418 724 1419
rect 1402 1419 1408 1420
rect 723 1416 745 1418
rect 723 1415 724 1416
rect 718 1414 724 1415
rect 1186 1415 1192 1416
rect 506 1410 512 1411
rect 1186 1411 1187 1415
rect 1191 1411 1192 1415
rect 1402 1415 1403 1419
rect 1407 1418 1408 1419
rect 1407 1416 1457 1418
rect 1407 1415 1408 1416
rect 1402 1414 1408 1415
rect 1882 1415 1888 1416
rect 1186 1410 1192 1411
rect 1882 1411 1883 1415
rect 1887 1411 1888 1415
rect 1882 1410 1888 1411
rect 2122 1407 2128 1408
rect 2092 1398 2094 1405
rect 2122 1403 2123 1407
rect 2127 1406 2128 1407
rect 2258 1407 2264 1408
rect 2127 1404 2137 1406
rect 2127 1403 2128 1404
rect 2122 1402 2128 1403
rect 2258 1403 2259 1407
rect 2263 1406 2264 1407
rect 2394 1407 2400 1408
rect 2263 1404 2273 1406
rect 2263 1403 2264 1404
rect 2258 1402 2264 1403
rect 2394 1403 2395 1407
rect 2399 1406 2400 1407
rect 2530 1407 2536 1408
rect 2399 1404 2409 1406
rect 2399 1403 2400 1404
rect 2394 1402 2400 1403
rect 2530 1403 2531 1407
rect 2535 1406 2536 1407
rect 2770 1407 2776 1408
rect 2535 1404 2545 1406
rect 2535 1403 2536 1404
rect 2530 1402 2536 1403
rect 2770 1403 2771 1407
rect 2775 1403 2776 1407
rect 2770 1402 2776 1403
rect 2802 1407 2808 1408
rect 2802 1403 2803 1407
rect 2807 1406 2808 1407
rect 3298 1407 3304 1408
rect 3298 1406 3299 1407
rect 2807 1404 2817 1406
rect 3045 1404 3299 1406
rect 2807 1403 2808 1404
rect 2802 1402 2808 1403
rect 3298 1403 3299 1404
rect 3303 1403 3304 1407
rect 3298 1402 3304 1403
rect 2298 1399 2304 1400
rect 2298 1398 2299 1399
rect 2092 1396 2299 1398
rect 506 1395 512 1396
rect 506 1391 507 1395
rect 511 1394 512 1395
rect 862 1395 868 1396
rect 862 1394 863 1395
rect 511 1392 863 1394
rect 511 1391 512 1392
rect 506 1390 512 1391
rect 862 1391 863 1392
rect 867 1391 868 1395
rect 862 1390 868 1391
rect 1186 1395 1192 1396
rect 1186 1391 1187 1395
rect 1191 1394 1192 1395
rect 1574 1395 1580 1396
rect 1574 1394 1575 1395
rect 1191 1392 1575 1394
rect 1191 1391 1192 1392
rect 1186 1390 1192 1391
rect 1574 1391 1575 1392
rect 1579 1391 1580 1395
rect 2298 1395 2299 1396
rect 2303 1395 2304 1399
rect 2298 1394 2304 1395
rect 1574 1390 1580 1391
rect 3778 1391 3784 1392
rect 3778 1387 3779 1391
rect 3783 1390 3784 1391
rect 4154 1391 4160 1392
rect 3783 1388 3865 1390
rect 3783 1387 3784 1388
rect 3778 1386 3784 1387
rect 4154 1387 4155 1391
rect 4159 1387 4160 1391
rect 5582 1391 5588 1392
rect 4154 1386 4160 1387
rect 4314 1387 4320 1388
rect 4314 1383 4315 1387
rect 4319 1383 4320 1387
rect 4314 1382 4320 1383
rect 4586 1387 4592 1388
rect 4586 1383 4587 1387
rect 4591 1383 4592 1387
rect 4586 1382 4592 1383
rect 4882 1387 4888 1388
rect 4882 1383 4883 1387
rect 4887 1383 4888 1387
rect 4882 1382 4888 1383
rect 5194 1387 5200 1388
rect 5194 1383 5195 1387
rect 5199 1383 5200 1387
rect 5582 1387 5583 1391
rect 5587 1387 5588 1391
rect 5582 1386 5588 1387
rect 5194 1382 5200 1383
rect 255 1375 261 1376
rect 255 1371 256 1375
rect 260 1374 261 1375
rect 303 1375 309 1376
rect 303 1374 304 1375
rect 260 1372 304 1374
rect 260 1371 261 1372
rect 255 1370 261 1371
rect 303 1371 304 1372
rect 308 1371 309 1375
rect 303 1370 309 1371
rect 535 1375 541 1376
rect 535 1371 536 1375
rect 540 1374 541 1375
rect 543 1375 549 1376
rect 543 1374 544 1375
rect 540 1372 544 1374
rect 540 1371 541 1372
rect 535 1370 541 1371
rect 543 1371 544 1372
rect 548 1371 549 1375
rect 543 1370 549 1371
rect 862 1375 869 1376
rect 862 1371 863 1375
rect 868 1371 869 1375
rect 862 1370 869 1371
rect 1034 1375 1040 1376
rect 1034 1371 1035 1375
rect 1039 1374 1040 1375
rect 1215 1375 1221 1376
rect 1215 1374 1216 1375
rect 1039 1372 1216 1374
rect 1039 1371 1040 1372
rect 1034 1370 1040 1371
rect 1215 1371 1216 1372
rect 1220 1371 1221 1375
rect 1215 1370 1221 1371
rect 1574 1375 1581 1376
rect 1574 1371 1575 1375
rect 1580 1371 1581 1375
rect 1574 1370 1581 1371
rect 1911 1375 1917 1376
rect 1911 1371 1912 1375
rect 1916 1374 1917 1375
rect 1999 1375 2005 1376
rect 1999 1374 2000 1375
rect 1916 1372 2000 1374
rect 1916 1371 1917 1372
rect 1911 1370 1917 1371
rect 1999 1371 2000 1372
rect 2004 1371 2005 1375
rect 1999 1370 2005 1371
rect 110 1368 116 1369
rect 1934 1368 1940 1369
rect 110 1364 111 1368
rect 115 1364 116 1368
rect 110 1363 116 1364
rect 130 1367 136 1368
rect 130 1363 131 1367
rect 135 1363 136 1367
rect 130 1362 136 1363
rect 410 1367 416 1368
rect 410 1363 411 1367
rect 415 1363 416 1367
rect 410 1362 416 1363
rect 738 1367 744 1368
rect 738 1363 739 1367
rect 743 1363 744 1367
rect 738 1362 744 1363
rect 1090 1367 1096 1368
rect 1090 1363 1091 1367
rect 1095 1363 1096 1367
rect 1090 1362 1096 1363
rect 1450 1367 1456 1368
rect 1450 1363 1451 1367
rect 1455 1363 1456 1367
rect 1450 1362 1456 1363
rect 1786 1367 1792 1368
rect 1786 1363 1787 1367
rect 1791 1363 1792 1367
rect 1934 1364 1935 1368
rect 1939 1364 1940 1368
rect 2839 1367 2845 1368
rect 2839 1366 2840 1367
rect 2661 1364 2840 1366
rect 1934 1363 1940 1364
rect 2282 1363 2288 1364
rect 1786 1362 1792 1363
rect 2282 1359 2283 1363
rect 2287 1359 2288 1363
rect 2839 1363 2840 1364
rect 2844 1363 2845 1367
rect 2839 1362 2845 1363
rect 2934 1367 2940 1368
rect 2934 1363 2935 1367
rect 2939 1363 2940 1367
rect 3370 1367 3376 1368
rect 3370 1366 3371 1367
rect 3221 1364 3371 1366
rect 2934 1362 2940 1363
rect 3370 1363 3371 1364
rect 3375 1363 3376 1367
rect 3370 1362 3376 1363
rect 3402 1363 3408 1364
rect 2282 1358 2288 1359
rect 3402 1359 3403 1363
rect 3407 1359 3408 1363
rect 3402 1358 3408 1359
rect 3658 1363 3664 1364
rect 3658 1359 3659 1363
rect 3663 1359 3664 1363
rect 3658 1358 3664 1359
rect 4682 1355 4688 1356
rect 158 1352 164 1353
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 158 1348 159 1352
rect 163 1348 164 1352
rect 158 1347 164 1348
rect 438 1352 444 1353
rect 438 1348 439 1352
rect 443 1348 444 1352
rect 438 1347 444 1348
rect 766 1352 772 1353
rect 766 1348 767 1352
rect 771 1348 772 1352
rect 766 1347 772 1348
rect 1118 1352 1124 1353
rect 1118 1348 1119 1352
rect 1123 1348 1124 1352
rect 1118 1347 1124 1348
rect 1478 1352 1484 1353
rect 1478 1348 1479 1352
rect 1483 1348 1484 1352
rect 1478 1347 1484 1348
rect 1814 1352 1820 1353
rect 1814 1348 1815 1352
rect 1819 1348 1820 1352
rect 1814 1347 1820 1348
rect 1934 1351 1940 1352
rect 1934 1347 1935 1351
rect 1939 1347 1940 1351
rect 4682 1351 4683 1355
rect 4687 1354 4688 1355
rect 4687 1352 5301 1354
rect 4687 1351 4688 1352
rect 4682 1350 4688 1351
rect 110 1346 116 1347
rect 1934 1346 1940 1347
rect 3954 1347 3960 1348
rect 3954 1343 3955 1347
rect 3959 1346 3960 1347
rect 3983 1347 3989 1348
rect 3983 1346 3984 1347
rect 3959 1344 3984 1346
rect 3959 1343 3960 1344
rect 3954 1342 3960 1343
rect 3983 1343 3984 1344
rect 3988 1343 3989 1347
rect 3983 1342 3989 1343
rect 4183 1347 4189 1348
rect 4183 1343 4184 1347
rect 4188 1346 4189 1347
rect 4314 1347 4320 1348
rect 4314 1346 4315 1347
rect 4188 1344 4315 1346
rect 4188 1343 4189 1344
rect 4183 1342 4189 1343
rect 4314 1343 4315 1344
rect 4319 1343 4320 1347
rect 4314 1342 4320 1343
rect 4431 1347 4437 1348
rect 4431 1343 4432 1347
rect 4436 1346 4437 1347
rect 4586 1347 4592 1348
rect 4586 1346 4587 1347
rect 4436 1344 4587 1346
rect 4436 1343 4437 1344
rect 4431 1342 4437 1343
rect 4586 1343 4587 1344
rect 4591 1343 4592 1347
rect 4586 1342 4592 1343
rect 4703 1347 4709 1348
rect 4703 1343 4704 1347
rect 4708 1346 4709 1347
rect 4882 1347 4888 1348
rect 4882 1346 4883 1347
rect 4708 1344 4883 1346
rect 4708 1343 4709 1344
rect 4703 1342 4709 1343
rect 4882 1343 4883 1344
rect 4887 1343 4888 1347
rect 4882 1342 4888 1343
rect 4999 1347 5005 1348
rect 4999 1343 5000 1347
rect 5004 1346 5005 1347
rect 5194 1347 5200 1348
rect 5194 1346 5195 1347
rect 5004 1344 5195 1346
rect 5004 1343 5005 1344
rect 4999 1342 5005 1343
rect 5194 1343 5195 1344
rect 5199 1343 5200 1347
rect 5299 1346 5301 1352
rect 5311 1347 5317 1348
rect 5311 1346 5312 1347
rect 5299 1344 5312 1346
rect 5194 1342 5200 1343
rect 5311 1343 5312 1344
rect 5316 1343 5317 1347
rect 5311 1342 5317 1343
rect 5610 1347 5616 1348
rect 5610 1343 5611 1347
rect 5615 1346 5616 1347
rect 5623 1347 5629 1348
rect 5623 1346 5624 1347
rect 5615 1344 5624 1346
rect 5615 1343 5616 1344
rect 5610 1342 5616 1343
rect 5623 1343 5624 1344
rect 5628 1343 5629 1347
rect 5623 1342 5629 1343
rect 3838 1340 3844 1341
rect 5662 1340 5668 1341
rect 3838 1336 3839 1340
rect 3843 1336 3844 1340
rect 3838 1335 3844 1336
rect 3858 1339 3864 1340
rect 3858 1335 3859 1339
rect 3863 1335 3864 1339
rect 3858 1334 3864 1335
rect 4058 1339 4064 1340
rect 4058 1335 4059 1339
rect 4063 1335 4064 1339
rect 4058 1334 4064 1335
rect 4306 1339 4312 1340
rect 4306 1335 4307 1339
rect 4311 1335 4312 1339
rect 4306 1334 4312 1335
rect 4578 1339 4584 1340
rect 4578 1335 4579 1339
rect 4583 1335 4584 1339
rect 4578 1334 4584 1335
rect 4874 1339 4880 1340
rect 4874 1335 4875 1339
rect 4879 1335 4880 1339
rect 4874 1334 4880 1335
rect 5186 1339 5192 1340
rect 5186 1335 5187 1339
rect 5191 1335 5192 1339
rect 5186 1334 5192 1335
rect 5498 1339 5504 1340
rect 5498 1335 5499 1339
rect 5503 1335 5504 1339
rect 5662 1336 5663 1340
rect 5667 1336 5668 1340
rect 5662 1335 5668 1336
rect 5498 1334 5504 1335
rect 3886 1324 3892 1325
rect 2119 1323 2125 1324
rect 2119 1319 2120 1323
rect 2124 1322 2125 1323
rect 2282 1323 2288 1324
rect 2282 1322 2283 1323
rect 2124 1320 2283 1322
rect 2124 1319 2125 1320
rect 2119 1318 2125 1319
rect 2282 1319 2283 1320
rect 2287 1319 2288 1323
rect 2282 1318 2288 1319
rect 2298 1323 2304 1324
rect 2298 1319 2299 1323
rect 2303 1322 2304 1323
rect 2399 1323 2405 1324
rect 2399 1322 2400 1323
rect 2303 1320 2400 1322
rect 2303 1319 2304 1320
rect 2298 1318 2304 1319
rect 2399 1319 2400 1320
rect 2404 1319 2405 1323
rect 2399 1318 2405 1319
rect 2686 1323 2693 1324
rect 2686 1319 2687 1323
rect 2692 1319 2693 1323
rect 2686 1318 2693 1319
rect 2839 1323 2845 1324
rect 2839 1319 2840 1323
rect 2844 1322 2845 1323
rect 2967 1323 2973 1324
rect 2967 1322 2968 1323
rect 2844 1320 2968 1322
rect 2844 1319 2845 1320
rect 2839 1318 2845 1319
rect 2967 1319 2968 1320
rect 2972 1319 2973 1323
rect 2967 1318 2973 1319
rect 3247 1323 3253 1324
rect 3247 1319 3248 1323
rect 3252 1322 3253 1323
rect 3402 1323 3408 1324
rect 3402 1322 3403 1323
rect 3252 1320 3403 1322
rect 3252 1319 3253 1320
rect 3247 1318 3253 1319
rect 3402 1319 3403 1320
rect 3407 1319 3408 1323
rect 3402 1318 3408 1319
rect 3519 1323 3525 1324
rect 3519 1319 3520 1323
rect 3524 1322 3525 1323
rect 3658 1323 3664 1324
rect 3658 1322 3659 1323
rect 3524 1320 3659 1322
rect 3524 1319 3525 1320
rect 3519 1318 3525 1319
rect 3658 1319 3659 1320
rect 3663 1319 3664 1323
rect 3658 1318 3664 1319
rect 3775 1323 3784 1324
rect 3775 1319 3776 1323
rect 3783 1319 3784 1323
rect 3775 1318 3784 1319
rect 3838 1323 3844 1324
rect 3838 1319 3839 1323
rect 3843 1319 3844 1323
rect 3886 1320 3887 1324
rect 3891 1320 3892 1324
rect 3886 1319 3892 1320
rect 4086 1324 4092 1325
rect 4086 1320 4087 1324
rect 4091 1320 4092 1324
rect 4086 1319 4092 1320
rect 4334 1324 4340 1325
rect 4334 1320 4335 1324
rect 4339 1320 4340 1324
rect 4334 1319 4340 1320
rect 4606 1324 4612 1325
rect 4606 1320 4607 1324
rect 4611 1320 4612 1324
rect 4606 1319 4612 1320
rect 4902 1324 4908 1325
rect 4902 1320 4903 1324
rect 4907 1320 4908 1324
rect 4902 1319 4908 1320
rect 5214 1324 5220 1325
rect 5214 1320 5215 1324
rect 5219 1320 5220 1324
rect 5214 1319 5220 1320
rect 5526 1324 5532 1325
rect 5526 1320 5527 1324
rect 5531 1320 5532 1324
rect 5526 1319 5532 1320
rect 5662 1323 5668 1324
rect 5662 1319 5663 1323
rect 5667 1319 5668 1323
rect 3838 1318 3844 1319
rect 5662 1318 5668 1319
rect 1974 1316 1980 1317
rect 3798 1316 3804 1317
rect 1974 1312 1975 1316
rect 1979 1312 1980 1316
rect 1974 1311 1980 1312
rect 1994 1315 2000 1316
rect 1994 1311 1995 1315
rect 1999 1311 2000 1315
rect 1994 1310 2000 1311
rect 2274 1315 2280 1316
rect 2274 1311 2275 1315
rect 2279 1311 2280 1315
rect 2274 1310 2280 1311
rect 2562 1315 2568 1316
rect 2562 1311 2563 1315
rect 2567 1311 2568 1315
rect 2562 1310 2568 1311
rect 2842 1315 2848 1316
rect 2842 1311 2843 1315
rect 2847 1311 2848 1315
rect 2842 1310 2848 1311
rect 3122 1315 3128 1316
rect 3122 1311 3123 1315
rect 3127 1311 3128 1315
rect 3122 1310 3128 1311
rect 3394 1315 3400 1316
rect 3394 1311 3395 1315
rect 3399 1311 3400 1315
rect 3394 1310 3400 1311
rect 3650 1315 3656 1316
rect 3650 1311 3651 1315
rect 3655 1311 3656 1315
rect 3798 1312 3799 1316
rect 3803 1312 3804 1316
rect 3798 1311 3804 1312
rect 3650 1310 3656 1311
rect 2022 1300 2028 1301
rect 1974 1299 1980 1300
rect 1974 1295 1975 1299
rect 1979 1295 1980 1299
rect 2022 1296 2023 1300
rect 2027 1296 2028 1300
rect 2022 1295 2028 1296
rect 2302 1300 2308 1301
rect 2302 1296 2303 1300
rect 2307 1296 2308 1300
rect 2302 1295 2308 1296
rect 2590 1300 2596 1301
rect 2590 1296 2591 1300
rect 2595 1296 2596 1300
rect 2590 1295 2596 1296
rect 2870 1300 2876 1301
rect 2870 1296 2871 1300
rect 2875 1296 2876 1300
rect 2870 1295 2876 1296
rect 3150 1300 3156 1301
rect 3150 1296 3151 1300
rect 3155 1296 3156 1300
rect 3150 1295 3156 1296
rect 3422 1300 3428 1301
rect 3422 1296 3423 1300
rect 3427 1296 3428 1300
rect 3422 1295 3428 1296
rect 3678 1300 3684 1301
rect 3678 1296 3679 1300
rect 3683 1296 3684 1300
rect 3678 1295 3684 1296
rect 3798 1299 3804 1300
rect 3798 1295 3799 1299
rect 3803 1295 3804 1299
rect 1974 1294 1980 1295
rect 3798 1294 3804 1295
rect 110 1293 116 1294
rect 1934 1293 1940 1294
rect 110 1289 111 1293
rect 115 1289 116 1293
rect 110 1288 116 1289
rect 158 1292 164 1293
rect 158 1288 159 1292
rect 163 1288 164 1292
rect 158 1287 164 1288
rect 358 1292 364 1293
rect 358 1288 359 1292
rect 363 1288 364 1292
rect 358 1287 364 1288
rect 574 1292 580 1293
rect 574 1288 575 1292
rect 579 1288 580 1292
rect 574 1287 580 1288
rect 774 1292 780 1293
rect 774 1288 775 1292
rect 779 1288 780 1292
rect 774 1287 780 1288
rect 966 1292 972 1293
rect 966 1288 967 1292
rect 971 1288 972 1292
rect 966 1287 972 1288
rect 1150 1292 1156 1293
rect 1150 1288 1151 1292
rect 1155 1288 1156 1292
rect 1150 1287 1156 1288
rect 1326 1292 1332 1293
rect 1326 1288 1327 1292
rect 1331 1288 1332 1292
rect 1326 1287 1332 1288
rect 1494 1292 1500 1293
rect 1494 1288 1495 1292
rect 1499 1288 1500 1292
rect 1494 1287 1500 1288
rect 1662 1292 1668 1293
rect 1662 1288 1663 1292
rect 1667 1288 1668 1292
rect 1662 1287 1668 1288
rect 1814 1292 1820 1293
rect 1814 1288 1815 1292
rect 1819 1288 1820 1292
rect 1934 1289 1935 1293
rect 1939 1289 1940 1293
rect 1934 1288 1940 1289
rect 1814 1287 1820 1288
rect 130 1277 136 1278
rect 110 1276 116 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 130 1273 131 1277
rect 135 1273 136 1277
rect 130 1272 136 1273
rect 330 1277 336 1278
rect 330 1273 331 1277
rect 335 1273 336 1277
rect 330 1272 336 1273
rect 546 1277 552 1278
rect 546 1273 547 1277
rect 551 1273 552 1277
rect 546 1272 552 1273
rect 746 1277 752 1278
rect 746 1273 747 1277
rect 751 1273 752 1277
rect 746 1272 752 1273
rect 938 1277 944 1278
rect 938 1273 939 1277
rect 943 1273 944 1277
rect 938 1272 944 1273
rect 1122 1277 1128 1278
rect 1122 1273 1123 1277
rect 1127 1273 1128 1277
rect 1122 1272 1128 1273
rect 1298 1277 1304 1278
rect 1298 1273 1299 1277
rect 1303 1273 1304 1277
rect 1298 1272 1304 1273
rect 1466 1277 1472 1278
rect 1466 1273 1467 1277
rect 1471 1273 1472 1277
rect 1466 1272 1472 1273
rect 1634 1277 1640 1278
rect 1634 1273 1635 1277
rect 1639 1273 1640 1277
rect 1634 1272 1640 1273
rect 1786 1277 1792 1278
rect 1786 1273 1787 1277
rect 1791 1273 1792 1277
rect 1786 1272 1792 1273
rect 1934 1276 1940 1277
rect 1934 1272 1935 1276
rect 1939 1272 1940 1276
rect 110 1271 116 1272
rect 1934 1271 1940 1272
rect 226 1267 232 1268
rect 226 1263 227 1267
rect 231 1266 232 1267
rect 255 1267 261 1268
rect 255 1266 256 1267
rect 231 1264 256 1266
rect 231 1263 232 1264
rect 226 1262 232 1263
rect 255 1263 256 1264
rect 260 1263 261 1267
rect 255 1262 261 1263
rect 386 1267 392 1268
rect 386 1263 387 1267
rect 391 1266 392 1267
rect 455 1267 461 1268
rect 455 1266 456 1267
rect 391 1264 456 1266
rect 391 1263 392 1264
rect 386 1262 392 1263
rect 455 1263 456 1264
rect 460 1263 461 1267
rect 455 1262 461 1263
rect 535 1267 541 1268
rect 535 1263 536 1267
rect 540 1266 541 1267
rect 671 1267 677 1268
rect 671 1266 672 1267
rect 540 1264 672 1266
rect 540 1263 541 1264
rect 535 1262 541 1263
rect 671 1263 672 1264
rect 676 1263 677 1267
rect 671 1262 677 1263
rect 870 1267 877 1268
rect 870 1263 871 1267
rect 876 1263 877 1267
rect 870 1262 877 1263
rect 903 1267 909 1268
rect 903 1263 904 1267
rect 908 1266 909 1267
rect 1063 1267 1069 1268
rect 1063 1266 1064 1267
rect 908 1264 1064 1266
rect 908 1263 909 1264
rect 903 1262 909 1263
rect 1063 1263 1064 1264
rect 1068 1263 1069 1267
rect 1063 1262 1069 1263
rect 1247 1267 1256 1268
rect 1247 1263 1248 1267
rect 1255 1263 1256 1267
rect 1247 1262 1256 1263
rect 1423 1267 1432 1268
rect 1423 1263 1424 1267
rect 1431 1263 1432 1267
rect 1423 1262 1432 1263
rect 1591 1267 1600 1268
rect 1591 1263 1592 1267
rect 1599 1263 1600 1267
rect 1591 1262 1600 1263
rect 1759 1267 1768 1268
rect 1759 1263 1760 1267
rect 1767 1263 1768 1267
rect 1759 1262 1768 1263
rect 1882 1267 1888 1268
rect 1882 1263 1883 1267
rect 1887 1266 1888 1267
rect 1911 1267 1917 1268
rect 1911 1266 1912 1267
rect 1887 1264 1912 1266
rect 1887 1263 1888 1264
rect 1882 1262 1888 1263
rect 1911 1263 1912 1264
rect 1916 1263 1917 1267
rect 1911 1262 1917 1263
rect 3838 1257 3844 1258
rect 5662 1257 5668 1258
rect 3838 1253 3839 1257
rect 3843 1253 3844 1257
rect 3838 1252 3844 1253
rect 4614 1256 4620 1257
rect 4614 1252 4615 1256
rect 4619 1252 4620 1256
rect 4614 1251 4620 1252
rect 4790 1256 4796 1257
rect 4790 1252 4791 1256
rect 4795 1252 4796 1256
rect 4790 1251 4796 1252
rect 4974 1256 4980 1257
rect 4974 1252 4975 1256
rect 4979 1252 4980 1256
rect 4974 1251 4980 1252
rect 5166 1256 5172 1257
rect 5166 1252 5167 1256
rect 5171 1252 5172 1256
rect 5166 1251 5172 1252
rect 5366 1256 5372 1257
rect 5366 1252 5367 1256
rect 5371 1252 5372 1256
rect 5366 1251 5372 1252
rect 5542 1256 5548 1257
rect 5542 1252 5543 1256
rect 5547 1252 5548 1256
rect 5662 1253 5663 1257
rect 5667 1253 5668 1257
rect 5662 1252 5668 1253
rect 5542 1251 5548 1252
rect 4586 1241 4592 1242
rect 3838 1240 3844 1241
rect 3838 1236 3839 1240
rect 3843 1236 3844 1240
rect 4586 1237 4587 1241
rect 4591 1237 4592 1241
rect 4586 1236 4592 1237
rect 4762 1241 4768 1242
rect 4762 1237 4763 1241
rect 4767 1237 4768 1241
rect 4762 1236 4768 1237
rect 4946 1241 4952 1242
rect 4946 1237 4947 1241
rect 4951 1237 4952 1241
rect 4946 1236 4952 1237
rect 5138 1241 5144 1242
rect 5138 1237 5139 1241
rect 5143 1237 5144 1241
rect 5138 1236 5144 1237
rect 5338 1241 5344 1242
rect 5338 1237 5339 1241
rect 5343 1237 5344 1241
rect 5338 1236 5344 1237
rect 5514 1241 5520 1242
rect 5514 1237 5515 1241
rect 5519 1237 5520 1241
rect 5514 1236 5520 1237
rect 5662 1240 5668 1241
rect 5662 1236 5663 1240
rect 5667 1236 5668 1240
rect 3838 1235 3844 1236
rect 5662 1235 5668 1236
rect 4711 1231 4720 1232
rect 226 1227 232 1228
rect 226 1223 227 1227
rect 231 1223 232 1227
rect 535 1227 541 1228
rect 535 1226 536 1227
rect 429 1224 536 1226
rect 226 1222 232 1223
rect 535 1223 536 1224
rect 540 1223 541 1227
rect 535 1222 541 1223
rect 543 1227 549 1228
rect 543 1223 544 1227
rect 548 1226 549 1227
rect 903 1227 909 1228
rect 903 1226 904 1227
rect 548 1224 553 1226
rect 845 1224 904 1226
rect 548 1223 549 1224
rect 543 1222 549 1223
rect 903 1223 904 1224
rect 908 1223 909 1227
rect 903 1222 909 1223
rect 1034 1227 1040 1228
rect 1034 1223 1035 1227
rect 1039 1223 1040 1227
rect 1034 1222 1040 1223
rect 1218 1227 1224 1228
rect 1218 1223 1219 1227
rect 1223 1223 1224 1227
rect 1218 1222 1224 1223
rect 1250 1227 1256 1228
rect 1250 1223 1251 1227
rect 1255 1226 1256 1227
rect 1426 1227 1432 1228
rect 1255 1224 1305 1226
rect 1255 1223 1256 1224
rect 1250 1222 1256 1223
rect 1426 1223 1427 1227
rect 1431 1226 1432 1227
rect 1594 1227 1600 1228
rect 1431 1224 1473 1226
rect 1431 1223 1432 1224
rect 1426 1222 1432 1223
rect 1594 1223 1595 1227
rect 1599 1226 1600 1227
rect 1762 1227 1768 1228
rect 1599 1224 1641 1226
rect 1599 1223 1600 1224
rect 1594 1222 1600 1223
rect 1762 1223 1763 1227
rect 1767 1226 1768 1227
rect 4711 1227 4712 1231
rect 4719 1227 4720 1231
rect 4711 1226 4720 1227
rect 4887 1231 4896 1232
rect 4887 1227 4888 1231
rect 4895 1227 4896 1231
rect 4887 1226 4896 1227
rect 5071 1231 5080 1232
rect 5071 1227 5072 1231
rect 5079 1227 5080 1231
rect 5071 1226 5080 1227
rect 5082 1231 5088 1232
rect 5082 1227 5083 1231
rect 5087 1230 5088 1231
rect 5263 1231 5269 1232
rect 5263 1230 5264 1231
rect 5087 1228 5264 1230
rect 5087 1227 5088 1228
rect 5082 1226 5088 1227
rect 5263 1227 5264 1228
rect 5268 1227 5269 1231
rect 5263 1226 5269 1227
rect 5463 1231 5472 1232
rect 5463 1227 5464 1231
rect 5471 1227 5472 1231
rect 5463 1226 5472 1227
rect 5618 1231 5624 1232
rect 5618 1227 5619 1231
rect 5623 1230 5624 1231
rect 5639 1231 5645 1232
rect 5639 1230 5640 1231
rect 5623 1228 5640 1230
rect 5623 1227 5624 1228
rect 5618 1226 5624 1227
rect 5639 1227 5640 1228
rect 5644 1227 5645 1231
rect 5639 1226 5645 1227
rect 1767 1224 1793 1226
rect 1767 1223 1768 1224
rect 1762 1222 1768 1223
rect 1974 1217 1980 1218
rect 3798 1217 3804 1218
rect 1974 1213 1975 1217
rect 1979 1213 1980 1217
rect 1974 1212 1980 1213
rect 2654 1216 2660 1217
rect 2654 1212 2655 1216
rect 2659 1212 2660 1216
rect 2654 1211 2660 1212
rect 2830 1216 2836 1217
rect 2830 1212 2831 1216
rect 2835 1212 2836 1216
rect 2830 1211 2836 1212
rect 3006 1216 3012 1217
rect 3006 1212 3007 1216
rect 3011 1212 3012 1216
rect 3006 1211 3012 1212
rect 3182 1216 3188 1217
rect 3182 1212 3183 1216
rect 3187 1212 3188 1216
rect 3182 1211 3188 1212
rect 3358 1216 3364 1217
rect 3358 1212 3359 1216
rect 3363 1212 3364 1216
rect 3358 1211 3364 1212
rect 3542 1216 3548 1217
rect 3542 1212 3543 1216
rect 3547 1212 3548 1216
rect 3798 1213 3799 1217
rect 3803 1213 3804 1217
rect 3798 1212 3804 1213
rect 3542 1211 3548 1212
rect 2626 1201 2632 1202
rect 1974 1200 1980 1201
rect 1974 1196 1975 1200
rect 1979 1196 1980 1200
rect 2626 1197 2627 1201
rect 2631 1197 2632 1201
rect 2626 1196 2632 1197
rect 2802 1201 2808 1202
rect 2802 1197 2803 1201
rect 2807 1197 2808 1201
rect 2802 1196 2808 1197
rect 2978 1201 2984 1202
rect 2978 1197 2979 1201
rect 2983 1197 2984 1201
rect 2978 1196 2984 1197
rect 3154 1201 3160 1202
rect 3154 1197 3155 1201
rect 3159 1197 3160 1201
rect 3154 1196 3160 1197
rect 3330 1201 3336 1202
rect 3330 1197 3331 1201
rect 3335 1197 3336 1201
rect 3330 1196 3336 1197
rect 3514 1201 3520 1202
rect 3514 1197 3515 1201
rect 3519 1197 3520 1201
rect 3514 1196 3520 1197
rect 3798 1200 3804 1201
rect 3798 1196 3799 1200
rect 3803 1196 3804 1200
rect 1974 1195 1980 1196
rect 3798 1195 3804 1196
rect 2751 1191 2760 1192
rect 2751 1187 2752 1191
rect 2759 1187 2760 1191
rect 2927 1191 2933 1192
rect 2927 1190 2928 1191
rect 2751 1186 2760 1187
rect 2779 1188 2928 1190
rect 270 1183 276 1184
rect 270 1182 271 1183
rect 229 1180 271 1182
rect 270 1179 271 1180
rect 275 1179 276 1183
rect 270 1178 276 1179
rect 386 1183 392 1184
rect 386 1179 387 1183
rect 391 1179 392 1183
rect 870 1183 876 1184
rect 386 1178 392 1179
rect 482 1179 488 1180
rect 482 1175 483 1179
rect 487 1175 488 1179
rect 482 1174 488 1175
rect 666 1179 672 1180
rect 666 1175 667 1179
rect 671 1175 672 1179
rect 870 1179 871 1183
rect 875 1179 876 1183
rect 1327 1183 1333 1184
rect 1327 1182 1328 1183
rect 1269 1180 1328 1182
rect 870 1178 876 1179
rect 1010 1179 1016 1180
rect 666 1174 672 1175
rect 1010 1175 1011 1179
rect 1015 1175 1016 1179
rect 1327 1179 1328 1180
rect 1332 1179 1333 1183
rect 1482 1183 1488 1184
rect 1482 1182 1483 1183
rect 1429 1180 1483 1182
rect 1327 1178 1333 1179
rect 1482 1179 1483 1180
rect 1487 1179 1488 1183
rect 1647 1183 1653 1184
rect 1647 1182 1648 1183
rect 1589 1180 1648 1182
rect 1482 1178 1488 1179
rect 1647 1179 1648 1180
rect 1652 1179 1653 1183
rect 2118 1183 2124 1184
rect 2118 1182 2119 1183
rect 1885 1180 2119 1182
rect 1647 1178 1653 1179
rect 1746 1179 1752 1180
rect 1010 1174 1016 1175
rect 1746 1175 1747 1179
rect 1751 1175 1752 1179
rect 2118 1179 2119 1180
rect 2123 1179 2124 1183
rect 2118 1178 2124 1179
rect 2266 1183 2272 1184
rect 2266 1179 2267 1183
rect 2271 1182 2272 1183
rect 2779 1182 2781 1188
rect 2927 1187 2928 1188
rect 2932 1187 2933 1191
rect 2927 1186 2933 1187
rect 3103 1191 3109 1192
rect 3103 1187 3104 1191
rect 3108 1190 3109 1191
rect 3119 1191 3125 1192
rect 3119 1190 3120 1191
rect 3108 1188 3120 1190
rect 3108 1187 3109 1188
rect 3103 1186 3109 1187
rect 3119 1187 3120 1188
rect 3124 1187 3125 1191
rect 3119 1186 3125 1187
rect 3279 1191 3288 1192
rect 3279 1187 3280 1191
rect 3287 1187 3288 1191
rect 3279 1186 3288 1187
rect 3455 1191 3464 1192
rect 3455 1187 3456 1191
rect 3463 1187 3464 1191
rect 3639 1191 3645 1192
rect 3639 1190 3640 1191
rect 3455 1186 3464 1187
rect 3619 1188 3640 1190
rect 2271 1180 2781 1182
rect 3370 1183 3376 1184
rect 2271 1179 2272 1180
rect 2266 1178 2272 1179
rect 3370 1179 3371 1183
rect 3375 1182 3376 1183
rect 3619 1182 3621 1188
rect 3639 1187 3640 1188
rect 3644 1187 3645 1191
rect 3639 1186 3645 1187
rect 4682 1191 4688 1192
rect 4682 1187 4683 1191
rect 4687 1187 4688 1191
rect 4682 1186 4688 1187
rect 4714 1191 4720 1192
rect 4714 1187 4715 1191
rect 4719 1190 4720 1191
rect 4890 1191 4896 1192
rect 4719 1188 4769 1190
rect 4719 1187 4720 1188
rect 4714 1186 4720 1187
rect 4890 1187 4891 1191
rect 4895 1190 4896 1191
rect 5074 1191 5080 1192
rect 4895 1188 4953 1190
rect 4895 1187 4896 1188
rect 4890 1186 4896 1187
rect 5074 1187 5075 1191
rect 5079 1190 5080 1191
rect 5478 1191 5484 1192
rect 5478 1190 5479 1191
rect 5079 1188 5145 1190
rect 5437 1188 5479 1190
rect 5079 1187 5080 1188
rect 5074 1186 5080 1187
rect 5478 1187 5479 1188
rect 5483 1187 5484 1191
rect 5478 1186 5484 1187
rect 5610 1191 5616 1192
rect 5610 1187 5611 1191
rect 5615 1187 5616 1191
rect 5610 1186 5616 1187
rect 3375 1180 3621 1182
rect 3375 1179 3376 1180
rect 3370 1178 3376 1179
rect 1746 1174 1752 1175
rect 5082 1159 5088 1160
rect 5082 1158 5083 1159
rect 4972 1156 5083 1158
rect 4972 1154 4974 1156
rect 5082 1155 5083 1156
rect 5087 1155 5088 1159
rect 5082 1154 5088 1155
rect 5618 1155 5624 1156
rect 5618 1154 5619 1155
rect 4933 1152 4974 1154
rect 5613 1152 5619 1154
rect 2686 1151 2692 1152
rect 1746 1147 1752 1148
rect 1746 1143 1747 1147
rect 1751 1146 1752 1147
rect 2686 1147 2687 1151
rect 2691 1147 2692 1151
rect 2686 1146 2692 1147
rect 2754 1151 2760 1152
rect 2754 1147 2755 1151
rect 2759 1150 2760 1151
rect 3119 1151 3125 1152
rect 2759 1148 2809 1150
rect 2759 1147 2760 1148
rect 2754 1146 2760 1147
rect 1751 1144 1834 1146
rect 1751 1143 1752 1144
rect 1746 1142 1752 1143
rect 226 1139 232 1140
rect 226 1135 227 1139
rect 231 1138 232 1139
rect 255 1139 261 1140
rect 255 1138 256 1139
rect 231 1136 256 1138
rect 231 1135 232 1136
rect 226 1134 232 1135
rect 255 1135 256 1136
rect 260 1135 261 1139
rect 255 1134 261 1135
rect 415 1139 421 1140
rect 415 1135 416 1139
rect 420 1138 421 1139
rect 482 1139 488 1140
rect 482 1138 483 1139
rect 420 1136 483 1138
rect 420 1135 421 1136
rect 415 1134 421 1135
rect 482 1135 483 1136
rect 487 1135 488 1139
rect 482 1134 488 1135
rect 599 1139 605 1140
rect 599 1135 600 1139
rect 604 1138 605 1139
rect 666 1139 672 1140
rect 666 1138 667 1139
rect 604 1136 667 1138
rect 604 1135 605 1136
rect 599 1134 605 1135
rect 666 1135 667 1136
rect 671 1135 672 1139
rect 666 1134 672 1135
rect 754 1139 760 1140
rect 754 1135 755 1139
rect 759 1138 760 1139
rect 783 1139 789 1140
rect 783 1138 784 1139
rect 759 1136 784 1138
rect 759 1135 760 1136
rect 754 1134 760 1135
rect 783 1135 784 1136
rect 788 1135 789 1139
rect 783 1134 789 1135
rect 959 1139 965 1140
rect 959 1135 960 1139
rect 964 1138 965 1139
rect 1010 1139 1016 1140
rect 1010 1138 1011 1139
rect 964 1136 1011 1138
rect 964 1135 965 1136
rect 959 1134 965 1135
rect 1010 1135 1011 1136
rect 1015 1135 1016 1139
rect 1010 1134 1016 1135
rect 1127 1139 1133 1140
rect 1127 1135 1128 1139
rect 1132 1138 1133 1139
rect 1142 1139 1148 1140
rect 1142 1138 1143 1139
rect 1132 1136 1143 1138
rect 1132 1135 1133 1136
rect 1127 1134 1133 1135
rect 1142 1135 1143 1136
rect 1147 1135 1148 1139
rect 1142 1134 1148 1135
rect 1218 1139 1224 1140
rect 1218 1135 1219 1139
rect 1223 1138 1224 1139
rect 1295 1139 1301 1140
rect 1295 1138 1296 1139
rect 1223 1136 1296 1138
rect 1223 1135 1224 1136
rect 1218 1134 1224 1135
rect 1295 1135 1296 1136
rect 1300 1135 1301 1139
rect 1295 1134 1301 1135
rect 1327 1139 1333 1140
rect 1327 1135 1328 1139
rect 1332 1138 1333 1139
rect 1455 1139 1461 1140
rect 1455 1138 1456 1139
rect 1332 1136 1456 1138
rect 1332 1135 1333 1136
rect 1327 1134 1333 1135
rect 1455 1135 1456 1136
rect 1460 1135 1461 1139
rect 1455 1134 1461 1135
rect 1482 1139 1488 1140
rect 1482 1135 1483 1139
rect 1487 1138 1488 1139
rect 1615 1139 1621 1140
rect 1615 1138 1616 1139
rect 1487 1136 1616 1138
rect 1487 1135 1488 1136
rect 1482 1134 1488 1135
rect 1615 1135 1616 1136
rect 1620 1135 1621 1139
rect 1615 1134 1621 1135
rect 1647 1139 1653 1140
rect 1647 1135 1648 1139
rect 1652 1138 1653 1139
rect 1775 1139 1781 1140
rect 1775 1138 1776 1139
rect 1652 1136 1776 1138
rect 1652 1135 1653 1136
rect 1647 1134 1653 1135
rect 1775 1135 1776 1136
rect 1780 1135 1781 1139
rect 1832 1138 1834 1144
rect 3076 1142 3078 1149
rect 3119 1147 3120 1151
rect 3124 1150 3125 1151
rect 3282 1151 3288 1152
rect 3124 1148 3161 1150
rect 3124 1147 3125 1148
rect 3119 1146 3125 1147
rect 3282 1147 3283 1151
rect 3287 1150 3288 1151
rect 3458 1151 3464 1152
rect 3287 1148 3337 1150
rect 3287 1147 3288 1148
rect 3282 1146 3288 1147
rect 3458 1147 3459 1151
rect 3463 1150 3464 1151
rect 4978 1151 4984 1152
rect 3463 1148 3521 1150
rect 3463 1147 3464 1148
rect 3458 1146 3464 1147
rect 4978 1147 4979 1151
rect 4983 1147 4984 1151
rect 4978 1146 4984 1147
rect 5114 1151 5120 1152
rect 5114 1147 5115 1151
rect 5119 1147 5120 1151
rect 5114 1146 5120 1147
rect 5250 1151 5256 1152
rect 5250 1147 5251 1151
rect 5255 1147 5256 1151
rect 5250 1146 5256 1147
rect 5386 1151 5392 1152
rect 5386 1147 5387 1151
rect 5391 1147 5392 1151
rect 5618 1151 5619 1152
rect 5623 1151 5624 1155
rect 5618 1150 5624 1151
rect 5386 1146 5392 1147
rect 3234 1143 3240 1144
rect 3234 1142 3235 1143
rect 3076 1140 3235 1142
rect 1911 1139 1917 1140
rect 1911 1138 1912 1139
rect 1832 1136 1912 1138
rect 1775 1134 1781 1135
rect 1911 1135 1912 1136
rect 1916 1135 1917 1139
rect 3234 1139 3235 1140
rect 3239 1139 3240 1143
rect 3234 1138 3240 1139
rect 1911 1134 1917 1135
rect 110 1132 116 1133
rect 1934 1132 1940 1133
rect 110 1128 111 1132
rect 115 1128 116 1132
rect 110 1127 116 1128
rect 130 1131 136 1132
rect 130 1127 131 1131
rect 135 1127 136 1131
rect 130 1126 136 1127
rect 290 1131 296 1132
rect 290 1127 291 1131
rect 295 1127 296 1131
rect 290 1126 296 1127
rect 474 1131 480 1132
rect 474 1127 475 1131
rect 479 1127 480 1131
rect 474 1126 480 1127
rect 658 1131 664 1132
rect 658 1127 659 1131
rect 663 1127 664 1131
rect 658 1126 664 1127
rect 834 1131 840 1132
rect 834 1127 835 1131
rect 839 1127 840 1131
rect 834 1126 840 1127
rect 1002 1131 1008 1132
rect 1002 1127 1003 1131
rect 1007 1127 1008 1131
rect 1002 1126 1008 1127
rect 1170 1131 1176 1132
rect 1170 1127 1171 1131
rect 1175 1127 1176 1131
rect 1170 1126 1176 1127
rect 1330 1131 1336 1132
rect 1330 1127 1331 1131
rect 1335 1127 1336 1131
rect 1330 1126 1336 1127
rect 1490 1131 1496 1132
rect 1490 1127 1491 1131
rect 1495 1127 1496 1131
rect 1490 1126 1496 1127
rect 1650 1131 1656 1132
rect 1650 1127 1651 1131
rect 1655 1127 1656 1131
rect 1650 1126 1656 1127
rect 1786 1131 1792 1132
rect 1786 1127 1787 1131
rect 1791 1127 1792 1131
rect 1934 1128 1935 1132
rect 1939 1128 1940 1132
rect 1934 1127 1940 1128
rect 1786 1126 1792 1127
rect 158 1116 164 1117
rect 110 1115 116 1116
rect 110 1111 111 1115
rect 115 1111 116 1115
rect 158 1112 159 1116
rect 163 1112 164 1116
rect 158 1111 164 1112
rect 318 1116 324 1117
rect 318 1112 319 1116
rect 323 1112 324 1116
rect 318 1111 324 1112
rect 502 1116 508 1117
rect 502 1112 503 1116
rect 507 1112 508 1116
rect 502 1111 508 1112
rect 686 1116 692 1117
rect 686 1112 687 1116
rect 691 1112 692 1116
rect 686 1111 692 1112
rect 862 1116 868 1117
rect 862 1112 863 1116
rect 867 1112 868 1116
rect 862 1111 868 1112
rect 1030 1116 1036 1117
rect 1030 1112 1031 1116
rect 1035 1112 1036 1116
rect 1030 1111 1036 1112
rect 1198 1116 1204 1117
rect 1198 1112 1199 1116
rect 1203 1112 1204 1116
rect 1198 1111 1204 1112
rect 1358 1116 1364 1117
rect 1358 1112 1359 1116
rect 1363 1112 1364 1116
rect 1358 1111 1364 1112
rect 1518 1116 1524 1117
rect 1518 1112 1519 1116
rect 1523 1112 1524 1116
rect 1518 1111 1524 1112
rect 1678 1116 1684 1117
rect 1678 1112 1679 1116
rect 1683 1112 1684 1116
rect 1678 1111 1684 1112
rect 1814 1116 1820 1117
rect 1814 1112 1815 1116
rect 1819 1112 1820 1116
rect 1814 1111 1820 1112
rect 1934 1115 1940 1116
rect 1934 1111 1935 1115
rect 1939 1111 1940 1115
rect 110 1110 116 1111
rect 1934 1110 1940 1111
rect 4959 1111 4965 1112
rect 4959 1107 4960 1111
rect 4964 1110 4965 1111
rect 4978 1111 4984 1112
rect 4978 1110 4979 1111
rect 4964 1108 4979 1110
rect 4964 1107 4965 1108
rect 4959 1106 4965 1107
rect 4978 1107 4979 1108
rect 4983 1107 4984 1111
rect 4978 1106 4984 1107
rect 5095 1111 5101 1112
rect 5095 1107 5096 1111
rect 5100 1110 5101 1111
rect 5114 1111 5120 1112
rect 5114 1110 5115 1111
rect 5100 1108 5115 1110
rect 5100 1107 5101 1108
rect 5095 1106 5101 1107
rect 5114 1107 5115 1108
rect 5119 1107 5120 1111
rect 5114 1106 5120 1107
rect 5231 1111 5237 1112
rect 5231 1107 5232 1111
rect 5236 1110 5237 1111
rect 5250 1111 5256 1112
rect 5250 1110 5251 1111
rect 5236 1108 5251 1110
rect 5236 1107 5237 1108
rect 5231 1106 5237 1107
rect 5250 1107 5251 1108
rect 5255 1107 5256 1111
rect 5250 1106 5256 1107
rect 5367 1111 5373 1112
rect 5367 1107 5368 1111
rect 5372 1110 5373 1111
rect 5386 1111 5392 1112
rect 5386 1110 5387 1111
rect 5372 1108 5387 1110
rect 5372 1107 5373 1108
rect 5367 1106 5373 1107
rect 5386 1107 5387 1108
rect 5391 1107 5392 1111
rect 5386 1106 5392 1107
rect 5418 1111 5424 1112
rect 5418 1107 5419 1111
rect 5423 1110 5424 1111
rect 5503 1111 5509 1112
rect 5503 1110 5504 1111
rect 5423 1108 5504 1110
rect 5423 1107 5424 1108
rect 5418 1106 5424 1107
rect 5503 1107 5504 1108
rect 5508 1107 5509 1111
rect 5503 1106 5509 1107
rect 5610 1111 5616 1112
rect 5610 1107 5611 1111
rect 5615 1110 5616 1111
rect 5639 1111 5645 1112
rect 5639 1110 5640 1111
rect 5615 1108 5640 1110
rect 5615 1107 5616 1108
rect 5610 1106 5616 1107
rect 5639 1107 5640 1108
rect 5644 1107 5645 1111
rect 5639 1106 5645 1107
rect 3838 1104 3844 1105
rect 5662 1104 5668 1105
rect 2266 1103 2272 1104
rect 2090 1099 2096 1100
rect 2090 1095 2091 1099
rect 2095 1095 2096 1099
rect 2266 1099 2267 1103
rect 2271 1099 2272 1103
rect 3406 1103 3412 1104
rect 2266 1098 2272 1099
rect 2370 1099 2376 1100
rect 2090 1094 2096 1095
rect 2370 1095 2371 1099
rect 2375 1095 2376 1099
rect 2370 1094 2376 1095
rect 2642 1099 2648 1100
rect 2642 1095 2643 1099
rect 2647 1095 2648 1099
rect 2642 1094 2648 1095
rect 2730 1099 2736 1100
rect 2730 1095 2731 1099
rect 2735 1095 2736 1099
rect 2730 1094 2736 1095
rect 2898 1099 2904 1100
rect 2898 1095 2899 1099
rect 2903 1095 2904 1099
rect 2898 1094 2904 1095
rect 3066 1099 3072 1100
rect 3066 1095 3067 1099
rect 3071 1095 3072 1099
rect 3066 1094 3072 1095
rect 3226 1099 3232 1100
rect 3226 1095 3227 1099
rect 3231 1095 3232 1099
rect 3406 1099 3407 1103
rect 3411 1099 3412 1103
rect 3838 1100 3839 1104
rect 3843 1100 3844 1104
rect 3838 1099 3844 1100
rect 4834 1103 4840 1104
rect 4834 1099 4835 1103
rect 4839 1099 4840 1103
rect 3406 1098 3412 1099
rect 4834 1098 4840 1099
rect 4970 1103 4976 1104
rect 4970 1099 4971 1103
rect 4975 1099 4976 1103
rect 4970 1098 4976 1099
rect 5106 1103 5112 1104
rect 5106 1099 5107 1103
rect 5111 1099 5112 1103
rect 5106 1098 5112 1099
rect 5242 1103 5248 1104
rect 5242 1099 5243 1103
rect 5247 1099 5248 1103
rect 5242 1098 5248 1099
rect 5378 1103 5384 1104
rect 5378 1099 5379 1103
rect 5383 1099 5384 1103
rect 5378 1098 5384 1099
rect 5514 1103 5520 1104
rect 5514 1099 5515 1103
rect 5519 1099 5520 1103
rect 5662 1100 5663 1104
rect 5667 1100 5668 1104
rect 5662 1099 5668 1100
rect 5514 1098 5520 1099
rect 3226 1094 3232 1095
rect 4862 1088 4868 1089
rect 3838 1087 3844 1088
rect 3838 1083 3839 1087
rect 3843 1083 3844 1087
rect 4862 1084 4863 1088
rect 4867 1084 4868 1088
rect 4862 1083 4868 1084
rect 4998 1088 5004 1089
rect 4998 1084 4999 1088
rect 5003 1084 5004 1088
rect 4998 1083 5004 1084
rect 5134 1088 5140 1089
rect 5134 1084 5135 1088
rect 5139 1084 5140 1088
rect 5134 1083 5140 1084
rect 5270 1088 5276 1089
rect 5270 1084 5271 1088
rect 5275 1084 5276 1088
rect 5270 1083 5276 1084
rect 5406 1088 5412 1089
rect 5406 1084 5407 1088
rect 5411 1084 5412 1088
rect 5406 1083 5412 1084
rect 5542 1088 5548 1089
rect 5542 1084 5543 1088
rect 5547 1084 5548 1088
rect 5542 1083 5548 1084
rect 5662 1087 5668 1088
rect 5662 1083 5663 1087
rect 5667 1083 5668 1087
rect 3838 1082 3844 1083
rect 5662 1082 5668 1083
rect 2642 1067 2648 1068
rect 2642 1063 2643 1067
rect 2647 1066 2648 1067
rect 2647 1064 3354 1066
rect 2647 1063 2648 1064
rect 2642 1062 2648 1063
rect 2118 1059 2125 1060
rect 2118 1055 2119 1059
rect 2124 1055 2125 1059
rect 2118 1054 2125 1055
rect 2295 1059 2301 1060
rect 2295 1055 2296 1059
rect 2300 1058 2301 1059
rect 2370 1059 2376 1060
rect 2370 1058 2371 1059
rect 2300 1056 2371 1058
rect 2300 1055 2301 1056
rect 2295 1054 2301 1055
rect 2370 1055 2371 1056
rect 2375 1055 2376 1059
rect 2370 1054 2376 1055
rect 2487 1059 2496 1060
rect 2487 1055 2488 1059
rect 2495 1055 2496 1059
rect 2487 1054 2496 1055
rect 2671 1059 2677 1060
rect 2671 1055 2672 1059
rect 2676 1058 2677 1059
rect 2730 1059 2736 1060
rect 2730 1058 2731 1059
rect 2676 1056 2731 1058
rect 2676 1055 2677 1056
rect 2671 1054 2677 1055
rect 2730 1055 2731 1056
rect 2735 1055 2736 1059
rect 2730 1054 2736 1055
rect 2847 1059 2853 1060
rect 2847 1055 2848 1059
rect 2852 1058 2853 1059
rect 2898 1059 2904 1060
rect 2898 1058 2899 1059
rect 2852 1056 2899 1058
rect 2852 1055 2853 1056
rect 2847 1054 2853 1055
rect 2898 1055 2899 1056
rect 2903 1055 2904 1059
rect 2898 1054 2904 1055
rect 3015 1059 3021 1060
rect 3015 1055 3016 1059
rect 3020 1058 3021 1059
rect 3066 1059 3072 1060
rect 3066 1058 3067 1059
rect 3020 1056 3067 1058
rect 3020 1055 3021 1056
rect 3015 1054 3021 1055
rect 3066 1055 3067 1056
rect 3071 1055 3072 1059
rect 3066 1054 3072 1055
rect 3183 1059 3189 1060
rect 3183 1055 3184 1059
rect 3188 1058 3189 1059
rect 3226 1059 3232 1060
rect 3226 1058 3227 1059
rect 3188 1056 3227 1058
rect 3188 1055 3189 1056
rect 3183 1054 3189 1055
rect 3226 1055 3227 1056
rect 3231 1055 3232 1059
rect 3226 1054 3232 1055
rect 3234 1059 3240 1060
rect 3234 1055 3235 1059
rect 3239 1058 3240 1059
rect 3343 1059 3349 1060
rect 3343 1058 3344 1059
rect 3239 1056 3344 1058
rect 3239 1055 3240 1056
rect 3234 1054 3240 1055
rect 3343 1055 3344 1056
rect 3348 1055 3349 1059
rect 3352 1058 3354 1064
rect 3511 1059 3517 1060
rect 3511 1058 3512 1059
rect 3352 1056 3512 1058
rect 3343 1054 3349 1055
rect 3511 1055 3512 1056
rect 3516 1055 3517 1059
rect 3511 1054 3517 1055
rect 1974 1052 1980 1053
rect 3798 1052 3804 1053
rect 1974 1048 1975 1052
rect 1979 1048 1980 1052
rect 1974 1047 1980 1048
rect 1994 1051 2000 1052
rect 1994 1047 1995 1051
rect 1999 1047 2000 1051
rect 1994 1046 2000 1047
rect 2170 1051 2176 1052
rect 2170 1047 2171 1051
rect 2175 1047 2176 1051
rect 2170 1046 2176 1047
rect 2362 1051 2368 1052
rect 2362 1047 2363 1051
rect 2367 1047 2368 1051
rect 2362 1046 2368 1047
rect 2546 1051 2552 1052
rect 2546 1047 2547 1051
rect 2551 1047 2552 1051
rect 2546 1046 2552 1047
rect 2722 1051 2728 1052
rect 2722 1047 2723 1051
rect 2727 1047 2728 1051
rect 2722 1046 2728 1047
rect 2890 1051 2896 1052
rect 2890 1047 2891 1051
rect 2895 1047 2896 1051
rect 2890 1046 2896 1047
rect 3058 1051 3064 1052
rect 3058 1047 3059 1051
rect 3063 1047 3064 1051
rect 3058 1046 3064 1047
rect 3218 1051 3224 1052
rect 3218 1047 3219 1051
rect 3223 1047 3224 1051
rect 3218 1046 3224 1047
rect 3386 1051 3392 1052
rect 3386 1047 3387 1051
rect 3391 1047 3392 1051
rect 3798 1048 3799 1052
rect 3803 1048 3804 1052
rect 3798 1047 3804 1048
rect 3386 1046 3392 1047
rect 110 1045 116 1046
rect 1934 1045 1940 1046
rect 110 1041 111 1045
rect 115 1041 116 1045
rect 110 1040 116 1041
rect 174 1044 180 1045
rect 174 1040 175 1044
rect 179 1040 180 1044
rect 174 1039 180 1040
rect 430 1044 436 1045
rect 430 1040 431 1044
rect 435 1040 436 1044
rect 430 1039 436 1040
rect 686 1044 692 1045
rect 686 1040 687 1044
rect 691 1040 692 1044
rect 686 1039 692 1040
rect 950 1044 956 1045
rect 950 1040 951 1044
rect 955 1040 956 1044
rect 950 1039 956 1040
rect 1214 1044 1220 1045
rect 1214 1040 1215 1044
rect 1219 1040 1220 1044
rect 1934 1041 1935 1045
rect 1939 1041 1940 1045
rect 1934 1040 1940 1041
rect 1214 1039 1220 1040
rect 2022 1036 2028 1037
rect 1974 1035 1980 1036
rect 1974 1031 1975 1035
rect 1979 1031 1980 1035
rect 2022 1032 2023 1036
rect 2027 1032 2028 1036
rect 2022 1031 2028 1032
rect 2198 1036 2204 1037
rect 2198 1032 2199 1036
rect 2203 1032 2204 1036
rect 2198 1031 2204 1032
rect 2390 1036 2396 1037
rect 2390 1032 2391 1036
rect 2395 1032 2396 1036
rect 2390 1031 2396 1032
rect 2574 1036 2580 1037
rect 2574 1032 2575 1036
rect 2579 1032 2580 1036
rect 2574 1031 2580 1032
rect 2750 1036 2756 1037
rect 2750 1032 2751 1036
rect 2755 1032 2756 1036
rect 2750 1031 2756 1032
rect 2918 1036 2924 1037
rect 2918 1032 2919 1036
rect 2923 1032 2924 1036
rect 2918 1031 2924 1032
rect 3086 1036 3092 1037
rect 3086 1032 3087 1036
rect 3091 1032 3092 1036
rect 3086 1031 3092 1032
rect 3246 1036 3252 1037
rect 3246 1032 3247 1036
rect 3251 1032 3252 1036
rect 3246 1031 3252 1032
rect 3414 1036 3420 1037
rect 3414 1032 3415 1036
rect 3419 1032 3420 1036
rect 3414 1031 3420 1032
rect 3798 1035 3804 1036
rect 3798 1031 3799 1035
rect 3803 1031 3804 1035
rect 1974 1030 1980 1031
rect 3798 1030 3804 1031
rect 146 1029 152 1030
rect 110 1028 116 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 146 1025 147 1029
rect 151 1025 152 1029
rect 146 1024 152 1025
rect 402 1029 408 1030
rect 402 1025 403 1029
rect 407 1025 408 1029
rect 402 1024 408 1025
rect 658 1029 664 1030
rect 658 1025 659 1029
rect 663 1025 664 1029
rect 658 1024 664 1025
rect 922 1029 928 1030
rect 922 1025 923 1029
rect 927 1025 928 1029
rect 922 1024 928 1025
rect 1186 1029 1192 1030
rect 1186 1025 1187 1029
rect 1191 1025 1192 1029
rect 1186 1024 1192 1025
rect 1934 1028 1940 1029
rect 1934 1024 1935 1028
rect 1939 1024 1940 1028
rect 110 1023 116 1024
rect 1934 1023 1940 1024
rect 3838 1025 3844 1026
rect 5662 1025 5668 1026
rect 3838 1021 3839 1025
rect 3843 1021 3844 1025
rect 3838 1020 3844 1021
rect 4806 1024 4812 1025
rect 4806 1020 4807 1024
rect 4811 1020 4812 1024
rect 270 1019 277 1020
rect 270 1015 271 1019
rect 276 1015 277 1019
rect 270 1014 277 1015
rect 354 1019 360 1020
rect 354 1015 355 1019
rect 359 1018 360 1019
rect 527 1019 533 1020
rect 527 1018 528 1019
rect 359 1016 528 1018
rect 359 1015 360 1016
rect 354 1014 360 1015
rect 527 1015 528 1016
rect 532 1015 533 1019
rect 527 1014 533 1015
rect 778 1019 789 1020
rect 778 1015 779 1019
rect 783 1015 784 1019
rect 788 1015 789 1019
rect 778 1014 789 1015
rect 1002 1019 1008 1020
rect 1002 1015 1003 1019
rect 1007 1018 1008 1019
rect 1047 1019 1053 1020
rect 1047 1018 1048 1019
rect 1007 1016 1048 1018
rect 1007 1015 1008 1016
rect 1002 1014 1008 1015
rect 1047 1015 1048 1016
rect 1052 1015 1053 1019
rect 1047 1014 1053 1015
rect 1134 1019 1140 1020
rect 1134 1015 1135 1019
rect 1139 1018 1140 1019
rect 1311 1019 1317 1020
rect 4806 1019 4812 1020
rect 4942 1024 4948 1025
rect 4942 1020 4943 1024
rect 4947 1020 4948 1024
rect 4942 1019 4948 1020
rect 5078 1024 5084 1025
rect 5078 1020 5079 1024
rect 5083 1020 5084 1024
rect 5078 1019 5084 1020
rect 5214 1024 5220 1025
rect 5214 1020 5215 1024
rect 5219 1020 5220 1024
rect 5214 1019 5220 1020
rect 5350 1024 5356 1025
rect 5350 1020 5351 1024
rect 5355 1020 5356 1024
rect 5350 1019 5356 1020
rect 5486 1024 5492 1025
rect 5486 1020 5487 1024
rect 5491 1020 5492 1024
rect 5662 1021 5663 1025
rect 5667 1021 5668 1025
rect 5662 1020 5668 1021
rect 5486 1019 5492 1020
rect 1311 1018 1312 1019
rect 1139 1016 1312 1018
rect 1139 1015 1140 1016
rect 1134 1014 1140 1015
rect 1311 1015 1312 1016
rect 1316 1015 1317 1019
rect 1311 1014 1317 1015
rect 4778 1009 4784 1010
rect 3838 1008 3844 1009
rect 3838 1004 3839 1008
rect 3843 1004 3844 1008
rect 4778 1005 4779 1009
rect 4783 1005 4784 1009
rect 4778 1004 4784 1005
rect 4914 1009 4920 1010
rect 4914 1005 4915 1009
rect 4919 1005 4920 1009
rect 4914 1004 4920 1005
rect 5050 1009 5056 1010
rect 5050 1005 5051 1009
rect 5055 1005 5056 1009
rect 5050 1004 5056 1005
rect 5186 1009 5192 1010
rect 5186 1005 5187 1009
rect 5191 1005 5192 1009
rect 5186 1004 5192 1005
rect 5322 1009 5328 1010
rect 5322 1005 5323 1009
rect 5327 1005 5328 1009
rect 5322 1004 5328 1005
rect 5458 1009 5464 1010
rect 5458 1005 5459 1009
rect 5463 1005 5464 1009
rect 5458 1004 5464 1005
rect 5662 1008 5668 1009
rect 5662 1004 5663 1008
rect 5667 1004 5668 1008
rect 3838 1003 3844 1004
rect 5662 1003 5668 1004
rect 4903 999 4912 1000
rect 4903 995 4904 999
rect 4911 995 4912 999
rect 4903 994 4912 995
rect 5039 999 5048 1000
rect 5039 995 5040 999
rect 5047 995 5048 999
rect 5039 994 5048 995
rect 5175 999 5184 1000
rect 5175 995 5176 999
rect 5183 995 5184 999
rect 5311 999 5317 1000
rect 5311 998 5312 999
rect 5175 994 5184 995
rect 5299 996 5312 998
rect 4874 991 4880 992
rect 4874 987 4875 991
rect 4879 990 4880 991
rect 5299 990 5301 996
rect 5311 995 5312 996
rect 5316 995 5317 999
rect 5311 994 5317 995
rect 5330 999 5336 1000
rect 5330 995 5331 999
rect 5335 998 5336 999
rect 5447 999 5453 1000
rect 5447 998 5448 999
rect 5335 996 5448 998
rect 5335 995 5336 996
rect 5330 994 5336 995
rect 5447 995 5448 996
rect 5452 995 5453 999
rect 5447 994 5453 995
rect 5478 999 5484 1000
rect 5478 995 5479 999
rect 5483 998 5484 999
rect 5583 999 5589 1000
rect 5583 998 5584 999
rect 5483 996 5584 998
rect 5483 995 5484 996
rect 5478 994 5484 995
rect 5583 995 5584 996
rect 5588 995 5589 999
rect 5583 994 5589 995
rect 4879 988 5301 990
rect 4879 987 4880 988
rect 4874 986 4880 987
rect 354 979 360 980
rect 354 978 355 979
rect 245 976 355 978
rect 354 975 355 976
rect 359 975 360 979
rect 354 974 360 975
rect 362 979 368 980
rect 362 975 363 979
rect 367 978 368 979
rect 754 979 760 980
rect 367 976 409 978
rect 367 975 368 976
rect 362 974 368 975
rect 754 975 755 979
rect 759 975 760 979
rect 1134 979 1140 980
rect 1134 978 1135 979
rect 1021 976 1135 978
rect 754 974 760 975
rect 1134 975 1135 976
rect 1139 975 1140 979
rect 1134 974 1140 975
rect 1142 979 1148 980
rect 1142 975 1143 979
rect 1147 978 1148 979
rect 1147 976 1193 978
rect 1974 977 1980 978
rect 3798 977 3804 978
rect 1147 975 1148 976
rect 1142 974 1148 975
rect 1974 973 1975 977
rect 1979 973 1980 977
rect 1974 972 1980 973
rect 2022 976 2028 977
rect 2022 972 2023 976
rect 2027 972 2028 976
rect 2022 971 2028 972
rect 2190 976 2196 977
rect 2190 972 2191 976
rect 2195 972 2196 976
rect 2190 971 2196 972
rect 2374 976 2380 977
rect 2374 972 2375 976
rect 2379 972 2380 976
rect 2374 971 2380 972
rect 2566 976 2572 977
rect 2566 972 2567 976
rect 2571 972 2572 976
rect 2566 971 2572 972
rect 2758 976 2764 977
rect 2758 972 2759 976
rect 2763 972 2764 976
rect 2758 971 2764 972
rect 2942 976 2948 977
rect 2942 972 2943 976
rect 2947 972 2948 976
rect 2942 971 2948 972
rect 3126 976 3132 977
rect 3126 972 3127 976
rect 3131 972 3132 976
rect 3126 971 3132 972
rect 3310 976 3316 977
rect 3310 972 3311 976
rect 3315 972 3316 976
rect 3310 971 3316 972
rect 3494 976 3500 977
rect 3494 972 3495 976
rect 3499 972 3500 976
rect 3494 971 3500 972
rect 3678 976 3684 977
rect 3678 972 3679 976
rect 3683 972 3684 976
rect 3798 973 3799 977
rect 3803 973 3804 977
rect 3798 972 3804 973
rect 3678 971 3684 972
rect 5330 967 5336 968
rect 5330 966 5331 967
rect 5299 964 5331 966
rect 1994 961 2000 962
rect 1974 960 1980 961
rect 1974 956 1975 960
rect 1979 956 1980 960
rect 1994 957 1995 961
rect 1999 957 2000 961
rect 1994 956 2000 957
rect 2162 961 2168 962
rect 2162 957 2163 961
rect 2167 957 2168 961
rect 2162 956 2168 957
rect 2346 961 2352 962
rect 2346 957 2347 961
rect 2351 957 2352 961
rect 2346 956 2352 957
rect 2538 961 2544 962
rect 2538 957 2539 961
rect 2543 957 2544 961
rect 2538 956 2544 957
rect 2730 961 2736 962
rect 2730 957 2731 961
rect 2735 957 2736 961
rect 2730 956 2736 957
rect 2914 961 2920 962
rect 2914 957 2915 961
rect 2919 957 2920 961
rect 2914 956 2920 957
rect 3098 961 3104 962
rect 3098 957 3099 961
rect 3103 957 3104 961
rect 3098 956 3104 957
rect 3282 961 3288 962
rect 3282 957 3283 961
rect 3287 957 3288 961
rect 3282 956 3288 957
rect 3466 961 3472 962
rect 3466 957 3467 961
rect 3471 957 3472 961
rect 3466 956 3472 957
rect 3650 961 3656 962
rect 3650 957 3651 961
rect 3655 957 3656 961
rect 3650 956 3656 957
rect 3798 960 3804 961
rect 3798 956 3799 960
rect 3803 956 3804 960
rect 1974 955 1980 956
rect 3798 955 3804 956
rect 4874 959 4880 960
rect 4874 955 4875 959
rect 4879 955 4880 959
rect 4874 954 4880 955
rect 4906 959 4912 960
rect 4906 955 4907 959
rect 4911 958 4912 959
rect 5042 959 5048 960
rect 4911 956 4921 958
rect 4911 955 4912 956
rect 4906 954 4912 955
rect 5042 955 5043 959
rect 5047 958 5048 959
rect 5299 958 5301 964
rect 5330 963 5331 964
rect 5335 963 5336 967
rect 5330 962 5336 963
rect 5047 956 5057 958
rect 5285 956 5301 958
rect 5418 959 5424 960
rect 5047 955 5048 956
rect 5042 954 5048 955
rect 5418 955 5419 959
rect 5423 955 5424 959
rect 5418 954 5424 955
rect 5554 959 5560 960
rect 5554 955 5555 959
rect 5559 955 5560 959
rect 5554 954 5560 955
rect 2090 951 2096 952
rect 2090 947 2091 951
rect 2095 950 2096 951
rect 2119 951 2125 952
rect 2119 950 2120 951
rect 2095 948 2120 950
rect 2095 947 2096 948
rect 2090 946 2096 947
rect 2119 947 2120 948
rect 2124 947 2125 951
rect 2119 946 2125 947
rect 2154 951 2160 952
rect 2154 947 2155 951
rect 2159 950 2160 951
rect 2287 951 2293 952
rect 2287 950 2288 951
rect 2159 948 2288 950
rect 2159 947 2160 948
rect 2154 946 2160 947
rect 2287 947 2288 948
rect 2292 947 2293 951
rect 2287 946 2293 947
rect 2319 951 2325 952
rect 2319 947 2320 951
rect 2324 950 2325 951
rect 2471 951 2477 952
rect 2471 950 2472 951
rect 2324 948 2472 950
rect 2324 947 2325 948
rect 2319 946 2325 947
rect 2471 947 2472 948
rect 2476 947 2477 951
rect 2471 946 2477 947
rect 2663 951 2672 952
rect 2663 947 2664 951
rect 2671 947 2672 951
rect 2663 946 2672 947
rect 2855 951 2861 952
rect 2855 947 2856 951
rect 2860 950 2861 951
rect 2894 951 2900 952
rect 2894 950 2895 951
rect 2860 948 2895 950
rect 2860 947 2861 948
rect 2855 946 2861 947
rect 2894 947 2895 948
rect 2899 947 2900 951
rect 2894 946 2900 947
rect 3039 951 3048 952
rect 3039 947 3040 951
rect 3047 947 3048 951
rect 3039 946 3048 947
rect 3223 951 3232 952
rect 3223 947 3224 951
rect 3231 947 3232 951
rect 3223 946 3232 947
rect 3406 951 3413 952
rect 3406 947 3407 951
rect 3412 947 3413 951
rect 3591 951 3597 952
rect 3591 950 3592 951
rect 3406 946 3413 947
rect 3416 948 3592 950
rect 3010 943 3016 944
rect 3010 939 3011 943
rect 3015 942 3016 943
rect 3416 942 3418 948
rect 3591 947 3592 948
rect 3596 947 3597 951
rect 3591 946 3597 947
rect 3642 951 3648 952
rect 3642 947 3643 951
rect 3647 950 3648 951
rect 3775 951 3781 952
rect 3775 950 3776 951
rect 3647 948 3776 950
rect 3647 947 3648 948
rect 3642 946 3648 947
rect 3775 947 3776 948
rect 3780 947 3781 951
rect 3775 946 3781 947
rect 3015 940 3418 942
rect 3015 939 3016 940
rect 3010 938 3016 939
rect 270 935 276 936
rect 270 931 271 935
rect 275 931 276 935
rect 679 935 685 936
rect 679 934 680 935
rect 557 932 680 934
rect 270 930 276 931
rect 679 931 680 932
rect 684 931 685 935
rect 679 930 685 931
rect 778 935 784 936
rect 778 931 779 935
rect 783 931 784 935
rect 778 930 784 931
rect 1002 935 1008 936
rect 1002 931 1003 935
rect 1007 931 1008 935
rect 1002 930 1008 931
rect 1138 931 1144 932
rect 1138 927 1139 931
rect 1143 927 1144 931
rect 1138 926 1144 927
rect 1370 931 1376 932
rect 1370 927 1371 931
rect 1375 927 1376 931
rect 1370 926 1376 927
rect 4162 923 4168 924
rect 4162 922 4163 923
rect 4093 920 4163 922
rect 3954 919 3960 920
rect 3954 915 3955 919
rect 3959 915 3960 919
rect 4162 919 4163 920
rect 4167 919 4168 923
rect 4274 923 4280 924
rect 4274 922 4275 923
rect 4269 920 4275 922
rect 4162 918 4168 919
rect 4274 919 4275 920
rect 4279 919 4280 923
rect 5178 923 5184 924
rect 4274 918 4280 919
rect 4482 919 4488 920
rect 3954 914 3960 915
rect 4482 915 4483 919
rect 4487 915 4488 919
rect 4482 914 4488 915
rect 4650 919 4656 920
rect 4650 915 4651 919
rect 4655 915 4656 919
rect 4650 914 4656 915
rect 4938 919 4944 920
rect 4938 915 4939 919
rect 4943 915 4944 919
rect 5178 919 5179 923
rect 5183 922 5184 923
rect 5610 923 5616 924
rect 5183 920 5241 922
rect 5183 919 5184 920
rect 5178 918 5184 919
rect 5610 919 5611 923
rect 5615 919 5616 923
rect 5610 918 5616 919
rect 4938 914 4944 915
rect 2154 911 2160 912
rect 2154 910 2155 911
rect 2093 908 2155 910
rect 2154 907 2155 908
rect 2159 907 2160 911
rect 2319 911 2325 912
rect 2319 910 2320 911
rect 2261 908 2320 910
rect 2154 906 2160 907
rect 2319 907 2320 908
rect 2324 907 2325 911
rect 2319 906 2325 907
rect 2327 911 2333 912
rect 2327 907 2328 911
rect 2332 910 2333 911
rect 2490 911 2496 912
rect 2332 908 2353 910
rect 2332 907 2333 908
rect 2327 906 2333 907
rect 2490 907 2491 911
rect 2495 910 2496 911
rect 2666 911 2672 912
rect 2495 908 2545 910
rect 2495 907 2496 908
rect 2490 906 2496 907
rect 2666 907 2667 911
rect 2671 910 2672 911
rect 3010 911 3016 912
rect 2671 908 2737 910
rect 2671 907 2672 908
rect 2666 906 2672 907
rect 3010 907 3011 911
rect 3015 907 3016 911
rect 3010 906 3016 907
rect 3042 911 3048 912
rect 3042 907 3043 911
rect 3047 910 3048 911
rect 3226 911 3232 912
rect 3047 908 3105 910
rect 3047 907 3048 908
rect 3042 906 3048 907
rect 3226 907 3227 911
rect 3231 910 3232 911
rect 3642 911 3648 912
rect 3642 910 3643 911
rect 3231 908 3289 910
rect 3565 908 3643 910
rect 3231 907 3232 908
rect 3226 906 3232 907
rect 3642 907 3643 908
rect 3647 907 3648 911
rect 3642 906 3648 907
rect 3746 911 3752 912
rect 3746 907 3747 911
rect 3751 907 3752 911
rect 3746 906 3752 907
rect 359 891 368 892
rect 359 887 360 891
rect 367 887 368 891
rect 359 886 368 887
rect 498 891 504 892
rect 498 887 499 891
rect 503 890 504 891
rect 583 891 589 892
rect 583 890 584 891
rect 503 888 584 890
rect 503 887 504 888
rect 498 886 504 887
rect 583 887 584 888
rect 588 887 589 891
rect 583 886 589 887
rect 679 891 685 892
rect 679 887 680 891
rect 684 890 685 891
rect 807 891 813 892
rect 807 890 808 891
rect 684 888 808 890
rect 684 887 685 888
rect 679 886 685 887
rect 807 887 808 888
rect 812 887 813 891
rect 807 886 813 887
rect 1031 891 1037 892
rect 1031 887 1032 891
rect 1036 890 1037 891
rect 1138 891 1144 892
rect 1138 890 1139 891
rect 1036 888 1139 890
rect 1036 887 1037 888
rect 1031 886 1037 887
rect 1138 887 1139 888
rect 1143 887 1144 891
rect 1138 886 1144 887
rect 1255 891 1261 892
rect 1255 887 1256 891
rect 1260 890 1261 891
rect 1370 891 1376 892
rect 1370 890 1371 891
rect 1260 888 1371 890
rect 1260 887 1261 888
rect 1255 886 1261 887
rect 1370 887 1371 888
rect 1375 887 1376 891
rect 1370 886 1376 887
rect 1487 891 1496 892
rect 1487 887 1488 891
rect 1495 887 1496 891
rect 1487 886 1496 887
rect 4482 887 4488 888
rect 110 884 116 885
rect 1934 884 1940 885
rect 110 880 111 884
rect 115 880 116 884
rect 110 879 116 880
rect 234 883 240 884
rect 234 879 235 883
rect 239 879 240 883
rect 234 878 240 879
rect 458 883 464 884
rect 458 879 459 883
rect 463 879 464 883
rect 458 878 464 879
rect 682 883 688 884
rect 682 879 683 883
rect 687 879 688 883
rect 682 878 688 879
rect 906 883 912 884
rect 906 879 907 883
rect 911 879 912 883
rect 906 878 912 879
rect 1130 883 1136 884
rect 1130 879 1131 883
rect 1135 879 1136 883
rect 1130 878 1136 879
rect 1362 883 1368 884
rect 1362 879 1363 883
rect 1367 879 1368 883
rect 1934 880 1935 884
rect 1939 880 1940 884
rect 2526 883 2532 884
rect 2526 882 2527 883
rect 1934 879 1940 880
rect 2180 880 2527 882
rect 1362 878 1368 879
rect 2180 874 2182 880
rect 2526 879 2527 880
rect 2531 879 2532 883
rect 4482 883 4483 887
rect 4487 886 4488 887
rect 4487 884 5301 886
rect 4487 883 4488 884
rect 4482 882 4488 883
rect 2526 878 2532 879
rect 3983 879 3989 880
rect 3983 878 3984 879
rect 3820 876 3984 878
rect 2615 875 2621 876
rect 2615 874 2616 875
rect 2093 872 2182 874
rect 2501 872 2616 874
rect 2186 871 2192 872
rect 262 868 268 869
rect 110 867 116 868
rect 110 863 111 867
rect 115 863 116 867
rect 262 864 263 868
rect 267 864 268 868
rect 262 863 268 864
rect 486 868 492 869
rect 486 864 487 868
rect 491 864 492 868
rect 486 863 492 864
rect 710 868 716 869
rect 710 864 711 868
rect 715 864 716 868
rect 710 863 716 864
rect 934 868 940 869
rect 934 864 935 868
rect 939 864 940 868
rect 934 863 940 864
rect 1158 868 1164 869
rect 1158 864 1159 868
rect 1163 864 1164 868
rect 1158 863 1164 864
rect 1390 868 1396 869
rect 1390 864 1391 868
rect 1395 864 1396 868
rect 1390 863 1396 864
rect 1934 867 1940 868
rect 1934 863 1935 867
rect 1939 863 1940 867
rect 2186 867 2187 871
rect 2191 867 2192 871
rect 2615 871 2616 872
rect 2620 871 2621 875
rect 2894 875 2900 876
rect 2615 870 2621 871
rect 2770 871 2776 872
rect 2186 866 2192 867
rect 2770 867 2771 871
rect 2775 867 2776 871
rect 2894 871 2895 875
rect 2899 874 2900 875
rect 3820 874 3822 876
rect 3983 875 3984 876
rect 3988 875 3989 879
rect 3983 874 3989 875
rect 4090 879 4096 880
rect 4090 875 4091 879
rect 4095 878 4096 879
rect 4119 879 4125 880
rect 4119 878 4120 879
rect 4095 876 4120 878
rect 4095 875 4096 876
rect 4090 874 4096 875
rect 4119 875 4120 876
rect 4124 875 4125 879
rect 4119 874 4125 875
rect 4162 879 4168 880
rect 4162 875 4163 879
rect 4167 878 4168 879
rect 4295 879 4301 880
rect 4295 878 4296 879
rect 4167 876 4296 878
rect 4167 875 4168 876
rect 4162 874 4168 875
rect 4295 875 4296 876
rect 4300 875 4301 879
rect 4295 874 4301 875
rect 4511 879 4517 880
rect 4511 875 4512 879
rect 4516 878 4517 879
rect 4650 879 4656 880
rect 4650 878 4651 879
rect 4516 876 4651 878
rect 4516 875 4517 876
rect 4511 874 4517 875
rect 4650 875 4651 876
rect 4655 875 4656 879
rect 4650 874 4656 875
rect 4767 879 4773 880
rect 4767 875 4768 879
rect 4772 878 4773 879
rect 4938 879 4944 880
rect 4938 878 4939 879
rect 4772 876 4939 878
rect 4772 875 4773 876
rect 4767 874 4773 875
rect 4938 875 4939 876
rect 4943 875 4944 879
rect 4938 874 4944 875
rect 5055 879 5061 880
rect 5055 875 5056 879
rect 5060 878 5061 879
rect 5066 879 5072 880
rect 5066 878 5067 879
rect 5060 876 5067 878
rect 5060 875 5061 876
rect 5055 874 5061 875
rect 5066 875 5067 876
rect 5071 875 5072 879
rect 5299 878 5301 884
rect 5359 879 5365 880
rect 5359 878 5360 879
rect 5299 876 5360 878
rect 5066 874 5072 875
rect 5359 875 5360 876
rect 5364 875 5365 879
rect 5359 874 5365 875
rect 5610 879 5616 880
rect 5610 875 5611 879
rect 5615 878 5616 879
rect 5639 879 5645 880
rect 5639 878 5640 879
rect 5615 876 5640 878
rect 5615 875 5616 876
rect 5610 874 5616 875
rect 5639 875 5640 876
rect 5644 875 5645 879
rect 5639 874 5645 875
rect 2899 872 2993 874
rect 3749 872 3822 874
rect 3838 872 3844 873
rect 5662 872 5668 873
rect 2899 871 2900 872
rect 2894 870 2900 871
rect 3330 871 3336 872
rect 2770 866 2776 867
rect 3330 867 3331 871
rect 3335 867 3336 871
rect 3838 868 3839 872
rect 3843 868 3844 872
rect 3838 867 3844 868
rect 3858 871 3864 872
rect 3858 867 3859 871
rect 3863 867 3864 871
rect 3330 866 3336 867
rect 3858 866 3864 867
rect 3994 871 4000 872
rect 3994 867 3995 871
rect 3999 867 4000 871
rect 3994 866 4000 867
rect 4170 871 4176 872
rect 4170 867 4171 871
rect 4175 867 4176 871
rect 4170 866 4176 867
rect 4386 871 4392 872
rect 4386 867 4387 871
rect 4391 867 4392 871
rect 4386 866 4392 867
rect 4642 871 4648 872
rect 4642 867 4643 871
rect 4647 867 4648 871
rect 4642 866 4648 867
rect 4930 871 4936 872
rect 4930 867 4931 871
rect 4935 867 4936 871
rect 4930 866 4936 867
rect 5234 871 5240 872
rect 5234 867 5235 871
rect 5239 867 5240 871
rect 5234 866 5240 867
rect 5514 871 5520 872
rect 5514 867 5515 871
rect 5519 867 5520 871
rect 5662 868 5663 872
rect 5667 868 5668 872
rect 5662 867 5668 868
rect 5514 866 5520 867
rect 110 862 116 863
rect 1934 862 1940 863
rect 3886 856 3892 857
rect 3838 855 3844 856
rect 3838 851 3839 855
rect 3843 851 3844 855
rect 3886 852 3887 856
rect 3891 852 3892 856
rect 3886 851 3892 852
rect 4022 856 4028 857
rect 4022 852 4023 856
rect 4027 852 4028 856
rect 4022 851 4028 852
rect 4198 856 4204 857
rect 4198 852 4199 856
rect 4203 852 4204 856
rect 4198 851 4204 852
rect 4414 856 4420 857
rect 4414 852 4415 856
rect 4419 852 4420 856
rect 4414 851 4420 852
rect 4670 856 4676 857
rect 4670 852 4671 856
rect 4675 852 4676 856
rect 4670 851 4676 852
rect 4958 856 4964 857
rect 4958 852 4959 856
rect 4963 852 4964 856
rect 4958 851 4964 852
rect 5262 856 5268 857
rect 5262 852 5263 856
rect 5267 852 5268 856
rect 5262 851 5268 852
rect 5542 856 5548 857
rect 5542 852 5543 856
rect 5547 852 5548 856
rect 5542 851 5548 852
rect 5662 855 5668 856
rect 5662 851 5663 855
rect 5667 851 5668 855
rect 3838 850 3844 851
rect 5662 850 5668 851
rect 2770 839 2776 840
rect 2770 835 2771 839
rect 2775 838 2776 839
rect 2775 836 3342 838
rect 2775 835 2776 836
rect 2770 834 2776 835
rect 2119 831 2125 832
rect 2119 827 2120 831
rect 2124 830 2125 831
rect 2186 831 2192 832
rect 2186 830 2187 831
rect 2124 828 2187 830
rect 2124 827 2125 828
rect 2119 826 2125 827
rect 2186 827 2187 828
rect 2191 827 2192 831
rect 2186 826 2192 827
rect 2303 831 2309 832
rect 2303 827 2304 831
rect 2308 830 2309 831
rect 2327 831 2333 832
rect 2327 830 2328 831
rect 2308 828 2328 830
rect 2308 827 2309 828
rect 2303 826 2309 827
rect 2327 827 2328 828
rect 2332 827 2333 831
rect 2327 826 2333 827
rect 2526 831 2533 832
rect 2526 827 2527 831
rect 2532 827 2533 831
rect 2526 826 2533 827
rect 2615 831 2621 832
rect 2615 827 2616 831
rect 2620 830 2621 831
rect 2799 831 2805 832
rect 2799 830 2800 831
rect 2620 828 2800 830
rect 2620 827 2621 828
rect 2615 826 2621 827
rect 2799 827 2800 828
rect 2804 827 2805 831
rect 2799 826 2805 827
rect 3111 831 3117 832
rect 3111 827 3112 831
rect 3116 830 3117 831
rect 3330 831 3336 832
rect 3330 830 3331 831
rect 3116 828 3331 830
rect 3116 827 3117 828
rect 3111 826 3117 827
rect 3330 827 3331 828
rect 3335 827 3336 831
rect 3340 830 3342 836
rect 3447 831 3453 832
rect 3447 830 3448 831
rect 3340 828 3448 830
rect 3330 826 3336 827
rect 3447 827 3448 828
rect 3452 827 3453 831
rect 3447 826 3453 827
rect 3746 831 3752 832
rect 3746 827 3747 831
rect 3751 830 3752 831
rect 3775 831 3781 832
rect 3775 830 3776 831
rect 3751 828 3776 830
rect 3751 827 3752 828
rect 3746 826 3752 827
rect 3775 827 3776 828
rect 3780 827 3781 831
rect 3775 826 3781 827
rect 1974 824 1980 825
rect 3798 824 3804 825
rect 1974 820 1975 824
rect 1979 820 1980 824
rect 1974 819 1980 820
rect 1994 823 2000 824
rect 1994 819 1995 823
rect 1999 819 2000 823
rect 1994 818 2000 819
rect 2178 823 2184 824
rect 2178 819 2179 823
rect 2183 819 2184 823
rect 2178 818 2184 819
rect 2402 823 2408 824
rect 2402 819 2403 823
rect 2407 819 2408 823
rect 2402 818 2408 819
rect 2674 823 2680 824
rect 2674 819 2675 823
rect 2679 819 2680 823
rect 2674 818 2680 819
rect 2986 823 2992 824
rect 2986 819 2987 823
rect 2991 819 2992 823
rect 2986 818 2992 819
rect 3322 823 3328 824
rect 3322 819 3323 823
rect 3327 819 3328 823
rect 3322 818 3328 819
rect 3650 823 3656 824
rect 3650 819 3651 823
rect 3655 819 3656 823
rect 3798 820 3799 824
rect 3803 820 3804 824
rect 3798 819 3804 820
rect 3650 818 3656 819
rect 2022 808 2028 809
rect 1974 807 1980 808
rect 1974 803 1975 807
rect 1979 803 1980 807
rect 2022 804 2023 808
rect 2027 804 2028 808
rect 2022 803 2028 804
rect 2206 808 2212 809
rect 2206 804 2207 808
rect 2211 804 2212 808
rect 2206 803 2212 804
rect 2430 808 2436 809
rect 2430 804 2431 808
rect 2435 804 2436 808
rect 2430 803 2436 804
rect 2702 808 2708 809
rect 2702 804 2703 808
rect 2707 804 2708 808
rect 2702 803 2708 804
rect 3014 808 3020 809
rect 3014 804 3015 808
rect 3019 804 3020 808
rect 3014 803 3020 804
rect 3350 808 3356 809
rect 3350 804 3351 808
rect 3355 804 3356 808
rect 3350 803 3356 804
rect 3678 808 3684 809
rect 3678 804 3679 808
rect 3683 804 3684 808
rect 3678 803 3684 804
rect 3798 807 3804 808
rect 3798 803 3799 807
rect 3803 803 3804 807
rect 1974 802 1980 803
rect 3798 802 3804 803
rect 3838 797 3844 798
rect 5662 797 5668 798
rect 110 793 116 794
rect 1934 793 1940 794
rect 110 789 111 793
rect 115 789 116 793
rect 110 788 116 789
rect 174 792 180 793
rect 174 788 175 792
rect 179 788 180 792
rect 174 787 180 788
rect 430 792 436 793
rect 430 788 431 792
rect 435 788 436 792
rect 430 787 436 788
rect 670 792 676 793
rect 670 788 671 792
rect 675 788 676 792
rect 670 787 676 788
rect 902 792 908 793
rect 902 788 903 792
rect 907 788 908 792
rect 902 787 908 788
rect 1126 792 1132 793
rect 1126 788 1127 792
rect 1131 788 1132 792
rect 1126 787 1132 788
rect 1350 792 1356 793
rect 1350 788 1351 792
rect 1355 788 1356 792
rect 1350 787 1356 788
rect 1574 792 1580 793
rect 1574 788 1575 792
rect 1579 788 1580 792
rect 1934 789 1935 793
rect 1939 789 1940 793
rect 3838 793 3839 797
rect 3843 793 3844 797
rect 3838 792 3844 793
rect 3886 796 3892 797
rect 3886 792 3887 796
rect 3891 792 3892 796
rect 3886 791 3892 792
rect 4022 796 4028 797
rect 4022 792 4023 796
rect 4027 792 4028 796
rect 4022 791 4028 792
rect 4158 796 4164 797
rect 4158 792 4159 796
rect 4163 792 4164 796
rect 4158 791 4164 792
rect 4294 796 4300 797
rect 4294 792 4295 796
rect 4299 792 4300 796
rect 4294 791 4300 792
rect 4430 796 4436 797
rect 4430 792 4431 796
rect 4435 792 4436 796
rect 4430 791 4436 792
rect 4566 796 4572 797
rect 4566 792 4567 796
rect 4571 792 4572 796
rect 4566 791 4572 792
rect 4718 796 4724 797
rect 4718 792 4719 796
rect 4723 792 4724 796
rect 4718 791 4724 792
rect 4894 796 4900 797
rect 4894 792 4895 796
rect 4899 792 4900 796
rect 4894 791 4900 792
rect 5086 796 5092 797
rect 5086 792 5087 796
rect 5091 792 5092 796
rect 5086 791 5092 792
rect 5286 796 5292 797
rect 5286 792 5287 796
rect 5291 792 5292 796
rect 5286 791 5292 792
rect 5486 796 5492 797
rect 5486 792 5487 796
rect 5491 792 5492 796
rect 5662 793 5663 797
rect 5667 793 5668 797
rect 5662 792 5668 793
rect 5486 791 5492 792
rect 1934 788 1940 789
rect 1574 787 1580 788
rect 3858 781 3864 782
rect 3838 780 3844 781
rect 146 777 152 778
rect 110 776 116 777
rect 110 772 111 776
rect 115 772 116 776
rect 146 773 147 777
rect 151 773 152 777
rect 146 772 152 773
rect 402 777 408 778
rect 402 773 403 777
rect 407 773 408 777
rect 402 772 408 773
rect 642 777 648 778
rect 642 773 643 777
rect 647 773 648 777
rect 642 772 648 773
rect 874 777 880 778
rect 874 773 875 777
rect 879 773 880 777
rect 874 772 880 773
rect 1098 777 1104 778
rect 1098 773 1099 777
rect 1103 773 1104 777
rect 1098 772 1104 773
rect 1322 777 1328 778
rect 1322 773 1323 777
rect 1327 773 1328 777
rect 1322 772 1328 773
rect 1546 777 1552 778
rect 1546 773 1547 777
rect 1551 773 1552 777
rect 1546 772 1552 773
rect 1934 776 1940 777
rect 1934 772 1935 776
rect 1939 772 1940 776
rect 3838 776 3839 780
rect 3843 776 3844 780
rect 3858 777 3859 781
rect 3863 777 3864 781
rect 3858 776 3864 777
rect 3994 781 4000 782
rect 3994 777 3995 781
rect 3999 777 4000 781
rect 3994 776 4000 777
rect 4130 781 4136 782
rect 4130 777 4131 781
rect 4135 777 4136 781
rect 4130 776 4136 777
rect 4266 781 4272 782
rect 4266 777 4267 781
rect 4271 777 4272 781
rect 4266 776 4272 777
rect 4402 781 4408 782
rect 4402 777 4403 781
rect 4407 777 4408 781
rect 4402 776 4408 777
rect 4538 781 4544 782
rect 4538 777 4539 781
rect 4543 777 4544 781
rect 4538 776 4544 777
rect 4690 781 4696 782
rect 4690 777 4691 781
rect 4695 777 4696 781
rect 4690 776 4696 777
rect 4866 781 4872 782
rect 4866 777 4867 781
rect 4871 777 4872 781
rect 4866 776 4872 777
rect 5058 781 5064 782
rect 5058 777 5059 781
rect 5063 777 5064 781
rect 5058 776 5064 777
rect 5258 781 5264 782
rect 5258 777 5259 781
rect 5263 777 5264 781
rect 5258 776 5264 777
rect 5458 781 5464 782
rect 5458 777 5459 781
rect 5463 777 5464 781
rect 5458 776 5464 777
rect 5662 780 5668 781
rect 5662 776 5663 780
rect 5667 776 5668 780
rect 3838 775 3844 776
rect 5662 775 5668 776
rect 110 771 116 772
rect 1934 771 1940 772
rect 3954 771 3960 772
rect 270 767 277 768
rect 270 763 271 767
rect 276 763 277 767
rect 270 762 277 763
rect 527 767 536 768
rect 527 763 528 767
rect 535 763 536 767
rect 527 762 536 763
rect 766 767 773 768
rect 766 763 767 767
rect 772 763 773 767
rect 766 762 773 763
rect 999 767 1005 768
rect 999 763 1000 767
rect 1004 766 1005 767
rect 1007 767 1013 768
rect 1007 766 1008 767
rect 1004 764 1008 766
rect 1004 763 1005 764
rect 999 762 1005 763
rect 1007 763 1008 764
rect 1012 763 1013 767
rect 1007 762 1013 763
rect 1062 767 1068 768
rect 1062 763 1063 767
rect 1067 766 1068 767
rect 1223 767 1229 768
rect 1223 766 1224 767
rect 1067 764 1224 766
rect 1067 763 1068 764
rect 1062 762 1068 763
rect 1223 763 1224 764
rect 1228 763 1229 767
rect 1223 762 1229 763
rect 1319 767 1325 768
rect 1319 763 1320 767
rect 1324 766 1325 767
rect 1447 767 1453 768
rect 1447 766 1448 767
rect 1324 764 1448 766
rect 1324 763 1325 764
rect 1319 762 1325 763
rect 1447 763 1448 764
rect 1452 763 1453 767
rect 1447 762 1453 763
rect 1482 767 1488 768
rect 1482 763 1483 767
rect 1487 766 1488 767
rect 1671 767 1677 768
rect 1671 766 1672 767
rect 1487 764 1672 766
rect 1487 763 1488 764
rect 1482 762 1488 763
rect 1671 763 1672 764
rect 1676 763 1677 767
rect 3954 767 3955 771
rect 3959 770 3960 771
rect 3983 771 3989 772
rect 3983 770 3984 771
rect 3959 768 3984 770
rect 3959 767 3960 768
rect 3954 766 3960 767
rect 3983 767 3984 768
rect 3988 767 3989 771
rect 3983 766 3989 767
rect 4119 771 4128 772
rect 4119 767 4120 771
rect 4127 767 4128 771
rect 4119 766 4128 767
rect 4255 771 4264 772
rect 4255 767 4256 771
rect 4263 767 4264 771
rect 4255 766 4264 767
rect 4391 771 4400 772
rect 4391 767 4392 771
rect 4399 767 4400 771
rect 4391 766 4400 767
rect 4527 771 4536 772
rect 4527 767 4528 771
rect 4535 767 4536 771
rect 4527 766 4536 767
rect 4634 771 4640 772
rect 4634 767 4635 771
rect 4639 770 4640 771
rect 4663 771 4669 772
rect 4663 770 4664 771
rect 4639 768 4664 770
rect 4639 767 4640 768
rect 4634 766 4640 767
rect 4663 767 4664 768
rect 4668 767 4669 771
rect 4815 771 4821 772
rect 4815 770 4816 771
rect 4663 766 4669 767
rect 4672 768 4816 770
rect 1671 762 1677 763
rect 4274 763 4280 764
rect 4274 759 4275 763
rect 4279 762 4280 763
rect 4672 762 4674 768
rect 4815 767 4816 768
rect 4820 767 4821 771
rect 4815 766 4821 767
rect 4842 771 4848 772
rect 4842 767 4843 771
rect 4847 770 4848 771
rect 4991 771 4997 772
rect 4991 770 4992 771
rect 4847 768 4992 770
rect 4847 767 4848 768
rect 4842 766 4848 767
rect 4991 767 4992 768
rect 4996 767 4997 771
rect 4991 766 4997 767
rect 5183 771 5189 772
rect 5183 767 5184 771
rect 5188 770 5189 771
rect 5218 771 5224 772
rect 5218 770 5219 771
rect 5188 768 5219 770
rect 5188 767 5189 768
rect 5183 766 5189 767
rect 5218 767 5219 768
rect 5223 767 5224 771
rect 5383 771 5389 772
rect 5383 770 5384 771
rect 5218 766 5224 767
rect 5299 768 5384 770
rect 4279 760 4674 762
rect 4962 763 4968 764
rect 4279 759 4280 760
rect 4274 758 4280 759
rect 4962 759 4963 763
rect 4967 762 4968 763
rect 5299 762 5301 768
rect 5383 767 5384 768
rect 5388 767 5389 771
rect 5383 766 5389 767
rect 5554 771 5560 772
rect 5554 767 5555 771
rect 5559 770 5560 771
rect 5583 771 5589 772
rect 5583 770 5584 771
rect 5559 768 5584 770
rect 5559 767 5560 768
rect 5554 766 5560 767
rect 5583 767 5584 768
rect 5588 767 5589 771
rect 5583 766 5589 767
rect 4967 760 5301 762
rect 4967 759 4968 760
rect 4962 758 4968 759
rect 3954 731 3960 732
rect 242 727 248 728
rect 242 723 243 727
rect 247 723 248 727
rect 242 722 248 723
rect 498 727 504 728
rect 498 723 499 727
rect 503 723 504 727
rect 498 722 504 723
rect 530 727 536 728
rect 530 723 531 727
rect 535 726 536 727
rect 1062 727 1068 728
rect 1062 726 1063 727
rect 535 724 649 726
rect 973 724 1063 726
rect 535 723 536 724
rect 530 722 536 723
rect 1062 723 1063 724
rect 1067 723 1068 727
rect 1319 727 1325 728
rect 1319 726 1320 727
rect 1197 724 1320 726
rect 1062 722 1068 723
rect 1319 723 1320 724
rect 1324 723 1325 727
rect 1482 727 1488 728
rect 1482 726 1483 727
rect 1421 724 1483 726
rect 1319 722 1325 723
rect 1482 723 1483 724
rect 1487 723 1488 727
rect 1482 722 1488 723
rect 1490 727 1496 728
rect 1490 723 1491 727
rect 1495 726 1496 727
rect 3954 727 3955 731
rect 3959 727 3960 731
rect 3954 726 3960 727
rect 4090 731 4096 732
rect 4090 727 4091 731
rect 4095 727 4096 731
rect 4090 726 4096 727
rect 4122 731 4128 732
rect 4122 727 4123 731
rect 4127 730 4128 731
rect 4258 731 4264 732
rect 4127 728 4137 730
rect 4127 727 4128 728
rect 4122 726 4128 727
rect 4258 727 4259 731
rect 4263 730 4264 731
rect 4394 731 4400 732
rect 4263 728 4273 730
rect 4263 727 4264 728
rect 4258 726 4264 727
rect 4394 727 4395 731
rect 4399 730 4400 731
rect 4530 731 4536 732
rect 4399 728 4409 730
rect 4399 727 4400 728
rect 4394 726 4400 727
rect 4530 727 4531 731
rect 4535 730 4536 731
rect 4842 731 4848 732
rect 4842 730 4843 731
rect 4535 728 4545 730
rect 4789 728 4843 730
rect 4535 727 4536 728
rect 4530 726 4536 727
rect 4842 727 4843 728
rect 4847 727 4848 731
rect 4842 726 4848 727
rect 4962 731 4968 732
rect 4962 727 4963 731
rect 4967 727 4968 731
rect 4962 726 4968 727
rect 5066 731 5072 732
rect 5066 727 5067 731
rect 5071 727 5072 731
rect 5066 726 5072 727
rect 5218 731 5224 732
rect 5218 727 5219 731
rect 5223 730 5224 731
rect 5554 731 5560 732
rect 5223 728 5265 730
rect 5223 727 5224 728
rect 5218 726 5224 727
rect 5554 727 5555 731
rect 5559 727 5560 731
rect 5554 726 5560 727
rect 1495 724 1553 726
rect 1495 723 1496 724
rect 1490 722 1496 723
rect 306 695 312 696
rect 306 694 307 695
rect 229 692 307 694
rect 306 691 307 692
rect 311 691 312 695
rect 766 695 772 696
rect 306 690 312 691
rect 410 691 416 692
rect 410 687 411 691
rect 415 687 416 691
rect 410 686 416 687
rect 618 691 624 692
rect 618 687 619 691
rect 623 687 624 691
rect 766 691 767 695
rect 771 691 772 695
rect 1007 695 1013 696
rect 766 690 772 691
rect 914 691 920 692
rect 618 686 624 687
rect 914 687 915 691
rect 919 687 920 691
rect 1007 691 1008 695
rect 1012 694 1013 695
rect 3991 695 3997 696
rect 3991 694 3992 695
rect 1012 692 1089 694
rect 3957 692 3992 694
rect 1012 691 1013 692
rect 1007 690 1013 691
rect 1266 691 1272 692
rect 914 686 920 687
rect 1266 687 1267 691
rect 1271 687 1272 691
rect 1266 686 1272 687
rect 1434 691 1440 692
rect 1434 687 1435 691
rect 1439 687 1440 691
rect 1434 686 1440 687
rect 1602 691 1608 692
rect 1602 687 1603 691
rect 1607 687 1608 691
rect 1602 686 1608 687
rect 1778 691 1784 692
rect 1778 687 1779 691
rect 1783 687 1784 691
rect 3991 691 3992 692
rect 3996 691 3997 695
rect 4634 695 4640 696
rect 3991 690 3997 691
rect 4002 691 4008 692
rect 1778 686 1784 687
rect 4002 687 4003 691
rect 4007 687 4008 691
rect 4002 686 4008 687
rect 4138 691 4144 692
rect 4138 687 4139 691
rect 4143 687 4144 691
rect 4138 686 4144 687
rect 4274 691 4280 692
rect 4274 687 4275 691
rect 4279 687 4280 691
rect 4274 686 4280 687
rect 4410 691 4416 692
rect 4410 687 4411 691
rect 4415 687 4416 691
rect 4634 691 4635 695
rect 4639 691 4640 695
rect 5610 695 5616 696
rect 4634 690 4640 691
rect 4706 691 4712 692
rect 4410 686 4416 687
rect 4706 687 4707 691
rect 4711 687 4712 691
rect 4706 686 4712 687
rect 4898 691 4904 692
rect 4898 687 4899 691
rect 4903 687 4904 691
rect 4898 686 4904 687
rect 5106 691 5112 692
rect 5106 687 5107 691
rect 5111 687 5112 691
rect 5106 686 5112 687
rect 5322 691 5328 692
rect 5322 687 5323 691
rect 5327 687 5328 691
rect 5610 691 5611 695
rect 5615 691 5616 695
rect 5610 690 5616 691
rect 5322 686 5328 687
rect 618 659 624 660
rect 618 655 619 659
rect 623 658 624 659
rect 3991 659 3997 660
rect 623 656 926 658
rect 623 655 624 656
rect 618 654 624 655
rect 242 651 248 652
rect 242 647 243 651
rect 247 650 248 651
rect 255 651 261 652
rect 255 650 256 651
rect 247 648 256 650
rect 247 647 248 648
rect 242 646 248 647
rect 255 647 256 648
rect 260 647 261 651
rect 255 646 261 647
rect 306 651 312 652
rect 306 647 307 651
rect 311 650 312 651
rect 439 651 445 652
rect 439 650 440 651
rect 311 648 440 650
rect 311 647 312 648
rect 306 646 312 647
rect 439 647 440 648
rect 444 647 445 651
rect 439 646 445 647
rect 646 651 653 652
rect 646 647 647 651
rect 652 647 653 651
rect 646 646 653 647
rect 847 651 853 652
rect 847 647 848 651
rect 852 650 853 651
rect 914 651 920 652
rect 914 650 915 651
rect 852 648 915 650
rect 852 647 853 648
rect 847 646 853 647
rect 914 647 915 648
rect 919 647 920 651
rect 924 650 926 656
rect 3991 655 3992 659
rect 3996 658 3997 659
rect 3996 656 4461 658
rect 3996 655 3997 656
rect 3991 654 3997 655
rect 1031 651 1037 652
rect 1031 650 1032 651
rect 924 648 1032 650
rect 914 646 920 647
rect 1031 647 1032 648
rect 1036 647 1037 651
rect 1031 646 1037 647
rect 1207 651 1213 652
rect 1207 647 1208 651
rect 1212 650 1213 651
rect 1266 651 1272 652
rect 1266 650 1267 651
rect 1212 648 1267 650
rect 1212 647 1213 648
rect 1207 646 1213 647
rect 1266 647 1267 648
rect 1271 647 1272 651
rect 1266 646 1272 647
rect 1383 651 1389 652
rect 1383 647 1384 651
rect 1388 650 1389 651
rect 1434 651 1440 652
rect 1434 650 1435 651
rect 1388 648 1435 650
rect 1388 647 1389 648
rect 1383 646 1389 647
rect 1434 647 1435 648
rect 1439 647 1440 651
rect 1434 646 1440 647
rect 1551 651 1557 652
rect 1551 647 1552 651
rect 1556 650 1557 651
rect 1602 651 1608 652
rect 1602 650 1603 651
rect 1556 648 1603 650
rect 1556 647 1557 648
rect 1551 646 1557 647
rect 1602 647 1603 648
rect 1607 647 1608 651
rect 1602 646 1608 647
rect 1719 651 1725 652
rect 1719 647 1720 651
rect 1724 650 1725 651
rect 1778 651 1784 652
rect 1778 650 1779 651
rect 1724 648 1779 650
rect 1724 647 1725 648
rect 1719 646 1725 647
rect 1778 647 1779 648
rect 1783 647 1784 651
rect 1778 646 1784 647
rect 1894 651 1901 652
rect 1894 647 1895 651
rect 1900 647 1901 651
rect 1894 646 1901 647
rect 3954 651 3960 652
rect 3954 647 3955 651
rect 3959 650 3960 651
rect 3983 651 3989 652
rect 3983 650 3984 651
rect 3959 648 3984 650
rect 3959 647 3960 648
rect 3954 646 3960 647
rect 3983 647 3984 648
rect 3988 647 3989 651
rect 3983 646 3989 647
rect 4119 651 4125 652
rect 4119 647 4120 651
rect 4124 650 4125 651
rect 4138 651 4144 652
rect 4138 650 4139 651
rect 4124 648 4139 650
rect 4124 647 4125 648
rect 4119 646 4125 647
rect 4138 647 4139 648
rect 4143 647 4144 651
rect 4138 646 4144 647
rect 4255 651 4261 652
rect 4255 647 4256 651
rect 4260 650 4261 651
rect 4274 651 4280 652
rect 4274 650 4275 651
rect 4260 648 4275 650
rect 4260 647 4261 648
rect 4255 646 4261 647
rect 4274 647 4275 648
rect 4279 647 4280 651
rect 4274 646 4280 647
rect 4391 651 4397 652
rect 4391 647 4392 651
rect 4396 650 4397 651
rect 4410 651 4416 652
rect 4410 650 4411 651
rect 4396 648 4411 650
rect 4396 647 4397 648
rect 4391 646 4397 647
rect 4410 647 4411 648
rect 4415 647 4416 651
rect 4459 650 4461 656
rect 4527 651 4533 652
rect 4527 650 4528 651
rect 4459 648 4528 650
rect 4410 646 4416 647
rect 4527 647 4528 648
rect 4532 647 4533 651
rect 4527 646 4533 647
rect 4663 651 4669 652
rect 4663 647 4664 651
rect 4668 650 4669 651
rect 4706 651 4712 652
rect 4706 650 4707 651
rect 4668 648 4707 650
rect 4668 647 4669 648
rect 4663 646 4669 647
rect 4706 647 4707 648
rect 4711 647 4712 651
rect 4706 646 4712 647
rect 4823 651 4829 652
rect 4823 647 4824 651
rect 4828 650 4829 651
rect 4898 651 4904 652
rect 4898 650 4899 651
rect 4828 648 4899 650
rect 4828 647 4829 648
rect 4823 646 4829 647
rect 4898 647 4899 648
rect 4903 647 4904 651
rect 4898 646 4904 647
rect 5015 651 5021 652
rect 5015 647 5016 651
rect 5020 650 5021 651
rect 5106 651 5112 652
rect 5106 650 5107 651
rect 5020 648 5107 650
rect 5020 647 5021 648
rect 5015 646 5021 647
rect 5106 647 5107 648
rect 5111 647 5112 651
rect 5106 646 5112 647
rect 5223 651 5229 652
rect 5223 647 5224 651
rect 5228 650 5229 651
rect 5322 651 5328 652
rect 5322 650 5323 651
rect 5228 648 5323 650
rect 5228 647 5229 648
rect 5223 646 5229 647
rect 5322 647 5323 648
rect 5327 647 5328 651
rect 5322 646 5328 647
rect 5366 651 5372 652
rect 5366 647 5367 651
rect 5371 650 5372 651
rect 5439 651 5445 652
rect 5439 650 5440 651
rect 5371 648 5440 650
rect 5371 647 5372 648
rect 5366 646 5372 647
rect 5439 647 5440 648
rect 5444 647 5445 651
rect 5439 646 5445 647
rect 5554 651 5560 652
rect 5554 647 5555 651
rect 5559 650 5560 651
rect 5639 651 5645 652
rect 5639 650 5640 651
rect 5559 648 5640 650
rect 5559 647 5560 648
rect 5554 646 5560 647
rect 5639 647 5640 648
rect 5644 647 5645 651
rect 5639 646 5645 647
rect 110 644 116 645
rect 1934 644 1940 645
rect 110 640 111 644
rect 115 640 116 644
rect 110 639 116 640
rect 130 643 136 644
rect 130 639 131 643
rect 135 639 136 643
rect 130 638 136 639
rect 314 643 320 644
rect 314 639 315 643
rect 319 639 320 643
rect 314 638 320 639
rect 522 643 528 644
rect 522 639 523 643
rect 527 639 528 643
rect 522 638 528 639
rect 722 643 728 644
rect 722 639 723 643
rect 727 639 728 643
rect 722 638 728 639
rect 906 643 912 644
rect 906 639 907 643
rect 911 639 912 643
rect 906 638 912 639
rect 1082 643 1088 644
rect 1082 639 1083 643
rect 1087 639 1088 643
rect 1082 638 1088 639
rect 1258 643 1264 644
rect 1258 639 1259 643
rect 1263 639 1264 643
rect 1258 638 1264 639
rect 1426 643 1432 644
rect 1426 639 1427 643
rect 1431 639 1432 643
rect 1426 638 1432 639
rect 1594 643 1600 644
rect 1594 639 1595 643
rect 1599 639 1600 643
rect 1594 638 1600 639
rect 1770 643 1776 644
rect 1770 639 1771 643
rect 1775 639 1776 643
rect 1934 640 1935 644
rect 1939 640 1940 644
rect 1934 639 1940 640
rect 3838 644 3844 645
rect 5662 644 5668 645
rect 3838 640 3839 644
rect 3843 640 3844 644
rect 3838 639 3844 640
rect 3858 643 3864 644
rect 3858 639 3859 643
rect 3863 639 3864 643
rect 1770 638 1776 639
rect 3858 638 3864 639
rect 3994 643 4000 644
rect 3994 639 3995 643
rect 3999 639 4000 643
rect 3994 638 4000 639
rect 4130 643 4136 644
rect 4130 639 4131 643
rect 4135 639 4136 643
rect 4130 638 4136 639
rect 4266 643 4272 644
rect 4266 639 4267 643
rect 4271 639 4272 643
rect 4266 638 4272 639
rect 4402 643 4408 644
rect 4402 639 4403 643
rect 4407 639 4408 643
rect 4402 638 4408 639
rect 4538 643 4544 644
rect 4538 639 4539 643
rect 4543 639 4544 643
rect 4538 638 4544 639
rect 4698 643 4704 644
rect 4698 639 4699 643
rect 4703 639 4704 643
rect 4698 638 4704 639
rect 4890 643 4896 644
rect 4890 639 4891 643
rect 4895 639 4896 643
rect 4890 638 4896 639
rect 5098 643 5104 644
rect 5098 639 5099 643
rect 5103 639 5104 643
rect 5098 638 5104 639
rect 5314 643 5320 644
rect 5314 639 5315 643
rect 5319 639 5320 643
rect 5314 638 5320 639
rect 5514 643 5520 644
rect 5514 639 5515 643
rect 5519 639 5520 643
rect 5662 640 5663 644
rect 5667 640 5668 644
rect 5662 639 5668 640
rect 5514 638 5520 639
rect 158 628 164 629
rect 110 627 116 628
rect 110 623 111 627
rect 115 623 116 627
rect 158 624 159 628
rect 163 624 164 628
rect 158 623 164 624
rect 342 628 348 629
rect 342 624 343 628
rect 347 624 348 628
rect 342 623 348 624
rect 550 628 556 629
rect 550 624 551 628
rect 555 624 556 628
rect 550 623 556 624
rect 750 628 756 629
rect 750 624 751 628
rect 755 624 756 628
rect 750 623 756 624
rect 934 628 940 629
rect 934 624 935 628
rect 939 624 940 628
rect 934 623 940 624
rect 1110 628 1116 629
rect 1110 624 1111 628
rect 1115 624 1116 628
rect 1110 623 1116 624
rect 1286 628 1292 629
rect 1286 624 1287 628
rect 1291 624 1292 628
rect 1286 623 1292 624
rect 1454 628 1460 629
rect 1454 624 1455 628
rect 1459 624 1460 628
rect 1454 623 1460 624
rect 1622 628 1628 629
rect 1622 624 1623 628
rect 1627 624 1628 628
rect 1622 623 1628 624
rect 1798 628 1804 629
rect 3886 628 3892 629
rect 1798 624 1799 628
rect 1803 624 1804 628
rect 1798 623 1804 624
rect 1934 627 1940 628
rect 1934 623 1935 627
rect 1939 623 1940 627
rect 110 622 116 623
rect 1934 622 1940 623
rect 3838 627 3844 628
rect 3838 623 3839 627
rect 3843 623 3844 627
rect 3886 624 3887 628
rect 3891 624 3892 628
rect 3886 623 3892 624
rect 4022 628 4028 629
rect 4022 624 4023 628
rect 4027 624 4028 628
rect 4022 623 4028 624
rect 4158 628 4164 629
rect 4158 624 4159 628
rect 4163 624 4164 628
rect 4158 623 4164 624
rect 4294 628 4300 629
rect 4294 624 4295 628
rect 4299 624 4300 628
rect 4294 623 4300 624
rect 4430 628 4436 629
rect 4430 624 4431 628
rect 4435 624 4436 628
rect 4430 623 4436 624
rect 4566 628 4572 629
rect 4566 624 4567 628
rect 4571 624 4572 628
rect 4566 623 4572 624
rect 4726 628 4732 629
rect 4726 624 4727 628
rect 4731 624 4732 628
rect 4726 623 4732 624
rect 4918 628 4924 629
rect 4918 624 4919 628
rect 4923 624 4924 628
rect 4918 623 4924 624
rect 5126 628 5132 629
rect 5126 624 5127 628
rect 5131 624 5132 628
rect 5126 623 5132 624
rect 5342 628 5348 629
rect 5342 624 5343 628
rect 5347 624 5348 628
rect 5342 623 5348 624
rect 5542 628 5548 629
rect 5542 624 5543 628
rect 5547 624 5548 628
rect 5542 623 5548 624
rect 5662 627 5668 628
rect 5662 623 5663 627
rect 5667 623 5668 627
rect 3838 622 3844 623
rect 5662 622 5668 623
rect 110 569 116 570
rect 1934 569 1940 570
rect 110 565 111 569
rect 115 565 116 569
rect 110 564 116 565
rect 158 568 164 569
rect 158 564 159 568
rect 163 564 164 568
rect 158 563 164 564
rect 374 568 380 569
rect 374 564 375 568
rect 379 564 380 568
rect 374 563 380 564
rect 598 568 604 569
rect 598 564 599 568
rect 603 564 604 568
rect 598 563 604 564
rect 806 568 812 569
rect 806 564 807 568
rect 811 564 812 568
rect 806 563 812 564
rect 998 568 1004 569
rect 998 564 999 568
rect 1003 564 1004 568
rect 998 563 1004 564
rect 1174 568 1180 569
rect 1174 564 1175 568
rect 1179 564 1180 568
rect 1174 563 1180 564
rect 1342 568 1348 569
rect 1342 564 1343 568
rect 1347 564 1348 568
rect 1342 563 1348 564
rect 1510 568 1516 569
rect 1510 564 1511 568
rect 1515 564 1516 568
rect 1510 563 1516 564
rect 1670 568 1676 569
rect 1670 564 1671 568
rect 1675 564 1676 568
rect 1670 563 1676 564
rect 1814 568 1820 569
rect 1814 564 1815 568
rect 1819 564 1820 568
rect 1934 565 1935 569
rect 1939 565 1940 569
rect 1934 564 1940 565
rect 3838 569 3844 570
rect 5662 569 5668 570
rect 3838 565 3839 569
rect 3843 565 3844 569
rect 3838 564 3844 565
rect 3886 568 3892 569
rect 3886 564 3887 568
rect 3891 564 3892 568
rect 1814 563 1820 564
rect 3886 563 3892 564
rect 4070 568 4076 569
rect 4070 564 4071 568
rect 4075 564 4076 568
rect 4070 563 4076 564
rect 4310 568 4316 569
rect 4310 564 4311 568
rect 4315 564 4316 568
rect 4310 563 4316 564
rect 4574 568 4580 569
rect 4574 564 4575 568
rect 4579 564 4580 568
rect 4574 563 4580 564
rect 4854 568 4860 569
rect 4854 564 4855 568
rect 4859 564 4860 568
rect 4854 563 4860 564
rect 5150 568 5156 569
rect 5150 564 5151 568
rect 5155 564 5156 568
rect 5150 563 5156 564
rect 5446 568 5452 569
rect 5446 564 5447 568
rect 5451 564 5452 568
rect 5662 565 5663 569
rect 5667 565 5668 569
rect 5662 564 5668 565
rect 5446 563 5452 564
rect 130 553 136 554
rect 110 552 116 553
rect 110 548 111 552
rect 115 548 116 552
rect 130 549 131 553
rect 135 549 136 553
rect 130 548 136 549
rect 346 553 352 554
rect 346 549 347 553
rect 351 549 352 553
rect 346 548 352 549
rect 570 553 576 554
rect 570 549 571 553
rect 575 549 576 553
rect 570 548 576 549
rect 778 553 784 554
rect 778 549 779 553
rect 783 549 784 553
rect 778 548 784 549
rect 970 553 976 554
rect 970 549 971 553
rect 975 549 976 553
rect 970 548 976 549
rect 1146 553 1152 554
rect 1146 549 1147 553
rect 1151 549 1152 553
rect 1146 548 1152 549
rect 1314 553 1320 554
rect 1314 549 1315 553
rect 1319 549 1320 553
rect 1314 548 1320 549
rect 1482 553 1488 554
rect 1482 549 1483 553
rect 1487 549 1488 553
rect 1482 548 1488 549
rect 1642 553 1648 554
rect 1642 549 1643 553
rect 1647 549 1648 553
rect 1642 548 1648 549
rect 1786 553 1792 554
rect 3858 553 3864 554
rect 1786 549 1787 553
rect 1791 549 1792 553
rect 1786 548 1792 549
rect 1934 552 1940 553
rect 1934 548 1935 552
rect 1939 548 1940 552
rect 3838 552 3844 553
rect 110 547 116 548
rect 1934 547 1940 548
rect 1974 549 1980 550
rect 3798 549 3804 550
rect 1974 545 1975 549
rect 1979 545 1980 549
rect 1974 544 1980 545
rect 3134 548 3140 549
rect 3134 544 3135 548
rect 3139 544 3140 548
rect 254 543 261 544
rect 254 539 255 543
rect 260 539 261 543
rect 254 538 261 539
rect 410 543 416 544
rect 410 539 411 543
rect 415 542 416 543
rect 471 543 477 544
rect 471 542 472 543
rect 415 540 472 542
rect 415 539 416 540
rect 410 538 416 539
rect 471 539 472 540
rect 476 539 477 543
rect 471 538 477 539
rect 695 543 701 544
rect 695 539 696 543
rect 700 542 701 543
rect 742 543 748 544
rect 742 542 743 543
rect 700 540 743 542
rect 700 539 701 540
rect 695 538 701 539
rect 742 539 743 540
rect 747 539 748 543
rect 742 538 748 539
rect 903 543 912 544
rect 903 539 904 543
rect 911 539 912 543
rect 903 538 912 539
rect 1095 543 1101 544
rect 1095 539 1096 543
rect 1100 542 1101 543
rect 1119 543 1125 544
rect 1119 542 1120 543
rect 1100 540 1120 542
rect 1100 539 1101 540
rect 1095 538 1101 539
rect 1119 539 1120 540
rect 1124 539 1125 543
rect 1119 538 1125 539
rect 1271 543 1280 544
rect 1271 539 1272 543
rect 1279 539 1280 543
rect 1271 538 1280 539
rect 1439 543 1448 544
rect 1439 539 1440 543
rect 1447 539 1448 543
rect 1439 538 1448 539
rect 1607 543 1613 544
rect 1607 539 1608 543
rect 1612 542 1613 543
rect 1630 543 1636 544
rect 1630 542 1631 543
rect 1612 540 1631 542
rect 1612 539 1613 540
rect 1607 538 1613 539
rect 1630 539 1631 540
rect 1635 539 1636 543
rect 1630 538 1636 539
rect 1767 543 1776 544
rect 1767 539 1768 543
rect 1775 539 1776 543
rect 1767 538 1776 539
rect 1882 543 1888 544
rect 1882 539 1883 543
rect 1887 542 1888 543
rect 1911 543 1917 544
rect 3134 543 3140 544
rect 3270 548 3276 549
rect 3270 544 3271 548
rect 3275 544 3276 548
rect 3270 543 3276 544
rect 3406 548 3412 549
rect 3406 544 3407 548
rect 3411 544 3412 548
rect 3406 543 3412 544
rect 3542 548 3548 549
rect 3542 544 3543 548
rect 3547 544 3548 548
rect 3542 543 3548 544
rect 3678 548 3684 549
rect 3678 544 3679 548
rect 3683 544 3684 548
rect 3798 545 3799 549
rect 3803 545 3804 549
rect 3838 548 3839 552
rect 3843 548 3844 552
rect 3858 549 3859 553
rect 3863 549 3864 553
rect 3858 548 3864 549
rect 4042 553 4048 554
rect 4042 549 4043 553
rect 4047 549 4048 553
rect 4042 548 4048 549
rect 4282 553 4288 554
rect 4282 549 4283 553
rect 4287 549 4288 553
rect 4282 548 4288 549
rect 4546 553 4552 554
rect 4546 549 4547 553
rect 4551 549 4552 553
rect 4546 548 4552 549
rect 4826 553 4832 554
rect 4826 549 4827 553
rect 4831 549 4832 553
rect 4826 548 4832 549
rect 5122 553 5128 554
rect 5122 549 5123 553
rect 5127 549 5128 553
rect 5122 548 5128 549
rect 5418 553 5424 554
rect 5418 549 5419 553
rect 5423 549 5424 553
rect 5418 548 5424 549
rect 5662 552 5668 553
rect 5662 548 5663 552
rect 5667 548 5668 552
rect 3838 547 3844 548
rect 5662 547 5668 548
rect 3798 544 3804 545
rect 3678 543 3684 544
rect 3983 543 3989 544
rect 1911 542 1912 543
rect 1887 540 1912 542
rect 1887 539 1888 540
rect 1882 538 1888 539
rect 1911 539 1912 540
rect 1916 539 1917 543
rect 1911 538 1917 539
rect 3983 539 3984 543
rect 3988 542 3989 543
rect 4002 543 4008 544
rect 4002 542 4003 543
rect 3988 540 4003 542
rect 3988 539 3989 540
rect 3983 538 3989 539
rect 4002 539 4003 540
rect 4007 539 4008 543
rect 4002 538 4008 539
rect 4167 543 4176 544
rect 4167 539 4168 543
rect 4175 539 4176 543
rect 4167 538 4176 539
rect 4407 543 4413 544
rect 4407 539 4408 543
rect 4412 542 4413 543
rect 4431 543 4437 544
rect 4431 542 4432 543
rect 4412 540 4432 542
rect 4412 539 4413 540
rect 4407 538 4413 539
rect 4431 539 4432 540
rect 4436 539 4437 543
rect 4431 538 4437 539
rect 4671 543 4680 544
rect 4671 539 4672 543
rect 4679 539 4680 543
rect 4671 538 4680 539
rect 4951 543 4957 544
rect 4951 539 4952 543
rect 4956 542 4957 543
rect 4999 543 5005 544
rect 4999 542 5000 543
rect 4956 540 5000 542
rect 4956 539 4957 540
rect 4951 538 4957 539
rect 4999 539 5000 540
rect 5004 539 5005 543
rect 5247 543 5253 544
rect 5247 542 5248 543
rect 4999 538 5005 539
rect 5008 540 5248 542
rect 4634 535 4640 536
rect 3106 533 3112 534
rect 1974 532 1980 533
rect 1974 528 1975 532
rect 1979 528 1980 532
rect 3106 529 3107 533
rect 3111 529 3112 533
rect 3106 528 3112 529
rect 3242 533 3248 534
rect 3242 529 3243 533
rect 3247 529 3248 533
rect 3242 528 3248 529
rect 3378 533 3384 534
rect 3378 529 3379 533
rect 3383 529 3384 533
rect 3378 528 3384 529
rect 3514 533 3520 534
rect 3514 529 3515 533
rect 3519 529 3520 533
rect 3514 528 3520 529
rect 3650 533 3656 534
rect 3650 529 3651 533
rect 3655 529 3656 533
rect 3650 528 3656 529
rect 3798 532 3804 533
rect 3798 528 3799 532
rect 3803 528 3804 532
rect 4634 531 4635 535
rect 4639 534 4640 535
rect 5008 534 5010 540
rect 5247 539 5248 540
rect 5252 539 5253 543
rect 5247 538 5253 539
rect 5542 543 5549 544
rect 5542 539 5543 543
rect 5548 539 5549 543
rect 5542 538 5549 539
rect 4639 532 5010 534
rect 4639 531 4640 532
rect 4634 530 4640 531
rect 1974 527 1980 528
rect 3798 527 3804 528
rect 3231 523 3240 524
rect 3231 519 3232 523
rect 3239 519 3240 523
rect 3231 518 3240 519
rect 3367 523 3376 524
rect 3367 519 3368 523
rect 3375 519 3376 523
rect 3367 518 3376 519
rect 3503 523 3512 524
rect 3503 519 3504 523
rect 3511 519 3512 523
rect 3503 518 3512 519
rect 3639 523 3648 524
rect 3639 519 3640 523
rect 3647 519 3648 523
rect 3639 518 3648 519
rect 3775 523 3784 524
rect 3775 519 3776 523
rect 3783 519 3784 523
rect 3775 518 3784 519
rect 226 503 232 504
rect 226 499 227 503
rect 231 499 232 503
rect 226 498 232 499
rect 254 503 260 504
rect 254 499 255 503
rect 259 502 260 503
rect 646 503 652 504
rect 259 500 353 502
rect 259 499 260 500
rect 254 498 260 499
rect 646 499 647 503
rect 651 499 652 503
rect 646 498 652 499
rect 742 503 748 504
rect 742 499 743 503
rect 747 502 748 503
rect 906 503 912 504
rect 747 500 785 502
rect 747 499 748 500
rect 742 498 748 499
rect 906 499 907 503
rect 911 502 912 503
rect 1274 503 1280 504
rect 911 500 977 502
rect 911 499 912 500
rect 906 498 912 499
rect 1244 494 1246 501
rect 1274 499 1275 503
rect 1279 502 1280 503
rect 1442 503 1448 504
rect 1279 500 1321 502
rect 1279 499 1280 500
rect 1274 498 1280 499
rect 1442 499 1443 503
rect 1447 502 1448 503
rect 1630 503 1636 504
rect 1447 500 1489 502
rect 1447 499 1448 500
rect 1442 498 1448 499
rect 1630 499 1631 503
rect 1635 502 1636 503
rect 1770 503 1776 504
rect 1635 500 1649 502
rect 1635 499 1636 500
rect 1630 498 1636 499
rect 1770 499 1771 503
rect 1775 502 1776 503
rect 3778 503 3784 504
rect 1775 500 1793 502
rect 1775 499 1776 500
rect 1770 498 1776 499
rect 3778 499 3779 503
rect 3783 502 3784 503
rect 4170 503 4176 504
rect 3783 500 3865 502
rect 3783 499 3784 500
rect 3778 498 3784 499
rect 1894 495 1900 496
rect 1894 494 1895 495
rect 1244 492 1895 494
rect 1894 491 1895 492
rect 1899 491 1900 495
rect 1894 490 1900 491
rect 4140 486 4142 501
rect 4170 499 4171 503
rect 4175 502 4176 503
rect 4431 503 4437 504
rect 4175 500 4289 502
rect 4175 499 4176 500
rect 4170 498 4176 499
rect 4431 499 4432 503
rect 4436 502 4437 503
rect 4674 503 4680 504
rect 4436 500 4553 502
rect 4436 499 4437 500
rect 4431 498 4437 499
rect 4674 499 4675 503
rect 4679 502 4680 503
rect 4999 503 5005 504
rect 4679 500 4833 502
rect 4679 499 4680 500
rect 4674 498 4680 499
rect 4999 499 5000 503
rect 5004 502 5005 503
rect 5394 503 5400 504
rect 5004 500 5129 502
rect 5004 499 5005 500
rect 4999 498 5005 499
rect 5394 499 5395 503
rect 5399 502 5400 503
rect 5399 500 5425 502
rect 5399 499 5400 500
rect 5394 498 5400 499
rect 5366 487 5372 488
rect 5366 486 5367 487
rect 4140 484 5367 486
rect 3202 483 3208 484
rect 3202 479 3203 483
rect 3207 479 3208 483
rect 3202 478 3208 479
rect 3234 483 3240 484
rect 3234 479 3235 483
rect 3239 482 3240 483
rect 3370 483 3376 484
rect 3239 480 3249 482
rect 3239 479 3240 480
rect 3234 478 3240 479
rect 3370 479 3371 483
rect 3375 482 3376 483
rect 3506 483 3512 484
rect 3375 480 3385 482
rect 3375 479 3376 480
rect 3370 478 3376 479
rect 3506 479 3507 483
rect 3511 482 3512 483
rect 3642 483 3648 484
rect 3511 480 3521 482
rect 3511 479 3512 480
rect 3506 478 3512 479
rect 3642 479 3643 483
rect 3647 482 3648 483
rect 5366 483 5367 484
rect 5371 483 5372 487
rect 5366 482 5372 483
rect 3647 480 3657 482
rect 3647 479 3648 480
rect 3642 478 3648 479
rect 1119 471 1125 472
rect 250 467 256 468
rect 250 463 251 467
rect 255 463 256 467
rect 250 462 256 463
rect 578 467 584 468
rect 578 463 579 467
rect 583 463 584 467
rect 578 462 584 463
rect 906 467 912 468
rect 906 463 907 467
rect 911 463 912 467
rect 1119 467 1120 471
rect 1124 470 1125 471
rect 1882 471 1888 472
rect 1124 468 1145 470
rect 1124 467 1125 468
rect 1119 466 1125 467
rect 1482 467 1488 468
rect 906 462 912 463
rect 1482 463 1483 467
rect 1487 463 1488 467
rect 1882 467 1883 471
rect 1887 467 1888 471
rect 1882 466 1888 467
rect 1482 462 1488 463
rect 4634 459 4640 460
rect 4634 458 4635 459
rect 4549 456 4635 458
rect 4634 455 4635 456
rect 4639 455 4640 459
rect 5542 459 5548 460
rect 4634 454 4640 455
rect 4650 455 4656 456
rect 1914 451 1920 452
rect 1914 447 1915 451
rect 1919 450 1920 451
rect 3634 451 3640 452
rect 1919 448 2001 450
rect 1919 447 1920 448
rect 1914 446 1920 447
rect 2210 447 2216 448
rect 2210 443 2211 447
rect 2215 443 2216 447
rect 2210 442 2216 443
rect 2434 447 2440 448
rect 2434 443 2435 447
rect 2439 443 2440 447
rect 2434 442 2440 443
rect 2658 447 2664 448
rect 2658 443 2659 447
rect 2663 443 2664 447
rect 2658 442 2664 443
rect 2954 447 2960 448
rect 2954 443 2955 447
rect 2959 443 2960 447
rect 2954 442 2960 443
rect 3074 447 3080 448
rect 3074 443 3075 447
rect 3079 443 3080 447
rect 3074 442 3080 443
rect 3274 447 3280 448
rect 3274 443 3275 447
rect 3279 443 3280 447
rect 3274 442 3280 443
rect 3474 447 3480 448
rect 3474 443 3475 447
rect 3479 443 3480 447
rect 3634 447 3635 451
rect 3639 450 3640 451
rect 4650 451 4651 455
rect 4655 451 4656 455
rect 4650 450 4656 451
rect 4850 455 4856 456
rect 4850 451 4851 455
rect 4855 451 4856 455
rect 4850 450 4856 451
rect 5058 455 5064 456
rect 5058 451 5059 455
rect 5063 451 5064 455
rect 5058 450 5064 451
rect 5362 455 5368 456
rect 5362 451 5363 455
rect 5367 451 5368 455
rect 5542 455 5543 459
rect 5547 455 5548 459
rect 5542 454 5548 455
rect 5362 450 5368 451
rect 3639 448 3657 450
rect 3639 447 3640 448
rect 3634 446 3640 447
rect 3474 442 3480 443
rect 250 435 256 436
rect 250 431 251 435
rect 255 434 256 435
rect 906 435 912 436
rect 255 432 502 434
rect 255 431 256 432
rect 250 430 256 431
rect 226 427 232 428
rect 226 423 227 427
rect 231 426 232 427
rect 279 427 285 428
rect 279 426 280 427
rect 231 424 280 426
rect 231 423 232 424
rect 226 422 232 423
rect 279 423 280 424
rect 284 423 285 427
rect 500 426 502 432
rect 906 431 907 435
rect 911 434 912 435
rect 911 432 1494 434
rect 911 431 912 432
rect 906 430 912 431
rect 607 427 613 428
rect 607 426 608 427
rect 500 424 608 426
rect 279 422 285 423
rect 607 423 608 424
rect 612 423 613 427
rect 607 422 613 423
rect 934 427 941 428
rect 934 423 935 427
rect 940 423 941 427
rect 934 422 941 423
rect 1263 427 1269 428
rect 1263 423 1264 427
rect 1268 426 1269 427
rect 1482 427 1488 428
rect 1482 426 1483 427
rect 1268 424 1483 426
rect 1268 423 1269 424
rect 1263 422 1269 423
rect 1482 423 1483 424
rect 1487 423 1488 427
rect 1492 426 1494 432
rect 1599 427 1605 428
rect 1599 426 1600 427
rect 1492 424 1600 426
rect 1482 422 1488 423
rect 1599 423 1600 424
rect 1604 423 1605 427
rect 1599 422 1605 423
rect 1911 427 1920 428
rect 1911 423 1912 427
rect 1919 423 1920 427
rect 1911 422 1920 423
rect 110 420 116 421
rect 1934 420 1940 421
rect 110 416 111 420
rect 115 416 116 420
rect 110 415 116 416
rect 154 419 160 420
rect 154 415 155 419
rect 159 415 160 419
rect 154 414 160 415
rect 482 419 488 420
rect 482 415 483 419
rect 487 415 488 419
rect 482 414 488 415
rect 810 419 816 420
rect 810 415 811 419
rect 815 415 816 419
rect 810 414 816 415
rect 1138 419 1144 420
rect 1138 415 1139 419
rect 1143 415 1144 419
rect 1138 414 1144 415
rect 1474 419 1480 420
rect 1474 415 1475 419
rect 1479 415 1480 419
rect 1474 414 1480 415
rect 1786 419 1792 420
rect 1786 415 1787 419
rect 1791 415 1792 419
rect 1934 416 1935 420
rect 1939 416 1940 420
rect 1934 415 1940 416
rect 3202 415 3208 416
rect 1786 414 1792 415
rect 3202 411 3203 415
rect 3207 414 3208 415
rect 4575 415 4581 416
rect 3207 412 3621 414
rect 3207 411 3208 412
rect 3202 410 3208 411
rect 3619 410 3621 412
rect 4575 411 4576 415
rect 4580 414 4581 415
rect 4650 415 4656 416
rect 4650 414 4651 415
rect 4580 412 4651 414
rect 4580 411 4581 412
rect 4575 410 4581 411
rect 4650 411 4651 412
rect 4655 411 4656 415
rect 4650 410 4656 411
rect 4767 415 4773 416
rect 4767 411 4768 415
rect 4772 414 4773 415
rect 4850 415 4856 416
rect 4850 414 4851 415
rect 4772 412 4851 414
rect 4772 411 4773 412
rect 4767 410 4773 411
rect 4850 411 4851 412
rect 4855 411 4856 415
rect 4850 410 4856 411
rect 4967 415 4973 416
rect 4967 411 4968 415
rect 4972 414 4973 415
rect 5058 415 5064 416
rect 5058 414 5059 415
rect 4972 412 5059 414
rect 4972 411 4973 412
rect 4967 410 4973 411
rect 5058 411 5059 412
rect 5063 411 5064 415
rect 5058 410 5064 411
rect 5118 415 5124 416
rect 5118 411 5119 415
rect 5123 414 5124 415
rect 5175 415 5181 416
rect 5175 414 5176 415
rect 5123 412 5176 414
rect 5123 411 5124 412
rect 5118 410 5124 411
rect 5175 411 5176 412
rect 5180 411 5181 415
rect 5175 410 5181 411
rect 5391 415 5400 416
rect 5391 411 5392 415
rect 5399 411 5400 415
rect 5391 410 5400 411
rect 5594 415 5600 416
rect 5594 411 5595 415
rect 5599 414 5600 415
rect 5607 415 5613 416
rect 5607 414 5608 415
rect 5599 412 5608 414
rect 5599 411 5600 412
rect 5594 410 5600 411
rect 5607 411 5608 412
rect 5612 411 5613 415
rect 5607 410 5613 411
rect 3619 408 3758 410
rect 3838 408 3844 409
rect 5662 408 5668 409
rect 2119 407 2125 408
rect 182 404 188 405
rect 110 403 116 404
rect 110 399 111 403
rect 115 399 116 403
rect 182 400 183 404
rect 187 400 188 404
rect 182 399 188 400
rect 510 404 516 405
rect 510 400 511 404
rect 515 400 516 404
rect 510 399 516 400
rect 838 404 844 405
rect 838 400 839 404
rect 843 400 844 404
rect 838 399 844 400
rect 1166 404 1172 405
rect 1166 400 1167 404
rect 1171 400 1172 404
rect 1166 399 1172 400
rect 1502 404 1508 405
rect 1502 400 1503 404
rect 1507 400 1508 404
rect 1502 399 1508 400
rect 1814 404 1820 405
rect 1814 400 1815 404
rect 1819 400 1820 404
rect 1814 399 1820 400
rect 1934 403 1940 404
rect 1934 399 1935 403
rect 1939 399 1940 403
rect 2119 403 2120 407
rect 2124 406 2125 407
rect 2210 407 2216 408
rect 2210 406 2211 407
rect 2124 404 2211 406
rect 2124 403 2125 404
rect 2119 402 2125 403
rect 2210 403 2211 404
rect 2215 403 2216 407
rect 2210 402 2216 403
rect 2327 407 2333 408
rect 2327 403 2328 407
rect 2332 406 2333 407
rect 2434 407 2440 408
rect 2434 406 2435 407
rect 2332 404 2435 406
rect 2332 403 2333 404
rect 2327 402 2333 403
rect 2434 403 2435 404
rect 2439 403 2440 407
rect 2434 402 2440 403
rect 2551 407 2557 408
rect 2551 403 2552 407
rect 2556 406 2557 407
rect 2658 407 2664 408
rect 2658 406 2659 407
rect 2556 404 2659 406
rect 2556 403 2557 404
rect 2551 402 2557 403
rect 2658 403 2659 404
rect 2663 403 2664 407
rect 2658 402 2664 403
rect 2686 407 2692 408
rect 2686 403 2687 407
rect 2691 406 2692 407
rect 2775 407 2781 408
rect 2775 406 2776 407
rect 2691 404 2776 406
rect 2691 403 2692 404
rect 2686 402 2692 403
rect 2775 403 2776 404
rect 2780 403 2781 407
rect 2775 402 2781 403
rect 2983 407 2989 408
rect 2983 403 2984 407
rect 2988 406 2989 407
rect 3074 407 3080 408
rect 3074 406 3075 407
rect 2988 404 3075 406
rect 2988 403 2989 404
rect 2983 402 2989 403
rect 3074 403 3075 404
rect 3079 403 3080 407
rect 3074 402 3080 403
rect 3191 407 3197 408
rect 3191 403 3192 407
rect 3196 406 3197 407
rect 3274 407 3280 408
rect 3274 406 3275 407
rect 3196 404 3275 406
rect 3196 403 3197 404
rect 3191 402 3197 403
rect 3274 403 3275 404
rect 3279 403 3280 407
rect 3274 402 3280 403
rect 3391 407 3397 408
rect 3391 403 3392 407
rect 3396 406 3397 407
rect 3474 407 3480 408
rect 3474 406 3475 407
rect 3396 404 3475 406
rect 3396 403 3397 404
rect 3391 402 3397 403
rect 3474 403 3475 404
rect 3479 403 3480 407
rect 3474 402 3480 403
rect 3591 407 3597 408
rect 3591 403 3592 407
rect 3596 406 3597 407
rect 3756 406 3758 408
rect 3775 407 3781 408
rect 3775 406 3776 407
rect 3596 404 3638 406
rect 3756 404 3776 406
rect 3596 403 3597 404
rect 3591 402 3597 403
rect 3634 403 3640 404
rect 110 398 116 399
rect 1934 398 1940 399
rect 1974 400 1980 401
rect 1974 396 1975 400
rect 1979 396 1980 400
rect 1974 395 1980 396
rect 1994 399 2000 400
rect 1994 395 1995 399
rect 1999 395 2000 399
rect 1994 394 2000 395
rect 2202 399 2208 400
rect 2202 395 2203 399
rect 2207 395 2208 399
rect 2202 394 2208 395
rect 2426 399 2432 400
rect 2426 395 2427 399
rect 2431 395 2432 399
rect 2426 394 2432 395
rect 2650 399 2656 400
rect 2650 395 2651 399
rect 2655 395 2656 399
rect 2650 394 2656 395
rect 2858 399 2864 400
rect 2858 395 2859 399
rect 2863 395 2864 399
rect 2858 394 2864 395
rect 3066 399 3072 400
rect 3066 395 3067 399
rect 3071 395 3072 399
rect 3066 394 3072 395
rect 3266 399 3272 400
rect 3266 395 3267 399
rect 3271 395 3272 399
rect 3266 394 3272 395
rect 3466 399 3472 400
rect 3466 395 3467 399
rect 3471 395 3472 399
rect 3634 399 3635 403
rect 3639 399 3640 403
rect 3775 403 3776 404
rect 3780 403 3781 407
rect 3838 404 3839 408
rect 3843 404 3844 408
rect 3838 403 3844 404
rect 4450 407 4456 408
rect 4450 403 4451 407
rect 4455 403 4456 407
rect 3775 402 3781 403
rect 4450 402 4456 403
rect 4642 407 4648 408
rect 4642 403 4643 407
rect 4647 403 4648 407
rect 4642 402 4648 403
rect 4842 407 4848 408
rect 4842 403 4843 407
rect 4847 403 4848 407
rect 4842 402 4848 403
rect 5050 407 5056 408
rect 5050 403 5051 407
rect 5055 403 5056 407
rect 5050 402 5056 403
rect 5266 407 5272 408
rect 5266 403 5267 407
rect 5271 403 5272 407
rect 5266 402 5272 403
rect 5482 407 5488 408
rect 5482 403 5483 407
rect 5487 403 5488 407
rect 5662 404 5663 408
rect 5667 404 5668 408
rect 5662 403 5668 404
rect 5482 402 5488 403
rect 3798 400 3804 401
rect 3634 398 3640 399
rect 3650 399 3656 400
rect 3466 394 3472 395
rect 3650 395 3651 399
rect 3655 395 3656 399
rect 3798 396 3799 400
rect 3803 396 3804 400
rect 3798 395 3804 396
rect 3650 394 3656 395
rect 4478 392 4484 393
rect 3838 391 3844 392
rect 3838 387 3839 391
rect 3843 387 3844 391
rect 4478 388 4479 392
rect 4483 388 4484 392
rect 4478 387 4484 388
rect 4670 392 4676 393
rect 4670 388 4671 392
rect 4675 388 4676 392
rect 4670 387 4676 388
rect 4870 392 4876 393
rect 4870 388 4871 392
rect 4875 388 4876 392
rect 4870 387 4876 388
rect 5078 392 5084 393
rect 5078 388 5079 392
rect 5083 388 5084 392
rect 5078 387 5084 388
rect 5294 392 5300 393
rect 5294 388 5295 392
rect 5299 388 5300 392
rect 5294 387 5300 388
rect 5510 392 5516 393
rect 5510 388 5511 392
rect 5515 388 5516 392
rect 5510 387 5516 388
rect 5662 391 5668 392
rect 5662 387 5663 391
rect 5667 387 5668 391
rect 3838 386 3844 387
rect 5662 386 5668 387
rect 2022 384 2028 385
rect 1974 383 1980 384
rect 1974 379 1975 383
rect 1979 379 1980 383
rect 2022 380 2023 384
rect 2027 380 2028 384
rect 2022 379 2028 380
rect 2230 384 2236 385
rect 2230 380 2231 384
rect 2235 380 2236 384
rect 2230 379 2236 380
rect 2454 384 2460 385
rect 2454 380 2455 384
rect 2459 380 2460 384
rect 2454 379 2460 380
rect 2678 384 2684 385
rect 2678 380 2679 384
rect 2683 380 2684 384
rect 2678 379 2684 380
rect 2886 384 2892 385
rect 2886 380 2887 384
rect 2891 380 2892 384
rect 2886 379 2892 380
rect 3094 384 3100 385
rect 3094 380 3095 384
rect 3099 380 3100 384
rect 3094 379 3100 380
rect 3294 384 3300 385
rect 3294 380 3295 384
rect 3299 380 3300 384
rect 3294 379 3300 380
rect 3494 384 3500 385
rect 3494 380 3495 384
rect 3499 380 3500 384
rect 3494 379 3500 380
rect 3678 384 3684 385
rect 3678 380 3679 384
rect 3683 380 3684 384
rect 3678 379 3684 380
rect 3798 383 3804 384
rect 3798 379 3799 383
rect 3803 379 3804 383
rect 1974 378 1980 379
rect 3798 378 3804 379
rect 110 333 116 334
rect 1934 333 1940 334
rect 110 329 111 333
rect 115 329 116 333
rect 110 328 116 329
rect 278 332 284 333
rect 278 328 279 332
rect 283 328 284 332
rect 278 327 284 328
rect 486 332 492 333
rect 486 328 487 332
rect 491 328 492 332
rect 486 327 492 328
rect 702 332 708 333
rect 702 328 703 332
rect 707 328 708 332
rect 702 327 708 328
rect 918 332 924 333
rect 918 328 919 332
rect 923 328 924 332
rect 918 327 924 328
rect 1134 332 1140 333
rect 1134 328 1135 332
rect 1139 328 1140 332
rect 1934 329 1935 333
rect 1939 329 1940 333
rect 1934 328 1940 329
rect 3838 329 3844 330
rect 5662 329 5668 330
rect 1134 327 1140 328
rect 3838 325 3839 329
rect 3843 325 3844 329
rect 3838 324 3844 325
rect 4614 328 4620 329
rect 4614 324 4615 328
rect 4619 324 4620 328
rect 4614 323 4620 324
rect 4774 328 4780 329
rect 4774 324 4775 328
rect 4779 324 4780 328
rect 4774 323 4780 324
rect 4950 328 4956 329
rect 4950 324 4951 328
rect 4955 324 4956 328
rect 4950 323 4956 324
rect 5134 328 5140 329
rect 5134 324 5135 328
rect 5139 324 5140 328
rect 5134 323 5140 324
rect 5326 328 5332 329
rect 5326 324 5327 328
rect 5331 324 5332 328
rect 5326 323 5332 324
rect 5526 328 5532 329
rect 5526 324 5527 328
rect 5531 324 5532 328
rect 5662 325 5663 329
rect 5667 325 5668 329
rect 5662 324 5668 325
rect 5526 323 5532 324
rect 250 317 256 318
rect 110 316 116 317
rect 110 312 111 316
rect 115 312 116 316
rect 250 313 251 317
rect 255 313 256 317
rect 250 312 256 313
rect 458 317 464 318
rect 458 313 459 317
rect 463 313 464 317
rect 458 312 464 313
rect 674 317 680 318
rect 674 313 675 317
rect 679 313 680 317
rect 674 312 680 313
rect 890 317 896 318
rect 890 313 891 317
rect 895 313 896 317
rect 890 312 896 313
rect 1106 317 1112 318
rect 1106 313 1107 317
rect 1111 313 1112 317
rect 1106 312 1112 313
rect 1934 316 1940 317
rect 1934 312 1935 316
rect 1939 312 1940 316
rect 4586 313 4592 314
rect 110 311 116 312
rect 1934 311 1940 312
rect 3838 312 3844 313
rect 1974 309 1980 310
rect 3798 309 3804 310
rect 375 307 381 308
rect 375 303 376 307
rect 380 306 381 307
rect 407 307 413 308
rect 407 306 408 307
rect 380 304 408 306
rect 380 303 381 304
rect 375 302 381 303
rect 407 303 408 304
rect 412 303 413 307
rect 407 302 413 303
rect 578 307 589 308
rect 578 303 579 307
rect 583 303 584 307
rect 588 303 589 307
rect 578 302 589 303
rect 799 307 805 308
rect 799 303 800 307
rect 804 306 805 307
rect 807 307 813 308
rect 807 306 808 307
rect 804 304 808 306
rect 804 303 805 304
rect 799 302 805 303
rect 807 303 808 304
rect 812 303 813 307
rect 807 302 813 303
rect 1015 307 1021 308
rect 1015 303 1016 307
rect 1020 306 1021 307
rect 1062 307 1068 308
rect 1062 306 1063 307
rect 1020 304 1063 306
rect 1020 303 1021 304
rect 1015 302 1021 303
rect 1062 303 1063 304
rect 1067 303 1068 307
rect 1231 307 1237 308
rect 1231 306 1232 307
rect 1062 302 1068 303
rect 1099 304 1232 306
rect 770 299 776 300
rect 770 295 771 299
rect 775 298 776 299
rect 1099 298 1101 304
rect 1231 303 1232 304
rect 1236 303 1237 307
rect 1974 305 1975 309
rect 1979 305 1980 309
rect 1974 304 1980 305
rect 2022 308 2028 309
rect 2022 304 2023 308
rect 2027 304 2028 308
rect 2022 303 2028 304
rect 2158 308 2164 309
rect 2158 304 2159 308
rect 2163 304 2164 308
rect 2158 303 2164 304
rect 2294 308 2300 309
rect 2294 304 2295 308
rect 2299 304 2300 308
rect 2294 303 2300 304
rect 2430 308 2436 309
rect 2430 304 2431 308
rect 2435 304 2436 308
rect 2430 303 2436 304
rect 2566 308 2572 309
rect 2566 304 2567 308
rect 2571 304 2572 308
rect 2566 303 2572 304
rect 2702 308 2708 309
rect 2702 304 2703 308
rect 2707 304 2708 308
rect 2702 303 2708 304
rect 2838 308 2844 309
rect 2838 304 2839 308
rect 2843 304 2844 308
rect 2838 303 2844 304
rect 2974 308 2980 309
rect 2974 304 2975 308
rect 2979 304 2980 308
rect 2974 303 2980 304
rect 3110 308 3116 309
rect 3110 304 3111 308
rect 3115 304 3116 308
rect 3110 303 3116 304
rect 3246 308 3252 309
rect 3246 304 3247 308
rect 3251 304 3252 308
rect 3246 303 3252 304
rect 3382 308 3388 309
rect 3382 304 3383 308
rect 3387 304 3388 308
rect 3382 303 3388 304
rect 3518 308 3524 309
rect 3518 304 3519 308
rect 3523 304 3524 308
rect 3518 303 3524 304
rect 3654 308 3660 309
rect 3654 304 3655 308
rect 3659 304 3660 308
rect 3798 305 3799 309
rect 3803 305 3804 309
rect 3838 308 3839 312
rect 3843 308 3844 312
rect 4586 309 4587 313
rect 4591 309 4592 313
rect 4586 308 4592 309
rect 4746 313 4752 314
rect 4746 309 4747 313
rect 4751 309 4752 313
rect 4746 308 4752 309
rect 4922 313 4928 314
rect 4922 309 4923 313
rect 4927 309 4928 313
rect 4922 308 4928 309
rect 5106 313 5112 314
rect 5106 309 5107 313
rect 5111 309 5112 313
rect 5106 308 5112 309
rect 5298 313 5304 314
rect 5298 309 5299 313
rect 5303 309 5304 313
rect 5298 308 5304 309
rect 5498 313 5504 314
rect 5498 309 5499 313
rect 5503 309 5504 313
rect 5498 308 5504 309
rect 5662 312 5668 313
rect 5662 308 5663 312
rect 5667 308 5668 312
rect 3838 307 3844 308
rect 5662 307 5668 308
rect 3798 304 3804 305
rect 3654 303 3660 304
rect 4711 303 4717 304
rect 1231 302 1237 303
rect 4711 299 4712 303
rect 4716 302 4717 303
rect 4734 303 4740 304
rect 4734 302 4735 303
rect 4716 300 4735 302
rect 4716 299 4717 300
rect 4711 298 4717 299
rect 4734 299 4735 300
rect 4739 299 4740 303
rect 4734 298 4740 299
rect 4871 303 4880 304
rect 4871 299 4872 303
rect 4879 299 4880 303
rect 4871 298 4880 299
rect 5047 303 5056 304
rect 5047 299 5048 303
rect 5055 299 5056 303
rect 5047 298 5056 299
rect 5231 303 5237 304
rect 5231 299 5232 303
rect 5236 302 5237 303
rect 5263 303 5269 304
rect 5263 302 5264 303
rect 5236 300 5264 302
rect 5236 299 5237 300
rect 5231 298 5237 299
rect 5263 299 5264 300
rect 5268 299 5269 303
rect 5423 303 5429 304
rect 5423 302 5424 303
rect 5263 298 5269 299
rect 5299 300 5424 302
rect 775 296 1101 298
rect 775 295 776 296
rect 770 294 776 295
rect 4674 295 4680 296
rect 1994 293 2000 294
rect 1974 292 1980 293
rect 1974 288 1975 292
rect 1979 288 1980 292
rect 1994 289 1995 293
rect 1999 289 2000 293
rect 1994 288 2000 289
rect 2130 293 2136 294
rect 2130 289 2131 293
rect 2135 289 2136 293
rect 2130 288 2136 289
rect 2266 293 2272 294
rect 2266 289 2267 293
rect 2271 289 2272 293
rect 2266 288 2272 289
rect 2402 293 2408 294
rect 2402 289 2403 293
rect 2407 289 2408 293
rect 2402 288 2408 289
rect 2538 293 2544 294
rect 2538 289 2539 293
rect 2543 289 2544 293
rect 2538 288 2544 289
rect 2674 293 2680 294
rect 2674 289 2675 293
rect 2679 289 2680 293
rect 2674 288 2680 289
rect 2810 293 2816 294
rect 2810 289 2811 293
rect 2815 289 2816 293
rect 2810 288 2816 289
rect 2946 293 2952 294
rect 2946 289 2947 293
rect 2951 289 2952 293
rect 2946 288 2952 289
rect 3082 293 3088 294
rect 3082 289 3083 293
rect 3087 289 3088 293
rect 3082 288 3088 289
rect 3218 293 3224 294
rect 3218 289 3219 293
rect 3223 289 3224 293
rect 3218 288 3224 289
rect 3354 293 3360 294
rect 3354 289 3355 293
rect 3359 289 3360 293
rect 3354 288 3360 289
rect 3490 293 3496 294
rect 3490 289 3491 293
rect 3495 289 3496 293
rect 3490 288 3496 289
rect 3626 293 3632 294
rect 3626 289 3627 293
rect 3631 289 3632 293
rect 3626 288 3632 289
rect 3798 292 3804 293
rect 3798 288 3799 292
rect 3803 288 3804 292
rect 4674 291 4675 295
rect 4679 294 4680 295
rect 5299 294 5301 300
rect 5423 299 5424 300
rect 5428 299 5429 303
rect 5423 298 5429 299
rect 5610 303 5616 304
rect 5610 299 5611 303
rect 5615 302 5616 303
rect 5623 303 5629 304
rect 5623 302 5624 303
rect 5615 300 5624 302
rect 5615 299 5616 300
rect 5610 298 5616 299
rect 5623 299 5624 300
rect 5628 299 5629 303
rect 5623 298 5629 299
rect 4679 292 5301 294
rect 4679 291 4680 292
rect 4674 290 4680 291
rect 1974 287 1980 288
rect 3798 287 3804 288
rect 2119 283 2128 284
rect 2119 279 2120 283
rect 2127 279 2128 283
rect 2119 278 2128 279
rect 2255 283 2264 284
rect 2255 279 2256 283
rect 2263 279 2264 283
rect 2255 278 2264 279
rect 2391 283 2400 284
rect 2391 279 2392 283
rect 2399 279 2400 283
rect 2391 278 2400 279
rect 2527 283 2536 284
rect 2527 279 2528 283
rect 2535 279 2536 283
rect 2527 278 2536 279
rect 2663 283 2672 284
rect 2663 279 2664 283
rect 2671 279 2672 283
rect 2663 278 2672 279
rect 2799 283 2808 284
rect 2799 279 2800 283
rect 2807 279 2808 283
rect 2799 278 2808 279
rect 2854 283 2860 284
rect 2854 279 2855 283
rect 2859 282 2860 283
rect 2935 283 2941 284
rect 2935 282 2936 283
rect 2859 280 2936 282
rect 2859 279 2860 280
rect 2854 278 2860 279
rect 2935 279 2936 280
rect 2940 279 2941 283
rect 2935 278 2941 279
rect 3071 283 3080 284
rect 3071 279 3072 283
rect 3079 279 3080 283
rect 3071 278 3080 279
rect 3207 283 3216 284
rect 3207 279 3208 283
rect 3215 279 3216 283
rect 3207 278 3216 279
rect 3343 283 3352 284
rect 3343 279 3344 283
rect 3351 279 3352 283
rect 3343 278 3352 279
rect 3479 283 3488 284
rect 3479 279 3480 283
rect 3487 279 3488 283
rect 3479 278 3488 279
rect 3615 283 3621 284
rect 3615 279 3616 283
rect 3620 282 3621 283
rect 3623 283 3629 284
rect 3623 282 3624 283
rect 3620 280 3624 282
rect 3620 279 3621 280
rect 3615 278 3621 279
rect 3623 279 3624 280
rect 3628 279 3629 283
rect 3751 283 3757 284
rect 3751 282 3752 283
rect 3623 278 3629 279
rect 3684 280 3752 282
rect 2090 275 2096 276
rect 2090 271 2091 275
rect 2095 274 2096 275
rect 2686 275 2692 276
rect 2686 274 2687 275
rect 2095 272 2687 274
rect 2095 271 2096 272
rect 2090 270 2096 271
rect 2686 271 2687 272
rect 2691 271 2692 275
rect 2686 270 2692 271
rect 346 267 352 268
rect 346 263 347 267
rect 351 263 352 267
rect 346 262 352 263
rect 407 267 413 268
rect 407 263 408 267
rect 412 266 413 267
rect 770 267 776 268
rect 412 264 465 266
rect 412 263 413 264
rect 407 262 413 263
rect 770 263 771 267
rect 775 263 776 267
rect 770 262 776 263
rect 934 267 940 268
rect 934 263 935 267
rect 939 263 940 267
rect 934 262 940 263
rect 1062 267 1068 268
rect 1062 263 1063 267
rect 1067 266 1068 267
rect 2954 267 2960 268
rect 1067 264 1113 266
rect 1067 263 1068 264
rect 1062 262 1068 263
rect 2954 263 2955 267
rect 2959 266 2960 267
rect 3684 266 3686 280
rect 3751 279 3752 280
rect 3756 279 3757 283
rect 3751 278 3757 279
rect 2959 264 3686 266
rect 2959 263 2960 264
rect 2954 262 2960 263
rect 4734 263 4740 264
rect 4386 255 4392 256
rect 4386 251 4387 255
rect 4391 254 4392 255
rect 4674 255 4680 256
rect 4674 254 4675 255
rect 4391 252 4675 254
rect 4391 251 4392 252
rect 4386 250 4392 251
rect 4674 251 4675 252
rect 4679 251 4680 255
rect 4684 254 4686 261
rect 4734 259 4735 263
rect 4739 262 4740 263
rect 4874 263 4880 264
rect 4739 260 4753 262
rect 4739 259 4740 260
rect 4734 258 4740 259
rect 4874 259 4875 263
rect 4879 262 4880 263
rect 5050 263 5056 264
rect 4879 260 4929 262
rect 4879 259 4880 260
rect 4874 258 4880 259
rect 5050 259 5051 263
rect 5055 262 5056 263
rect 5263 263 5269 264
rect 5055 260 5113 262
rect 5055 259 5056 260
rect 5050 258 5056 259
rect 5263 259 5264 263
rect 5268 262 5269 263
rect 5594 263 5600 264
rect 5268 260 5305 262
rect 5268 259 5269 260
rect 5263 258 5269 259
rect 5594 259 5595 263
rect 5599 259 5600 263
rect 5594 258 5600 259
rect 5118 255 5124 256
rect 5118 254 5119 255
rect 4684 252 5119 254
rect 4674 250 4680 251
rect 5118 251 5119 252
rect 5123 251 5124 255
rect 5118 250 5124 251
rect 2090 243 2096 244
rect 2090 239 2091 243
rect 2095 239 2096 243
rect 2090 238 2096 239
rect 2122 243 2128 244
rect 2122 239 2123 243
rect 2127 242 2128 243
rect 2258 243 2264 244
rect 2127 240 2137 242
rect 2127 239 2128 240
rect 2122 238 2128 239
rect 2258 239 2259 243
rect 2263 242 2264 243
rect 2394 243 2400 244
rect 2263 240 2273 242
rect 2263 239 2264 240
rect 2258 238 2264 239
rect 2394 239 2395 243
rect 2399 242 2400 243
rect 2530 243 2536 244
rect 2399 240 2409 242
rect 2399 239 2400 240
rect 2394 238 2400 239
rect 2530 239 2531 243
rect 2535 242 2536 243
rect 2666 243 2672 244
rect 2535 240 2545 242
rect 2535 239 2536 240
rect 2530 238 2536 239
rect 2666 239 2667 243
rect 2671 242 2672 243
rect 2802 243 2808 244
rect 2671 240 2681 242
rect 2671 239 2672 240
rect 2666 238 2672 239
rect 2802 239 2803 243
rect 2807 242 2808 243
rect 3042 243 3048 244
rect 2807 240 2817 242
rect 2807 239 2808 240
rect 2802 238 2808 239
rect 3042 239 3043 243
rect 3047 239 3048 243
rect 3042 238 3048 239
rect 3074 243 3080 244
rect 3074 239 3075 243
rect 3079 242 3080 243
rect 3210 243 3216 244
rect 3079 240 3089 242
rect 3079 239 3080 240
rect 3074 238 3080 239
rect 3210 239 3211 243
rect 3215 242 3216 243
rect 3346 243 3352 244
rect 3215 240 3225 242
rect 3215 239 3216 240
rect 3210 238 3216 239
rect 3346 239 3347 243
rect 3351 242 3352 243
rect 3482 243 3488 244
rect 3351 240 3361 242
rect 3351 239 3352 240
rect 3346 238 3352 239
rect 3482 239 3483 243
rect 3487 242 3488 243
rect 3623 243 3629 244
rect 3487 240 3497 242
rect 3487 239 3488 240
rect 3482 238 3488 239
rect 3623 239 3624 243
rect 3628 242 3629 243
rect 3628 240 3633 242
rect 3628 239 3629 240
rect 3623 238 3629 239
rect 2090 235 2096 236
rect 2090 231 2091 235
rect 2095 234 2096 235
rect 2854 235 2860 236
rect 2854 234 2855 235
rect 2095 232 2855 234
rect 2095 231 2096 232
rect 2090 230 2096 231
rect 2854 231 2855 232
rect 2859 231 2860 235
rect 2854 230 2860 231
rect 1206 203 1212 204
rect 1206 202 1207 203
rect 800 200 1207 202
rect 535 195 541 196
rect 535 194 536 195
rect 501 192 536 194
rect 226 191 232 192
rect 226 187 227 191
rect 231 187 232 191
rect 226 186 232 187
rect 274 191 280 192
rect 274 187 275 191
rect 279 187 280 191
rect 535 191 536 192
rect 540 191 541 195
rect 800 194 802 200
rect 1206 199 1207 200
rect 1211 199 1212 203
rect 1206 198 1212 199
rect 773 192 802 194
rect 807 195 813 196
rect 535 190 541 191
rect 634 191 640 192
rect 274 186 280 187
rect 634 187 635 191
rect 639 187 640 191
rect 807 191 808 195
rect 812 194 813 195
rect 812 192 817 194
rect 812 191 813 192
rect 807 190 813 191
rect 954 191 960 192
rect 634 186 640 187
rect 954 187 955 191
rect 959 187 960 191
rect 954 186 960 187
rect 1090 191 1096 192
rect 1090 187 1091 191
rect 1095 187 1096 191
rect 1090 186 1096 187
rect 4386 191 4392 192
rect 4386 187 4387 191
rect 4391 187 4392 191
rect 5610 191 5616 192
rect 4386 186 4392 187
rect 4434 187 4440 188
rect 4434 183 4435 187
rect 4439 183 4440 187
rect 4434 182 4440 183
rect 4570 187 4576 188
rect 4570 183 4571 187
rect 4575 183 4576 187
rect 4570 182 4576 183
rect 4706 187 4712 188
rect 4706 183 4707 187
rect 4711 183 4712 187
rect 4706 182 4712 183
rect 4842 187 4848 188
rect 4842 183 4843 187
rect 4847 183 4848 187
rect 4842 182 4848 183
rect 4978 187 4984 188
rect 4978 183 4979 187
rect 4983 183 4984 187
rect 4978 182 4984 183
rect 5114 187 5120 188
rect 5114 183 5115 187
rect 5119 183 5120 187
rect 5114 182 5120 183
rect 5250 187 5256 188
rect 5250 183 5251 187
rect 5255 183 5256 187
rect 5250 182 5256 183
rect 5474 187 5480 188
rect 5474 183 5475 187
rect 5479 183 5480 187
rect 5610 187 5611 191
rect 5615 187 5616 191
rect 5610 186 5616 187
rect 5474 182 5480 183
rect 2090 175 2096 176
rect 2090 171 2091 175
rect 2095 171 2096 175
rect 2090 170 2096 171
rect 2138 171 2144 172
rect 2138 167 2139 171
rect 2143 167 2144 171
rect 2138 166 2144 167
rect 2274 171 2280 172
rect 2274 167 2275 171
rect 2279 167 2280 171
rect 2274 166 2280 167
rect 2410 171 2416 172
rect 2410 167 2411 171
rect 2415 167 2416 171
rect 2410 166 2416 167
rect 2546 171 2552 172
rect 2546 167 2547 171
rect 2551 167 2552 171
rect 2546 166 2552 167
rect 2682 171 2688 172
rect 2682 167 2683 171
rect 2687 167 2688 171
rect 2682 166 2688 167
rect 2818 171 2824 172
rect 2818 167 2819 171
rect 2823 167 2824 171
rect 2818 166 2824 167
rect 2954 171 2960 172
rect 2954 167 2955 171
rect 2959 167 2960 171
rect 2954 166 2960 167
rect 3090 171 3096 172
rect 3090 167 3091 171
rect 3095 167 3096 171
rect 3090 166 3096 167
rect 3226 171 3232 172
rect 3226 167 3227 171
rect 3231 167 3232 171
rect 3226 166 3232 167
rect 3362 171 3368 172
rect 3362 167 3363 171
rect 3367 167 3368 171
rect 3362 166 3368 167
rect 3498 171 3504 172
rect 3498 167 3499 171
rect 3503 167 3504 171
rect 3498 166 3504 167
rect 3634 171 3640 172
rect 3634 167 3635 171
rect 3639 167 3640 171
rect 3634 166 3640 167
rect 226 159 232 160
rect 226 155 227 159
rect 231 158 232 159
rect 634 159 640 160
rect 231 156 402 158
rect 231 155 232 156
rect 226 154 232 155
rect 255 151 261 152
rect 255 147 256 151
rect 260 150 261 151
rect 274 151 280 152
rect 274 150 275 151
rect 260 148 275 150
rect 260 147 261 148
rect 255 146 261 147
rect 274 147 275 148
rect 279 147 280 151
rect 274 146 280 147
rect 346 151 352 152
rect 346 147 347 151
rect 351 150 352 151
rect 391 151 397 152
rect 391 150 392 151
rect 351 148 392 150
rect 351 147 352 148
rect 346 146 352 147
rect 391 147 392 148
rect 396 147 397 151
rect 400 150 402 156
rect 634 155 635 159
rect 639 158 640 159
rect 639 156 674 158
rect 639 155 640 156
rect 634 154 640 155
rect 527 151 533 152
rect 527 150 528 151
rect 400 148 528 150
rect 391 146 397 147
rect 527 147 528 148
rect 532 147 533 151
rect 527 146 533 147
rect 535 151 541 152
rect 535 147 536 151
rect 540 150 541 151
rect 663 151 669 152
rect 663 150 664 151
rect 540 148 664 150
rect 540 147 541 148
rect 535 146 541 147
rect 663 147 664 148
rect 668 147 669 151
rect 672 150 674 156
rect 799 151 805 152
rect 799 150 800 151
rect 672 148 800 150
rect 663 146 669 147
rect 799 147 800 148
rect 804 147 805 151
rect 799 146 805 147
rect 935 151 941 152
rect 935 147 936 151
rect 940 150 941 151
rect 954 151 960 152
rect 954 150 955 151
rect 940 148 955 150
rect 940 147 941 148
rect 935 146 941 147
rect 954 147 955 148
rect 959 147 960 151
rect 954 146 960 147
rect 1071 151 1077 152
rect 1071 147 1072 151
rect 1076 150 1077 151
rect 1090 151 1096 152
rect 1090 150 1091 151
rect 1076 148 1091 150
rect 1076 147 1077 148
rect 1071 146 1077 147
rect 1090 147 1091 148
rect 1095 147 1096 151
rect 1090 146 1096 147
rect 1206 151 1213 152
rect 1206 147 1207 151
rect 1212 147 1213 151
rect 1206 146 1213 147
rect 4415 147 4421 148
rect 110 144 116 145
rect 1934 144 1940 145
rect 110 140 111 144
rect 115 140 116 144
rect 110 139 116 140
rect 130 143 136 144
rect 130 139 131 143
rect 135 139 136 143
rect 130 138 136 139
rect 266 143 272 144
rect 266 139 267 143
rect 271 139 272 143
rect 266 138 272 139
rect 402 143 408 144
rect 402 139 403 143
rect 407 139 408 143
rect 402 138 408 139
rect 538 143 544 144
rect 538 139 539 143
rect 543 139 544 143
rect 538 138 544 139
rect 674 143 680 144
rect 674 139 675 143
rect 679 139 680 143
rect 674 138 680 139
rect 810 143 816 144
rect 810 139 811 143
rect 815 139 816 143
rect 810 138 816 139
rect 946 143 952 144
rect 946 139 947 143
rect 951 139 952 143
rect 946 138 952 139
rect 1082 143 1088 144
rect 1082 139 1083 143
rect 1087 139 1088 143
rect 1934 140 1935 144
rect 1939 140 1940 144
rect 4415 143 4416 147
rect 4420 146 4421 147
rect 4434 147 4440 148
rect 4434 146 4435 147
rect 4420 144 4435 146
rect 4420 143 4421 144
rect 4415 142 4421 143
rect 4434 143 4435 144
rect 4439 143 4440 147
rect 4434 142 4440 143
rect 4551 147 4557 148
rect 4551 143 4552 147
rect 4556 146 4557 147
rect 4570 147 4576 148
rect 4570 146 4571 147
rect 4556 144 4571 146
rect 4556 143 4557 144
rect 4551 142 4557 143
rect 4570 143 4571 144
rect 4575 143 4576 147
rect 4570 142 4576 143
rect 4687 147 4693 148
rect 4687 143 4688 147
rect 4692 146 4693 147
rect 4706 147 4712 148
rect 4706 146 4707 147
rect 4692 144 4707 146
rect 4692 143 4693 144
rect 4687 142 4693 143
rect 4706 143 4707 144
rect 4711 143 4712 147
rect 4706 142 4712 143
rect 4823 147 4829 148
rect 4823 143 4824 147
rect 4828 146 4829 147
rect 4842 147 4848 148
rect 4842 146 4843 147
rect 4828 144 4843 146
rect 4828 143 4829 144
rect 4823 142 4829 143
rect 4842 143 4843 144
rect 4847 143 4848 147
rect 4842 142 4848 143
rect 4959 147 4965 148
rect 4959 143 4960 147
rect 4964 146 4965 147
rect 4978 147 4984 148
rect 4978 146 4979 147
rect 4964 144 4979 146
rect 4964 143 4965 144
rect 4959 142 4965 143
rect 4978 143 4979 144
rect 4983 143 4984 147
rect 4978 142 4984 143
rect 5095 147 5101 148
rect 5095 143 5096 147
rect 5100 146 5101 147
rect 5114 147 5120 148
rect 5114 146 5115 147
rect 5100 144 5115 146
rect 5100 143 5101 144
rect 5095 142 5101 143
rect 5114 143 5115 144
rect 5119 143 5120 147
rect 5114 142 5120 143
rect 5231 147 5237 148
rect 5231 143 5232 147
rect 5236 146 5237 147
rect 5250 147 5256 148
rect 5250 146 5251 147
rect 5236 144 5251 146
rect 5236 143 5237 144
rect 5231 142 5237 143
rect 5250 143 5251 144
rect 5255 143 5256 147
rect 5250 142 5256 143
rect 5362 147 5373 148
rect 5362 143 5363 147
rect 5367 143 5368 147
rect 5372 143 5373 147
rect 5362 142 5373 143
rect 5474 147 5480 148
rect 5474 143 5475 147
rect 5479 146 5480 147
rect 5639 147 5645 148
rect 5639 146 5640 147
rect 5479 144 5640 146
rect 5479 143 5480 144
rect 5474 142 5480 143
rect 5639 143 5640 144
rect 5644 143 5645 147
rect 5639 142 5645 143
rect 1934 139 1940 140
rect 3838 140 3844 141
rect 5662 140 5668 141
rect 1082 138 1088 139
rect 3838 136 3839 140
rect 3843 136 3844 140
rect 3838 135 3844 136
rect 4290 139 4296 140
rect 4290 135 4291 139
rect 4295 135 4296 139
rect 4290 134 4296 135
rect 4426 139 4432 140
rect 4426 135 4427 139
rect 4431 135 4432 139
rect 4426 134 4432 135
rect 4562 139 4568 140
rect 4562 135 4563 139
rect 4567 135 4568 139
rect 4562 134 4568 135
rect 4698 139 4704 140
rect 4698 135 4699 139
rect 4703 135 4704 139
rect 4698 134 4704 135
rect 4834 139 4840 140
rect 4834 135 4835 139
rect 4839 135 4840 139
rect 4834 134 4840 135
rect 4970 139 4976 140
rect 4970 135 4971 139
rect 4975 135 4976 139
rect 4970 134 4976 135
rect 5106 139 5112 140
rect 5106 135 5107 139
rect 5111 135 5112 139
rect 5106 134 5112 135
rect 5242 139 5248 140
rect 5242 135 5243 139
rect 5247 135 5248 139
rect 5242 134 5248 135
rect 5378 139 5384 140
rect 5378 135 5379 139
rect 5383 135 5384 139
rect 5378 134 5384 135
rect 5514 139 5520 140
rect 5514 135 5515 139
rect 5519 135 5520 139
rect 5662 136 5663 140
rect 5667 136 5668 140
rect 5662 135 5668 136
rect 5514 134 5520 135
rect 2119 131 2125 132
rect 158 128 164 129
rect 110 127 116 128
rect 110 123 111 127
rect 115 123 116 127
rect 158 124 159 128
rect 163 124 164 128
rect 158 123 164 124
rect 294 128 300 129
rect 294 124 295 128
rect 299 124 300 128
rect 294 123 300 124
rect 430 128 436 129
rect 430 124 431 128
rect 435 124 436 128
rect 430 123 436 124
rect 566 128 572 129
rect 566 124 567 128
rect 571 124 572 128
rect 566 123 572 124
rect 702 128 708 129
rect 702 124 703 128
rect 707 124 708 128
rect 702 123 708 124
rect 838 128 844 129
rect 838 124 839 128
rect 843 124 844 128
rect 838 123 844 124
rect 974 128 980 129
rect 974 124 975 128
rect 979 124 980 128
rect 974 123 980 124
rect 1110 128 1116 129
rect 1110 124 1111 128
rect 1115 124 1116 128
rect 1110 123 1116 124
rect 1934 127 1940 128
rect 1934 123 1935 127
rect 1939 123 1940 127
rect 2119 127 2120 131
rect 2124 130 2125 131
rect 2138 131 2144 132
rect 2138 130 2139 131
rect 2124 128 2139 130
rect 2124 127 2125 128
rect 2119 126 2125 127
rect 2138 127 2139 128
rect 2143 127 2144 131
rect 2138 126 2144 127
rect 2255 131 2261 132
rect 2255 127 2256 131
rect 2260 130 2261 131
rect 2274 131 2280 132
rect 2274 130 2275 131
rect 2260 128 2275 130
rect 2260 127 2261 128
rect 2255 126 2261 127
rect 2274 127 2275 128
rect 2279 127 2280 131
rect 2274 126 2280 127
rect 2391 131 2397 132
rect 2391 127 2392 131
rect 2396 130 2397 131
rect 2410 131 2416 132
rect 2410 130 2411 131
rect 2396 128 2411 130
rect 2396 127 2397 128
rect 2391 126 2397 127
rect 2410 127 2411 128
rect 2415 127 2416 131
rect 2410 126 2416 127
rect 2527 131 2533 132
rect 2527 127 2528 131
rect 2532 130 2533 131
rect 2546 131 2552 132
rect 2546 130 2547 131
rect 2532 128 2547 130
rect 2532 127 2533 128
rect 2527 126 2533 127
rect 2546 127 2547 128
rect 2551 127 2552 131
rect 2546 126 2552 127
rect 2663 131 2669 132
rect 2663 127 2664 131
rect 2668 130 2669 131
rect 2682 131 2688 132
rect 2682 130 2683 131
rect 2668 128 2683 130
rect 2668 127 2669 128
rect 2663 126 2669 127
rect 2682 127 2683 128
rect 2687 127 2688 131
rect 2682 126 2688 127
rect 2799 131 2805 132
rect 2799 127 2800 131
rect 2804 130 2805 131
rect 2818 131 2824 132
rect 2818 130 2819 131
rect 2804 128 2819 130
rect 2804 127 2805 128
rect 2799 126 2805 127
rect 2818 127 2819 128
rect 2823 127 2824 131
rect 2818 126 2824 127
rect 2935 131 2941 132
rect 2935 127 2936 131
rect 2940 130 2941 131
rect 2954 131 2960 132
rect 2954 130 2955 131
rect 2940 128 2955 130
rect 2940 127 2941 128
rect 2935 126 2941 127
rect 2954 127 2955 128
rect 2959 127 2960 131
rect 2954 126 2960 127
rect 3071 131 3077 132
rect 3071 127 3072 131
rect 3076 130 3077 131
rect 3090 131 3096 132
rect 3090 130 3091 131
rect 3076 128 3091 130
rect 3076 127 3077 128
rect 3071 126 3077 127
rect 3090 127 3091 128
rect 3095 127 3096 131
rect 3090 126 3096 127
rect 3207 131 3213 132
rect 3207 127 3208 131
rect 3212 130 3213 131
rect 3226 131 3232 132
rect 3226 130 3227 131
rect 3212 128 3227 130
rect 3212 127 3213 128
rect 3207 126 3213 127
rect 3226 127 3227 128
rect 3231 127 3232 131
rect 3226 126 3232 127
rect 3343 131 3349 132
rect 3343 127 3344 131
rect 3348 130 3349 131
rect 3362 131 3368 132
rect 3362 130 3363 131
rect 3348 128 3363 130
rect 3348 127 3349 128
rect 3343 126 3349 127
rect 3362 127 3363 128
rect 3367 127 3368 131
rect 3362 126 3368 127
rect 3479 131 3485 132
rect 3479 127 3480 131
rect 3484 130 3485 131
rect 3498 131 3504 132
rect 3498 130 3499 131
rect 3484 128 3499 130
rect 3484 127 3485 128
rect 3479 126 3485 127
rect 3498 127 3499 128
rect 3503 127 3504 131
rect 3498 126 3504 127
rect 3615 131 3621 132
rect 3615 127 3616 131
rect 3620 130 3621 131
rect 3634 131 3640 132
rect 3634 130 3635 131
rect 3620 128 3635 130
rect 3620 127 3621 128
rect 3615 126 3621 127
rect 3634 127 3635 128
rect 3639 127 3640 131
rect 3634 126 3640 127
rect 3646 131 3652 132
rect 3646 127 3647 131
rect 3651 130 3652 131
rect 3751 131 3757 132
rect 3751 130 3752 131
rect 3651 128 3752 130
rect 3651 127 3652 128
rect 3646 126 3652 127
rect 3751 127 3752 128
rect 3756 127 3757 131
rect 3751 126 3757 127
rect 110 122 116 123
rect 1934 122 1940 123
rect 1974 124 1980 125
rect 3798 124 3804 125
rect 4318 124 4324 125
rect 1974 120 1975 124
rect 1979 120 1980 124
rect 1974 119 1980 120
rect 1994 123 2000 124
rect 1994 119 1995 123
rect 1999 119 2000 123
rect 1994 118 2000 119
rect 2130 123 2136 124
rect 2130 119 2131 123
rect 2135 119 2136 123
rect 2130 118 2136 119
rect 2266 123 2272 124
rect 2266 119 2267 123
rect 2271 119 2272 123
rect 2266 118 2272 119
rect 2402 123 2408 124
rect 2402 119 2403 123
rect 2407 119 2408 123
rect 2402 118 2408 119
rect 2538 123 2544 124
rect 2538 119 2539 123
rect 2543 119 2544 123
rect 2538 118 2544 119
rect 2674 123 2680 124
rect 2674 119 2675 123
rect 2679 119 2680 123
rect 2674 118 2680 119
rect 2810 123 2816 124
rect 2810 119 2811 123
rect 2815 119 2816 123
rect 2810 118 2816 119
rect 2946 123 2952 124
rect 2946 119 2947 123
rect 2951 119 2952 123
rect 2946 118 2952 119
rect 3082 123 3088 124
rect 3082 119 3083 123
rect 3087 119 3088 123
rect 3082 118 3088 119
rect 3218 123 3224 124
rect 3218 119 3219 123
rect 3223 119 3224 123
rect 3218 118 3224 119
rect 3354 123 3360 124
rect 3354 119 3355 123
rect 3359 119 3360 123
rect 3354 118 3360 119
rect 3490 123 3496 124
rect 3490 119 3491 123
rect 3495 119 3496 123
rect 3490 118 3496 119
rect 3626 123 3632 124
rect 3626 119 3627 123
rect 3631 119 3632 123
rect 3798 120 3799 124
rect 3803 120 3804 124
rect 3798 119 3804 120
rect 3838 123 3844 124
rect 3838 119 3839 123
rect 3843 119 3844 123
rect 4318 120 4319 124
rect 4323 120 4324 124
rect 4318 119 4324 120
rect 4454 124 4460 125
rect 4454 120 4455 124
rect 4459 120 4460 124
rect 4454 119 4460 120
rect 4590 124 4596 125
rect 4590 120 4591 124
rect 4595 120 4596 124
rect 4590 119 4596 120
rect 4726 124 4732 125
rect 4726 120 4727 124
rect 4731 120 4732 124
rect 4726 119 4732 120
rect 4862 124 4868 125
rect 4862 120 4863 124
rect 4867 120 4868 124
rect 4862 119 4868 120
rect 4998 124 5004 125
rect 4998 120 4999 124
rect 5003 120 5004 124
rect 4998 119 5004 120
rect 5134 124 5140 125
rect 5134 120 5135 124
rect 5139 120 5140 124
rect 5134 119 5140 120
rect 5270 124 5276 125
rect 5270 120 5271 124
rect 5275 120 5276 124
rect 5270 119 5276 120
rect 5406 124 5412 125
rect 5406 120 5407 124
rect 5411 120 5412 124
rect 5406 119 5412 120
rect 5542 124 5548 125
rect 5542 120 5543 124
rect 5547 120 5548 124
rect 5542 119 5548 120
rect 5662 123 5668 124
rect 5662 119 5663 123
rect 5667 119 5668 123
rect 3626 118 3632 119
rect 3838 118 3844 119
rect 5662 118 5668 119
rect 2022 108 2028 109
rect 1974 107 1980 108
rect 1974 103 1975 107
rect 1979 103 1980 107
rect 2022 104 2023 108
rect 2027 104 2028 108
rect 2022 103 2028 104
rect 2158 108 2164 109
rect 2158 104 2159 108
rect 2163 104 2164 108
rect 2158 103 2164 104
rect 2294 108 2300 109
rect 2294 104 2295 108
rect 2299 104 2300 108
rect 2294 103 2300 104
rect 2430 108 2436 109
rect 2430 104 2431 108
rect 2435 104 2436 108
rect 2430 103 2436 104
rect 2566 108 2572 109
rect 2566 104 2567 108
rect 2571 104 2572 108
rect 2566 103 2572 104
rect 2702 108 2708 109
rect 2702 104 2703 108
rect 2707 104 2708 108
rect 2702 103 2708 104
rect 2838 108 2844 109
rect 2838 104 2839 108
rect 2843 104 2844 108
rect 2838 103 2844 104
rect 2974 108 2980 109
rect 2974 104 2975 108
rect 2979 104 2980 108
rect 2974 103 2980 104
rect 3110 108 3116 109
rect 3110 104 3111 108
rect 3115 104 3116 108
rect 3110 103 3116 104
rect 3246 108 3252 109
rect 3246 104 3247 108
rect 3251 104 3252 108
rect 3246 103 3252 104
rect 3382 108 3388 109
rect 3382 104 3383 108
rect 3387 104 3388 108
rect 3382 103 3388 104
rect 3518 108 3524 109
rect 3518 104 3519 108
rect 3523 104 3524 108
rect 3518 103 3524 104
rect 3654 108 3660 109
rect 3654 104 3655 108
rect 3659 104 3660 108
rect 3654 103 3660 104
rect 3798 107 3804 108
rect 3798 103 3799 107
rect 3803 103 3804 107
rect 1974 102 1980 103
rect 3798 102 3804 103
<< m3c >>
rect 111 5725 115 5729
rect 159 5724 163 5728
rect 295 5724 299 5728
rect 1935 5725 1939 5729
rect 111 5708 115 5712
rect 131 5709 135 5713
rect 267 5709 271 5713
rect 1935 5708 1939 5712
rect 379 5699 383 5703
rect 379 5631 383 5635
rect 283 5623 287 5627
rect 483 5623 487 5627
rect 707 5623 711 5627
rect 963 5623 967 5627
rect 1235 5623 1239 5627
rect 1779 5627 1783 5631
rect 1795 5623 1799 5627
rect 1975 5625 1979 5629
rect 2023 5624 2027 5628
rect 2183 5624 2187 5628
rect 2367 5624 2371 5628
rect 2551 5624 2555 5628
rect 2727 5624 2731 5628
rect 2895 5624 2899 5628
rect 3063 5624 3067 5628
rect 3223 5624 3227 5628
rect 3383 5624 3387 5628
rect 3543 5624 3547 5628
rect 3679 5624 3683 5628
rect 3799 5625 3803 5629
rect 3839 5621 3843 5625
rect 4335 5620 4339 5624
rect 4471 5620 4475 5624
rect 4607 5620 4611 5624
rect 4743 5620 4747 5624
rect 4879 5620 4883 5624
rect 5015 5620 5019 5624
rect 5663 5621 5667 5625
rect 1975 5608 1979 5612
rect 1995 5609 1999 5613
rect 2155 5609 2159 5613
rect 2339 5609 2343 5613
rect 2523 5609 2527 5613
rect 2699 5609 2703 5613
rect 2867 5609 2871 5613
rect 3035 5609 3039 5613
rect 3195 5609 3199 5613
rect 3355 5609 3359 5613
rect 3515 5609 3519 5613
rect 3651 5609 3655 5613
rect 3799 5608 3803 5612
rect 3839 5604 3843 5608
rect 4307 5605 4311 5609
rect 4443 5605 4447 5609
rect 4579 5605 4583 5609
rect 4715 5605 4719 5609
rect 4851 5605 4855 5609
rect 4987 5605 4991 5609
rect 5663 5604 5667 5608
rect 2143 5599 2147 5603
rect 2283 5599 2284 5603
rect 2284 5599 2287 5603
rect 2467 5599 2468 5603
rect 2468 5599 2471 5603
rect 2647 5599 2648 5603
rect 2648 5599 2651 5603
rect 2827 5599 2828 5603
rect 2828 5599 2831 5603
rect 2995 5599 2996 5603
rect 2996 5599 2999 5603
rect 3183 5599 3187 5603
rect 3343 5599 3347 5603
rect 3503 5599 3507 5603
rect 3643 5599 3644 5603
rect 3644 5599 3647 5603
rect 3739 5599 3743 5603
rect 4435 5595 4436 5599
rect 4436 5595 4439 5599
rect 4571 5595 4572 5599
rect 4572 5595 4575 5599
rect 4707 5595 4708 5599
rect 4708 5595 4711 5599
rect 4843 5595 4844 5599
rect 4844 5595 4847 5599
rect 4979 5595 4980 5599
rect 4980 5595 4983 5599
rect 5111 5595 5112 5599
rect 5112 5595 5115 5599
rect 283 5583 287 5587
rect 483 5583 487 5587
rect 707 5583 711 5587
rect 963 5583 967 5587
rect 1235 5583 1239 5587
rect 1279 5583 1283 5587
rect 1795 5583 1799 5587
rect 1963 5583 1967 5587
rect 111 5576 115 5580
rect 131 5575 135 5579
rect 275 5575 279 5579
rect 475 5575 479 5579
rect 699 5575 703 5579
rect 955 5575 959 5579
rect 1227 5575 1231 5579
rect 1515 5575 1519 5579
rect 1787 5575 1791 5579
rect 1935 5576 1939 5580
rect 111 5559 115 5563
rect 159 5560 163 5564
rect 303 5560 307 5564
rect 503 5560 507 5564
rect 727 5560 731 5564
rect 983 5560 987 5564
rect 1255 5560 1259 5564
rect 1543 5560 1547 5564
rect 1815 5560 1819 5564
rect 1935 5559 1939 5563
rect 1963 5559 1967 5563
rect 2143 5559 2147 5563
rect 2283 5559 2287 5563
rect 2467 5559 2471 5563
rect 2795 5559 2799 5563
rect 2827 5559 2831 5563
rect 2995 5559 2999 5563
rect 3183 5559 3187 5563
rect 3343 5559 3347 5563
rect 3503 5559 3507 5563
rect 3643 5559 3647 5563
rect 4375 5555 4379 5559
rect 4435 5555 4439 5559
rect 4571 5555 4575 5559
rect 4707 5555 4711 5559
rect 4843 5555 4847 5559
rect 4979 5555 4983 5559
rect 2647 5527 2651 5531
rect 3167 5527 3171 5531
rect 3635 5527 3639 5531
rect 3739 5527 3743 5531
rect 4575 5523 4579 5527
rect 4851 5523 4855 5527
rect 5111 5523 5115 5527
rect 111 5501 115 5505
rect 279 5500 283 5504
rect 519 5500 523 5504
rect 767 5500 771 5504
rect 1015 5500 1019 5504
rect 1263 5500 1267 5504
rect 1511 5500 1515 5504
rect 1767 5500 1771 5504
rect 1935 5501 1939 5505
rect 111 5484 115 5488
rect 251 5485 255 5489
rect 491 5485 495 5489
rect 739 5485 743 5489
rect 987 5485 991 5489
rect 1235 5485 1239 5489
rect 1483 5485 1487 5489
rect 1739 5485 1743 5489
rect 1935 5484 1939 5488
rect 2263 5483 2264 5487
rect 2264 5483 2267 5487
rect 2795 5483 2799 5487
rect 3327 5483 3331 5487
rect 3635 5483 3639 5487
rect 379 5475 380 5479
rect 380 5475 383 5479
rect 619 5475 620 5479
rect 620 5475 623 5479
rect 867 5475 868 5479
rect 868 5475 871 5479
rect 507 5467 511 5471
rect 1363 5475 1364 5479
rect 1364 5475 1367 5479
rect 1611 5475 1612 5479
rect 1612 5475 1615 5479
rect 1779 5475 1783 5479
rect 1975 5476 1979 5480
rect 2139 5475 2143 5479
rect 2355 5475 2359 5479
rect 2563 5475 2567 5479
rect 2755 5475 2759 5479
rect 2939 5475 2943 5479
rect 3115 5475 3119 5479
rect 3291 5475 3295 5479
rect 3467 5475 3471 5479
rect 3643 5475 3647 5479
rect 3799 5476 3803 5480
rect 4375 5479 4376 5483
rect 4376 5479 4379 5483
rect 4763 5479 4767 5483
rect 4851 5479 4855 5483
rect 3839 5472 3843 5476
rect 4251 5471 4255 5475
rect 4403 5471 4407 5475
rect 4555 5471 4559 5475
rect 4707 5471 4711 5475
rect 4859 5471 4863 5475
rect 5019 5471 5023 5475
rect 5663 5472 5667 5476
rect 1975 5459 1979 5463
rect 2167 5460 2171 5464
rect 2383 5460 2387 5464
rect 2591 5460 2595 5464
rect 2783 5460 2787 5464
rect 2967 5460 2971 5464
rect 3143 5460 3147 5464
rect 3319 5460 3323 5464
rect 3495 5460 3499 5464
rect 3671 5460 3675 5464
rect 3799 5459 3803 5463
rect 3839 5455 3843 5459
rect 4279 5456 4283 5460
rect 4431 5456 4435 5460
rect 4583 5456 4587 5460
rect 4735 5456 4739 5460
rect 4887 5456 4891 5460
rect 5047 5456 5051 5460
rect 5663 5455 5667 5459
rect 379 5435 383 5439
rect 619 5435 623 5439
rect 867 5435 871 5439
rect 1331 5435 1335 5439
rect 1363 5435 1367 5439
rect 1611 5435 1615 5439
rect 1279 5427 1283 5431
rect 507 5403 511 5407
rect 619 5399 623 5403
rect 827 5399 831 5403
rect 1043 5399 1047 5403
rect 1587 5399 1591 5403
rect 1975 5393 1979 5397
rect 2311 5392 2315 5396
rect 2511 5392 2515 5396
rect 2703 5392 2707 5396
rect 2887 5392 2891 5396
rect 3071 5392 3075 5396
rect 3247 5392 3251 5396
rect 3423 5392 3427 5396
rect 3607 5392 3611 5396
rect 3799 5393 3803 5397
rect 1975 5376 1979 5380
rect 2283 5377 2287 5381
rect 2483 5377 2487 5381
rect 2675 5377 2679 5381
rect 2859 5377 2863 5381
rect 3043 5377 3047 5381
rect 3219 5377 3223 5381
rect 3395 5377 3399 5381
rect 3579 5377 3583 5381
rect 3799 5376 3803 5380
rect 3839 5377 3843 5381
rect 4279 5376 4283 5380
rect 4487 5376 4491 5380
rect 4695 5376 4699 5380
rect 4911 5376 4915 5380
rect 5127 5376 5131 5380
rect 5663 5377 5667 5381
rect 659 5367 663 5371
rect 619 5359 623 5363
rect 827 5359 831 5363
rect 1043 5359 1047 5363
rect 2443 5367 2447 5371
rect 2611 5367 2612 5371
rect 2612 5367 2615 5371
rect 2811 5367 2815 5371
rect 2987 5367 2988 5371
rect 2988 5367 2991 5371
rect 3167 5367 3168 5371
rect 3168 5367 3171 5371
rect 3347 5367 3348 5371
rect 3348 5367 3351 5371
rect 3523 5367 3524 5371
rect 3524 5367 3527 5371
rect 3675 5367 3679 5371
rect 1331 5359 1335 5363
rect 3839 5360 3843 5364
rect 4251 5361 4255 5365
rect 4459 5361 4463 5365
rect 4667 5361 4671 5365
rect 4883 5361 4887 5365
rect 5099 5361 5103 5365
rect 5663 5360 5667 5364
rect 111 5352 115 5356
rect 411 5351 415 5355
rect 611 5351 615 5355
rect 819 5351 823 5355
rect 1035 5351 1039 5355
rect 1259 5351 1263 5355
rect 1491 5351 1495 5355
rect 1935 5352 1939 5356
rect 4419 5351 4423 5355
rect 4575 5351 4579 5355
rect 4807 5351 4811 5355
rect 5011 5351 5012 5355
rect 5012 5351 5015 5355
rect 5223 5351 5224 5355
rect 5224 5351 5227 5355
rect 111 5335 115 5339
rect 439 5336 443 5340
rect 639 5336 643 5340
rect 847 5336 851 5340
rect 1063 5336 1067 5340
rect 1287 5336 1291 5340
rect 1519 5336 1523 5340
rect 1935 5335 1939 5339
rect 2263 5327 2267 5331
rect 2443 5327 2447 5331
rect 2611 5327 2615 5331
rect 2955 5327 2959 5331
rect 2987 5327 2991 5331
rect 3327 5327 3331 5331
rect 3347 5327 3351 5331
rect 3523 5327 3527 5331
rect 4347 5311 4351 5315
rect 4419 5311 4423 5315
rect 4763 5311 4767 5315
rect 4807 5311 4811 5315
rect 5011 5311 5015 5315
rect 2331 5295 2335 5299
rect 2483 5295 2487 5299
rect 2803 5295 2807 5299
rect 2811 5295 2815 5299
rect 3195 5291 3199 5295
rect 3675 5295 3679 5299
rect 111 5277 115 5281
rect 591 5276 595 5280
rect 727 5276 731 5280
rect 863 5276 867 5280
rect 999 5276 1003 5280
rect 1135 5276 1139 5280
rect 1271 5276 1275 5280
rect 1407 5276 1411 5280
rect 1543 5276 1547 5280
rect 1935 5277 1939 5281
rect 111 5260 115 5264
rect 563 5261 567 5265
rect 699 5261 703 5265
rect 835 5261 839 5265
rect 971 5261 975 5265
rect 1107 5261 1111 5265
rect 1243 5261 1247 5265
rect 1379 5261 1383 5265
rect 1515 5261 1519 5265
rect 1935 5260 1939 5264
rect 4503 5263 4507 5267
rect 5223 5263 5227 5267
rect 691 5251 692 5255
rect 692 5251 695 5255
rect 827 5251 828 5255
rect 828 5251 831 5255
rect 963 5251 964 5255
rect 964 5251 967 5255
rect 1235 5251 1236 5255
rect 1236 5251 1239 5255
rect 1371 5251 1372 5255
rect 1372 5251 1375 5255
rect 1507 5251 1508 5255
rect 1508 5251 1511 5255
rect 1587 5251 1591 5255
rect 2319 5251 2320 5255
rect 2320 5251 2323 5255
rect 2331 5251 2335 5255
rect 2483 5251 2487 5255
rect 2803 5251 2807 5255
rect 2955 5251 2959 5255
rect 3355 5251 3359 5255
rect 1975 5244 1979 5248
rect 2195 5243 2199 5247
rect 2339 5243 2343 5247
rect 2491 5243 2495 5247
rect 2651 5243 2655 5247
rect 2819 5243 2823 5247
rect 3003 5243 3007 5247
rect 3187 5243 3191 5247
rect 3379 5243 3383 5247
rect 3579 5243 3583 5247
rect 3799 5244 3803 5248
rect 1975 5227 1979 5231
rect 2223 5228 2227 5232
rect 2367 5228 2371 5232
rect 2519 5228 2523 5232
rect 2679 5228 2683 5232
rect 2847 5228 2851 5232
rect 3031 5228 3035 5232
rect 3215 5228 3219 5232
rect 3407 5228 3411 5232
rect 3607 5228 3611 5232
rect 3799 5227 3803 5231
rect 4347 5219 4351 5223
rect 4843 5219 4844 5223
rect 4844 5219 4847 5223
rect 659 5211 663 5215
rect 691 5211 695 5215
rect 827 5211 831 5215
rect 963 5211 967 5215
rect 1235 5211 1239 5215
rect 1371 5211 1375 5215
rect 1507 5211 1511 5215
rect 3839 5212 3843 5216
rect 4251 5211 4255 5215
rect 4483 5211 4487 5215
rect 4715 5211 4719 5215
rect 4947 5211 4951 5215
rect 5187 5211 5191 5215
rect 5663 5212 5667 5216
rect 3839 5195 3843 5199
rect 4279 5196 4283 5200
rect 4511 5196 4515 5200
rect 4743 5196 4747 5200
rect 4975 5196 4979 5200
rect 5215 5196 5219 5200
rect 5663 5195 5667 5199
rect 1975 5169 1979 5173
rect 2023 5168 2027 5172
rect 2159 5168 2163 5172
rect 2327 5168 2331 5172
rect 2511 5168 2515 5172
rect 2695 5168 2699 5172
rect 2887 5168 2891 5172
rect 3087 5168 3091 5172
rect 3287 5168 3291 5172
rect 3495 5168 3499 5172
rect 3679 5168 3683 5172
rect 3799 5169 3803 5173
rect 1975 5152 1979 5156
rect 1995 5153 1999 5157
rect 2131 5153 2135 5157
rect 2299 5153 2303 5157
rect 2483 5153 2487 5157
rect 2667 5153 2671 5157
rect 2859 5153 2863 5157
rect 3059 5153 3063 5157
rect 3259 5153 3263 5157
rect 3467 5153 3471 5157
rect 3651 5153 3655 5157
rect 3799 5152 3803 5156
rect 2091 5143 2095 5147
rect 2139 5143 2143 5147
rect 2427 5143 2428 5147
rect 2428 5143 2431 5147
rect 2611 5143 2612 5147
rect 2612 5143 2615 5147
rect 2227 5135 2231 5139
rect 2999 5143 3003 5147
rect 3195 5143 3199 5147
rect 3427 5143 3431 5147
rect 3607 5143 3611 5147
rect 3747 5143 3751 5147
rect 2139 5111 2143 5115
rect 3839 5109 3843 5113
rect 3887 5108 3891 5112
rect 2227 5103 2231 5107
rect 2319 5103 2323 5107
rect 2427 5103 2431 5107
rect 2611 5103 2615 5107
rect 2999 5103 3003 5107
rect 3355 5103 3359 5107
rect 3427 5103 3431 5107
rect 4135 5108 4139 5112
rect 4407 5108 4411 5112
rect 4679 5108 4683 5112
rect 4959 5108 4963 5112
rect 5239 5108 5243 5112
rect 5663 5109 5667 5113
rect 3607 5103 3611 5107
rect 3839 5092 3843 5096
rect 3859 5093 3863 5097
rect 4107 5093 4111 5097
rect 4379 5093 4383 5097
rect 4651 5093 4655 5097
rect 4931 5093 4935 5097
rect 5211 5093 5215 5097
rect 5663 5092 5667 5096
rect 3955 5083 3959 5087
rect 4235 5083 4236 5087
rect 4236 5083 4239 5087
rect 4503 5083 4504 5087
rect 4504 5083 4507 5087
rect 443 5071 447 5075
rect 491 5071 495 5075
rect 1131 5071 1135 5075
rect 1223 5075 1227 5079
rect 1347 5071 1351 5075
rect 1587 5071 1591 5075
rect 1659 5071 1663 5075
rect 2119 5075 2123 5079
rect 2091 5067 2095 5071
rect 2955 5071 2959 5075
rect 3019 5071 3023 5075
rect 3747 5071 3751 5075
rect 4203 5075 4207 5079
rect 5059 5083 5060 5087
rect 5060 5083 5063 5087
rect 5335 5083 5336 5087
rect 5336 5083 5339 5087
rect 1131 5051 1135 5055
rect 1587 5051 1591 5055
rect 1911 5051 1915 5055
rect 443 5039 447 5043
rect 4203 5043 4207 5047
rect 4235 5043 4239 5047
rect 4747 5043 4751 5047
rect 4843 5043 4847 5047
rect 5059 5043 5063 5047
rect 491 5031 495 5035
rect 607 5031 608 5035
rect 608 5031 611 5035
rect 1347 5031 1351 5035
rect 1659 5031 1663 5035
rect 1779 5031 1780 5035
rect 1780 5031 1783 5035
rect 1911 5031 1912 5035
rect 1912 5031 1915 5035
rect 111 5024 115 5028
rect 347 5023 351 5027
rect 483 5023 487 5027
rect 619 5023 623 5027
rect 755 5023 759 5027
rect 891 5023 895 5027
rect 1035 5023 1039 5027
rect 1187 5023 1191 5027
rect 1339 5023 1343 5027
rect 1491 5023 1495 5027
rect 1651 5023 1655 5027
rect 1787 5023 1791 5027
rect 1935 5024 1939 5028
rect 2119 5027 2120 5031
rect 2120 5027 2123 5031
rect 2955 5027 2959 5031
rect 1975 5020 1979 5024
rect 1995 5019 1999 5023
rect 2531 5019 2535 5023
rect 3099 5019 3103 5023
rect 3651 5019 3655 5023
rect 3799 5020 3803 5024
rect 111 5007 115 5011
rect 375 5008 379 5012
rect 511 5008 515 5012
rect 647 5008 651 5012
rect 783 5008 787 5012
rect 919 5008 923 5012
rect 1063 5008 1067 5012
rect 1215 5008 1219 5012
rect 1367 5008 1371 5012
rect 1519 5008 1523 5012
rect 1679 5008 1683 5012
rect 1815 5008 1819 5012
rect 1935 5007 1939 5011
rect 1975 5003 1979 5007
rect 2023 5004 2027 5008
rect 2559 5004 2563 5008
rect 3127 5004 3131 5008
rect 3679 5004 3683 5008
rect 3799 5003 3803 5007
rect 3955 4999 3959 5003
rect 4819 5003 4823 5007
rect 4027 4995 4031 4999
rect 4219 4995 4223 4999
rect 4635 4995 4639 4999
rect 4851 4995 4855 4999
rect 5335 4999 5339 5003
rect 4027 4955 4031 4959
rect 4219 4955 4223 4959
rect 4335 4955 4336 4959
rect 4336 4955 4339 4959
rect 4635 4955 4639 4959
rect 4747 4955 4751 4959
rect 4819 4955 4823 4959
rect 5191 4955 5192 4959
rect 5192 4955 5195 4959
rect 111 4949 115 4953
rect 159 4948 163 4952
rect 343 4948 347 4952
rect 551 4948 555 4952
rect 751 4948 755 4952
rect 943 4948 947 4952
rect 1127 4948 1131 4952
rect 1311 4948 1315 4952
rect 1487 4948 1491 4952
rect 1663 4948 1667 4952
rect 1815 4948 1819 4952
rect 1935 4949 1939 4953
rect 3839 4948 3843 4952
rect 3859 4947 3863 4951
rect 4019 4947 4023 4951
rect 4211 4947 4215 4951
rect 4411 4947 4415 4951
rect 4627 4947 4631 4951
rect 4843 4947 4847 4951
rect 5067 4947 5071 4951
rect 5299 4947 5303 4951
rect 5663 4948 5667 4952
rect 111 4932 115 4936
rect 131 4933 135 4937
rect 315 4933 319 4937
rect 523 4933 527 4937
rect 723 4933 727 4937
rect 915 4933 919 4937
rect 1099 4933 1103 4937
rect 1283 4933 1287 4937
rect 1459 4933 1463 4937
rect 1635 4933 1639 4937
rect 1787 4933 1791 4937
rect 1935 4932 1939 4936
rect 3839 4931 3843 4935
rect 3887 4932 3891 4936
rect 4047 4932 4051 4936
rect 4239 4932 4243 4936
rect 4439 4932 4443 4936
rect 4655 4932 4659 4936
rect 4871 4932 4875 4936
rect 5095 4932 5099 4936
rect 5327 4932 5331 4936
rect 5663 4931 5667 4935
rect 227 4923 231 4927
rect 275 4923 279 4927
rect 687 4923 691 4927
rect 411 4915 415 4919
rect 1071 4923 1075 4927
rect 1223 4923 1224 4927
rect 1224 4923 1227 4927
rect 1011 4915 1015 4919
rect 1435 4923 1439 4927
rect 1611 4923 1615 4927
rect 1771 4923 1775 4927
rect 1975 4913 1979 4917
rect 2871 4912 2875 4916
rect 3007 4912 3011 4916
rect 3799 4913 3803 4917
rect 1975 4896 1979 4900
rect 2843 4897 2847 4901
rect 2979 4897 2983 4901
rect 3799 4896 3803 4900
rect 275 4883 279 4887
rect 411 4883 415 4887
rect 607 4883 611 4887
rect 687 4883 691 4887
rect 1011 4883 1015 4887
rect 1071 4883 1075 4887
rect 1435 4883 1439 4887
rect 1611 4883 1615 4887
rect 1771 4883 1775 4887
rect 1779 4883 1783 4887
rect 3019 4887 3023 4891
rect 2939 4879 2943 4883
rect 3839 4853 3843 4857
rect 3887 4852 3891 4856
rect 227 4843 231 4847
rect 2939 4847 2943 4851
rect 4071 4852 4075 4856
rect 4287 4852 4291 4856
rect 4511 4852 4515 4856
rect 4735 4852 4739 4856
rect 4959 4852 4963 4856
rect 5183 4852 5187 4856
rect 5407 4852 5411 4856
rect 5663 4853 5667 4857
rect 3147 4847 3151 4851
rect 275 4839 279 4843
rect 411 4839 415 4843
rect 547 4839 551 4843
rect 683 4839 687 4843
rect 3839 4836 3843 4840
rect 3859 4837 3863 4841
rect 4043 4837 4047 4841
rect 4259 4837 4263 4841
rect 4483 4837 4487 4841
rect 4707 4837 4711 4841
rect 4931 4837 4935 4841
rect 5155 4837 5159 4841
rect 5379 4837 5383 4841
rect 5663 4836 5667 4840
rect 3983 4827 3984 4831
rect 3984 4827 3987 4831
rect 4611 4827 4612 4831
rect 4612 4827 4615 4831
rect 4851 4827 4855 4831
rect 4579 4819 4583 4823
rect 5467 4827 5471 4831
rect 275 4799 279 4803
rect 411 4799 415 4803
rect 547 4799 551 4803
rect 683 4799 687 4803
rect 691 4799 695 4803
rect 111 4792 115 4796
rect 131 4791 135 4795
rect 267 4791 271 4795
rect 403 4791 407 4795
rect 539 4791 543 4795
rect 675 4791 679 4795
rect 1935 4792 1939 4796
rect 1967 4791 1971 4795
rect 2163 4787 2167 4791
rect 2355 4787 2359 4791
rect 2547 4787 2551 4791
rect 2791 4791 2795 4795
rect 2939 4787 2943 4791
rect 3139 4787 3143 4791
rect 4335 4787 4339 4791
rect 4579 4787 4583 4791
rect 4611 4787 4615 4791
rect 5083 4787 5087 4791
rect 5191 4787 5195 4791
rect 111 4775 115 4779
rect 159 4776 163 4780
rect 295 4776 299 4780
rect 431 4776 435 4780
rect 567 4776 571 4780
rect 703 4776 707 4780
rect 1935 4775 1939 4779
rect 2163 4747 2167 4751
rect 2355 4747 2359 4751
rect 2547 4747 2551 4751
rect 2659 4747 2663 4751
rect 2939 4747 2943 4751
rect 3139 4747 3143 4751
rect 3147 4747 3151 4751
rect 3983 4751 3987 4755
rect 4195 4747 4199 4751
rect 4475 4747 4479 4751
rect 4859 4747 4863 4751
rect 5075 4747 5079 4751
rect 5467 4751 5471 4755
rect 227 4739 231 4743
rect 691 4739 695 4743
rect 1975 4740 1979 4744
rect 1995 4739 1999 4743
rect 2155 4739 2159 4743
rect 2347 4739 2351 4743
rect 2539 4739 2543 4743
rect 2731 4739 2735 4743
rect 2931 4739 2935 4743
rect 3131 4739 3135 4743
rect 3799 4740 3803 4744
rect 1975 4723 1979 4727
rect 2023 4724 2027 4728
rect 2183 4724 2187 4728
rect 2375 4724 2379 4728
rect 2567 4724 2571 4728
rect 2759 4724 2763 4728
rect 2959 4724 2963 4728
rect 3159 4724 3163 4728
rect 3799 4723 3803 4727
rect 111 4709 115 4713
rect 159 4708 163 4712
rect 343 4708 347 4712
rect 567 4708 571 4712
rect 807 4708 811 4712
rect 1055 4708 1059 4712
rect 1311 4708 1315 4712
rect 1575 4708 1579 4712
rect 1815 4708 1819 4712
rect 1935 4709 1939 4713
rect 4195 4707 4199 4711
rect 4475 4707 4479 4711
rect 4591 4707 4592 4711
rect 4592 4707 4595 4711
rect 5075 4707 5079 4711
rect 5083 4707 5087 4711
rect 5495 4707 5496 4711
rect 5496 4707 5499 4711
rect 3839 4700 3843 4704
rect 3915 4699 3919 4703
rect 4187 4699 4191 4703
rect 4467 4699 4471 4703
rect 4763 4699 4767 4703
rect 5067 4699 5071 4703
rect 5371 4699 5375 4703
rect 5663 4700 5667 4704
rect 111 4692 115 4696
rect 131 4693 135 4697
rect 315 4693 319 4697
rect 539 4693 543 4697
rect 779 4693 783 4697
rect 1027 4693 1031 4697
rect 1283 4693 1287 4697
rect 1547 4693 1551 4697
rect 1787 4693 1791 4697
rect 1935 4692 1939 4696
rect 443 4683 444 4687
rect 444 4683 447 4687
rect 667 4683 668 4687
rect 668 4683 671 4687
rect 907 4683 908 4687
rect 908 4683 911 4687
rect 1011 4683 1015 4687
rect 1411 4683 1412 4687
rect 1412 4683 1415 4687
rect 1675 4683 1676 4687
rect 1676 4683 1679 4687
rect 1967 4683 1971 4687
rect 3839 4683 3843 4687
rect 3943 4684 3947 4688
rect 4215 4684 4219 4688
rect 4495 4684 4499 4688
rect 4791 4684 4795 4688
rect 5095 4684 5099 4688
rect 5399 4684 5403 4688
rect 5663 4683 5667 4687
rect 1975 4661 1979 4665
rect 2023 4660 2027 4664
rect 2239 4660 2243 4664
rect 2471 4660 2475 4664
rect 2695 4660 2699 4664
rect 2919 4660 2923 4664
rect 3143 4660 3147 4664
rect 3367 4660 3371 4664
rect 3799 4661 3803 4665
rect 227 4643 231 4647
rect 443 4643 447 4647
rect 667 4643 671 4647
rect 907 4643 911 4647
rect 1411 4643 1415 4647
rect 1675 4643 1679 4647
rect 1975 4644 1979 4648
rect 1995 4645 1999 4649
rect 2211 4645 2215 4649
rect 2443 4645 2447 4649
rect 2667 4645 2671 4649
rect 2891 4645 2895 4649
rect 3115 4645 3119 4649
rect 3339 4645 3343 4649
rect 3799 4644 3803 4648
rect 1519 4635 1523 4639
rect 2339 4635 2340 4639
rect 2340 4635 2343 4639
rect 2791 4635 2792 4639
rect 2792 4635 2795 4639
rect 2883 4635 2887 4639
rect 3243 4635 3244 4639
rect 3244 4635 3247 4639
rect 2987 4627 2991 4631
rect 3839 4625 3843 4629
rect 4063 4624 4067 4628
rect 4327 4624 4331 4628
rect 4599 4624 4603 4628
rect 4871 4624 4875 4628
rect 5151 4624 5155 4628
rect 5439 4624 5443 4628
rect 5663 4625 5667 4629
rect 3839 4608 3843 4612
rect 4035 4609 4039 4613
rect 4299 4609 4303 4613
rect 4571 4609 4575 4613
rect 4843 4609 4847 4613
rect 5123 4609 5127 4613
rect 5411 4609 5415 4613
rect 5663 4608 5667 4612
rect 1011 4599 1015 4603
rect 1907 4599 1911 4603
rect 403 4591 407 4595
rect 651 4591 655 4595
rect 915 4591 919 4595
rect 1203 4591 1207 4595
rect 1795 4591 1799 4595
rect 2339 4595 2343 4599
rect 2883 4595 2887 4599
rect 2987 4595 2991 4599
rect 3127 4595 3131 4599
rect 3243 4595 3247 4599
rect 4171 4599 4175 4603
rect 4543 4599 4547 4603
rect 4859 4599 4863 4603
rect 5067 4599 5071 4603
rect 5535 4599 5536 4603
rect 5536 4599 5539 4603
rect 2659 4587 2663 4591
rect 403 4551 407 4555
rect 651 4551 655 4555
rect 915 4551 919 4555
rect 1203 4551 1207 4555
rect 1231 4551 1235 4555
rect 1519 4551 1523 4555
rect 1907 4551 1911 4555
rect 2891 4555 2895 4559
rect 3011 4555 3015 4559
rect 3707 4555 3711 4559
rect 4543 4559 4547 4563
rect 4591 4559 4595 4563
rect 5067 4559 5071 4563
rect 5219 4559 5223 4563
rect 5495 4559 5499 4563
rect 111 4544 115 4548
rect 171 4543 175 4547
rect 395 4543 399 4547
rect 643 4543 647 4547
rect 907 4543 911 4547
rect 1195 4543 1199 4547
rect 1491 4543 1495 4547
rect 1787 4543 1791 4547
rect 1935 4544 1939 4548
rect 111 4527 115 4531
rect 199 4528 203 4532
rect 423 4528 427 4532
rect 671 4528 675 4532
rect 935 4528 939 4532
rect 1223 4528 1227 4532
rect 1519 4528 1523 4532
rect 1815 4528 1819 4532
rect 1935 4527 1939 4531
rect 2891 4523 2895 4527
rect 4171 4527 4175 4531
rect 2223 4515 2224 4519
rect 2224 4515 2227 4519
rect 3011 4515 3015 4519
rect 3127 4515 3128 4519
rect 3128 4515 3131 4519
rect 4419 4523 4423 4527
rect 4667 4523 4671 4527
rect 4975 4527 4979 4531
rect 5187 4523 5191 4527
rect 5535 4527 5539 4531
rect 1975 4508 1979 4512
rect 2099 4507 2103 4511
rect 2347 4507 2351 4511
rect 2579 4507 2583 4511
rect 2795 4507 2799 4511
rect 3003 4507 3007 4511
rect 3203 4507 3207 4511
rect 3403 4507 3407 4511
rect 3611 4507 3615 4511
rect 3799 4508 3803 4512
rect 1975 4491 1979 4495
rect 2127 4492 2131 4496
rect 2375 4492 2379 4496
rect 2607 4492 2611 4496
rect 2823 4492 2827 4496
rect 3031 4492 3035 4496
rect 3231 4492 3235 4496
rect 3431 4492 3435 4496
rect 3639 4492 3643 4496
rect 3799 4491 3803 4495
rect 4419 4483 4423 4487
rect 4667 4483 4671 4487
rect 4755 4483 4759 4487
rect 5187 4483 5191 4487
rect 5219 4483 5223 4487
rect 5567 4483 5568 4487
rect 5568 4483 5571 4487
rect 3839 4476 3843 4480
rect 4179 4475 4183 4479
rect 4411 4475 4415 4479
rect 4659 4475 4663 4479
rect 4915 4475 4919 4479
rect 5179 4475 5183 4479
rect 5443 4475 5447 4479
rect 5663 4476 5667 4480
rect 111 4465 115 4469
rect 447 4464 451 4468
rect 655 4464 659 4468
rect 887 4464 891 4468
rect 1143 4464 1147 4468
rect 1407 4464 1411 4468
rect 1679 4464 1683 4468
rect 1935 4465 1939 4469
rect 3839 4459 3843 4463
rect 4207 4460 4211 4464
rect 4439 4460 4443 4464
rect 4687 4460 4691 4464
rect 4943 4460 4947 4464
rect 5207 4460 5211 4464
rect 5471 4460 5475 4464
rect 5663 4459 5667 4463
rect 111 4448 115 4452
rect 419 4449 423 4453
rect 627 4449 631 4453
rect 859 4449 863 4453
rect 1115 4449 1119 4453
rect 1379 4449 1383 4453
rect 1651 4449 1655 4453
rect 1935 4448 1939 4452
rect 587 4439 591 4443
rect 755 4439 756 4443
rect 756 4439 759 4443
rect 1079 4439 1083 4443
rect 1243 4439 1244 4443
rect 1244 4439 1247 4443
rect 1275 4439 1279 4443
rect 1795 4439 1799 4443
rect 515 4431 519 4435
rect 1231 4431 1235 4435
rect 1975 4425 1979 4429
rect 2231 4424 2235 4428
rect 2447 4424 2451 4428
rect 2663 4424 2667 4428
rect 2871 4424 2875 4428
rect 3079 4424 3083 4428
rect 3287 4424 3291 4428
rect 3495 4424 3499 4428
rect 3679 4424 3683 4428
rect 3799 4425 3803 4429
rect 1975 4408 1979 4412
rect 2203 4409 2207 4413
rect 2419 4409 2423 4413
rect 2635 4409 2639 4413
rect 2843 4409 2847 4413
rect 3051 4409 3055 4413
rect 3259 4409 3263 4413
rect 3467 4409 3471 4413
rect 3651 4409 3655 4413
rect 3799 4408 3803 4412
rect 515 4399 519 4403
rect 587 4399 591 4403
rect 755 4399 759 4403
rect 1079 4399 1083 4403
rect 1243 4399 1247 4403
rect 1747 4399 1751 4403
rect 2331 4399 2332 4403
rect 2332 4399 2335 4403
rect 2547 4399 2548 4403
rect 2548 4399 2551 4403
rect 2787 4399 2791 4403
rect 2915 4399 2919 4403
rect 3191 4399 3195 4403
rect 3431 4399 3435 4403
rect 3607 4399 3611 4403
rect 3707 4399 3711 4403
rect 3839 4393 3843 4397
rect 4359 4392 4363 4396
rect 4519 4392 4523 4396
rect 4687 4392 4691 4396
rect 4879 4392 4883 4396
rect 5079 4392 5083 4396
rect 5287 4392 5291 4396
rect 5503 4392 5507 4396
rect 5663 4393 5667 4397
rect 3839 4376 3843 4380
rect 4331 4377 4335 4381
rect 4491 4377 4495 4381
rect 4659 4377 4663 4381
rect 4851 4377 4855 4381
rect 5051 4377 5055 4381
rect 5259 4377 5263 4381
rect 5475 4377 5479 4381
rect 5663 4376 5667 4380
rect 1275 4367 1279 4371
rect 4347 4367 4351 4371
rect 4483 4367 4487 4371
rect 4975 4367 4976 4371
rect 4976 4367 4979 4371
rect 5011 4367 5015 4371
rect 5595 4367 5599 4371
rect 819 4359 823 4363
rect 971 4359 975 4363
rect 1131 4359 1135 4363
rect 1299 4359 1303 4363
rect 1563 4359 1567 4363
rect 1659 4359 1663 4363
rect 2223 4359 2227 4363
rect 2331 4359 2335 4363
rect 2547 4359 2551 4363
rect 2787 4359 2791 4363
rect 3191 4359 3195 4363
rect 3431 4359 3435 4363
rect 3607 4359 3611 4363
rect 3439 4351 3443 4355
rect 819 4319 823 4323
rect 971 4319 975 4323
rect 1131 4319 1135 4323
rect 1299 4319 1303 4323
rect 1307 4319 1311 4323
rect 1659 4319 1663 4323
rect 1747 4319 1751 4323
rect 2915 4323 2919 4327
rect 4483 4327 4487 4331
rect 4755 4327 4759 4331
rect 5011 4327 5015 4331
rect 5355 4327 5359 4331
rect 5567 4327 5571 4331
rect 111 4312 115 4316
rect 667 4311 671 4315
rect 811 4311 815 4315
rect 963 4311 967 4315
rect 1123 4311 1127 4315
rect 1291 4311 1295 4315
rect 1467 4311 1471 4315
rect 1651 4311 1655 4315
rect 1935 4312 1939 4316
rect 2467 4315 2471 4319
rect 2635 4315 2639 4319
rect 2819 4315 2823 4319
rect 3019 4315 3023 4319
rect 3235 4315 3239 4319
rect 3643 4319 3647 4323
rect 3983 4319 3987 4323
rect 111 4295 115 4299
rect 695 4296 699 4300
rect 839 4296 843 4300
rect 991 4296 995 4300
rect 1151 4296 1155 4300
rect 1319 4296 1323 4300
rect 1495 4296 1499 4300
rect 1679 4296 1683 4300
rect 1935 4295 1939 4299
rect 4051 4291 4055 4295
rect 4347 4295 4351 4299
rect 4483 4291 4487 4295
rect 4723 4291 4727 4295
rect 4979 4291 4983 4295
rect 5243 4291 5247 4295
rect 5595 4295 5599 4299
rect 2467 4275 2471 4279
rect 2635 4275 2639 4279
rect 2819 4275 2823 4279
rect 3019 4275 3023 4279
rect 3235 4275 3239 4279
rect 3351 4275 3352 4279
rect 3352 4275 3355 4279
rect 3439 4275 3443 4279
rect 3643 4275 3647 4279
rect 1975 4268 1979 4272
rect 2307 4267 2311 4271
rect 2459 4267 2463 4271
rect 2627 4267 2631 4271
rect 2811 4267 2815 4271
rect 3011 4267 3015 4271
rect 3227 4267 3231 4271
rect 3451 4267 3455 4271
rect 3651 4267 3655 4271
rect 3799 4268 3803 4272
rect 1975 4251 1979 4255
rect 2335 4252 2339 4256
rect 2487 4252 2491 4256
rect 2655 4252 2659 4256
rect 2839 4252 2843 4256
rect 3039 4252 3043 4256
rect 3255 4252 3259 4256
rect 3479 4252 3483 4256
rect 3679 4252 3683 4256
rect 3799 4251 3803 4255
rect 3983 4251 3984 4255
rect 3984 4251 3987 4255
rect 4483 4251 4487 4255
rect 4723 4251 4727 4255
rect 4979 4251 4983 4255
rect 5243 4251 5247 4255
rect 5355 4251 5359 4255
rect 5611 4251 5615 4255
rect 3839 4244 3843 4248
rect 3859 4243 3863 4247
rect 4043 4243 4047 4247
rect 4251 4243 4255 4247
rect 4475 4243 4479 4247
rect 4715 4243 4719 4247
rect 4971 4243 4975 4247
rect 5235 4243 5239 4247
rect 5499 4243 5503 4247
rect 5663 4244 5667 4248
rect 3839 4227 3843 4231
rect 3887 4228 3891 4232
rect 4071 4228 4075 4232
rect 4279 4228 4283 4232
rect 4503 4228 4507 4232
rect 4743 4228 4747 4232
rect 4999 4228 5003 4232
rect 5263 4228 5267 4232
rect 5527 4228 5531 4232
rect 5663 4227 5667 4231
rect 111 4221 115 4225
rect 815 4220 819 4224
rect 951 4220 955 4224
rect 1087 4220 1091 4224
rect 1223 4220 1227 4224
rect 1359 4220 1363 4224
rect 1495 4220 1499 4224
rect 1631 4220 1635 4224
rect 1767 4220 1771 4224
rect 1935 4221 1939 4225
rect 111 4204 115 4208
rect 787 4205 791 4209
rect 923 4205 927 4209
rect 1059 4205 1063 4209
rect 1195 4205 1199 4209
rect 1331 4205 1335 4209
rect 1467 4205 1471 4209
rect 1603 4205 1607 4209
rect 1739 4205 1743 4209
rect 1935 4204 1939 4208
rect 915 4195 916 4199
rect 916 4195 919 4199
rect 1051 4195 1052 4199
rect 1052 4195 1055 4199
rect 1187 4195 1188 4199
rect 1188 4195 1191 4199
rect 1323 4195 1324 4199
rect 1324 4195 1327 4199
rect 1379 4195 1383 4199
rect 1563 4195 1567 4199
rect 1731 4195 1732 4199
rect 1732 4195 1735 4199
rect 1563 4187 1567 4191
rect 1975 4185 1979 4189
rect 2567 4184 2571 4188
rect 2703 4184 2707 4188
rect 2839 4184 2843 4188
rect 2975 4184 2979 4188
rect 3799 4185 3803 4189
rect 1975 4168 1979 4172
rect 2539 4169 2543 4173
rect 2675 4169 2679 4173
rect 2811 4169 2815 4173
rect 2947 4169 2951 4173
rect 3799 4168 3803 4172
rect 915 4155 919 4159
rect 1051 4155 1055 4159
rect 1187 4155 1191 4159
rect 1323 4155 1327 4159
rect 1563 4155 1567 4159
rect 1671 4155 1675 4159
rect 1731 4155 1735 4159
rect 2659 4159 2663 4163
rect 2955 4159 2959 4163
rect 1307 4147 1311 4151
rect 3839 4133 3843 4137
rect 3887 4132 3891 4136
rect 4415 4132 4419 4136
rect 4975 4132 4979 4136
rect 5543 4132 5547 4136
rect 5663 4133 5667 4137
rect 1379 4123 1383 4127
rect 1099 4115 1103 4119
rect 1371 4115 1375 4119
rect 1419 4115 1423 4119
rect 1555 4115 1559 4119
rect 2955 4127 2959 4131
rect 3351 4119 3355 4123
rect 3839 4116 3843 4120
rect 3859 4117 3863 4121
rect 4387 4117 4391 4121
rect 4947 4117 4951 4121
rect 5515 4117 5519 4121
rect 5663 4116 5667 4120
rect 4051 4107 4055 4111
rect 4879 4107 4883 4111
rect 3955 4099 3959 4103
rect 5619 4107 5623 4111
rect 1099 4083 1103 4087
rect 855 4075 856 4079
rect 856 4075 859 4079
rect 1419 4075 1423 4079
rect 1555 4075 1559 4079
rect 1671 4075 1672 4079
rect 1672 4075 1675 4079
rect 111 4068 115 4072
rect 731 4067 735 4071
rect 867 4067 871 4071
rect 1003 4067 1007 4071
rect 1139 4067 1143 4071
rect 1275 4067 1279 4071
rect 1411 4067 1415 4071
rect 1547 4067 1551 4071
rect 1935 4068 1939 4072
rect 2387 4063 2391 4067
rect 2435 4063 2439 4067
rect 2659 4067 2663 4071
rect 2707 4063 2711 4067
rect 2843 4063 2847 4067
rect 3955 4067 3959 4071
rect 4879 4067 4883 4071
rect 5611 4067 5615 4071
rect 111 4051 115 4055
rect 759 4052 763 4056
rect 895 4052 899 4056
rect 1031 4052 1035 4056
rect 1167 4052 1171 4056
rect 1303 4052 1307 4056
rect 1439 4052 1443 4056
rect 1575 4052 1579 4056
rect 1935 4051 1939 4055
rect 3867 4031 3871 4035
rect 4011 4031 4015 4035
rect 4179 4031 4183 4035
rect 5399 4035 5403 4039
rect 5619 4035 5623 4039
rect 2435 4023 2439 4027
rect 2551 4023 2552 4027
rect 2552 4023 2555 4027
rect 2707 4023 2711 4027
rect 2843 4023 2847 4027
rect 2959 4023 2960 4027
rect 2960 4023 2963 4027
rect 1975 4016 1979 4020
rect 2291 4015 2295 4019
rect 2427 4015 2431 4019
rect 2563 4015 2567 4019
rect 2699 4015 2703 4019
rect 2835 4015 2839 4019
rect 3799 4016 3803 4020
rect 1975 3999 1979 4003
rect 2319 4000 2323 4004
rect 2455 4000 2459 4004
rect 2591 4000 2595 4004
rect 2727 4000 2731 4004
rect 2863 4000 2867 4004
rect 3799 3999 3803 4003
rect 4011 3991 4015 3995
rect 4179 3991 4183 3995
rect 4451 3991 4455 3995
rect 5635 3991 5639 3995
rect 3839 3984 3843 3988
rect 3859 3983 3863 3987
rect 4003 3983 4007 3987
rect 4171 3983 4175 3987
rect 4339 3983 4343 3987
rect 4499 3983 4503 3987
rect 4651 3983 4655 3987
rect 4803 3983 4807 3987
rect 4947 3983 4951 3987
rect 5091 3983 5095 3987
rect 5235 3983 5239 3987
rect 5379 3983 5383 3987
rect 5515 3983 5519 3987
rect 5663 3984 5667 3988
rect 111 3969 115 3973
rect 511 3968 515 3972
rect 663 3968 667 3972
rect 823 3968 827 3972
rect 983 3968 987 3972
rect 1151 3968 1155 3972
rect 1319 3968 1323 3972
rect 1935 3969 1939 3973
rect 3839 3967 3843 3971
rect 3887 3968 3891 3972
rect 4031 3968 4035 3972
rect 4199 3968 4203 3972
rect 4367 3968 4371 3972
rect 4527 3968 4531 3972
rect 4679 3968 4683 3972
rect 4831 3968 4835 3972
rect 4975 3968 4979 3972
rect 5119 3968 5123 3972
rect 5263 3968 5267 3972
rect 5407 3968 5411 3972
rect 5543 3968 5547 3972
rect 5663 3967 5667 3971
rect 111 3952 115 3956
rect 483 3953 487 3957
rect 635 3953 639 3957
rect 795 3953 799 3957
rect 955 3953 959 3957
rect 1123 3953 1127 3957
rect 1291 3953 1295 3957
rect 1935 3952 1939 3956
rect 611 3943 612 3947
rect 612 3943 615 3947
rect 759 3943 760 3947
rect 760 3943 763 3947
rect 943 3943 947 3947
rect 579 3935 583 3939
rect 1251 3943 1252 3947
rect 1252 3943 1255 3947
rect 1371 3943 1375 3947
rect 1975 3937 1979 3941
rect 2119 3936 2123 3940
rect 2327 3936 2331 3940
rect 2535 3936 2539 3940
rect 2743 3936 2747 3940
rect 2943 3936 2947 3940
rect 3135 3936 3139 3940
rect 3319 3936 3323 3940
rect 3511 3936 3515 3940
rect 3679 3936 3683 3940
rect 3799 3937 3803 3941
rect 1975 3920 1979 3924
rect 2091 3921 2095 3925
rect 2299 3921 2303 3925
rect 2507 3921 2511 3925
rect 2715 3921 2719 3925
rect 2915 3921 2919 3925
rect 3107 3921 3111 3925
rect 3291 3921 3295 3925
rect 3483 3921 3487 3925
rect 3651 3921 3655 3925
rect 3799 3920 3803 3924
rect 2215 3911 2216 3915
rect 2216 3911 2219 3915
rect 2291 3911 2295 3915
rect 579 3903 583 3907
rect 611 3903 615 3907
rect 855 3903 859 3907
rect 943 3903 947 3907
rect 1219 3903 1223 3907
rect 1251 3903 1255 3907
rect 2395 3903 2399 3907
rect 3043 3911 3044 3915
rect 3044 3911 3047 3915
rect 3235 3911 3236 3915
rect 3236 3911 3239 3915
rect 3419 3911 3420 3915
rect 3420 3911 3423 3915
rect 3611 3911 3612 3915
rect 3612 3911 3615 3915
rect 3867 3911 3871 3915
rect 3839 3885 3843 3889
rect 4383 3884 4387 3888
rect 4599 3884 4603 3888
rect 4823 3884 4827 3888
rect 5063 3884 5067 3888
rect 5311 3884 5315 3888
rect 5543 3884 5547 3888
rect 5663 3885 5667 3889
rect 2291 3871 2295 3875
rect 2395 3871 2399 3875
rect 2551 3871 2555 3875
rect 3011 3871 3015 3875
rect 3043 3871 3047 3875
rect 3235 3871 3239 3875
rect 3419 3871 3423 3875
rect 3611 3871 3615 3875
rect 3839 3868 3843 3872
rect 4355 3869 4359 3873
rect 4571 3869 4575 3873
rect 4795 3869 4799 3873
rect 5035 3869 5039 3873
rect 5283 3869 5287 3873
rect 5515 3869 5519 3873
rect 5663 3868 5667 3872
rect 4483 3859 4484 3863
rect 4484 3859 4487 3863
rect 4699 3859 4700 3863
rect 4700 3859 4703 3863
rect 4923 3859 4924 3863
rect 4924 3859 4927 3863
rect 5059 3859 5063 3863
rect 5399 3859 5403 3863
rect 5611 3859 5615 3863
rect 627 3851 631 3855
rect 315 3839 319 3843
rect 759 3843 763 3847
rect 1151 3843 1155 3847
rect 1171 3839 1175 3843
rect 2215 3827 2219 3831
rect 2379 3823 2383 3827
rect 2595 3823 2599 3827
rect 2803 3823 2807 3827
rect 3003 3823 3007 3827
rect 3203 3823 3207 3827
rect 3411 3823 3415 3827
rect 4451 3819 4455 3823
rect 4483 3819 4487 3823
rect 4699 3819 4703 3823
rect 4923 3819 4927 3823
rect 5375 3819 5379 3823
rect 5635 3819 5639 3823
rect 315 3799 319 3803
rect 403 3799 407 3803
rect 627 3799 631 3803
rect 1171 3799 1175 3803
rect 1219 3799 1223 3803
rect 111 3792 115 3796
rect 131 3791 135 3795
rect 307 3791 311 3795
rect 515 3791 519 3795
rect 723 3791 727 3795
rect 939 3791 943 3795
rect 1163 3791 1167 3795
rect 1935 3792 1939 3796
rect 2379 3783 2383 3787
rect 2391 3783 2395 3787
rect 2803 3783 2807 3787
rect 3003 3783 3007 3787
rect 3203 3783 3207 3787
rect 3411 3783 3415 3787
rect 3419 3783 3423 3787
rect 111 3775 115 3779
rect 159 3776 163 3780
rect 335 3776 339 3780
rect 543 3776 547 3780
rect 751 3776 755 3780
rect 967 3776 971 3780
rect 1191 3776 1195 3780
rect 1935 3775 1939 3779
rect 1975 3776 1979 3780
rect 2139 3775 2143 3779
rect 2371 3775 2375 3779
rect 2587 3775 2591 3779
rect 2795 3775 2799 3779
rect 2995 3775 2999 3779
rect 3195 3775 3199 3779
rect 3403 3775 3407 3779
rect 3799 3776 3803 3780
rect 4091 3767 4095 3771
rect 4211 3767 4215 3771
rect 4443 3767 4447 3771
rect 4699 3767 4703 3771
rect 5059 3771 5063 3775
rect 5347 3767 5351 3771
rect 5611 3771 5615 3775
rect 1975 3759 1979 3763
rect 2167 3760 2171 3764
rect 2399 3760 2403 3764
rect 2615 3760 2619 3764
rect 2823 3760 2827 3764
rect 3023 3760 3027 3764
rect 3223 3760 3227 3764
rect 3431 3760 3435 3764
rect 3799 3759 3803 3763
rect 4211 3727 4215 3731
rect 4443 3727 4447 3731
rect 4699 3727 4703 3731
rect 4815 3727 4816 3731
rect 4816 3727 4819 3731
rect 4939 3727 4943 3731
rect 5375 3727 5376 3731
rect 5376 3727 5379 3731
rect 5627 3727 5631 3731
rect 111 3717 115 3721
rect 159 3716 163 3720
rect 335 3716 339 3720
rect 527 3716 531 3720
rect 711 3716 715 3720
rect 887 3716 891 3720
rect 1055 3716 1059 3720
rect 1215 3716 1219 3720
rect 1367 3716 1371 3720
rect 1519 3716 1523 3720
rect 1679 3716 1683 3720
rect 1815 3716 1819 3720
rect 1935 3717 1939 3721
rect 3839 3720 3843 3724
rect 3995 3719 3999 3723
rect 4203 3719 4207 3723
rect 4435 3719 4439 3723
rect 4691 3719 4695 3723
rect 4963 3719 4967 3723
rect 5251 3719 5255 3723
rect 5515 3719 5519 3723
rect 5663 3720 5667 3724
rect 111 3700 115 3704
rect 131 3701 135 3705
rect 307 3701 311 3705
rect 499 3701 503 3705
rect 683 3701 687 3705
rect 859 3701 863 3705
rect 1027 3701 1031 3705
rect 1187 3701 1191 3705
rect 1339 3701 1343 3705
rect 1491 3701 1495 3705
rect 1651 3701 1655 3705
rect 1787 3701 1791 3705
rect 1935 3700 1939 3704
rect 3839 3703 3843 3707
rect 4023 3704 4027 3708
rect 4231 3704 4235 3708
rect 4463 3704 4467 3708
rect 4719 3704 4723 3708
rect 4991 3704 4995 3708
rect 5279 3704 5283 3708
rect 5543 3704 5547 3708
rect 5663 3703 5667 3707
rect 1975 3697 1979 3701
rect 2279 3696 2283 3700
rect 243 3691 247 3695
rect 435 3691 436 3695
rect 436 3691 439 3695
rect 227 3683 231 3687
rect 811 3691 812 3695
rect 812 3691 815 3695
rect 1131 3691 1135 3695
rect 1151 3691 1152 3695
rect 1152 3691 1155 3695
rect 1315 3691 1316 3695
rect 1316 3691 1319 3695
rect 1467 3691 1468 3695
rect 1468 3691 1471 3695
rect 1639 3691 1643 3695
rect 1779 3691 1780 3695
rect 1780 3691 1783 3695
rect 1883 3691 1887 3695
rect 2479 3696 2483 3700
rect 2679 3696 2683 3700
rect 2879 3696 2883 3700
rect 3079 3696 3083 3700
rect 3279 3696 3283 3700
rect 3799 3697 3803 3701
rect 1975 3680 1979 3684
rect 2251 3681 2255 3685
rect 2451 3681 2455 3685
rect 2651 3681 2655 3685
rect 2851 3681 2855 3685
rect 3051 3681 3055 3685
rect 3251 3681 3255 3685
rect 3799 3680 3803 3684
rect 2347 3671 2351 3675
rect 2595 3671 2599 3675
rect 2947 3663 2951 3667
rect 227 3651 231 3655
rect 403 3651 407 3655
rect 435 3651 439 3655
rect 811 3651 815 3655
rect 1123 3651 1127 3655
rect 1131 3651 1135 3655
rect 1315 3651 1319 3655
rect 1467 3651 1471 3655
rect 1639 3651 1643 3655
rect 1779 3651 1783 3655
rect 1415 3643 1419 3647
rect 2391 3631 2395 3635
rect 2947 3631 2951 3635
rect 3103 3631 3107 3635
rect 243 3607 247 3611
rect 1671 3615 1675 3619
rect 3839 3617 3843 3621
rect 4215 3616 4219 3620
rect 4399 3616 4403 3620
rect 4607 3616 4611 3620
rect 4831 3616 4835 3620
rect 5071 3616 5075 3620
rect 5319 3616 5323 3620
rect 5543 3616 5547 3620
rect 5663 3617 5667 3621
rect 363 3603 367 3607
rect 579 3603 583 3607
rect 811 3603 815 3607
rect 1139 3603 1143 3607
rect 1583 3607 1587 3611
rect 1883 3607 1887 3611
rect 3839 3600 3843 3604
rect 4187 3601 4191 3605
rect 4371 3601 4375 3605
rect 4579 3601 4583 3605
rect 4803 3601 4807 3605
rect 5043 3601 5047 3605
rect 5291 3601 5295 3605
rect 5515 3601 5519 3605
rect 5663 3600 5667 3604
rect 1923 3587 1927 3591
rect 2347 3587 2351 3591
rect 2523 3583 2527 3587
rect 2851 3583 2855 3587
rect 2987 3583 2991 3587
rect 4327 3591 4331 3595
rect 4539 3591 4543 3595
rect 4707 3591 4708 3595
rect 4708 3591 4711 3595
rect 4931 3591 4932 3595
rect 4932 3591 4935 3595
rect 3635 3583 3639 3587
rect 4627 3583 4631 3587
rect 5347 3591 5351 3595
rect 5611 3591 5615 3595
rect 363 3563 367 3567
rect 579 3563 583 3567
rect 811 3563 815 3567
rect 927 3563 928 3567
rect 928 3563 931 3567
rect 1123 3563 1127 3567
rect 1415 3563 1416 3567
rect 1416 3563 1419 3567
rect 1671 3563 1672 3567
rect 1672 3563 1675 3567
rect 1923 3563 1927 3567
rect 111 3556 115 3560
rect 147 3555 151 3559
rect 355 3555 359 3559
rect 571 3555 575 3559
rect 803 3555 807 3559
rect 1043 3555 1047 3559
rect 1291 3555 1295 3559
rect 1547 3555 1551 3559
rect 1787 3555 1791 3559
rect 1935 3556 1939 3560
rect 2851 3551 2855 3555
rect 111 3539 115 3543
rect 175 3540 179 3544
rect 383 3540 387 3544
rect 599 3540 603 3544
rect 831 3540 835 3544
rect 1071 3540 1075 3544
rect 1319 3540 1323 3544
rect 1575 3540 1579 3544
rect 1815 3540 1819 3544
rect 1935 3539 1939 3543
rect 2091 3543 2095 3547
rect 2523 3543 2527 3547
rect 2639 3543 2640 3547
rect 2640 3543 2643 3547
rect 2987 3543 2991 3547
rect 3103 3543 3104 3547
rect 3104 3543 3107 3547
rect 4327 3551 4331 3555
rect 4539 3551 4543 3555
rect 4707 3551 4711 3555
rect 4931 3551 4935 3555
rect 5387 3551 5391 3555
rect 5627 3551 5631 3555
rect 4815 3543 4819 3547
rect 1975 3536 1979 3540
rect 1995 3535 1999 3539
rect 2251 3535 2255 3539
rect 2515 3535 2519 3539
rect 2755 3535 2759 3539
rect 2979 3535 2983 3539
rect 3195 3535 3199 3539
rect 3411 3535 3415 3539
rect 3627 3535 3631 3539
rect 3799 3536 3803 3540
rect 1975 3519 1979 3523
rect 2023 3520 2027 3524
rect 2279 3520 2283 3524
rect 2543 3520 2547 3524
rect 2783 3520 2787 3524
rect 3007 3520 3011 3524
rect 3223 3520 3227 3524
rect 3439 3520 3443 3524
rect 3655 3520 3659 3524
rect 3799 3519 3803 3523
rect 4627 3495 4631 3499
rect 4691 3491 4695 3495
rect 4851 3491 4855 3495
rect 5011 3491 5015 3495
rect 5179 3491 5183 3495
rect 5319 3495 5323 3499
rect 5611 3495 5615 3499
rect 111 3457 115 3461
rect 303 3456 307 3460
rect 447 3456 451 3460
rect 599 3456 603 3460
rect 759 3456 763 3460
rect 935 3456 939 3460
rect 1111 3456 1115 3460
rect 1295 3456 1299 3460
rect 1487 3456 1491 3460
rect 1935 3457 1939 3461
rect 1975 3453 1979 3457
rect 2023 3452 2027 3456
rect 2191 3452 2195 3456
rect 2399 3452 2403 3456
rect 2615 3452 2619 3456
rect 2831 3452 2835 3456
rect 3047 3452 3051 3456
rect 3263 3452 3267 3456
rect 3479 3452 3483 3456
rect 3679 3452 3683 3456
rect 3799 3453 3803 3457
rect 4691 3451 4695 3455
rect 4851 3451 4855 3455
rect 5011 3451 5015 3455
rect 5179 3451 5183 3455
rect 5239 3451 5243 3455
rect 5387 3451 5391 3455
rect 5639 3451 5640 3455
rect 5640 3451 5643 3455
rect 111 3440 115 3444
rect 275 3441 279 3445
rect 419 3441 423 3445
rect 571 3441 575 3445
rect 731 3441 735 3445
rect 907 3441 911 3445
rect 1083 3441 1087 3445
rect 1267 3441 1271 3445
rect 1459 3441 1463 3445
rect 1935 3440 1939 3444
rect 3839 3444 3843 3448
rect 4531 3443 4535 3447
rect 4683 3443 4687 3447
rect 4843 3443 4847 3447
rect 5003 3443 5007 3447
rect 5171 3443 5175 3447
rect 5347 3443 5351 3447
rect 5515 3443 5519 3447
rect 5663 3444 5667 3448
rect 1975 3436 1979 3440
rect 1995 3437 1999 3441
rect 2163 3437 2167 3441
rect 2371 3437 2375 3441
rect 2587 3437 2591 3441
rect 2803 3437 2807 3441
rect 3019 3437 3023 3441
rect 3235 3437 3239 3441
rect 3451 3437 3455 3441
rect 3651 3437 3655 3441
rect 3799 3436 3803 3440
rect 403 3431 404 3435
rect 404 3431 407 3435
rect 547 3431 548 3435
rect 548 3431 551 3435
rect 719 3431 723 3435
rect 763 3431 767 3435
rect 1035 3431 1036 3435
rect 1036 3431 1039 3435
rect 1139 3431 1143 3435
rect 1395 3431 1396 3435
rect 1396 3431 1399 3435
rect 1583 3431 1584 3435
rect 1584 3431 1587 3435
rect 2123 3427 2124 3431
rect 2124 3427 2127 3431
rect 2335 3427 2339 3431
rect 2347 3427 2351 3431
rect 3147 3427 3148 3431
rect 3148 3427 3151 3431
rect 3363 3427 3364 3431
rect 3364 3427 3367 3431
rect 3635 3427 3639 3431
rect 3691 3427 3695 3431
rect 3839 3427 3843 3431
rect 4559 3428 4563 3432
rect 4711 3428 4715 3432
rect 4871 3428 4875 3432
rect 5031 3428 5035 3432
rect 5199 3428 5203 3432
rect 5375 3428 5379 3432
rect 5543 3428 5547 3432
rect 5663 3427 5667 3431
rect 403 3391 407 3395
rect 547 3391 551 3395
rect 719 3391 723 3395
rect 835 3391 839 3395
rect 1035 3391 1039 3395
rect 1363 3391 1367 3395
rect 1395 3391 1399 3395
rect 927 3383 931 3387
rect 2091 3387 2095 3391
rect 2123 3387 2127 3391
rect 2335 3387 2339 3391
rect 2639 3387 2643 3391
rect 3147 3387 3151 3391
rect 3363 3387 3367 3391
rect 3747 3387 3751 3391
rect 3691 3371 3695 3375
rect 3839 3365 3843 3369
rect 3887 3364 3891 3368
rect 4151 3364 4155 3368
rect 4423 3364 4427 3368
rect 4671 3364 4675 3368
rect 4895 3364 4899 3368
rect 5111 3364 5115 3368
rect 5327 3364 5331 3368
rect 5543 3364 5547 3368
rect 5663 3365 5667 3369
rect 3839 3348 3843 3352
rect 3859 3349 3863 3353
rect 4123 3349 4127 3353
rect 4395 3349 4399 3353
rect 4643 3349 4647 3353
rect 4867 3349 4871 3353
rect 5083 3349 5087 3353
rect 5299 3349 5303 3353
rect 5515 3349 5519 3353
rect 5663 3348 5667 3352
rect 563 3339 567 3343
rect 763 3343 767 3347
rect 883 3339 887 3343
rect 1099 3339 1103 3343
rect 1391 3343 1395 3347
rect 3747 3339 3751 3343
rect 4131 3339 4135 3343
rect 4523 3339 4524 3343
rect 4524 3339 4527 3343
rect 4771 3339 4772 3343
rect 4772 3339 4775 3343
rect 5255 3339 5259 3343
rect 5143 3331 5147 3335
rect 5611 3339 5615 3343
rect 2187 3315 2191 3319
rect 2347 3315 2351 3319
rect 835 3307 839 3311
rect 2627 3311 2631 3315
rect 2907 3311 2911 3315
rect 3011 3311 3015 3315
rect 3195 3311 3199 3315
rect 3379 3311 3383 3315
rect 3563 3311 3567 3315
rect 883 3299 887 3303
rect 1099 3299 1103 3303
rect 1155 3299 1159 3303
rect 1363 3299 1367 3303
rect 4131 3307 4135 3311
rect 3987 3299 3991 3303
rect 111 3292 115 3296
rect 467 3291 471 3295
rect 667 3291 671 3295
rect 875 3291 879 3295
rect 1091 3291 1095 3295
rect 1315 3291 1319 3295
rect 1935 3292 1939 3296
rect 4523 3299 4527 3303
rect 4771 3299 4775 3303
rect 5255 3299 5259 3303
rect 5639 3299 5643 3303
rect 5239 3291 5243 3295
rect 111 3275 115 3279
rect 495 3276 499 3280
rect 695 3276 699 3280
rect 903 3276 907 3280
rect 1119 3276 1123 3280
rect 1343 3276 1347 3280
rect 1935 3275 1939 3279
rect 1951 3271 1955 3275
rect 2187 3271 2191 3275
rect 2627 3271 2631 3275
rect 2731 3271 2735 3275
rect 3011 3271 3015 3275
rect 3195 3271 3199 3275
rect 3379 3271 3383 3275
rect 3563 3271 3567 3275
rect 3679 3271 3680 3275
rect 3680 3271 3683 3275
rect 1975 3264 1979 3268
rect 1995 3263 1999 3267
rect 2195 3263 2199 3267
rect 2411 3263 2415 3267
rect 2619 3263 2623 3267
rect 2811 3263 2815 3267
rect 3003 3263 3007 3267
rect 3187 3263 3191 3267
rect 3371 3263 3375 3267
rect 3555 3263 3559 3267
rect 3799 3264 3803 3268
rect 3955 3263 3959 3267
rect 4195 3263 4199 3267
rect 4355 3263 4359 3267
rect 4979 3267 4983 3271
rect 5143 3267 5147 3271
rect 5347 3267 5351 3271
rect 5611 3267 5615 3271
rect 1975 3247 1979 3251
rect 2023 3248 2027 3252
rect 2223 3248 2227 3252
rect 2439 3248 2443 3252
rect 2647 3248 2651 3252
rect 2839 3248 2843 3252
rect 3031 3248 3035 3252
rect 3215 3248 3219 3252
rect 3399 3248 3403 3252
rect 3583 3248 3587 3252
rect 3799 3247 3803 3251
rect 4195 3231 4199 3235
rect 3987 3223 3988 3227
rect 3988 3223 3991 3227
rect 4355 3223 4359 3227
rect 4475 3223 4476 3227
rect 4476 3223 4479 3227
rect 4979 3223 4983 3227
rect 5319 3223 5323 3227
rect 5347 3223 5351 3227
rect 111 3217 115 3221
rect 535 3216 539 3220
rect 727 3216 731 3220
rect 919 3216 923 3220
rect 1111 3216 1115 3220
rect 1295 3216 1299 3220
rect 1471 3216 1475 3220
rect 1655 3216 1659 3220
rect 1815 3216 1819 3220
rect 1935 3217 1939 3221
rect 3839 3216 3843 3220
rect 3859 3215 3863 3219
rect 4099 3215 4103 3219
rect 4347 3215 4351 3219
rect 4579 3215 4583 3219
rect 4787 3215 4791 3219
rect 4987 3215 4991 3219
rect 5171 3215 5175 3219
rect 5355 3215 5359 3219
rect 5515 3215 5519 3219
rect 5663 3216 5667 3220
rect 111 3200 115 3204
rect 507 3201 511 3205
rect 699 3201 703 3205
rect 891 3201 895 3205
rect 1083 3201 1087 3205
rect 1267 3201 1271 3205
rect 1443 3201 1447 3205
rect 1627 3201 1631 3205
rect 1787 3201 1791 3205
rect 1935 3200 1939 3204
rect 3839 3199 3843 3203
rect 3887 3200 3891 3204
rect 4127 3200 4131 3204
rect 4375 3200 4379 3204
rect 4607 3200 4611 3204
rect 4815 3200 4819 3204
rect 5015 3200 5019 3204
rect 5199 3200 5203 3204
rect 5383 3200 5387 3204
rect 5543 3200 5547 3204
rect 5663 3199 5667 3203
rect 563 3191 567 3195
rect 659 3191 663 3195
rect 1211 3191 1212 3195
rect 1212 3191 1215 3195
rect 1391 3191 1392 3195
rect 1392 3191 1395 3195
rect 1567 3191 1568 3195
rect 1568 3191 1571 3195
rect 1595 3191 1599 3195
rect 1975 3189 1979 3193
rect 2463 3188 2467 3192
rect 2663 3188 2667 3192
rect 2863 3188 2867 3192
rect 3055 3188 3059 3192
rect 3239 3188 3243 3192
rect 3431 3188 3435 3192
rect 3623 3188 3627 3192
rect 3799 3189 3803 3193
rect 1975 3172 1979 3176
rect 2435 3173 2439 3177
rect 2635 3173 2639 3177
rect 2835 3173 2839 3177
rect 3027 3173 3031 3177
rect 3211 3173 3215 3177
rect 3403 3173 3407 3177
rect 3595 3173 3599 3177
rect 3799 3172 3803 3176
rect 2427 3163 2431 3167
rect 2907 3163 2911 3167
rect 3339 3163 3340 3167
rect 3340 3163 3343 3167
rect 3527 3163 3528 3167
rect 3528 3163 3531 3167
rect 551 3151 555 3155
rect 1155 3143 1159 3147
rect 1211 3151 1215 3155
rect 1595 3151 1599 3155
rect 1951 3151 1955 3155
rect 3307 3155 3311 3159
rect 1399 3143 1403 3147
rect 2731 3123 2735 3127
rect 3123 3123 3127 3127
rect 3307 3123 3311 3127
rect 3339 3123 3343 3127
rect 3679 3123 3683 3127
rect 3839 3125 3843 3129
rect 3903 3124 3907 3128
rect 4135 3124 4139 3128
rect 4359 3124 4363 3128
rect 4583 3124 4587 3128
rect 4807 3124 4811 3128
rect 5031 3124 5035 3128
rect 5663 3125 5667 3129
rect 435 3107 439 3111
rect 659 3111 663 3115
rect 707 3107 711 3111
rect 843 3107 847 3111
rect 979 3107 983 3111
rect 1115 3107 1119 3111
rect 1251 3107 1255 3111
rect 1387 3107 1391 3111
rect 1567 3111 1571 3115
rect 1659 3107 1663 3111
rect 1795 3107 1799 3111
rect 3839 3108 3843 3112
rect 3875 3109 3879 3113
rect 4107 3109 4111 3113
rect 4331 3109 4335 3113
rect 4555 3109 4559 3113
rect 4779 3109 4783 3113
rect 5003 3109 5007 3113
rect 5663 3108 5667 3112
rect 3955 3099 3959 3103
rect 4235 3099 4236 3103
rect 4236 3099 4239 3103
rect 4455 3099 4456 3103
rect 4456 3099 4459 3103
rect 4683 3099 4684 3103
rect 4684 3099 4687 3103
rect 4907 3099 4908 3103
rect 4908 3099 4911 3103
rect 4203 3091 4207 3095
rect 2427 3079 2431 3083
rect 2563 3075 2567 3079
rect 2839 3079 2843 3083
rect 3011 3075 3015 3079
rect 3527 3079 3531 3083
rect 551 3067 552 3071
rect 552 3067 555 3071
rect 707 3067 711 3071
rect 843 3067 847 3071
rect 979 3067 983 3071
rect 1115 3067 1119 3071
rect 1251 3067 1255 3071
rect 1387 3067 1391 3071
rect 1399 3067 1403 3071
rect 1659 3067 1663 3071
rect 1795 3067 1799 3071
rect 1907 3067 1911 3071
rect 111 3060 115 3064
rect 427 3059 431 3063
rect 563 3059 567 3063
rect 699 3059 703 3063
rect 835 3059 839 3063
rect 971 3059 975 3063
rect 1107 3059 1111 3063
rect 1243 3059 1247 3063
rect 1379 3059 1383 3063
rect 1515 3059 1519 3063
rect 1651 3059 1655 3063
rect 1787 3059 1791 3063
rect 1935 3060 1939 3064
rect 3971 3059 3975 3063
rect 4203 3059 4207 3063
rect 4235 3059 4239 3063
rect 4475 3059 4479 3063
rect 4683 3059 4687 3063
rect 4907 3059 4911 3063
rect 111 3043 115 3047
rect 455 3044 459 3048
rect 591 3044 595 3048
rect 727 3044 731 3048
rect 863 3044 867 3048
rect 999 3044 1003 3048
rect 1135 3044 1139 3048
rect 1271 3044 1275 3048
rect 1407 3044 1411 3048
rect 1543 3044 1547 3048
rect 1679 3044 1683 3048
rect 1815 3044 1819 3048
rect 1935 3043 1939 3047
rect 2563 3035 2567 3039
rect 2611 3035 2615 3039
rect 3011 3035 3015 3039
rect 3123 3035 3127 3039
rect 3359 3035 3360 3039
rect 3360 3035 3363 3039
rect 1975 3028 1979 3032
rect 2331 3027 2335 3031
rect 2555 3027 2559 3031
rect 2779 3027 2783 3031
rect 3003 3027 3007 3031
rect 3235 3027 3239 3031
rect 3467 3027 3471 3031
rect 3799 3028 3803 3032
rect 3991 3027 3995 3031
rect 4879 3035 4883 3039
rect 4251 3023 4255 3027
rect 4455 3027 4459 3031
rect 4587 3023 4591 3027
rect 4763 3023 4767 3027
rect 1975 3011 1979 3015
rect 2359 3012 2363 3016
rect 2583 3012 2587 3016
rect 2807 3012 2811 3016
rect 3031 3012 3035 3016
rect 3263 3012 3267 3016
rect 3495 3012 3499 3016
rect 3799 3011 3803 3015
rect 3971 2983 3975 2987
rect 4251 2983 4255 2987
rect 4367 2983 4368 2987
rect 4368 2983 4371 2987
rect 4587 2983 4591 2987
rect 4763 2983 4767 2987
rect 4879 2983 4880 2987
rect 4880 2983 4883 2987
rect 3839 2976 3843 2980
rect 3907 2975 3911 2979
rect 4075 2975 4079 2979
rect 4243 2975 4247 2979
rect 4411 2975 4415 2979
rect 4579 2975 4583 2979
rect 4755 2975 4759 2979
rect 5663 2976 5667 2980
rect 111 2957 115 2961
rect 199 2956 203 2960
rect 511 2956 515 2960
rect 815 2956 819 2960
rect 1111 2956 1115 2960
rect 1415 2956 1419 2960
rect 1719 2956 1723 2960
rect 1935 2957 1939 2961
rect 3839 2959 3843 2963
rect 3935 2960 3939 2964
rect 4103 2960 4107 2964
rect 4271 2960 4275 2964
rect 4439 2960 4443 2964
rect 4607 2960 4611 2964
rect 4783 2960 4787 2964
rect 5663 2959 5667 2963
rect 111 2940 115 2944
rect 171 2941 175 2945
rect 483 2941 487 2945
rect 787 2941 791 2945
rect 1083 2941 1087 2945
rect 1387 2941 1391 2945
rect 1691 2941 1695 2945
rect 1935 2940 1939 2944
rect 1975 2941 1979 2945
rect 2143 2940 2147 2944
rect 2343 2940 2347 2944
rect 2543 2940 2547 2944
rect 2743 2940 2747 2944
rect 2935 2940 2939 2944
rect 3135 2940 3139 2944
rect 3335 2940 3339 2944
rect 3799 2941 3803 2945
rect 435 2931 439 2935
rect 443 2931 447 2935
rect 723 2931 727 2935
rect 1211 2931 1212 2935
rect 1212 2931 1215 2935
rect 1671 2931 1675 2935
rect 1975 2924 1979 2928
rect 2115 2925 2119 2929
rect 2315 2925 2319 2929
rect 2515 2925 2519 2929
rect 2715 2925 2719 2929
rect 2907 2925 2911 2929
rect 3107 2925 3111 2929
rect 3307 2925 3311 2929
rect 3799 2924 3803 2928
rect 2251 2915 2255 2919
rect 2275 2915 2279 2919
rect 2475 2915 2479 2919
rect 2839 2915 2840 2919
rect 2840 2915 2843 2919
rect 3031 2915 3032 2919
rect 3032 2915 3035 2919
rect 3067 2915 3071 2919
rect 3267 2915 3271 2919
rect 3839 2897 3843 2901
rect 3895 2896 3899 2900
rect 443 2891 447 2895
rect 723 2891 727 2895
rect 1027 2891 1031 2895
rect 1671 2891 1675 2895
rect 4031 2896 4035 2900
rect 4167 2896 4171 2900
rect 4303 2896 4307 2900
rect 4439 2896 4443 2900
rect 4575 2896 4579 2900
rect 5663 2897 5667 2901
rect 1907 2891 1911 2895
rect 3839 2880 3843 2884
rect 3867 2881 3871 2885
rect 4003 2881 4007 2885
rect 4139 2881 4143 2885
rect 4275 2881 4279 2885
rect 4411 2881 4415 2885
rect 4547 2881 4551 2885
rect 5663 2880 5667 2884
rect 2275 2875 2279 2879
rect 2475 2875 2479 2879
rect 2611 2875 2615 2879
rect 2635 2875 2639 2879
rect 3067 2875 3071 2879
rect 3267 2875 3271 2879
rect 3359 2875 3363 2879
rect 3991 2871 3992 2875
rect 3992 2871 3995 2875
rect 4123 2871 4127 2875
rect 4403 2871 4404 2875
rect 4404 2871 4407 2875
rect 4539 2871 4540 2875
rect 4540 2871 4543 2875
rect 299 2859 303 2863
rect 315 2855 319 2859
rect 531 2855 535 2859
rect 771 2855 775 2859
rect 1019 2855 1023 2859
rect 1211 2859 1215 2863
rect 4235 2863 4239 2867
rect 1547 2855 1551 2859
rect 2155 2835 2159 2839
rect 2251 2835 2255 2839
rect 2515 2831 2519 2835
rect 3031 2835 3035 2839
rect 3963 2831 3967 2835
rect 4235 2831 4239 2835
rect 4367 2831 4371 2835
rect 4403 2831 4407 2835
rect 4539 2831 4543 2835
rect 315 2815 319 2819
rect 531 2815 535 2819
rect 771 2815 775 2819
rect 1019 2815 1023 2819
rect 1027 2815 1031 2819
rect 1547 2815 1551 2819
rect 1619 2815 1623 2819
rect 111 2808 115 2812
rect 131 2807 135 2811
rect 307 2807 311 2811
rect 523 2807 527 2811
rect 763 2807 767 2811
rect 1011 2807 1015 2811
rect 1275 2807 1279 2811
rect 1539 2807 1543 2811
rect 1935 2808 1939 2812
rect 111 2791 115 2795
rect 159 2792 163 2796
rect 335 2792 339 2796
rect 551 2792 555 2796
rect 791 2792 795 2796
rect 1039 2792 1043 2796
rect 1303 2792 1307 2796
rect 1567 2792 1571 2796
rect 1935 2791 1939 2795
rect 2091 2791 2095 2795
rect 2155 2791 2159 2795
rect 2635 2791 2636 2795
rect 2636 2791 2639 2795
rect 2807 2791 2811 2795
rect 4055 2791 4059 2795
rect 4123 2791 4127 2795
rect 1975 2784 1979 2788
rect 2011 2783 2015 2787
rect 2259 2783 2263 2787
rect 2507 2783 2511 2787
rect 2755 2783 2759 2787
rect 3003 2783 3007 2787
rect 3799 2784 3803 2788
rect 4275 2787 4279 2791
rect 4411 2787 4415 2791
rect 4547 2787 4551 2791
rect 4683 2787 4687 2791
rect 4819 2787 4823 2791
rect 1975 2767 1979 2771
rect 2039 2768 2043 2772
rect 2287 2768 2291 2772
rect 2535 2768 2539 2772
rect 2783 2768 2787 2772
rect 3031 2768 3035 2772
rect 3799 2767 3803 2771
rect 3963 2747 3967 2751
rect 4275 2747 4279 2751
rect 4411 2747 4415 2751
rect 4547 2747 4551 2751
rect 4683 2747 4687 2751
rect 4819 2747 4823 2751
rect 4831 2747 4835 2751
rect 3839 2740 3843 2744
rect 3859 2739 3863 2743
rect 3995 2739 3999 2743
rect 4131 2739 4135 2743
rect 4267 2739 4271 2743
rect 4403 2739 4407 2743
rect 4539 2739 4543 2743
rect 4675 2739 4679 2743
rect 4811 2739 4815 2743
rect 5663 2740 5667 2744
rect 111 2729 115 2733
rect 279 2728 283 2732
rect 455 2728 459 2732
rect 647 2728 651 2732
rect 855 2728 859 2732
rect 1079 2728 1083 2732
rect 1311 2728 1315 2732
rect 1551 2728 1555 2732
rect 1799 2728 1803 2732
rect 1935 2729 1939 2733
rect 3839 2723 3843 2727
rect 3887 2724 3891 2728
rect 4023 2724 4027 2728
rect 4159 2724 4163 2728
rect 4295 2724 4299 2728
rect 4431 2724 4435 2728
rect 4567 2724 4571 2728
rect 4703 2724 4707 2728
rect 4839 2724 4843 2728
rect 5663 2723 5667 2727
rect 111 2712 115 2716
rect 251 2713 255 2717
rect 427 2713 431 2717
rect 619 2713 623 2717
rect 827 2713 831 2717
rect 1051 2713 1055 2717
rect 1283 2713 1287 2717
rect 1523 2713 1527 2717
rect 1771 2713 1775 2717
rect 1935 2712 1939 2716
rect 299 2703 303 2707
rect 407 2703 411 2707
rect 1407 2703 1408 2707
rect 1408 2703 1411 2707
rect 1787 2703 1791 2707
rect 1975 2705 1979 2709
rect 2023 2704 2027 2708
rect 2247 2704 2251 2708
rect 2503 2704 2507 2708
rect 2759 2704 2763 2708
rect 3015 2704 3019 2708
rect 3799 2705 3803 2709
rect 1975 2688 1979 2692
rect 1995 2689 1999 2693
rect 2219 2689 2223 2693
rect 2475 2689 2479 2693
rect 2731 2689 2735 2693
rect 2987 2689 2991 2693
rect 3799 2688 3803 2692
rect 407 2663 411 2667
rect 1019 2663 1023 2667
rect 1619 2663 1623 2667
rect 2515 2679 2519 2683
rect 2603 2679 2604 2683
rect 2604 2679 2607 2683
rect 2859 2679 2860 2683
rect 2860 2679 2863 2683
rect 3111 2679 3112 2683
rect 3112 2679 3115 2683
rect 3839 2665 3843 2669
rect 3959 2664 3963 2668
rect 4255 2664 4259 2668
rect 4543 2664 4547 2668
rect 4823 2664 4827 2668
rect 5111 2664 5115 2668
rect 5399 2664 5403 2668
rect 5663 2665 5667 2669
rect 3839 2648 3843 2652
rect 3931 2649 3935 2653
rect 4227 2649 4231 2653
rect 4515 2649 4519 2653
rect 4795 2649 4799 2653
rect 5083 2649 5087 2653
rect 5371 2649 5375 2653
rect 5663 2648 5667 2652
rect 883 2635 887 2639
rect 2091 2639 2095 2643
rect 739 2627 743 2631
rect 899 2627 903 2631
rect 1187 2631 1191 2635
rect 1407 2631 1411 2635
rect 1787 2631 1791 2635
rect 2539 2631 2543 2635
rect 2603 2639 2607 2643
rect 2859 2639 2863 2643
rect 4055 2639 4056 2643
rect 4056 2639 4059 2643
rect 4443 2639 4447 2643
rect 4639 2639 4640 2643
rect 4640 2639 4643 2643
rect 4975 2639 4979 2643
rect 5267 2639 5271 2643
rect 5419 2639 5423 2643
rect 2807 2631 2811 2635
rect 4323 2623 4327 2627
rect 4831 2623 4835 2627
rect 2775 2595 2779 2599
rect 3111 2595 3115 2599
rect 3983 2599 3987 2603
rect 4323 2599 4327 2603
rect 4443 2599 4447 2603
rect 4891 2599 4895 2603
rect 4975 2599 4979 2603
rect 5267 2599 5271 2603
rect 739 2587 743 2591
rect 899 2587 903 2591
rect 1019 2587 1020 2591
rect 1020 2587 1023 2591
rect 1091 2587 1095 2591
rect 1187 2587 1191 2591
rect 1499 2587 1503 2591
rect 111 2580 115 2584
rect 571 2579 575 2583
rect 731 2579 735 2583
rect 891 2579 895 2583
rect 1043 2579 1047 2583
rect 1195 2579 1199 2583
rect 1355 2579 1359 2583
rect 1515 2579 1519 2583
rect 1675 2579 1679 2583
rect 1935 2580 1939 2584
rect 111 2563 115 2567
rect 599 2564 603 2568
rect 759 2564 763 2568
rect 919 2564 923 2568
rect 1071 2564 1075 2568
rect 1223 2564 1227 2568
rect 1383 2564 1387 2568
rect 1543 2564 1547 2568
rect 1703 2564 1707 2568
rect 1935 2563 1939 2567
rect 4179 2563 4183 2567
rect 4639 2567 4643 2571
rect 5171 2563 5175 2567
rect 5419 2567 5423 2571
rect 2539 2551 2543 2555
rect 2951 2551 2952 2555
rect 2952 2551 2955 2555
rect 1975 2544 1979 2548
rect 2555 2543 2559 2547
rect 2691 2543 2695 2547
rect 2827 2543 2831 2547
rect 2963 2543 2967 2547
rect 3099 2543 3103 2547
rect 3799 2544 3803 2548
rect 1975 2527 1979 2531
rect 2583 2528 2587 2532
rect 2719 2528 2723 2532
rect 2855 2528 2859 2532
rect 2991 2528 2995 2532
rect 3127 2528 3131 2532
rect 3799 2527 3803 2531
rect 3983 2523 3984 2527
rect 3984 2523 3987 2527
rect 4395 2523 4399 2527
rect 4891 2523 4895 2527
rect 5447 2523 5448 2527
rect 5448 2523 5451 2527
rect 3839 2516 3843 2520
rect 3859 2515 3863 2519
rect 4083 2515 4087 2519
rect 4331 2515 4335 2519
rect 4579 2515 4583 2519
rect 4827 2515 4831 2519
rect 5075 2515 5079 2519
rect 5323 2515 5327 2519
rect 5663 2516 5667 2520
rect 111 2505 115 2509
rect 383 2504 387 2508
rect 599 2504 603 2508
rect 815 2504 819 2508
rect 1023 2504 1027 2508
rect 1231 2504 1235 2508
rect 1431 2504 1435 2508
rect 1631 2504 1635 2508
rect 1815 2504 1819 2508
rect 1935 2505 1939 2509
rect 3839 2499 3843 2503
rect 3887 2500 3891 2504
rect 4111 2500 4115 2504
rect 4359 2500 4363 2504
rect 4607 2500 4611 2504
rect 4855 2500 4859 2504
rect 5103 2500 5107 2504
rect 5351 2500 5355 2504
rect 5663 2499 5667 2503
rect 111 2488 115 2492
rect 355 2489 359 2493
rect 571 2489 575 2493
rect 787 2489 791 2493
rect 995 2489 999 2493
rect 1203 2489 1207 2493
rect 1403 2489 1407 2493
rect 1603 2489 1607 2493
rect 1787 2489 1791 2493
rect 1935 2488 1939 2492
rect 883 2479 887 2483
rect 1167 2479 1171 2483
rect 1563 2479 1567 2483
rect 1731 2479 1732 2483
rect 1732 2479 1735 2483
rect 1883 2479 1887 2483
rect 1975 2445 1979 2449
rect 2023 2444 2027 2448
rect 363 2439 367 2443
rect 1091 2439 1095 2443
rect 1167 2439 1171 2443
rect 1499 2439 1503 2443
rect 1563 2439 1567 2443
rect 2223 2444 2227 2448
rect 2447 2444 2451 2448
rect 2679 2444 2683 2448
rect 2927 2444 2931 2448
rect 3183 2444 3187 2448
rect 3439 2444 3443 2448
rect 3679 2444 3683 2448
rect 3799 2445 3803 2449
rect 1731 2439 1735 2443
rect 3839 2437 3843 2441
rect 3887 2436 3891 2440
rect 4087 2436 4091 2440
rect 4327 2436 4331 2440
rect 4583 2436 4587 2440
rect 4847 2436 4851 2440
rect 5119 2436 5123 2440
rect 5399 2436 5403 2440
rect 5663 2437 5667 2441
rect 1975 2428 1979 2432
rect 1995 2429 1999 2433
rect 2195 2429 2199 2433
rect 2419 2429 2423 2433
rect 2651 2429 2655 2433
rect 2899 2429 2903 2433
rect 3155 2429 3159 2433
rect 3411 2429 3415 2433
rect 3651 2429 3655 2433
rect 3799 2428 3803 2432
rect 2091 2419 2095 2423
rect 2323 2419 2324 2423
rect 2324 2419 2327 2423
rect 2547 2419 2548 2423
rect 2548 2419 2551 2423
rect 2775 2419 2776 2423
rect 2776 2419 2779 2423
rect 3027 2419 3028 2423
rect 3028 2419 3031 2423
rect 3283 2419 3284 2423
rect 3284 2419 3287 2423
rect 3535 2419 3536 2423
rect 3536 2419 3539 2423
rect 3823 2419 3827 2423
rect 3839 2420 3843 2424
rect 3859 2421 3863 2425
rect 4059 2421 4063 2425
rect 4299 2421 4303 2425
rect 4555 2421 4559 2425
rect 4819 2421 4823 2425
rect 5091 2421 5095 2425
rect 5371 2421 5375 2425
rect 5663 2420 5667 2424
rect 455 2403 459 2407
rect 1279 2411 1283 2415
rect 1595 2411 1599 2415
rect 4023 2411 4027 2415
rect 4179 2411 4183 2415
rect 4683 2411 4684 2415
rect 4684 2411 4687 2415
rect 4891 2411 4895 2415
rect 5171 2411 5175 2415
rect 5435 2411 5439 2415
rect 619 2399 623 2403
rect 1883 2403 1887 2407
rect 2323 2379 2327 2383
rect 2547 2379 2551 2383
rect 2951 2379 2955 2383
rect 3027 2379 3031 2383
rect 3283 2379 3287 2383
rect 3747 2379 3751 2383
rect 363 2359 367 2363
rect 455 2359 459 2363
rect 899 2359 903 2363
rect 1279 2359 1280 2363
rect 1280 2359 1283 2363
rect 1595 2359 1599 2363
rect 2547 2371 2551 2375
rect 3823 2371 3827 2375
rect 4023 2371 4027 2375
rect 4395 2371 4399 2375
rect 4683 2371 4687 2375
rect 5099 2371 5103 2375
rect 5447 2371 5451 2375
rect 111 2352 115 2356
rect 227 2351 231 2355
rect 523 2351 527 2355
rect 835 2351 839 2355
rect 1155 2351 1159 2355
rect 1483 2351 1487 2355
rect 1787 2351 1791 2355
rect 1935 2352 1939 2356
rect 111 2335 115 2339
rect 255 2336 259 2340
rect 551 2336 555 2340
rect 863 2336 867 2340
rect 1183 2336 1187 2340
rect 1511 2336 1515 2340
rect 1815 2336 1819 2340
rect 1935 2335 1939 2339
rect 2091 2339 2095 2343
rect 2163 2335 2167 2339
rect 2355 2335 2359 2339
rect 2807 2339 2811 2343
rect 3019 2335 3023 2339
rect 3123 2335 3127 2339
rect 3395 2335 3399 2339
rect 3535 2339 3539 2343
rect 3659 2335 3663 2339
rect 4891 2331 4895 2335
rect 4619 2323 4623 2327
rect 4795 2323 4799 2327
rect 5327 2327 5331 2331
rect 5435 2327 5439 2331
rect 5523 2323 5527 2327
rect 3019 2303 3023 2307
rect 2163 2295 2167 2299
rect 2355 2295 2359 2299
rect 2471 2295 2472 2299
rect 2472 2295 2475 2299
rect 2547 2295 2551 2299
rect 3123 2295 3127 2299
rect 3239 2295 3240 2299
rect 3240 2295 3243 2299
rect 3659 2295 3663 2299
rect 3747 2295 3751 2299
rect 1975 2288 1979 2292
rect 1995 2287 1999 2291
rect 2155 2287 2159 2291
rect 2347 2287 2351 2291
rect 2539 2287 2543 2291
rect 2731 2287 2735 2291
rect 2923 2287 2927 2291
rect 3115 2287 3119 2291
rect 3299 2287 3303 2291
rect 3483 2287 3487 2291
rect 3651 2287 3655 2291
rect 3799 2288 3803 2292
rect 4619 2283 4623 2287
rect 4795 2283 4799 2287
rect 4903 2283 4907 2287
rect 5099 2283 5103 2287
rect 5523 2283 5527 2287
rect 5611 2283 5615 2287
rect 1975 2271 1979 2275
rect 2023 2272 2027 2276
rect 2183 2272 2187 2276
rect 2375 2272 2379 2276
rect 2567 2272 2571 2276
rect 2759 2272 2763 2276
rect 2951 2272 2955 2276
rect 3143 2272 3147 2276
rect 3327 2272 3331 2276
rect 3511 2272 3515 2276
rect 3839 2276 3843 2280
rect 3679 2272 3683 2276
rect 4443 2275 4447 2279
rect 3799 2271 3803 2275
rect 4611 2275 4615 2279
rect 4787 2275 4791 2279
rect 4963 2275 4967 2279
rect 5147 2275 5151 2279
rect 5339 2275 5343 2279
rect 5515 2275 5519 2279
rect 5663 2276 5667 2280
rect 111 2261 115 2265
rect 159 2260 163 2264
rect 367 2260 371 2264
rect 599 2260 603 2264
rect 831 2260 835 2264
rect 1063 2260 1067 2264
rect 1935 2261 1939 2265
rect 3839 2259 3843 2263
rect 4471 2260 4475 2264
rect 4639 2260 4643 2264
rect 4815 2260 4819 2264
rect 4991 2260 4995 2264
rect 5175 2260 5179 2264
rect 5367 2260 5371 2264
rect 5543 2260 5547 2264
rect 5663 2259 5667 2263
rect 111 2244 115 2248
rect 131 2245 135 2249
rect 339 2245 343 2249
rect 571 2245 575 2249
rect 803 2245 807 2249
rect 1035 2245 1039 2249
rect 1935 2244 1939 2248
rect 279 2235 283 2239
rect 467 2235 468 2239
rect 468 2235 471 2239
rect 619 2235 623 2239
rect 931 2235 932 2239
rect 932 2235 935 2239
rect 1159 2235 1160 2239
rect 1160 2235 1163 2239
rect 1975 2205 1979 2209
rect 2023 2204 2027 2208
rect 2191 2204 2195 2208
rect 2359 2204 2363 2208
rect 2535 2204 2539 2208
rect 2711 2204 2715 2208
rect 2879 2204 2883 2208
rect 3047 2204 3051 2208
rect 3207 2204 3211 2208
rect 3367 2204 3371 2208
rect 3535 2204 3539 2208
rect 3679 2204 3683 2208
rect 3799 2205 3803 2209
rect 227 2195 231 2199
rect 279 2195 283 2199
rect 467 2195 471 2199
rect 899 2195 903 2199
rect 931 2195 935 2199
rect 1975 2188 1979 2192
rect 1995 2189 1999 2193
rect 2163 2189 2167 2193
rect 2331 2189 2335 2193
rect 2507 2189 2511 2193
rect 2683 2189 2687 2193
rect 2851 2189 2855 2193
rect 3019 2189 3023 2193
rect 3179 2189 3183 2193
rect 3339 2189 3343 2193
rect 3507 2189 3511 2193
rect 3651 2189 3655 2193
rect 3799 2188 3803 2192
rect 3839 2189 3843 2193
rect 4543 2188 4547 2192
rect 4719 2188 4723 2192
rect 4911 2188 4915 2192
rect 5119 2188 5123 2192
rect 5335 2188 5339 2192
rect 5543 2188 5547 2192
rect 5663 2189 5667 2193
rect 2123 2179 2124 2183
rect 2124 2179 2127 2183
rect 2291 2179 2292 2183
rect 2292 2179 2295 2183
rect 2459 2179 2460 2183
rect 2460 2179 2463 2183
rect 2635 2179 2636 2183
rect 2636 2179 2639 2183
rect 2807 2179 2808 2183
rect 2808 2179 2811 2183
rect 2979 2179 2980 2183
rect 2980 2179 2983 2183
rect 3143 2179 3144 2183
rect 3144 2179 3147 2183
rect 2947 2171 2951 2175
rect 3395 2179 3399 2183
rect 3479 2179 3483 2183
rect 3839 2172 3843 2176
rect 4515 2173 4519 2177
rect 4691 2173 4695 2177
rect 4883 2173 4887 2177
rect 5091 2173 5095 2177
rect 5307 2173 5311 2177
rect 5515 2173 5519 2177
rect 5663 2172 5667 2176
rect 4643 2163 4644 2167
rect 4644 2163 4647 2167
rect 4671 2163 4675 2167
rect 5279 2163 5283 2167
rect 5327 2163 5331 2167
rect 5639 2163 5640 2167
rect 5640 2163 5643 2167
rect 339 2151 343 2155
rect 639 2151 643 2155
rect 1159 2151 1163 2155
rect 1795 2147 1799 2151
rect 2123 2139 2127 2143
rect 2291 2139 2295 2143
rect 2459 2139 2463 2143
rect 2635 2139 2639 2143
rect 2947 2139 2951 2143
rect 2979 2139 2983 2143
rect 3239 2139 3243 2143
rect 3479 2139 3483 2143
rect 3747 2139 3751 2143
rect 2471 2131 2475 2135
rect 4671 2123 4675 2127
rect 4903 2123 4907 2127
rect 5167 2123 5171 2127
rect 5279 2123 5283 2127
rect 5611 2123 5615 2127
rect 227 2107 231 2111
rect 339 2107 343 2111
rect 959 2107 960 2111
rect 960 2107 963 2111
rect 1439 2107 1440 2111
rect 1440 2107 1443 2111
rect 111 2100 115 2104
rect 131 2099 135 2103
rect 347 2099 351 2103
rect 595 2099 599 2103
rect 835 2099 839 2103
rect 1075 2099 1079 2103
rect 1315 2099 1319 2103
rect 1563 2099 1567 2103
rect 1787 2099 1791 2103
rect 1935 2100 1939 2104
rect 3143 2091 3147 2095
rect 3767 2095 3771 2099
rect 111 2083 115 2087
rect 159 2084 163 2088
rect 375 2084 379 2088
rect 623 2084 627 2088
rect 863 2084 867 2088
rect 1103 2084 1107 2088
rect 1343 2084 1347 2088
rect 1591 2084 1595 2088
rect 1815 2084 1819 2088
rect 1935 2083 1939 2087
rect 3251 2087 3255 2091
rect 3387 2087 3391 2091
rect 3659 2087 3663 2091
rect 4643 2091 4647 2095
rect 4779 2087 4783 2091
rect 4915 2087 4919 2091
rect 5051 2087 5055 2091
rect 5367 2091 5371 2095
rect 3251 2047 3255 2051
rect 3387 2047 3391 2051
rect 3467 2047 3471 2051
rect 3659 2047 3663 2051
rect 3747 2047 3751 2051
rect 4779 2047 4783 2051
rect 4915 2047 4919 2051
rect 5051 2047 5055 2051
rect 5167 2047 5168 2051
rect 5168 2047 5171 2051
rect 5219 2047 5223 2051
rect 1975 2040 1979 2044
rect 3107 2039 3111 2043
rect 3243 2039 3247 2043
rect 3379 2039 3383 2043
rect 3515 2039 3519 2043
rect 3651 2039 3655 2043
rect 3799 2040 3803 2044
rect 3839 2040 3843 2044
rect 4635 2039 4639 2043
rect 4771 2039 4775 2043
rect 4907 2039 4911 2043
rect 5043 2039 5047 2043
rect 5179 2039 5183 2043
rect 5663 2040 5667 2044
rect 111 2021 115 2025
rect 271 2020 275 2024
rect 407 2020 411 2024
rect 543 2020 547 2024
rect 687 2020 691 2024
rect 831 2020 835 2024
rect 975 2020 979 2024
rect 1119 2020 1123 2024
rect 1263 2020 1267 2024
rect 1407 2020 1411 2024
rect 1543 2020 1547 2024
rect 1679 2020 1683 2024
rect 1815 2020 1819 2024
rect 1935 2021 1939 2025
rect 1975 2023 1979 2027
rect 3135 2024 3139 2028
rect 3271 2024 3275 2028
rect 3407 2024 3411 2028
rect 3543 2024 3547 2028
rect 3679 2024 3683 2028
rect 3799 2023 3803 2027
rect 3839 2023 3843 2027
rect 4663 2024 4667 2028
rect 4799 2024 4803 2028
rect 4935 2024 4939 2028
rect 5071 2024 5075 2028
rect 5207 2024 5211 2028
rect 5663 2023 5667 2027
rect 111 2004 115 2008
rect 243 2005 247 2009
rect 379 2005 383 2009
rect 515 2005 519 2009
rect 659 2005 663 2009
rect 803 2005 807 2009
rect 947 2005 951 2009
rect 1091 2005 1095 2009
rect 1235 2005 1239 2009
rect 1379 2005 1383 2009
rect 1515 2005 1519 2009
rect 1651 2005 1655 2009
rect 1787 2005 1791 2009
rect 1935 2004 1939 2008
rect 371 1995 372 1999
rect 372 1995 375 1999
rect 507 1995 508 1999
rect 508 1995 511 1999
rect 639 1995 640 1999
rect 640 1995 643 1999
rect 683 1995 687 1999
rect 1219 1995 1220 1999
rect 1220 1995 1223 1999
rect 1359 1995 1360 1999
rect 1360 1995 1363 1999
rect 1507 1995 1508 1999
rect 1508 1995 1511 1999
rect 1187 1987 1191 1991
rect 1795 1995 1799 1999
rect 1747 1987 1751 1991
rect 1975 1965 1979 1969
rect 3127 1964 3131 1968
rect 3263 1964 3267 1968
rect 3399 1964 3403 1968
rect 3535 1964 3539 1968
rect 3671 1964 3675 1968
rect 3799 1965 3803 1969
rect 3839 1965 3843 1969
rect 4863 1964 4867 1968
rect 4999 1964 5003 1968
rect 5135 1964 5139 1968
rect 5271 1964 5275 1968
rect 5407 1964 5411 1968
rect 5543 1964 5547 1968
rect 5663 1965 5667 1969
rect 311 1955 315 1959
rect 371 1955 375 1959
rect 507 1955 511 1959
rect 959 1955 963 1959
rect 1187 1955 1191 1959
rect 1219 1955 1223 1959
rect 1439 1955 1443 1959
rect 1507 1955 1511 1959
rect 1747 1955 1751 1959
rect 1883 1955 1887 1959
rect 1975 1948 1979 1952
rect 3099 1949 3103 1953
rect 3235 1949 3239 1953
rect 3371 1949 3375 1953
rect 3507 1949 3511 1953
rect 3643 1949 3647 1953
rect 3799 1948 3803 1952
rect 3839 1948 3843 1952
rect 4835 1949 4839 1953
rect 4971 1949 4975 1953
rect 5107 1949 5111 1953
rect 5243 1949 5247 1953
rect 5379 1949 5383 1953
rect 5515 1949 5519 1953
rect 5663 1948 5667 1952
rect 3203 1939 3207 1943
rect 3635 1939 3636 1943
rect 3636 1939 3639 1943
rect 3767 1939 3768 1943
rect 3768 1939 3771 1943
rect 4771 1939 4775 1943
rect 5367 1939 5368 1943
rect 5368 1939 5371 1943
rect 5387 1939 5391 1943
rect 5611 1939 5615 1943
rect 475 1915 479 1919
rect 683 1919 687 1923
rect 819 1915 823 1919
rect 1059 1915 1063 1919
rect 1359 1919 1363 1923
rect 1563 1915 1567 1919
rect 2119 1919 2123 1923
rect 3467 1899 3471 1903
rect 3603 1899 3607 1903
rect 3635 1899 3639 1903
rect 5219 1899 5223 1903
rect 5387 1907 5391 1911
rect 5639 1899 5643 1903
rect 311 1875 312 1879
rect 312 1875 315 1879
rect 819 1875 823 1879
rect 1059 1875 1063 1879
rect 1135 1875 1139 1879
rect 1563 1875 1567 1879
rect 1643 1875 1647 1879
rect 1883 1875 1887 1879
rect 111 1868 115 1872
rect 187 1867 191 1871
rect 379 1867 383 1871
rect 587 1867 591 1871
rect 811 1867 815 1871
rect 1051 1867 1055 1871
rect 1299 1867 1303 1871
rect 1555 1867 1559 1871
rect 1787 1867 1791 1871
rect 1935 1868 1939 1872
rect 111 1851 115 1855
rect 215 1852 219 1856
rect 407 1852 411 1856
rect 615 1852 619 1856
rect 839 1852 843 1856
rect 1079 1852 1083 1856
rect 1327 1852 1331 1856
rect 1583 1852 1587 1856
rect 1815 1852 1819 1856
rect 1935 1851 1939 1855
rect 2219 1855 2223 1859
rect 2403 1855 2407 1859
rect 2411 1855 2415 1859
rect 2787 1851 2791 1855
rect 2915 1851 2919 1855
rect 3203 1855 3207 1859
rect 3395 1851 3399 1855
rect 3491 1851 3495 1855
rect 3983 1855 3987 1859
rect 4771 1855 4775 1859
rect 4827 1851 4831 1855
rect 4971 1851 4975 1855
rect 5251 1851 5255 1855
rect 5611 1855 5615 1859
rect 2787 1819 2791 1823
rect 2119 1811 2120 1815
rect 2120 1811 2123 1815
rect 2219 1811 2223 1815
rect 2403 1811 2407 1815
rect 2915 1811 2919 1815
rect 3031 1811 3032 1815
rect 3032 1811 3035 1815
rect 3395 1819 3399 1823
rect 3491 1811 3495 1815
rect 3603 1811 3607 1815
rect 4827 1811 4831 1815
rect 4971 1811 4975 1815
rect 5087 1811 5088 1815
rect 5088 1811 5091 1815
rect 5251 1811 5255 1815
rect 5499 1811 5503 1815
rect 1975 1804 1979 1808
rect 1995 1803 1999 1807
rect 2227 1803 2231 1807
rect 2467 1803 2471 1807
rect 2691 1803 2695 1807
rect 2907 1803 2911 1807
rect 3107 1803 3111 1807
rect 3299 1803 3303 1807
rect 3483 1803 3487 1807
rect 3651 1803 3655 1807
rect 3799 1804 3803 1808
rect 3839 1804 3843 1808
rect 4675 1803 4679 1807
rect 4819 1803 4823 1807
rect 4963 1803 4967 1807
rect 5107 1803 5111 1807
rect 5243 1803 5247 1807
rect 5379 1803 5383 1807
rect 5515 1803 5519 1807
rect 5663 1804 5667 1808
rect 111 1785 115 1789
rect 159 1784 163 1788
rect 375 1784 379 1788
rect 591 1784 595 1788
rect 799 1784 803 1788
rect 999 1784 1003 1788
rect 1191 1784 1195 1788
rect 1383 1784 1387 1788
rect 1575 1784 1579 1788
rect 1935 1785 1939 1789
rect 1975 1787 1979 1791
rect 2023 1788 2027 1792
rect 2255 1788 2259 1792
rect 2495 1788 2499 1792
rect 2719 1788 2723 1792
rect 2935 1788 2939 1792
rect 3135 1788 3139 1792
rect 3327 1788 3331 1792
rect 3511 1788 3515 1792
rect 3679 1788 3683 1792
rect 3799 1787 3803 1791
rect 3839 1787 3843 1791
rect 4703 1788 4707 1792
rect 4847 1788 4851 1792
rect 4991 1788 4995 1792
rect 5135 1788 5139 1792
rect 5271 1788 5275 1792
rect 5407 1788 5411 1792
rect 5543 1788 5547 1792
rect 5663 1787 5667 1791
rect 111 1768 115 1772
rect 131 1769 135 1773
rect 347 1769 351 1773
rect 563 1769 567 1773
rect 771 1769 775 1773
rect 971 1769 975 1773
rect 1163 1769 1167 1773
rect 1355 1769 1359 1773
rect 1547 1769 1551 1773
rect 1935 1768 1939 1772
rect 291 1759 295 1763
rect 475 1759 476 1763
rect 476 1759 479 1763
rect 491 1759 495 1763
rect 1107 1759 1111 1763
rect 1287 1759 1288 1763
rect 1288 1759 1291 1763
rect 1067 1751 1071 1755
rect 227 1719 231 1723
rect 291 1719 295 1723
rect 1067 1719 1071 1723
rect 1107 1719 1111 1723
rect 1643 1719 1647 1723
rect 1975 1721 1979 1725
rect 2023 1720 2027 1724
rect 2159 1720 2163 1724
rect 2311 1720 2315 1724
rect 2471 1720 2475 1724
rect 2639 1720 2643 1724
rect 2807 1720 2811 1724
rect 2975 1720 2979 1724
rect 3151 1720 3155 1724
rect 3799 1721 3803 1725
rect 1135 1711 1139 1715
rect 3839 1713 3843 1717
rect 3887 1712 3891 1716
rect 4079 1712 4083 1716
rect 4303 1712 4307 1716
rect 4535 1712 4539 1716
rect 4775 1712 4779 1716
rect 5023 1712 5027 1716
rect 5279 1712 5283 1716
rect 5535 1712 5539 1716
rect 5663 1713 5667 1717
rect 1975 1704 1979 1708
rect 1995 1705 1999 1709
rect 2131 1705 2135 1709
rect 2283 1705 2287 1709
rect 2443 1705 2447 1709
rect 2611 1705 2615 1709
rect 2779 1705 2783 1709
rect 2947 1705 2951 1709
rect 3123 1705 3127 1709
rect 3799 1704 3803 1708
rect 2123 1695 2124 1699
rect 2124 1695 2127 1699
rect 2259 1695 2260 1699
rect 2260 1695 2263 1699
rect 2411 1695 2412 1699
rect 2412 1695 2415 1699
rect 2091 1687 2095 1691
rect 2603 1695 2607 1699
rect 2915 1695 2919 1699
rect 3075 1695 3076 1699
rect 3076 1695 3079 1699
rect 2875 1687 2879 1691
rect 3839 1696 3843 1700
rect 3859 1697 3863 1701
rect 4051 1697 4055 1701
rect 4275 1697 4279 1701
rect 4507 1697 4511 1701
rect 4747 1697 4751 1701
rect 4995 1697 4999 1701
rect 5251 1697 5255 1701
rect 5507 1697 5511 1701
rect 5663 1696 5667 1700
rect 3983 1687 3984 1691
rect 3984 1687 3987 1691
rect 4435 1687 4439 1691
rect 4635 1687 4636 1691
rect 4636 1687 4639 1691
rect 4871 1687 4872 1691
rect 4872 1687 4875 1691
rect 4371 1679 4375 1683
rect 5555 1687 5559 1691
rect 239 1663 243 1667
rect 491 1663 495 1667
rect 691 1659 695 1663
rect 1075 1659 1079 1663
rect 1287 1663 1291 1667
rect 2091 1655 2095 1659
rect 2123 1655 2127 1659
rect 2259 1655 2263 1659
rect 2603 1655 2607 1659
rect 2707 1655 2711 1659
rect 2875 1655 2879 1659
rect 3031 1655 3035 1659
rect 3075 1655 3079 1659
rect 4147 1647 4151 1651
rect 4371 1647 4375 1651
rect 4435 1647 4439 1651
rect 4635 1647 4639 1651
rect 5087 1647 5091 1651
rect 5347 1647 5351 1651
rect 5499 1647 5503 1651
rect 1075 1631 1079 1635
rect 227 1619 231 1623
rect 691 1619 695 1623
rect 987 1619 991 1623
rect 995 1619 999 1623
rect 111 1612 115 1616
rect 131 1611 135 1615
rect 395 1611 399 1615
rect 683 1611 687 1615
rect 979 1611 983 1615
rect 1275 1611 1279 1615
rect 1935 1612 1939 1616
rect 2187 1611 2191 1615
rect 2235 1611 2239 1615
rect 2371 1611 2375 1615
rect 2507 1611 2511 1615
rect 2643 1611 2647 1615
rect 2779 1611 2783 1615
rect 2915 1615 2919 1619
rect 3051 1611 3055 1615
rect 3187 1611 3191 1615
rect 3955 1611 3959 1615
rect 4003 1611 4007 1615
rect 4251 1611 4255 1615
rect 4399 1615 4403 1619
rect 4683 1611 4687 1615
rect 4871 1615 4875 1619
rect 5139 1611 5143 1615
rect 5467 1615 5471 1619
rect 111 1595 115 1599
rect 159 1596 163 1600
rect 423 1596 427 1600
rect 711 1596 715 1600
rect 1007 1596 1011 1600
rect 1303 1596 1307 1600
rect 1935 1595 1939 1599
rect 2707 1579 2711 1583
rect 2235 1571 2239 1575
rect 2371 1571 2375 1575
rect 2507 1571 2511 1575
rect 2643 1571 2647 1575
rect 2779 1571 2783 1575
rect 3955 1579 3959 1583
rect 3051 1571 3055 1575
rect 3187 1571 3191 1575
rect 3299 1571 3303 1575
rect 4003 1571 4007 1575
rect 4123 1571 4124 1575
rect 4124 1571 4127 1575
rect 4147 1571 4151 1575
rect 4479 1571 4480 1575
rect 4480 1571 4483 1575
rect 4683 1579 4687 1583
rect 5139 1571 5143 1575
rect 5347 1571 5351 1575
rect 1975 1564 1979 1568
rect 2091 1563 2095 1567
rect 2227 1563 2231 1567
rect 2363 1563 2367 1567
rect 2499 1563 2503 1567
rect 2635 1563 2639 1567
rect 2771 1563 2775 1567
rect 2907 1563 2911 1567
rect 3043 1563 3047 1567
rect 3179 1563 3183 1567
rect 3799 1564 3803 1568
rect 3839 1564 3843 1568
rect 3859 1563 3863 1567
rect 3995 1563 3999 1567
rect 4155 1563 4159 1567
rect 4355 1563 4359 1567
rect 4587 1563 4591 1567
rect 4851 1563 4855 1567
rect 5131 1563 5135 1567
rect 5419 1563 5423 1567
rect 5663 1564 5667 1568
rect 1975 1547 1979 1551
rect 2119 1548 2123 1552
rect 2255 1548 2259 1552
rect 2391 1548 2395 1552
rect 2527 1548 2531 1552
rect 2663 1548 2667 1552
rect 2799 1548 2803 1552
rect 2935 1548 2939 1552
rect 3071 1548 3075 1552
rect 3207 1548 3211 1552
rect 3799 1547 3803 1551
rect 3839 1547 3843 1551
rect 3887 1548 3891 1552
rect 4023 1548 4027 1552
rect 4183 1548 4187 1552
rect 4383 1548 4387 1552
rect 4615 1548 4619 1552
rect 4879 1548 4883 1552
rect 5159 1548 5163 1552
rect 5447 1548 5451 1552
rect 5663 1547 5667 1551
rect 111 1525 115 1529
rect 159 1524 163 1528
rect 375 1524 379 1528
rect 607 1524 611 1528
rect 839 1524 843 1528
rect 1071 1524 1075 1528
rect 1303 1524 1307 1528
rect 1935 1525 1939 1529
rect 111 1508 115 1512
rect 131 1509 135 1513
rect 347 1509 351 1513
rect 579 1509 583 1513
rect 811 1509 815 1513
rect 1043 1509 1047 1513
rect 1275 1509 1279 1513
rect 1935 1508 1939 1512
rect 2187 1507 2191 1511
rect 2655 1507 2659 1511
rect 239 1499 243 1503
rect 355 1499 359 1503
rect 719 1499 723 1503
rect 803 1499 807 1503
rect 1171 1499 1172 1503
rect 1172 1499 1175 1503
rect 1403 1499 1404 1503
rect 1404 1499 1407 1503
rect 4123 1503 4127 1507
rect 4259 1503 4263 1507
rect 3839 1489 3843 1493
rect 3887 1488 3891 1492
rect 4023 1488 4027 1492
rect 4159 1488 4163 1492
rect 4303 1488 4307 1492
rect 4495 1488 4499 1492
rect 4719 1488 4723 1492
rect 4967 1488 4971 1492
rect 5223 1488 5227 1492
rect 5487 1488 5491 1492
rect 5663 1489 5667 1493
rect 355 1467 359 1471
rect 803 1459 807 1463
rect 995 1467 999 1471
rect 1975 1469 1979 1473
rect 2023 1468 2027 1472
rect 2159 1468 2163 1472
rect 2295 1468 2299 1472
rect 2431 1468 2435 1472
rect 2567 1468 2571 1472
rect 2703 1468 2707 1472
rect 2839 1468 2843 1472
rect 2975 1468 2979 1472
rect 3799 1469 3803 1473
rect 3839 1472 3843 1476
rect 3859 1473 3863 1477
rect 3995 1473 3999 1477
rect 4131 1473 4135 1477
rect 4275 1473 4279 1477
rect 4467 1473 4471 1477
rect 4691 1473 4695 1477
rect 4939 1473 4943 1477
rect 5195 1473 5199 1477
rect 5459 1473 5463 1477
rect 5663 1472 5667 1476
rect 987 1459 991 1463
rect 1171 1459 1175 1463
rect 3987 1463 3988 1467
rect 3988 1463 3991 1467
rect 4123 1463 4124 1467
rect 4124 1463 4127 1467
rect 4251 1463 4255 1467
rect 4399 1463 4400 1467
rect 4400 1463 4403 1467
rect 4595 1463 4596 1467
rect 4596 1463 4599 1467
rect 4819 1463 4820 1467
rect 4820 1463 4823 1467
rect 5067 1463 5068 1467
rect 5068 1463 5071 1467
rect 1975 1452 1979 1456
rect 1995 1453 1999 1457
rect 2131 1453 2135 1457
rect 2267 1453 2271 1457
rect 2403 1453 2407 1457
rect 2539 1453 2543 1457
rect 2675 1453 2679 1457
rect 2811 1453 2815 1457
rect 2947 1453 2951 1457
rect 3799 1452 3803 1456
rect 4155 1455 4159 1459
rect 5583 1463 5584 1467
rect 5584 1463 5587 1467
rect 2123 1443 2124 1447
rect 2124 1443 2127 1447
rect 2259 1443 2260 1447
rect 2260 1443 2263 1447
rect 2395 1443 2396 1447
rect 2396 1443 2399 1447
rect 2531 1443 2532 1447
rect 2532 1443 2535 1447
rect 2655 1443 2659 1447
rect 2803 1443 2804 1447
rect 2804 1443 2807 1447
rect 2935 1443 2936 1447
rect 2936 1443 2939 1447
rect 2771 1435 2775 1439
rect 3955 1423 3959 1427
rect 3987 1423 3991 1427
rect 4123 1423 4127 1427
rect 4259 1423 4263 1427
rect 4479 1423 4483 1427
rect 4595 1423 4599 1427
rect 4819 1423 4823 1427
rect 5067 1423 5071 1427
rect 5555 1423 5559 1427
rect 227 1411 231 1415
rect 507 1411 511 1415
rect 719 1415 723 1419
rect 1187 1411 1191 1415
rect 1403 1415 1407 1419
rect 1883 1411 1887 1415
rect 2123 1403 2127 1407
rect 2259 1403 2263 1407
rect 2395 1403 2399 1407
rect 2531 1403 2535 1407
rect 2771 1403 2775 1407
rect 2803 1403 2807 1407
rect 3299 1403 3303 1407
rect 507 1391 511 1395
rect 863 1391 867 1395
rect 1187 1391 1191 1395
rect 1575 1391 1579 1395
rect 2299 1395 2303 1399
rect 3779 1387 3783 1391
rect 4155 1387 4159 1391
rect 4315 1383 4319 1387
rect 4587 1383 4591 1387
rect 4883 1383 4887 1387
rect 5195 1383 5199 1387
rect 5583 1387 5587 1391
rect 863 1371 864 1375
rect 864 1371 867 1375
rect 1035 1371 1039 1375
rect 1575 1371 1576 1375
rect 1576 1371 1579 1375
rect 111 1364 115 1368
rect 131 1363 135 1367
rect 411 1363 415 1367
rect 739 1363 743 1367
rect 1091 1363 1095 1367
rect 1451 1363 1455 1367
rect 1787 1363 1791 1367
rect 1935 1364 1939 1368
rect 2283 1359 2287 1363
rect 2935 1363 2939 1367
rect 3371 1363 3375 1367
rect 3403 1359 3407 1363
rect 3659 1359 3663 1363
rect 111 1347 115 1351
rect 159 1348 163 1352
rect 439 1348 443 1352
rect 767 1348 771 1352
rect 1119 1348 1123 1352
rect 1479 1348 1483 1352
rect 1815 1348 1819 1352
rect 1935 1347 1939 1351
rect 4683 1351 4687 1355
rect 3955 1343 3959 1347
rect 4315 1343 4319 1347
rect 4587 1343 4591 1347
rect 4883 1343 4887 1347
rect 5195 1343 5199 1347
rect 5611 1343 5615 1347
rect 3839 1336 3843 1340
rect 3859 1335 3863 1339
rect 4059 1335 4063 1339
rect 4307 1335 4311 1339
rect 4579 1335 4583 1339
rect 4875 1335 4879 1339
rect 5187 1335 5191 1339
rect 5499 1335 5503 1339
rect 5663 1336 5667 1340
rect 2283 1319 2287 1323
rect 2299 1319 2303 1323
rect 2687 1319 2688 1323
rect 2688 1319 2691 1323
rect 3403 1319 3407 1323
rect 3659 1319 3663 1323
rect 3779 1319 3780 1323
rect 3780 1319 3783 1323
rect 3839 1319 3843 1323
rect 3887 1320 3891 1324
rect 4087 1320 4091 1324
rect 4335 1320 4339 1324
rect 4607 1320 4611 1324
rect 4903 1320 4907 1324
rect 5215 1320 5219 1324
rect 5527 1320 5531 1324
rect 5663 1319 5667 1323
rect 1975 1312 1979 1316
rect 1995 1311 1999 1315
rect 2275 1311 2279 1315
rect 2563 1311 2567 1315
rect 2843 1311 2847 1315
rect 3123 1311 3127 1315
rect 3395 1311 3399 1315
rect 3651 1311 3655 1315
rect 3799 1312 3803 1316
rect 1975 1295 1979 1299
rect 2023 1296 2027 1300
rect 2303 1296 2307 1300
rect 2591 1296 2595 1300
rect 2871 1296 2875 1300
rect 3151 1296 3155 1300
rect 3423 1296 3427 1300
rect 3679 1296 3683 1300
rect 3799 1295 3803 1299
rect 111 1289 115 1293
rect 159 1288 163 1292
rect 359 1288 363 1292
rect 575 1288 579 1292
rect 775 1288 779 1292
rect 967 1288 971 1292
rect 1151 1288 1155 1292
rect 1327 1288 1331 1292
rect 1495 1288 1499 1292
rect 1663 1288 1667 1292
rect 1815 1288 1819 1292
rect 1935 1289 1939 1293
rect 111 1272 115 1276
rect 131 1273 135 1277
rect 331 1273 335 1277
rect 547 1273 551 1277
rect 747 1273 751 1277
rect 939 1273 943 1277
rect 1123 1273 1127 1277
rect 1299 1273 1303 1277
rect 1467 1273 1471 1277
rect 1635 1273 1639 1277
rect 1787 1273 1791 1277
rect 1935 1272 1939 1276
rect 227 1263 231 1267
rect 387 1263 391 1267
rect 871 1263 872 1267
rect 872 1263 875 1267
rect 1251 1263 1252 1267
rect 1252 1263 1255 1267
rect 1427 1263 1428 1267
rect 1428 1263 1431 1267
rect 1595 1263 1596 1267
rect 1596 1263 1599 1267
rect 1763 1263 1764 1267
rect 1764 1263 1767 1267
rect 1883 1263 1887 1267
rect 3839 1253 3843 1257
rect 4615 1252 4619 1256
rect 4791 1252 4795 1256
rect 4975 1252 4979 1256
rect 5167 1252 5171 1256
rect 5367 1252 5371 1256
rect 5543 1252 5547 1256
rect 5663 1253 5667 1257
rect 3839 1236 3843 1240
rect 4587 1237 4591 1241
rect 4763 1237 4767 1241
rect 4947 1237 4951 1241
rect 5139 1237 5143 1241
rect 5339 1237 5343 1241
rect 5515 1237 5519 1241
rect 5663 1236 5667 1240
rect 227 1223 231 1227
rect 1035 1223 1039 1227
rect 1219 1223 1223 1227
rect 1251 1223 1255 1227
rect 1427 1223 1431 1227
rect 1595 1223 1599 1227
rect 1763 1223 1767 1227
rect 4715 1227 4716 1231
rect 4716 1227 4719 1231
rect 4891 1227 4892 1231
rect 4892 1227 4895 1231
rect 5075 1227 5076 1231
rect 5076 1227 5079 1231
rect 5083 1227 5087 1231
rect 5467 1227 5468 1231
rect 5468 1227 5471 1231
rect 5619 1227 5623 1231
rect 1975 1213 1979 1217
rect 2655 1212 2659 1216
rect 2831 1212 2835 1216
rect 3007 1212 3011 1216
rect 3183 1212 3187 1216
rect 3359 1212 3363 1216
rect 3543 1212 3547 1216
rect 3799 1213 3803 1217
rect 1975 1196 1979 1200
rect 2627 1197 2631 1201
rect 2803 1197 2807 1201
rect 2979 1197 2983 1201
rect 3155 1197 3159 1201
rect 3331 1197 3335 1201
rect 3515 1197 3519 1201
rect 3799 1196 3803 1200
rect 2755 1187 2756 1191
rect 2756 1187 2759 1191
rect 271 1179 275 1183
rect 387 1179 391 1183
rect 483 1175 487 1179
rect 667 1175 671 1179
rect 871 1179 875 1183
rect 1011 1175 1015 1179
rect 1483 1179 1487 1183
rect 1747 1175 1751 1179
rect 2119 1179 2123 1183
rect 2267 1179 2271 1183
rect 3283 1187 3284 1191
rect 3284 1187 3287 1191
rect 3459 1187 3460 1191
rect 3460 1187 3463 1191
rect 3371 1179 3375 1183
rect 4683 1187 4687 1191
rect 4715 1187 4719 1191
rect 4891 1187 4895 1191
rect 5075 1187 5079 1191
rect 5479 1187 5483 1191
rect 5611 1187 5615 1191
rect 5083 1155 5087 1159
rect 1747 1143 1751 1147
rect 2687 1147 2691 1151
rect 2755 1147 2759 1151
rect 227 1135 231 1139
rect 483 1135 487 1139
rect 667 1135 671 1139
rect 755 1135 759 1139
rect 1011 1135 1015 1139
rect 1143 1135 1147 1139
rect 1219 1135 1223 1139
rect 1483 1135 1487 1139
rect 3283 1147 3287 1151
rect 3459 1147 3463 1151
rect 4979 1147 4983 1151
rect 5115 1147 5119 1151
rect 5251 1147 5255 1151
rect 5387 1147 5391 1151
rect 5619 1151 5623 1155
rect 3235 1139 3239 1143
rect 111 1128 115 1132
rect 131 1127 135 1131
rect 291 1127 295 1131
rect 475 1127 479 1131
rect 659 1127 663 1131
rect 835 1127 839 1131
rect 1003 1127 1007 1131
rect 1171 1127 1175 1131
rect 1331 1127 1335 1131
rect 1491 1127 1495 1131
rect 1651 1127 1655 1131
rect 1787 1127 1791 1131
rect 1935 1128 1939 1132
rect 111 1111 115 1115
rect 159 1112 163 1116
rect 319 1112 323 1116
rect 503 1112 507 1116
rect 687 1112 691 1116
rect 863 1112 867 1116
rect 1031 1112 1035 1116
rect 1199 1112 1203 1116
rect 1359 1112 1363 1116
rect 1519 1112 1523 1116
rect 1679 1112 1683 1116
rect 1815 1112 1819 1116
rect 1935 1111 1939 1115
rect 4979 1107 4983 1111
rect 5115 1107 5119 1111
rect 5251 1107 5255 1111
rect 5387 1107 5391 1111
rect 5419 1107 5423 1111
rect 5611 1107 5615 1111
rect 2091 1095 2095 1099
rect 2267 1099 2271 1103
rect 2371 1095 2375 1099
rect 2643 1095 2647 1099
rect 2731 1095 2735 1099
rect 2899 1095 2903 1099
rect 3067 1095 3071 1099
rect 3227 1095 3231 1099
rect 3407 1099 3411 1103
rect 3839 1100 3843 1104
rect 4835 1099 4839 1103
rect 4971 1099 4975 1103
rect 5107 1099 5111 1103
rect 5243 1099 5247 1103
rect 5379 1099 5383 1103
rect 5515 1099 5519 1103
rect 5663 1100 5667 1104
rect 3839 1083 3843 1087
rect 4863 1084 4867 1088
rect 4999 1084 5003 1088
rect 5135 1084 5139 1088
rect 5271 1084 5275 1088
rect 5407 1084 5411 1088
rect 5543 1084 5547 1088
rect 5663 1083 5667 1087
rect 2643 1063 2647 1067
rect 2119 1055 2120 1059
rect 2120 1055 2123 1059
rect 2371 1055 2375 1059
rect 2491 1055 2492 1059
rect 2492 1055 2495 1059
rect 2731 1055 2735 1059
rect 2899 1055 2903 1059
rect 3067 1055 3071 1059
rect 3227 1055 3231 1059
rect 3235 1055 3239 1059
rect 1975 1048 1979 1052
rect 1995 1047 1999 1051
rect 2171 1047 2175 1051
rect 2363 1047 2367 1051
rect 2547 1047 2551 1051
rect 2723 1047 2727 1051
rect 2891 1047 2895 1051
rect 3059 1047 3063 1051
rect 3219 1047 3223 1051
rect 3387 1047 3391 1051
rect 3799 1048 3803 1052
rect 111 1041 115 1045
rect 175 1040 179 1044
rect 431 1040 435 1044
rect 687 1040 691 1044
rect 951 1040 955 1044
rect 1215 1040 1219 1044
rect 1935 1041 1939 1045
rect 1975 1031 1979 1035
rect 2023 1032 2027 1036
rect 2199 1032 2203 1036
rect 2391 1032 2395 1036
rect 2575 1032 2579 1036
rect 2751 1032 2755 1036
rect 2919 1032 2923 1036
rect 3087 1032 3091 1036
rect 3247 1032 3251 1036
rect 3415 1032 3419 1036
rect 3799 1031 3803 1035
rect 111 1024 115 1028
rect 147 1025 151 1029
rect 403 1025 407 1029
rect 659 1025 663 1029
rect 923 1025 927 1029
rect 1187 1025 1191 1029
rect 1935 1024 1939 1028
rect 3839 1021 3843 1025
rect 4807 1020 4811 1024
rect 271 1015 272 1019
rect 272 1015 275 1019
rect 355 1015 359 1019
rect 779 1015 783 1019
rect 1003 1015 1007 1019
rect 1135 1015 1139 1019
rect 4943 1020 4947 1024
rect 5079 1020 5083 1024
rect 5215 1020 5219 1024
rect 5351 1020 5355 1024
rect 5487 1020 5491 1024
rect 5663 1021 5667 1025
rect 3839 1004 3843 1008
rect 4779 1005 4783 1009
rect 4915 1005 4919 1009
rect 5051 1005 5055 1009
rect 5187 1005 5191 1009
rect 5323 1005 5327 1009
rect 5459 1005 5463 1009
rect 5663 1004 5667 1008
rect 4907 995 4908 999
rect 4908 995 4911 999
rect 5043 995 5044 999
rect 5044 995 5047 999
rect 5179 995 5180 999
rect 5180 995 5183 999
rect 4875 987 4879 991
rect 5331 995 5335 999
rect 5479 995 5483 999
rect 355 975 359 979
rect 363 975 367 979
rect 755 975 759 979
rect 1135 975 1139 979
rect 1143 975 1147 979
rect 1975 973 1979 977
rect 2023 972 2027 976
rect 2191 972 2195 976
rect 2375 972 2379 976
rect 2567 972 2571 976
rect 2759 972 2763 976
rect 2943 972 2947 976
rect 3127 972 3131 976
rect 3311 972 3315 976
rect 3495 972 3499 976
rect 3679 972 3683 976
rect 3799 973 3803 977
rect 1975 956 1979 960
rect 1995 957 1999 961
rect 2163 957 2167 961
rect 2347 957 2351 961
rect 2539 957 2543 961
rect 2731 957 2735 961
rect 2915 957 2919 961
rect 3099 957 3103 961
rect 3283 957 3287 961
rect 3467 957 3471 961
rect 3651 957 3655 961
rect 3799 956 3803 960
rect 4875 955 4879 959
rect 4907 955 4911 959
rect 5043 955 5047 959
rect 5331 963 5335 967
rect 5419 955 5423 959
rect 5555 955 5559 959
rect 2091 947 2095 951
rect 2155 947 2159 951
rect 2667 947 2668 951
rect 2668 947 2671 951
rect 2895 947 2899 951
rect 3043 947 3044 951
rect 3044 947 3047 951
rect 3227 947 3228 951
rect 3228 947 3231 951
rect 3407 947 3408 951
rect 3408 947 3411 951
rect 3011 939 3015 943
rect 3643 947 3647 951
rect 271 931 275 935
rect 779 931 783 935
rect 1003 931 1007 935
rect 1139 927 1143 931
rect 1371 927 1375 931
rect 3955 915 3959 919
rect 4163 919 4167 923
rect 4275 919 4279 923
rect 4483 915 4487 919
rect 4651 915 4655 919
rect 4939 915 4943 919
rect 5179 919 5183 923
rect 5611 919 5615 923
rect 2155 907 2159 911
rect 2491 907 2495 911
rect 2667 907 2671 911
rect 3011 907 3015 911
rect 3043 907 3047 911
rect 3227 907 3231 911
rect 3643 907 3647 911
rect 3747 907 3751 911
rect 363 887 364 891
rect 364 887 367 891
rect 499 887 503 891
rect 1139 887 1143 891
rect 1371 887 1375 891
rect 1491 887 1492 891
rect 1492 887 1495 891
rect 111 880 115 884
rect 235 879 239 883
rect 459 879 463 883
rect 683 879 687 883
rect 907 879 911 883
rect 1131 879 1135 883
rect 1363 879 1367 883
rect 1935 880 1939 884
rect 2527 879 2531 883
rect 4483 883 4487 887
rect 111 863 115 867
rect 263 864 267 868
rect 487 864 491 868
rect 711 864 715 868
rect 935 864 939 868
rect 1159 864 1163 868
rect 1391 864 1395 868
rect 1935 863 1939 867
rect 2187 867 2191 871
rect 2771 867 2775 871
rect 2895 871 2899 875
rect 4091 875 4095 879
rect 4163 875 4167 879
rect 4651 875 4655 879
rect 4939 875 4943 879
rect 5067 875 5071 879
rect 5611 875 5615 879
rect 3331 867 3335 871
rect 3839 868 3843 872
rect 3859 867 3863 871
rect 3995 867 3999 871
rect 4171 867 4175 871
rect 4387 867 4391 871
rect 4643 867 4647 871
rect 4931 867 4935 871
rect 5235 867 5239 871
rect 5515 867 5519 871
rect 5663 868 5667 872
rect 3839 851 3843 855
rect 3887 852 3891 856
rect 4023 852 4027 856
rect 4199 852 4203 856
rect 4415 852 4419 856
rect 4671 852 4675 856
rect 4959 852 4963 856
rect 5263 852 5267 856
rect 5543 852 5547 856
rect 5663 851 5667 855
rect 2771 835 2775 839
rect 2187 827 2191 831
rect 2527 827 2528 831
rect 2528 827 2531 831
rect 3331 827 3335 831
rect 3747 827 3751 831
rect 1975 820 1979 824
rect 1995 819 1999 823
rect 2179 819 2183 823
rect 2403 819 2407 823
rect 2675 819 2679 823
rect 2987 819 2991 823
rect 3323 819 3327 823
rect 3651 819 3655 823
rect 3799 820 3803 824
rect 1975 803 1979 807
rect 2023 804 2027 808
rect 2207 804 2211 808
rect 2431 804 2435 808
rect 2703 804 2707 808
rect 3015 804 3019 808
rect 3351 804 3355 808
rect 3679 804 3683 808
rect 3799 803 3803 807
rect 111 789 115 793
rect 175 788 179 792
rect 431 788 435 792
rect 671 788 675 792
rect 903 788 907 792
rect 1127 788 1131 792
rect 1351 788 1355 792
rect 1575 788 1579 792
rect 1935 789 1939 793
rect 3839 793 3843 797
rect 3887 792 3891 796
rect 4023 792 4027 796
rect 4159 792 4163 796
rect 4295 792 4299 796
rect 4431 792 4435 796
rect 4567 792 4571 796
rect 4719 792 4723 796
rect 4895 792 4899 796
rect 5087 792 5091 796
rect 5287 792 5291 796
rect 5487 792 5491 796
rect 5663 793 5667 797
rect 111 772 115 776
rect 147 773 151 777
rect 403 773 407 777
rect 643 773 647 777
rect 875 773 879 777
rect 1099 773 1103 777
rect 1323 773 1327 777
rect 1547 773 1551 777
rect 1935 772 1939 776
rect 3839 776 3843 780
rect 3859 777 3863 781
rect 3995 777 3999 781
rect 4131 777 4135 781
rect 4267 777 4271 781
rect 4403 777 4407 781
rect 4539 777 4543 781
rect 4691 777 4695 781
rect 4867 777 4871 781
rect 5059 777 5063 781
rect 5259 777 5263 781
rect 5459 777 5463 781
rect 5663 776 5667 780
rect 271 763 272 767
rect 272 763 275 767
rect 531 763 532 767
rect 532 763 535 767
rect 767 763 768 767
rect 768 763 771 767
rect 1063 763 1067 767
rect 1483 763 1487 767
rect 3955 767 3959 771
rect 4123 767 4124 771
rect 4124 767 4127 771
rect 4259 767 4260 771
rect 4260 767 4263 771
rect 4395 767 4396 771
rect 4396 767 4399 771
rect 4531 767 4532 771
rect 4532 767 4535 771
rect 4635 767 4639 771
rect 4275 759 4279 763
rect 4843 767 4847 771
rect 5219 767 5223 771
rect 4963 759 4967 763
rect 5555 767 5559 771
rect 243 723 247 727
rect 499 723 503 727
rect 531 723 535 727
rect 1063 723 1067 727
rect 1483 723 1487 727
rect 1491 723 1495 727
rect 3955 727 3959 731
rect 4091 727 4095 731
rect 4123 727 4127 731
rect 4259 727 4263 731
rect 4395 727 4399 731
rect 4531 727 4535 731
rect 4843 727 4847 731
rect 4963 727 4967 731
rect 5067 727 5071 731
rect 5219 727 5223 731
rect 5555 727 5559 731
rect 307 691 311 695
rect 411 687 415 691
rect 619 687 623 691
rect 767 691 771 695
rect 915 687 919 691
rect 1267 687 1271 691
rect 1435 687 1439 691
rect 1603 687 1607 691
rect 1779 687 1783 691
rect 4003 687 4007 691
rect 4139 687 4143 691
rect 4275 687 4279 691
rect 4411 687 4415 691
rect 4635 691 4639 695
rect 4707 687 4711 691
rect 4899 687 4903 691
rect 5107 687 5111 691
rect 5323 687 5327 691
rect 5611 691 5615 695
rect 619 655 623 659
rect 243 647 247 651
rect 307 647 311 651
rect 647 647 648 651
rect 648 647 651 651
rect 915 647 919 651
rect 1267 647 1271 651
rect 1435 647 1439 651
rect 1603 647 1607 651
rect 1779 647 1783 651
rect 1895 647 1896 651
rect 1896 647 1899 651
rect 3955 647 3959 651
rect 4139 647 4143 651
rect 4275 647 4279 651
rect 4411 647 4415 651
rect 4707 647 4711 651
rect 4899 647 4903 651
rect 5107 647 5111 651
rect 5323 647 5327 651
rect 5367 647 5371 651
rect 5555 647 5559 651
rect 111 640 115 644
rect 131 639 135 643
rect 315 639 319 643
rect 523 639 527 643
rect 723 639 727 643
rect 907 639 911 643
rect 1083 639 1087 643
rect 1259 639 1263 643
rect 1427 639 1431 643
rect 1595 639 1599 643
rect 1771 639 1775 643
rect 1935 640 1939 644
rect 3839 640 3843 644
rect 3859 639 3863 643
rect 3995 639 3999 643
rect 4131 639 4135 643
rect 4267 639 4271 643
rect 4403 639 4407 643
rect 4539 639 4543 643
rect 4699 639 4703 643
rect 4891 639 4895 643
rect 5099 639 5103 643
rect 5315 639 5319 643
rect 5515 639 5519 643
rect 5663 640 5667 644
rect 111 623 115 627
rect 159 624 163 628
rect 343 624 347 628
rect 551 624 555 628
rect 751 624 755 628
rect 935 624 939 628
rect 1111 624 1115 628
rect 1287 624 1291 628
rect 1455 624 1459 628
rect 1623 624 1627 628
rect 1799 624 1803 628
rect 1935 623 1939 627
rect 3839 623 3843 627
rect 3887 624 3891 628
rect 4023 624 4027 628
rect 4159 624 4163 628
rect 4295 624 4299 628
rect 4431 624 4435 628
rect 4567 624 4571 628
rect 4727 624 4731 628
rect 4919 624 4923 628
rect 5127 624 5131 628
rect 5343 624 5347 628
rect 5543 624 5547 628
rect 5663 623 5667 627
rect 111 565 115 569
rect 159 564 163 568
rect 375 564 379 568
rect 599 564 603 568
rect 807 564 811 568
rect 999 564 1003 568
rect 1175 564 1179 568
rect 1343 564 1347 568
rect 1511 564 1515 568
rect 1671 564 1675 568
rect 1815 564 1819 568
rect 1935 565 1939 569
rect 3839 565 3843 569
rect 3887 564 3891 568
rect 4071 564 4075 568
rect 4311 564 4315 568
rect 4575 564 4579 568
rect 4855 564 4859 568
rect 5151 564 5155 568
rect 5447 564 5451 568
rect 5663 565 5667 569
rect 111 548 115 552
rect 131 549 135 553
rect 347 549 351 553
rect 571 549 575 553
rect 779 549 783 553
rect 971 549 975 553
rect 1147 549 1151 553
rect 1315 549 1319 553
rect 1483 549 1487 553
rect 1643 549 1647 553
rect 1787 549 1791 553
rect 1935 548 1939 552
rect 1975 545 1979 549
rect 3135 544 3139 548
rect 255 539 256 543
rect 256 539 259 543
rect 411 539 415 543
rect 743 539 747 543
rect 907 539 908 543
rect 908 539 911 543
rect 1275 539 1276 543
rect 1276 539 1279 543
rect 1443 539 1444 543
rect 1444 539 1447 543
rect 1631 539 1635 543
rect 1771 539 1772 543
rect 1772 539 1775 543
rect 1883 539 1887 543
rect 3271 544 3275 548
rect 3407 544 3411 548
rect 3543 544 3547 548
rect 3679 544 3683 548
rect 3799 545 3803 549
rect 3839 548 3843 552
rect 3859 549 3863 553
rect 4043 549 4047 553
rect 4283 549 4287 553
rect 4547 549 4551 553
rect 4827 549 4831 553
rect 5123 549 5127 553
rect 5419 549 5423 553
rect 5663 548 5667 552
rect 4003 539 4007 543
rect 4171 539 4172 543
rect 4172 539 4175 543
rect 4675 539 4676 543
rect 4676 539 4679 543
rect 1975 528 1979 532
rect 3107 529 3111 533
rect 3243 529 3247 533
rect 3379 529 3383 533
rect 3515 529 3519 533
rect 3651 529 3655 533
rect 3799 528 3803 532
rect 4635 531 4639 535
rect 5543 539 5544 543
rect 5544 539 5547 543
rect 3235 519 3236 523
rect 3236 519 3239 523
rect 3371 519 3372 523
rect 3372 519 3375 523
rect 3507 519 3508 523
rect 3508 519 3511 523
rect 3643 519 3644 523
rect 3644 519 3647 523
rect 3779 519 3780 523
rect 3780 519 3783 523
rect 227 499 231 503
rect 255 499 259 503
rect 647 499 651 503
rect 743 499 747 503
rect 907 499 911 503
rect 1275 499 1279 503
rect 1443 499 1447 503
rect 1631 499 1635 503
rect 1771 499 1775 503
rect 3779 499 3783 503
rect 1895 491 1899 495
rect 4171 499 4175 503
rect 4675 499 4679 503
rect 5395 499 5399 503
rect 3203 479 3207 483
rect 3235 479 3239 483
rect 3371 479 3375 483
rect 3507 479 3511 483
rect 3643 479 3647 483
rect 5367 483 5371 487
rect 251 463 255 467
rect 579 463 583 467
rect 907 463 911 467
rect 1483 463 1487 467
rect 1883 467 1887 471
rect 4635 455 4639 459
rect 1915 447 1919 451
rect 2211 443 2215 447
rect 2435 443 2439 447
rect 2659 443 2663 447
rect 2955 443 2959 447
rect 3075 443 3079 447
rect 3275 443 3279 447
rect 3475 443 3479 447
rect 3635 447 3639 451
rect 4651 451 4655 455
rect 4851 451 4855 455
rect 5059 451 5063 455
rect 5363 451 5367 455
rect 5543 455 5547 459
rect 251 431 255 435
rect 227 423 231 427
rect 907 431 911 435
rect 935 423 936 427
rect 936 423 939 427
rect 1483 423 1487 427
rect 1915 423 1916 427
rect 1916 423 1919 427
rect 111 416 115 420
rect 155 415 159 419
rect 483 415 487 419
rect 811 415 815 419
rect 1139 415 1143 419
rect 1475 415 1479 419
rect 1787 415 1791 419
rect 1935 416 1939 420
rect 3203 411 3207 415
rect 4651 411 4655 415
rect 4851 411 4855 415
rect 5059 411 5063 415
rect 5119 411 5123 415
rect 5395 411 5396 415
rect 5396 411 5399 415
rect 5595 411 5599 415
rect 111 399 115 403
rect 183 400 187 404
rect 511 400 515 404
rect 839 400 843 404
rect 1167 400 1171 404
rect 1503 400 1507 404
rect 1815 400 1819 404
rect 1935 399 1939 403
rect 2211 403 2215 407
rect 2435 403 2439 407
rect 2659 403 2663 407
rect 2687 403 2691 407
rect 3075 403 3079 407
rect 3275 403 3279 407
rect 3475 403 3479 407
rect 1975 396 1979 400
rect 1995 395 1999 399
rect 2203 395 2207 399
rect 2427 395 2431 399
rect 2651 395 2655 399
rect 2859 395 2863 399
rect 3067 395 3071 399
rect 3267 395 3271 399
rect 3467 395 3471 399
rect 3635 399 3639 403
rect 3839 404 3843 408
rect 4451 403 4455 407
rect 4643 403 4647 407
rect 4843 403 4847 407
rect 5051 403 5055 407
rect 5267 403 5271 407
rect 5483 403 5487 407
rect 5663 404 5667 408
rect 3651 395 3655 399
rect 3799 396 3803 400
rect 3839 387 3843 391
rect 4479 388 4483 392
rect 4671 388 4675 392
rect 4871 388 4875 392
rect 5079 388 5083 392
rect 5295 388 5299 392
rect 5511 388 5515 392
rect 5663 387 5667 391
rect 1975 379 1979 383
rect 2023 380 2027 384
rect 2231 380 2235 384
rect 2455 380 2459 384
rect 2679 380 2683 384
rect 2887 380 2891 384
rect 3095 380 3099 384
rect 3295 380 3299 384
rect 3495 380 3499 384
rect 3679 380 3683 384
rect 3799 379 3803 383
rect 111 329 115 333
rect 279 328 283 332
rect 487 328 491 332
rect 703 328 707 332
rect 919 328 923 332
rect 1135 328 1139 332
rect 1935 329 1939 333
rect 3839 325 3843 329
rect 4615 324 4619 328
rect 4775 324 4779 328
rect 4951 324 4955 328
rect 5135 324 5139 328
rect 5327 324 5331 328
rect 5527 324 5531 328
rect 5663 325 5667 329
rect 111 312 115 316
rect 251 313 255 317
rect 459 313 463 317
rect 675 313 679 317
rect 891 313 895 317
rect 1107 313 1111 317
rect 1935 312 1939 316
rect 579 303 583 307
rect 1063 303 1067 307
rect 771 295 775 299
rect 1975 305 1979 309
rect 2023 304 2027 308
rect 2159 304 2163 308
rect 2295 304 2299 308
rect 2431 304 2435 308
rect 2567 304 2571 308
rect 2703 304 2707 308
rect 2839 304 2843 308
rect 2975 304 2979 308
rect 3111 304 3115 308
rect 3247 304 3251 308
rect 3383 304 3387 308
rect 3519 304 3523 308
rect 3655 304 3659 308
rect 3799 305 3803 309
rect 3839 308 3843 312
rect 4587 309 4591 313
rect 4747 309 4751 313
rect 4923 309 4927 313
rect 5107 309 5111 313
rect 5299 309 5303 313
rect 5499 309 5503 313
rect 5663 308 5667 312
rect 4735 299 4739 303
rect 4875 299 4876 303
rect 4876 299 4879 303
rect 5051 299 5052 303
rect 5052 299 5055 303
rect 1975 288 1979 292
rect 1995 289 1999 293
rect 2131 289 2135 293
rect 2267 289 2271 293
rect 2403 289 2407 293
rect 2539 289 2543 293
rect 2675 289 2679 293
rect 2811 289 2815 293
rect 2947 289 2951 293
rect 3083 289 3087 293
rect 3219 289 3223 293
rect 3355 289 3359 293
rect 3491 289 3495 293
rect 3627 289 3631 293
rect 3799 288 3803 292
rect 4675 291 4679 295
rect 5611 299 5615 303
rect 2123 279 2124 283
rect 2124 279 2127 283
rect 2259 279 2260 283
rect 2260 279 2263 283
rect 2395 279 2396 283
rect 2396 279 2399 283
rect 2531 279 2532 283
rect 2532 279 2535 283
rect 2667 279 2668 283
rect 2668 279 2671 283
rect 2803 279 2804 283
rect 2804 279 2807 283
rect 2855 279 2859 283
rect 3075 279 3076 283
rect 3076 279 3079 283
rect 3211 279 3212 283
rect 3212 279 3215 283
rect 3347 279 3348 283
rect 3348 279 3351 283
rect 3483 279 3484 283
rect 3484 279 3487 283
rect 2091 271 2095 275
rect 2687 271 2691 275
rect 347 263 351 267
rect 771 263 775 267
rect 935 263 939 267
rect 1063 263 1067 267
rect 2955 263 2959 267
rect 4387 251 4391 255
rect 4675 251 4679 255
rect 4735 259 4739 263
rect 4875 259 4879 263
rect 5051 259 5055 263
rect 5595 259 5599 263
rect 5119 251 5123 255
rect 2091 239 2095 243
rect 2123 239 2127 243
rect 2259 239 2263 243
rect 2395 239 2399 243
rect 2531 239 2535 243
rect 2667 239 2671 243
rect 2803 239 2807 243
rect 3043 239 3047 243
rect 3075 239 3079 243
rect 3211 239 3215 243
rect 3347 239 3351 243
rect 3483 239 3487 243
rect 2091 231 2095 235
rect 2855 231 2859 235
rect 227 187 231 191
rect 275 187 279 191
rect 1207 199 1211 203
rect 635 187 639 191
rect 955 187 959 191
rect 1091 187 1095 191
rect 4387 187 4391 191
rect 4435 183 4439 187
rect 4571 183 4575 187
rect 4707 183 4711 187
rect 4843 183 4847 187
rect 4979 183 4983 187
rect 5115 183 5119 187
rect 5251 183 5255 187
rect 5475 183 5479 187
rect 5611 187 5615 191
rect 2091 171 2095 175
rect 2139 167 2143 171
rect 2275 167 2279 171
rect 2411 167 2415 171
rect 2547 167 2551 171
rect 2683 167 2687 171
rect 2819 167 2823 171
rect 2955 167 2959 171
rect 3091 167 3095 171
rect 3227 167 3231 171
rect 3363 167 3367 171
rect 3499 167 3503 171
rect 3635 167 3639 171
rect 227 155 231 159
rect 275 147 279 151
rect 347 147 351 151
rect 635 155 639 159
rect 955 147 959 151
rect 1091 147 1095 151
rect 1207 147 1208 151
rect 1208 147 1211 151
rect 111 140 115 144
rect 131 139 135 143
rect 267 139 271 143
rect 403 139 407 143
rect 539 139 543 143
rect 675 139 679 143
rect 811 139 815 143
rect 947 139 951 143
rect 1083 139 1087 143
rect 1935 140 1939 144
rect 4435 143 4439 147
rect 4571 143 4575 147
rect 4707 143 4711 147
rect 4843 143 4847 147
rect 4979 143 4983 147
rect 5115 143 5119 147
rect 5251 143 5255 147
rect 5363 143 5367 147
rect 5475 143 5479 147
rect 3839 136 3843 140
rect 4291 135 4295 139
rect 4427 135 4431 139
rect 4563 135 4567 139
rect 4699 135 4703 139
rect 4835 135 4839 139
rect 4971 135 4975 139
rect 5107 135 5111 139
rect 5243 135 5247 139
rect 5379 135 5383 139
rect 5515 135 5519 139
rect 5663 136 5667 140
rect 111 123 115 127
rect 159 124 163 128
rect 295 124 299 128
rect 431 124 435 128
rect 567 124 571 128
rect 703 124 707 128
rect 839 124 843 128
rect 975 124 979 128
rect 1111 124 1115 128
rect 1935 123 1939 127
rect 2139 127 2143 131
rect 2275 127 2279 131
rect 2411 127 2415 131
rect 2547 127 2551 131
rect 2683 127 2687 131
rect 2819 127 2823 131
rect 2955 127 2959 131
rect 3091 127 3095 131
rect 3227 127 3231 131
rect 3363 127 3367 131
rect 3499 127 3503 131
rect 3635 127 3639 131
rect 3647 127 3651 131
rect 1975 120 1979 124
rect 1995 119 1999 123
rect 2131 119 2135 123
rect 2267 119 2271 123
rect 2403 119 2407 123
rect 2539 119 2543 123
rect 2675 119 2679 123
rect 2811 119 2815 123
rect 2947 119 2951 123
rect 3083 119 3087 123
rect 3219 119 3223 123
rect 3355 119 3359 123
rect 3491 119 3495 123
rect 3627 119 3631 123
rect 3799 120 3803 124
rect 3839 119 3843 123
rect 4319 120 4323 124
rect 4455 120 4459 124
rect 4591 120 4595 124
rect 4727 120 4731 124
rect 4863 120 4867 124
rect 4999 120 5003 124
rect 5135 120 5139 124
rect 5271 120 5275 124
rect 5407 120 5411 124
rect 5543 120 5547 124
rect 5663 119 5667 123
rect 1975 103 1979 107
rect 2023 104 2027 108
rect 2159 104 2163 108
rect 2295 104 2299 108
rect 2431 104 2435 108
rect 2567 104 2571 108
rect 2703 104 2707 108
rect 2839 104 2843 108
rect 2975 104 2979 108
rect 3111 104 3115 108
rect 3247 104 3251 108
rect 3383 104 3387 108
rect 3519 104 3523 108
rect 3655 104 3659 108
rect 3799 103 3803 107
<< m3 >>
rect 111 5758 115 5759
rect 111 5753 115 5754
rect 159 5758 163 5759
rect 159 5753 163 5754
rect 295 5758 299 5759
rect 295 5753 299 5754
rect 1935 5758 1939 5759
rect 1935 5753 1939 5754
rect 112 5730 114 5753
rect 110 5729 116 5730
rect 160 5729 162 5753
rect 296 5729 298 5753
rect 1936 5730 1938 5753
rect 1934 5729 1940 5730
rect 110 5725 111 5729
rect 115 5725 116 5729
rect 110 5724 116 5725
rect 158 5728 164 5729
rect 158 5724 159 5728
rect 163 5724 164 5728
rect 158 5723 164 5724
rect 294 5728 300 5729
rect 294 5724 295 5728
rect 299 5724 300 5728
rect 1934 5725 1935 5729
rect 1939 5725 1940 5729
rect 1934 5724 1940 5725
rect 294 5723 300 5724
rect 130 5713 136 5714
rect 110 5712 116 5713
rect 110 5708 111 5712
rect 115 5708 116 5712
rect 130 5709 131 5713
rect 135 5709 136 5713
rect 130 5708 136 5709
rect 266 5713 272 5714
rect 266 5709 267 5713
rect 271 5709 272 5713
rect 266 5708 272 5709
rect 1934 5712 1940 5713
rect 1934 5708 1935 5712
rect 1939 5708 1940 5712
rect 110 5707 116 5708
rect 112 5647 114 5707
rect 132 5647 134 5708
rect 268 5647 270 5708
rect 1934 5707 1940 5708
rect 378 5703 384 5704
rect 378 5699 379 5703
rect 383 5699 384 5703
rect 378 5698 384 5699
rect 111 5646 115 5647
rect 111 5641 115 5642
rect 131 5646 135 5647
rect 131 5641 135 5642
rect 267 5646 271 5647
rect 267 5641 271 5642
rect 275 5646 279 5647
rect 275 5641 279 5642
rect 112 5581 114 5641
rect 110 5580 116 5581
rect 132 5580 134 5641
rect 276 5580 278 5641
rect 380 5636 382 5698
rect 1936 5647 1938 5707
rect 1975 5658 1979 5659
rect 1975 5653 1979 5654
rect 2023 5658 2027 5659
rect 2023 5653 2027 5654
rect 2183 5658 2187 5659
rect 2183 5653 2187 5654
rect 2367 5658 2371 5659
rect 2367 5653 2371 5654
rect 2551 5658 2555 5659
rect 2551 5653 2555 5654
rect 2727 5658 2731 5659
rect 2727 5653 2731 5654
rect 2895 5658 2899 5659
rect 2895 5653 2899 5654
rect 3063 5658 3067 5659
rect 3063 5653 3067 5654
rect 3223 5658 3227 5659
rect 3223 5653 3227 5654
rect 3383 5658 3387 5659
rect 3383 5653 3387 5654
rect 3543 5658 3547 5659
rect 3543 5653 3547 5654
rect 3679 5658 3683 5659
rect 3679 5653 3683 5654
rect 3799 5658 3803 5659
rect 3799 5653 3803 5654
rect 3839 5654 3843 5655
rect 475 5646 479 5647
rect 475 5641 479 5642
rect 699 5646 703 5647
rect 699 5641 703 5642
rect 955 5646 959 5647
rect 955 5641 959 5642
rect 1227 5646 1231 5647
rect 1227 5641 1231 5642
rect 1515 5646 1519 5647
rect 1515 5641 1519 5642
rect 1787 5646 1791 5647
rect 1787 5641 1791 5642
rect 1935 5646 1939 5647
rect 1935 5641 1939 5642
rect 378 5635 384 5636
rect 378 5631 379 5635
rect 383 5631 384 5635
rect 378 5630 384 5631
rect 282 5627 288 5628
rect 282 5623 283 5627
rect 287 5623 288 5627
rect 282 5622 288 5623
rect 284 5588 286 5622
rect 282 5587 288 5588
rect 282 5583 283 5587
rect 287 5583 288 5587
rect 282 5582 288 5583
rect 476 5580 478 5641
rect 482 5627 488 5628
rect 482 5623 483 5627
rect 487 5623 488 5627
rect 482 5622 488 5623
rect 484 5588 486 5622
rect 482 5587 488 5588
rect 482 5583 483 5587
rect 487 5583 488 5587
rect 482 5582 488 5583
rect 700 5580 702 5641
rect 706 5627 712 5628
rect 706 5623 707 5627
rect 711 5623 712 5627
rect 706 5622 712 5623
rect 708 5588 710 5622
rect 706 5587 712 5588
rect 706 5583 707 5587
rect 711 5583 712 5587
rect 706 5582 712 5583
rect 956 5580 958 5641
rect 962 5627 968 5628
rect 962 5623 963 5627
rect 967 5623 968 5627
rect 962 5622 968 5623
rect 964 5588 966 5622
rect 962 5587 968 5588
rect 962 5583 963 5587
rect 967 5583 968 5587
rect 962 5582 968 5583
rect 1228 5580 1230 5641
rect 1234 5627 1240 5628
rect 1234 5623 1235 5627
rect 1239 5623 1240 5627
rect 1234 5622 1240 5623
rect 1236 5588 1238 5622
rect 1234 5587 1240 5588
rect 1234 5583 1235 5587
rect 1239 5583 1240 5587
rect 1234 5582 1240 5583
rect 1278 5587 1284 5588
rect 1278 5583 1279 5587
rect 1283 5583 1284 5587
rect 1278 5582 1284 5583
rect 110 5576 111 5580
rect 115 5576 116 5580
rect 110 5575 116 5576
rect 130 5579 136 5580
rect 130 5575 131 5579
rect 135 5575 136 5579
rect 130 5574 136 5575
rect 274 5579 280 5580
rect 274 5575 275 5579
rect 279 5575 280 5579
rect 274 5574 280 5575
rect 474 5579 480 5580
rect 474 5575 475 5579
rect 479 5575 480 5579
rect 474 5574 480 5575
rect 698 5579 704 5580
rect 698 5575 699 5579
rect 703 5575 704 5579
rect 698 5574 704 5575
rect 954 5579 960 5580
rect 954 5575 955 5579
rect 959 5575 960 5579
rect 954 5574 960 5575
rect 1226 5579 1232 5580
rect 1226 5575 1227 5579
rect 1231 5575 1232 5579
rect 1226 5574 1232 5575
rect 158 5564 164 5565
rect 110 5563 116 5564
rect 110 5559 111 5563
rect 115 5559 116 5563
rect 158 5560 159 5564
rect 163 5560 164 5564
rect 158 5559 164 5560
rect 302 5564 308 5565
rect 302 5560 303 5564
rect 307 5560 308 5564
rect 302 5559 308 5560
rect 502 5564 508 5565
rect 502 5560 503 5564
rect 507 5560 508 5564
rect 502 5559 508 5560
rect 726 5564 732 5565
rect 726 5560 727 5564
rect 731 5560 732 5564
rect 726 5559 732 5560
rect 982 5564 988 5565
rect 982 5560 983 5564
rect 987 5560 988 5564
rect 982 5559 988 5560
rect 1254 5564 1260 5565
rect 1254 5560 1255 5564
rect 1259 5560 1260 5564
rect 1254 5559 1260 5560
rect 110 5558 116 5559
rect 112 5535 114 5558
rect 160 5535 162 5559
rect 304 5535 306 5559
rect 504 5535 506 5559
rect 728 5535 730 5559
rect 984 5535 986 5559
rect 1256 5535 1258 5559
rect 111 5534 115 5535
rect 111 5529 115 5530
rect 159 5534 163 5535
rect 159 5529 163 5530
rect 279 5534 283 5535
rect 279 5529 283 5530
rect 303 5534 307 5535
rect 303 5529 307 5530
rect 503 5534 507 5535
rect 503 5529 507 5530
rect 519 5534 523 5535
rect 519 5529 523 5530
rect 727 5534 731 5535
rect 727 5529 731 5530
rect 767 5534 771 5535
rect 767 5529 771 5530
rect 983 5534 987 5535
rect 983 5529 987 5530
rect 1015 5534 1019 5535
rect 1015 5529 1019 5530
rect 1255 5534 1259 5535
rect 1255 5529 1259 5530
rect 1263 5534 1267 5535
rect 1263 5529 1267 5530
rect 112 5506 114 5529
rect 110 5505 116 5506
rect 280 5505 282 5529
rect 520 5505 522 5529
rect 768 5505 770 5529
rect 1016 5505 1018 5529
rect 1264 5505 1266 5529
rect 110 5501 111 5505
rect 115 5501 116 5505
rect 110 5500 116 5501
rect 278 5504 284 5505
rect 278 5500 279 5504
rect 283 5500 284 5504
rect 278 5499 284 5500
rect 518 5504 524 5505
rect 518 5500 519 5504
rect 523 5500 524 5504
rect 518 5499 524 5500
rect 766 5504 772 5505
rect 766 5500 767 5504
rect 771 5500 772 5504
rect 766 5499 772 5500
rect 1014 5504 1020 5505
rect 1014 5500 1015 5504
rect 1019 5500 1020 5504
rect 1014 5499 1020 5500
rect 1262 5504 1268 5505
rect 1262 5500 1263 5504
rect 1267 5500 1268 5504
rect 1262 5499 1268 5500
rect 250 5489 256 5490
rect 110 5488 116 5489
rect 110 5484 111 5488
rect 115 5484 116 5488
rect 250 5485 251 5489
rect 255 5485 256 5489
rect 250 5484 256 5485
rect 490 5489 496 5490
rect 490 5485 491 5489
rect 495 5485 496 5489
rect 490 5484 496 5485
rect 738 5489 744 5490
rect 738 5485 739 5489
rect 743 5485 744 5489
rect 738 5484 744 5485
rect 986 5489 992 5490
rect 986 5485 987 5489
rect 991 5485 992 5489
rect 986 5484 992 5485
rect 1234 5489 1240 5490
rect 1234 5485 1235 5489
rect 1239 5485 1240 5489
rect 1234 5484 1240 5485
rect 110 5483 116 5484
rect 112 5423 114 5483
rect 252 5423 254 5484
rect 378 5479 384 5480
rect 378 5475 379 5479
rect 383 5475 384 5479
rect 378 5474 384 5475
rect 380 5440 382 5474
rect 378 5439 384 5440
rect 378 5435 379 5439
rect 383 5435 384 5439
rect 378 5434 384 5435
rect 492 5423 494 5484
rect 618 5479 624 5480
rect 618 5475 619 5479
rect 623 5475 624 5479
rect 618 5474 624 5475
rect 506 5471 512 5472
rect 506 5467 507 5471
rect 511 5467 512 5471
rect 506 5466 512 5467
rect 111 5422 115 5423
rect 111 5417 115 5418
rect 251 5422 255 5423
rect 251 5417 255 5418
rect 411 5422 415 5423
rect 411 5417 415 5418
rect 491 5422 495 5423
rect 491 5417 495 5418
rect 112 5357 114 5417
rect 110 5356 116 5357
rect 412 5356 414 5417
rect 508 5408 510 5466
rect 620 5440 622 5474
rect 618 5439 624 5440
rect 618 5435 619 5439
rect 623 5435 624 5439
rect 618 5434 624 5435
rect 740 5423 742 5484
rect 866 5479 872 5480
rect 866 5475 867 5479
rect 871 5475 872 5479
rect 866 5474 872 5475
rect 868 5440 870 5474
rect 866 5439 872 5440
rect 866 5435 867 5439
rect 871 5435 872 5439
rect 866 5434 872 5435
rect 988 5423 990 5484
rect 1236 5423 1238 5484
rect 1280 5432 1282 5582
rect 1516 5580 1518 5641
rect 1778 5631 1784 5632
rect 1778 5627 1779 5631
rect 1783 5627 1784 5631
rect 1778 5626 1784 5627
rect 1514 5579 1520 5580
rect 1514 5575 1515 5579
rect 1519 5575 1520 5579
rect 1514 5574 1520 5575
rect 1542 5564 1548 5565
rect 1542 5560 1543 5564
rect 1547 5560 1548 5564
rect 1542 5559 1548 5560
rect 1544 5535 1546 5559
rect 1511 5534 1515 5535
rect 1511 5529 1515 5530
rect 1543 5534 1547 5535
rect 1543 5529 1547 5530
rect 1767 5534 1771 5535
rect 1767 5529 1771 5530
rect 1512 5505 1514 5529
rect 1768 5505 1770 5529
rect 1510 5504 1516 5505
rect 1510 5500 1511 5504
rect 1515 5500 1516 5504
rect 1510 5499 1516 5500
rect 1766 5504 1772 5505
rect 1766 5500 1767 5504
rect 1771 5500 1772 5504
rect 1766 5499 1772 5500
rect 1482 5489 1488 5490
rect 1482 5485 1483 5489
rect 1487 5485 1488 5489
rect 1482 5484 1488 5485
rect 1738 5489 1744 5490
rect 1738 5485 1739 5489
rect 1743 5485 1744 5489
rect 1738 5484 1744 5485
rect 1362 5479 1368 5480
rect 1362 5475 1363 5479
rect 1367 5475 1368 5479
rect 1362 5474 1368 5475
rect 1364 5440 1366 5474
rect 1330 5439 1336 5440
rect 1330 5435 1331 5439
rect 1335 5435 1336 5439
rect 1330 5434 1336 5435
rect 1362 5439 1368 5440
rect 1362 5435 1363 5439
rect 1367 5435 1368 5439
rect 1362 5434 1368 5435
rect 1278 5431 1284 5432
rect 1278 5427 1279 5431
rect 1283 5427 1284 5431
rect 1278 5426 1284 5427
rect 611 5422 615 5423
rect 611 5417 615 5418
rect 739 5422 743 5423
rect 739 5417 743 5418
rect 819 5422 823 5423
rect 819 5417 823 5418
rect 987 5422 991 5423
rect 987 5417 991 5418
rect 1035 5422 1039 5423
rect 1035 5417 1039 5418
rect 1235 5422 1239 5423
rect 1235 5417 1239 5418
rect 1259 5422 1263 5423
rect 1259 5417 1263 5418
rect 506 5407 512 5408
rect 506 5403 507 5407
rect 511 5403 512 5407
rect 506 5402 512 5403
rect 612 5356 614 5417
rect 618 5403 624 5404
rect 618 5399 619 5403
rect 623 5399 624 5403
rect 618 5398 624 5399
rect 620 5364 622 5398
rect 658 5371 664 5372
rect 658 5367 659 5371
rect 663 5367 664 5371
rect 658 5366 664 5367
rect 618 5363 624 5364
rect 618 5359 619 5363
rect 623 5359 624 5363
rect 618 5358 624 5359
rect 110 5352 111 5356
rect 115 5352 116 5356
rect 110 5351 116 5352
rect 410 5355 416 5356
rect 410 5351 411 5355
rect 415 5351 416 5355
rect 410 5350 416 5351
rect 610 5355 616 5356
rect 610 5351 611 5355
rect 615 5351 616 5355
rect 610 5350 616 5351
rect 438 5340 444 5341
rect 110 5339 116 5340
rect 110 5335 111 5339
rect 115 5335 116 5339
rect 438 5336 439 5340
rect 443 5336 444 5340
rect 438 5335 444 5336
rect 638 5340 644 5341
rect 638 5336 639 5340
rect 643 5336 644 5340
rect 638 5335 644 5336
rect 110 5334 116 5335
rect 112 5311 114 5334
rect 440 5311 442 5335
rect 640 5311 642 5335
rect 111 5310 115 5311
rect 111 5305 115 5306
rect 439 5310 443 5311
rect 439 5305 443 5306
rect 591 5310 595 5311
rect 591 5305 595 5306
rect 639 5310 643 5311
rect 639 5305 643 5306
rect 112 5282 114 5305
rect 110 5281 116 5282
rect 592 5281 594 5305
rect 110 5277 111 5281
rect 115 5277 116 5281
rect 110 5276 116 5277
rect 590 5280 596 5281
rect 590 5276 591 5280
rect 595 5276 596 5280
rect 590 5275 596 5276
rect 562 5265 568 5266
rect 110 5264 116 5265
rect 110 5260 111 5264
rect 115 5260 116 5264
rect 562 5261 563 5265
rect 567 5261 568 5265
rect 562 5260 568 5261
rect 110 5259 116 5260
rect 112 5095 114 5259
rect 564 5095 566 5260
rect 660 5216 662 5366
rect 820 5356 822 5417
rect 826 5403 832 5404
rect 826 5399 827 5403
rect 831 5399 832 5403
rect 826 5398 832 5399
rect 828 5364 830 5398
rect 826 5363 832 5364
rect 826 5359 827 5363
rect 831 5359 832 5363
rect 826 5358 832 5359
rect 1036 5356 1038 5417
rect 1042 5403 1048 5404
rect 1042 5399 1043 5403
rect 1047 5399 1048 5403
rect 1042 5398 1048 5399
rect 1044 5364 1046 5398
rect 1042 5363 1048 5364
rect 1042 5359 1043 5363
rect 1047 5359 1048 5363
rect 1042 5358 1048 5359
rect 1260 5356 1262 5417
rect 1332 5364 1334 5434
rect 1484 5423 1486 5484
rect 1610 5479 1616 5480
rect 1610 5475 1611 5479
rect 1615 5475 1616 5479
rect 1610 5474 1616 5475
rect 1612 5440 1614 5474
rect 1610 5439 1616 5440
rect 1610 5435 1611 5439
rect 1615 5435 1616 5439
rect 1610 5434 1616 5435
rect 1740 5423 1742 5484
rect 1780 5480 1782 5626
rect 1788 5580 1790 5641
rect 1794 5627 1800 5628
rect 1794 5623 1795 5627
rect 1799 5623 1800 5627
rect 1794 5622 1800 5623
rect 1796 5588 1798 5622
rect 1794 5587 1800 5588
rect 1794 5583 1795 5587
rect 1799 5583 1800 5587
rect 1794 5582 1800 5583
rect 1936 5581 1938 5641
rect 1976 5630 1978 5653
rect 1974 5629 1980 5630
rect 2024 5629 2026 5653
rect 2184 5629 2186 5653
rect 2368 5629 2370 5653
rect 2552 5629 2554 5653
rect 2728 5629 2730 5653
rect 2896 5629 2898 5653
rect 3064 5629 3066 5653
rect 3224 5629 3226 5653
rect 3384 5629 3386 5653
rect 3544 5629 3546 5653
rect 3680 5629 3682 5653
rect 3800 5630 3802 5653
rect 3839 5649 3843 5650
rect 4335 5654 4339 5655
rect 4335 5649 4339 5650
rect 4471 5654 4475 5655
rect 4471 5649 4475 5650
rect 4607 5654 4611 5655
rect 4607 5649 4611 5650
rect 4743 5654 4747 5655
rect 4743 5649 4747 5650
rect 4879 5654 4883 5655
rect 4879 5649 4883 5650
rect 5015 5654 5019 5655
rect 5015 5649 5019 5650
rect 5663 5654 5667 5655
rect 5663 5649 5667 5650
rect 3798 5629 3804 5630
rect 1974 5625 1975 5629
rect 1979 5625 1980 5629
rect 1974 5624 1980 5625
rect 2022 5628 2028 5629
rect 2022 5624 2023 5628
rect 2027 5624 2028 5628
rect 2022 5623 2028 5624
rect 2182 5628 2188 5629
rect 2182 5624 2183 5628
rect 2187 5624 2188 5628
rect 2182 5623 2188 5624
rect 2366 5628 2372 5629
rect 2366 5624 2367 5628
rect 2371 5624 2372 5628
rect 2366 5623 2372 5624
rect 2550 5628 2556 5629
rect 2550 5624 2551 5628
rect 2555 5624 2556 5628
rect 2550 5623 2556 5624
rect 2726 5628 2732 5629
rect 2726 5624 2727 5628
rect 2731 5624 2732 5628
rect 2726 5623 2732 5624
rect 2894 5628 2900 5629
rect 2894 5624 2895 5628
rect 2899 5624 2900 5628
rect 2894 5623 2900 5624
rect 3062 5628 3068 5629
rect 3062 5624 3063 5628
rect 3067 5624 3068 5628
rect 3062 5623 3068 5624
rect 3222 5628 3228 5629
rect 3222 5624 3223 5628
rect 3227 5624 3228 5628
rect 3222 5623 3228 5624
rect 3382 5628 3388 5629
rect 3382 5624 3383 5628
rect 3387 5624 3388 5628
rect 3382 5623 3388 5624
rect 3542 5628 3548 5629
rect 3542 5624 3543 5628
rect 3547 5624 3548 5628
rect 3542 5623 3548 5624
rect 3678 5628 3684 5629
rect 3678 5624 3679 5628
rect 3683 5624 3684 5628
rect 3798 5625 3799 5629
rect 3803 5625 3804 5629
rect 3840 5626 3842 5649
rect 3798 5624 3804 5625
rect 3838 5625 3844 5626
rect 4336 5625 4338 5649
rect 4472 5625 4474 5649
rect 4608 5625 4610 5649
rect 4744 5625 4746 5649
rect 4880 5625 4882 5649
rect 5016 5625 5018 5649
rect 5664 5626 5666 5649
rect 5662 5625 5668 5626
rect 3678 5623 3684 5624
rect 3838 5621 3839 5625
rect 3843 5621 3844 5625
rect 3838 5620 3844 5621
rect 4334 5624 4340 5625
rect 4334 5620 4335 5624
rect 4339 5620 4340 5624
rect 4334 5619 4340 5620
rect 4470 5624 4476 5625
rect 4470 5620 4471 5624
rect 4475 5620 4476 5624
rect 4470 5619 4476 5620
rect 4606 5624 4612 5625
rect 4606 5620 4607 5624
rect 4611 5620 4612 5624
rect 4606 5619 4612 5620
rect 4742 5624 4748 5625
rect 4742 5620 4743 5624
rect 4747 5620 4748 5624
rect 4742 5619 4748 5620
rect 4878 5624 4884 5625
rect 4878 5620 4879 5624
rect 4883 5620 4884 5624
rect 4878 5619 4884 5620
rect 5014 5624 5020 5625
rect 5014 5620 5015 5624
rect 5019 5620 5020 5624
rect 5662 5621 5663 5625
rect 5667 5621 5668 5625
rect 5662 5620 5668 5621
rect 5014 5619 5020 5620
rect 1994 5613 2000 5614
rect 1974 5612 1980 5613
rect 1974 5608 1975 5612
rect 1979 5608 1980 5612
rect 1994 5609 1995 5613
rect 1999 5609 2000 5613
rect 1994 5608 2000 5609
rect 2154 5613 2160 5614
rect 2154 5609 2155 5613
rect 2159 5609 2160 5613
rect 2154 5608 2160 5609
rect 2338 5613 2344 5614
rect 2338 5609 2339 5613
rect 2343 5609 2344 5613
rect 2338 5608 2344 5609
rect 2522 5613 2528 5614
rect 2522 5609 2523 5613
rect 2527 5609 2528 5613
rect 2522 5608 2528 5609
rect 2698 5613 2704 5614
rect 2698 5609 2699 5613
rect 2703 5609 2704 5613
rect 2698 5608 2704 5609
rect 2866 5613 2872 5614
rect 2866 5609 2867 5613
rect 2871 5609 2872 5613
rect 2866 5608 2872 5609
rect 3034 5613 3040 5614
rect 3034 5609 3035 5613
rect 3039 5609 3040 5613
rect 3034 5608 3040 5609
rect 3194 5613 3200 5614
rect 3194 5609 3195 5613
rect 3199 5609 3200 5613
rect 3194 5608 3200 5609
rect 3354 5613 3360 5614
rect 3354 5609 3355 5613
rect 3359 5609 3360 5613
rect 3354 5608 3360 5609
rect 3514 5613 3520 5614
rect 3514 5609 3515 5613
rect 3519 5609 3520 5613
rect 3514 5608 3520 5609
rect 3650 5613 3656 5614
rect 3650 5609 3651 5613
rect 3655 5609 3656 5613
rect 3650 5608 3656 5609
rect 3798 5612 3804 5613
rect 3798 5608 3799 5612
rect 3803 5608 3804 5612
rect 4306 5609 4312 5610
rect 1974 5607 1980 5608
rect 1962 5587 1968 5588
rect 1962 5583 1963 5587
rect 1967 5583 1968 5587
rect 1962 5582 1968 5583
rect 1934 5580 1940 5581
rect 1786 5579 1792 5580
rect 1786 5575 1787 5579
rect 1791 5575 1792 5579
rect 1934 5576 1935 5580
rect 1939 5576 1940 5580
rect 1934 5575 1940 5576
rect 1786 5574 1792 5575
rect 1814 5564 1820 5565
rect 1964 5564 1966 5582
rect 1814 5560 1815 5564
rect 1819 5560 1820 5564
rect 1814 5559 1820 5560
rect 1934 5563 1940 5564
rect 1934 5559 1935 5563
rect 1939 5559 1940 5563
rect 1816 5535 1818 5559
rect 1934 5558 1940 5559
rect 1962 5563 1968 5564
rect 1962 5559 1963 5563
rect 1967 5559 1968 5563
rect 1962 5558 1968 5559
rect 1936 5535 1938 5558
rect 1976 5547 1978 5607
rect 1996 5547 1998 5608
rect 2142 5603 2148 5604
rect 2142 5599 2143 5603
rect 2147 5599 2148 5603
rect 2142 5598 2148 5599
rect 2144 5564 2146 5598
rect 2142 5563 2148 5564
rect 2142 5559 2143 5563
rect 2147 5559 2148 5563
rect 2142 5558 2148 5559
rect 2156 5547 2158 5608
rect 2282 5603 2288 5604
rect 2282 5599 2283 5603
rect 2287 5599 2288 5603
rect 2282 5598 2288 5599
rect 2284 5564 2286 5598
rect 2282 5563 2288 5564
rect 2282 5559 2283 5563
rect 2287 5559 2288 5563
rect 2282 5558 2288 5559
rect 2340 5547 2342 5608
rect 2466 5603 2472 5604
rect 2466 5599 2467 5603
rect 2471 5599 2472 5603
rect 2466 5598 2472 5599
rect 2468 5564 2470 5598
rect 2466 5563 2472 5564
rect 2466 5559 2467 5563
rect 2471 5559 2472 5563
rect 2466 5558 2472 5559
rect 2524 5547 2526 5608
rect 2646 5603 2652 5604
rect 2646 5599 2647 5603
rect 2651 5599 2652 5603
rect 2646 5598 2652 5599
rect 1975 5546 1979 5547
rect 1975 5541 1979 5542
rect 1995 5546 1999 5547
rect 1995 5541 1999 5542
rect 2139 5546 2143 5547
rect 2139 5541 2143 5542
rect 2155 5546 2159 5547
rect 2155 5541 2159 5542
rect 2339 5546 2343 5547
rect 2339 5541 2343 5542
rect 2355 5546 2359 5547
rect 2355 5541 2359 5542
rect 2523 5546 2527 5547
rect 2523 5541 2527 5542
rect 2563 5546 2567 5547
rect 2563 5541 2567 5542
rect 1815 5534 1819 5535
rect 1815 5529 1819 5530
rect 1935 5534 1939 5535
rect 1935 5529 1939 5530
rect 1936 5506 1938 5529
rect 1934 5505 1940 5506
rect 1934 5501 1935 5505
rect 1939 5501 1940 5505
rect 1934 5500 1940 5501
rect 1934 5488 1940 5489
rect 1934 5484 1935 5488
rect 1939 5484 1940 5488
rect 1934 5483 1940 5484
rect 1778 5479 1784 5480
rect 1778 5475 1779 5479
rect 1783 5475 1784 5479
rect 1778 5474 1784 5475
rect 1936 5423 1938 5483
rect 1976 5481 1978 5541
rect 1974 5480 1980 5481
rect 2140 5480 2142 5541
rect 2262 5487 2268 5488
rect 2262 5483 2263 5487
rect 2267 5483 2268 5487
rect 2262 5482 2268 5483
rect 1974 5476 1975 5480
rect 1979 5476 1980 5480
rect 1974 5475 1980 5476
rect 2138 5479 2144 5480
rect 2138 5475 2139 5479
rect 2143 5475 2144 5479
rect 2138 5474 2144 5475
rect 2166 5464 2172 5465
rect 1974 5463 1980 5464
rect 1974 5459 1975 5463
rect 1979 5459 1980 5463
rect 2166 5460 2167 5464
rect 2171 5460 2172 5464
rect 2166 5459 2172 5460
rect 1974 5458 1980 5459
rect 1976 5427 1978 5458
rect 2168 5427 2170 5459
rect 1975 5426 1979 5427
rect 1483 5422 1487 5423
rect 1483 5417 1487 5418
rect 1491 5422 1495 5423
rect 1491 5417 1495 5418
rect 1739 5422 1743 5423
rect 1739 5417 1743 5418
rect 1935 5422 1939 5423
rect 1975 5421 1979 5422
rect 2167 5426 2171 5427
rect 2167 5421 2171 5422
rect 1935 5417 1939 5418
rect 1330 5363 1336 5364
rect 1330 5359 1331 5363
rect 1335 5359 1336 5363
rect 1330 5358 1336 5359
rect 1492 5356 1494 5417
rect 1586 5403 1592 5404
rect 1586 5399 1587 5403
rect 1591 5399 1592 5403
rect 1586 5398 1592 5399
rect 818 5355 824 5356
rect 818 5351 819 5355
rect 823 5351 824 5355
rect 818 5350 824 5351
rect 1034 5355 1040 5356
rect 1034 5351 1035 5355
rect 1039 5351 1040 5355
rect 1034 5350 1040 5351
rect 1258 5355 1264 5356
rect 1258 5351 1259 5355
rect 1263 5351 1264 5355
rect 1258 5350 1264 5351
rect 1490 5355 1496 5356
rect 1490 5351 1491 5355
rect 1495 5351 1496 5355
rect 1490 5350 1496 5351
rect 846 5340 852 5341
rect 846 5336 847 5340
rect 851 5336 852 5340
rect 846 5335 852 5336
rect 1062 5340 1068 5341
rect 1062 5336 1063 5340
rect 1067 5336 1068 5340
rect 1062 5335 1068 5336
rect 1286 5340 1292 5341
rect 1286 5336 1287 5340
rect 1291 5336 1292 5340
rect 1286 5335 1292 5336
rect 1518 5340 1524 5341
rect 1518 5336 1519 5340
rect 1523 5336 1524 5340
rect 1518 5335 1524 5336
rect 848 5311 850 5335
rect 1064 5311 1066 5335
rect 1288 5311 1290 5335
rect 1520 5311 1522 5335
rect 727 5310 731 5311
rect 727 5305 731 5306
rect 847 5310 851 5311
rect 847 5305 851 5306
rect 863 5310 867 5311
rect 863 5305 867 5306
rect 999 5310 1003 5311
rect 999 5305 1003 5306
rect 1063 5310 1067 5311
rect 1063 5305 1067 5306
rect 1135 5310 1139 5311
rect 1135 5305 1139 5306
rect 1271 5310 1275 5311
rect 1271 5305 1275 5306
rect 1287 5310 1291 5311
rect 1287 5305 1291 5306
rect 1407 5310 1411 5311
rect 1407 5305 1411 5306
rect 1519 5310 1523 5311
rect 1519 5305 1523 5306
rect 1543 5310 1547 5311
rect 1543 5305 1547 5306
rect 728 5281 730 5305
rect 864 5281 866 5305
rect 1000 5281 1002 5305
rect 1136 5281 1138 5305
rect 1272 5281 1274 5305
rect 1408 5281 1410 5305
rect 1544 5281 1546 5305
rect 726 5280 732 5281
rect 726 5276 727 5280
rect 731 5276 732 5280
rect 726 5275 732 5276
rect 862 5280 868 5281
rect 862 5276 863 5280
rect 867 5276 868 5280
rect 862 5275 868 5276
rect 998 5280 1004 5281
rect 998 5276 999 5280
rect 1003 5276 1004 5280
rect 998 5275 1004 5276
rect 1134 5280 1140 5281
rect 1134 5276 1135 5280
rect 1139 5276 1140 5280
rect 1134 5275 1140 5276
rect 1270 5280 1276 5281
rect 1270 5276 1271 5280
rect 1275 5276 1276 5280
rect 1270 5275 1276 5276
rect 1406 5280 1412 5281
rect 1406 5276 1407 5280
rect 1411 5276 1412 5280
rect 1406 5275 1412 5276
rect 1542 5280 1548 5281
rect 1542 5276 1543 5280
rect 1547 5276 1548 5280
rect 1542 5275 1548 5276
rect 698 5265 704 5266
rect 698 5261 699 5265
rect 703 5261 704 5265
rect 698 5260 704 5261
rect 834 5265 840 5266
rect 834 5261 835 5265
rect 839 5261 840 5265
rect 834 5260 840 5261
rect 970 5265 976 5266
rect 970 5261 971 5265
rect 975 5261 976 5265
rect 970 5260 976 5261
rect 1106 5265 1112 5266
rect 1106 5261 1107 5265
rect 1111 5261 1112 5265
rect 1106 5260 1112 5261
rect 1242 5265 1248 5266
rect 1242 5261 1243 5265
rect 1247 5261 1248 5265
rect 1242 5260 1248 5261
rect 1378 5265 1384 5266
rect 1378 5261 1379 5265
rect 1383 5261 1384 5265
rect 1378 5260 1384 5261
rect 1514 5265 1520 5266
rect 1514 5261 1515 5265
rect 1519 5261 1520 5265
rect 1514 5260 1520 5261
rect 690 5255 696 5256
rect 690 5251 691 5255
rect 695 5251 696 5255
rect 690 5250 696 5251
rect 692 5216 694 5250
rect 658 5215 664 5216
rect 658 5211 659 5215
rect 663 5211 664 5215
rect 658 5210 664 5211
rect 690 5215 696 5216
rect 690 5211 691 5215
rect 695 5211 696 5215
rect 690 5210 696 5211
rect 700 5095 702 5260
rect 826 5255 832 5256
rect 826 5251 827 5255
rect 831 5251 832 5255
rect 826 5250 832 5251
rect 828 5216 830 5250
rect 826 5215 832 5216
rect 826 5211 827 5215
rect 831 5211 832 5215
rect 826 5210 832 5211
rect 836 5095 838 5260
rect 962 5255 968 5256
rect 962 5251 963 5255
rect 967 5251 968 5255
rect 962 5250 968 5251
rect 964 5216 966 5250
rect 962 5215 968 5216
rect 962 5211 963 5215
rect 967 5211 968 5215
rect 962 5210 968 5211
rect 972 5095 974 5260
rect 1108 5095 1110 5260
rect 1234 5255 1240 5256
rect 1234 5251 1235 5255
rect 1239 5251 1240 5255
rect 1234 5250 1240 5251
rect 1236 5216 1238 5250
rect 1234 5215 1240 5216
rect 1234 5211 1235 5215
rect 1239 5211 1240 5215
rect 1234 5210 1240 5211
rect 1244 5095 1246 5260
rect 1370 5255 1376 5256
rect 1370 5251 1371 5255
rect 1375 5251 1376 5255
rect 1370 5250 1376 5251
rect 1372 5216 1374 5250
rect 1370 5215 1376 5216
rect 1370 5211 1371 5215
rect 1375 5211 1376 5215
rect 1370 5210 1376 5211
rect 1380 5095 1382 5260
rect 1506 5255 1512 5256
rect 1506 5251 1507 5255
rect 1511 5251 1512 5255
rect 1506 5250 1512 5251
rect 1508 5216 1510 5250
rect 1506 5215 1512 5216
rect 1506 5211 1507 5215
rect 1511 5211 1512 5215
rect 1506 5210 1512 5211
rect 1516 5095 1518 5260
rect 1588 5256 1590 5398
rect 1936 5357 1938 5417
rect 1976 5398 1978 5421
rect 1974 5397 1980 5398
rect 1974 5393 1975 5397
rect 1979 5393 1980 5397
rect 1974 5392 1980 5393
rect 1974 5380 1980 5381
rect 1974 5376 1975 5380
rect 1979 5376 1980 5380
rect 1974 5375 1980 5376
rect 1934 5356 1940 5357
rect 1934 5352 1935 5356
rect 1939 5352 1940 5356
rect 1934 5351 1940 5352
rect 1934 5339 1940 5340
rect 1934 5335 1935 5339
rect 1939 5335 1940 5339
rect 1934 5334 1940 5335
rect 1936 5311 1938 5334
rect 1976 5315 1978 5375
rect 2264 5332 2266 5482
rect 2356 5480 2358 5541
rect 2564 5480 2566 5541
rect 2648 5532 2650 5598
rect 2700 5547 2702 5608
rect 2826 5603 2832 5604
rect 2826 5599 2827 5603
rect 2831 5599 2832 5603
rect 2826 5598 2832 5599
rect 2828 5564 2830 5598
rect 2794 5563 2800 5564
rect 2794 5559 2795 5563
rect 2799 5559 2800 5563
rect 2794 5558 2800 5559
rect 2826 5563 2832 5564
rect 2826 5559 2827 5563
rect 2831 5559 2832 5563
rect 2826 5558 2832 5559
rect 2699 5546 2703 5547
rect 2699 5541 2703 5542
rect 2755 5546 2759 5547
rect 2755 5541 2759 5542
rect 2646 5531 2652 5532
rect 2646 5527 2647 5531
rect 2651 5527 2652 5531
rect 2646 5526 2652 5527
rect 2756 5480 2758 5541
rect 2796 5488 2798 5558
rect 2868 5547 2870 5608
rect 2994 5603 3000 5604
rect 2994 5599 2995 5603
rect 2999 5599 3000 5603
rect 2994 5598 3000 5599
rect 2996 5564 2998 5598
rect 2994 5563 3000 5564
rect 2994 5559 2995 5563
rect 2999 5559 3000 5563
rect 2994 5558 3000 5559
rect 3036 5547 3038 5608
rect 3182 5603 3188 5604
rect 3182 5599 3183 5603
rect 3187 5599 3188 5603
rect 3182 5598 3188 5599
rect 3184 5564 3186 5598
rect 3182 5563 3188 5564
rect 3182 5559 3183 5563
rect 3187 5559 3188 5563
rect 3182 5558 3188 5559
rect 3196 5547 3198 5608
rect 3342 5603 3348 5604
rect 3342 5599 3343 5603
rect 3347 5599 3348 5603
rect 3342 5598 3348 5599
rect 3344 5564 3346 5598
rect 3342 5563 3348 5564
rect 3342 5559 3343 5563
rect 3347 5559 3348 5563
rect 3342 5558 3348 5559
rect 3356 5547 3358 5608
rect 3502 5603 3508 5604
rect 3502 5599 3503 5603
rect 3507 5599 3508 5603
rect 3502 5598 3508 5599
rect 3504 5564 3506 5598
rect 3502 5563 3508 5564
rect 3502 5559 3503 5563
rect 3507 5559 3508 5563
rect 3502 5558 3508 5559
rect 3516 5547 3518 5608
rect 3642 5603 3648 5604
rect 3642 5599 3643 5603
rect 3647 5599 3648 5603
rect 3642 5598 3648 5599
rect 3644 5564 3646 5598
rect 3642 5563 3648 5564
rect 3642 5559 3643 5563
rect 3647 5559 3648 5563
rect 3642 5558 3648 5559
rect 3652 5547 3654 5608
rect 3798 5607 3804 5608
rect 3838 5608 3844 5609
rect 3738 5603 3744 5604
rect 3738 5599 3739 5603
rect 3743 5599 3744 5603
rect 3738 5598 3744 5599
rect 2867 5546 2871 5547
rect 2867 5541 2871 5542
rect 2939 5546 2943 5547
rect 2939 5541 2943 5542
rect 3035 5546 3039 5547
rect 3035 5541 3039 5542
rect 3115 5546 3119 5547
rect 3115 5541 3119 5542
rect 3195 5546 3199 5547
rect 3195 5541 3199 5542
rect 3291 5546 3295 5547
rect 3291 5541 3295 5542
rect 3355 5546 3359 5547
rect 3355 5541 3359 5542
rect 3467 5546 3471 5547
rect 3467 5541 3471 5542
rect 3515 5546 3519 5547
rect 3515 5541 3519 5542
rect 3643 5546 3647 5547
rect 3643 5541 3647 5542
rect 3651 5546 3655 5547
rect 3651 5541 3655 5542
rect 2794 5487 2800 5488
rect 2794 5483 2795 5487
rect 2799 5483 2800 5487
rect 2794 5482 2800 5483
rect 2940 5480 2942 5541
rect 3116 5480 3118 5541
rect 3166 5531 3172 5532
rect 3166 5527 3167 5531
rect 3171 5527 3172 5531
rect 3166 5526 3172 5527
rect 2354 5479 2360 5480
rect 2354 5475 2355 5479
rect 2359 5475 2360 5479
rect 2354 5474 2360 5475
rect 2562 5479 2568 5480
rect 2562 5475 2563 5479
rect 2567 5475 2568 5479
rect 2562 5474 2568 5475
rect 2754 5479 2760 5480
rect 2754 5475 2755 5479
rect 2759 5475 2760 5479
rect 2754 5474 2760 5475
rect 2938 5479 2944 5480
rect 2938 5475 2939 5479
rect 2943 5475 2944 5479
rect 2938 5474 2944 5475
rect 3114 5479 3120 5480
rect 3114 5475 3115 5479
rect 3119 5475 3120 5479
rect 3114 5474 3120 5475
rect 2382 5464 2388 5465
rect 2382 5460 2383 5464
rect 2387 5460 2388 5464
rect 2382 5459 2388 5460
rect 2590 5464 2596 5465
rect 2590 5460 2591 5464
rect 2595 5460 2596 5464
rect 2590 5459 2596 5460
rect 2782 5464 2788 5465
rect 2782 5460 2783 5464
rect 2787 5460 2788 5464
rect 2782 5459 2788 5460
rect 2966 5464 2972 5465
rect 2966 5460 2967 5464
rect 2971 5460 2972 5464
rect 2966 5459 2972 5460
rect 3142 5464 3148 5465
rect 3142 5460 3143 5464
rect 3147 5460 3148 5464
rect 3142 5459 3148 5460
rect 2384 5427 2386 5459
rect 2592 5427 2594 5459
rect 2784 5427 2786 5459
rect 2968 5427 2970 5459
rect 3144 5427 3146 5459
rect 2311 5426 2315 5427
rect 2311 5421 2315 5422
rect 2383 5426 2387 5427
rect 2383 5421 2387 5422
rect 2511 5426 2515 5427
rect 2511 5421 2515 5422
rect 2591 5426 2595 5427
rect 2591 5421 2595 5422
rect 2703 5426 2707 5427
rect 2703 5421 2707 5422
rect 2783 5426 2787 5427
rect 2783 5421 2787 5422
rect 2887 5426 2891 5427
rect 2887 5421 2891 5422
rect 2967 5426 2971 5427
rect 2967 5421 2971 5422
rect 3071 5426 3075 5427
rect 3071 5421 3075 5422
rect 3143 5426 3147 5427
rect 3143 5421 3147 5422
rect 2312 5397 2314 5421
rect 2512 5397 2514 5421
rect 2704 5397 2706 5421
rect 2888 5397 2890 5421
rect 3072 5397 3074 5421
rect 2310 5396 2316 5397
rect 2310 5392 2311 5396
rect 2315 5392 2316 5396
rect 2310 5391 2316 5392
rect 2510 5396 2516 5397
rect 2510 5392 2511 5396
rect 2515 5392 2516 5396
rect 2510 5391 2516 5392
rect 2702 5396 2708 5397
rect 2702 5392 2703 5396
rect 2707 5392 2708 5396
rect 2702 5391 2708 5392
rect 2886 5396 2892 5397
rect 2886 5392 2887 5396
rect 2891 5392 2892 5396
rect 2886 5391 2892 5392
rect 3070 5396 3076 5397
rect 3070 5392 3071 5396
rect 3075 5392 3076 5396
rect 3070 5391 3076 5392
rect 2282 5381 2288 5382
rect 2282 5377 2283 5381
rect 2287 5377 2288 5381
rect 2282 5376 2288 5377
rect 2482 5381 2488 5382
rect 2482 5377 2483 5381
rect 2487 5377 2488 5381
rect 2482 5376 2488 5377
rect 2674 5381 2680 5382
rect 2674 5377 2675 5381
rect 2679 5377 2680 5381
rect 2674 5376 2680 5377
rect 2858 5381 2864 5382
rect 2858 5377 2859 5381
rect 2863 5377 2864 5381
rect 2858 5376 2864 5377
rect 3042 5381 3048 5382
rect 3042 5377 3043 5381
rect 3047 5377 3048 5381
rect 3042 5376 3048 5377
rect 2262 5331 2268 5332
rect 2262 5327 2263 5331
rect 2267 5327 2268 5331
rect 2262 5326 2268 5327
rect 2284 5315 2286 5376
rect 2442 5371 2448 5372
rect 2442 5367 2443 5371
rect 2447 5367 2448 5371
rect 2442 5366 2448 5367
rect 2444 5332 2446 5366
rect 2442 5331 2448 5332
rect 2442 5327 2443 5331
rect 2447 5327 2448 5331
rect 2442 5326 2448 5327
rect 2484 5315 2486 5376
rect 2610 5371 2616 5372
rect 2610 5367 2611 5371
rect 2615 5367 2616 5371
rect 2610 5366 2616 5367
rect 2612 5332 2614 5366
rect 2610 5331 2616 5332
rect 2610 5327 2611 5331
rect 2615 5327 2616 5331
rect 2610 5326 2616 5327
rect 2676 5315 2678 5376
rect 2810 5371 2816 5372
rect 2810 5367 2811 5371
rect 2815 5367 2816 5371
rect 2810 5366 2816 5367
rect 1975 5314 1979 5315
rect 1935 5310 1939 5311
rect 1975 5309 1979 5310
rect 2195 5314 2199 5315
rect 2195 5309 2199 5310
rect 2283 5314 2287 5315
rect 2283 5309 2287 5310
rect 2339 5314 2343 5315
rect 2339 5309 2343 5310
rect 2483 5314 2487 5315
rect 2483 5309 2487 5310
rect 2491 5314 2495 5315
rect 2491 5309 2495 5310
rect 2651 5314 2655 5315
rect 2651 5309 2655 5310
rect 2675 5314 2679 5315
rect 2675 5309 2679 5310
rect 1935 5305 1939 5306
rect 1936 5282 1938 5305
rect 1934 5281 1940 5282
rect 1934 5277 1935 5281
rect 1939 5277 1940 5281
rect 1934 5276 1940 5277
rect 1934 5264 1940 5265
rect 1934 5260 1935 5264
rect 1939 5260 1940 5264
rect 1934 5259 1940 5260
rect 1586 5255 1592 5256
rect 1586 5251 1587 5255
rect 1591 5251 1592 5255
rect 1586 5250 1592 5251
rect 1936 5095 1938 5259
rect 1976 5249 1978 5309
rect 1974 5248 1980 5249
rect 2196 5248 2198 5309
rect 2330 5299 2336 5300
rect 2330 5295 2331 5299
rect 2335 5295 2336 5299
rect 2330 5294 2336 5295
rect 2332 5256 2334 5294
rect 2318 5255 2324 5256
rect 2318 5251 2319 5255
rect 2323 5251 2324 5255
rect 2318 5250 2324 5251
rect 2330 5255 2336 5256
rect 2330 5251 2331 5255
rect 2335 5251 2336 5255
rect 2330 5250 2336 5251
rect 1974 5244 1975 5248
rect 1979 5244 1980 5248
rect 1974 5243 1980 5244
rect 2194 5247 2200 5248
rect 2194 5243 2195 5247
rect 2199 5243 2200 5247
rect 2194 5242 2200 5243
rect 2222 5232 2228 5233
rect 1974 5231 1980 5232
rect 1974 5227 1975 5231
rect 1979 5227 1980 5231
rect 2222 5228 2223 5232
rect 2227 5228 2228 5232
rect 2222 5227 2228 5228
rect 1974 5226 1980 5227
rect 1976 5203 1978 5226
rect 2224 5203 2226 5227
rect 1975 5202 1979 5203
rect 1975 5197 1979 5198
rect 2023 5202 2027 5203
rect 2023 5197 2027 5198
rect 2159 5202 2163 5203
rect 2159 5197 2163 5198
rect 2223 5202 2227 5203
rect 2223 5197 2227 5198
rect 1976 5174 1978 5197
rect 1974 5173 1980 5174
rect 2024 5173 2026 5197
rect 2160 5173 2162 5197
rect 1974 5169 1975 5173
rect 1979 5169 1980 5173
rect 1974 5168 1980 5169
rect 2022 5172 2028 5173
rect 2022 5168 2023 5172
rect 2027 5168 2028 5172
rect 2022 5167 2028 5168
rect 2158 5172 2164 5173
rect 2158 5168 2159 5172
rect 2163 5168 2164 5172
rect 2158 5167 2164 5168
rect 1994 5157 2000 5158
rect 1974 5156 1980 5157
rect 1974 5152 1975 5156
rect 1979 5152 1980 5156
rect 1994 5153 1995 5157
rect 1999 5153 2000 5157
rect 1994 5152 2000 5153
rect 2130 5157 2136 5158
rect 2130 5153 2131 5157
rect 2135 5153 2136 5157
rect 2130 5152 2136 5153
rect 2298 5157 2304 5158
rect 2298 5153 2299 5157
rect 2303 5153 2304 5157
rect 2298 5152 2304 5153
rect 1974 5151 1980 5152
rect 111 5094 115 5095
rect 111 5089 115 5090
rect 347 5094 351 5095
rect 347 5089 351 5090
rect 483 5094 487 5095
rect 483 5089 487 5090
rect 563 5094 567 5095
rect 563 5089 567 5090
rect 619 5094 623 5095
rect 619 5089 623 5090
rect 699 5094 703 5095
rect 699 5089 703 5090
rect 755 5094 759 5095
rect 755 5089 759 5090
rect 835 5094 839 5095
rect 835 5089 839 5090
rect 891 5094 895 5095
rect 891 5089 895 5090
rect 971 5094 975 5095
rect 971 5089 975 5090
rect 1035 5094 1039 5095
rect 1035 5089 1039 5090
rect 1107 5094 1111 5095
rect 1107 5089 1111 5090
rect 1187 5094 1191 5095
rect 1187 5089 1191 5090
rect 1243 5094 1247 5095
rect 1243 5089 1247 5090
rect 1339 5094 1343 5095
rect 1339 5089 1343 5090
rect 1379 5094 1383 5095
rect 1379 5089 1383 5090
rect 1491 5094 1495 5095
rect 1491 5089 1495 5090
rect 1515 5094 1519 5095
rect 1515 5089 1519 5090
rect 1651 5094 1655 5095
rect 1651 5089 1655 5090
rect 1787 5094 1791 5095
rect 1787 5089 1791 5090
rect 1935 5094 1939 5095
rect 1976 5091 1978 5151
rect 1996 5091 1998 5152
rect 2090 5147 2096 5148
rect 2090 5143 2091 5147
rect 2095 5143 2096 5147
rect 2090 5142 2096 5143
rect 1935 5089 1939 5090
rect 1975 5090 1979 5091
rect 112 5029 114 5089
rect 110 5028 116 5029
rect 348 5028 350 5089
rect 442 5075 448 5076
rect 442 5071 443 5075
rect 447 5071 448 5075
rect 442 5070 448 5071
rect 444 5044 446 5070
rect 442 5043 448 5044
rect 442 5039 443 5043
rect 447 5039 448 5043
rect 442 5038 448 5039
rect 484 5028 486 5089
rect 490 5075 496 5076
rect 490 5071 491 5075
rect 495 5071 496 5075
rect 490 5070 496 5071
rect 492 5036 494 5070
rect 490 5035 496 5036
rect 490 5031 491 5035
rect 495 5031 496 5035
rect 490 5030 496 5031
rect 606 5035 612 5036
rect 606 5031 607 5035
rect 611 5031 612 5035
rect 606 5030 612 5031
rect 110 5024 111 5028
rect 115 5024 116 5028
rect 110 5023 116 5024
rect 346 5027 352 5028
rect 346 5023 347 5027
rect 351 5023 352 5027
rect 346 5022 352 5023
rect 482 5027 488 5028
rect 482 5023 483 5027
rect 487 5023 488 5027
rect 482 5022 488 5023
rect 374 5012 380 5013
rect 110 5011 116 5012
rect 110 5007 111 5011
rect 115 5007 116 5011
rect 374 5008 375 5012
rect 379 5008 380 5012
rect 374 5007 380 5008
rect 510 5012 516 5013
rect 510 5008 511 5012
rect 515 5008 516 5012
rect 510 5007 516 5008
rect 110 5006 116 5007
rect 112 4983 114 5006
rect 376 4983 378 5007
rect 512 4983 514 5007
rect 111 4982 115 4983
rect 111 4977 115 4978
rect 159 4982 163 4983
rect 159 4977 163 4978
rect 343 4982 347 4983
rect 343 4977 347 4978
rect 375 4982 379 4983
rect 375 4977 379 4978
rect 511 4982 515 4983
rect 511 4977 515 4978
rect 551 4982 555 4983
rect 551 4977 555 4978
rect 112 4954 114 4977
rect 110 4953 116 4954
rect 160 4953 162 4977
rect 344 4953 346 4977
rect 552 4953 554 4977
rect 110 4949 111 4953
rect 115 4949 116 4953
rect 110 4948 116 4949
rect 158 4952 164 4953
rect 158 4948 159 4952
rect 163 4948 164 4952
rect 158 4947 164 4948
rect 342 4952 348 4953
rect 342 4948 343 4952
rect 347 4948 348 4952
rect 342 4947 348 4948
rect 550 4952 556 4953
rect 550 4948 551 4952
rect 555 4948 556 4952
rect 550 4947 556 4948
rect 130 4937 136 4938
rect 110 4936 116 4937
rect 110 4932 111 4936
rect 115 4932 116 4936
rect 130 4933 131 4937
rect 135 4933 136 4937
rect 130 4932 136 4933
rect 314 4937 320 4938
rect 314 4933 315 4937
rect 319 4933 320 4937
rect 314 4932 320 4933
rect 522 4937 528 4938
rect 522 4933 523 4937
rect 527 4933 528 4937
rect 522 4932 528 4933
rect 110 4931 116 4932
rect 112 4863 114 4931
rect 132 4863 134 4932
rect 226 4927 232 4928
rect 226 4923 227 4927
rect 231 4923 232 4927
rect 226 4922 232 4923
rect 274 4927 280 4928
rect 274 4923 275 4927
rect 279 4923 280 4927
rect 274 4922 280 4923
rect 111 4862 115 4863
rect 111 4857 115 4858
rect 131 4862 135 4863
rect 131 4857 135 4858
rect 112 4797 114 4857
rect 110 4796 116 4797
rect 132 4796 134 4857
rect 228 4848 230 4922
rect 276 4888 278 4922
rect 274 4887 280 4888
rect 274 4883 275 4887
rect 279 4883 280 4887
rect 274 4882 280 4883
rect 316 4863 318 4932
rect 410 4919 416 4920
rect 410 4915 411 4919
rect 415 4915 416 4919
rect 410 4914 416 4915
rect 412 4888 414 4914
rect 410 4887 416 4888
rect 410 4883 411 4887
rect 415 4883 416 4887
rect 410 4882 416 4883
rect 524 4863 526 4932
rect 608 4888 610 5030
rect 620 5028 622 5089
rect 756 5028 758 5089
rect 892 5028 894 5089
rect 1036 5028 1038 5089
rect 1130 5075 1136 5076
rect 1130 5071 1131 5075
rect 1135 5071 1136 5075
rect 1130 5070 1136 5071
rect 1132 5056 1134 5070
rect 1130 5055 1136 5056
rect 1130 5051 1131 5055
rect 1135 5051 1136 5055
rect 1130 5050 1136 5051
rect 1188 5028 1190 5089
rect 1222 5079 1228 5080
rect 1222 5075 1223 5079
rect 1227 5075 1228 5079
rect 1222 5074 1228 5075
rect 618 5027 624 5028
rect 618 5023 619 5027
rect 623 5023 624 5027
rect 618 5022 624 5023
rect 754 5027 760 5028
rect 754 5023 755 5027
rect 759 5023 760 5027
rect 754 5022 760 5023
rect 890 5027 896 5028
rect 890 5023 891 5027
rect 895 5023 896 5027
rect 890 5022 896 5023
rect 1034 5027 1040 5028
rect 1034 5023 1035 5027
rect 1039 5023 1040 5027
rect 1034 5022 1040 5023
rect 1186 5027 1192 5028
rect 1186 5023 1187 5027
rect 1191 5023 1192 5027
rect 1186 5022 1192 5023
rect 646 5012 652 5013
rect 646 5008 647 5012
rect 651 5008 652 5012
rect 646 5007 652 5008
rect 782 5012 788 5013
rect 782 5008 783 5012
rect 787 5008 788 5012
rect 782 5007 788 5008
rect 918 5012 924 5013
rect 918 5008 919 5012
rect 923 5008 924 5012
rect 918 5007 924 5008
rect 1062 5012 1068 5013
rect 1062 5008 1063 5012
rect 1067 5008 1068 5012
rect 1062 5007 1068 5008
rect 1214 5012 1220 5013
rect 1214 5008 1215 5012
rect 1219 5008 1220 5012
rect 1214 5007 1220 5008
rect 648 4983 650 5007
rect 784 4983 786 5007
rect 920 4983 922 5007
rect 1064 4983 1066 5007
rect 1216 4983 1218 5007
rect 647 4982 651 4983
rect 647 4977 651 4978
rect 751 4982 755 4983
rect 751 4977 755 4978
rect 783 4982 787 4983
rect 783 4977 787 4978
rect 919 4982 923 4983
rect 919 4977 923 4978
rect 943 4982 947 4983
rect 943 4977 947 4978
rect 1063 4982 1067 4983
rect 1063 4977 1067 4978
rect 1127 4982 1131 4983
rect 1127 4977 1131 4978
rect 1215 4982 1219 4983
rect 1215 4977 1219 4978
rect 752 4953 754 4977
rect 944 4953 946 4977
rect 1128 4953 1130 4977
rect 750 4952 756 4953
rect 750 4948 751 4952
rect 755 4948 756 4952
rect 750 4947 756 4948
rect 942 4952 948 4953
rect 942 4948 943 4952
rect 947 4948 948 4952
rect 942 4947 948 4948
rect 1126 4952 1132 4953
rect 1126 4948 1127 4952
rect 1131 4948 1132 4952
rect 1126 4947 1132 4948
rect 722 4937 728 4938
rect 722 4933 723 4937
rect 727 4933 728 4937
rect 722 4932 728 4933
rect 914 4937 920 4938
rect 914 4933 915 4937
rect 919 4933 920 4937
rect 914 4932 920 4933
rect 1098 4937 1104 4938
rect 1098 4933 1099 4937
rect 1103 4933 1104 4937
rect 1098 4932 1104 4933
rect 686 4927 692 4928
rect 686 4923 687 4927
rect 691 4923 692 4927
rect 686 4922 692 4923
rect 688 4888 690 4922
rect 606 4887 612 4888
rect 606 4883 607 4887
rect 611 4883 612 4887
rect 606 4882 612 4883
rect 686 4887 692 4888
rect 686 4883 687 4887
rect 691 4883 692 4887
rect 686 4882 692 4883
rect 724 4863 726 4932
rect 916 4863 918 4932
rect 1070 4927 1076 4928
rect 1070 4923 1071 4927
rect 1075 4923 1076 4927
rect 1070 4922 1076 4923
rect 1010 4919 1016 4920
rect 1010 4915 1011 4919
rect 1015 4915 1016 4919
rect 1010 4914 1016 4915
rect 1012 4888 1014 4914
rect 1072 4888 1074 4922
rect 1010 4887 1016 4888
rect 1010 4883 1011 4887
rect 1015 4883 1016 4887
rect 1010 4882 1016 4883
rect 1070 4887 1076 4888
rect 1070 4883 1071 4887
rect 1075 4883 1076 4887
rect 1070 4882 1076 4883
rect 1100 4863 1102 4932
rect 1224 4928 1226 5074
rect 1340 5028 1342 5089
rect 1346 5075 1352 5076
rect 1346 5071 1347 5075
rect 1351 5071 1352 5075
rect 1346 5070 1352 5071
rect 1348 5036 1350 5070
rect 1346 5035 1352 5036
rect 1346 5031 1347 5035
rect 1351 5031 1352 5035
rect 1346 5030 1352 5031
rect 1492 5028 1494 5089
rect 1586 5075 1592 5076
rect 1586 5071 1587 5075
rect 1591 5071 1592 5075
rect 1586 5070 1592 5071
rect 1588 5056 1590 5070
rect 1586 5055 1592 5056
rect 1586 5051 1587 5055
rect 1591 5051 1592 5055
rect 1586 5050 1592 5051
rect 1652 5028 1654 5089
rect 1658 5075 1664 5076
rect 1658 5071 1659 5075
rect 1663 5071 1664 5075
rect 1658 5070 1664 5071
rect 1660 5036 1662 5070
rect 1658 5035 1664 5036
rect 1658 5031 1659 5035
rect 1663 5031 1664 5035
rect 1658 5030 1664 5031
rect 1778 5035 1784 5036
rect 1778 5031 1779 5035
rect 1783 5031 1784 5035
rect 1778 5030 1784 5031
rect 1338 5027 1344 5028
rect 1338 5023 1339 5027
rect 1343 5023 1344 5027
rect 1338 5022 1344 5023
rect 1490 5027 1496 5028
rect 1490 5023 1491 5027
rect 1495 5023 1496 5027
rect 1490 5022 1496 5023
rect 1650 5027 1656 5028
rect 1650 5023 1651 5027
rect 1655 5023 1656 5027
rect 1650 5022 1656 5023
rect 1366 5012 1372 5013
rect 1366 5008 1367 5012
rect 1371 5008 1372 5012
rect 1366 5007 1372 5008
rect 1518 5012 1524 5013
rect 1518 5008 1519 5012
rect 1523 5008 1524 5012
rect 1518 5007 1524 5008
rect 1678 5012 1684 5013
rect 1678 5008 1679 5012
rect 1683 5008 1684 5012
rect 1678 5007 1684 5008
rect 1368 4983 1370 5007
rect 1520 4983 1522 5007
rect 1680 4983 1682 5007
rect 1311 4982 1315 4983
rect 1311 4977 1315 4978
rect 1367 4982 1371 4983
rect 1367 4977 1371 4978
rect 1487 4982 1491 4983
rect 1487 4977 1491 4978
rect 1519 4982 1523 4983
rect 1519 4977 1523 4978
rect 1663 4982 1667 4983
rect 1663 4977 1667 4978
rect 1679 4982 1683 4983
rect 1679 4977 1683 4978
rect 1312 4953 1314 4977
rect 1488 4953 1490 4977
rect 1664 4953 1666 4977
rect 1310 4952 1316 4953
rect 1310 4948 1311 4952
rect 1315 4948 1316 4952
rect 1310 4947 1316 4948
rect 1486 4952 1492 4953
rect 1486 4948 1487 4952
rect 1491 4948 1492 4952
rect 1486 4947 1492 4948
rect 1662 4952 1668 4953
rect 1662 4948 1663 4952
rect 1667 4948 1668 4952
rect 1662 4947 1668 4948
rect 1282 4937 1288 4938
rect 1282 4933 1283 4937
rect 1287 4933 1288 4937
rect 1282 4932 1288 4933
rect 1458 4937 1464 4938
rect 1458 4933 1459 4937
rect 1463 4933 1464 4937
rect 1458 4932 1464 4933
rect 1634 4937 1640 4938
rect 1634 4933 1635 4937
rect 1639 4933 1640 4937
rect 1634 4932 1640 4933
rect 1222 4927 1228 4928
rect 1222 4923 1223 4927
rect 1227 4923 1228 4927
rect 1222 4922 1228 4923
rect 1284 4863 1286 4932
rect 1434 4927 1440 4928
rect 1434 4923 1435 4927
rect 1439 4923 1440 4927
rect 1434 4922 1440 4923
rect 1436 4888 1438 4922
rect 1434 4887 1440 4888
rect 1434 4883 1435 4887
rect 1439 4883 1440 4887
rect 1434 4882 1440 4883
rect 1460 4863 1462 4932
rect 1610 4927 1616 4928
rect 1610 4923 1611 4927
rect 1615 4923 1616 4927
rect 1610 4922 1616 4923
rect 1612 4888 1614 4922
rect 1610 4887 1616 4888
rect 1610 4883 1611 4887
rect 1615 4883 1616 4887
rect 1610 4882 1616 4883
rect 1636 4863 1638 4932
rect 1770 4927 1776 4928
rect 1770 4923 1771 4927
rect 1775 4923 1776 4927
rect 1770 4922 1776 4923
rect 1772 4888 1774 4922
rect 1780 4888 1782 5030
rect 1788 5028 1790 5089
rect 1910 5055 1916 5056
rect 1910 5051 1911 5055
rect 1915 5051 1916 5055
rect 1910 5050 1916 5051
rect 1912 5036 1914 5050
rect 1910 5035 1916 5036
rect 1910 5031 1911 5035
rect 1915 5031 1916 5035
rect 1910 5030 1916 5031
rect 1936 5029 1938 5089
rect 1975 5085 1979 5086
rect 1995 5090 1999 5091
rect 1995 5085 1999 5086
rect 1934 5028 1940 5029
rect 1786 5027 1792 5028
rect 1786 5023 1787 5027
rect 1791 5023 1792 5027
rect 1934 5024 1935 5028
rect 1939 5024 1940 5028
rect 1976 5025 1978 5085
rect 1934 5023 1940 5024
rect 1974 5024 1980 5025
rect 1996 5024 1998 5085
rect 2092 5072 2094 5142
rect 2132 5091 2134 5152
rect 2138 5147 2144 5148
rect 2138 5143 2139 5147
rect 2143 5143 2144 5147
rect 2138 5142 2144 5143
rect 2140 5116 2142 5142
rect 2226 5139 2232 5140
rect 2226 5135 2227 5139
rect 2231 5135 2232 5139
rect 2226 5134 2232 5135
rect 2138 5115 2144 5116
rect 2138 5111 2139 5115
rect 2143 5111 2144 5115
rect 2138 5110 2144 5111
rect 2228 5108 2230 5134
rect 2226 5107 2232 5108
rect 2226 5103 2227 5107
rect 2231 5103 2232 5107
rect 2226 5102 2232 5103
rect 2300 5091 2302 5152
rect 2320 5108 2322 5250
rect 2340 5248 2342 5309
rect 2482 5299 2488 5300
rect 2482 5295 2483 5299
rect 2487 5295 2488 5299
rect 2482 5294 2488 5295
rect 2484 5256 2486 5294
rect 2482 5255 2488 5256
rect 2482 5251 2483 5255
rect 2487 5251 2488 5255
rect 2482 5250 2488 5251
rect 2492 5248 2494 5309
rect 2652 5248 2654 5309
rect 2812 5300 2814 5366
rect 2860 5315 2862 5376
rect 2986 5371 2992 5372
rect 2986 5367 2987 5371
rect 2991 5367 2992 5371
rect 2986 5366 2992 5367
rect 2988 5332 2990 5366
rect 2954 5331 2960 5332
rect 2954 5327 2955 5331
rect 2959 5327 2960 5331
rect 2954 5326 2960 5327
rect 2986 5331 2992 5332
rect 2986 5327 2987 5331
rect 2991 5327 2992 5331
rect 2986 5326 2992 5327
rect 2819 5314 2823 5315
rect 2819 5309 2823 5310
rect 2859 5314 2863 5315
rect 2859 5309 2863 5310
rect 2802 5299 2808 5300
rect 2802 5295 2803 5299
rect 2807 5295 2808 5299
rect 2802 5294 2808 5295
rect 2810 5299 2816 5300
rect 2810 5295 2811 5299
rect 2815 5295 2816 5299
rect 2810 5294 2816 5295
rect 2804 5256 2806 5294
rect 2802 5255 2808 5256
rect 2802 5251 2803 5255
rect 2807 5251 2808 5255
rect 2802 5250 2808 5251
rect 2820 5248 2822 5309
rect 2956 5256 2958 5326
rect 3044 5315 3046 5376
rect 3168 5372 3170 5526
rect 3292 5480 3294 5541
rect 3326 5487 3332 5488
rect 3326 5483 3327 5487
rect 3331 5483 3332 5487
rect 3326 5482 3332 5483
rect 3290 5479 3296 5480
rect 3290 5475 3291 5479
rect 3295 5475 3296 5479
rect 3290 5474 3296 5475
rect 3318 5464 3324 5465
rect 3318 5460 3319 5464
rect 3323 5460 3324 5464
rect 3318 5459 3324 5460
rect 3320 5427 3322 5459
rect 3247 5426 3251 5427
rect 3247 5421 3251 5422
rect 3319 5426 3323 5427
rect 3319 5421 3323 5422
rect 3248 5397 3250 5421
rect 3246 5396 3252 5397
rect 3246 5392 3247 5396
rect 3251 5392 3252 5396
rect 3246 5391 3252 5392
rect 3218 5381 3224 5382
rect 3218 5377 3219 5381
rect 3223 5377 3224 5381
rect 3218 5376 3224 5377
rect 3166 5371 3172 5372
rect 3166 5367 3167 5371
rect 3171 5367 3172 5371
rect 3166 5366 3172 5367
rect 3220 5315 3222 5376
rect 3328 5332 3330 5482
rect 3468 5480 3470 5541
rect 3634 5531 3640 5532
rect 3634 5527 3635 5531
rect 3639 5527 3640 5531
rect 3634 5526 3640 5527
rect 3636 5488 3638 5526
rect 3634 5487 3640 5488
rect 3634 5483 3635 5487
rect 3639 5483 3640 5487
rect 3634 5482 3640 5483
rect 3644 5480 3646 5541
rect 3740 5532 3742 5598
rect 3800 5547 3802 5607
rect 3838 5604 3839 5608
rect 3843 5604 3844 5608
rect 4306 5605 4307 5609
rect 4311 5605 4312 5609
rect 4306 5604 4312 5605
rect 4442 5609 4448 5610
rect 4442 5605 4443 5609
rect 4447 5605 4448 5609
rect 4442 5604 4448 5605
rect 4578 5609 4584 5610
rect 4578 5605 4579 5609
rect 4583 5605 4584 5609
rect 4578 5604 4584 5605
rect 4714 5609 4720 5610
rect 4714 5605 4715 5609
rect 4719 5605 4720 5609
rect 4714 5604 4720 5605
rect 4850 5609 4856 5610
rect 4850 5605 4851 5609
rect 4855 5605 4856 5609
rect 4850 5604 4856 5605
rect 4986 5609 4992 5610
rect 4986 5605 4987 5609
rect 4991 5605 4992 5609
rect 4986 5604 4992 5605
rect 5662 5608 5668 5609
rect 5662 5604 5663 5608
rect 5667 5604 5668 5608
rect 3838 5603 3844 5604
rect 3799 5546 3803 5547
rect 3840 5543 3842 5603
rect 4308 5543 4310 5604
rect 4434 5599 4440 5600
rect 4434 5595 4435 5599
rect 4439 5595 4440 5599
rect 4434 5594 4440 5595
rect 4436 5560 4438 5594
rect 4374 5559 4380 5560
rect 4374 5555 4375 5559
rect 4379 5555 4380 5559
rect 4374 5554 4380 5555
rect 4434 5559 4440 5560
rect 4434 5555 4435 5559
rect 4439 5555 4440 5559
rect 4434 5554 4440 5555
rect 3799 5541 3803 5542
rect 3839 5542 3843 5543
rect 3738 5531 3744 5532
rect 3738 5527 3739 5531
rect 3743 5527 3744 5531
rect 3738 5526 3744 5527
rect 3800 5481 3802 5541
rect 3839 5537 3843 5538
rect 4251 5542 4255 5543
rect 4251 5537 4255 5538
rect 4307 5542 4311 5543
rect 4307 5537 4311 5538
rect 3798 5480 3804 5481
rect 3466 5479 3472 5480
rect 3466 5475 3467 5479
rect 3471 5475 3472 5479
rect 3466 5474 3472 5475
rect 3642 5479 3648 5480
rect 3642 5475 3643 5479
rect 3647 5475 3648 5479
rect 3798 5476 3799 5480
rect 3803 5476 3804 5480
rect 3840 5477 3842 5537
rect 3798 5475 3804 5476
rect 3838 5476 3844 5477
rect 4252 5476 4254 5537
rect 4376 5484 4378 5554
rect 4444 5543 4446 5604
rect 4570 5599 4576 5600
rect 4570 5595 4571 5599
rect 4575 5595 4576 5599
rect 4570 5594 4576 5595
rect 4572 5560 4574 5594
rect 4570 5559 4576 5560
rect 4570 5555 4571 5559
rect 4575 5555 4576 5559
rect 4570 5554 4576 5555
rect 4580 5543 4582 5604
rect 4706 5599 4712 5600
rect 4706 5595 4707 5599
rect 4711 5595 4712 5599
rect 4706 5594 4712 5595
rect 4708 5560 4710 5594
rect 4706 5559 4712 5560
rect 4706 5555 4707 5559
rect 4711 5555 4712 5559
rect 4706 5554 4712 5555
rect 4716 5543 4718 5604
rect 4842 5599 4848 5600
rect 4842 5595 4843 5599
rect 4847 5595 4848 5599
rect 4842 5594 4848 5595
rect 4844 5560 4846 5594
rect 4842 5559 4848 5560
rect 4842 5555 4843 5559
rect 4847 5555 4848 5559
rect 4842 5554 4848 5555
rect 4852 5543 4854 5604
rect 4978 5599 4984 5600
rect 4978 5595 4979 5599
rect 4983 5595 4984 5599
rect 4978 5594 4984 5595
rect 4980 5560 4982 5594
rect 4978 5559 4984 5560
rect 4978 5555 4979 5559
rect 4983 5555 4984 5559
rect 4978 5554 4984 5555
rect 4988 5543 4990 5604
rect 5662 5603 5668 5604
rect 5110 5599 5116 5600
rect 5110 5595 5111 5599
rect 5115 5595 5116 5599
rect 5110 5594 5116 5595
rect 4403 5542 4407 5543
rect 4403 5537 4407 5538
rect 4443 5542 4447 5543
rect 4443 5537 4447 5538
rect 4555 5542 4559 5543
rect 4555 5537 4559 5538
rect 4579 5542 4583 5543
rect 4579 5537 4583 5538
rect 4707 5542 4711 5543
rect 4707 5537 4711 5538
rect 4715 5542 4719 5543
rect 4715 5537 4719 5538
rect 4851 5542 4855 5543
rect 4851 5537 4855 5538
rect 4859 5542 4863 5543
rect 4859 5537 4863 5538
rect 4987 5542 4991 5543
rect 4987 5537 4991 5538
rect 5019 5542 5023 5543
rect 5019 5537 5023 5538
rect 4374 5483 4380 5484
rect 4374 5479 4375 5483
rect 4379 5479 4380 5483
rect 4374 5478 4380 5479
rect 4404 5476 4406 5537
rect 4556 5476 4558 5537
rect 4574 5527 4580 5528
rect 4574 5523 4575 5527
rect 4579 5523 4580 5527
rect 4574 5522 4580 5523
rect 3642 5474 3648 5475
rect 3838 5472 3839 5476
rect 3843 5472 3844 5476
rect 3838 5471 3844 5472
rect 4250 5475 4256 5476
rect 4250 5471 4251 5475
rect 4255 5471 4256 5475
rect 4250 5470 4256 5471
rect 4402 5475 4408 5476
rect 4402 5471 4403 5475
rect 4407 5471 4408 5475
rect 4402 5470 4408 5471
rect 4554 5475 4560 5476
rect 4554 5471 4555 5475
rect 4559 5471 4560 5475
rect 4554 5470 4560 5471
rect 3494 5464 3500 5465
rect 3494 5460 3495 5464
rect 3499 5460 3500 5464
rect 3494 5459 3500 5460
rect 3670 5464 3676 5465
rect 3670 5460 3671 5464
rect 3675 5460 3676 5464
rect 3670 5459 3676 5460
rect 3798 5463 3804 5464
rect 3798 5459 3799 5463
rect 3803 5459 3804 5463
rect 4278 5460 4284 5461
rect 3496 5427 3498 5459
rect 3672 5427 3674 5459
rect 3798 5458 3804 5459
rect 3838 5459 3844 5460
rect 3800 5427 3802 5458
rect 3838 5455 3839 5459
rect 3843 5455 3844 5459
rect 4278 5456 4279 5460
rect 4283 5456 4284 5460
rect 4278 5455 4284 5456
rect 4430 5460 4436 5461
rect 4430 5456 4431 5460
rect 4435 5456 4436 5460
rect 4430 5455 4436 5456
rect 3838 5454 3844 5455
rect 3423 5426 3427 5427
rect 3423 5421 3427 5422
rect 3495 5426 3499 5427
rect 3495 5421 3499 5422
rect 3607 5426 3611 5427
rect 3607 5421 3611 5422
rect 3671 5426 3675 5427
rect 3671 5421 3675 5422
rect 3799 5426 3803 5427
rect 3799 5421 3803 5422
rect 3424 5397 3426 5421
rect 3608 5397 3610 5421
rect 3800 5398 3802 5421
rect 3840 5411 3842 5454
rect 4280 5411 4282 5455
rect 4432 5411 4434 5455
rect 3839 5410 3843 5411
rect 3839 5405 3843 5406
rect 4279 5410 4283 5411
rect 4279 5405 4283 5406
rect 4431 5410 4435 5411
rect 4431 5405 4435 5406
rect 4487 5410 4491 5411
rect 4487 5405 4491 5406
rect 3798 5397 3804 5398
rect 3422 5396 3428 5397
rect 3422 5392 3423 5396
rect 3427 5392 3428 5396
rect 3422 5391 3428 5392
rect 3606 5396 3612 5397
rect 3606 5392 3607 5396
rect 3611 5392 3612 5396
rect 3798 5393 3799 5397
rect 3803 5393 3804 5397
rect 3798 5392 3804 5393
rect 3606 5391 3612 5392
rect 3840 5382 3842 5405
rect 3394 5381 3400 5382
rect 3394 5377 3395 5381
rect 3399 5377 3400 5381
rect 3394 5376 3400 5377
rect 3578 5381 3584 5382
rect 3838 5381 3844 5382
rect 4280 5381 4282 5405
rect 4488 5381 4490 5405
rect 3578 5377 3579 5381
rect 3583 5377 3584 5381
rect 3578 5376 3584 5377
rect 3798 5380 3804 5381
rect 3798 5376 3799 5380
rect 3803 5376 3804 5380
rect 3838 5377 3839 5381
rect 3843 5377 3844 5381
rect 3838 5376 3844 5377
rect 4278 5380 4284 5381
rect 4278 5376 4279 5380
rect 4283 5376 4284 5380
rect 3346 5371 3352 5372
rect 3346 5367 3347 5371
rect 3351 5367 3352 5371
rect 3346 5366 3352 5367
rect 3348 5332 3350 5366
rect 3326 5331 3332 5332
rect 3326 5327 3327 5331
rect 3331 5327 3332 5331
rect 3326 5326 3332 5327
rect 3346 5331 3352 5332
rect 3346 5327 3347 5331
rect 3351 5327 3352 5331
rect 3346 5326 3352 5327
rect 3396 5315 3398 5376
rect 3522 5371 3528 5372
rect 3522 5367 3523 5371
rect 3527 5367 3528 5371
rect 3522 5366 3528 5367
rect 3524 5332 3526 5366
rect 3522 5331 3528 5332
rect 3522 5327 3523 5331
rect 3527 5327 3528 5331
rect 3522 5326 3528 5327
rect 3580 5315 3582 5376
rect 3798 5375 3804 5376
rect 4278 5375 4284 5376
rect 4486 5380 4492 5381
rect 4486 5376 4487 5380
rect 4491 5376 4492 5380
rect 4486 5375 4492 5376
rect 3674 5371 3680 5372
rect 3674 5367 3675 5371
rect 3679 5367 3680 5371
rect 3674 5366 3680 5367
rect 3003 5314 3007 5315
rect 3003 5309 3007 5310
rect 3043 5314 3047 5315
rect 3043 5309 3047 5310
rect 3187 5314 3191 5315
rect 3187 5309 3191 5310
rect 3219 5314 3223 5315
rect 3219 5309 3223 5310
rect 3379 5314 3383 5315
rect 3379 5309 3383 5310
rect 3395 5314 3399 5315
rect 3395 5309 3399 5310
rect 3579 5314 3583 5315
rect 3579 5309 3583 5310
rect 2954 5255 2960 5256
rect 2954 5251 2955 5255
rect 2959 5251 2960 5255
rect 2954 5250 2960 5251
rect 3004 5248 3006 5309
rect 3188 5248 3190 5309
rect 3194 5295 3200 5296
rect 3194 5291 3195 5295
rect 3199 5291 3200 5295
rect 3194 5290 3200 5291
rect 2338 5247 2344 5248
rect 2338 5243 2339 5247
rect 2343 5243 2344 5247
rect 2338 5242 2344 5243
rect 2490 5247 2496 5248
rect 2490 5243 2491 5247
rect 2495 5243 2496 5247
rect 2490 5242 2496 5243
rect 2650 5247 2656 5248
rect 2650 5243 2651 5247
rect 2655 5243 2656 5247
rect 2650 5242 2656 5243
rect 2818 5247 2824 5248
rect 2818 5243 2819 5247
rect 2823 5243 2824 5247
rect 2818 5242 2824 5243
rect 3002 5247 3008 5248
rect 3002 5243 3003 5247
rect 3007 5243 3008 5247
rect 3002 5242 3008 5243
rect 3186 5247 3192 5248
rect 3186 5243 3187 5247
rect 3191 5243 3192 5247
rect 3186 5242 3192 5243
rect 2366 5232 2372 5233
rect 2366 5228 2367 5232
rect 2371 5228 2372 5232
rect 2366 5227 2372 5228
rect 2518 5232 2524 5233
rect 2518 5228 2519 5232
rect 2523 5228 2524 5232
rect 2518 5227 2524 5228
rect 2678 5232 2684 5233
rect 2678 5228 2679 5232
rect 2683 5228 2684 5232
rect 2678 5227 2684 5228
rect 2846 5232 2852 5233
rect 2846 5228 2847 5232
rect 2851 5228 2852 5232
rect 2846 5227 2852 5228
rect 3030 5232 3036 5233
rect 3030 5228 3031 5232
rect 3035 5228 3036 5232
rect 3030 5227 3036 5228
rect 2368 5203 2370 5227
rect 2520 5203 2522 5227
rect 2680 5203 2682 5227
rect 2848 5203 2850 5227
rect 3032 5203 3034 5227
rect 2327 5202 2331 5203
rect 2327 5197 2331 5198
rect 2367 5202 2371 5203
rect 2367 5197 2371 5198
rect 2511 5202 2515 5203
rect 2511 5197 2515 5198
rect 2519 5202 2523 5203
rect 2519 5197 2523 5198
rect 2679 5202 2683 5203
rect 2679 5197 2683 5198
rect 2695 5202 2699 5203
rect 2695 5197 2699 5198
rect 2847 5202 2851 5203
rect 2847 5197 2851 5198
rect 2887 5202 2891 5203
rect 2887 5197 2891 5198
rect 3031 5202 3035 5203
rect 3031 5197 3035 5198
rect 3087 5202 3091 5203
rect 3087 5197 3091 5198
rect 2328 5173 2330 5197
rect 2512 5173 2514 5197
rect 2696 5173 2698 5197
rect 2888 5173 2890 5197
rect 3088 5173 3090 5197
rect 2326 5172 2332 5173
rect 2326 5168 2327 5172
rect 2331 5168 2332 5172
rect 2326 5167 2332 5168
rect 2510 5172 2516 5173
rect 2510 5168 2511 5172
rect 2515 5168 2516 5172
rect 2510 5167 2516 5168
rect 2694 5172 2700 5173
rect 2694 5168 2695 5172
rect 2699 5168 2700 5172
rect 2694 5167 2700 5168
rect 2886 5172 2892 5173
rect 2886 5168 2887 5172
rect 2891 5168 2892 5172
rect 2886 5167 2892 5168
rect 3086 5172 3092 5173
rect 3086 5168 3087 5172
rect 3091 5168 3092 5172
rect 3086 5167 3092 5168
rect 2482 5157 2488 5158
rect 2482 5153 2483 5157
rect 2487 5153 2488 5157
rect 2482 5152 2488 5153
rect 2666 5157 2672 5158
rect 2666 5153 2667 5157
rect 2671 5153 2672 5157
rect 2666 5152 2672 5153
rect 2858 5157 2864 5158
rect 2858 5153 2859 5157
rect 2863 5153 2864 5157
rect 2858 5152 2864 5153
rect 3058 5157 3064 5158
rect 3058 5153 3059 5157
rect 3063 5153 3064 5157
rect 3058 5152 3064 5153
rect 2426 5147 2432 5148
rect 2426 5143 2427 5147
rect 2431 5143 2432 5147
rect 2426 5142 2432 5143
rect 2428 5108 2430 5142
rect 2318 5107 2324 5108
rect 2318 5103 2319 5107
rect 2323 5103 2324 5107
rect 2318 5102 2324 5103
rect 2426 5107 2432 5108
rect 2426 5103 2427 5107
rect 2431 5103 2432 5107
rect 2426 5102 2432 5103
rect 2484 5091 2486 5152
rect 2610 5147 2616 5148
rect 2610 5143 2611 5147
rect 2615 5143 2616 5147
rect 2610 5142 2616 5143
rect 2612 5108 2614 5142
rect 2610 5107 2616 5108
rect 2610 5103 2611 5107
rect 2615 5103 2616 5107
rect 2610 5102 2616 5103
rect 2668 5091 2670 5152
rect 2860 5091 2862 5152
rect 2998 5147 3004 5148
rect 2998 5143 2999 5147
rect 3003 5143 3004 5147
rect 2998 5142 3004 5143
rect 3000 5108 3002 5142
rect 2998 5107 3004 5108
rect 2998 5103 2999 5107
rect 3003 5103 3004 5107
rect 2998 5102 3004 5103
rect 3060 5091 3062 5152
rect 3196 5148 3198 5290
rect 3354 5255 3360 5256
rect 3354 5251 3355 5255
rect 3359 5251 3360 5255
rect 3354 5250 3360 5251
rect 3214 5232 3220 5233
rect 3214 5228 3215 5232
rect 3219 5228 3220 5232
rect 3214 5227 3220 5228
rect 3216 5203 3218 5227
rect 3215 5202 3219 5203
rect 3215 5197 3219 5198
rect 3287 5202 3291 5203
rect 3287 5197 3291 5198
rect 3288 5173 3290 5197
rect 3286 5172 3292 5173
rect 3286 5168 3287 5172
rect 3291 5168 3292 5172
rect 3286 5167 3292 5168
rect 3258 5157 3264 5158
rect 3258 5153 3259 5157
rect 3263 5153 3264 5157
rect 3258 5152 3264 5153
rect 3194 5147 3200 5148
rect 3194 5143 3195 5147
rect 3199 5143 3200 5147
rect 3194 5142 3200 5143
rect 3260 5091 3262 5152
rect 3356 5108 3358 5250
rect 3380 5248 3382 5309
rect 3580 5248 3582 5309
rect 3676 5300 3678 5366
rect 3800 5315 3802 5375
rect 4250 5365 4256 5366
rect 3838 5364 3844 5365
rect 3838 5360 3839 5364
rect 3843 5360 3844 5364
rect 4250 5361 4251 5365
rect 4255 5361 4256 5365
rect 4250 5360 4256 5361
rect 4458 5365 4464 5366
rect 4458 5361 4459 5365
rect 4463 5361 4464 5365
rect 4458 5360 4464 5361
rect 3838 5359 3844 5360
rect 3799 5314 3803 5315
rect 3799 5309 3803 5310
rect 3674 5299 3680 5300
rect 3674 5295 3675 5299
rect 3679 5295 3680 5299
rect 3674 5294 3680 5295
rect 3800 5249 3802 5309
rect 3840 5283 3842 5359
rect 4252 5283 4254 5360
rect 4418 5355 4424 5356
rect 4418 5351 4419 5355
rect 4423 5351 4424 5355
rect 4418 5350 4424 5351
rect 4420 5316 4422 5350
rect 4346 5315 4352 5316
rect 4346 5311 4347 5315
rect 4351 5311 4352 5315
rect 4346 5310 4352 5311
rect 4418 5315 4424 5316
rect 4418 5311 4419 5315
rect 4423 5311 4424 5315
rect 4418 5310 4424 5311
rect 3839 5282 3843 5283
rect 3839 5277 3843 5278
rect 4251 5282 4255 5283
rect 4251 5277 4255 5278
rect 3798 5248 3804 5249
rect 3378 5247 3384 5248
rect 3378 5243 3379 5247
rect 3383 5243 3384 5247
rect 3378 5242 3384 5243
rect 3578 5247 3584 5248
rect 3578 5243 3579 5247
rect 3583 5243 3584 5247
rect 3798 5244 3799 5248
rect 3803 5244 3804 5248
rect 3798 5243 3804 5244
rect 3578 5242 3584 5243
rect 3406 5232 3412 5233
rect 3406 5228 3407 5232
rect 3411 5228 3412 5232
rect 3406 5227 3412 5228
rect 3606 5232 3612 5233
rect 3606 5228 3607 5232
rect 3611 5228 3612 5232
rect 3606 5227 3612 5228
rect 3798 5231 3804 5232
rect 3798 5227 3799 5231
rect 3803 5227 3804 5231
rect 3408 5203 3410 5227
rect 3608 5203 3610 5227
rect 3798 5226 3804 5227
rect 3800 5203 3802 5226
rect 3840 5217 3842 5277
rect 3838 5216 3844 5217
rect 4252 5216 4254 5277
rect 4348 5224 4350 5310
rect 4460 5283 4462 5360
rect 4576 5356 4578 5522
rect 4708 5476 4710 5537
rect 4850 5527 4856 5528
rect 4850 5523 4851 5527
rect 4855 5523 4856 5527
rect 4850 5522 4856 5523
rect 4852 5484 4854 5522
rect 4762 5483 4768 5484
rect 4762 5479 4763 5483
rect 4767 5479 4768 5483
rect 4762 5478 4768 5479
rect 4850 5483 4856 5484
rect 4850 5479 4851 5483
rect 4855 5479 4856 5483
rect 4850 5478 4856 5479
rect 4706 5475 4712 5476
rect 4706 5471 4707 5475
rect 4711 5471 4712 5475
rect 4706 5470 4712 5471
rect 4582 5460 4588 5461
rect 4582 5456 4583 5460
rect 4587 5456 4588 5460
rect 4582 5455 4588 5456
rect 4734 5460 4740 5461
rect 4734 5456 4735 5460
rect 4739 5456 4740 5460
rect 4734 5455 4740 5456
rect 4584 5411 4586 5455
rect 4736 5411 4738 5455
rect 4583 5410 4587 5411
rect 4583 5405 4587 5406
rect 4695 5410 4699 5411
rect 4695 5405 4699 5406
rect 4735 5410 4739 5411
rect 4735 5405 4739 5406
rect 4696 5381 4698 5405
rect 4694 5380 4700 5381
rect 4694 5376 4695 5380
rect 4699 5376 4700 5380
rect 4694 5375 4700 5376
rect 4666 5365 4672 5366
rect 4666 5361 4667 5365
rect 4671 5361 4672 5365
rect 4666 5360 4672 5361
rect 4574 5355 4580 5356
rect 4574 5351 4575 5355
rect 4579 5351 4580 5355
rect 4574 5350 4580 5351
rect 4668 5283 4670 5360
rect 4764 5316 4766 5478
rect 4860 5476 4862 5537
rect 5020 5476 5022 5537
rect 5112 5528 5114 5594
rect 5664 5543 5666 5603
rect 5663 5542 5667 5543
rect 5663 5537 5667 5538
rect 5110 5527 5116 5528
rect 5110 5523 5111 5527
rect 5115 5523 5116 5527
rect 5110 5522 5116 5523
rect 5664 5477 5666 5537
rect 5662 5476 5668 5477
rect 4858 5475 4864 5476
rect 4858 5471 4859 5475
rect 4863 5471 4864 5475
rect 4858 5470 4864 5471
rect 5018 5475 5024 5476
rect 5018 5471 5019 5475
rect 5023 5471 5024 5475
rect 5662 5472 5663 5476
rect 5667 5472 5668 5476
rect 5662 5471 5668 5472
rect 5018 5470 5024 5471
rect 4886 5460 4892 5461
rect 4886 5456 4887 5460
rect 4891 5456 4892 5460
rect 4886 5455 4892 5456
rect 5046 5460 5052 5461
rect 5046 5456 5047 5460
rect 5051 5456 5052 5460
rect 5046 5455 5052 5456
rect 5662 5459 5668 5460
rect 5662 5455 5663 5459
rect 5667 5455 5668 5459
rect 4888 5411 4890 5455
rect 5048 5411 5050 5455
rect 5662 5454 5668 5455
rect 5664 5411 5666 5454
rect 4887 5410 4891 5411
rect 4887 5405 4891 5406
rect 4911 5410 4915 5411
rect 4911 5405 4915 5406
rect 5047 5410 5051 5411
rect 5047 5405 5051 5406
rect 5127 5410 5131 5411
rect 5127 5405 5131 5406
rect 5663 5410 5667 5411
rect 5663 5405 5667 5406
rect 4912 5381 4914 5405
rect 5128 5381 5130 5405
rect 5664 5382 5666 5405
rect 5662 5381 5668 5382
rect 4910 5380 4916 5381
rect 4910 5376 4911 5380
rect 4915 5376 4916 5380
rect 4910 5375 4916 5376
rect 5126 5380 5132 5381
rect 5126 5376 5127 5380
rect 5131 5376 5132 5380
rect 5662 5377 5663 5381
rect 5667 5377 5668 5381
rect 5662 5376 5668 5377
rect 5126 5375 5132 5376
rect 4882 5365 4888 5366
rect 4882 5361 4883 5365
rect 4887 5361 4888 5365
rect 4882 5360 4888 5361
rect 5098 5365 5104 5366
rect 5098 5361 5099 5365
rect 5103 5361 5104 5365
rect 5098 5360 5104 5361
rect 5662 5364 5668 5365
rect 5662 5360 5663 5364
rect 5667 5360 5668 5364
rect 4806 5355 4812 5356
rect 4806 5351 4807 5355
rect 4811 5351 4812 5355
rect 4806 5350 4812 5351
rect 4808 5316 4810 5350
rect 4762 5315 4768 5316
rect 4762 5311 4763 5315
rect 4767 5311 4768 5315
rect 4762 5310 4768 5311
rect 4806 5315 4812 5316
rect 4806 5311 4807 5315
rect 4811 5311 4812 5315
rect 4806 5310 4812 5311
rect 4884 5283 4886 5360
rect 5010 5355 5016 5356
rect 5010 5351 5011 5355
rect 5015 5351 5016 5355
rect 5010 5350 5016 5351
rect 5012 5316 5014 5350
rect 5010 5315 5016 5316
rect 5010 5311 5011 5315
rect 5015 5311 5016 5315
rect 5010 5310 5016 5311
rect 5100 5283 5102 5360
rect 5662 5359 5668 5360
rect 5222 5355 5228 5356
rect 5222 5351 5223 5355
rect 5227 5351 5228 5355
rect 5222 5350 5228 5351
rect 4459 5282 4463 5283
rect 4459 5277 4463 5278
rect 4483 5282 4487 5283
rect 4483 5277 4487 5278
rect 4667 5282 4671 5283
rect 4667 5277 4671 5278
rect 4715 5282 4719 5283
rect 4715 5277 4719 5278
rect 4883 5282 4887 5283
rect 4883 5277 4887 5278
rect 4947 5282 4951 5283
rect 4947 5277 4951 5278
rect 5099 5282 5103 5283
rect 5099 5277 5103 5278
rect 5187 5282 5191 5283
rect 5187 5277 5191 5278
rect 4346 5223 4352 5224
rect 4346 5219 4347 5223
rect 4351 5219 4352 5223
rect 4346 5218 4352 5219
rect 4484 5216 4486 5277
rect 4502 5267 4508 5268
rect 4502 5263 4503 5267
rect 4507 5263 4508 5267
rect 4502 5262 4508 5263
rect 3838 5212 3839 5216
rect 3843 5212 3844 5216
rect 3838 5211 3844 5212
rect 4250 5215 4256 5216
rect 4250 5211 4251 5215
rect 4255 5211 4256 5215
rect 4250 5210 4256 5211
rect 4482 5215 4488 5216
rect 4482 5211 4483 5215
rect 4487 5211 4488 5215
rect 4482 5210 4488 5211
rect 3407 5202 3411 5203
rect 3407 5197 3411 5198
rect 3495 5202 3499 5203
rect 3495 5197 3499 5198
rect 3607 5202 3611 5203
rect 3607 5197 3611 5198
rect 3679 5202 3683 5203
rect 3679 5197 3683 5198
rect 3799 5202 3803 5203
rect 4278 5200 4284 5201
rect 3799 5197 3803 5198
rect 3838 5199 3844 5200
rect 3496 5173 3498 5197
rect 3680 5173 3682 5197
rect 3800 5174 3802 5197
rect 3838 5195 3839 5199
rect 3843 5195 3844 5199
rect 4278 5196 4279 5200
rect 4283 5196 4284 5200
rect 4278 5195 4284 5196
rect 3838 5194 3844 5195
rect 3798 5173 3804 5174
rect 3494 5172 3500 5173
rect 3494 5168 3495 5172
rect 3499 5168 3500 5172
rect 3494 5167 3500 5168
rect 3678 5172 3684 5173
rect 3678 5168 3679 5172
rect 3683 5168 3684 5172
rect 3798 5169 3799 5173
rect 3803 5169 3804 5173
rect 3798 5168 3804 5169
rect 3678 5167 3684 5168
rect 3466 5157 3472 5158
rect 3466 5153 3467 5157
rect 3471 5153 3472 5157
rect 3466 5152 3472 5153
rect 3650 5157 3656 5158
rect 3650 5153 3651 5157
rect 3655 5153 3656 5157
rect 3650 5152 3656 5153
rect 3798 5156 3804 5157
rect 3798 5152 3799 5156
rect 3803 5152 3804 5156
rect 3426 5147 3432 5148
rect 3426 5143 3427 5147
rect 3431 5143 3432 5147
rect 3426 5142 3432 5143
rect 3428 5108 3430 5142
rect 3354 5107 3360 5108
rect 3354 5103 3355 5107
rect 3359 5103 3360 5107
rect 3354 5102 3360 5103
rect 3426 5107 3432 5108
rect 3426 5103 3427 5107
rect 3431 5103 3432 5107
rect 3426 5102 3432 5103
rect 3468 5091 3470 5152
rect 3606 5147 3612 5148
rect 3606 5143 3607 5147
rect 3611 5143 3612 5147
rect 3606 5142 3612 5143
rect 3608 5108 3610 5142
rect 3606 5107 3612 5108
rect 3606 5103 3607 5107
rect 3611 5103 3612 5107
rect 3606 5102 3612 5103
rect 3652 5091 3654 5152
rect 3798 5151 3804 5152
rect 3746 5147 3752 5148
rect 3746 5143 3747 5147
rect 3751 5143 3752 5147
rect 3746 5142 3752 5143
rect 2131 5090 2135 5091
rect 2131 5085 2135 5086
rect 2299 5090 2303 5091
rect 2299 5085 2303 5086
rect 2483 5090 2487 5091
rect 2483 5085 2487 5086
rect 2531 5090 2535 5091
rect 2531 5085 2535 5086
rect 2667 5090 2671 5091
rect 2667 5085 2671 5086
rect 2859 5090 2863 5091
rect 2859 5085 2863 5086
rect 3059 5090 3063 5091
rect 3059 5085 3063 5086
rect 3099 5090 3103 5091
rect 3099 5085 3103 5086
rect 3259 5090 3263 5091
rect 3259 5085 3263 5086
rect 3467 5090 3471 5091
rect 3467 5085 3471 5086
rect 3651 5090 3655 5091
rect 3651 5085 3655 5086
rect 2118 5079 2124 5080
rect 2118 5075 2119 5079
rect 2123 5075 2124 5079
rect 2118 5074 2124 5075
rect 2090 5071 2096 5072
rect 2090 5067 2091 5071
rect 2095 5067 2096 5071
rect 2090 5066 2096 5067
rect 2120 5032 2122 5074
rect 2118 5031 2124 5032
rect 2118 5027 2119 5031
rect 2123 5027 2124 5031
rect 2118 5026 2124 5027
rect 2532 5024 2534 5085
rect 2954 5075 2960 5076
rect 2954 5071 2955 5075
rect 2959 5071 2960 5075
rect 2954 5070 2960 5071
rect 3018 5075 3024 5076
rect 3018 5071 3019 5075
rect 3023 5071 3024 5075
rect 3018 5070 3024 5071
rect 2956 5032 2958 5070
rect 2954 5031 2960 5032
rect 2954 5027 2955 5031
rect 2959 5027 2960 5031
rect 2954 5026 2960 5027
rect 1786 5022 1792 5023
rect 1974 5020 1975 5024
rect 1979 5020 1980 5024
rect 1974 5019 1980 5020
rect 1994 5023 2000 5024
rect 1994 5019 1995 5023
rect 1999 5019 2000 5023
rect 1994 5018 2000 5019
rect 2530 5023 2536 5024
rect 2530 5019 2531 5023
rect 2535 5019 2536 5023
rect 2530 5018 2536 5019
rect 1814 5012 1820 5013
rect 1814 5008 1815 5012
rect 1819 5008 1820 5012
rect 1814 5007 1820 5008
rect 1934 5011 1940 5012
rect 1934 5007 1935 5011
rect 1939 5007 1940 5011
rect 2022 5008 2028 5009
rect 1816 4983 1818 5007
rect 1934 5006 1940 5007
rect 1974 5007 1980 5008
rect 1936 4983 1938 5006
rect 1974 5003 1975 5007
rect 1979 5003 1980 5007
rect 2022 5004 2023 5008
rect 2027 5004 2028 5008
rect 2022 5003 2028 5004
rect 2558 5008 2564 5009
rect 2558 5004 2559 5008
rect 2563 5004 2564 5008
rect 2558 5003 2564 5004
rect 1974 5002 1980 5003
rect 1815 4982 1819 4983
rect 1815 4977 1819 4978
rect 1935 4982 1939 4983
rect 1935 4977 1939 4978
rect 1816 4953 1818 4977
rect 1936 4954 1938 4977
rect 1934 4953 1940 4954
rect 1814 4952 1820 4953
rect 1814 4948 1815 4952
rect 1819 4948 1820 4952
rect 1934 4949 1935 4953
rect 1939 4949 1940 4953
rect 1934 4948 1940 4949
rect 1814 4947 1820 4948
rect 1976 4947 1978 5002
rect 2024 4947 2026 5003
rect 2560 4947 2562 5003
rect 1975 4946 1979 4947
rect 1975 4941 1979 4942
rect 2023 4946 2027 4947
rect 2023 4941 2027 4942
rect 2559 4946 2563 4947
rect 2559 4941 2563 4942
rect 2871 4946 2875 4947
rect 2871 4941 2875 4942
rect 3007 4946 3011 4947
rect 3007 4941 3011 4942
rect 1786 4937 1792 4938
rect 1786 4933 1787 4937
rect 1791 4933 1792 4937
rect 1786 4932 1792 4933
rect 1934 4936 1940 4937
rect 1934 4932 1935 4936
rect 1939 4932 1940 4936
rect 1770 4887 1776 4888
rect 1770 4883 1771 4887
rect 1775 4883 1776 4887
rect 1770 4882 1776 4883
rect 1778 4887 1784 4888
rect 1778 4883 1779 4887
rect 1783 4883 1784 4887
rect 1778 4882 1784 4883
rect 1788 4863 1790 4932
rect 1934 4931 1940 4932
rect 1936 4863 1938 4931
rect 1976 4918 1978 4941
rect 1974 4917 1980 4918
rect 2872 4917 2874 4941
rect 3008 4917 3010 4941
rect 1974 4913 1975 4917
rect 1979 4913 1980 4917
rect 1974 4912 1980 4913
rect 2870 4916 2876 4917
rect 2870 4912 2871 4916
rect 2875 4912 2876 4916
rect 2870 4911 2876 4912
rect 3006 4916 3012 4917
rect 3006 4912 3007 4916
rect 3011 4912 3012 4916
rect 3006 4911 3012 4912
rect 2842 4901 2848 4902
rect 1974 4900 1980 4901
rect 1974 4896 1975 4900
rect 1979 4896 1980 4900
rect 2842 4897 2843 4901
rect 2847 4897 2848 4901
rect 2842 4896 2848 4897
rect 2978 4901 2984 4902
rect 2978 4897 2979 4901
rect 2983 4897 2984 4901
rect 2978 4896 2984 4897
rect 1974 4895 1980 4896
rect 267 4862 271 4863
rect 267 4857 271 4858
rect 315 4862 319 4863
rect 315 4857 319 4858
rect 403 4862 407 4863
rect 403 4857 407 4858
rect 523 4862 527 4863
rect 523 4857 527 4858
rect 539 4862 543 4863
rect 539 4857 543 4858
rect 675 4862 679 4863
rect 675 4857 679 4858
rect 723 4862 727 4863
rect 723 4857 727 4858
rect 915 4862 919 4863
rect 915 4857 919 4858
rect 1099 4862 1103 4863
rect 1099 4857 1103 4858
rect 1283 4862 1287 4863
rect 1283 4857 1287 4858
rect 1459 4862 1463 4863
rect 1459 4857 1463 4858
rect 1635 4862 1639 4863
rect 1635 4857 1639 4858
rect 1787 4862 1791 4863
rect 1787 4857 1791 4858
rect 1935 4862 1939 4863
rect 1935 4857 1939 4858
rect 226 4847 232 4848
rect 226 4843 227 4847
rect 231 4843 232 4847
rect 226 4842 232 4843
rect 268 4796 270 4857
rect 274 4843 280 4844
rect 274 4839 275 4843
rect 279 4839 280 4843
rect 274 4838 280 4839
rect 276 4804 278 4838
rect 274 4803 280 4804
rect 274 4799 275 4803
rect 279 4799 280 4803
rect 274 4798 280 4799
rect 404 4796 406 4857
rect 410 4843 416 4844
rect 410 4839 411 4843
rect 415 4839 416 4843
rect 410 4838 416 4839
rect 412 4804 414 4838
rect 410 4803 416 4804
rect 410 4799 411 4803
rect 415 4799 416 4803
rect 410 4798 416 4799
rect 540 4796 542 4857
rect 546 4843 552 4844
rect 546 4839 547 4843
rect 551 4839 552 4843
rect 546 4838 552 4839
rect 548 4804 550 4838
rect 546 4803 552 4804
rect 546 4799 547 4803
rect 551 4799 552 4803
rect 546 4798 552 4799
rect 676 4796 678 4857
rect 682 4843 688 4844
rect 682 4839 683 4843
rect 687 4839 688 4843
rect 682 4838 688 4839
rect 684 4804 686 4838
rect 682 4803 688 4804
rect 682 4799 683 4803
rect 687 4799 688 4803
rect 682 4798 688 4799
rect 690 4803 696 4804
rect 690 4799 691 4803
rect 695 4799 696 4803
rect 690 4798 696 4799
rect 110 4792 111 4796
rect 115 4792 116 4796
rect 110 4791 116 4792
rect 130 4795 136 4796
rect 130 4791 131 4795
rect 135 4791 136 4795
rect 130 4790 136 4791
rect 266 4795 272 4796
rect 266 4791 267 4795
rect 271 4791 272 4795
rect 266 4790 272 4791
rect 402 4795 408 4796
rect 402 4791 403 4795
rect 407 4791 408 4795
rect 402 4790 408 4791
rect 538 4795 544 4796
rect 538 4791 539 4795
rect 543 4791 544 4795
rect 538 4790 544 4791
rect 674 4795 680 4796
rect 674 4791 675 4795
rect 679 4791 680 4795
rect 674 4790 680 4791
rect 158 4780 164 4781
rect 110 4779 116 4780
rect 110 4775 111 4779
rect 115 4775 116 4779
rect 158 4776 159 4780
rect 163 4776 164 4780
rect 158 4775 164 4776
rect 294 4780 300 4781
rect 294 4776 295 4780
rect 299 4776 300 4780
rect 294 4775 300 4776
rect 430 4780 436 4781
rect 430 4776 431 4780
rect 435 4776 436 4780
rect 430 4775 436 4776
rect 566 4780 572 4781
rect 566 4776 567 4780
rect 571 4776 572 4780
rect 566 4775 572 4776
rect 110 4774 116 4775
rect 112 4743 114 4774
rect 160 4743 162 4775
rect 226 4743 232 4744
rect 296 4743 298 4775
rect 432 4743 434 4775
rect 568 4743 570 4775
rect 692 4744 694 4798
rect 1936 4797 1938 4857
rect 1976 4811 1978 4895
rect 2844 4811 2846 4896
rect 2938 4883 2944 4884
rect 2938 4879 2939 4883
rect 2943 4879 2944 4883
rect 2938 4878 2944 4879
rect 2940 4852 2942 4878
rect 2938 4851 2944 4852
rect 2938 4847 2939 4851
rect 2943 4847 2944 4851
rect 2938 4846 2944 4847
rect 2980 4811 2982 4896
rect 3020 4892 3022 5070
rect 3100 5024 3102 5085
rect 3652 5024 3654 5085
rect 3748 5076 3750 5142
rect 3800 5091 3802 5151
rect 3840 5143 3842 5194
rect 4280 5143 4282 5195
rect 3839 5142 3843 5143
rect 3839 5137 3843 5138
rect 3887 5142 3891 5143
rect 3887 5137 3891 5138
rect 4135 5142 4139 5143
rect 4135 5137 4139 5138
rect 4279 5142 4283 5143
rect 4279 5137 4283 5138
rect 4407 5142 4411 5143
rect 4407 5137 4411 5138
rect 3840 5114 3842 5137
rect 3838 5113 3844 5114
rect 3888 5113 3890 5137
rect 4136 5113 4138 5137
rect 4408 5113 4410 5137
rect 3838 5109 3839 5113
rect 3843 5109 3844 5113
rect 3838 5108 3844 5109
rect 3886 5112 3892 5113
rect 3886 5108 3887 5112
rect 3891 5108 3892 5112
rect 3886 5107 3892 5108
rect 4134 5112 4140 5113
rect 4134 5108 4135 5112
rect 4139 5108 4140 5112
rect 4134 5107 4140 5108
rect 4406 5112 4412 5113
rect 4406 5108 4407 5112
rect 4411 5108 4412 5112
rect 4406 5107 4412 5108
rect 3858 5097 3864 5098
rect 3838 5096 3844 5097
rect 3838 5092 3839 5096
rect 3843 5092 3844 5096
rect 3858 5093 3859 5097
rect 3863 5093 3864 5097
rect 3858 5092 3864 5093
rect 4106 5097 4112 5098
rect 4106 5093 4107 5097
rect 4111 5093 4112 5097
rect 4106 5092 4112 5093
rect 4378 5097 4384 5098
rect 4378 5093 4379 5097
rect 4383 5093 4384 5097
rect 4378 5092 4384 5093
rect 3838 5091 3844 5092
rect 3799 5090 3803 5091
rect 3799 5085 3803 5086
rect 3746 5075 3752 5076
rect 3746 5071 3747 5075
rect 3751 5071 3752 5075
rect 3746 5070 3752 5071
rect 3800 5025 3802 5085
rect 3798 5024 3804 5025
rect 3098 5023 3104 5024
rect 3098 5019 3099 5023
rect 3103 5019 3104 5023
rect 3098 5018 3104 5019
rect 3650 5023 3656 5024
rect 3650 5019 3651 5023
rect 3655 5019 3656 5023
rect 3798 5020 3799 5024
rect 3803 5020 3804 5024
rect 3798 5019 3804 5020
rect 3840 5019 3842 5091
rect 3860 5019 3862 5092
rect 3954 5087 3960 5088
rect 3954 5083 3955 5087
rect 3959 5083 3960 5087
rect 3954 5082 3960 5083
rect 3650 5018 3656 5019
rect 3839 5018 3843 5019
rect 3839 5013 3843 5014
rect 3859 5018 3863 5019
rect 3859 5013 3863 5014
rect 3126 5008 3132 5009
rect 3126 5004 3127 5008
rect 3131 5004 3132 5008
rect 3126 5003 3132 5004
rect 3678 5008 3684 5009
rect 3678 5004 3679 5008
rect 3683 5004 3684 5008
rect 3678 5003 3684 5004
rect 3798 5007 3804 5008
rect 3798 5003 3799 5007
rect 3803 5003 3804 5007
rect 3128 4947 3130 5003
rect 3680 4947 3682 5003
rect 3798 5002 3804 5003
rect 3800 4947 3802 5002
rect 3840 4953 3842 5013
rect 3838 4952 3844 4953
rect 3860 4952 3862 5013
rect 3956 5004 3958 5082
rect 4108 5019 4110 5092
rect 4234 5087 4240 5088
rect 4234 5083 4235 5087
rect 4239 5083 4240 5087
rect 4234 5082 4240 5083
rect 4202 5079 4208 5080
rect 4202 5075 4203 5079
rect 4207 5075 4208 5079
rect 4202 5074 4208 5075
rect 4204 5048 4206 5074
rect 4236 5048 4238 5082
rect 4202 5047 4208 5048
rect 4202 5043 4203 5047
rect 4207 5043 4208 5047
rect 4202 5042 4208 5043
rect 4234 5047 4240 5048
rect 4234 5043 4235 5047
rect 4239 5043 4240 5047
rect 4234 5042 4240 5043
rect 4380 5019 4382 5092
rect 4504 5088 4506 5262
rect 4716 5216 4718 5277
rect 4842 5223 4848 5224
rect 4842 5219 4843 5223
rect 4847 5219 4848 5223
rect 4842 5218 4848 5219
rect 4714 5215 4720 5216
rect 4714 5211 4715 5215
rect 4719 5211 4720 5215
rect 4714 5210 4720 5211
rect 4510 5200 4516 5201
rect 4510 5196 4511 5200
rect 4515 5196 4516 5200
rect 4510 5195 4516 5196
rect 4742 5200 4748 5201
rect 4742 5196 4743 5200
rect 4747 5196 4748 5200
rect 4742 5195 4748 5196
rect 4512 5143 4514 5195
rect 4744 5143 4746 5195
rect 4511 5142 4515 5143
rect 4511 5137 4515 5138
rect 4679 5142 4683 5143
rect 4679 5137 4683 5138
rect 4743 5142 4747 5143
rect 4743 5137 4747 5138
rect 4680 5113 4682 5137
rect 4678 5112 4684 5113
rect 4678 5108 4679 5112
rect 4683 5108 4684 5112
rect 4678 5107 4684 5108
rect 4650 5097 4656 5098
rect 4650 5093 4651 5097
rect 4655 5093 4656 5097
rect 4650 5092 4656 5093
rect 4502 5087 4508 5088
rect 4502 5083 4503 5087
rect 4507 5083 4508 5087
rect 4502 5082 4508 5083
rect 4652 5019 4654 5092
rect 4844 5048 4846 5218
rect 4948 5216 4950 5277
rect 5188 5216 5190 5277
rect 5224 5268 5226 5350
rect 5664 5283 5666 5359
rect 5663 5282 5667 5283
rect 5663 5277 5667 5278
rect 5222 5267 5228 5268
rect 5222 5263 5223 5267
rect 5227 5263 5228 5267
rect 5222 5262 5228 5263
rect 5664 5217 5666 5277
rect 5662 5216 5668 5217
rect 4946 5215 4952 5216
rect 4946 5211 4947 5215
rect 4951 5211 4952 5215
rect 4946 5210 4952 5211
rect 5186 5215 5192 5216
rect 5186 5211 5187 5215
rect 5191 5211 5192 5215
rect 5662 5212 5663 5216
rect 5667 5212 5668 5216
rect 5662 5211 5668 5212
rect 5186 5210 5192 5211
rect 4974 5200 4980 5201
rect 4974 5196 4975 5200
rect 4979 5196 4980 5200
rect 4974 5195 4980 5196
rect 5214 5200 5220 5201
rect 5214 5196 5215 5200
rect 5219 5196 5220 5200
rect 5214 5195 5220 5196
rect 5662 5199 5668 5200
rect 5662 5195 5663 5199
rect 5667 5195 5668 5199
rect 4976 5143 4978 5195
rect 5216 5143 5218 5195
rect 5662 5194 5668 5195
rect 5664 5143 5666 5194
rect 4959 5142 4963 5143
rect 4959 5137 4963 5138
rect 4975 5142 4979 5143
rect 4975 5137 4979 5138
rect 5215 5142 5219 5143
rect 5215 5137 5219 5138
rect 5239 5142 5243 5143
rect 5239 5137 5243 5138
rect 5663 5142 5667 5143
rect 5663 5137 5667 5138
rect 4960 5113 4962 5137
rect 5240 5113 5242 5137
rect 5664 5114 5666 5137
rect 5662 5113 5668 5114
rect 4958 5112 4964 5113
rect 4958 5108 4959 5112
rect 4963 5108 4964 5112
rect 4958 5107 4964 5108
rect 5238 5112 5244 5113
rect 5238 5108 5239 5112
rect 5243 5108 5244 5112
rect 5662 5109 5663 5113
rect 5667 5109 5668 5113
rect 5662 5108 5668 5109
rect 5238 5107 5244 5108
rect 4930 5097 4936 5098
rect 4930 5093 4931 5097
rect 4935 5093 4936 5097
rect 4930 5092 4936 5093
rect 5210 5097 5216 5098
rect 5210 5093 5211 5097
rect 5215 5093 5216 5097
rect 5210 5092 5216 5093
rect 5662 5096 5668 5097
rect 5662 5092 5663 5096
rect 5667 5092 5668 5096
rect 4746 5047 4752 5048
rect 4746 5043 4747 5047
rect 4751 5043 4752 5047
rect 4746 5042 4752 5043
rect 4842 5047 4848 5048
rect 4842 5043 4843 5047
rect 4847 5043 4848 5047
rect 4842 5042 4848 5043
rect 4019 5018 4023 5019
rect 4019 5013 4023 5014
rect 4107 5018 4111 5019
rect 4107 5013 4111 5014
rect 4211 5018 4215 5019
rect 4211 5013 4215 5014
rect 4379 5018 4383 5019
rect 4379 5013 4383 5014
rect 4411 5018 4415 5019
rect 4411 5013 4415 5014
rect 4627 5018 4631 5019
rect 4627 5013 4631 5014
rect 4651 5018 4655 5019
rect 4651 5013 4655 5014
rect 3954 5003 3960 5004
rect 3954 4999 3955 5003
rect 3959 4999 3960 5003
rect 3954 4998 3960 4999
rect 4020 4952 4022 5013
rect 4026 4999 4032 5000
rect 4026 4995 4027 4999
rect 4031 4995 4032 4999
rect 4026 4994 4032 4995
rect 4028 4960 4030 4994
rect 4026 4959 4032 4960
rect 4026 4955 4027 4959
rect 4031 4955 4032 4959
rect 4026 4954 4032 4955
rect 4212 4952 4214 5013
rect 4218 4999 4224 5000
rect 4218 4995 4219 4999
rect 4223 4995 4224 4999
rect 4218 4994 4224 4995
rect 4220 4960 4222 4994
rect 4218 4959 4224 4960
rect 4218 4955 4219 4959
rect 4223 4955 4224 4959
rect 4218 4954 4224 4955
rect 4334 4959 4340 4960
rect 4334 4955 4335 4959
rect 4339 4955 4340 4959
rect 4334 4954 4340 4955
rect 3838 4948 3839 4952
rect 3843 4948 3844 4952
rect 3838 4947 3844 4948
rect 3858 4951 3864 4952
rect 3858 4947 3859 4951
rect 3863 4947 3864 4951
rect 3127 4946 3131 4947
rect 3127 4941 3131 4942
rect 3679 4946 3683 4947
rect 3679 4941 3683 4942
rect 3799 4946 3803 4947
rect 3858 4946 3864 4947
rect 4018 4951 4024 4952
rect 4018 4947 4019 4951
rect 4023 4947 4024 4951
rect 4018 4946 4024 4947
rect 4210 4951 4216 4952
rect 4210 4947 4211 4951
rect 4215 4947 4216 4951
rect 4210 4946 4216 4947
rect 3799 4941 3803 4942
rect 3800 4918 3802 4941
rect 3886 4936 3892 4937
rect 3838 4935 3844 4936
rect 3838 4931 3839 4935
rect 3843 4931 3844 4935
rect 3886 4932 3887 4936
rect 3891 4932 3892 4936
rect 3886 4931 3892 4932
rect 4046 4936 4052 4937
rect 4046 4932 4047 4936
rect 4051 4932 4052 4936
rect 4046 4931 4052 4932
rect 4238 4936 4244 4937
rect 4238 4932 4239 4936
rect 4243 4932 4244 4936
rect 4238 4931 4244 4932
rect 3838 4930 3844 4931
rect 3798 4917 3804 4918
rect 3798 4913 3799 4917
rect 3803 4913 3804 4917
rect 3798 4912 3804 4913
rect 3798 4900 3804 4901
rect 3798 4896 3799 4900
rect 3803 4896 3804 4900
rect 3798 4895 3804 4896
rect 3018 4891 3024 4892
rect 3018 4887 3019 4891
rect 3023 4887 3024 4891
rect 3018 4886 3024 4887
rect 3146 4851 3152 4852
rect 3146 4847 3147 4851
rect 3151 4847 3152 4851
rect 3146 4846 3152 4847
rect 1975 4810 1979 4811
rect 1975 4805 1979 4806
rect 1995 4810 1999 4811
rect 1995 4805 1999 4806
rect 2155 4810 2159 4811
rect 2155 4805 2159 4806
rect 2347 4810 2351 4811
rect 2347 4805 2351 4806
rect 2539 4810 2543 4811
rect 2539 4805 2543 4806
rect 2731 4810 2735 4811
rect 2731 4805 2735 4806
rect 2843 4810 2847 4811
rect 2843 4805 2847 4806
rect 2931 4810 2935 4811
rect 2931 4805 2935 4806
rect 2979 4810 2983 4811
rect 2979 4805 2983 4806
rect 3131 4810 3135 4811
rect 3131 4805 3135 4806
rect 1934 4796 1940 4797
rect 1934 4792 1935 4796
rect 1939 4792 1940 4796
rect 1934 4791 1940 4792
rect 1966 4795 1972 4796
rect 1966 4791 1967 4795
rect 1971 4791 1972 4795
rect 1966 4790 1972 4791
rect 702 4780 708 4781
rect 702 4776 703 4780
rect 707 4776 708 4780
rect 702 4775 708 4776
rect 1934 4779 1940 4780
rect 1934 4775 1935 4779
rect 1939 4775 1940 4779
rect 690 4743 696 4744
rect 704 4743 706 4775
rect 1934 4774 1940 4775
rect 1936 4743 1938 4774
rect 111 4742 115 4743
rect 111 4737 115 4738
rect 159 4742 163 4743
rect 226 4739 227 4743
rect 231 4739 232 4743
rect 226 4738 232 4739
rect 295 4742 299 4743
rect 159 4737 163 4738
rect 112 4714 114 4737
rect 110 4713 116 4714
rect 160 4713 162 4737
rect 110 4709 111 4713
rect 115 4709 116 4713
rect 110 4708 116 4709
rect 158 4712 164 4713
rect 158 4708 159 4712
rect 163 4708 164 4712
rect 158 4707 164 4708
rect 130 4697 136 4698
rect 110 4696 116 4697
rect 110 4692 111 4696
rect 115 4692 116 4696
rect 130 4693 131 4697
rect 135 4693 136 4697
rect 130 4692 136 4693
rect 110 4691 116 4692
rect 112 4615 114 4691
rect 132 4615 134 4692
rect 228 4648 230 4738
rect 295 4737 299 4738
rect 343 4742 347 4743
rect 343 4737 347 4738
rect 431 4742 435 4743
rect 431 4737 435 4738
rect 567 4742 571 4743
rect 690 4739 691 4743
rect 695 4739 696 4743
rect 690 4738 696 4739
rect 703 4742 707 4743
rect 567 4737 571 4738
rect 703 4737 707 4738
rect 807 4742 811 4743
rect 807 4737 811 4738
rect 1055 4742 1059 4743
rect 1055 4737 1059 4738
rect 1311 4742 1315 4743
rect 1311 4737 1315 4738
rect 1575 4742 1579 4743
rect 1575 4737 1579 4738
rect 1815 4742 1819 4743
rect 1815 4737 1819 4738
rect 1935 4742 1939 4743
rect 1935 4737 1939 4738
rect 344 4713 346 4737
rect 568 4713 570 4737
rect 808 4713 810 4737
rect 1056 4713 1058 4737
rect 1312 4713 1314 4737
rect 1576 4713 1578 4737
rect 1816 4713 1818 4737
rect 1936 4714 1938 4737
rect 1934 4713 1940 4714
rect 342 4712 348 4713
rect 342 4708 343 4712
rect 347 4708 348 4712
rect 342 4707 348 4708
rect 566 4712 572 4713
rect 566 4708 567 4712
rect 571 4708 572 4712
rect 566 4707 572 4708
rect 806 4712 812 4713
rect 806 4708 807 4712
rect 811 4708 812 4712
rect 806 4707 812 4708
rect 1054 4712 1060 4713
rect 1054 4708 1055 4712
rect 1059 4708 1060 4712
rect 1054 4707 1060 4708
rect 1310 4712 1316 4713
rect 1310 4708 1311 4712
rect 1315 4708 1316 4712
rect 1310 4707 1316 4708
rect 1574 4712 1580 4713
rect 1574 4708 1575 4712
rect 1579 4708 1580 4712
rect 1574 4707 1580 4708
rect 1814 4712 1820 4713
rect 1814 4708 1815 4712
rect 1819 4708 1820 4712
rect 1934 4709 1935 4713
rect 1939 4709 1940 4713
rect 1934 4708 1940 4709
rect 1814 4707 1820 4708
rect 314 4697 320 4698
rect 314 4693 315 4697
rect 319 4693 320 4697
rect 314 4692 320 4693
rect 538 4697 544 4698
rect 538 4693 539 4697
rect 543 4693 544 4697
rect 538 4692 544 4693
rect 778 4697 784 4698
rect 778 4693 779 4697
rect 783 4693 784 4697
rect 778 4692 784 4693
rect 1026 4697 1032 4698
rect 1026 4693 1027 4697
rect 1031 4693 1032 4697
rect 1026 4692 1032 4693
rect 1282 4697 1288 4698
rect 1282 4693 1283 4697
rect 1287 4693 1288 4697
rect 1282 4692 1288 4693
rect 1546 4697 1552 4698
rect 1546 4693 1547 4697
rect 1551 4693 1552 4697
rect 1546 4692 1552 4693
rect 1786 4697 1792 4698
rect 1786 4693 1787 4697
rect 1791 4693 1792 4697
rect 1786 4692 1792 4693
rect 1934 4696 1940 4697
rect 1934 4692 1935 4696
rect 1939 4692 1940 4696
rect 226 4647 232 4648
rect 226 4643 227 4647
rect 231 4643 232 4647
rect 226 4642 232 4643
rect 316 4615 318 4692
rect 442 4687 448 4688
rect 442 4683 443 4687
rect 447 4683 448 4687
rect 442 4682 448 4683
rect 444 4648 446 4682
rect 442 4647 448 4648
rect 442 4643 443 4647
rect 447 4643 448 4647
rect 442 4642 448 4643
rect 540 4615 542 4692
rect 666 4687 672 4688
rect 666 4683 667 4687
rect 671 4683 672 4687
rect 666 4682 672 4683
rect 668 4648 670 4682
rect 666 4647 672 4648
rect 666 4643 667 4647
rect 671 4643 672 4647
rect 666 4642 672 4643
rect 780 4615 782 4692
rect 906 4687 912 4688
rect 906 4683 907 4687
rect 911 4683 912 4687
rect 906 4682 912 4683
rect 1010 4687 1016 4688
rect 1010 4683 1011 4687
rect 1015 4683 1016 4687
rect 1010 4682 1016 4683
rect 908 4648 910 4682
rect 906 4647 912 4648
rect 906 4643 907 4647
rect 911 4643 912 4647
rect 906 4642 912 4643
rect 111 4614 115 4615
rect 111 4609 115 4610
rect 131 4614 135 4615
rect 131 4609 135 4610
rect 171 4614 175 4615
rect 171 4609 175 4610
rect 315 4614 319 4615
rect 315 4609 319 4610
rect 395 4614 399 4615
rect 395 4609 399 4610
rect 539 4614 543 4615
rect 539 4609 543 4610
rect 643 4614 647 4615
rect 643 4609 647 4610
rect 779 4614 783 4615
rect 779 4609 783 4610
rect 907 4614 911 4615
rect 907 4609 911 4610
rect 112 4549 114 4609
rect 110 4548 116 4549
rect 172 4548 174 4609
rect 396 4548 398 4609
rect 402 4595 408 4596
rect 402 4591 403 4595
rect 407 4591 408 4595
rect 402 4590 408 4591
rect 404 4556 406 4590
rect 402 4555 408 4556
rect 402 4551 403 4555
rect 407 4551 408 4555
rect 402 4550 408 4551
rect 644 4548 646 4609
rect 650 4595 656 4596
rect 650 4591 651 4595
rect 655 4591 656 4595
rect 650 4590 656 4591
rect 652 4556 654 4590
rect 650 4555 656 4556
rect 650 4551 651 4555
rect 655 4551 656 4555
rect 650 4550 656 4551
rect 908 4548 910 4609
rect 1012 4604 1014 4682
rect 1028 4615 1030 4692
rect 1284 4615 1286 4692
rect 1410 4687 1416 4688
rect 1410 4683 1411 4687
rect 1415 4683 1416 4687
rect 1410 4682 1416 4683
rect 1412 4648 1414 4682
rect 1410 4647 1416 4648
rect 1410 4643 1411 4647
rect 1415 4643 1416 4647
rect 1410 4642 1416 4643
rect 1518 4639 1524 4640
rect 1518 4635 1519 4639
rect 1523 4635 1524 4639
rect 1518 4634 1524 4635
rect 1027 4614 1031 4615
rect 1027 4609 1031 4610
rect 1195 4614 1199 4615
rect 1195 4609 1199 4610
rect 1283 4614 1287 4615
rect 1283 4609 1287 4610
rect 1491 4614 1495 4615
rect 1491 4609 1495 4610
rect 1010 4603 1016 4604
rect 1010 4599 1011 4603
rect 1015 4599 1016 4603
rect 1010 4598 1016 4599
rect 914 4595 920 4596
rect 914 4591 915 4595
rect 919 4591 920 4595
rect 914 4590 920 4591
rect 916 4556 918 4590
rect 914 4555 920 4556
rect 914 4551 915 4555
rect 919 4551 920 4555
rect 914 4550 920 4551
rect 1196 4548 1198 4609
rect 1202 4595 1208 4596
rect 1202 4591 1203 4595
rect 1207 4591 1208 4595
rect 1202 4590 1208 4591
rect 1204 4556 1206 4590
rect 1202 4555 1208 4556
rect 1202 4551 1203 4555
rect 1207 4551 1208 4555
rect 1202 4550 1208 4551
rect 1230 4555 1236 4556
rect 1230 4551 1231 4555
rect 1235 4551 1236 4555
rect 1230 4550 1236 4551
rect 110 4544 111 4548
rect 115 4544 116 4548
rect 110 4543 116 4544
rect 170 4547 176 4548
rect 170 4543 171 4547
rect 175 4543 176 4547
rect 170 4542 176 4543
rect 394 4547 400 4548
rect 394 4543 395 4547
rect 399 4543 400 4547
rect 394 4542 400 4543
rect 642 4547 648 4548
rect 642 4543 643 4547
rect 647 4543 648 4547
rect 642 4542 648 4543
rect 906 4547 912 4548
rect 906 4543 907 4547
rect 911 4543 912 4547
rect 906 4542 912 4543
rect 1194 4547 1200 4548
rect 1194 4543 1195 4547
rect 1199 4543 1200 4547
rect 1194 4542 1200 4543
rect 198 4532 204 4533
rect 110 4531 116 4532
rect 110 4527 111 4531
rect 115 4527 116 4531
rect 198 4528 199 4532
rect 203 4528 204 4532
rect 198 4527 204 4528
rect 422 4532 428 4533
rect 422 4528 423 4532
rect 427 4528 428 4532
rect 422 4527 428 4528
rect 670 4532 676 4533
rect 670 4528 671 4532
rect 675 4528 676 4532
rect 670 4527 676 4528
rect 934 4532 940 4533
rect 934 4528 935 4532
rect 939 4528 940 4532
rect 934 4527 940 4528
rect 1222 4532 1228 4533
rect 1222 4528 1223 4532
rect 1227 4528 1228 4532
rect 1222 4527 1228 4528
rect 110 4526 116 4527
rect 112 4499 114 4526
rect 200 4499 202 4527
rect 424 4499 426 4527
rect 672 4499 674 4527
rect 936 4499 938 4527
rect 1224 4499 1226 4527
rect 111 4498 115 4499
rect 111 4493 115 4494
rect 199 4498 203 4499
rect 199 4493 203 4494
rect 423 4498 427 4499
rect 423 4493 427 4494
rect 447 4498 451 4499
rect 447 4493 451 4494
rect 655 4498 659 4499
rect 655 4493 659 4494
rect 671 4498 675 4499
rect 671 4493 675 4494
rect 887 4498 891 4499
rect 887 4493 891 4494
rect 935 4498 939 4499
rect 935 4493 939 4494
rect 1143 4498 1147 4499
rect 1143 4493 1147 4494
rect 1223 4498 1227 4499
rect 1223 4493 1227 4494
rect 112 4470 114 4493
rect 110 4469 116 4470
rect 448 4469 450 4493
rect 656 4469 658 4493
rect 888 4469 890 4493
rect 1144 4469 1146 4493
rect 110 4465 111 4469
rect 115 4465 116 4469
rect 110 4464 116 4465
rect 446 4468 452 4469
rect 446 4464 447 4468
rect 451 4464 452 4468
rect 446 4463 452 4464
rect 654 4468 660 4469
rect 654 4464 655 4468
rect 659 4464 660 4468
rect 654 4463 660 4464
rect 886 4468 892 4469
rect 886 4464 887 4468
rect 891 4464 892 4468
rect 886 4463 892 4464
rect 1142 4468 1148 4469
rect 1142 4464 1143 4468
rect 1147 4464 1148 4468
rect 1142 4463 1148 4464
rect 418 4453 424 4454
rect 110 4452 116 4453
rect 110 4448 111 4452
rect 115 4448 116 4452
rect 418 4449 419 4453
rect 423 4449 424 4453
rect 418 4448 424 4449
rect 626 4453 632 4454
rect 626 4449 627 4453
rect 631 4449 632 4453
rect 626 4448 632 4449
rect 858 4453 864 4454
rect 858 4449 859 4453
rect 863 4449 864 4453
rect 858 4448 864 4449
rect 1114 4453 1120 4454
rect 1114 4449 1115 4453
rect 1119 4449 1120 4453
rect 1114 4448 1120 4449
rect 110 4447 116 4448
rect 112 4383 114 4447
rect 420 4383 422 4448
rect 586 4443 592 4444
rect 586 4439 587 4443
rect 591 4439 592 4443
rect 586 4438 592 4439
rect 514 4435 520 4436
rect 514 4431 515 4435
rect 519 4431 520 4435
rect 514 4430 520 4431
rect 516 4404 518 4430
rect 588 4404 590 4438
rect 514 4403 520 4404
rect 514 4399 515 4403
rect 519 4399 520 4403
rect 514 4398 520 4399
rect 586 4403 592 4404
rect 586 4399 587 4403
rect 591 4399 592 4403
rect 586 4398 592 4399
rect 628 4383 630 4448
rect 754 4443 760 4444
rect 754 4439 755 4443
rect 759 4439 760 4443
rect 754 4438 760 4439
rect 756 4404 758 4438
rect 754 4403 760 4404
rect 754 4399 755 4403
rect 759 4399 760 4403
rect 754 4398 760 4399
rect 860 4383 862 4448
rect 1078 4443 1084 4444
rect 1078 4439 1079 4443
rect 1083 4439 1084 4443
rect 1078 4438 1084 4439
rect 1080 4404 1082 4438
rect 1078 4403 1084 4404
rect 1078 4399 1079 4403
rect 1083 4399 1084 4403
rect 1078 4398 1084 4399
rect 1116 4383 1118 4448
rect 1232 4436 1234 4550
rect 1492 4548 1494 4609
rect 1520 4556 1522 4634
rect 1548 4615 1550 4692
rect 1674 4687 1680 4688
rect 1674 4683 1675 4687
rect 1679 4683 1680 4687
rect 1674 4682 1680 4683
rect 1676 4648 1678 4682
rect 1674 4647 1680 4648
rect 1674 4643 1675 4647
rect 1679 4643 1680 4647
rect 1674 4642 1680 4643
rect 1788 4615 1790 4692
rect 1934 4691 1940 4692
rect 1936 4615 1938 4691
rect 1968 4688 1970 4790
rect 1976 4745 1978 4805
rect 1974 4744 1980 4745
rect 1996 4744 1998 4805
rect 2156 4744 2158 4805
rect 2162 4791 2168 4792
rect 2162 4787 2163 4791
rect 2167 4787 2168 4791
rect 2162 4786 2168 4787
rect 2164 4752 2166 4786
rect 2162 4751 2168 4752
rect 2162 4747 2163 4751
rect 2167 4747 2168 4751
rect 2162 4746 2168 4747
rect 2348 4744 2350 4805
rect 2354 4791 2360 4792
rect 2354 4787 2355 4791
rect 2359 4787 2360 4791
rect 2354 4786 2360 4787
rect 2356 4752 2358 4786
rect 2354 4751 2360 4752
rect 2354 4747 2355 4751
rect 2359 4747 2360 4751
rect 2354 4746 2360 4747
rect 2540 4744 2542 4805
rect 2546 4791 2552 4792
rect 2546 4787 2547 4791
rect 2551 4787 2552 4791
rect 2546 4786 2552 4787
rect 2548 4752 2550 4786
rect 2546 4751 2552 4752
rect 2546 4747 2547 4751
rect 2551 4747 2552 4751
rect 2546 4746 2552 4747
rect 2658 4751 2664 4752
rect 2658 4747 2659 4751
rect 2663 4747 2664 4751
rect 2658 4746 2664 4747
rect 1974 4740 1975 4744
rect 1979 4740 1980 4744
rect 1974 4739 1980 4740
rect 1994 4743 2000 4744
rect 1994 4739 1995 4743
rect 1999 4739 2000 4743
rect 1994 4738 2000 4739
rect 2154 4743 2160 4744
rect 2154 4739 2155 4743
rect 2159 4739 2160 4743
rect 2154 4738 2160 4739
rect 2346 4743 2352 4744
rect 2346 4739 2347 4743
rect 2351 4739 2352 4743
rect 2346 4738 2352 4739
rect 2538 4743 2544 4744
rect 2538 4739 2539 4743
rect 2543 4739 2544 4743
rect 2538 4738 2544 4739
rect 2022 4728 2028 4729
rect 1974 4727 1980 4728
rect 1974 4723 1975 4727
rect 1979 4723 1980 4727
rect 2022 4724 2023 4728
rect 2027 4724 2028 4728
rect 2022 4723 2028 4724
rect 2182 4728 2188 4729
rect 2182 4724 2183 4728
rect 2187 4724 2188 4728
rect 2182 4723 2188 4724
rect 2374 4728 2380 4729
rect 2374 4724 2375 4728
rect 2379 4724 2380 4728
rect 2374 4723 2380 4724
rect 2566 4728 2572 4729
rect 2566 4724 2567 4728
rect 2571 4724 2572 4728
rect 2566 4723 2572 4724
rect 1974 4722 1980 4723
rect 1976 4695 1978 4722
rect 2024 4695 2026 4723
rect 2184 4695 2186 4723
rect 2376 4695 2378 4723
rect 2568 4695 2570 4723
rect 1975 4694 1979 4695
rect 1975 4689 1979 4690
rect 2023 4694 2027 4695
rect 2023 4689 2027 4690
rect 2183 4694 2187 4695
rect 2183 4689 2187 4690
rect 2239 4694 2243 4695
rect 2239 4689 2243 4690
rect 2375 4694 2379 4695
rect 2375 4689 2379 4690
rect 2471 4694 2475 4695
rect 2471 4689 2475 4690
rect 2567 4694 2571 4695
rect 2567 4689 2571 4690
rect 1966 4687 1972 4688
rect 1966 4683 1967 4687
rect 1971 4683 1972 4687
rect 1966 4682 1972 4683
rect 1976 4666 1978 4689
rect 1974 4665 1980 4666
rect 2024 4665 2026 4689
rect 2240 4665 2242 4689
rect 2472 4665 2474 4689
rect 1974 4661 1975 4665
rect 1979 4661 1980 4665
rect 1974 4660 1980 4661
rect 2022 4664 2028 4665
rect 2022 4660 2023 4664
rect 2027 4660 2028 4664
rect 2022 4659 2028 4660
rect 2238 4664 2244 4665
rect 2238 4660 2239 4664
rect 2243 4660 2244 4664
rect 2238 4659 2244 4660
rect 2470 4664 2476 4665
rect 2470 4660 2471 4664
rect 2475 4660 2476 4664
rect 2470 4659 2476 4660
rect 1994 4649 2000 4650
rect 1974 4648 1980 4649
rect 1974 4644 1975 4648
rect 1979 4644 1980 4648
rect 1994 4645 1995 4649
rect 1999 4645 2000 4649
rect 1994 4644 2000 4645
rect 2210 4649 2216 4650
rect 2210 4645 2211 4649
rect 2215 4645 2216 4649
rect 2210 4644 2216 4645
rect 2442 4649 2448 4650
rect 2442 4645 2443 4649
rect 2447 4645 2448 4649
rect 2442 4644 2448 4645
rect 1974 4643 1980 4644
rect 1547 4614 1551 4615
rect 1547 4609 1551 4610
rect 1787 4614 1791 4615
rect 1787 4609 1791 4610
rect 1935 4614 1939 4615
rect 1935 4609 1939 4610
rect 1518 4555 1524 4556
rect 1518 4551 1519 4555
rect 1523 4551 1524 4555
rect 1518 4550 1524 4551
rect 1788 4548 1790 4609
rect 1906 4603 1912 4604
rect 1906 4599 1907 4603
rect 1911 4599 1912 4603
rect 1906 4598 1912 4599
rect 1794 4595 1800 4596
rect 1794 4591 1795 4595
rect 1799 4591 1800 4595
rect 1794 4590 1800 4591
rect 1490 4547 1496 4548
rect 1490 4543 1491 4547
rect 1495 4543 1496 4547
rect 1490 4542 1496 4543
rect 1786 4547 1792 4548
rect 1786 4543 1787 4547
rect 1791 4543 1792 4547
rect 1786 4542 1792 4543
rect 1518 4532 1524 4533
rect 1518 4528 1519 4532
rect 1523 4528 1524 4532
rect 1518 4527 1524 4528
rect 1520 4499 1522 4527
rect 1407 4498 1411 4499
rect 1407 4493 1411 4494
rect 1519 4498 1523 4499
rect 1519 4493 1523 4494
rect 1679 4498 1683 4499
rect 1679 4493 1683 4494
rect 1408 4469 1410 4493
rect 1680 4469 1682 4493
rect 1406 4468 1412 4469
rect 1406 4464 1407 4468
rect 1411 4464 1412 4468
rect 1406 4463 1412 4464
rect 1678 4468 1684 4469
rect 1678 4464 1679 4468
rect 1683 4464 1684 4468
rect 1678 4463 1684 4464
rect 1378 4453 1384 4454
rect 1378 4449 1379 4453
rect 1383 4449 1384 4453
rect 1378 4448 1384 4449
rect 1650 4453 1656 4454
rect 1650 4449 1651 4453
rect 1655 4449 1656 4453
rect 1650 4448 1656 4449
rect 1242 4443 1248 4444
rect 1242 4439 1243 4443
rect 1247 4439 1248 4443
rect 1242 4438 1248 4439
rect 1274 4443 1280 4444
rect 1274 4439 1275 4443
rect 1279 4439 1280 4443
rect 1274 4438 1280 4439
rect 1230 4435 1236 4436
rect 1230 4431 1231 4435
rect 1235 4431 1236 4435
rect 1230 4430 1236 4431
rect 1244 4404 1246 4438
rect 1242 4403 1248 4404
rect 1242 4399 1243 4403
rect 1247 4399 1248 4403
rect 1242 4398 1248 4399
rect 111 4382 115 4383
rect 111 4377 115 4378
rect 419 4382 423 4383
rect 419 4377 423 4378
rect 627 4382 631 4383
rect 627 4377 631 4378
rect 667 4382 671 4383
rect 667 4377 671 4378
rect 811 4382 815 4383
rect 811 4377 815 4378
rect 859 4382 863 4383
rect 859 4377 863 4378
rect 963 4382 967 4383
rect 963 4377 967 4378
rect 1115 4382 1119 4383
rect 1115 4377 1119 4378
rect 1123 4382 1127 4383
rect 1123 4377 1127 4378
rect 112 4317 114 4377
rect 110 4316 116 4317
rect 668 4316 670 4377
rect 812 4316 814 4377
rect 818 4363 824 4364
rect 818 4359 819 4363
rect 823 4359 824 4363
rect 818 4358 824 4359
rect 820 4324 822 4358
rect 818 4323 824 4324
rect 818 4319 819 4323
rect 823 4319 824 4323
rect 818 4318 824 4319
rect 964 4316 966 4377
rect 970 4363 976 4364
rect 970 4359 971 4363
rect 975 4359 976 4363
rect 970 4358 976 4359
rect 972 4324 974 4358
rect 970 4323 976 4324
rect 970 4319 971 4323
rect 975 4319 976 4323
rect 970 4318 976 4319
rect 1124 4316 1126 4377
rect 1276 4372 1278 4438
rect 1380 4383 1382 4448
rect 1652 4383 1654 4448
rect 1796 4444 1798 4590
rect 1908 4556 1910 4598
rect 1906 4555 1912 4556
rect 1906 4551 1907 4555
rect 1911 4551 1912 4555
rect 1906 4550 1912 4551
rect 1936 4549 1938 4609
rect 1976 4579 1978 4643
rect 1996 4579 1998 4644
rect 2212 4579 2214 4644
rect 2338 4639 2344 4640
rect 2338 4635 2339 4639
rect 2343 4635 2344 4639
rect 2338 4634 2344 4635
rect 2340 4600 2342 4634
rect 2338 4599 2344 4600
rect 2338 4595 2339 4599
rect 2343 4595 2344 4599
rect 2338 4594 2344 4595
rect 2444 4579 2446 4644
rect 2660 4592 2662 4746
rect 2732 4744 2734 4805
rect 2790 4795 2796 4796
rect 2790 4791 2791 4795
rect 2795 4791 2796 4795
rect 2790 4790 2796 4791
rect 2730 4743 2736 4744
rect 2730 4739 2731 4743
rect 2735 4739 2736 4743
rect 2730 4738 2736 4739
rect 2758 4728 2764 4729
rect 2758 4724 2759 4728
rect 2763 4724 2764 4728
rect 2758 4723 2764 4724
rect 2760 4695 2762 4723
rect 2695 4694 2699 4695
rect 2695 4689 2699 4690
rect 2759 4694 2763 4695
rect 2759 4689 2763 4690
rect 2696 4665 2698 4689
rect 2694 4664 2700 4665
rect 2694 4660 2695 4664
rect 2699 4660 2700 4664
rect 2694 4659 2700 4660
rect 2666 4649 2672 4650
rect 2666 4645 2667 4649
rect 2671 4645 2672 4649
rect 2666 4644 2672 4645
rect 2658 4591 2664 4592
rect 2658 4587 2659 4591
rect 2663 4587 2664 4591
rect 2658 4586 2664 4587
rect 2668 4579 2670 4644
rect 2792 4640 2794 4790
rect 2932 4744 2934 4805
rect 2938 4791 2944 4792
rect 2938 4787 2939 4791
rect 2943 4787 2944 4791
rect 2938 4786 2944 4787
rect 2940 4752 2942 4786
rect 2938 4751 2944 4752
rect 2938 4747 2939 4751
rect 2943 4747 2944 4751
rect 2938 4746 2944 4747
rect 3132 4744 3134 4805
rect 3138 4791 3144 4792
rect 3138 4787 3139 4791
rect 3143 4787 3144 4791
rect 3138 4786 3144 4787
rect 3140 4752 3142 4786
rect 3148 4752 3150 4846
rect 3800 4811 3802 4895
rect 3840 4887 3842 4930
rect 3888 4887 3890 4931
rect 4048 4887 4050 4931
rect 4240 4887 4242 4931
rect 3839 4886 3843 4887
rect 3839 4881 3843 4882
rect 3887 4886 3891 4887
rect 3887 4881 3891 4882
rect 4047 4886 4051 4887
rect 4047 4881 4051 4882
rect 4071 4886 4075 4887
rect 4071 4881 4075 4882
rect 4239 4886 4243 4887
rect 4239 4881 4243 4882
rect 4287 4886 4291 4887
rect 4287 4881 4291 4882
rect 3840 4858 3842 4881
rect 3838 4857 3844 4858
rect 3888 4857 3890 4881
rect 4072 4857 4074 4881
rect 4288 4857 4290 4881
rect 3838 4853 3839 4857
rect 3843 4853 3844 4857
rect 3838 4852 3844 4853
rect 3886 4856 3892 4857
rect 3886 4852 3887 4856
rect 3891 4852 3892 4856
rect 3886 4851 3892 4852
rect 4070 4856 4076 4857
rect 4070 4852 4071 4856
rect 4075 4852 4076 4856
rect 4070 4851 4076 4852
rect 4286 4856 4292 4857
rect 4286 4852 4287 4856
rect 4291 4852 4292 4856
rect 4286 4851 4292 4852
rect 3858 4841 3864 4842
rect 3838 4840 3844 4841
rect 3838 4836 3839 4840
rect 3843 4836 3844 4840
rect 3858 4837 3859 4841
rect 3863 4837 3864 4841
rect 3858 4836 3864 4837
rect 4042 4841 4048 4842
rect 4042 4837 4043 4841
rect 4047 4837 4048 4841
rect 4042 4836 4048 4837
rect 4258 4841 4264 4842
rect 4258 4837 4259 4841
rect 4263 4837 4264 4841
rect 4258 4836 4264 4837
rect 3838 4835 3844 4836
rect 3799 4810 3803 4811
rect 3799 4805 3803 4806
rect 3138 4751 3144 4752
rect 3138 4747 3139 4751
rect 3143 4747 3144 4751
rect 3138 4746 3144 4747
rect 3146 4751 3152 4752
rect 3146 4747 3147 4751
rect 3151 4747 3152 4751
rect 3146 4746 3152 4747
rect 3800 4745 3802 4805
rect 3840 4771 3842 4835
rect 3860 4771 3862 4836
rect 3982 4831 3988 4832
rect 3982 4827 3983 4831
rect 3987 4827 3988 4831
rect 3982 4826 3988 4827
rect 3839 4770 3843 4771
rect 3839 4765 3843 4766
rect 3859 4770 3863 4771
rect 3859 4765 3863 4766
rect 3915 4770 3919 4771
rect 3915 4765 3919 4766
rect 3798 4744 3804 4745
rect 2930 4743 2936 4744
rect 2930 4739 2931 4743
rect 2935 4739 2936 4743
rect 2930 4738 2936 4739
rect 3130 4743 3136 4744
rect 3130 4739 3131 4743
rect 3135 4739 3136 4743
rect 3798 4740 3799 4744
rect 3803 4740 3804 4744
rect 3798 4739 3804 4740
rect 3130 4738 3136 4739
rect 2958 4728 2964 4729
rect 2958 4724 2959 4728
rect 2963 4724 2964 4728
rect 2958 4723 2964 4724
rect 3158 4728 3164 4729
rect 3158 4724 3159 4728
rect 3163 4724 3164 4728
rect 3158 4723 3164 4724
rect 3798 4727 3804 4728
rect 3798 4723 3799 4727
rect 3803 4723 3804 4727
rect 2960 4695 2962 4723
rect 3160 4695 3162 4723
rect 3798 4722 3804 4723
rect 3800 4695 3802 4722
rect 3840 4705 3842 4765
rect 3838 4704 3844 4705
rect 3916 4704 3918 4765
rect 3984 4756 3986 4826
rect 4044 4771 4046 4836
rect 4260 4771 4262 4836
rect 4336 4792 4338 4954
rect 4412 4952 4414 5013
rect 4628 4952 4630 5013
rect 4634 4999 4640 5000
rect 4634 4995 4635 4999
rect 4639 4995 4640 4999
rect 4634 4994 4640 4995
rect 4636 4960 4638 4994
rect 4748 4960 4750 5042
rect 4932 5019 4934 5092
rect 5058 5087 5064 5088
rect 5058 5083 5059 5087
rect 5063 5083 5064 5087
rect 5058 5082 5064 5083
rect 5060 5048 5062 5082
rect 5058 5047 5064 5048
rect 5058 5043 5059 5047
rect 5063 5043 5064 5047
rect 5058 5042 5064 5043
rect 5212 5019 5214 5092
rect 5662 5091 5668 5092
rect 5334 5087 5340 5088
rect 5334 5083 5335 5087
rect 5339 5083 5340 5087
rect 5334 5082 5340 5083
rect 4843 5018 4847 5019
rect 4843 5013 4847 5014
rect 4931 5018 4935 5019
rect 4931 5013 4935 5014
rect 5067 5018 5071 5019
rect 5067 5013 5071 5014
rect 5211 5018 5215 5019
rect 5211 5013 5215 5014
rect 5299 5018 5303 5019
rect 5299 5013 5303 5014
rect 4818 5007 4824 5008
rect 4818 5003 4819 5007
rect 4823 5003 4824 5007
rect 4818 5002 4824 5003
rect 4820 4960 4822 5002
rect 4634 4959 4640 4960
rect 4634 4955 4635 4959
rect 4639 4955 4640 4959
rect 4634 4954 4640 4955
rect 4746 4959 4752 4960
rect 4746 4955 4747 4959
rect 4751 4955 4752 4959
rect 4746 4954 4752 4955
rect 4818 4959 4824 4960
rect 4818 4955 4819 4959
rect 4823 4955 4824 4959
rect 4818 4954 4824 4955
rect 4844 4952 4846 5013
rect 4850 4999 4856 5000
rect 4850 4995 4851 4999
rect 4855 4995 4856 4999
rect 4850 4994 4856 4995
rect 4410 4951 4416 4952
rect 4410 4947 4411 4951
rect 4415 4947 4416 4951
rect 4410 4946 4416 4947
rect 4626 4951 4632 4952
rect 4626 4947 4627 4951
rect 4631 4947 4632 4951
rect 4626 4946 4632 4947
rect 4842 4951 4848 4952
rect 4842 4947 4843 4951
rect 4847 4947 4848 4951
rect 4842 4946 4848 4947
rect 4438 4936 4444 4937
rect 4438 4932 4439 4936
rect 4443 4932 4444 4936
rect 4438 4931 4444 4932
rect 4654 4936 4660 4937
rect 4654 4932 4655 4936
rect 4659 4932 4660 4936
rect 4654 4931 4660 4932
rect 4440 4887 4442 4931
rect 4656 4887 4658 4931
rect 4439 4886 4443 4887
rect 4439 4881 4443 4882
rect 4511 4886 4515 4887
rect 4511 4881 4515 4882
rect 4655 4886 4659 4887
rect 4655 4881 4659 4882
rect 4735 4886 4739 4887
rect 4735 4881 4739 4882
rect 4512 4857 4514 4881
rect 4736 4857 4738 4881
rect 4510 4856 4516 4857
rect 4510 4852 4511 4856
rect 4515 4852 4516 4856
rect 4510 4851 4516 4852
rect 4734 4856 4740 4857
rect 4734 4852 4735 4856
rect 4739 4852 4740 4856
rect 4734 4851 4740 4852
rect 4482 4841 4488 4842
rect 4482 4837 4483 4841
rect 4487 4837 4488 4841
rect 4482 4836 4488 4837
rect 4706 4841 4712 4842
rect 4706 4837 4707 4841
rect 4711 4837 4712 4841
rect 4706 4836 4712 4837
rect 4334 4791 4340 4792
rect 4334 4787 4335 4791
rect 4339 4787 4340 4791
rect 4334 4786 4340 4787
rect 4484 4771 4486 4836
rect 4610 4831 4616 4832
rect 4610 4827 4611 4831
rect 4615 4827 4616 4831
rect 4610 4826 4616 4827
rect 4578 4823 4584 4824
rect 4578 4819 4579 4823
rect 4583 4819 4584 4823
rect 4578 4818 4584 4819
rect 4580 4792 4582 4818
rect 4612 4792 4614 4826
rect 4578 4791 4584 4792
rect 4578 4787 4579 4791
rect 4583 4787 4584 4791
rect 4578 4786 4584 4787
rect 4610 4791 4616 4792
rect 4610 4787 4611 4791
rect 4615 4787 4616 4791
rect 4610 4786 4616 4787
rect 4708 4771 4710 4836
rect 4852 4832 4854 4994
rect 5068 4952 5070 5013
rect 5190 4959 5196 4960
rect 5190 4955 5191 4959
rect 5195 4955 5196 4959
rect 5190 4954 5196 4955
rect 5066 4951 5072 4952
rect 5066 4947 5067 4951
rect 5071 4947 5072 4951
rect 5066 4946 5072 4947
rect 4870 4936 4876 4937
rect 4870 4932 4871 4936
rect 4875 4932 4876 4936
rect 4870 4931 4876 4932
rect 5094 4936 5100 4937
rect 5094 4932 5095 4936
rect 5099 4932 5100 4936
rect 5094 4931 5100 4932
rect 4872 4887 4874 4931
rect 5096 4887 5098 4931
rect 4871 4886 4875 4887
rect 4871 4881 4875 4882
rect 4959 4886 4963 4887
rect 4959 4881 4963 4882
rect 5095 4886 5099 4887
rect 5095 4881 5099 4882
rect 5183 4886 5187 4887
rect 5183 4881 5187 4882
rect 4960 4857 4962 4881
rect 5184 4857 5186 4881
rect 4958 4856 4964 4857
rect 4958 4852 4959 4856
rect 4963 4852 4964 4856
rect 4958 4851 4964 4852
rect 5182 4856 5188 4857
rect 5182 4852 5183 4856
rect 5187 4852 5188 4856
rect 5182 4851 5188 4852
rect 4930 4841 4936 4842
rect 4930 4837 4931 4841
rect 4935 4837 4936 4841
rect 4930 4836 4936 4837
rect 5154 4841 5160 4842
rect 5154 4837 5155 4841
rect 5159 4837 5160 4841
rect 5154 4836 5160 4837
rect 4850 4831 4856 4832
rect 4850 4827 4851 4831
rect 4855 4827 4856 4831
rect 4850 4826 4856 4827
rect 4932 4771 4934 4836
rect 5082 4791 5088 4792
rect 5082 4787 5083 4791
rect 5087 4787 5088 4791
rect 5082 4786 5088 4787
rect 4043 4770 4047 4771
rect 4043 4765 4047 4766
rect 4187 4770 4191 4771
rect 4187 4765 4191 4766
rect 4259 4770 4263 4771
rect 4259 4765 4263 4766
rect 4467 4770 4471 4771
rect 4467 4765 4471 4766
rect 4483 4770 4487 4771
rect 4483 4765 4487 4766
rect 4707 4770 4711 4771
rect 4707 4765 4711 4766
rect 4763 4770 4767 4771
rect 4763 4765 4767 4766
rect 4931 4770 4935 4771
rect 4931 4765 4935 4766
rect 5067 4770 5071 4771
rect 5067 4765 5071 4766
rect 3982 4755 3988 4756
rect 3982 4751 3983 4755
rect 3987 4751 3988 4755
rect 3982 4750 3988 4751
rect 4188 4704 4190 4765
rect 4194 4751 4200 4752
rect 4194 4747 4195 4751
rect 4199 4747 4200 4751
rect 4194 4746 4200 4747
rect 4196 4712 4198 4746
rect 4194 4711 4200 4712
rect 4194 4707 4195 4711
rect 4199 4707 4200 4711
rect 4194 4706 4200 4707
rect 4468 4704 4470 4765
rect 4474 4751 4480 4752
rect 4474 4747 4475 4751
rect 4479 4747 4480 4751
rect 4474 4746 4480 4747
rect 4476 4712 4478 4746
rect 4474 4711 4480 4712
rect 4474 4707 4475 4711
rect 4479 4707 4480 4711
rect 4474 4706 4480 4707
rect 4590 4711 4596 4712
rect 4590 4707 4591 4711
rect 4595 4707 4596 4711
rect 4590 4706 4596 4707
rect 3838 4700 3839 4704
rect 3843 4700 3844 4704
rect 3838 4699 3844 4700
rect 3914 4703 3920 4704
rect 3914 4699 3915 4703
rect 3919 4699 3920 4703
rect 3914 4698 3920 4699
rect 4186 4703 4192 4704
rect 4186 4699 4187 4703
rect 4191 4699 4192 4703
rect 4186 4698 4192 4699
rect 4466 4703 4472 4704
rect 4466 4699 4467 4703
rect 4471 4699 4472 4703
rect 4466 4698 4472 4699
rect 2919 4694 2923 4695
rect 2919 4689 2923 4690
rect 2959 4694 2963 4695
rect 2959 4689 2963 4690
rect 3143 4694 3147 4695
rect 3143 4689 3147 4690
rect 3159 4694 3163 4695
rect 3159 4689 3163 4690
rect 3367 4694 3371 4695
rect 3367 4689 3371 4690
rect 3799 4694 3803 4695
rect 3799 4689 3803 4690
rect 2920 4665 2922 4689
rect 3144 4665 3146 4689
rect 3368 4665 3370 4689
rect 3800 4666 3802 4689
rect 3942 4688 3948 4689
rect 3838 4687 3844 4688
rect 3838 4683 3839 4687
rect 3843 4683 3844 4687
rect 3942 4684 3943 4688
rect 3947 4684 3948 4688
rect 3942 4683 3948 4684
rect 4214 4688 4220 4689
rect 4214 4684 4215 4688
rect 4219 4684 4220 4688
rect 4214 4683 4220 4684
rect 4494 4688 4500 4689
rect 4494 4684 4495 4688
rect 4499 4684 4500 4688
rect 4494 4683 4500 4684
rect 3838 4682 3844 4683
rect 3798 4665 3804 4666
rect 2918 4664 2924 4665
rect 2918 4660 2919 4664
rect 2923 4660 2924 4664
rect 2918 4659 2924 4660
rect 3142 4664 3148 4665
rect 3142 4660 3143 4664
rect 3147 4660 3148 4664
rect 3142 4659 3148 4660
rect 3366 4664 3372 4665
rect 3366 4660 3367 4664
rect 3371 4660 3372 4664
rect 3798 4661 3799 4665
rect 3803 4661 3804 4665
rect 3798 4660 3804 4661
rect 3366 4659 3372 4660
rect 3840 4659 3842 4682
rect 3944 4659 3946 4683
rect 4216 4659 4218 4683
rect 4496 4659 4498 4683
rect 3839 4658 3843 4659
rect 3839 4653 3843 4654
rect 3943 4658 3947 4659
rect 3943 4653 3947 4654
rect 4063 4658 4067 4659
rect 4063 4653 4067 4654
rect 4215 4658 4219 4659
rect 4215 4653 4219 4654
rect 4327 4658 4331 4659
rect 4327 4653 4331 4654
rect 4495 4658 4499 4659
rect 4495 4653 4499 4654
rect 2890 4649 2896 4650
rect 2890 4645 2891 4649
rect 2895 4645 2896 4649
rect 2890 4644 2896 4645
rect 3114 4649 3120 4650
rect 3114 4645 3115 4649
rect 3119 4645 3120 4649
rect 3114 4644 3120 4645
rect 3338 4649 3344 4650
rect 3338 4645 3339 4649
rect 3343 4645 3344 4649
rect 3338 4644 3344 4645
rect 3798 4648 3804 4649
rect 3798 4644 3799 4648
rect 3803 4644 3804 4648
rect 2790 4639 2796 4640
rect 2790 4635 2791 4639
rect 2795 4635 2796 4639
rect 2790 4634 2796 4635
rect 2882 4639 2888 4640
rect 2882 4635 2883 4639
rect 2887 4635 2888 4639
rect 2882 4634 2888 4635
rect 2884 4600 2886 4634
rect 2882 4599 2888 4600
rect 2882 4595 2883 4599
rect 2887 4595 2888 4599
rect 2882 4594 2888 4595
rect 2892 4579 2894 4644
rect 2986 4631 2992 4632
rect 2986 4627 2987 4631
rect 2991 4627 2992 4631
rect 2986 4626 2992 4627
rect 2988 4600 2990 4626
rect 2986 4599 2992 4600
rect 2986 4595 2987 4599
rect 2991 4595 2992 4599
rect 2986 4594 2992 4595
rect 3116 4579 3118 4644
rect 3242 4639 3248 4640
rect 3242 4635 3243 4639
rect 3247 4635 3248 4639
rect 3242 4634 3248 4635
rect 3244 4600 3246 4634
rect 3126 4599 3132 4600
rect 3126 4595 3127 4599
rect 3131 4595 3132 4599
rect 3126 4594 3132 4595
rect 3242 4599 3248 4600
rect 3242 4595 3243 4599
rect 3247 4595 3248 4599
rect 3242 4594 3248 4595
rect 1975 4578 1979 4579
rect 1975 4573 1979 4574
rect 1995 4578 1999 4579
rect 1995 4573 1999 4574
rect 2099 4578 2103 4579
rect 2099 4573 2103 4574
rect 2211 4578 2215 4579
rect 2211 4573 2215 4574
rect 2347 4578 2351 4579
rect 2347 4573 2351 4574
rect 2443 4578 2447 4579
rect 2443 4573 2447 4574
rect 2579 4578 2583 4579
rect 2579 4573 2583 4574
rect 2667 4578 2671 4579
rect 2667 4573 2671 4574
rect 2795 4578 2799 4579
rect 2795 4573 2799 4574
rect 2891 4578 2895 4579
rect 2891 4573 2895 4574
rect 3003 4578 3007 4579
rect 3003 4573 3007 4574
rect 3115 4578 3119 4579
rect 3115 4573 3119 4574
rect 1934 4548 1940 4549
rect 1934 4544 1935 4548
rect 1939 4544 1940 4548
rect 1934 4543 1940 4544
rect 1814 4532 1820 4533
rect 1814 4528 1815 4532
rect 1819 4528 1820 4532
rect 1814 4527 1820 4528
rect 1934 4531 1940 4532
rect 1934 4527 1935 4531
rect 1939 4527 1940 4531
rect 1816 4499 1818 4527
rect 1934 4526 1940 4527
rect 1936 4499 1938 4526
rect 1976 4513 1978 4573
rect 1974 4512 1980 4513
rect 2100 4512 2102 4573
rect 2222 4519 2228 4520
rect 2222 4515 2223 4519
rect 2227 4515 2228 4519
rect 2222 4514 2228 4515
rect 1974 4508 1975 4512
rect 1979 4508 1980 4512
rect 1974 4507 1980 4508
rect 2098 4511 2104 4512
rect 2098 4507 2099 4511
rect 2103 4507 2104 4511
rect 2098 4506 2104 4507
rect 1815 4498 1819 4499
rect 1815 4493 1819 4494
rect 1935 4498 1939 4499
rect 2126 4496 2132 4497
rect 1935 4493 1939 4494
rect 1974 4495 1980 4496
rect 1936 4470 1938 4493
rect 1974 4491 1975 4495
rect 1979 4491 1980 4495
rect 2126 4492 2127 4496
rect 2131 4492 2132 4496
rect 2126 4491 2132 4492
rect 1974 4490 1980 4491
rect 1934 4469 1940 4470
rect 1934 4465 1935 4469
rect 1939 4465 1940 4469
rect 1934 4464 1940 4465
rect 1976 4459 1978 4490
rect 2128 4459 2130 4491
rect 1975 4458 1979 4459
rect 1975 4453 1979 4454
rect 2127 4458 2131 4459
rect 2127 4453 2131 4454
rect 1934 4452 1940 4453
rect 1934 4448 1935 4452
rect 1939 4448 1940 4452
rect 1934 4447 1940 4448
rect 1794 4443 1800 4444
rect 1794 4439 1795 4443
rect 1799 4439 1800 4443
rect 1794 4438 1800 4439
rect 1746 4403 1752 4404
rect 1746 4399 1747 4403
rect 1751 4399 1752 4403
rect 1746 4398 1752 4399
rect 1291 4382 1295 4383
rect 1291 4377 1295 4378
rect 1379 4382 1383 4383
rect 1379 4377 1383 4378
rect 1467 4382 1471 4383
rect 1467 4377 1471 4378
rect 1651 4382 1655 4383
rect 1651 4377 1655 4378
rect 1274 4371 1280 4372
rect 1274 4367 1275 4371
rect 1279 4367 1280 4371
rect 1274 4366 1280 4367
rect 1130 4363 1136 4364
rect 1130 4359 1131 4363
rect 1135 4359 1136 4363
rect 1130 4358 1136 4359
rect 1132 4324 1134 4358
rect 1130 4323 1136 4324
rect 1130 4319 1131 4323
rect 1135 4319 1136 4323
rect 1130 4318 1136 4319
rect 1292 4316 1294 4377
rect 1298 4363 1304 4364
rect 1298 4359 1299 4363
rect 1303 4359 1304 4363
rect 1298 4358 1304 4359
rect 1300 4324 1302 4358
rect 1298 4323 1304 4324
rect 1298 4319 1299 4323
rect 1303 4319 1304 4323
rect 1298 4318 1304 4319
rect 1306 4323 1312 4324
rect 1306 4319 1307 4323
rect 1311 4319 1312 4323
rect 1306 4318 1312 4319
rect 110 4312 111 4316
rect 115 4312 116 4316
rect 110 4311 116 4312
rect 666 4315 672 4316
rect 666 4311 667 4315
rect 671 4311 672 4315
rect 666 4310 672 4311
rect 810 4315 816 4316
rect 810 4311 811 4315
rect 815 4311 816 4315
rect 810 4310 816 4311
rect 962 4315 968 4316
rect 962 4311 963 4315
rect 967 4311 968 4315
rect 962 4310 968 4311
rect 1122 4315 1128 4316
rect 1122 4311 1123 4315
rect 1127 4311 1128 4315
rect 1122 4310 1128 4311
rect 1290 4315 1296 4316
rect 1290 4311 1291 4315
rect 1295 4311 1296 4315
rect 1290 4310 1296 4311
rect 694 4300 700 4301
rect 110 4299 116 4300
rect 110 4295 111 4299
rect 115 4295 116 4299
rect 694 4296 695 4300
rect 699 4296 700 4300
rect 694 4295 700 4296
rect 838 4300 844 4301
rect 838 4296 839 4300
rect 843 4296 844 4300
rect 838 4295 844 4296
rect 990 4300 996 4301
rect 990 4296 991 4300
rect 995 4296 996 4300
rect 990 4295 996 4296
rect 1150 4300 1156 4301
rect 1150 4296 1151 4300
rect 1155 4296 1156 4300
rect 1150 4295 1156 4296
rect 110 4294 116 4295
rect 112 4255 114 4294
rect 696 4255 698 4295
rect 840 4255 842 4295
rect 992 4255 994 4295
rect 1152 4255 1154 4295
rect 111 4254 115 4255
rect 111 4249 115 4250
rect 695 4254 699 4255
rect 695 4249 699 4250
rect 815 4254 819 4255
rect 815 4249 819 4250
rect 839 4254 843 4255
rect 839 4249 843 4250
rect 951 4254 955 4255
rect 951 4249 955 4250
rect 991 4254 995 4255
rect 991 4249 995 4250
rect 1087 4254 1091 4255
rect 1087 4249 1091 4250
rect 1151 4254 1155 4255
rect 1151 4249 1155 4250
rect 1223 4254 1227 4255
rect 1223 4249 1227 4250
rect 112 4226 114 4249
rect 110 4225 116 4226
rect 816 4225 818 4249
rect 952 4225 954 4249
rect 1088 4225 1090 4249
rect 1224 4225 1226 4249
rect 110 4221 111 4225
rect 115 4221 116 4225
rect 110 4220 116 4221
rect 814 4224 820 4225
rect 814 4220 815 4224
rect 819 4220 820 4224
rect 814 4219 820 4220
rect 950 4224 956 4225
rect 950 4220 951 4224
rect 955 4220 956 4224
rect 950 4219 956 4220
rect 1086 4224 1092 4225
rect 1086 4220 1087 4224
rect 1091 4220 1092 4224
rect 1086 4219 1092 4220
rect 1222 4224 1228 4225
rect 1222 4220 1223 4224
rect 1227 4220 1228 4224
rect 1222 4219 1228 4220
rect 786 4209 792 4210
rect 110 4208 116 4209
rect 110 4204 111 4208
rect 115 4204 116 4208
rect 786 4205 787 4209
rect 791 4205 792 4209
rect 786 4204 792 4205
rect 922 4209 928 4210
rect 922 4205 923 4209
rect 927 4205 928 4209
rect 922 4204 928 4205
rect 1058 4209 1064 4210
rect 1058 4205 1059 4209
rect 1063 4205 1064 4209
rect 1058 4204 1064 4205
rect 1194 4209 1200 4210
rect 1194 4205 1195 4209
rect 1199 4205 1200 4209
rect 1194 4204 1200 4205
rect 110 4203 116 4204
rect 112 4139 114 4203
rect 788 4139 790 4204
rect 914 4199 920 4200
rect 914 4195 915 4199
rect 919 4195 920 4199
rect 914 4194 920 4195
rect 916 4160 918 4194
rect 914 4159 920 4160
rect 914 4155 915 4159
rect 919 4155 920 4159
rect 914 4154 920 4155
rect 924 4139 926 4204
rect 1050 4199 1056 4200
rect 1050 4195 1051 4199
rect 1055 4195 1056 4199
rect 1050 4194 1056 4195
rect 1052 4160 1054 4194
rect 1050 4159 1056 4160
rect 1050 4155 1051 4159
rect 1055 4155 1056 4159
rect 1050 4154 1056 4155
rect 1060 4139 1062 4204
rect 1186 4199 1192 4200
rect 1186 4195 1187 4199
rect 1191 4195 1192 4199
rect 1186 4194 1192 4195
rect 1188 4160 1190 4194
rect 1186 4159 1192 4160
rect 1186 4155 1187 4159
rect 1191 4155 1192 4159
rect 1186 4154 1192 4155
rect 1196 4139 1198 4204
rect 1308 4152 1310 4318
rect 1468 4316 1470 4377
rect 1562 4363 1568 4364
rect 1562 4359 1563 4363
rect 1567 4359 1568 4363
rect 1562 4358 1568 4359
rect 1466 4315 1472 4316
rect 1466 4311 1467 4315
rect 1471 4311 1472 4315
rect 1466 4310 1472 4311
rect 1318 4300 1324 4301
rect 1318 4296 1319 4300
rect 1323 4296 1324 4300
rect 1318 4295 1324 4296
rect 1494 4300 1500 4301
rect 1494 4296 1495 4300
rect 1499 4296 1500 4300
rect 1494 4295 1500 4296
rect 1320 4255 1322 4295
rect 1496 4255 1498 4295
rect 1319 4254 1323 4255
rect 1319 4249 1323 4250
rect 1359 4254 1363 4255
rect 1359 4249 1363 4250
rect 1495 4254 1499 4255
rect 1495 4249 1499 4250
rect 1360 4225 1362 4249
rect 1496 4225 1498 4249
rect 1358 4224 1364 4225
rect 1358 4220 1359 4224
rect 1363 4220 1364 4224
rect 1358 4219 1364 4220
rect 1494 4224 1500 4225
rect 1494 4220 1495 4224
rect 1499 4220 1500 4224
rect 1494 4219 1500 4220
rect 1330 4209 1336 4210
rect 1330 4205 1331 4209
rect 1335 4205 1336 4209
rect 1330 4204 1336 4205
rect 1466 4209 1472 4210
rect 1466 4205 1467 4209
rect 1471 4205 1472 4209
rect 1466 4204 1472 4205
rect 1322 4199 1328 4200
rect 1322 4195 1323 4199
rect 1327 4195 1328 4199
rect 1322 4194 1328 4195
rect 1324 4160 1326 4194
rect 1322 4159 1328 4160
rect 1322 4155 1323 4159
rect 1327 4155 1328 4159
rect 1322 4154 1328 4155
rect 1306 4151 1312 4152
rect 1306 4147 1307 4151
rect 1311 4147 1312 4151
rect 1306 4146 1312 4147
rect 1332 4139 1334 4204
rect 1378 4199 1384 4200
rect 1378 4195 1379 4199
rect 1383 4195 1384 4199
rect 1378 4194 1384 4195
rect 111 4138 115 4139
rect 111 4133 115 4134
rect 731 4138 735 4139
rect 731 4133 735 4134
rect 787 4138 791 4139
rect 787 4133 791 4134
rect 867 4138 871 4139
rect 867 4133 871 4134
rect 923 4138 927 4139
rect 923 4133 927 4134
rect 1003 4138 1007 4139
rect 1003 4133 1007 4134
rect 1059 4138 1063 4139
rect 1059 4133 1063 4134
rect 1139 4138 1143 4139
rect 1139 4133 1143 4134
rect 1195 4138 1199 4139
rect 1195 4133 1199 4134
rect 1275 4138 1279 4139
rect 1275 4133 1279 4134
rect 1331 4138 1335 4139
rect 1331 4133 1335 4134
rect 112 4073 114 4133
rect 110 4072 116 4073
rect 732 4072 734 4133
rect 854 4079 860 4080
rect 854 4075 855 4079
rect 859 4075 860 4079
rect 854 4074 860 4075
rect 110 4068 111 4072
rect 115 4068 116 4072
rect 110 4067 116 4068
rect 730 4071 736 4072
rect 730 4067 731 4071
rect 735 4067 736 4071
rect 730 4066 736 4067
rect 758 4056 764 4057
rect 110 4055 116 4056
rect 110 4051 111 4055
rect 115 4051 116 4055
rect 758 4052 759 4056
rect 763 4052 764 4056
rect 758 4051 764 4052
rect 110 4050 116 4051
rect 112 4003 114 4050
rect 760 4003 762 4051
rect 111 4002 115 4003
rect 111 3997 115 3998
rect 511 4002 515 4003
rect 511 3997 515 3998
rect 663 4002 667 4003
rect 663 3997 667 3998
rect 759 4002 763 4003
rect 759 3997 763 3998
rect 823 4002 827 4003
rect 823 3997 827 3998
rect 112 3974 114 3997
rect 110 3973 116 3974
rect 512 3973 514 3997
rect 664 3973 666 3997
rect 824 3973 826 3997
rect 110 3969 111 3973
rect 115 3969 116 3973
rect 110 3968 116 3969
rect 510 3972 516 3973
rect 510 3968 511 3972
rect 515 3968 516 3972
rect 510 3967 516 3968
rect 662 3972 668 3973
rect 662 3968 663 3972
rect 667 3968 668 3972
rect 662 3967 668 3968
rect 822 3972 828 3973
rect 822 3968 823 3972
rect 827 3968 828 3972
rect 822 3967 828 3968
rect 482 3957 488 3958
rect 110 3956 116 3957
rect 110 3952 111 3956
rect 115 3952 116 3956
rect 482 3953 483 3957
rect 487 3953 488 3957
rect 482 3952 488 3953
rect 634 3957 640 3958
rect 634 3953 635 3957
rect 639 3953 640 3957
rect 634 3952 640 3953
rect 794 3957 800 3958
rect 794 3953 795 3957
rect 799 3953 800 3957
rect 794 3952 800 3953
rect 110 3951 116 3952
rect 112 3863 114 3951
rect 484 3863 486 3952
rect 610 3947 616 3948
rect 610 3943 611 3947
rect 615 3943 616 3947
rect 610 3942 616 3943
rect 578 3939 584 3940
rect 578 3935 579 3939
rect 583 3935 584 3939
rect 578 3934 584 3935
rect 580 3908 582 3934
rect 612 3908 614 3942
rect 578 3907 584 3908
rect 578 3903 579 3907
rect 583 3903 584 3907
rect 578 3902 584 3903
rect 610 3907 616 3908
rect 610 3903 611 3907
rect 615 3903 616 3907
rect 610 3902 616 3903
rect 636 3863 638 3952
rect 758 3947 764 3948
rect 758 3943 759 3947
rect 763 3943 764 3947
rect 758 3942 764 3943
rect 111 3862 115 3863
rect 111 3857 115 3858
rect 131 3862 135 3863
rect 131 3857 135 3858
rect 307 3862 311 3863
rect 307 3857 311 3858
rect 483 3862 487 3863
rect 483 3857 487 3858
rect 515 3862 519 3863
rect 515 3857 519 3858
rect 635 3862 639 3863
rect 635 3857 639 3858
rect 723 3862 727 3863
rect 723 3857 727 3858
rect 112 3797 114 3857
rect 110 3796 116 3797
rect 132 3796 134 3857
rect 308 3796 310 3857
rect 314 3843 320 3844
rect 314 3839 315 3843
rect 319 3839 320 3843
rect 314 3838 320 3839
rect 316 3804 318 3838
rect 314 3803 320 3804
rect 314 3799 315 3803
rect 319 3799 320 3803
rect 314 3798 320 3799
rect 402 3803 408 3804
rect 402 3799 403 3803
rect 407 3799 408 3803
rect 402 3798 408 3799
rect 110 3792 111 3796
rect 115 3792 116 3796
rect 110 3791 116 3792
rect 130 3795 136 3796
rect 130 3791 131 3795
rect 135 3791 136 3795
rect 130 3790 136 3791
rect 306 3795 312 3796
rect 306 3791 307 3795
rect 311 3791 312 3795
rect 306 3790 312 3791
rect 158 3780 164 3781
rect 110 3779 116 3780
rect 110 3775 111 3779
rect 115 3775 116 3779
rect 158 3776 159 3780
rect 163 3776 164 3780
rect 158 3775 164 3776
rect 334 3780 340 3781
rect 334 3776 335 3780
rect 339 3776 340 3780
rect 334 3775 340 3776
rect 110 3774 116 3775
rect 112 3751 114 3774
rect 160 3751 162 3775
rect 336 3751 338 3775
rect 111 3750 115 3751
rect 111 3745 115 3746
rect 159 3750 163 3751
rect 159 3745 163 3746
rect 335 3750 339 3751
rect 335 3745 339 3746
rect 112 3722 114 3745
rect 110 3721 116 3722
rect 160 3721 162 3745
rect 336 3721 338 3745
rect 110 3717 111 3721
rect 115 3717 116 3721
rect 110 3716 116 3717
rect 158 3720 164 3721
rect 158 3716 159 3720
rect 163 3716 164 3720
rect 158 3715 164 3716
rect 334 3720 340 3721
rect 334 3716 335 3720
rect 339 3716 340 3720
rect 334 3715 340 3716
rect 130 3705 136 3706
rect 110 3704 116 3705
rect 110 3700 111 3704
rect 115 3700 116 3704
rect 130 3701 131 3705
rect 135 3701 136 3705
rect 130 3700 136 3701
rect 306 3705 312 3706
rect 306 3701 307 3705
rect 311 3701 312 3705
rect 306 3700 312 3701
rect 110 3699 116 3700
rect 112 3627 114 3699
rect 132 3627 134 3700
rect 242 3695 248 3696
rect 242 3691 243 3695
rect 247 3691 248 3695
rect 242 3690 248 3691
rect 226 3687 232 3688
rect 226 3683 227 3687
rect 231 3683 232 3687
rect 226 3682 232 3683
rect 228 3656 230 3682
rect 226 3655 232 3656
rect 226 3651 227 3655
rect 231 3651 232 3655
rect 226 3650 232 3651
rect 111 3626 115 3627
rect 111 3621 115 3622
rect 131 3626 135 3627
rect 131 3621 135 3622
rect 147 3626 151 3627
rect 147 3621 151 3622
rect 112 3561 114 3621
rect 110 3560 116 3561
rect 148 3560 150 3621
rect 244 3612 246 3690
rect 308 3627 310 3700
rect 404 3656 406 3798
rect 516 3796 518 3857
rect 626 3855 632 3856
rect 626 3851 627 3855
rect 631 3851 632 3855
rect 626 3850 632 3851
rect 628 3804 630 3850
rect 626 3803 632 3804
rect 626 3799 627 3803
rect 631 3799 632 3803
rect 626 3798 632 3799
rect 724 3796 726 3857
rect 760 3848 762 3942
rect 796 3863 798 3952
rect 856 3908 858 4074
rect 868 4072 870 4133
rect 1004 4072 1006 4133
rect 1098 4119 1104 4120
rect 1098 4115 1099 4119
rect 1103 4115 1104 4119
rect 1098 4114 1104 4115
rect 1100 4088 1102 4114
rect 1098 4087 1104 4088
rect 1098 4083 1099 4087
rect 1103 4083 1104 4087
rect 1098 4082 1104 4083
rect 1140 4072 1142 4133
rect 1276 4072 1278 4133
rect 1380 4128 1382 4194
rect 1468 4139 1470 4204
rect 1564 4200 1566 4358
rect 1652 4316 1654 4377
rect 1658 4363 1664 4364
rect 1658 4359 1659 4363
rect 1663 4359 1664 4363
rect 1658 4358 1664 4359
rect 1660 4324 1662 4358
rect 1748 4324 1750 4398
rect 1936 4383 1938 4447
rect 1976 4430 1978 4453
rect 1974 4429 1980 4430
rect 1974 4425 1975 4429
rect 1979 4425 1980 4429
rect 1974 4424 1980 4425
rect 2202 4413 2208 4414
rect 1974 4412 1980 4413
rect 1974 4408 1975 4412
rect 1979 4408 1980 4412
rect 2202 4409 2203 4413
rect 2207 4409 2208 4413
rect 2202 4408 2208 4409
rect 1974 4407 1980 4408
rect 1935 4382 1939 4383
rect 1935 4377 1939 4378
rect 1658 4323 1664 4324
rect 1658 4319 1659 4323
rect 1663 4319 1664 4323
rect 1658 4318 1664 4319
rect 1746 4323 1752 4324
rect 1746 4319 1747 4323
rect 1751 4319 1752 4323
rect 1746 4318 1752 4319
rect 1936 4317 1938 4377
rect 1976 4339 1978 4407
rect 2204 4339 2206 4408
rect 2224 4364 2226 4514
rect 2348 4512 2350 4573
rect 2580 4512 2582 4573
rect 2796 4512 2798 4573
rect 2890 4559 2896 4560
rect 2890 4555 2891 4559
rect 2895 4555 2896 4559
rect 2890 4554 2896 4555
rect 2892 4528 2894 4554
rect 2890 4527 2896 4528
rect 2890 4523 2891 4527
rect 2895 4523 2896 4527
rect 2890 4522 2896 4523
rect 3004 4512 3006 4573
rect 3010 4559 3016 4560
rect 3010 4555 3011 4559
rect 3015 4555 3016 4559
rect 3010 4554 3016 4555
rect 3012 4520 3014 4554
rect 3128 4520 3130 4594
rect 3340 4579 3342 4644
rect 3798 4643 3804 4644
rect 3800 4579 3802 4643
rect 3840 4630 3842 4653
rect 3838 4629 3844 4630
rect 4064 4629 4066 4653
rect 4328 4629 4330 4653
rect 3838 4625 3839 4629
rect 3843 4625 3844 4629
rect 3838 4624 3844 4625
rect 4062 4628 4068 4629
rect 4062 4624 4063 4628
rect 4067 4624 4068 4628
rect 4062 4623 4068 4624
rect 4326 4628 4332 4629
rect 4326 4624 4327 4628
rect 4331 4624 4332 4628
rect 4326 4623 4332 4624
rect 4034 4613 4040 4614
rect 3838 4612 3844 4613
rect 3838 4608 3839 4612
rect 3843 4608 3844 4612
rect 4034 4609 4035 4613
rect 4039 4609 4040 4613
rect 4034 4608 4040 4609
rect 4298 4613 4304 4614
rect 4298 4609 4299 4613
rect 4303 4609 4304 4613
rect 4298 4608 4304 4609
rect 4570 4613 4576 4614
rect 4570 4609 4571 4613
rect 4575 4609 4576 4613
rect 4570 4608 4576 4609
rect 3838 4607 3844 4608
rect 3203 4578 3207 4579
rect 3203 4573 3207 4574
rect 3339 4578 3343 4579
rect 3339 4573 3343 4574
rect 3403 4578 3407 4579
rect 3403 4573 3407 4574
rect 3611 4578 3615 4579
rect 3611 4573 3615 4574
rect 3799 4578 3803 4579
rect 3799 4573 3803 4574
rect 3010 4519 3016 4520
rect 3010 4515 3011 4519
rect 3015 4515 3016 4519
rect 3010 4514 3016 4515
rect 3126 4519 3132 4520
rect 3126 4515 3127 4519
rect 3131 4515 3132 4519
rect 3126 4514 3132 4515
rect 3204 4512 3206 4573
rect 3404 4512 3406 4573
rect 3612 4512 3614 4573
rect 3706 4559 3712 4560
rect 3706 4555 3707 4559
rect 3711 4555 3712 4559
rect 3706 4554 3712 4555
rect 2346 4511 2352 4512
rect 2346 4507 2347 4511
rect 2351 4507 2352 4511
rect 2346 4506 2352 4507
rect 2578 4511 2584 4512
rect 2578 4507 2579 4511
rect 2583 4507 2584 4511
rect 2578 4506 2584 4507
rect 2794 4511 2800 4512
rect 2794 4507 2795 4511
rect 2799 4507 2800 4511
rect 2794 4506 2800 4507
rect 3002 4511 3008 4512
rect 3002 4507 3003 4511
rect 3007 4507 3008 4511
rect 3002 4506 3008 4507
rect 3202 4511 3208 4512
rect 3202 4507 3203 4511
rect 3207 4507 3208 4511
rect 3202 4506 3208 4507
rect 3402 4511 3408 4512
rect 3402 4507 3403 4511
rect 3407 4507 3408 4511
rect 3402 4506 3408 4507
rect 3610 4511 3616 4512
rect 3610 4507 3611 4511
rect 3615 4507 3616 4511
rect 3610 4506 3616 4507
rect 2374 4496 2380 4497
rect 2374 4492 2375 4496
rect 2379 4492 2380 4496
rect 2374 4491 2380 4492
rect 2606 4496 2612 4497
rect 2606 4492 2607 4496
rect 2611 4492 2612 4496
rect 2606 4491 2612 4492
rect 2822 4496 2828 4497
rect 2822 4492 2823 4496
rect 2827 4492 2828 4496
rect 2822 4491 2828 4492
rect 3030 4496 3036 4497
rect 3030 4492 3031 4496
rect 3035 4492 3036 4496
rect 3030 4491 3036 4492
rect 3230 4496 3236 4497
rect 3230 4492 3231 4496
rect 3235 4492 3236 4496
rect 3230 4491 3236 4492
rect 3430 4496 3436 4497
rect 3430 4492 3431 4496
rect 3435 4492 3436 4496
rect 3430 4491 3436 4492
rect 3638 4496 3644 4497
rect 3638 4492 3639 4496
rect 3643 4492 3644 4496
rect 3638 4491 3644 4492
rect 2376 4459 2378 4491
rect 2608 4459 2610 4491
rect 2824 4459 2826 4491
rect 3032 4459 3034 4491
rect 3232 4459 3234 4491
rect 3432 4459 3434 4491
rect 3640 4459 3642 4491
rect 2231 4458 2235 4459
rect 2231 4453 2235 4454
rect 2375 4458 2379 4459
rect 2375 4453 2379 4454
rect 2447 4458 2451 4459
rect 2447 4453 2451 4454
rect 2607 4458 2611 4459
rect 2607 4453 2611 4454
rect 2663 4458 2667 4459
rect 2663 4453 2667 4454
rect 2823 4458 2827 4459
rect 2823 4453 2827 4454
rect 2871 4458 2875 4459
rect 2871 4453 2875 4454
rect 3031 4458 3035 4459
rect 3031 4453 3035 4454
rect 3079 4458 3083 4459
rect 3079 4453 3083 4454
rect 3231 4458 3235 4459
rect 3231 4453 3235 4454
rect 3287 4458 3291 4459
rect 3287 4453 3291 4454
rect 3431 4458 3435 4459
rect 3431 4453 3435 4454
rect 3495 4458 3499 4459
rect 3495 4453 3499 4454
rect 3639 4458 3643 4459
rect 3639 4453 3643 4454
rect 3679 4458 3683 4459
rect 3679 4453 3683 4454
rect 2232 4429 2234 4453
rect 2448 4429 2450 4453
rect 2664 4429 2666 4453
rect 2872 4429 2874 4453
rect 3080 4429 3082 4453
rect 3288 4429 3290 4453
rect 3496 4429 3498 4453
rect 3680 4429 3682 4453
rect 2230 4428 2236 4429
rect 2230 4424 2231 4428
rect 2235 4424 2236 4428
rect 2230 4423 2236 4424
rect 2446 4428 2452 4429
rect 2446 4424 2447 4428
rect 2451 4424 2452 4428
rect 2446 4423 2452 4424
rect 2662 4428 2668 4429
rect 2662 4424 2663 4428
rect 2667 4424 2668 4428
rect 2662 4423 2668 4424
rect 2870 4428 2876 4429
rect 2870 4424 2871 4428
rect 2875 4424 2876 4428
rect 2870 4423 2876 4424
rect 3078 4428 3084 4429
rect 3078 4424 3079 4428
rect 3083 4424 3084 4428
rect 3078 4423 3084 4424
rect 3286 4428 3292 4429
rect 3286 4424 3287 4428
rect 3291 4424 3292 4428
rect 3286 4423 3292 4424
rect 3494 4428 3500 4429
rect 3494 4424 3495 4428
rect 3499 4424 3500 4428
rect 3494 4423 3500 4424
rect 3678 4428 3684 4429
rect 3678 4424 3679 4428
rect 3683 4424 3684 4428
rect 3678 4423 3684 4424
rect 2418 4413 2424 4414
rect 2418 4409 2419 4413
rect 2423 4409 2424 4413
rect 2418 4408 2424 4409
rect 2634 4413 2640 4414
rect 2634 4409 2635 4413
rect 2639 4409 2640 4413
rect 2634 4408 2640 4409
rect 2842 4413 2848 4414
rect 2842 4409 2843 4413
rect 2847 4409 2848 4413
rect 2842 4408 2848 4409
rect 3050 4413 3056 4414
rect 3050 4409 3051 4413
rect 3055 4409 3056 4413
rect 3050 4408 3056 4409
rect 3258 4413 3264 4414
rect 3258 4409 3259 4413
rect 3263 4409 3264 4413
rect 3258 4408 3264 4409
rect 3466 4413 3472 4414
rect 3466 4409 3467 4413
rect 3471 4409 3472 4413
rect 3466 4408 3472 4409
rect 3650 4413 3656 4414
rect 3650 4409 3651 4413
rect 3655 4409 3656 4413
rect 3650 4408 3656 4409
rect 2330 4403 2336 4404
rect 2330 4399 2331 4403
rect 2335 4399 2336 4403
rect 2330 4398 2336 4399
rect 2332 4364 2334 4398
rect 2222 4363 2228 4364
rect 2222 4359 2223 4363
rect 2227 4359 2228 4363
rect 2222 4358 2228 4359
rect 2330 4363 2336 4364
rect 2330 4359 2331 4363
rect 2335 4359 2336 4363
rect 2330 4358 2336 4359
rect 2420 4339 2422 4408
rect 2546 4403 2552 4404
rect 2546 4399 2547 4403
rect 2551 4399 2552 4403
rect 2546 4398 2552 4399
rect 2548 4364 2550 4398
rect 2546 4363 2552 4364
rect 2546 4359 2547 4363
rect 2551 4359 2552 4363
rect 2546 4358 2552 4359
rect 2636 4339 2638 4408
rect 2786 4403 2792 4404
rect 2786 4399 2787 4403
rect 2791 4399 2792 4403
rect 2786 4398 2792 4399
rect 2788 4364 2790 4398
rect 2786 4363 2792 4364
rect 2786 4359 2787 4363
rect 2791 4359 2792 4363
rect 2786 4358 2792 4359
rect 2844 4339 2846 4408
rect 2914 4403 2920 4404
rect 2914 4399 2915 4403
rect 2919 4399 2920 4403
rect 2914 4398 2920 4399
rect 1975 4338 1979 4339
rect 1975 4333 1979 4334
rect 2203 4338 2207 4339
rect 2203 4333 2207 4334
rect 2307 4338 2311 4339
rect 2307 4333 2311 4334
rect 2419 4338 2423 4339
rect 2419 4333 2423 4334
rect 2459 4338 2463 4339
rect 2459 4333 2463 4334
rect 2627 4338 2631 4339
rect 2627 4333 2631 4334
rect 2635 4338 2639 4339
rect 2635 4333 2639 4334
rect 2811 4338 2815 4339
rect 2811 4333 2815 4334
rect 2843 4338 2847 4339
rect 2843 4333 2847 4334
rect 1934 4316 1940 4317
rect 1650 4315 1656 4316
rect 1650 4311 1651 4315
rect 1655 4311 1656 4315
rect 1934 4312 1935 4316
rect 1939 4312 1940 4316
rect 1934 4311 1940 4312
rect 1650 4310 1656 4311
rect 1678 4300 1684 4301
rect 1678 4296 1679 4300
rect 1683 4296 1684 4300
rect 1678 4295 1684 4296
rect 1934 4299 1940 4300
rect 1934 4295 1935 4299
rect 1939 4295 1940 4299
rect 1680 4255 1682 4295
rect 1934 4294 1940 4295
rect 1936 4255 1938 4294
rect 1976 4273 1978 4333
rect 1974 4272 1980 4273
rect 2308 4272 2310 4333
rect 2460 4272 2462 4333
rect 2466 4319 2472 4320
rect 2466 4315 2467 4319
rect 2471 4315 2472 4319
rect 2466 4314 2472 4315
rect 2468 4280 2470 4314
rect 2466 4279 2472 4280
rect 2466 4275 2467 4279
rect 2471 4275 2472 4279
rect 2466 4274 2472 4275
rect 2628 4272 2630 4333
rect 2634 4319 2640 4320
rect 2634 4315 2635 4319
rect 2639 4315 2640 4319
rect 2634 4314 2640 4315
rect 2636 4280 2638 4314
rect 2634 4279 2640 4280
rect 2634 4275 2635 4279
rect 2639 4275 2640 4279
rect 2634 4274 2640 4275
rect 2812 4272 2814 4333
rect 2916 4328 2918 4398
rect 3052 4339 3054 4408
rect 3190 4403 3196 4404
rect 3190 4399 3191 4403
rect 3195 4399 3196 4403
rect 3190 4398 3196 4399
rect 3192 4364 3194 4398
rect 3190 4363 3196 4364
rect 3190 4359 3191 4363
rect 3195 4359 3196 4363
rect 3190 4358 3196 4359
rect 3260 4339 3262 4408
rect 3430 4403 3436 4404
rect 3430 4399 3431 4403
rect 3435 4399 3436 4403
rect 3430 4398 3436 4399
rect 3432 4364 3434 4398
rect 3430 4363 3436 4364
rect 3430 4359 3431 4363
rect 3435 4359 3436 4363
rect 3430 4358 3436 4359
rect 3438 4355 3444 4356
rect 3438 4351 3439 4355
rect 3443 4351 3444 4355
rect 3438 4350 3444 4351
rect 3011 4338 3015 4339
rect 3011 4333 3015 4334
rect 3051 4338 3055 4339
rect 3051 4333 3055 4334
rect 3227 4338 3231 4339
rect 3227 4333 3231 4334
rect 3259 4338 3263 4339
rect 3259 4333 3263 4334
rect 2914 4327 2920 4328
rect 2914 4323 2915 4327
rect 2919 4323 2920 4327
rect 2914 4322 2920 4323
rect 2818 4319 2824 4320
rect 2818 4315 2819 4319
rect 2823 4315 2824 4319
rect 2818 4314 2824 4315
rect 2820 4280 2822 4314
rect 2818 4279 2824 4280
rect 2818 4275 2819 4279
rect 2823 4275 2824 4279
rect 2818 4274 2824 4275
rect 3012 4272 3014 4333
rect 3018 4319 3024 4320
rect 3018 4315 3019 4319
rect 3023 4315 3024 4319
rect 3018 4314 3024 4315
rect 3020 4280 3022 4314
rect 3018 4279 3024 4280
rect 3018 4275 3019 4279
rect 3023 4275 3024 4279
rect 3018 4274 3024 4275
rect 3228 4272 3230 4333
rect 3234 4319 3240 4320
rect 3234 4315 3235 4319
rect 3239 4315 3240 4319
rect 3234 4314 3240 4315
rect 3236 4280 3238 4314
rect 3440 4280 3442 4350
rect 3468 4339 3470 4408
rect 3606 4403 3612 4404
rect 3606 4399 3607 4403
rect 3611 4399 3612 4403
rect 3606 4398 3612 4399
rect 3608 4364 3610 4398
rect 3606 4363 3612 4364
rect 3606 4359 3607 4363
rect 3611 4359 3612 4363
rect 3606 4358 3612 4359
rect 3652 4339 3654 4408
rect 3708 4404 3710 4554
rect 3800 4513 3802 4573
rect 3840 4547 3842 4607
rect 4036 4547 4038 4608
rect 4170 4603 4176 4604
rect 4170 4599 4171 4603
rect 4175 4599 4176 4603
rect 4170 4598 4176 4599
rect 3839 4546 3843 4547
rect 3839 4541 3843 4542
rect 4035 4546 4039 4547
rect 4035 4541 4039 4542
rect 3798 4512 3804 4513
rect 3798 4508 3799 4512
rect 3803 4508 3804 4512
rect 3798 4507 3804 4508
rect 3798 4495 3804 4496
rect 3798 4491 3799 4495
rect 3803 4491 3804 4495
rect 3798 4490 3804 4491
rect 3800 4459 3802 4490
rect 3840 4481 3842 4541
rect 4172 4532 4174 4598
rect 4300 4547 4302 4608
rect 4542 4603 4548 4604
rect 4542 4599 4543 4603
rect 4547 4599 4548 4603
rect 4542 4598 4548 4599
rect 4544 4564 4546 4598
rect 4542 4563 4548 4564
rect 4542 4559 4543 4563
rect 4547 4559 4548 4563
rect 4542 4558 4548 4559
rect 4572 4547 4574 4608
rect 4592 4564 4594 4706
rect 4764 4704 4766 4765
rect 4858 4751 4864 4752
rect 4858 4747 4859 4751
rect 4863 4747 4864 4751
rect 4858 4746 4864 4747
rect 4762 4703 4768 4704
rect 4762 4699 4763 4703
rect 4767 4699 4768 4703
rect 4762 4698 4768 4699
rect 4790 4688 4796 4689
rect 4790 4684 4791 4688
rect 4795 4684 4796 4688
rect 4790 4683 4796 4684
rect 4792 4659 4794 4683
rect 4599 4658 4603 4659
rect 4599 4653 4603 4654
rect 4791 4658 4795 4659
rect 4791 4653 4795 4654
rect 4600 4629 4602 4653
rect 4598 4628 4604 4629
rect 4598 4624 4599 4628
rect 4603 4624 4604 4628
rect 4598 4623 4604 4624
rect 4842 4613 4848 4614
rect 4842 4609 4843 4613
rect 4847 4609 4848 4613
rect 4842 4608 4848 4609
rect 4590 4563 4596 4564
rect 4590 4559 4591 4563
rect 4595 4559 4596 4563
rect 4590 4558 4596 4559
rect 4844 4547 4846 4608
rect 4860 4604 4862 4746
rect 5068 4704 5070 4765
rect 5074 4751 5080 4752
rect 5074 4747 5075 4751
rect 5079 4747 5080 4751
rect 5074 4746 5080 4747
rect 5076 4712 5078 4746
rect 5084 4712 5086 4786
rect 5156 4771 5158 4836
rect 5192 4792 5194 4954
rect 5300 4952 5302 5013
rect 5336 5004 5338 5082
rect 5664 5019 5666 5091
rect 5663 5018 5667 5019
rect 5663 5013 5667 5014
rect 5334 5003 5340 5004
rect 5334 4999 5335 5003
rect 5339 4999 5340 5003
rect 5334 4998 5340 4999
rect 5664 4953 5666 5013
rect 5662 4952 5668 4953
rect 5298 4951 5304 4952
rect 5298 4947 5299 4951
rect 5303 4947 5304 4951
rect 5662 4948 5663 4952
rect 5667 4948 5668 4952
rect 5662 4947 5668 4948
rect 5298 4946 5304 4947
rect 5326 4936 5332 4937
rect 5326 4932 5327 4936
rect 5331 4932 5332 4936
rect 5326 4931 5332 4932
rect 5662 4935 5668 4936
rect 5662 4931 5663 4935
rect 5667 4931 5668 4935
rect 5328 4887 5330 4931
rect 5662 4930 5668 4931
rect 5664 4887 5666 4930
rect 5327 4886 5331 4887
rect 5327 4881 5331 4882
rect 5407 4886 5411 4887
rect 5407 4881 5411 4882
rect 5663 4886 5667 4887
rect 5663 4881 5667 4882
rect 5408 4857 5410 4881
rect 5664 4858 5666 4881
rect 5662 4857 5668 4858
rect 5406 4856 5412 4857
rect 5406 4852 5407 4856
rect 5411 4852 5412 4856
rect 5662 4853 5663 4857
rect 5667 4853 5668 4857
rect 5662 4852 5668 4853
rect 5406 4851 5412 4852
rect 5378 4841 5384 4842
rect 5378 4837 5379 4841
rect 5383 4837 5384 4841
rect 5378 4836 5384 4837
rect 5662 4840 5668 4841
rect 5662 4836 5663 4840
rect 5667 4836 5668 4840
rect 5190 4791 5196 4792
rect 5190 4787 5191 4791
rect 5195 4787 5196 4791
rect 5190 4786 5196 4787
rect 5380 4771 5382 4836
rect 5662 4835 5668 4836
rect 5466 4831 5472 4832
rect 5466 4827 5467 4831
rect 5471 4827 5472 4831
rect 5466 4826 5472 4827
rect 5155 4770 5159 4771
rect 5155 4765 5159 4766
rect 5371 4770 5375 4771
rect 5371 4765 5375 4766
rect 5379 4770 5383 4771
rect 5379 4765 5383 4766
rect 5074 4711 5080 4712
rect 5074 4707 5075 4711
rect 5079 4707 5080 4711
rect 5074 4706 5080 4707
rect 5082 4711 5088 4712
rect 5082 4707 5083 4711
rect 5087 4707 5088 4711
rect 5082 4706 5088 4707
rect 5372 4704 5374 4765
rect 5468 4756 5470 4826
rect 5664 4771 5666 4835
rect 5663 4770 5667 4771
rect 5663 4765 5667 4766
rect 5466 4755 5472 4756
rect 5466 4751 5467 4755
rect 5471 4751 5472 4755
rect 5466 4750 5472 4751
rect 5494 4711 5500 4712
rect 5494 4707 5495 4711
rect 5499 4707 5500 4711
rect 5494 4706 5500 4707
rect 5066 4703 5072 4704
rect 5066 4699 5067 4703
rect 5071 4699 5072 4703
rect 5066 4698 5072 4699
rect 5370 4703 5376 4704
rect 5370 4699 5371 4703
rect 5375 4699 5376 4703
rect 5370 4698 5376 4699
rect 5094 4688 5100 4689
rect 5094 4684 5095 4688
rect 5099 4684 5100 4688
rect 5094 4683 5100 4684
rect 5398 4688 5404 4689
rect 5398 4684 5399 4688
rect 5403 4684 5404 4688
rect 5398 4683 5404 4684
rect 5096 4659 5098 4683
rect 5400 4659 5402 4683
rect 4871 4658 4875 4659
rect 4871 4653 4875 4654
rect 5095 4658 5099 4659
rect 5095 4653 5099 4654
rect 5151 4658 5155 4659
rect 5151 4653 5155 4654
rect 5399 4658 5403 4659
rect 5399 4653 5403 4654
rect 5439 4658 5443 4659
rect 5439 4653 5443 4654
rect 4872 4629 4874 4653
rect 5152 4629 5154 4653
rect 5440 4629 5442 4653
rect 4870 4628 4876 4629
rect 4870 4624 4871 4628
rect 4875 4624 4876 4628
rect 4870 4623 4876 4624
rect 5150 4628 5156 4629
rect 5150 4624 5151 4628
rect 5155 4624 5156 4628
rect 5150 4623 5156 4624
rect 5438 4628 5444 4629
rect 5438 4624 5439 4628
rect 5443 4624 5444 4628
rect 5438 4623 5444 4624
rect 5122 4613 5128 4614
rect 5122 4609 5123 4613
rect 5127 4609 5128 4613
rect 5122 4608 5128 4609
rect 5410 4613 5416 4614
rect 5410 4609 5411 4613
rect 5415 4609 5416 4613
rect 5410 4608 5416 4609
rect 4858 4603 4864 4604
rect 4858 4599 4859 4603
rect 4863 4599 4864 4603
rect 4858 4598 4864 4599
rect 5066 4603 5072 4604
rect 5066 4599 5067 4603
rect 5071 4599 5072 4603
rect 5066 4598 5072 4599
rect 5068 4564 5070 4598
rect 5066 4563 5072 4564
rect 5066 4559 5067 4563
rect 5071 4559 5072 4563
rect 5066 4558 5072 4559
rect 5124 4547 5126 4608
rect 5218 4563 5224 4564
rect 5218 4559 5219 4563
rect 5223 4559 5224 4563
rect 5218 4558 5224 4559
rect 4179 4546 4183 4547
rect 4179 4541 4183 4542
rect 4299 4546 4303 4547
rect 4299 4541 4303 4542
rect 4411 4546 4415 4547
rect 4411 4541 4415 4542
rect 4571 4546 4575 4547
rect 4571 4541 4575 4542
rect 4659 4546 4663 4547
rect 4659 4541 4663 4542
rect 4843 4546 4847 4547
rect 4843 4541 4847 4542
rect 4915 4546 4919 4547
rect 4915 4541 4919 4542
rect 5123 4546 5127 4547
rect 5123 4541 5127 4542
rect 5179 4546 5183 4547
rect 5179 4541 5183 4542
rect 4170 4531 4176 4532
rect 4170 4527 4171 4531
rect 4175 4527 4176 4531
rect 4170 4526 4176 4527
rect 3838 4480 3844 4481
rect 4180 4480 4182 4541
rect 4412 4480 4414 4541
rect 4418 4527 4424 4528
rect 4418 4523 4419 4527
rect 4423 4523 4424 4527
rect 4418 4522 4424 4523
rect 4420 4488 4422 4522
rect 4418 4487 4424 4488
rect 4418 4483 4419 4487
rect 4423 4483 4424 4487
rect 4418 4482 4424 4483
rect 4660 4480 4662 4541
rect 4666 4527 4672 4528
rect 4666 4523 4667 4527
rect 4671 4523 4672 4527
rect 4666 4522 4672 4523
rect 4668 4488 4670 4522
rect 4666 4487 4672 4488
rect 4666 4483 4667 4487
rect 4671 4483 4672 4487
rect 4666 4482 4672 4483
rect 4754 4487 4760 4488
rect 4754 4483 4755 4487
rect 4759 4483 4760 4487
rect 4754 4482 4760 4483
rect 3838 4476 3839 4480
rect 3843 4476 3844 4480
rect 3838 4475 3844 4476
rect 4178 4479 4184 4480
rect 4178 4475 4179 4479
rect 4183 4475 4184 4479
rect 4178 4474 4184 4475
rect 4410 4479 4416 4480
rect 4410 4475 4411 4479
rect 4415 4475 4416 4479
rect 4410 4474 4416 4475
rect 4658 4479 4664 4480
rect 4658 4475 4659 4479
rect 4663 4475 4664 4479
rect 4658 4474 4664 4475
rect 4206 4464 4212 4465
rect 3838 4463 3844 4464
rect 3838 4459 3839 4463
rect 3843 4459 3844 4463
rect 4206 4460 4207 4464
rect 4211 4460 4212 4464
rect 4206 4459 4212 4460
rect 4438 4464 4444 4465
rect 4438 4460 4439 4464
rect 4443 4460 4444 4464
rect 4438 4459 4444 4460
rect 4686 4464 4692 4465
rect 4686 4460 4687 4464
rect 4691 4460 4692 4464
rect 4686 4459 4692 4460
rect 3799 4458 3803 4459
rect 3838 4458 3844 4459
rect 3799 4453 3803 4454
rect 3800 4430 3802 4453
rect 3798 4429 3804 4430
rect 3798 4425 3799 4429
rect 3803 4425 3804 4429
rect 3840 4427 3842 4458
rect 4208 4427 4210 4459
rect 4440 4427 4442 4459
rect 4688 4427 4690 4459
rect 3798 4424 3804 4425
rect 3839 4426 3843 4427
rect 3839 4421 3843 4422
rect 4207 4426 4211 4427
rect 4207 4421 4211 4422
rect 4359 4426 4363 4427
rect 4359 4421 4363 4422
rect 4439 4426 4443 4427
rect 4439 4421 4443 4422
rect 4519 4426 4523 4427
rect 4519 4421 4523 4422
rect 4687 4426 4691 4427
rect 4687 4421 4691 4422
rect 3798 4412 3804 4413
rect 3798 4408 3799 4412
rect 3803 4408 3804 4412
rect 3798 4407 3804 4408
rect 3706 4403 3712 4404
rect 3706 4399 3707 4403
rect 3711 4399 3712 4403
rect 3706 4398 3712 4399
rect 3800 4339 3802 4407
rect 3840 4398 3842 4421
rect 3838 4397 3844 4398
rect 4360 4397 4362 4421
rect 4520 4397 4522 4421
rect 4688 4397 4690 4421
rect 3838 4393 3839 4397
rect 3843 4393 3844 4397
rect 3838 4392 3844 4393
rect 4358 4396 4364 4397
rect 4358 4392 4359 4396
rect 4363 4392 4364 4396
rect 4358 4391 4364 4392
rect 4518 4396 4524 4397
rect 4518 4392 4519 4396
rect 4523 4392 4524 4396
rect 4518 4391 4524 4392
rect 4686 4396 4692 4397
rect 4686 4392 4687 4396
rect 4691 4392 4692 4396
rect 4686 4391 4692 4392
rect 4330 4381 4336 4382
rect 3838 4380 3844 4381
rect 3838 4376 3839 4380
rect 3843 4376 3844 4380
rect 4330 4377 4331 4381
rect 4335 4377 4336 4381
rect 4330 4376 4336 4377
rect 4490 4381 4496 4382
rect 4490 4377 4491 4381
rect 4495 4377 4496 4381
rect 4490 4376 4496 4377
rect 4658 4381 4664 4382
rect 4658 4377 4659 4381
rect 4663 4377 4664 4381
rect 4658 4376 4664 4377
rect 3838 4375 3844 4376
rect 3451 4338 3455 4339
rect 3451 4333 3455 4334
rect 3467 4338 3471 4339
rect 3467 4333 3471 4334
rect 3651 4338 3655 4339
rect 3651 4333 3655 4334
rect 3799 4338 3803 4339
rect 3799 4333 3803 4334
rect 3234 4279 3240 4280
rect 3234 4275 3235 4279
rect 3239 4275 3240 4279
rect 3234 4274 3240 4275
rect 3350 4279 3356 4280
rect 3350 4275 3351 4279
rect 3355 4275 3356 4279
rect 3350 4274 3356 4275
rect 3438 4279 3444 4280
rect 3438 4275 3439 4279
rect 3443 4275 3444 4279
rect 3438 4274 3444 4275
rect 1974 4268 1975 4272
rect 1979 4268 1980 4272
rect 1974 4267 1980 4268
rect 2306 4271 2312 4272
rect 2306 4267 2307 4271
rect 2311 4267 2312 4271
rect 2306 4266 2312 4267
rect 2458 4271 2464 4272
rect 2458 4267 2459 4271
rect 2463 4267 2464 4271
rect 2458 4266 2464 4267
rect 2626 4271 2632 4272
rect 2626 4267 2627 4271
rect 2631 4267 2632 4271
rect 2626 4266 2632 4267
rect 2810 4271 2816 4272
rect 2810 4267 2811 4271
rect 2815 4267 2816 4271
rect 2810 4266 2816 4267
rect 3010 4271 3016 4272
rect 3010 4267 3011 4271
rect 3015 4267 3016 4271
rect 3010 4266 3016 4267
rect 3226 4271 3232 4272
rect 3226 4267 3227 4271
rect 3231 4267 3232 4271
rect 3226 4266 3232 4267
rect 2334 4256 2340 4257
rect 1974 4255 1980 4256
rect 1631 4254 1635 4255
rect 1631 4249 1635 4250
rect 1679 4254 1683 4255
rect 1679 4249 1683 4250
rect 1767 4254 1771 4255
rect 1767 4249 1771 4250
rect 1935 4254 1939 4255
rect 1974 4251 1975 4255
rect 1979 4251 1980 4255
rect 2334 4252 2335 4256
rect 2339 4252 2340 4256
rect 2334 4251 2340 4252
rect 2486 4256 2492 4257
rect 2486 4252 2487 4256
rect 2491 4252 2492 4256
rect 2486 4251 2492 4252
rect 2654 4256 2660 4257
rect 2654 4252 2655 4256
rect 2659 4252 2660 4256
rect 2654 4251 2660 4252
rect 2838 4256 2844 4257
rect 2838 4252 2839 4256
rect 2843 4252 2844 4256
rect 2838 4251 2844 4252
rect 3038 4256 3044 4257
rect 3038 4252 3039 4256
rect 3043 4252 3044 4256
rect 3038 4251 3044 4252
rect 3254 4256 3260 4257
rect 3254 4252 3255 4256
rect 3259 4252 3260 4256
rect 3254 4251 3260 4252
rect 1974 4250 1980 4251
rect 1935 4249 1939 4250
rect 1632 4225 1634 4249
rect 1768 4225 1770 4249
rect 1936 4226 1938 4249
rect 1934 4225 1940 4226
rect 1630 4224 1636 4225
rect 1630 4220 1631 4224
rect 1635 4220 1636 4224
rect 1630 4219 1636 4220
rect 1766 4224 1772 4225
rect 1766 4220 1767 4224
rect 1771 4220 1772 4224
rect 1934 4221 1935 4225
rect 1939 4221 1940 4225
rect 1934 4220 1940 4221
rect 1766 4219 1772 4220
rect 1976 4219 1978 4250
rect 2336 4219 2338 4251
rect 2488 4219 2490 4251
rect 2656 4219 2658 4251
rect 2840 4219 2842 4251
rect 3040 4219 3042 4251
rect 3256 4219 3258 4251
rect 1975 4218 1979 4219
rect 1975 4213 1979 4214
rect 2335 4218 2339 4219
rect 2335 4213 2339 4214
rect 2487 4218 2491 4219
rect 2487 4213 2491 4214
rect 2567 4218 2571 4219
rect 2567 4213 2571 4214
rect 2655 4218 2659 4219
rect 2655 4213 2659 4214
rect 2703 4218 2707 4219
rect 2703 4213 2707 4214
rect 2839 4218 2843 4219
rect 2839 4213 2843 4214
rect 2975 4218 2979 4219
rect 2975 4213 2979 4214
rect 3039 4218 3043 4219
rect 3039 4213 3043 4214
rect 3255 4218 3259 4219
rect 3255 4213 3259 4214
rect 1602 4209 1608 4210
rect 1602 4205 1603 4209
rect 1607 4205 1608 4209
rect 1602 4204 1608 4205
rect 1738 4209 1744 4210
rect 1738 4205 1739 4209
rect 1743 4205 1744 4209
rect 1738 4204 1744 4205
rect 1934 4208 1940 4209
rect 1934 4204 1935 4208
rect 1939 4204 1940 4208
rect 1562 4199 1568 4200
rect 1562 4195 1563 4199
rect 1567 4195 1568 4199
rect 1562 4194 1568 4195
rect 1562 4191 1568 4192
rect 1562 4187 1563 4191
rect 1567 4187 1568 4191
rect 1562 4186 1568 4187
rect 1564 4160 1566 4186
rect 1562 4159 1568 4160
rect 1562 4155 1563 4159
rect 1567 4155 1568 4159
rect 1562 4154 1568 4155
rect 1604 4139 1606 4204
rect 1730 4199 1736 4200
rect 1730 4195 1731 4199
rect 1735 4195 1736 4199
rect 1730 4194 1736 4195
rect 1732 4160 1734 4194
rect 1670 4159 1676 4160
rect 1670 4155 1671 4159
rect 1675 4155 1676 4159
rect 1670 4154 1676 4155
rect 1730 4159 1736 4160
rect 1730 4155 1731 4159
rect 1735 4155 1736 4159
rect 1730 4154 1736 4155
rect 1411 4138 1415 4139
rect 1411 4133 1415 4134
rect 1467 4138 1471 4139
rect 1467 4133 1471 4134
rect 1547 4138 1551 4139
rect 1547 4133 1551 4134
rect 1603 4138 1607 4139
rect 1603 4133 1607 4134
rect 1378 4127 1384 4128
rect 1378 4123 1379 4127
rect 1383 4123 1384 4127
rect 1378 4122 1384 4123
rect 1370 4119 1376 4120
rect 1370 4115 1371 4119
rect 1375 4115 1376 4119
rect 1370 4114 1376 4115
rect 866 4071 872 4072
rect 866 4067 867 4071
rect 871 4067 872 4071
rect 866 4066 872 4067
rect 1002 4071 1008 4072
rect 1002 4067 1003 4071
rect 1007 4067 1008 4071
rect 1002 4066 1008 4067
rect 1138 4071 1144 4072
rect 1138 4067 1139 4071
rect 1143 4067 1144 4071
rect 1138 4066 1144 4067
rect 1274 4071 1280 4072
rect 1274 4067 1275 4071
rect 1279 4067 1280 4071
rect 1274 4066 1280 4067
rect 894 4056 900 4057
rect 894 4052 895 4056
rect 899 4052 900 4056
rect 894 4051 900 4052
rect 1030 4056 1036 4057
rect 1030 4052 1031 4056
rect 1035 4052 1036 4056
rect 1030 4051 1036 4052
rect 1166 4056 1172 4057
rect 1166 4052 1167 4056
rect 1171 4052 1172 4056
rect 1166 4051 1172 4052
rect 1302 4056 1308 4057
rect 1302 4052 1303 4056
rect 1307 4052 1308 4056
rect 1302 4051 1308 4052
rect 896 4003 898 4051
rect 1032 4003 1034 4051
rect 1168 4003 1170 4051
rect 1304 4003 1306 4051
rect 895 4002 899 4003
rect 895 3997 899 3998
rect 983 4002 987 4003
rect 983 3997 987 3998
rect 1031 4002 1035 4003
rect 1031 3997 1035 3998
rect 1151 4002 1155 4003
rect 1151 3997 1155 3998
rect 1167 4002 1171 4003
rect 1167 3997 1171 3998
rect 1303 4002 1307 4003
rect 1303 3997 1307 3998
rect 1319 4002 1323 4003
rect 1319 3997 1323 3998
rect 984 3973 986 3997
rect 1152 3973 1154 3997
rect 1320 3973 1322 3997
rect 982 3972 988 3973
rect 982 3968 983 3972
rect 987 3968 988 3972
rect 982 3967 988 3968
rect 1150 3972 1156 3973
rect 1150 3968 1151 3972
rect 1155 3968 1156 3972
rect 1150 3967 1156 3968
rect 1318 3972 1324 3973
rect 1318 3968 1319 3972
rect 1323 3968 1324 3972
rect 1318 3967 1324 3968
rect 954 3957 960 3958
rect 954 3953 955 3957
rect 959 3953 960 3957
rect 954 3952 960 3953
rect 1122 3957 1128 3958
rect 1122 3953 1123 3957
rect 1127 3953 1128 3957
rect 1122 3952 1128 3953
rect 1290 3957 1296 3958
rect 1290 3953 1291 3957
rect 1295 3953 1296 3957
rect 1290 3952 1296 3953
rect 942 3947 948 3948
rect 942 3943 943 3947
rect 947 3943 948 3947
rect 942 3942 948 3943
rect 944 3908 946 3942
rect 854 3907 860 3908
rect 854 3903 855 3907
rect 859 3903 860 3907
rect 854 3902 860 3903
rect 942 3907 948 3908
rect 942 3903 943 3907
rect 947 3903 948 3907
rect 942 3902 948 3903
rect 956 3863 958 3952
rect 1124 3863 1126 3952
rect 1250 3947 1256 3948
rect 1250 3943 1251 3947
rect 1255 3943 1256 3947
rect 1250 3942 1256 3943
rect 1252 3908 1254 3942
rect 1218 3907 1224 3908
rect 1218 3903 1219 3907
rect 1223 3903 1224 3907
rect 1218 3902 1224 3903
rect 1250 3907 1256 3908
rect 1250 3903 1251 3907
rect 1255 3903 1256 3907
rect 1250 3902 1256 3903
rect 795 3862 799 3863
rect 795 3857 799 3858
rect 939 3862 943 3863
rect 939 3857 943 3858
rect 955 3862 959 3863
rect 955 3857 959 3858
rect 1123 3862 1127 3863
rect 1123 3857 1127 3858
rect 1163 3862 1167 3863
rect 1163 3857 1167 3858
rect 758 3847 764 3848
rect 758 3843 759 3847
rect 763 3843 764 3847
rect 758 3842 764 3843
rect 940 3796 942 3857
rect 1150 3847 1156 3848
rect 1150 3843 1151 3847
rect 1155 3843 1156 3847
rect 1150 3842 1156 3843
rect 514 3795 520 3796
rect 514 3791 515 3795
rect 519 3791 520 3795
rect 514 3790 520 3791
rect 722 3795 728 3796
rect 722 3791 723 3795
rect 727 3791 728 3795
rect 722 3790 728 3791
rect 938 3795 944 3796
rect 938 3791 939 3795
rect 943 3791 944 3795
rect 938 3790 944 3791
rect 542 3780 548 3781
rect 542 3776 543 3780
rect 547 3776 548 3780
rect 542 3775 548 3776
rect 750 3780 756 3781
rect 750 3776 751 3780
rect 755 3776 756 3780
rect 750 3775 756 3776
rect 966 3780 972 3781
rect 966 3776 967 3780
rect 971 3776 972 3780
rect 966 3775 972 3776
rect 544 3751 546 3775
rect 752 3751 754 3775
rect 968 3751 970 3775
rect 527 3750 531 3751
rect 527 3745 531 3746
rect 543 3750 547 3751
rect 543 3745 547 3746
rect 711 3750 715 3751
rect 711 3745 715 3746
rect 751 3750 755 3751
rect 751 3745 755 3746
rect 887 3750 891 3751
rect 887 3745 891 3746
rect 967 3750 971 3751
rect 967 3745 971 3746
rect 1055 3750 1059 3751
rect 1055 3745 1059 3746
rect 528 3721 530 3745
rect 712 3721 714 3745
rect 888 3721 890 3745
rect 1056 3721 1058 3745
rect 526 3720 532 3721
rect 526 3716 527 3720
rect 531 3716 532 3720
rect 526 3715 532 3716
rect 710 3720 716 3721
rect 710 3716 711 3720
rect 715 3716 716 3720
rect 710 3715 716 3716
rect 886 3720 892 3721
rect 886 3716 887 3720
rect 891 3716 892 3720
rect 886 3715 892 3716
rect 1054 3720 1060 3721
rect 1054 3716 1055 3720
rect 1059 3716 1060 3720
rect 1054 3715 1060 3716
rect 498 3705 504 3706
rect 498 3701 499 3705
rect 503 3701 504 3705
rect 498 3700 504 3701
rect 682 3705 688 3706
rect 682 3701 683 3705
rect 687 3701 688 3705
rect 682 3700 688 3701
rect 858 3705 864 3706
rect 858 3701 859 3705
rect 863 3701 864 3705
rect 858 3700 864 3701
rect 1026 3705 1032 3706
rect 1026 3701 1027 3705
rect 1031 3701 1032 3705
rect 1026 3700 1032 3701
rect 434 3695 440 3696
rect 434 3691 435 3695
rect 439 3691 440 3695
rect 434 3690 440 3691
rect 436 3656 438 3690
rect 402 3655 408 3656
rect 402 3651 403 3655
rect 407 3651 408 3655
rect 402 3650 408 3651
rect 434 3655 440 3656
rect 434 3651 435 3655
rect 439 3651 440 3655
rect 434 3650 440 3651
rect 500 3627 502 3700
rect 684 3627 686 3700
rect 810 3695 816 3696
rect 810 3691 811 3695
rect 815 3691 816 3695
rect 810 3690 816 3691
rect 812 3656 814 3690
rect 810 3655 816 3656
rect 810 3651 811 3655
rect 815 3651 816 3655
rect 810 3650 816 3651
rect 860 3627 862 3700
rect 1028 3627 1030 3700
rect 1152 3696 1154 3842
rect 1164 3796 1166 3857
rect 1170 3843 1176 3844
rect 1170 3839 1171 3843
rect 1175 3839 1176 3843
rect 1170 3838 1176 3839
rect 1172 3804 1174 3838
rect 1220 3804 1222 3902
rect 1292 3863 1294 3952
rect 1372 3948 1374 4114
rect 1412 4072 1414 4133
rect 1418 4119 1424 4120
rect 1418 4115 1419 4119
rect 1423 4115 1424 4119
rect 1418 4114 1424 4115
rect 1420 4080 1422 4114
rect 1418 4079 1424 4080
rect 1418 4075 1419 4079
rect 1423 4075 1424 4079
rect 1418 4074 1424 4075
rect 1548 4072 1550 4133
rect 1554 4119 1560 4120
rect 1554 4115 1555 4119
rect 1559 4115 1560 4119
rect 1554 4114 1560 4115
rect 1556 4080 1558 4114
rect 1672 4080 1674 4154
rect 1740 4139 1742 4204
rect 1934 4203 1940 4204
rect 1936 4139 1938 4203
rect 1976 4190 1978 4213
rect 1974 4189 1980 4190
rect 2568 4189 2570 4213
rect 2704 4189 2706 4213
rect 2840 4189 2842 4213
rect 2976 4189 2978 4213
rect 1974 4185 1975 4189
rect 1979 4185 1980 4189
rect 1974 4184 1980 4185
rect 2566 4188 2572 4189
rect 2566 4184 2567 4188
rect 2571 4184 2572 4188
rect 2566 4183 2572 4184
rect 2702 4188 2708 4189
rect 2702 4184 2703 4188
rect 2707 4184 2708 4188
rect 2702 4183 2708 4184
rect 2838 4188 2844 4189
rect 2838 4184 2839 4188
rect 2843 4184 2844 4188
rect 2838 4183 2844 4184
rect 2974 4188 2980 4189
rect 2974 4184 2975 4188
rect 2979 4184 2980 4188
rect 2974 4183 2980 4184
rect 2538 4173 2544 4174
rect 1974 4172 1980 4173
rect 1974 4168 1975 4172
rect 1979 4168 1980 4172
rect 2538 4169 2539 4173
rect 2543 4169 2544 4173
rect 2538 4168 2544 4169
rect 2674 4173 2680 4174
rect 2674 4169 2675 4173
rect 2679 4169 2680 4173
rect 2674 4168 2680 4169
rect 2810 4173 2816 4174
rect 2810 4169 2811 4173
rect 2815 4169 2816 4173
rect 2810 4168 2816 4169
rect 2946 4173 2952 4174
rect 2946 4169 2947 4173
rect 2951 4169 2952 4173
rect 2946 4168 2952 4169
rect 1974 4167 1980 4168
rect 1739 4138 1743 4139
rect 1739 4133 1743 4134
rect 1935 4138 1939 4139
rect 1935 4133 1939 4134
rect 1554 4079 1560 4080
rect 1554 4075 1555 4079
rect 1559 4075 1560 4079
rect 1554 4074 1560 4075
rect 1670 4079 1676 4080
rect 1670 4075 1671 4079
rect 1675 4075 1676 4079
rect 1670 4074 1676 4075
rect 1936 4073 1938 4133
rect 1976 4087 1978 4167
rect 2540 4087 2542 4168
rect 2658 4163 2664 4164
rect 2658 4159 2659 4163
rect 2663 4159 2664 4163
rect 2658 4158 2664 4159
rect 1975 4086 1979 4087
rect 1975 4081 1979 4082
rect 2291 4086 2295 4087
rect 2291 4081 2295 4082
rect 2427 4086 2431 4087
rect 2427 4081 2431 4082
rect 2539 4086 2543 4087
rect 2539 4081 2543 4082
rect 2563 4086 2567 4087
rect 2563 4081 2567 4082
rect 1934 4072 1940 4073
rect 1410 4071 1416 4072
rect 1410 4067 1411 4071
rect 1415 4067 1416 4071
rect 1410 4066 1416 4067
rect 1546 4071 1552 4072
rect 1546 4067 1547 4071
rect 1551 4067 1552 4071
rect 1934 4068 1935 4072
rect 1939 4068 1940 4072
rect 1934 4067 1940 4068
rect 1546 4066 1552 4067
rect 1438 4056 1444 4057
rect 1438 4052 1439 4056
rect 1443 4052 1444 4056
rect 1438 4051 1444 4052
rect 1574 4056 1580 4057
rect 1574 4052 1575 4056
rect 1579 4052 1580 4056
rect 1574 4051 1580 4052
rect 1934 4055 1940 4056
rect 1934 4051 1935 4055
rect 1939 4051 1940 4055
rect 1440 4003 1442 4051
rect 1576 4003 1578 4051
rect 1934 4050 1940 4051
rect 1936 4003 1938 4050
rect 1976 4021 1978 4081
rect 1974 4020 1980 4021
rect 2292 4020 2294 4081
rect 2386 4067 2392 4068
rect 2386 4063 2387 4067
rect 2391 4063 2392 4067
rect 2386 4062 2392 4063
rect 2388 4053 2390 4062
rect 2387 4052 2391 4053
rect 2387 4047 2391 4048
rect 2428 4020 2430 4081
rect 2434 4067 2440 4068
rect 2434 4063 2435 4067
rect 2439 4063 2440 4067
rect 2434 4062 2440 4063
rect 2436 4028 2438 4062
rect 2434 4027 2440 4028
rect 2434 4023 2435 4027
rect 2439 4023 2440 4027
rect 2434 4022 2440 4023
rect 2550 4027 2556 4028
rect 2550 4023 2551 4027
rect 2555 4023 2556 4027
rect 2550 4022 2556 4023
rect 1974 4016 1975 4020
rect 1979 4016 1980 4020
rect 1974 4015 1980 4016
rect 2290 4019 2296 4020
rect 2290 4015 2291 4019
rect 2295 4015 2296 4019
rect 2290 4014 2296 4015
rect 2426 4019 2432 4020
rect 2426 4015 2427 4019
rect 2431 4015 2432 4019
rect 2426 4014 2432 4015
rect 2318 4004 2324 4005
rect 1974 4003 1980 4004
rect 1439 4002 1443 4003
rect 1439 3997 1443 3998
rect 1575 4002 1579 4003
rect 1575 3997 1579 3998
rect 1935 4002 1939 4003
rect 1974 3999 1975 4003
rect 1979 3999 1980 4003
rect 2318 4000 2319 4004
rect 2323 4000 2324 4004
rect 2318 3999 2324 4000
rect 2454 4004 2460 4005
rect 2454 4000 2455 4004
rect 2459 4000 2460 4004
rect 2454 3999 2460 4000
rect 1974 3998 1980 3999
rect 1935 3997 1939 3998
rect 1936 3974 1938 3997
rect 1934 3973 1940 3974
rect 1934 3969 1935 3973
rect 1939 3969 1940 3973
rect 1976 3971 1978 3998
rect 2320 3971 2322 3999
rect 2456 3971 2458 3999
rect 1934 3968 1940 3969
rect 1975 3970 1979 3971
rect 1975 3965 1979 3966
rect 2119 3970 2123 3971
rect 2119 3965 2123 3966
rect 2319 3970 2323 3971
rect 2319 3965 2323 3966
rect 2327 3970 2331 3971
rect 2327 3965 2331 3966
rect 2455 3970 2459 3971
rect 2455 3965 2459 3966
rect 2535 3970 2539 3971
rect 2535 3965 2539 3966
rect 1934 3956 1940 3957
rect 1934 3952 1935 3956
rect 1939 3952 1940 3956
rect 1934 3951 1940 3952
rect 1370 3947 1376 3948
rect 1370 3943 1371 3947
rect 1375 3943 1376 3947
rect 1370 3942 1376 3943
rect 1936 3863 1938 3951
rect 1976 3942 1978 3965
rect 1974 3941 1980 3942
rect 2120 3941 2122 3965
rect 2328 3941 2330 3965
rect 2536 3941 2538 3965
rect 1974 3937 1975 3941
rect 1979 3937 1980 3941
rect 1974 3936 1980 3937
rect 2118 3940 2124 3941
rect 2118 3936 2119 3940
rect 2123 3936 2124 3940
rect 2118 3935 2124 3936
rect 2326 3940 2332 3941
rect 2326 3936 2327 3940
rect 2331 3936 2332 3940
rect 2326 3935 2332 3936
rect 2534 3940 2540 3941
rect 2534 3936 2535 3940
rect 2539 3936 2540 3940
rect 2534 3935 2540 3936
rect 2090 3925 2096 3926
rect 1974 3924 1980 3925
rect 1974 3920 1975 3924
rect 1979 3920 1980 3924
rect 2090 3921 2091 3925
rect 2095 3921 2096 3925
rect 2090 3920 2096 3921
rect 2298 3925 2304 3926
rect 2298 3921 2299 3925
rect 2303 3921 2304 3925
rect 2298 3920 2304 3921
rect 2506 3925 2512 3926
rect 2506 3921 2507 3925
rect 2511 3921 2512 3925
rect 2506 3920 2512 3921
rect 1974 3919 1980 3920
rect 1291 3862 1295 3863
rect 1291 3857 1295 3858
rect 1935 3862 1939 3863
rect 1935 3857 1939 3858
rect 1170 3803 1176 3804
rect 1170 3799 1171 3803
rect 1175 3799 1176 3803
rect 1170 3798 1176 3799
rect 1218 3803 1224 3804
rect 1218 3799 1219 3803
rect 1223 3799 1224 3803
rect 1218 3798 1224 3799
rect 1936 3797 1938 3857
rect 1976 3847 1978 3919
rect 2092 3847 2094 3920
rect 2214 3915 2220 3916
rect 2214 3911 2215 3915
rect 2219 3911 2220 3915
rect 2214 3910 2220 3911
rect 2290 3915 2296 3916
rect 2290 3911 2291 3915
rect 2295 3911 2296 3915
rect 2290 3910 2296 3911
rect 1975 3846 1979 3847
rect 1975 3841 1979 3842
rect 2091 3846 2095 3847
rect 2091 3841 2095 3842
rect 2139 3846 2143 3847
rect 2139 3841 2143 3842
rect 1934 3796 1940 3797
rect 1162 3795 1168 3796
rect 1162 3791 1163 3795
rect 1167 3791 1168 3795
rect 1934 3792 1935 3796
rect 1939 3792 1940 3796
rect 1934 3791 1940 3792
rect 1162 3790 1168 3791
rect 1976 3781 1978 3841
rect 1190 3780 1196 3781
rect 1974 3780 1980 3781
rect 2140 3780 2142 3841
rect 2216 3832 2218 3910
rect 2292 3876 2294 3910
rect 2290 3875 2296 3876
rect 2290 3871 2291 3875
rect 2295 3871 2296 3875
rect 2290 3870 2296 3871
rect 2300 3847 2302 3920
rect 2394 3907 2400 3908
rect 2394 3903 2395 3907
rect 2399 3903 2400 3907
rect 2394 3902 2400 3903
rect 2396 3876 2398 3902
rect 2394 3875 2400 3876
rect 2394 3871 2395 3875
rect 2399 3871 2400 3875
rect 2394 3870 2400 3871
rect 2508 3847 2510 3920
rect 2552 3876 2554 4022
rect 2564 4020 2566 4081
rect 2660 4072 2662 4158
rect 2676 4087 2678 4168
rect 2812 4087 2814 4168
rect 2948 4087 2950 4168
rect 2954 4163 2960 4164
rect 2954 4159 2955 4163
rect 2959 4159 2960 4163
rect 2954 4158 2960 4159
rect 2956 4132 2958 4158
rect 2954 4131 2960 4132
rect 2954 4127 2955 4131
rect 2959 4127 2960 4131
rect 2954 4126 2960 4127
rect 3352 4124 3354 4274
rect 3452 4272 3454 4333
rect 3642 4323 3648 4324
rect 3642 4319 3643 4323
rect 3647 4319 3648 4323
rect 3642 4318 3648 4319
rect 3644 4280 3646 4318
rect 3642 4279 3648 4280
rect 3642 4275 3643 4279
rect 3647 4275 3648 4279
rect 3642 4274 3648 4275
rect 3652 4272 3654 4333
rect 3800 4273 3802 4333
rect 3840 4315 3842 4375
rect 3982 4323 3988 4324
rect 3982 4319 3983 4323
rect 3987 4319 3988 4323
rect 3982 4318 3988 4319
rect 3839 4314 3843 4315
rect 3839 4309 3843 4310
rect 3859 4314 3863 4315
rect 3859 4309 3863 4310
rect 3798 4272 3804 4273
rect 3450 4271 3456 4272
rect 3450 4267 3451 4271
rect 3455 4267 3456 4271
rect 3450 4266 3456 4267
rect 3650 4271 3656 4272
rect 3650 4267 3651 4271
rect 3655 4267 3656 4271
rect 3798 4268 3799 4272
rect 3803 4268 3804 4272
rect 3798 4267 3804 4268
rect 3650 4266 3656 4267
rect 3478 4256 3484 4257
rect 3478 4252 3479 4256
rect 3483 4252 3484 4256
rect 3478 4251 3484 4252
rect 3678 4256 3684 4257
rect 3678 4252 3679 4256
rect 3683 4252 3684 4256
rect 3678 4251 3684 4252
rect 3798 4255 3804 4256
rect 3798 4251 3799 4255
rect 3803 4251 3804 4255
rect 3480 4219 3482 4251
rect 3680 4219 3682 4251
rect 3798 4250 3804 4251
rect 3800 4219 3802 4250
rect 3840 4249 3842 4309
rect 3838 4248 3844 4249
rect 3860 4248 3862 4309
rect 3984 4256 3986 4318
rect 4332 4315 4334 4376
rect 4346 4371 4352 4372
rect 4346 4367 4347 4371
rect 4351 4367 4352 4371
rect 4346 4366 4352 4367
rect 4482 4371 4488 4372
rect 4482 4367 4483 4371
rect 4487 4367 4488 4371
rect 4482 4366 4488 4367
rect 4043 4314 4047 4315
rect 4043 4309 4047 4310
rect 4251 4314 4255 4315
rect 4251 4309 4255 4310
rect 4331 4314 4335 4315
rect 4331 4309 4335 4310
rect 3982 4255 3988 4256
rect 3982 4251 3983 4255
rect 3987 4251 3988 4255
rect 3982 4250 3988 4251
rect 4044 4248 4046 4309
rect 4050 4295 4056 4296
rect 4050 4291 4051 4295
rect 4055 4291 4056 4295
rect 4050 4290 4056 4291
rect 3838 4244 3839 4248
rect 3843 4244 3844 4248
rect 3838 4243 3844 4244
rect 3858 4247 3864 4248
rect 3858 4243 3859 4247
rect 3863 4243 3864 4247
rect 3858 4242 3864 4243
rect 4042 4247 4048 4248
rect 4042 4243 4043 4247
rect 4047 4243 4048 4247
rect 4042 4242 4048 4243
rect 3886 4232 3892 4233
rect 3838 4231 3844 4232
rect 3838 4227 3839 4231
rect 3843 4227 3844 4231
rect 3886 4228 3887 4232
rect 3891 4228 3892 4232
rect 3886 4227 3892 4228
rect 3838 4226 3844 4227
rect 3479 4218 3483 4219
rect 3479 4213 3483 4214
rect 3679 4218 3683 4219
rect 3679 4213 3683 4214
rect 3799 4218 3803 4219
rect 3799 4213 3803 4214
rect 3800 4190 3802 4213
rect 3798 4189 3804 4190
rect 3798 4185 3799 4189
rect 3803 4185 3804 4189
rect 3798 4184 3804 4185
rect 3798 4172 3804 4173
rect 3798 4168 3799 4172
rect 3803 4168 3804 4172
rect 3798 4167 3804 4168
rect 3840 4167 3842 4226
rect 3888 4167 3890 4227
rect 3350 4123 3356 4124
rect 3350 4119 3351 4123
rect 3355 4119 3356 4123
rect 3350 4118 3356 4119
rect 3800 4087 3802 4167
rect 3839 4166 3843 4167
rect 3839 4161 3843 4162
rect 3887 4166 3891 4167
rect 3887 4161 3891 4162
rect 3840 4138 3842 4161
rect 3838 4137 3844 4138
rect 3888 4137 3890 4161
rect 3838 4133 3839 4137
rect 3843 4133 3844 4137
rect 3838 4132 3844 4133
rect 3886 4136 3892 4137
rect 3886 4132 3887 4136
rect 3891 4132 3892 4136
rect 3886 4131 3892 4132
rect 3858 4121 3864 4122
rect 3838 4120 3844 4121
rect 3838 4116 3839 4120
rect 3843 4116 3844 4120
rect 3858 4117 3859 4121
rect 3863 4117 3864 4121
rect 3858 4116 3864 4117
rect 3838 4115 3844 4116
rect 2675 4086 2679 4087
rect 2675 4081 2679 4082
rect 2699 4086 2703 4087
rect 2699 4081 2703 4082
rect 2811 4086 2815 4087
rect 2811 4081 2815 4082
rect 2835 4086 2839 4087
rect 2835 4081 2839 4082
rect 2947 4086 2951 4087
rect 2947 4081 2951 4082
rect 3799 4086 3803 4087
rect 3799 4081 3803 4082
rect 2658 4071 2664 4072
rect 2658 4067 2659 4071
rect 2663 4067 2664 4071
rect 2658 4066 2664 4067
rect 2700 4020 2702 4081
rect 2706 4067 2712 4068
rect 2706 4063 2707 4067
rect 2711 4063 2712 4067
rect 2706 4062 2712 4063
rect 2708 4028 2710 4062
rect 2706 4027 2712 4028
rect 2706 4023 2707 4027
rect 2711 4023 2712 4027
rect 2706 4022 2712 4023
rect 2836 4020 2838 4081
rect 2842 4067 2848 4068
rect 2842 4063 2843 4067
rect 2847 4063 2848 4067
rect 2842 4062 2848 4063
rect 2844 4028 2846 4062
rect 2959 4052 2963 4053
rect 2959 4047 2963 4048
rect 2960 4028 2962 4047
rect 2842 4027 2848 4028
rect 2842 4023 2843 4027
rect 2847 4023 2848 4027
rect 2842 4022 2848 4023
rect 2958 4027 2964 4028
rect 2958 4023 2959 4027
rect 2963 4023 2964 4027
rect 2958 4022 2964 4023
rect 3800 4021 3802 4081
rect 3840 4055 3842 4115
rect 3860 4055 3862 4116
rect 4052 4112 4054 4290
rect 4252 4248 4254 4309
rect 4348 4300 4350 4366
rect 4484 4332 4486 4366
rect 4482 4331 4488 4332
rect 4482 4327 4483 4331
rect 4487 4327 4488 4331
rect 4482 4326 4488 4327
rect 4492 4315 4494 4376
rect 4660 4315 4662 4376
rect 4756 4332 4758 4482
rect 4916 4480 4918 4541
rect 4974 4531 4980 4532
rect 4974 4527 4975 4531
rect 4979 4527 4980 4531
rect 4974 4526 4980 4527
rect 4914 4479 4920 4480
rect 4914 4475 4915 4479
rect 4919 4475 4920 4479
rect 4914 4474 4920 4475
rect 4942 4464 4948 4465
rect 4942 4460 4943 4464
rect 4947 4460 4948 4464
rect 4942 4459 4948 4460
rect 4944 4427 4946 4459
rect 4879 4426 4883 4427
rect 4879 4421 4883 4422
rect 4943 4426 4947 4427
rect 4943 4421 4947 4422
rect 4880 4397 4882 4421
rect 4878 4396 4884 4397
rect 4878 4392 4879 4396
rect 4883 4392 4884 4396
rect 4878 4391 4884 4392
rect 4850 4381 4856 4382
rect 4850 4377 4851 4381
rect 4855 4377 4856 4381
rect 4850 4376 4856 4377
rect 4754 4331 4760 4332
rect 4754 4327 4755 4331
rect 4759 4327 4760 4331
rect 4754 4326 4760 4327
rect 4852 4315 4854 4376
rect 4976 4372 4978 4526
rect 5180 4480 5182 4541
rect 5186 4527 5192 4528
rect 5186 4523 5187 4527
rect 5191 4523 5192 4527
rect 5186 4522 5192 4523
rect 5188 4488 5190 4522
rect 5220 4488 5222 4558
rect 5412 4547 5414 4608
rect 5496 4564 5498 4706
rect 5664 4705 5666 4765
rect 5662 4704 5668 4705
rect 5662 4700 5663 4704
rect 5667 4700 5668 4704
rect 5662 4699 5668 4700
rect 5662 4687 5668 4688
rect 5662 4683 5663 4687
rect 5667 4683 5668 4687
rect 5662 4682 5668 4683
rect 5664 4659 5666 4682
rect 5663 4658 5667 4659
rect 5663 4653 5667 4654
rect 5664 4630 5666 4653
rect 5662 4629 5668 4630
rect 5662 4625 5663 4629
rect 5667 4625 5668 4629
rect 5662 4624 5668 4625
rect 5662 4612 5668 4613
rect 5662 4608 5663 4612
rect 5667 4608 5668 4612
rect 5662 4607 5668 4608
rect 5534 4603 5540 4604
rect 5534 4599 5535 4603
rect 5539 4599 5540 4603
rect 5534 4598 5540 4599
rect 5494 4563 5500 4564
rect 5494 4559 5495 4563
rect 5499 4559 5500 4563
rect 5494 4558 5500 4559
rect 5411 4546 5415 4547
rect 5411 4541 5415 4542
rect 5443 4546 5447 4547
rect 5443 4541 5447 4542
rect 5186 4487 5192 4488
rect 5186 4483 5187 4487
rect 5191 4483 5192 4487
rect 5186 4482 5192 4483
rect 5218 4487 5224 4488
rect 5218 4483 5219 4487
rect 5223 4483 5224 4487
rect 5218 4482 5224 4483
rect 5444 4480 5446 4541
rect 5536 4532 5538 4598
rect 5664 4547 5666 4607
rect 5663 4546 5667 4547
rect 5663 4541 5667 4542
rect 5534 4531 5540 4532
rect 5534 4527 5535 4531
rect 5539 4527 5540 4531
rect 5534 4526 5540 4527
rect 5566 4487 5572 4488
rect 5566 4483 5567 4487
rect 5571 4483 5572 4487
rect 5566 4482 5572 4483
rect 5178 4479 5184 4480
rect 5178 4475 5179 4479
rect 5183 4475 5184 4479
rect 5178 4474 5184 4475
rect 5442 4479 5448 4480
rect 5442 4475 5443 4479
rect 5447 4475 5448 4479
rect 5442 4474 5448 4475
rect 5206 4464 5212 4465
rect 5206 4460 5207 4464
rect 5211 4460 5212 4464
rect 5206 4459 5212 4460
rect 5470 4464 5476 4465
rect 5470 4460 5471 4464
rect 5475 4460 5476 4464
rect 5470 4459 5476 4460
rect 5208 4427 5210 4459
rect 5472 4427 5474 4459
rect 5079 4426 5083 4427
rect 5079 4421 5083 4422
rect 5207 4426 5211 4427
rect 5207 4421 5211 4422
rect 5287 4426 5291 4427
rect 5287 4421 5291 4422
rect 5471 4426 5475 4427
rect 5471 4421 5475 4422
rect 5503 4426 5507 4427
rect 5503 4421 5507 4422
rect 5080 4397 5082 4421
rect 5288 4397 5290 4421
rect 5504 4397 5506 4421
rect 5078 4396 5084 4397
rect 5078 4392 5079 4396
rect 5083 4392 5084 4396
rect 5078 4391 5084 4392
rect 5286 4396 5292 4397
rect 5286 4392 5287 4396
rect 5291 4392 5292 4396
rect 5286 4391 5292 4392
rect 5502 4396 5508 4397
rect 5502 4392 5503 4396
rect 5507 4392 5508 4396
rect 5502 4391 5508 4392
rect 5050 4381 5056 4382
rect 5050 4377 5051 4381
rect 5055 4377 5056 4381
rect 5050 4376 5056 4377
rect 5258 4381 5264 4382
rect 5258 4377 5259 4381
rect 5263 4377 5264 4381
rect 5258 4376 5264 4377
rect 5474 4381 5480 4382
rect 5474 4377 5475 4381
rect 5479 4377 5480 4381
rect 5474 4376 5480 4377
rect 4974 4371 4980 4372
rect 4974 4367 4975 4371
rect 4979 4367 4980 4371
rect 4974 4366 4980 4367
rect 5010 4371 5016 4372
rect 5010 4367 5011 4371
rect 5015 4367 5016 4371
rect 5010 4366 5016 4367
rect 5012 4332 5014 4366
rect 5010 4331 5016 4332
rect 5010 4327 5011 4331
rect 5015 4327 5016 4331
rect 5010 4326 5016 4327
rect 5052 4315 5054 4376
rect 5260 4315 5262 4376
rect 5354 4331 5360 4332
rect 5354 4327 5355 4331
rect 5359 4327 5360 4331
rect 5354 4326 5360 4327
rect 4475 4314 4479 4315
rect 4475 4309 4479 4310
rect 4491 4314 4495 4315
rect 4491 4309 4495 4310
rect 4659 4314 4663 4315
rect 4659 4309 4663 4310
rect 4715 4314 4719 4315
rect 4715 4309 4719 4310
rect 4851 4314 4855 4315
rect 4851 4309 4855 4310
rect 4971 4314 4975 4315
rect 4971 4309 4975 4310
rect 5051 4314 5055 4315
rect 5051 4309 5055 4310
rect 5235 4314 5239 4315
rect 5235 4309 5239 4310
rect 5259 4314 5263 4315
rect 5259 4309 5263 4310
rect 4346 4299 4352 4300
rect 4346 4295 4347 4299
rect 4351 4295 4352 4299
rect 4346 4294 4352 4295
rect 4476 4248 4478 4309
rect 4482 4295 4488 4296
rect 4482 4291 4483 4295
rect 4487 4291 4488 4295
rect 4482 4290 4488 4291
rect 4484 4256 4486 4290
rect 4482 4255 4488 4256
rect 4482 4251 4483 4255
rect 4487 4251 4488 4255
rect 4482 4250 4488 4251
rect 4716 4248 4718 4309
rect 4722 4295 4728 4296
rect 4722 4291 4723 4295
rect 4727 4291 4728 4295
rect 4722 4290 4728 4291
rect 4724 4256 4726 4290
rect 4722 4255 4728 4256
rect 4722 4251 4723 4255
rect 4727 4251 4728 4255
rect 4722 4250 4728 4251
rect 4972 4248 4974 4309
rect 4978 4295 4984 4296
rect 4978 4291 4979 4295
rect 4983 4291 4984 4295
rect 4978 4290 4984 4291
rect 4980 4256 4982 4290
rect 4978 4255 4984 4256
rect 4978 4251 4979 4255
rect 4983 4251 4984 4255
rect 4978 4250 4984 4251
rect 5236 4248 5238 4309
rect 5242 4295 5248 4296
rect 5242 4291 5243 4295
rect 5247 4291 5248 4295
rect 5242 4290 5248 4291
rect 5244 4256 5246 4290
rect 5356 4256 5358 4326
rect 5476 4315 5478 4376
rect 5568 4332 5570 4482
rect 5664 4481 5666 4541
rect 5662 4480 5668 4481
rect 5662 4476 5663 4480
rect 5667 4476 5668 4480
rect 5662 4475 5668 4476
rect 5662 4463 5668 4464
rect 5662 4459 5663 4463
rect 5667 4459 5668 4463
rect 5662 4458 5668 4459
rect 5664 4427 5666 4458
rect 5663 4426 5667 4427
rect 5663 4421 5667 4422
rect 5664 4398 5666 4421
rect 5662 4397 5668 4398
rect 5662 4393 5663 4397
rect 5667 4393 5668 4397
rect 5662 4392 5668 4393
rect 5662 4380 5668 4381
rect 5662 4376 5663 4380
rect 5667 4376 5668 4380
rect 5662 4375 5668 4376
rect 5594 4371 5600 4372
rect 5594 4367 5595 4371
rect 5599 4367 5600 4371
rect 5594 4366 5600 4367
rect 5566 4331 5572 4332
rect 5566 4327 5567 4331
rect 5571 4327 5572 4331
rect 5566 4326 5572 4327
rect 5475 4314 5479 4315
rect 5475 4309 5479 4310
rect 5499 4314 5503 4315
rect 5499 4309 5503 4310
rect 5242 4255 5248 4256
rect 5242 4251 5243 4255
rect 5247 4251 5248 4255
rect 5242 4250 5248 4251
rect 5354 4255 5360 4256
rect 5354 4251 5355 4255
rect 5359 4251 5360 4255
rect 5354 4250 5360 4251
rect 5500 4248 5502 4309
rect 5596 4300 5598 4366
rect 5664 4315 5666 4375
rect 5663 4314 5667 4315
rect 5663 4309 5667 4310
rect 5594 4299 5600 4300
rect 5594 4295 5595 4299
rect 5599 4295 5600 4299
rect 5594 4294 5600 4295
rect 5610 4255 5616 4256
rect 5610 4251 5611 4255
rect 5615 4251 5616 4255
rect 5610 4250 5616 4251
rect 4250 4247 4256 4248
rect 4250 4243 4251 4247
rect 4255 4243 4256 4247
rect 4250 4242 4256 4243
rect 4474 4247 4480 4248
rect 4474 4243 4475 4247
rect 4479 4243 4480 4247
rect 4474 4242 4480 4243
rect 4714 4247 4720 4248
rect 4714 4243 4715 4247
rect 4719 4243 4720 4247
rect 4714 4242 4720 4243
rect 4970 4247 4976 4248
rect 4970 4243 4971 4247
rect 4975 4243 4976 4247
rect 4970 4242 4976 4243
rect 5234 4247 5240 4248
rect 5234 4243 5235 4247
rect 5239 4243 5240 4247
rect 5234 4242 5240 4243
rect 5498 4247 5504 4248
rect 5498 4243 5499 4247
rect 5503 4243 5504 4247
rect 5498 4242 5504 4243
rect 4070 4232 4076 4233
rect 4070 4228 4071 4232
rect 4075 4228 4076 4232
rect 4070 4227 4076 4228
rect 4278 4232 4284 4233
rect 4278 4228 4279 4232
rect 4283 4228 4284 4232
rect 4278 4227 4284 4228
rect 4502 4232 4508 4233
rect 4502 4228 4503 4232
rect 4507 4228 4508 4232
rect 4502 4227 4508 4228
rect 4742 4232 4748 4233
rect 4742 4228 4743 4232
rect 4747 4228 4748 4232
rect 4742 4227 4748 4228
rect 4998 4232 5004 4233
rect 4998 4228 4999 4232
rect 5003 4228 5004 4232
rect 4998 4227 5004 4228
rect 5262 4232 5268 4233
rect 5262 4228 5263 4232
rect 5267 4228 5268 4232
rect 5262 4227 5268 4228
rect 5526 4232 5532 4233
rect 5526 4228 5527 4232
rect 5531 4228 5532 4232
rect 5526 4227 5532 4228
rect 4072 4167 4074 4227
rect 4280 4167 4282 4227
rect 4504 4167 4506 4227
rect 4744 4167 4746 4227
rect 5000 4167 5002 4227
rect 5264 4167 5266 4227
rect 5528 4167 5530 4227
rect 4071 4166 4075 4167
rect 4071 4161 4075 4162
rect 4279 4166 4283 4167
rect 4279 4161 4283 4162
rect 4415 4166 4419 4167
rect 4415 4161 4419 4162
rect 4503 4166 4507 4167
rect 4503 4161 4507 4162
rect 4743 4166 4747 4167
rect 4743 4161 4747 4162
rect 4975 4166 4979 4167
rect 4975 4161 4979 4162
rect 4999 4166 5003 4167
rect 4999 4161 5003 4162
rect 5263 4166 5267 4167
rect 5263 4161 5267 4162
rect 5527 4166 5531 4167
rect 5527 4161 5531 4162
rect 5543 4166 5547 4167
rect 5543 4161 5547 4162
rect 4416 4137 4418 4161
rect 4976 4137 4978 4161
rect 5544 4137 5546 4161
rect 4414 4136 4420 4137
rect 4414 4132 4415 4136
rect 4419 4132 4420 4136
rect 4414 4131 4420 4132
rect 4974 4136 4980 4137
rect 4974 4132 4975 4136
rect 4979 4132 4980 4136
rect 4974 4131 4980 4132
rect 5542 4136 5548 4137
rect 5542 4132 5543 4136
rect 5547 4132 5548 4136
rect 5542 4131 5548 4132
rect 4386 4121 4392 4122
rect 4386 4117 4387 4121
rect 4391 4117 4392 4121
rect 4386 4116 4392 4117
rect 4946 4121 4952 4122
rect 4946 4117 4947 4121
rect 4951 4117 4952 4121
rect 4946 4116 4952 4117
rect 5514 4121 5520 4122
rect 5514 4117 5515 4121
rect 5519 4117 5520 4121
rect 5514 4116 5520 4117
rect 4050 4111 4056 4112
rect 4050 4107 4051 4111
rect 4055 4107 4056 4111
rect 4050 4106 4056 4107
rect 3954 4103 3960 4104
rect 3954 4099 3955 4103
rect 3959 4099 3960 4103
rect 3954 4098 3960 4099
rect 3956 4072 3958 4098
rect 3954 4071 3960 4072
rect 3954 4067 3955 4071
rect 3959 4067 3960 4071
rect 3954 4066 3960 4067
rect 4388 4055 4390 4116
rect 4878 4111 4884 4112
rect 4878 4107 4879 4111
rect 4883 4107 4884 4111
rect 4878 4106 4884 4107
rect 4880 4072 4882 4106
rect 4878 4071 4884 4072
rect 4878 4067 4879 4071
rect 4883 4067 4884 4071
rect 4878 4066 4884 4067
rect 4948 4055 4950 4116
rect 5516 4055 5518 4116
rect 5612 4072 5614 4250
rect 5664 4249 5666 4309
rect 5662 4248 5668 4249
rect 5662 4244 5663 4248
rect 5667 4244 5668 4248
rect 5662 4243 5668 4244
rect 5662 4231 5668 4232
rect 5662 4227 5663 4231
rect 5667 4227 5668 4231
rect 5662 4226 5668 4227
rect 5664 4167 5666 4226
rect 5663 4166 5667 4167
rect 5663 4161 5667 4162
rect 5664 4138 5666 4161
rect 5662 4137 5668 4138
rect 5662 4133 5663 4137
rect 5667 4133 5668 4137
rect 5662 4132 5668 4133
rect 5662 4120 5668 4121
rect 5662 4116 5663 4120
rect 5667 4116 5668 4120
rect 5662 4115 5668 4116
rect 5618 4111 5624 4112
rect 5618 4107 5619 4111
rect 5623 4107 5624 4111
rect 5618 4106 5624 4107
rect 5610 4071 5616 4072
rect 5610 4067 5611 4071
rect 5615 4067 5616 4071
rect 5610 4066 5616 4067
rect 3839 4054 3843 4055
rect 3839 4049 3843 4050
rect 3859 4054 3863 4055
rect 3859 4049 3863 4050
rect 4003 4054 4007 4055
rect 4003 4049 4007 4050
rect 4171 4054 4175 4055
rect 4171 4049 4175 4050
rect 4339 4054 4343 4055
rect 4339 4049 4343 4050
rect 4387 4054 4391 4055
rect 4387 4049 4391 4050
rect 4499 4054 4503 4055
rect 4499 4049 4503 4050
rect 4651 4054 4655 4055
rect 4651 4049 4655 4050
rect 4803 4054 4807 4055
rect 4803 4049 4807 4050
rect 4947 4054 4951 4055
rect 4947 4049 4951 4050
rect 5091 4054 5095 4055
rect 5091 4049 5095 4050
rect 5235 4054 5239 4055
rect 5235 4049 5239 4050
rect 5379 4054 5383 4055
rect 5379 4049 5383 4050
rect 5515 4054 5519 4055
rect 5515 4049 5519 4050
rect 3798 4020 3804 4021
rect 2562 4019 2568 4020
rect 2562 4015 2563 4019
rect 2567 4015 2568 4019
rect 2562 4014 2568 4015
rect 2698 4019 2704 4020
rect 2698 4015 2699 4019
rect 2703 4015 2704 4019
rect 2698 4014 2704 4015
rect 2834 4019 2840 4020
rect 2834 4015 2835 4019
rect 2839 4015 2840 4019
rect 3798 4016 3799 4020
rect 3803 4016 3804 4020
rect 3798 4015 3804 4016
rect 2834 4014 2840 4015
rect 2590 4004 2596 4005
rect 2590 4000 2591 4004
rect 2595 4000 2596 4004
rect 2590 3999 2596 4000
rect 2726 4004 2732 4005
rect 2726 4000 2727 4004
rect 2731 4000 2732 4004
rect 2726 3999 2732 4000
rect 2862 4004 2868 4005
rect 2862 4000 2863 4004
rect 2867 4000 2868 4004
rect 2862 3999 2868 4000
rect 3798 4003 3804 4004
rect 3798 3999 3799 4003
rect 3803 3999 3804 4003
rect 2592 3971 2594 3999
rect 2728 3971 2730 3999
rect 2864 3971 2866 3999
rect 3798 3998 3804 3999
rect 3800 3971 3802 3998
rect 3840 3989 3842 4049
rect 3838 3988 3844 3989
rect 3860 3988 3862 4049
rect 3866 4035 3872 4036
rect 3866 4031 3867 4035
rect 3871 4031 3872 4035
rect 3866 4030 3872 4031
rect 3838 3984 3839 3988
rect 3843 3984 3844 3988
rect 3838 3983 3844 3984
rect 3858 3987 3864 3988
rect 3858 3983 3859 3987
rect 3863 3983 3864 3987
rect 3858 3982 3864 3983
rect 3838 3971 3844 3972
rect 2591 3970 2595 3971
rect 2591 3965 2595 3966
rect 2727 3970 2731 3971
rect 2727 3965 2731 3966
rect 2743 3970 2747 3971
rect 2743 3965 2747 3966
rect 2863 3970 2867 3971
rect 2863 3965 2867 3966
rect 2943 3970 2947 3971
rect 2943 3965 2947 3966
rect 3135 3970 3139 3971
rect 3135 3965 3139 3966
rect 3319 3970 3323 3971
rect 3319 3965 3323 3966
rect 3511 3970 3515 3971
rect 3511 3965 3515 3966
rect 3679 3970 3683 3971
rect 3679 3965 3683 3966
rect 3799 3970 3803 3971
rect 3838 3967 3839 3971
rect 3843 3967 3844 3971
rect 3838 3966 3844 3967
rect 3799 3965 3803 3966
rect 2744 3941 2746 3965
rect 2944 3941 2946 3965
rect 3136 3941 3138 3965
rect 3320 3941 3322 3965
rect 3512 3941 3514 3965
rect 3680 3941 3682 3965
rect 3800 3942 3802 3965
rect 3798 3941 3804 3942
rect 2742 3940 2748 3941
rect 2742 3936 2743 3940
rect 2747 3936 2748 3940
rect 2742 3935 2748 3936
rect 2942 3940 2948 3941
rect 2942 3936 2943 3940
rect 2947 3936 2948 3940
rect 2942 3935 2948 3936
rect 3134 3940 3140 3941
rect 3134 3936 3135 3940
rect 3139 3936 3140 3940
rect 3134 3935 3140 3936
rect 3318 3940 3324 3941
rect 3318 3936 3319 3940
rect 3323 3936 3324 3940
rect 3318 3935 3324 3936
rect 3510 3940 3516 3941
rect 3510 3936 3511 3940
rect 3515 3936 3516 3940
rect 3510 3935 3516 3936
rect 3678 3940 3684 3941
rect 3678 3936 3679 3940
rect 3683 3936 3684 3940
rect 3798 3937 3799 3941
rect 3803 3937 3804 3941
rect 3798 3936 3804 3937
rect 3678 3935 3684 3936
rect 2714 3925 2720 3926
rect 2714 3921 2715 3925
rect 2719 3921 2720 3925
rect 2714 3920 2720 3921
rect 2914 3925 2920 3926
rect 2914 3921 2915 3925
rect 2919 3921 2920 3925
rect 2914 3920 2920 3921
rect 3106 3925 3112 3926
rect 3106 3921 3107 3925
rect 3111 3921 3112 3925
rect 3106 3920 3112 3921
rect 3290 3925 3296 3926
rect 3290 3921 3291 3925
rect 3295 3921 3296 3925
rect 3290 3920 3296 3921
rect 3482 3925 3488 3926
rect 3482 3921 3483 3925
rect 3487 3921 3488 3925
rect 3482 3920 3488 3921
rect 3650 3925 3656 3926
rect 3650 3921 3651 3925
rect 3655 3921 3656 3925
rect 3650 3920 3656 3921
rect 3798 3924 3804 3925
rect 3798 3920 3799 3924
rect 3803 3920 3804 3924
rect 2550 3875 2556 3876
rect 2550 3871 2551 3875
rect 2555 3871 2556 3875
rect 2550 3870 2556 3871
rect 2716 3847 2718 3920
rect 2916 3847 2918 3920
rect 3042 3915 3048 3916
rect 3042 3911 3043 3915
rect 3047 3911 3048 3915
rect 3042 3910 3048 3911
rect 3044 3876 3046 3910
rect 3010 3875 3016 3876
rect 3010 3871 3011 3875
rect 3015 3871 3016 3875
rect 3010 3870 3016 3871
rect 3042 3875 3048 3876
rect 3042 3871 3043 3875
rect 3047 3871 3048 3875
rect 3042 3870 3048 3871
rect 2299 3846 2303 3847
rect 2299 3841 2303 3842
rect 2371 3846 2375 3847
rect 2371 3841 2375 3842
rect 2507 3846 2511 3847
rect 2507 3841 2511 3842
rect 2587 3846 2591 3847
rect 2587 3841 2591 3842
rect 2715 3846 2719 3847
rect 2715 3841 2719 3842
rect 2795 3846 2799 3847
rect 2795 3841 2799 3842
rect 2915 3846 2919 3847
rect 2915 3841 2919 3842
rect 2995 3846 2999 3847
rect 2995 3841 2999 3842
rect 2214 3831 2220 3832
rect 2214 3827 2215 3831
rect 2219 3827 2220 3831
rect 2214 3826 2220 3827
rect 2372 3780 2374 3841
rect 2378 3827 2384 3828
rect 2378 3823 2379 3827
rect 2383 3823 2384 3827
rect 2378 3822 2384 3823
rect 2380 3788 2382 3822
rect 2378 3787 2384 3788
rect 2378 3783 2379 3787
rect 2383 3783 2384 3787
rect 2378 3782 2384 3783
rect 2390 3787 2396 3788
rect 2390 3783 2391 3787
rect 2395 3783 2396 3787
rect 2390 3782 2396 3783
rect 1190 3776 1191 3780
rect 1195 3776 1196 3780
rect 1190 3775 1196 3776
rect 1934 3779 1940 3780
rect 1934 3775 1935 3779
rect 1939 3775 1940 3779
rect 1974 3776 1975 3780
rect 1979 3776 1980 3780
rect 1974 3775 1980 3776
rect 2138 3779 2144 3780
rect 2138 3775 2139 3779
rect 2143 3775 2144 3779
rect 1192 3751 1194 3775
rect 1934 3774 1940 3775
rect 2138 3774 2144 3775
rect 2370 3779 2376 3780
rect 2370 3775 2371 3779
rect 2375 3775 2376 3779
rect 2370 3774 2376 3775
rect 1936 3751 1938 3774
rect 2166 3764 2172 3765
rect 1974 3763 1980 3764
rect 1974 3759 1975 3763
rect 1979 3759 1980 3763
rect 2166 3760 2167 3764
rect 2171 3760 2172 3764
rect 2166 3759 2172 3760
rect 1974 3758 1980 3759
rect 1191 3750 1195 3751
rect 1191 3745 1195 3746
rect 1215 3750 1219 3751
rect 1215 3745 1219 3746
rect 1367 3750 1371 3751
rect 1367 3745 1371 3746
rect 1519 3750 1523 3751
rect 1519 3745 1523 3746
rect 1679 3750 1683 3751
rect 1679 3745 1683 3746
rect 1815 3750 1819 3751
rect 1815 3745 1819 3746
rect 1935 3750 1939 3751
rect 1935 3745 1939 3746
rect 1216 3721 1218 3745
rect 1368 3721 1370 3745
rect 1520 3721 1522 3745
rect 1680 3721 1682 3745
rect 1816 3721 1818 3745
rect 1936 3722 1938 3745
rect 1976 3731 1978 3758
rect 2168 3731 2170 3759
rect 1975 3730 1979 3731
rect 1975 3725 1979 3726
rect 2167 3730 2171 3731
rect 2167 3725 2171 3726
rect 2279 3730 2283 3731
rect 2279 3725 2283 3726
rect 1934 3721 1940 3722
rect 1214 3720 1220 3721
rect 1214 3716 1215 3720
rect 1219 3716 1220 3720
rect 1214 3715 1220 3716
rect 1366 3720 1372 3721
rect 1366 3716 1367 3720
rect 1371 3716 1372 3720
rect 1366 3715 1372 3716
rect 1518 3720 1524 3721
rect 1518 3716 1519 3720
rect 1523 3716 1524 3720
rect 1518 3715 1524 3716
rect 1678 3720 1684 3721
rect 1678 3716 1679 3720
rect 1683 3716 1684 3720
rect 1678 3715 1684 3716
rect 1814 3720 1820 3721
rect 1814 3716 1815 3720
rect 1819 3716 1820 3720
rect 1934 3717 1935 3721
rect 1939 3717 1940 3721
rect 1934 3716 1940 3717
rect 1814 3715 1820 3716
rect 1186 3705 1192 3706
rect 1186 3701 1187 3705
rect 1191 3701 1192 3705
rect 1186 3700 1192 3701
rect 1338 3705 1344 3706
rect 1338 3701 1339 3705
rect 1343 3701 1344 3705
rect 1338 3700 1344 3701
rect 1490 3705 1496 3706
rect 1490 3701 1491 3705
rect 1495 3701 1496 3705
rect 1490 3700 1496 3701
rect 1650 3705 1656 3706
rect 1650 3701 1651 3705
rect 1655 3701 1656 3705
rect 1650 3700 1656 3701
rect 1786 3705 1792 3706
rect 1786 3701 1787 3705
rect 1791 3701 1792 3705
rect 1786 3700 1792 3701
rect 1934 3704 1940 3705
rect 1934 3700 1935 3704
rect 1939 3700 1940 3704
rect 1976 3702 1978 3725
rect 1130 3695 1136 3696
rect 1130 3691 1131 3695
rect 1135 3691 1136 3695
rect 1130 3690 1136 3691
rect 1150 3695 1156 3696
rect 1150 3691 1151 3695
rect 1155 3691 1156 3695
rect 1150 3690 1156 3691
rect 1132 3656 1134 3690
rect 1122 3655 1128 3656
rect 1122 3651 1123 3655
rect 1127 3651 1128 3655
rect 1122 3650 1128 3651
rect 1130 3655 1136 3656
rect 1130 3651 1131 3655
rect 1135 3651 1136 3655
rect 1130 3650 1136 3651
rect 307 3626 311 3627
rect 307 3621 311 3622
rect 355 3626 359 3627
rect 355 3621 359 3622
rect 499 3626 503 3627
rect 499 3621 503 3622
rect 571 3626 575 3627
rect 571 3621 575 3622
rect 683 3626 687 3627
rect 683 3621 687 3622
rect 803 3626 807 3627
rect 803 3621 807 3622
rect 859 3626 863 3627
rect 859 3621 863 3622
rect 1027 3626 1031 3627
rect 1027 3621 1031 3622
rect 1043 3626 1047 3627
rect 1043 3621 1047 3622
rect 242 3611 248 3612
rect 242 3607 243 3611
rect 247 3607 248 3611
rect 242 3606 248 3607
rect 356 3560 358 3621
rect 362 3607 368 3608
rect 362 3603 363 3607
rect 367 3603 368 3607
rect 362 3602 368 3603
rect 364 3568 366 3602
rect 362 3567 368 3568
rect 362 3563 363 3567
rect 367 3563 368 3567
rect 362 3562 368 3563
rect 572 3560 574 3621
rect 578 3607 584 3608
rect 578 3603 579 3607
rect 583 3603 584 3607
rect 578 3602 584 3603
rect 580 3568 582 3602
rect 578 3567 584 3568
rect 578 3563 579 3567
rect 583 3563 584 3567
rect 578 3562 584 3563
rect 804 3560 806 3621
rect 810 3607 816 3608
rect 810 3603 811 3607
rect 815 3603 816 3607
rect 810 3602 816 3603
rect 812 3568 814 3602
rect 810 3567 816 3568
rect 810 3563 811 3567
rect 815 3563 816 3567
rect 810 3562 816 3563
rect 926 3567 932 3568
rect 926 3563 927 3567
rect 931 3563 932 3567
rect 926 3562 932 3563
rect 110 3556 111 3560
rect 115 3556 116 3560
rect 110 3555 116 3556
rect 146 3559 152 3560
rect 146 3555 147 3559
rect 151 3555 152 3559
rect 146 3554 152 3555
rect 354 3559 360 3560
rect 354 3555 355 3559
rect 359 3555 360 3559
rect 354 3554 360 3555
rect 570 3559 576 3560
rect 570 3555 571 3559
rect 575 3555 576 3559
rect 570 3554 576 3555
rect 802 3559 808 3560
rect 802 3555 803 3559
rect 807 3555 808 3559
rect 802 3554 808 3555
rect 174 3544 180 3545
rect 110 3543 116 3544
rect 110 3539 111 3543
rect 115 3539 116 3543
rect 174 3540 175 3544
rect 179 3540 180 3544
rect 174 3539 180 3540
rect 382 3544 388 3545
rect 382 3540 383 3544
rect 387 3540 388 3544
rect 382 3539 388 3540
rect 598 3544 604 3545
rect 598 3540 599 3544
rect 603 3540 604 3544
rect 598 3539 604 3540
rect 830 3544 836 3545
rect 830 3540 831 3544
rect 835 3540 836 3544
rect 830 3539 836 3540
rect 110 3538 116 3539
rect 112 3491 114 3538
rect 176 3491 178 3539
rect 384 3491 386 3539
rect 600 3491 602 3539
rect 832 3491 834 3539
rect 111 3490 115 3491
rect 111 3485 115 3486
rect 175 3490 179 3491
rect 175 3485 179 3486
rect 303 3490 307 3491
rect 303 3485 307 3486
rect 383 3490 387 3491
rect 383 3485 387 3486
rect 447 3490 451 3491
rect 447 3485 451 3486
rect 599 3490 603 3491
rect 599 3485 603 3486
rect 759 3490 763 3491
rect 759 3485 763 3486
rect 831 3490 835 3491
rect 831 3485 835 3486
rect 112 3462 114 3485
rect 110 3461 116 3462
rect 304 3461 306 3485
rect 448 3461 450 3485
rect 600 3461 602 3485
rect 760 3461 762 3485
rect 110 3457 111 3461
rect 115 3457 116 3461
rect 110 3456 116 3457
rect 302 3460 308 3461
rect 302 3456 303 3460
rect 307 3456 308 3460
rect 302 3455 308 3456
rect 446 3460 452 3461
rect 446 3456 447 3460
rect 451 3456 452 3460
rect 446 3455 452 3456
rect 598 3460 604 3461
rect 598 3456 599 3460
rect 603 3456 604 3460
rect 598 3455 604 3456
rect 758 3460 764 3461
rect 758 3456 759 3460
rect 763 3456 764 3460
rect 758 3455 764 3456
rect 274 3445 280 3446
rect 110 3444 116 3445
rect 110 3440 111 3444
rect 115 3440 116 3444
rect 274 3441 275 3445
rect 279 3441 280 3445
rect 274 3440 280 3441
rect 418 3445 424 3446
rect 418 3441 419 3445
rect 423 3441 424 3445
rect 418 3440 424 3441
rect 570 3445 576 3446
rect 570 3441 571 3445
rect 575 3441 576 3445
rect 570 3440 576 3441
rect 730 3445 736 3446
rect 730 3441 731 3445
rect 735 3441 736 3445
rect 730 3440 736 3441
rect 906 3445 912 3446
rect 906 3441 907 3445
rect 911 3441 912 3445
rect 906 3440 912 3441
rect 110 3439 116 3440
rect 112 3363 114 3439
rect 276 3363 278 3440
rect 402 3435 408 3436
rect 402 3431 403 3435
rect 407 3431 408 3435
rect 402 3430 408 3431
rect 404 3396 406 3430
rect 402 3395 408 3396
rect 402 3391 403 3395
rect 407 3391 408 3395
rect 402 3390 408 3391
rect 420 3363 422 3440
rect 546 3435 552 3436
rect 546 3431 547 3435
rect 551 3431 552 3435
rect 546 3430 552 3431
rect 548 3396 550 3430
rect 546 3395 552 3396
rect 546 3391 547 3395
rect 551 3391 552 3395
rect 546 3390 552 3391
rect 572 3363 574 3440
rect 718 3435 724 3436
rect 718 3431 719 3435
rect 723 3431 724 3435
rect 718 3430 724 3431
rect 720 3396 722 3430
rect 718 3395 724 3396
rect 718 3391 719 3395
rect 723 3391 724 3395
rect 718 3390 724 3391
rect 732 3363 734 3440
rect 762 3435 768 3436
rect 762 3431 763 3435
rect 767 3431 768 3435
rect 762 3430 768 3431
rect 111 3362 115 3363
rect 111 3357 115 3358
rect 275 3362 279 3363
rect 275 3357 279 3358
rect 419 3362 423 3363
rect 419 3357 423 3358
rect 467 3362 471 3363
rect 467 3357 471 3358
rect 571 3362 575 3363
rect 571 3357 575 3358
rect 667 3362 671 3363
rect 667 3357 671 3358
rect 731 3362 735 3363
rect 731 3357 735 3358
rect 112 3297 114 3357
rect 110 3296 116 3297
rect 468 3296 470 3357
rect 562 3343 568 3344
rect 562 3339 563 3343
rect 567 3339 568 3343
rect 562 3338 568 3339
rect 110 3292 111 3296
rect 115 3292 116 3296
rect 110 3291 116 3292
rect 466 3295 472 3296
rect 466 3291 467 3295
rect 471 3291 472 3295
rect 466 3290 472 3291
rect 494 3280 500 3281
rect 110 3279 116 3280
rect 110 3275 111 3279
rect 115 3275 116 3279
rect 494 3276 495 3280
rect 499 3276 500 3280
rect 494 3275 500 3276
rect 110 3274 116 3275
rect 112 3251 114 3274
rect 496 3251 498 3275
rect 111 3250 115 3251
rect 111 3245 115 3246
rect 495 3250 499 3251
rect 495 3245 499 3246
rect 535 3250 539 3251
rect 535 3245 539 3246
rect 112 3222 114 3245
rect 110 3221 116 3222
rect 536 3221 538 3245
rect 110 3217 111 3221
rect 115 3217 116 3221
rect 110 3216 116 3217
rect 534 3220 540 3221
rect 534 3216 535 3220
rect 539 3216 540 3220
rect 534 3215 540 3216
rect 506 3205 512 3206
rect 110 3204 116 3205
rect 110 3200 111 3204
rect 115 3200 116 3204
rect 506 3201 507 3205
rect 511 3201 512 3205
rect 506 3200 512 3201
rect 110 3199 116 3200
rect 112 3131 114 3199
rect 508 3131 510 3200
rect 564 3196 566 3338
rect 668 3296 670 3357
rect 764 3348 766 3430
rect 834 3395 840 3396
rect 834 3391 835 3395
rect 839 3391 840 3395
rect 834 3390 840 3391
rect 762 3347 768 3348
rect 762 3343 763 3347
rect 767 3343 768 3347
rect 762 3342 768 3343
rect 836 3312 838 3390
rect 908 3363 910 3440
rect 928 3388 930 3562
rect 1044 3560 1046 3621
rect 1124 3568 1126 3650
rect 1188 3627 1190 3700
rect 1314 3695 1320 3696
rect 1314 3691 1315 3695
rect 1319 3691 1320 3695
rect 1314 3690 1320 3691
rect 1316 3656 1318 3690
rect 1314 3655 1320 3656
rect 1314 3651 1315 3655
rect 1319 3651 1320 3655
rect 1314 3650 1320 3651
rect 1340 3627 1342 3700
rect 1466 3695 1472 3696
rect 1466 3691 1467 3695
rect 1471 3691 1472 3695
rect 1466 3690 1472 3691
rect 1468 3656 1470 3690
rect 1466 3655 1472 3656
rect 1466 3651 1467 3655
rect 1471 3651 1472 3655
rect 1466 3650 1472 3651
rect 1414 3647 1420 3648
rect 1414 3643 1415 3647
rect 1419 3643 1420 3647
rect 1414 3642 1420 3643
rect 1187 3626 1191 3627
rect 1187 3621 1191 3622
rect 1291 3626 1295 3627
rect 1291 3621 1295 3622
rect 1339 3626 1343 3627
rect 1339 3621 1343 3622
rect 1138 3607 1144 3608
rect 1138 3603 1139 3607
rect 1143 3603 1144 3607
rect 1138 3602 1144 3603
rect 1122 3567 1128 3568
rect 1122 3563 1123 3567
rect 1127 3563 1128 3567
rect 1122 3562 1128 3563
rect 1042 3559 1048 3560
rect 1042 3555 1043 3559
rect 1047 3555 1048 3559
rect 1042 3554 1048 3555
rect 1070 3544 1076 3545
rect 1070 3540 1071 3544
rect 1075 3540 1076 3544
rect 1070 3539 1076 3540
rect 1072 3491 1074 3539
rect 935 3490 939 3491
rect 935 3485 939 3486
rect 1071 3490 1075 3491
rect 1071 3485 1075 3486
rect 1111 3490 1115 3491
rect 1111 3485 1115 3486
rect 936 3461 938 3485
rect 1112 3461 1114 3485
rect 934 3460 940 3461
rect 934 3456 935 3460
rect 939 3456 940 3460
rect 934 3455 940 3456
rect 1110 3460 1116 3461
rect 1110 3456 1111 3460
rect 1115 3456 1116 3460
rect 1110 3455 1116 3456
rect 1082 3445 1088 3446
rect 1082 3441 1083 3445
rect 1087 3441 1088 3445
rect 1082 3440 1088 3441
rect 1034 3435 1040 3436
rect 1034 3431 1035 3435
rect 1039 3431 1040 3435
rect 1034 3430 1040 3431
rect 1036 3396 1038 3430
rect 1034 3395 1040 3396
rect 1034 3391 1035 3395
rect 1039 3391 1040 3395
rect 1034 3390 1040 3391
rect 926 3387 932 3388
rect 926 3383 927 3387
rect 931 3383 932 3387
rect 926 3382 932 3383
rect 1084 3363 1086 3440
rect 1140 3436 1142 3602
rect 1292 3560 1294 3621
rect 1416 3568 1418 3642
rect 1492 3627 1494 3700
rect 1638 3695 1644 3696
rect 1638 3691 1639 3695
rect 1643 3691 1644 3695
rect 1638 3690 1644 3691
rect 1640 3656 1642 3690
rect 1638 3655 1644 3656
rect 1638 3651 1639 3655
rect 1643 3651 1644 3655
rect 1638 3650 1644 3651
rect 1652 3627 1654 3700
rect 1778 3695 1784 3696
rect 1778 3691 1779 3695
rect 1783 3691 1784 3695
rect 1778 3690 1784 3691
rect 1780 3656 1782 3690
rect 1778 3655 1784 3656
rect 1778 3651 1779 3655
rect 1783 3651 1784 3655
rect 1778 3650 1784 3651
rect 1788 3627 1790 3700
rect 1934 3699 1940 3700
rect 1974 3701 1980 3702
rect 2280 3701 2282 3725
rect 1882 3695 1888 3696
rect 1882 3691 1883 3695
rect 1887 3691 1888 3695
rect 1882 3690 1888 3691
rect 1491 3626 1495 3627
rect 1491 3621 1495 3622
rect 1547 3626 1551 3627
rect 1547 3621 1551 3622
rect 1651 3626 1655 3627
rect 1651 3621 1655 3622
rect 1787 3626 1791 3627
rect 1787 3621 1791 3622
rect 1414 3567 1420 3568
rect 1414 3563 1415 3567
rect 1419 3563 1420 3567
rect 1414 3562 1420 3563
rect 1548 3560 1550 3621
rect 1670 3619 1676 3620
rect 1670 3615 1671 3619
rect 1675 3615 1676 3619
rect 1670 3614 1676 3615
rect 1582 3611 1588 3612
rect 1582 3607 1583 3611
rect 1587 3607 1588 3611
rect 1582 3606 1588 3607
rect 1290 3559 1296 3560
rect 1290 3555 1291 3559
rect 1295 3555 1296 3559
rect 1290 3554 1296 3555
rect 1546 3559 1552 3560
rect 1546 3555 1547 3559
rect 1551 3555 1552 3559
rect 1546 3554 1552 3555
rect 1318 3544 1324 3545
rect 1318 3540 1319 3544
rect 1323 3540 1324 3544
rect 1318 3539 1324 3540
rect 1574 3544 1580 3545
rect 1574 3540 1575 3544
rect 1579 3540 1580 3544
rect 1574 3539 1580 3540
rect 1320 3491 1322 3539
rect 1576 3491 1578 3539
rect 1295 3490 1299 3491
rect 1295 3485 1299 3486
rect 1319 3490 1323 3491
rect 1319 3485 1323 3486
rect 1487 3490 1491 3491
rect 1487 3485 1491 3486
rect 1575 3490 1579 3491
rect 1575 3485 1579 3486
rect 1296 3461 1298 3485
rect 1488 3461 1490 3485
rect 1294 3460 1300 3461
rect 1294 3456 1295 3460
rect 1299 3456 1300 3460
rect 1294 3455 1300 3456
rect 1486 3460 1492 3461
rect 1486 3456 1487 3460
rect 1491 3456 1492 3460
rect 1486 3455 1492 3456
rect 1266 3445 1272 3446
rect 1266 3441 1267 3445
rect 1271 3441 1272 3445
rect 1266 3440 1272 3441
rect 1458 3445 1464 3446
rect 1458 3441 1459 3445
rect 1463 3441 1464 3445
rect 1458 3440 1464 3441
rect 1138 3435 1144 3436
rect 1138 3431 1139 3435
rect 1143 3431 1144 3435
rect 1138 3430 1144 3431
rect 1268 3363 1270 3440
rect 1394 3435 1400 3436
rect 1394 3431 1395 3435
rect 1399 3431 1400 3435
rect 1394 3430 1400 3431
rect 1396 3396 1398 3430
rect 1362 3395 1368 3396
rect 1362 3391 1363 3395
rect 1367 3391 1368 3395
rect 1362 3390 1368 3391
rect 1394 3395 1400 3396
rect 1394 3391 1395 3395
rect 1399 3391 1400 3395
rect 1394 3390 1400 3391
rect 875 3362 879 3363
rect 875 3357 879 3358
rect 907 3362 911 3363
rect 907 3357 911 3358
rect 1083 3362 1087 3363
rect 1083 3357 1087 3358
rect 1091 3362 1095 3363
rect 1091 3357 1095 3358
rect 1267 3362 1271 3363
rect 1267 3357 1271 3358
rect 1315 3362 1319 3363
rect 1315 3357 1319 3358
rect 834 3311 840 3312
rect 834 3307 835 3311
rect 839 3307 840 3311
rect 834 3306 840 3307
rect 876 3296 878 3357
rect 882 3343 888 3344
rect 882 3339 883 3343
rect 887 3339 888 3343
rect 882 3338 888 3339
rect 884 3304 886 3338
rect 882 3303 888 3304
rect 882 3299 883 3303
rect 887 3299 888 3303
rect 882 3298 888 3299
rect 1092 3296 1094 3357
rect 1098 3343 1104 3344
rect 1098 3339 1099 3343
rect 1103 3339 1104 3343
rect 1098 3338 1104 3339
rect 1100 3304 1102 3338
rect 1098 3303 1104 3304
rect 1098 3299 1099 3303
rect 1103 3299 1104 3303
rect 1098 3298 1104 3299
rect 1154 3303 1160 3304
rect 1154 3299 1155 3303
rect 1159 3299 1160 3303
rect 1154 3298 1160 3299
rect 666 3295 672 3296
rect 666 3291 667 3295
rect 671 3291 672 3295
rect 666 3290 672 3291
rect 874 3295 880 3296
rect 874 3291 875 3295
rect 879 3291 880 3295
rect 874 3290 880 3291
rect 1090 3295 1096 3296
rect 1090 3291 1091 3295
rect 1095 3291 1096 3295
rect 1090 3290 1096 3291
rect 694 3280 700 3281
rect 694 3276 695 3280
rect 699 3276 700 3280
rect 694 3275 700 3276
rect 902 3280 908 3281
rect 902 3276 903 3280
rect 907 3276 908 3280
rect 902 3275 908 3276
rect 1118 3280 1124 3281
rect 1118 3276 1119 3280
rect 1123 3276 1124 3280
rect 1118 3275 1124 3276
rect 696 3251 698 3275
rect 904 3251 906 3275
rect 1120 3251 1122 3275
rect 695 3250 699 3251
rect 695 3245 699 3246
rect 727 3250 731 3251
rect 727 3245 731 3246
rect 903 3250 907 3251
rect 903 3245 907 3246
rect 919 3250 923 3251
rect 919 3245 923 3246
rect 1111 3250 1115 3251
rect 1111 3245 1115 3246
rect 1119 3250 1123 3251
rect 1119 3245 1123 3246
rect 728 3221 730 3245
rect 920 3221 922 3245
rect 1112 3221 1114 3245
rect 726 3220 732 3221
rect 726 3216 727 3220
rect 731 3216 732 3220
rect 726 3215 732 3216
rect 918 3220 924 3221
rect 918 3216 919 3220
rect 923 3216 924 3220
rect 918 3215 924 3216
rect 1110 3220 1116 3221
rect 1110 3216 1111 3220
rect 1115 3216 1116 3220
rect 1110 3215 1116 3216
rect 698 3205 704 3206
rect 698 3201 699 3205
rect 703 3201 704 3205
rect 698 3200 704 3201
rect 890 3205 896 3206
rect 890 3201 891 3205
rect 895 3201 896 3205
rect 890 3200 896 3201
rect 1082 3205 1088 3206
rect 1082 3201 1083 3205
rect 1087 3201 1088 3205
rect 1082 3200 1088 3201
rect 562 3195 568 3196
rect 562 3191 563 3195
rect 567 3191 568 3195
rect 562 3190 568 3191
rect 658 3195 664 3196
rect 658 3191 659 3195
rect 663 3191 664 3195
rect 658 3190 664 3191
rect 550 3155 556 3156
rect 550 3151 551 3155
rect 555 3151 556 3155
rect 550 3150 556 3151
rect 111 3130 115 3131
rect 111 3125 115 3126
rect 427 3130 431 3131
rect 427 3125 431 3126
rect 507 3130 511 3131
rect 507 3125 511 3126
rect 112 3065 114 3125
rect 110 3064 116 3065
rect 428 3064 430 3125
rect 434 3111 440 3112
rect 434 3107 435 3111
rect 439 3107 440 3111
rect 434 3106 440 3107
rect 110 3060 111 3064
rect 115 3060 116 3064
rect 110 3059 116 3060
rect 426 3063 432 3064
rect 426 3059 427 3063
rect 431 3059 432 3063
rect 426 3058 432 3059
rect 110 3047 116 3048
rect 110 3043 111 3047
rect 115 3043 116 3047
rect 110 3042 116 3043
rect 112 2991 114 3042
rect 111 2990 115 2991
rect 111 2985 115 2986
rect 199 2990 203 2991
rect 199 2985 203 2986
rect 112 2962 114 2985
rect 110 2961 116 2962
rect 200 2961 202 2985
rect 110 2957 111 2961
rect 115 2957 116 2961
rect 110 2956 116 2957
rect 198 2960 204 2961
rect 198 2956 199 2960
rect 203 2956 204 2960
rect 198 2955 204 2956
rect 170 2945 176 2946
rect 110 2944 116 2945
rect 110 2940 111 2944
rect 115 2940 116 2944
rect 170 2941 171 2945
rect 175 2941 176 2945
rect 170 2940 176 2941
rect 110 2939 116 2940
rect 112 2879 114 2939
rect 172 2879 174 2940
rect 436 2936 438 3106
rect 552 3072 554 3150
rect 563 3130 567 3131
rect 563 3125 567 3126
rect 550 3071 556 3072
rect 550 3067 551 3071
rect 555 3067 556 3071
rect 550 3066 556 3067
rect 564 3064 566 3125
rect 660 3116 662 3190
rect 700 3131 702 3200
rect 892 3131 894 3200
rect 1084 3131 1086 3200
rect 1156 3148 1158 3298
rect 1316 3296 1318 3357
rect 1364 3304 1366 3390
rect 1460 3363 1462 3440
rect 1584 3436 1586 3606
rect 1672 3568 1674 3614
rect 1670 3567 1676 3568
rect 1670 3563 1671 3567
rect 1675 3563 1676 3567
rect 1670 3562 1676 3563
rect 1788 3560 1790 3621
rect 1884 3612 1886 3690
rect 1936 3627 1938 3699
rect 1974 3697 1975 3701
rect 1979 3697 1980 3701
rect 1974 3696 1980 3697
rect 2278 3700 2284 3701
rect 2278 3696 2279 3700
rect 2283 3696 2284 3700
rect 2278 3695 2284 3696
rect 2250 3685 2256 3686
rect 1974 3684 1980 3685
rect 1974 3680 1975 3684
rect 1979 3680 1980 3684
rect 2250 3681 2251 3685
rect 2255 3681 2256 3685
rect 2250 3680 2256 3681
rect 1974 3679 1980 3680
rect 1935 3626 1939 3627
rect 1935 3621 1939 3622
rect 1882 3611 1888 3612
rect 1882 3607 1883 3611
rect 1887 3607 1888 3611
rect 1882 3606 1888 3607
rect 1922 3591 1928 3592
rect 1922 3587 1923 3591
rect 1927 3587 1928 3591
rect 1922 3586 1928 3587
rect 1924 3568 1926 3586
rect 1922 3567 1928 3568
rect 1922 3563 1923 3567
rect 1927 3563 1928 3567
rect 1922 3562 1928 3563
rect 1936 3561 1938 3621
rect 1976 3607 1978 3679
rect 2252 3607 2254 3680
rect 2346 3675 2352 3676
rect 2346 3671 2347 3675
rect 2351 3671 2352 3675
rect 2346 3670 2352 3671
rect 1975 3606 1979 3607
rect 1975 3601 1979 3602
rect 1995 3606 1999 3607
rect 1995 3601 1999 3602
rect 2251 3606 2255 3607
rect 2251 3601 2255 3602
rect 1934 3560 1940 3561
rect 1786 3559 1792 3560
rect 1786 3555 1787 3559
rect 1791 3555 1792 3559
rect 1934 3556 1935 3560
rect 1939 3556 1940 3560
rect 1934 3555 1940 3556
rect 1786 3554 1792 3555
rect 1814 3544 1820 3545
rect 1814 3540 1815 3544
rect 1819 3540 1820 3544
rect 1814 3539 1820 3540
rect 1934 3543 1940 3544
rect 1934 3539 1935 3543
rect 1939 3539 1940 3543
rect 1976 3541 1978 3601
rect 1816 3491 1818 3539
rect 1934 3538 1940 3539
rect 1974 3540 1980 3541
rect 1996 3540 1998 3601
rect 2090 3547 2096 3548
rect 2090 3543 2091 3547
rect 2095 3543 2096 3547
rect 2090 3542 2096 3543
rect 1936 3491 1938 3538
rect 1974 3536 1975 3540
rect 1979 3536 1980 3540
rect 1974 3535 1980 3536
rect 1994 3539 2000 3540
rect 1994 3535 1995 3539
rect 1999 3535 2000 3539
rect 1994 3534 2000 3535
rect 2022 3524 2028 3525
rect 1974 3523 1980 3524
rect 1974 3519 1975 3523
rect 1979 3519 1980 3523
rect 2022 3520 2023 3524
rect 2027 3520 2028 3524
rect 2022 3519 2028 3520
rect 1974 3518 1980 3519
rect 1815 3490 1819 3491
rect 1815 3485 1819 3486
rect 1935 3490 1939 3491
rect 1976 3487 1978 3518
rect 2024 3487 2026 3519
rect 1935 3485 1939 3486
rect 1975 3486 1979 3487
rect 1936 3462 1938 3485
rect 1975 3481 1979 3482
rect 2023 3486 2027 3487
rect 2023 3481 2027 3482
rect 1934 3461 1940 3462
rect 1934 3457 1935 3461
rect 1939 3457 1940 3461
rect 1976 3458 1978 3481
rect 1934 3456 1940 3457
rect 1974 3457 1980 3458
rect 2024 3457 2026 3481
rect 1974 3453 1975 3457
rect 1979 3453 1980 3457
rect 1974 3452 1980 3453
rect 2022 3456 2028 3457
rect 2022 3452 2023 3456
rect 2027 3452 2028 3456
rect 2022 3451 2028 3452
rect 1934 3444 1940 3445
rect 1934 3440 1935 3444
rect 1939 3440 1940 3444
rect 1994 3441 2000 3442
rect 1934 3439 1940 3440
rect 1974 3440 1980 3441
rect 1582 3435 1588 3436
rect 1582 3431 1583 3435
rect 1587 3431 1588 3435
rect 1582 3430 1588 3431
rect 1936 3363 1938 3439
rect 1974 3436 1975 3440
rect 1979 3436 1980 3440
rect 1994 3437 1995 3441
rect 1999 3437 2000 3441
rect 1994 3436 2000 3437
rect 1974 3435 1980 3436
rect 1459 3362 1463 3363
rect 1459 3357 1463 3358
rect 1935 3362 1939 3363
rect 1935 3357 1939 3358
rect 1390 3347 1396 3348
rect 1390 3343 1391 3347
rect 1395 3343 1396 3347
rect 1390 3342 1396 3343
rect 1362 3303 1368 3304
rect 1362 3299 1363 3303
rect 1367 3299 1368 3303
rect 1362 3298 1368 3299
rect 1314 3295 1320 3296
rect 1314 3291 1315 3295
rect 1319 3291 1320 3295
rect 1314 3290 1320 3291
rect 1342 3280 1348 3281
rect 1342 3276 1343 3280
rect 1347 3276 1348 3280
rect 1342 3275 1348 3276
rect 1344 3251 1346 3275
rect 1295 3250 1299 3251
rect 1295 3245 1299 3246
rect 1343 3250 1347 3251
rect 1343 3245 1347 3246
rect 1296 3221 1298 3245
rect 1294 3220 1300 3221
rect 1294 3216 1295 3220
rect 1299 3216 1300 3220
rect 1294 3215 1300 3216
rect 1266 3205 1272 3206
rect 1266 3201 1267 3205
rect 1271 3201 1272 3205
rect 1266 3200 1272 3201
rect 1210 3195 1216 3196
rect 1210 3191 1211 3195
rect 1215 3191 1216 3195
rect 1210 3190 1216 3191
rect 1212 3156 1214 3190
rect 1210 3155 1216 3156
rect 1210 3151 1211 3155
rect 1215 3151 1216 3155
rect 1210 3150 1216 3151
rect 1154 3147 1160 3148
rect 1154 3143 1155 3147
rect 1159 3143 1160 3147
rect 1154 3142 1160 3143
rect 1268 3131 1270 3200
rect 1392 3196 1394 3342
rect 1936 3297 1938 3357
rect 1976 3335 1978 3435
rect 1996 3335 1998 3436
rect 2092 3392 2094 3542
rect 2252 3540 2254 3601
rect 2348 3592 2350 3670
rect 2392 3636 2394 3782
rect 2588 3780 2590 3841
rect 2594 3827 2600 3828
rect 2594 3823 2595 3827
rect 2599 3823 2600 3827
rect 2594 3822 2600 3823
rect 2586 3779 2592 3780
rect 2586 3775 2587 3779
rect 2591 3775 2592 3779
rect 2586 3774 2592 3775
rect 2398 3764 2404 3765
rect 2398 3760 2399 3764
rect 2403 3760 2404 3764
rect 2398 3759 2404 3760
rect 2400 3731 2402 3759
rect 2399 3730 2403 3731
rect 2399 3725 2403 3726
rect 2479 3730 2483 3731
rect 2479 3725 2483 3726
rect 2480 3701 2482 3725
rect 2478 3700 2484 3701
rect 2478 3696 2479 3700
rect 2483 3696 2484 3700
rect 2478 3695 2484 3696
rect 2450 3685 2456 3686
rect 2450 3681 2451 3685
rect 2455 3681 2456 3685
rect 2450 3680 2456 3681
rect 2390 3635 2396 3636
rect 2390 3631 2391 3635
rect 2395 3631 2396 3635
rect 2390 3630 2396 3631
rect 2452 3607 2454 3680
rect 2596 3676 2598 3822
rect 2796 3780 2798 3841
rect 2802 3827 2808 3828
rect 2802 3823 2803 3827
rect 2807 3823 2808 3827
rect 2802 3822 2808 3823
rect 2804 3788 2806 3822
rect 2802 3787 2808 3788
rect 2802 3783 2803 3787
rect 2807 3783 2808 3787
rect 2802 3782 2808 3783
rect 2996 3780 2998 3841
rect 3012 3829 3014 3870
rect 3108 3847 3110 3920
rect 3234 3915 3240 3916
rect 3234 3911 3235 3915
rect 3239 3911 3240 3915
rect 3234 3910 3240 3911
rect 3236 3876 3238 3910
rect 3234 3875 3240 3876
rect 3234 3871 3235 3875
rect 3239 3871 3240 3875
rect 3234 3870 3240 3871
rect 3292 3847 3294 3920
rect 3418 3915 3424 3916
rect 3418 3911 3419 3915
rect 3423 3911 3424 3915
rect 3418 3910 3424 3911
rect 3420 3876 3422 3910
rect 3418 3875 3424 3876
rect 3418 3871 3419 3875
rect 3423 3871 3424 3875
rect 3418 3870 3424 3871
rect 3484 3847 3486 3920
rect 3610 3915 3616 3916
rect 3610 3911 3611 3915
rect 3615 3911 3616 3915
rect 3610 3910 3616 3911
rect 3612 3876 3614 3910
rect 3610 3875 3616 3876
rect 3610 3871 3611 3875
rect 3615 3871 3616 3875
rect 3610 3870 3616 3871
rect 3652 3847 3654 3920
rect 3798 3919 3804 3920
rect 3840 3919 3842 3966
rect 3800 3847 3802 3919
rect 3839 3918 3843 3919
rect 3868 3916 3870 4030
rect 4004 3988 4006 4049
rect 4010 4035 4016 4036
rect 4010 4031 4011 4035
rect 4015 4031 4016 4035
rect 4010 4030 4016 4031
rect 4012 3996 4014 4030
rect 4010 3995 4016 3996
rect 4010 3991 4011 3995
rect 4015 3991 4016 3995
rect 4010 3990 4016 3991
rect 4172 3988 4174 4049
rect 4178 4035 4184 4036
rect 4178 4031 4179 4035
rect 4183 4031 4184 4035
rect 4178 4030 4184 4031
rect 4180 3996 4182 4030
rect 4178 3995 4184 3996
rect 4178 3991 4179 3995
rect 4183 3991 4184 3995
rect 4178 3990 4184 3991
rect 4340 3988 4342 4049
rect 4450 3995 4456 3996
rect 4450 3991 4451 3995
rect 4455 3991 4456 3995
rect 4450 3990 4456 3991
rect 4002 3987 4008 3988
rect 4002 3983 4003 3987
rect 4007 3983 4008 3987
rect 4002 3982 4008 3983
rect 4170 3987 4176 3988
rect 4170 3983 4171 3987
rect 4175 3983 4176 3987
rect 4170 3982 4176 3983
rect 4338 3987 4344 3988
rect 4338 3983 4339 3987
rect 4343 3983 4344 3987
rect 4338 3982 4344 3983
rect 3886 3972 3892 3973
rect 3886 3968 3887 3972
rect 3891 3968 3892 3972
rect 3886 3967 3892 3968
rect 4030 3972 4036 3973
rect 4030 3968 4031 3972
rect 4035 3968 4036 3972
rect 4030 3967 4036 3968
rect 4198 3972 4204 3973
rect 4198 3968 4199 3972
rect 4203 3968 4204 3972
rect 4198 3967 4204 3968
rect 4366 3972 4372 3973
rect 4366 3968 4367 3972
rect 4371 3968 4372 3972
rect 4366 3967 4372 3968
rect 3888 3919 3890 3967
rect 4032 3919 4034 3967
rect 4200 3919 4202 3967
rect 4368 3919 4370 3967
rect 3887 3918 3891 3919
rect 3839 3913 3843 3914
rect 3866 3915 3872 3916
rect 3840 3890 3842 3913
rect 3866 3911 3867 3915
rect 3871 3911 3872 3915
rect 3887 3913 3891 3914
rect 4031 3918 4035 3919
rect 4031 3913 4035 3914
rect 4199 3918 4203 3919
rect 4199 3913 4203 3914
rect 4367 3918 4371 3919
rect 4367 3913 4371 3914
rect 4383 3918 4387 3919
rect 4383 3913 4387 3914
rect 3866 3910 3872 3911
rect 3838 3889 3844 3890
rect 4384 3889 4386 3913
rect 3838 3885 3839 3889
rect 3843 3885 3844 3889
rect 3838 3884 3844 3885
rect 4382 3888 4388 3889
rect 4382 3884 4383 3888
rect 4387 3884 4388 3888
rect 4382 3883 4388 3884
rect 4354 3873 4360 3874
rect 3838 3872 3844 3873
rect 3838 3868 3839 3872
rect 3843 3868 3844 3872
rect 4354 3869 4355 3873
rect 4359 3869 4360 3873
rect 4354 3868 4360 3869
rect 3838 3867 3844 3868
rect 3107 3846 3111 3847
rect 3107 3841 3111 3842
rect 3195 3846 3199 3847
rect 3195 3841 3199 3842
rect 3291 3846 3295 3847
rect 3291 3841 3295 3842
rect 3403 3846 3407 3847
rect 3403 3841 3407 3842
rect 3483 3846 3487 3847
rect 3483 3841 3487 3842
rect 3651 3846 3655 3847
rect 3651 3841 3655 3842
rect 3799 3846 3803 3847
rect 3799 3841 3803 3842
rect 3011 3828 3015 3829
rect 3002 3827 3008 3828
rect 3002 3823 3003 3827
rect 3007 3823 3008 3827
rect 3011 3823 3015 3824
rect 3002 3822 3008 3823
rect 3004 3788 3006 3822
rect 3002 3787 3008 3788
rect 3002 3783 3003 3787
rect 3007 3783 3008 3787
rect 3002 3782 3008 3783
rect 3196 3780 3198 3841
rect 3202 3827 3208 3828
rect 3202 3823 3203 3827
rect 3207 3823 3208 3827
rect 3202 3822 3208 3823
rect 3204 3788 3206 3822
rect 3202 3787 3208 3788
rect 3202 3783 3203 3787
rect 3207 3783 3208 3787
rect 3202 3782 3208 3783
rect 3404 3780 3406 3841
rect 3419 3828 3423 3829
rect 3410 3827 3416 3828
rect 3410 3823 3411 3827
rect 3415 3823 3416 3827
rect 3419 3823 3423 3824
rect 3410 3822 3416 3823
rect 3412 3788 3414 3822
rect 3420 3788 3422 3823
rect 3410 3787 3416 3788
rect 3410 3783 3411 3787
rect 3415 3783 3416 3787
rect 3410 3782 3416 3783
rect 3418 3787 3424 3788
rect 3418 3783 3419 3787
rect 3423 3783 3424 3787
rect 3418 3782 3424 3783
rect 3800 3781 3802 3841
rect 3840 3791 3842 3867
rect 4356 3791 4358 3868
rect 4452 3824 4454 3990
rect 4500 3988 4502 4049
rect 4652 3988 4654 4049
rect 4804 3988 4806 4049
rect 4948 3988 4950 4049
rect 5092 3988 5094 4049
rect 5236 3988 5238 4049
rect 5380 3988 5382 4049
rect 5398 4039 5404 4040
rect 5398 4035 5399 4039
rect 5403 4035 5404 4039
rect 5398 4034 5404 4035
rect 4498 3987 4504 3988
rect 4498 3983 4499 3987
rect 4503 3983 4504 3987
rect 4498 3982 4504 3983
rect 4650 3987 4656 3988
rect 4650 3983 4651 3987
rect 4655 3983 4656 3987
rect 4650 3982 4656 3983
rect 4802 3987 4808 3988
rect 4802 3983 4803 3987
rect 4807 3983 4808 3987
rect 4802 3982 4808 3983
rect 4946 3987 4952 3988
rect 4946 3983 4947 3987
rect 4951 3983 4952 3987
rect 4946 3982 4952 3983
rect 5090 3987 5096 3988
rect 5090 3983 5091 3987
rect 5095 3983 5096 3987
rect 5090 3982 5096 3983
rect 5234 3987 5240 3988
rect 5234 3983 5235 3987
rect 5239 3983 5240 3987
rect 5234 3982 5240 3983
rect 5378 3987 5384 3988
rect 5378 3983 5379 3987
rect 5383 3983 5384 3987
rect 5378 3982 5384 3983
rect 4526 3972 4532 3973
rect 4526 3968 4527 3972
rect 4531 3968 4532 3972
rect 4526 3967 4532 3968
rect 4678 3972 4684 3973
rect 4678 3968 4679 3972
rect 4683 3968 4684 3972
rect 4678 3967 4684 3968
rect 4830 3972 4836 3973
rect 4830 3968 4831 3972
rect 4835 3968 4836 3972
rect 4830 3967 4836 3968
rect 4974 3972 4980 3973
rect 4974 3968 4975 3972
rect 4979 3968 4980 3972
rect 4974 3967 4980 3968
rect 5118 3972 5124 3973
rect 5118 3968 5119 3972
rect 5123 3968 5124 3972
rect 5118 3967 5124 3968
rect 5262 3972 5268 3973
rect 5262 3968 5263 3972
rect 5267 3968 5268 3972
rect 5262 3967 5268 3968
rect 4528 3919 4530 3967
rect 4680 3919 4682 3967
rect 4832 3919 4834 3967
rect 4976 3919 4978 3967
rect 5120 3919 5122 3967
rect 5264 3919 5266 3967
rect 4527 3918 4531 3919
rect 4527 3913 4531 3914
rect 4599 3918 4603 3919
rect 4599 3913 4603 3914
rect 4679 3918 4683 3919
rect 4679 3913 4683 3914
rect 4823 3918 4827 3919
rect 4823 3913 4827 3914
rect 4831 3918 4835 3919
rect 4831 3913 4835 3914
rect 4975 3918 4979 3919
rect 4975 3913 4979 3914
rect 5063 3918 5067 3919
rect 5063 3913 5067 3914
rect 5119 3918 5123 3919
rect 5119 3913 5123 3914
rect 5263 3918 5267 3919
rect 5263 3913 5267 3914
rect 5311 3918 5315 3919
rect 5311 3913 5315 3914
rect 4600 3889 4602 3913
rect 4824 3889 4826 3913
rect 5064 3889 5066 3913
rect 5312 3889 5314 3913
rect 4598 3888 4604 3889
rect 4598 3884 4599 3888
rect 4603 3884 4604 3888
rect 4598 3883 4604 3884
rect 4822 3888 4828 3889
rect 4822 3884 4823 3888
rect 4827 3884 4828 3888
rect 4822 3883 4828 3884
rect 5062 3888 5068 3889
rect 5062 3884 5063 3888
rect 5067 3884 5068 3888
rect 5062 3883 5068 3884
rect 5310 3888 5316 3889
rect 5310 3884 5311 3888
rect 5315 3884 5316 3888
rect 5310 3883 5316 3884
rect 4570 3873 4576 3874
rect 4570 3869 4571 3873
rect 4575 3869 4576 3873
rect 4570 3868 4576 3869
rect 4794 3873 4800 3874
rect 4794 3869 4795 3873
rect 4799 3869 4800 3873
rect 4794 3868 4800 3869
rect 5034 3873 5040 3874
rect 5034 3869 5035 3873
rect 5039 3869 5040 3873
rect 5034 3868 5040 3869
rect 5282 3873 5288 3874
rect 5282 3869 5283 3873
rect 5287 3869 5288 3873
rect 5282 3868 5288 3869
rect 4482 3863 4488 3864
rect 4482 3859 4483 3863
rect 4487 3859 4488 3863
rect 4482 3858 4488 3859
rect 4484 3824 4486 3858
rect 4450 3823 4456 3824
rect 4450 3819 4451 3823
rect 4455 3819 4456 3823
rect 4450 3818 4456 3819
rect 4482 3823 4488 3824
rect 4482 3819 4483 3823
rect 4487 3819 4488 3823
rect 4482 3818 4488 3819
rect 4572 3791 4574 3868
rect 4698 3863 4704 3864
rect 4698 3859 4699 3863
rect 4703 3859 4704 3863
rect 4698 3858 4704 3859
rect 4700 3824 4702 3858
rect 4698 3823 4704 3824
rect 4698 3819 4699 3823
rect 4703 3819 4704 3823
rect 4698 3818 4704 3819
rect 4796 3791 4798 3868
rect 4922 3863 4928 3864
rect 4922 3859 4923 3863
rect 4927 3859 4928 3863
rect 4922 3858 4928 3859
rect 4924 3824 4926 3858
rect 4922 3823 4928 3824
rect 4922 3819 4923 3823
rect 4927 3819 4928 3823
rect 4922 3818 4928 3819
rect 5036 3791 5038 3868
rect 5058 3863 5064 3864
rect 5058 3859 5059 3863
rect 5063 3859 5064 3863
rect 5058 3858 5064 3859
rect 3839 3790 3843 3791
rect 3839 3785 3843 3786
rect 3995 3790 3999 3791
rect 3995 3785 3999 3786
rect 4203 3790 4207 3791
rect 4203 3785 4207 3786
rect 4355 3790 4359 3791
rect 4355 3785 4359 3786
rect 4435 3790 4439 3791
rect 4435 3785 4439 3786
rect 4571 3790 4575 3791
rect 4571 3785 4575 3786
rect 4691 3790 4695 3791
rect 4691 3785 4695 3786
rect 4795 3790 4799 3791
rect 4795 3785 4799 3786
rect 4963 3790 4967 3791
rect 4963 3785 4967 3786
rect 5035 3790 5039 3791
rect 5035 3785 5039 3786
rect 3798 3780 3804 3781
rect 2794 3779 2800 3780
rect 2794 3775 2795 3779
rect 2799 3775 2800 3779
rect 2794 3774 2800 3775
rect 2994 3779 3000 3780
rect 2994 3775 2995 3779
rect 2999 3775 3000 3779
rect 2994 3774 3000 3775
rect 3194 3779 3200 3780
rect 3194 3775 3195 3779
rect 3199 3775 3200 3779
rect 3194 3774 3200 3775
rect 3402 3779 3408 3780
rect 3402 3775 3403 3779
rect 3407 3775 3408 3779
rect 3798 3776 3799 3780
rect 3803 3776 3804 3780
rect 3798 3775 3804 3776
rect 3402 3774 3408 3775
rect 2614 3764 2620 3765
rect 2614 3760 2615 3764
rect 2619 3760 2620 3764
rect 2614 3759 2620 3760
rect 2822 3764 2828 3765
rect 2822 3760 2823 3764
rect 2827 3760 2828 3764
rect 2822 3759 2828 3760
rect 3022 3764 3028 3765
rect 3022 3760 3023 3764
rect 3027 3760 3028 3764
rect 3022 3759 3028 3760
rect 3222 3764 3228 3765
rect 3222 3760 3223 3764
rect 3227 3760 3228 3764
rect 3222 3759 3228 3760
rect 3430 3764 3436 3765
rect 3430 3760 3431 3764
rect 3435 3760 3436 3764
rect 3430 3759 3436 3760
rect 3798 3763 3804 3764
rect 3798 3759 3799 3763
rect 3803 3759 3804 3763
rect 2616 3731 2618 3759
rect 2824 3731 2826 3759
rect 3024 3731 3026 3759
rect 3224 3731 3226 3759
rect 3432 3731 3434 3759
rect 3798 3758 3804 3759
rect 3800 3731 3802 3758
rect 2615 3730 2619 3731
rect 2615 3725 2619 3726
rect 2679 3730 2683 3731
rect 2679 3725 2683 3726
rect 2823 3730 2827 3731
rect 2823 3725 2827 3726
rect 2879 3730 2883 3731
rect 2879 3725 2883 3726
rect 3023 3730 3027 3731
rect 3023 3725 3027 3726
rect 3079 3730 3083 3731
rect 3079 3725 3083 3726
rect 3223 3730 3227 3731
rect 3223 3725 3227 3726
rect 3279 3730 3283 3731
rect 3279 3725 3283 3726
rect 3431 3730 3435 3731
rect 3431 3725 3435 3726
rect 3799 3730 3803 3731
rect 3799 3725 3803 3726
rect 3840 3725 3842 3785
rect 2680 3701 2682 3725
rect 2880 3701 2882 3725
rect 3080 3701 3082 3725
rect 3280 3701 3282 3725
rect 3800 3702 3802 3725
rect 3838 3724 3844 3725
rect 3996 3724 3998 3785
rect 4090 3771 4096 3772
rect 4090 3767 4091 3771
rect 4095 3767 4096 3771
rect 4090 3766 4096 3767
rect 4092 3733 4094 3766
rect 4091 3732 4095 3733
rect 4091 3727 4095 3728
rect 4204 3724 4206 3785
rect 4210 3771 4216 3772
rect 4210 3767 4211 3771
rect 4215 3767 4216 3771
rect 4210 3766 4216 3767
rect 4212 3732 4214 3766
rect 4210 3731 4216 3732
rect 4210 3727 4211 3731
rect 4215 3727 4216 3731
rect 4210 3726 4216 3727
rect 4436 3724 4438 3785
rect 4442 3771 4448 3772
rect 4442 3767 4443 3771
rect 4447 3767 4448 3771
rect 4442 3766 4448 3767
rect 4444 3732 4446 3766
rect 4442 3731 4448 3732
rect 4442 3727 4443 3731
rect 4447 3727 4448 3731
rect 4442 3726 4448 3727
rect 4692 3724 4694 3785
rect 4698 3771 4704 3772
rect 4698 3767 4699 3771
rect 4703 3767 4704 3771
rect 4698 3766 4704 3767
rect 4700 3732 4702 3766
rect 4939 3732 4943 3733
rect 4698 3731 4704 3732
rect 4698 3727 4699 3731
rect 4703 3727 4704 3731
rect 4698 3726 4704 3727
rect 4814 3731 4820 3732
rect 4814 3727 4815 3731
rect 4819 3727 4820 3731
rect 4814 3726 4820 3727
rect 4938 3727 4939 3732
rect 4943 3727 4944 3732
rect 4938 3726 4944 3727
rect 3838 3720 3839 3724
rect 3843 3720 3844 3724
rect 3838 3719 3844 3720
rect 3994 3723 4000 3724
rect 3994 3719 3995 3723
rect 3999 3719 4000 3723
rect 3994 3718 4000 3719
rect 4202 3723 4208 3724
rect 4202 3719 4203 3723
rect 4207 3719 4208 3723
rect 4202 3718 4208 3719
rect 4434 3723 4440 3724
rect 4434 3719 4435 3723
rect 4439 3719 4440 3723
rect 4434 3718 4440 3719
rect 4690 3723 4696 3724
rect 4690 3719 4691 3723
rect 4695 3719 4696 3723
rect 4690 3718 4696 3719
rect 4022 3708 4028 3709
rect 3838 3707 3844 3708
rect 3838 3703 3839 3707
rect 3843 3703 3844 3707
rect 4022 3704 4023 3708
rect 4027 3704 4028 3708
rect 4022 3703 4028 3704
rect 4230 3708 4236 3709
rect 4230 3704 4231 3708
rect 4235 3704 4236 3708
rect 4230 3703 4236 3704
rect 4462 3708 4468 3709
rect 4462 3704 4463 3708
rect 4467 3704 4468 3708
rect 4462 3703 4468 3704
rect 4718 3708 4724 3709
rect 4718 3704 4719 3708
rect 4723 3704 4724 3708
rect 4718 3703 4724 3704
rect 3838 3702 3844 3703
rect 3798 3701 3804 3702
rect 2678 3700 2684 3701
rect 2678 3696 2679 3700
rect 2683 3696 2684 3700
rect 2678 3695 2684 3696
rect 2878 3700 2884 3701
rect 2878 3696 2879 3700
rect 2883 3696 2884 3700
rect 2878 3695 2884 3696
rect 3078 3700 3084 3701
rect 3078 3696 3079 3700
rect 3083 3696 3084 3700
rect 3078 3695 3084 3696
rect 3278 3700 3284 3701
rect 3278 3696 3279 3700
rect 3283 3696 3284 3700
rect 3798 3697 3799 3701
rect 3803 3697 3804 3701
rect 3798 3696 3804 3697
rect 3278 3695 3284 3696
rect 2650 3685 2656 3686
rect 2650 3681 2651 3685
rect 2655 3681 2656 3685
rect 2650 3680 2656 3681
rect 2850 3685 2856 3686
rect 2850 3681 2851 3685
rect 2855 3681 2856 3685
rect 2850 3680 2856 3681
rect 3050 3685 3056 3686
rect 3050 3681 3051 3685
rect 3055 3681 3056 3685
rect 3050 3680 3056 3681
rect 3250 3685 3256 3686
rect 3250 3681 3251 3685
rect 3255 3681 3256 3685
rect 3250 3680 3256 3681
rect 3798 3684 3804 3685
rect 3798 3680 3799 3684
rect 3803 3680 3804 3684
rect 2594 3675 2600 3676
rect 2594 3671 2595 3675
rect 2599 3671 2600 3675
rect 2594 3670 2600 3671
rect 2652 3607 2654 3680
rect 2852 3607 2854 3680
rect 2946 3667 2952 3668
rect 2946 3663 2947 3667
rect 2951 3663 2952 3667
rect 2946 3662 2952 3663
rect 2948 3636 2950 3662
rect 2946 3635 2952 3636
rect 2946 3631 2947 3635
rect 2951 3631 2952 3635
rect 2946 3630 2952 3631
rect 3052 3607 3054 3680
rect 3102 3635 3108 3636
rect 3102 3631 3103 3635
rect 3107 3631 3108 3635
rect 3102 3630 3108 3631
rect 2451 3606 2455 3607
rect 2451 3601 2455 3602
rect 2515 3606 2519 3607
rect 2515 3601 2519 3602
rect 2651 3606 2655 3607
rect 2651 3601 2655 3602
rect 2755 3606 2759 3607
rect 2755 3601 2759 3602
rect 2851 3606 2855 3607
rect 2851 3601 2855 3602
rect 2979 3606 2983 3607
rect 2979 3601 2983 3602
rect 3051 3606 3055 3607
rect 3051 3601 3055 3602
rect 2346 3591 2352 3592
rect 2346 3587 2347 3591
rect 2351 3587 2352 3591
rect 2346 3586 2352 3587
rect 2516 3540 2518 3601
rect 2522 3587 2528 3588
rect 2522 3583 2523 3587
rect 2527 3583 2528 3587
rect 2522 3582 2528 3583
rect 2524 3548 2526 3582
rect 2522 3547 2528 3548
rect 2522 3543 2523 3547
rect 2527 3543 2528 3547
rect 2522 3542 2528 3543
rect 2638 3547 2644 3548
rect 2638 3543 2639 3547
rect 2643 3543 2644 3547
rect 2638 3542 2644 3543
rect 2250 3539 2256 3540
rect 2250 3535 2251 3539
rect 2255 3535 2256 3539
rect 2250 3534 2256 3535
rect 2514 3539 2520 3540
rect 2514 3535 2515 3539
rect 2519 3535 2520 3539
rect 2514 3534 2520 3535
rect 2278 3524 2284 3525
rect 2278 3520 2279 3524
rect 2283 3520 2284 3524
rect 2278 3519 2284 3520
rect 2542 3524 2548 3525
rect 2542 3520 2543 3524
rect 2547 3520 2548 3524
rect 2542 3519 2548 3520
rect 2280 3487 2282 3519
rect 2544 3487 2546 3519
rect 2191 3486 2195 3487
rect 2191 3481 2195 3482
rect 2279 3486 2283 3487
rect 2279 3481 2283 3482
rect 2399 3486 2403 3487
rect 2399 3481 2403 3482
rect 2543 3486 2547 3487
rect 2543 3481 2547 3482
rect 2615 3486 2619 3487
rect 2615 3481 2619 3482
rect 2192 3457 2194 3481
rect 2400 3457 2402 3481
rect 2616 3457 2618 3481
rect 2190 3456 2196 3457
rect 2190 3452 2191 3456
rect 2195 3452 2196 3456
rect 2190 3451 2196 3452
rect 2398 3456 2404 3457
rect 2398 3452 2399 3456
rect 2403 3452 2404 3456
rect 2398 3451 2404 3452
rect 2614 3456 2620 3457
rect 2614 3452 2615 3456
rect 2619 3452 2620 3456
rect 2614 3451 2620 3452
rect 2162 3441 2168 3442
rect 2162 3437 2163 3441
rect 2167 3437 2168 3441
rect 2162 3436 2168 3437
rect 2370 3441 2376 3442
rect 2370 3437 2371 3441
rect 2375 3437 2376 3441
rect 2370 3436 2376 3437
rect 2586 3441 2592 3442
rect 2586 3437 2587 3441
rect 2591 3437 2592 3441
rect 2586 3436 2592 3437
rect 2122 3431 2128 3432
rect 2122 3427 2123 3431
rect 2127 3427 2128 3431
rect 2122 3426 2128 3427
rect 2124 3392 2126 3426
rect 2090 3391 2096 3392
rect 2090 3387 2091 3391
rect 2095 3387 2096 3391
rect 2090 3386 2096 3387
rect 2122 3391 2128 3392
rect 2122 3387 2123 3391
rect 2127 3387 2128 3391
rect 2122 3386 2128 3387
rect 2164 3335 2166 3436
rect 2334 3431 2340 3432
rect 2334 3427 2335 3431
rect 2339 3427 2340 3431
rect 2334 3426 2340 3427
rect 2346 3431 2352 3432
rect 2346 3427 2347 3431
rect 2351 3427 2352 3431
rect 2346 3426 2352 3427
rect 2336 3392 2338 3426
rect 2334 3391 2340 3392
rect 2334 3387 2335 3391
rect 2339 3387 2340 3391
rect 2334 3386 2340 3387
rect 1975 3334 1979 3335
rect 1975 3329 1979 3330
rect 1995 3334 1999 3335
rect 1995 3329 1999 3330
rect 2163 3334 2167 3335
rect 2163 3329 2167 3330
rect 2195 3334 2199 3335
rect 2195 3329 2199 3330
rect 1934 3296 1940 3297
rect 1934 3292 1935 3296
rect 1939 3292 1940 3296
rect 1934 3291 1940 3292
rect 1934 3279 1940 3280
rect 1934 3275 1935 3279
rect 1939 3275 1940 3279
rect 1934 3274 1940 3275
rect 1950 3275 1956 3276
rect 1936 3251 1938 3274
rect 1950 3271 1951 3275
rect 1955 3271 1956 3275
rect 1950 3270 1956 3271
rect 1471 3250 1475 3251
rect 1471 3245 1475 3246
rect 1655 3250 1659 3251
rect 1655 3245 1659 3246
rect 1815 3250 1819 3251
rect 1815 3245 1819 3246
rect 1935 3250 1939 3251
rect 1935 3245 1939 3246
rect 1472 3221 1474 3245
rect 1656 3221 1658 3245
rect 1816 3221 1818 3245
rect 1936 3222 1938 3245
rect 1934 3221 1940 3222
rect 1470 3220 1476 3221
rect 1470 3216 1471 3220
rect 1475 3216 1476 3220
rect 1470 3215 1476 3216
rect 1654 3220 1660 3221
rect 1654 3216 1655 3220
rect 1659 3216 1660 3220
rect 1654 3215 1660 3216
rect 1814 3220 1820 3221
rect 1814 3216 1815 3220
rect 1819 3216 1820 3220
rect 1934 3217 1935 3221
rect 1939 3217 1940 3221
rect 1934 3216 1940 3217
rect 1814 3215 1820 3216
rect 1442 3205 1448 3206
rect 1442 3201 1443 3205
rect 1447 3201 1448 3205
rect 1442 3200 1448 3201
rect 1626 3205 1632 3206
rect 1626 3201 1627 3205
rect 1631 3201 1632 3205
rect 1626 3200 1632 3201
rect 1786 3205 1792 3206
rect 1786 3201 1787 3205
rect 1791 3201 1792 3205
rect 1786 3200 1792 3201
rect 1934 3204 1940 3205
rect 1934 3200 1935 3204
rect 1939 3200 1940 3204
rect 1390 3195 1396 3196
rect 1390 3191 1391 3195
rect 1395 3191 1396 3195
rect 1390 3190 1396 3191
rect 1398 3147 1404 3148
rect 1398 3143 1399 3147
rect 1403 3143 1404 3147
rect 1398 3142 1404 3143
rect 699 3130 703 3131
rect 699 3125 703 3126
rect 835 3130 839 3131
rect 835 3125 839 3126
rect 891 3130 895 3131
rect 891 3125 895 3126
rect 971 3130 975 3131
rect 971 3125 975 3126
rect 1083 3130 1087 3131
rect 1083 3125 1087 3126
rect 1107 3130 1111 3131
rect 1107 3125 1111 3126
rect 1243 3130 1247 3131
rect 1243 3125 1247 3126
rect 1267 3130 1271 3131
rect 1267 3125 1271 3126
rect 1379 3130 1383 3131
rect 1379 3125 1383 3126
rect 658 3115 664 3116
rect 658 3111 659 3115
rect 663 3111 664 3115
rect 658 3110 664 3111
rect 700 3064 702 3125
rect 706 3111 712 3112
rect 706 3107 707 3111
rect 711 3107 712 3111
rect 706 3106 712 3107
rect 708 3072 710 3106
rect 706 3071 712 3072
rect 706 3067 707 3071
rect 711 3067 712 3071
rect 706 3066 712 3067
rect 836 3064 838 3125
rect 842 3111 848 3112
rect 842 3107 843 3111
rect 847 3107 848 3111
rect 842 3106 848 3107
rect 844 3072 846 3106
rect 842 3071 848 3072
rect 842 3067 843 3071
rect 847 3067 848 3071
rect 842 3066 848 3067
rect 972 3064 974 3125
rect 978 3111 984 3112
rect 978 3107 979 3111
rect 983 3107 984 3111
rect 978 3106 984 3107
rect 980 3072 982 3106
rect 978 3071 984 3072
rect 978 3067 979 3071
rect 983 3067 984 3071
rect 978 3066 984 3067
rect 1108 3064 1110 3125
rect 1114 3111 1120 3112
rect 1114 3107 1115 3111
rect 1119 3107 1120 3111
rect 1114 3106 1120 3107
rect 1116 3072 1118 3106
rect 1114 3071 1120 3072
rect 1114 3067 1115 3071
rect 1119 3067 1120 3071
rect 1114 3066 1120 3067
rect 1244 3064 1246 3125
rect 1250 3111 1256 3112
rect 1250 3107 1251 3111
rect 1255 3107 1256 3111
rect 1250 3106 1256 3107
rect 1252 3072 1254 3106
rect 1250 3071 1256 3072
rect 1250 3067 1251 3071
rect 1255 3067 1256 3071
rect 1250 3066 1256 3067
rect 1380 3064 1382 3125
rect 1386 3111 1392 3112
rect 1386 3107 1387 3111
rect 1391 3107 1392 3111
rect 1386 3106 1392 3107
rect 1388 3072 1390 3106
rect 1400 3072 1402 3142
rect 1444 3131 1446 3200
rect 1566 3195 1572 3196
rect 1566 3191 1567 3195
rect 1571 3191 1572 3195
rect 1566 3190 1572 3191
rect 1594 3195 1600 3196
rect 1594 3191 1595 3195
rect 1599 3191 1600 3195
rect 1594 3190 1600 3191
rect 1443 3130 1447 3131
rect 1443 3125 1447 3126
rect 1515 3130 1519 3131
rect 1515 3125 1519 3126
rect 1386 3071 1392 3072
rect 1386 3067 1387 3071
rect 1391 3067 1392 3071
rect 1386 3066 1392 3067
rect 1398 3071 1404 3072
rect 1398 3067 1399 3071
rect 1403 3067 1404 3071
rect 1398 3066 1404 3067
rect 1516 3064 1518 3125
rect 1568 3116 1570 3190
rect 1596 3156 1598 3190
rect 1594 3155 1600 3156
rect 1594 3151 1595 3155
rect 1599 3151 1600 3155
rect 1594 3150 1600 3151
rect 1628 3131 1630 3200
rect 1788 3131 1790 3200
rect 1934 3199 1940 3200
rect 1936 3131 1938 3199
rect 1952 3156 1954 3270
rect 1976 3269 1978 3329
rect 1974 3268 1980 3269
rect 1996 3268 1998 3329
rect 2186 3319 2192 3320
rect 2186 3315 2187 3319
rect 2191 3315 2192 3319
rect 2186 3314 2192 3315
rect 2188 3276 2190 3314
rect 2186 3275 2192 3276
rect 2186 3271 2187 3275
rect 2191 3271 2192 3275
rect 2186 3270 2192 3271
rect 2196 3268 2198 3329
rect 2348 3320 2350 3426
rect 2372 3335 2374 3436
rect 2588 3335 2590 3436
rect 2640 3392 2642 3542
rect 2756 3540 2758 3601
rect 2850 3587 2856 3588
rect 2850 3583 2851 3587
rect 2855 3583 2856 3587
rect 2850 3582 2856 3583
rect 2852 3556 2854 3582
rect 2850 3555 2856 3556
rect 2850 3551 2851 3555
rect 2855 3551 2856 3555
rect 2850 3550 2856 3551
rect 2980 3540 2982 3601
rect 2986 3587 2992 3588
rect 2986 3583 2987 3587
rect 2991 3583 2992 3587
rect 2986 3582 2992 3583
rect 2988 3548 2990 3582
rect 3104 3548 3106 3630
rect 3252 3607 3254 3680
rect 3798 3679 3804 3680
rect 3800 3607 3802 3679
rect 3840 3651 3842 3702
rect 4024 3651 4026 3703
rect 4232 3651 4234 3703
rect 4464 3651 4466 3703
rect 4720 3651 4722 3703
rect 3839 3650 3843 3651
rect 3839 3645 3843 3646
rect 4023 3650 4027 3651
rect 4023 3645 4027 3646
rect 4215 3650 4219 3651
rect 4215 3645 4219 3646
rect 4231 3650 4235 3651
rect 4231 3645 4235 3646
rect 4399 3650 4403 3651
rect 4399 3645 4403 3646
rect 4463 3650 4467 3651
rect 4463 3645 4467 3646
rect 4607 3650 4611 3651
rect 4607 3645 4611 3646
rect 4719 3650 4723 3651
rect 4719 3645 4723 3646
rect 3840 3622 3842 3645
rect 3838 3621 3844 3622
rect 4216 3621 4218 3645
rect 4400 3621 4402 3645
rect 4608 3621 4610 3645
rect 3838 3617 3839 3621
rect 3843 3617 3844 3621
rect 3838 3616 3844 3617
rect 4214 3620 4220 3621
rect 4214 3616 4215 3620
rect 4219 3616 4220 3620
rect 4214 3615 4220 3616
rect 4398 3620 4404 3621
rect 4398 3616 4399 3620
rect 4403 3616 4404 3620
rect 4398 3615 4404 3616
rect 4606 3620 4612 3621
rect 4606 3616 4607 3620
rect 4611 3616 4612 3620
rect 4606 3615 4612 3616
rect 3195 3606 3199 3607
rect 3195 3601 3199 3602
rect 3251 3606 3255 3607
rect 3251 3601 3255 3602
rect 3411 3606 3415 3607
rect 3411 3601 3415 3602
rect 3627 3606 3631 3607
rect 3627 3601 3631 3602
rect 3799 3606 3803 3607
rect 4186 3605 4192 3606
rect 3799 3601 3803 3602
rect 3838 3604 3844 3605
rect 2986 3547 2992 3548
rect 2986 3543 2987 3547
rect 2991 3543 2992 3547
rect 2986 3542 2992 3543
rect 3102 3547 3108 3548
rect 3102 3543 3103 3547
rect 3107 3543 3108 3547
rect 3102 3542 3108 3543
rect 3196 3540 3198 3601
rect 3412 3540 3414 3601
rect 3628 3540 3630 3601
rect 3634 3587 3640 3588
rect 3634 3583 3635 3587
rect 3639 3583 3640 3587
rect 3634 3582 3640 3583
rect 2754 3539 2760 3540
rect 2754 3535 2755 3539
rect 2759 3535 2760 3539
rect 2754 3534 2760 3535
rect 2978 3539 2984 3540
rect 2978 3535 2979 3539
rect 2983 3535 2984 3539
rect 2978 3534 2984 3535
rect 3194 3539 3200 3540
rect 3194 3535 3195 3539
rect 3199 3535 3200 3539
rect 3194 3534 3200 3535
rect 3410 3539 3416 3540
rect 3410 3535 3411 3539
rect 3415 3535 3416 3539
rect 3410 3534 3416 3535
rect 3626 3539 3632 3540
rect 3626 3535 3627 3539
rect 3631 3535 3632 3539
rect 3626 3534 3632 3535
rect 2782 3524 2788 3525
rect 2782 3520 2783 3524
rect 2787 3520 2788 3524
rect 2782 3519 2788 3520
rect 3006 3524 3012 3525
rect 3006 3520 3007 3524
rect 3011 3520 3012 3524
rect 3006 3519 3012 3520
rect 3222 3524 3228 3525
rect 3222 3520 3223 3524
rect 3227 3520 3228 3524
rect 3222 3519 3228 3520
rect 3438 3524 3444 3525
rect 3438 3520 3439 3524
rect 3443 3520 3444 3524
rect 3438 3519 3444 3520
rect 2784 3487 2786 3519
rect 3008 3487 3010 3519
rect 3224 3487 3226 3519
rect 3440 3487 3442 3519
rect 2783 3486 2787 3487
rect 2783 3481 2787 3482
rect 2831 3486 2835 3487
rect 2831 3481 2835 3482
rect 3007 3486 3011 3487
rect 3007 3481 3011 3482
rect 3047 3486 3051 3487
rect 3047 3481 3051 3482
rect 3223 3486 3227 3487
rect 3223 3481 3227 3482
rect 3263 3486 3267 3487
rect 3263 3481 3267 3482
rect 3439 3486 3443 3487
rect 3439 3481 3443 3482
rect 3479 3486 3483 3487
rect 3479 3481 3483 3482
rect 2832 3457 2834 3481
rect 3048 3457 3050 3481
rect 3264 3457 3266 3481
rect 3480 3457 3482 3481
rect 2830 3456 2836 3457
rect 2830 3452 2831 3456
rect 2835 3452 2836 3456
rect 2830 3451 2836 3452
rect 3046 3456 3052 3457
rect 3046 3452 3047 3456
rect 3051 3452 3052 3456
rect 3046 3451 3052 3452
rect 3262 3456 3268 3457
rect 3262 3452 3263 3456
rect 3267 3452 3268 3456
rect 3262 3451 3268 3452
rect 3478 3456 3484 3457
rect 3478 3452 3479 3456
rect 3483 3452 3484 3456
rect 3478 3451 3484 3452
rect 2802 3441 2808 3442
rect 2802 3437 2803 3441
rect 2807 3437 2808 3441
rect 2802 3436 2808 3437
rect 3018 3441 3024 3442
rect 3018 3437 3019 3441
rect 3023 3437 3024 3441
rect 3018 3436 3024 3437
rect 3234 3441 3240 3442
rect 3234 3437 3235 3441
rect 3239 3437 3240 3441
rect 3234 3436 3240 3437
rect 3450 3441 3456 3442
rect 3450 3437 3451 3441
rect 3455 3437 3456 3441
rect 3450 3436 3456 3437
rect 2638 3391 2644 3392
rect 2638 3387 2639 3391
rect 2643 3387 2644 3391
rect 2638 3386 2644 3387
rect 2804 3335 2806 3436
rect 3020 3335 3022 3436
rect 3146 3431 3152 3432
rect 3146 3427 3147 3431
rect 3151 3427 3152 3431
rect 3146 3426 3152 3427
rect 3148 3392 3150 3426
rect 3146 3391 3152 3392
rect 3146 3387 3147 3391
rect 3151 3387 3152 3391
rect 3146 3386 3152 3387
rect 3236 3335 3238 3436
rect 3362 3431 3368 3432
rect 3362 3427 3363 3431
rect 3367 3427 3368 3431
rect 3362 3426 3368 3427
rect 3364 3392 3366 3426
rect 3362 3391 3368 3392
rect 3362 3387 3363 3391
rect 3367 3387 3368 3391
rect 3362 3386 3368 3387
rect 3452 3335 3454 3436
rect 3636 3432 3638 3582
rect 3800 3541 3802 3601
rect 3838 3600 3839 3604
rect 3843 3600 3844 3604
rect 4186 3601 4187 3605
rect 4191 3601 4192 3605
rect 4186 3600 4192 3601
rect 4370 3605 4376 3606
rect 4370 3601 4371 3605
rect 4375 3601 4376 3605
rect 4370 3600 4376 3601
rect 4578 3605 4584 3606
rect 4578 3601 4579 3605
rect 4583 3601 4584 3605
rect 4578 3600 4584 3601
rect 4802 3605 4808 3606
rect 4802 3601 4803 3605
rect 4807 3601 4808 3605
rect 4802 3600 4808 3601
rect 3838 3599 3844 3600
rect 3798 3540 3804 3541
rect 3798 3536 3799 3540
rect 3803 3536 3804 3540
rect 3798 3535 3804 3536
rect 3654 3524 3660 3525
rect 3654 3520 3655 3524
rect 3659 3520 3660 3524
rect 3654 3519 3660 3520
rect 3798 3523 3804 3524
rect 3798 3519 3799 3523
rect 3803 3519 3804 3523
rect 3656 3487 3658 3519
rect 3798 3518 3804 3519
rect 3800 3487 3802 3518
rect 3840 3515 3842 3599
rect 4188 3515 4190 3600
rect 4326 3595 4332 3596
rect 4326 3591 4327 3595
rect 4331 3591 4332 3595
rect 4326 3590 4332 3591
rect 4328 3556 4330 3590
rect 4326 3555 4332 3556
rect 4326 3551 4327 3555
rect 4331 3551 4332 3555
rect 4326 3550 4332 3551
rect 4372 3515 4374 3600
rect 4538 3595 4544 3596
rect 4538 3591 4539 3595
rect 4543 3591 4544 3595
rect 4538 3590 4544 3591
rect 4540 3556 4542 3590
rect 4538 3555 4544 3556
rect 4538 3551 4539 3555
rect 4543 3551 4544 3555
rect 4538 3550 4544 3551
rect 4580 3515 4582 3600
rect 4706 3595 4712 3596
rect 4706 3591 4707 3595
rect 4711 3591 4712 3595
rect 4706 3590 4712 3591
rect 4626 3587 4632 3588
rect 4626 3583 4627 3587
rect 4631 3583 4632 3587
rect 4626 3582 4632 3583
rect 3839 3514 3843 3515
rect 3839 3509 3843 3510
rect 4187 3514 4191 3515
rect 4187 3509 4191 3510
rect 4371 3514 4375 3515
rect 4371 3509 4375 3510
rect 4531 3514 4535 3515
rect 4531 3509 4535 3510
rect 4579 3514 4583 3515
rect 4579 3509 4583 3510
rect 3655 3486 3659 3487
rect 3655 3481 3659 3482
rect 3679 3486 3683 3487
rect 3679 3481 3683 3482
rect 3799 3486 3803 3487
rect 3799 3481 3803 3482
rect 3680 3457 3682 3481
rect 3800 3458 3802 3481
rect 3798 3457 3804 3458
rect 3678 3456 3684 3457
rect 3678 3452 3679 3456
rect 3683 3452 3684 3456
rect 3798 3453 3799 3457
rect 3803 3453 3804 3457
rect 3798 3452 3804 3453
rect 3678 3451 3684 3452
rect 3840 3449 3842 3509
rect 3838 3448 3844 3449
rect 4532 3448 4534 3509
rect 4628 3500 4630 3582
rect 4708 3556 4710 3590
rect 4706 3555 4712 3556
rect 4706 3551 4707 3555
rect 4711 3551 4712 3555
rect 4706 3550 4712 3551
rect 4804 3515 4806 3600
rect 4816 3548 4818 3726
rect 4964 3724 4966 3785
rect 5060 3776 5062 3858
rect 5284 3791 5286 3868
rect 5400 3864 5402 4034
rect 5516 3988 5518 4049
rect 5620 4040 5622 4106
rect 5664 4055 5666 4115
rect 5663 4054 5667 4055
rect 5663 4049 5667 4050
rect 5618 4039 5624 4040
rect 5618 4035 5619 4039
rect 5623 4035 5624 4039
rect 5618 4034 5624 4035
rect 5634 3995 5640 3996
rect 5634 3991 5635 3995
rect 5639 3991 5640 3995
rect 5634 3990 5640 3991
rect 5514 3987 5520 3988
rect 5514 3983 5515 3987
rect 5519 3983 5520 3987
rect 5514 3982 5520 3983
rect 5406 3972 5412 3973
rect 5406 3968 5407 3972
rect 5411 3968 5412 3972
rect 5406 3967 5412 3968
rect 5542 3972 5548 3973
rect 5542 3968 5543 3972
rect 5547 3968 5548 3972
rect 5542 3967 5548 3968
rect 5408 3919 5410 3967
rect 5544 3919 5546 3967
rect 5407 3918 5411 3919
rect 5407 3913 5411 3914
rect 5543 3918 5547 3919
rect 5543 3913 5547 3914
rect 5544 3889 5546 3913
rect 5542 3888 5548 3889
rect 5542 3884 5543 3888
rect 5547 3884 5548 3888
rect 5542 3883 5548 3884
rect 5514 3873 5520 3874
rect 5514 3869 5515 3873
rect 5519 3869 5520 3873
rect 5514 3868 5520 3869
rect 5398 3863 5404 3864
rect 5398 3859 5399 3863
rect 5403 3859 5404 3863
rect 5398 3858 5404 3859
rect 5374 3823 5380 3824
rect 5374 3819 5375 3823
rect 5379 3819 5380 3823
rect 5374 3818 5380 3819
rect 5251 3790 5255 3791
rect 5251 3785 5255 3786
rect 5283 3790 5287 3791
rect 5283 3785 5287 3786
rect 5058 3775 5064 3776
rect 5058 3771 5059 3775
rect 5063 3771 5064 3775
rect 5058 3770 5064 3771
rect 5252 3724 5254 3785
rect 5346 3771 5352 3772
rect 5346 3767 5347 3771
rect 5351 3767 5352 3771
rect 5346 3766 5352 3767
rect 4962 3723 4968 3724
rect 4962 3719 4963 3723
rect 4967 3719 4968 3723
rect 4962 3718 4968 3719
rect 5250 3723 5256 3724
rect 5250 3719 5251 3723
rect 5255 3719 5256 3723
rect 5250 3718 5256 3719
rect 4990 3708 4996 3709
rect 4990 3704 4991 3708
rect 4995 3704 4996 3708
rect 4990 3703 4996 3704
rect 5278 3708 5284 3709
rect 5278 3704 5279 3708
rect 5283 3704 5284 3708
rect 5278 3703 5284 3704
rect 4992 3651 4994 3703
rect 5280 3651 5282 3703
rect 4831 3650 4835 3651
rect 4831 3645 4835 3646
rect 4991 3650 4995 3651
rect 4991 3645 4995 3646
rect 5071 3650 5075 3651
rect 5071 3645 5075 3646
rect 5279 3650 5283 3651
rect 5279 3645 5283 3646
rect 5319 3650 5323 3651
rect 5319 3645 5323 3646
rect 4832 3621 4834 3645
rect 5072 3621 5074 3645
rect 5320 3621 5322 3645
rect 4830 3620 4836 3621
rect 4830 3616 4831 3620
rect 4835 3616 4836 3620
rect 4830 3615 4836 3616
rect 5070 3620 5076 3621
rect 5070 3616 5071 3620
rect 5075 3616 5076 3620
rect 5070 3615 5076 3616
rect 5318 3620 5324 3621
rect 5318 3616 5319 3620
rect 5323 3616 5324 3620
rect 5318 3615 5324 3616
rect 5042 3605 5048 3606
rect 5042 3601 5043 3605
rect 5047 3601 5048 3605
rect 5042 3600 5048 3601
rect 5290 3605 5296 3606
rect 5290 3601 5291 3605
rect 5295 3601 5296 3605
rect 5290 3600 5296 3601
rect 4930 3595 4936 3596
rect 4930 3591 4931 3595
rect 4935 3591 4936 3595
rect 4930 3590 4936 3591
rect 4932 3556 4934 3590
rect 4930 3555 4936 3556
rect 4930 3551 4931 3555
rect 4935 3551 4936 3555
rect 4930 3550 4936 3551
rect 4814 3547 4820 3548
rect 4814 3543 4815 3547
rect 4819 3543 4820 3547
rect 4814 3542 4820 3543
rect 5044 3515 5046 3600
rect 5292 3515 5294 3600
rect 5348 3596 5350 3766
rect 5376 3732 5378 3818
rect 5516 3791 5518 3868
rect 5610 3863 5616 3864
rect 5610 3859 5611 3863
rect 5615 3859 5616 3863
rect 5610 3858 5616 3859
rect 5515 3790 5519 3791
rect 5515 3785 5519 3786
rect 5374 3731 5380 3732
rect 5374 3727 5375 3731
rect 5379 3727 5380 3731
rect 5374 3726 5380 3727
rect 5516 3724 5518 3785
rect 5612 3776 5614 3858
rect 5636 3824 5638 3990
rect 5664 3989 5666 4049
rect 5662 3988 5668 3989
rect 5662 3984 5663 3988
rect 5667 3984 5668 3988
rect 5662 3983 5668 3984
rect 5662 3971 5668 3972
rect 5662 3967 5663 3971
rect 5667 3967 5668 3971
rect 5662 3966 5668 3967
rect 5664 3919 5666 3966
rect 5663 3918 5667 3919
rect 5663 3913 5667 3914
rect 5664 3890 5666 3913
rect 5662 3889 5668 3890
rect 5662 3885 5663 3889
rect 5667 3885 5668 3889
rect 5662 3884 5668 3885
rect 5662 3872 5668 3873
rect 5662 3868 5663 3872
rect 5667 3868 5668 3872
rect 5662 3867 5668 3868
rect 5634 3823 5640 3824
rect 5634 3819 5635 3823
rect 5639 3819 5640 3823
rect 5634 3818 5640 3819
rect 5664 3791 5666 3867
rect 5663 3790 5667 3791
rect 5663 3785 5667 3786
rect 5610 3775 5616 3776
rect 5610 3771 5611 3775
rect 5615 3771 5616 3775
rect 5610 3770 5616 3771
rect 5626 3731 5632 3732
rect 5626 3727 5627 3731
rect 5631 3727 5632 3731
rect 5626 3726 5632 3727
rect 5514 3723 5520 3724
rect 5514 3719 5515 3723
rect 5519 3719 5520 3723
rect 5514 3718 5520 3719
rect 5542 3708 5548 3709
rect 5542 3704 5543 3708
rect 5547 3704 5548 3708
rect 5542 3703 5548 3704
rect 5544 3651 5546 3703
rect 5543 3650 5547 3651
rect 5543 3645 5547 3646
rect 5544 3621 5546 3645
rect 5542 3620 5548 3621
rect 5542 3616 5543 3620
rect 5547 3616 5548 3620
rect 5542 3615 5548 3616
rect 5514 3605 5520 3606
rect 5514 3601 5515 3605
rect 5519 3601 5520 3605
rect 5514 3600 5520 3601
rect 5346 3595 5352 3596
rect 5346 3591 5347 3595
rect 5351 3591 5352 3595
rect 5346 3590 5352 3591
rect 5386 3555 5392 3556
rect 5386 3551 5387 3555
rect 5391 3551 5392 3555
rect 5386 3550 5392 3551
rect 4683 3514 4687 3515
rect 4683 3509 4687 3510
rect 4803 3514 4807 3515
rect 4803 3509 4807 3510
rect 4843 3514 4847 3515
rect 4843 3509 4847 3510
rect 5003 3514 5007 3515
rect 5003 3509 5007 3510
rect 5043 3514 5047 3515
rect 5043 3509 5047 3510
rect 5171 3514 5175 3515
rect 5171 3509 5175 3510
rect 5291 3514 5295 3515
rect 5291 3509 5295 3510
rect 5347 3514 5351 3515
rect 5347 3509 5351 3510
rect 4626 3499 4632 3500
rect 4626 3495 4627 3499
rect 4631 3495 4632 3499
rect 4626 3494 4632 3495
rect 4684 3448 4686 3509
rect 4690 3495 4696 3496
rect 4690 3491 4691 3495
rect 4695 3491 4696 3495
rect 4690 3490 4696 3491
rect 4692 3456 4694 3490
rect 4690 3455 4696 3456
rect 4690 3451 4691 3455
rect 4695 3451 4696 3455
rect 4690 3450 4696 3451
rect 4844 3448 4846 3509
rect 4850 3495 4856 3496
rect 4850 3491 4851 3495
rect 4855 3491 4856 3495
rect 4850 3490 4856 3491
rect 4852 3456 4854 3490
rect 4850 3455 4856 3456
rect 4850 3451 4851 3455
rect 4855 3451 4856 3455
rect 4850 3450 4856 3451
rect 5004 3448 5006 3509
rect 5010 3495 5016 3496
rect 5010 3491 5011 3495
rect 5015 3491 5016 3495
rect 5010 3490 5016 3491
rect 5012 3456 5014 3490
rect 5010 3455 5016 3456
rect 5010 3451 5011 3455
rect 5015 3451 5016 3455
rect 5010 3450 5016 3451
rect 5172 3448 5174 3509
rect 5318 3499 5324 3500
rect 5178 3495 5184 3496
rect 5178 3491 5179 3495
rect 5183 3491 5184 3495
rect 5318 3495 5319 3499
rect 5323 3495 5324 3499
rect 5318 3494 5324 3495
rect 5178 3490 5184 3491
rect 5180 3456 5182 3490
rect 5178 3455 5184 3456
rect 5178 3451 5179 3455
rect 5183 3451 5184 3455
rect 5178 3450 5184 3451
rect 5238 3455 5244 3456
rect 5238 3451 5239 3455
rect 5243 3451 5244 3455
rect 5238 3450 5244 3451
rect 3838 3444 3839 3448
rect 3843 3444 3844 3448
rect 3838 3443 3844 3444
rect 4530 3447 4536 3448
rect 4530 3443 4531 3447
rect 4535 3443 4536 3447
rect 4530 3442 4536 3443
rect 4682 3447 4688 3448
rect 4682 3443 4683 3447
rect 4687 3443 4688 3447
rect 4682 3442 4688 3443
rect 4842 3447 4848 3448
rect 4842 3443 4843 3447
rect 4847 3443 4848 3447
rect 4842 3442 4848 3443
rect 5002 3447 5008 3448
rect 5002 3443 5003 3447
rect 5007 3443 5008 3447
rect 5002 3442 5008 3443
rect 5170 3447 5176 3448
rect 5170 3443 5171 3447
rect 5175 3443 5176 3447
rect 5170 3442 5176 3443
rect 3650 3441 3656 3442
rect 3650 3437 3651 3441
rect 3655 3437 3656 3441
rect 3650 3436 3656 3437
rect 3798 3440 3804 3441
rect 3798 3436 3799 3440
rect 3803 3436 3804 3440
rect 3634 3431 3640 3432
rect 3634 3427 3635 3431
rect 3639 3427 3640 3431
rect 3634 3426 3640 3427
rect 3652 3335 3654 3436
rect 3798 3435 3804 3436
rect 3690 3431 3696 3432
rect 3690 3427 3691 3431
rect 3695 3427 3696 3431
rect 3690 3426 3696 3427
rect 3692 3376 3694 3426
rect 3746 3391 3752 3392
rect 3746 3387 3747 3391
rect 3751 3387 3752 3391
rect 3746 3386 3752 3387
rect 3690 3375 3696 3376
rect 3690 3371 3691 3375
rect 3695 3371 3696 3375
rect 3690 3370 3696 3371
rect 3748 3344 3750 3386
rect 3746 3343 3752 3344
rect 3746 3339 3747 3343
rect 3751 3339 3752 3343
rect 3746 3338 3752 3339
rect 3800 3335 3802 3435
rect 4558 3432 4564 3433
rect 3838 3431 3844 3432
rect 3838 3427 3839 3431
rect 3843 3427 3844 3431
rect 4558 3428 4559 3432
rect 4563 3428 4564 3432
rect 4558 3427 4564 3428
rect 4710 3432 4716 3433
rect 4710 3428 4711 3432
rect 4715 3428 4716 3432
rect 4710 3427 4716 3428
rect 4870 3432 4876 3433
rect 4870 3428 4871 3432
rect 4875 3428 4876 3432
rect 4870 3427 4876 3428
rect 5030 3432 5036 3433
rect 5030 3428 5031 3432
rect 5035 3428 5036 3432
rect 5030 3427 5036 3428
rect 5198 3432 5204 3433
rect 5198 3428 5199 3432
rect 5203 3428 5204 3432
rect 5198 3427 5204 3428
rect 3838 3426 3844 3427
rect 3840 3399 3842 3426
rect 4560 3399 4562 3427
rect 4712 3399 4714 3427
rect 4872 3399 4874 3427
rect 5032 3399 5034 3427
rect 5200 3399 5202 3427
rect 3839 3398 3843 3399
rect 3839 3393 3843 3394
rect 3887 3398 3891 3399
rect 3887 3393 3891 3394
rect 4151 3398 4155 3399
rect 4151 3393 4155 3394
rect 4423 3398 4427 3399
rect 4423 3393 4427 3394
rect 4559 3398 4563 3399
rect 4559 3393 4563 3394
rect 4671 3398 4675 3399
rect 4671 3393 4675 3394
rect 4711 3398 4715 3399
rect 4711 3393 4715 3394
rect 4871 3398 4875 3399
rect 4871 3393 4875 3394
rect 4895 3398 4899 3399
rect 4895 3393 4899 3394
rect 5031 3398 5035 3399
rect 5031 3393 5035 3394
rect 5111 3398 5115 3399
rect 5111 3393 5115 3394
rect 5199 3398 5203 3399
rect 5199 3393 5203 3394
rect 3840 3370 3842 3393
rect 3838 3369 3844 3370
rect 3888 3369 3890 3393
rect 4152 3369 4154 3393
rect 4424 3369 4426 3393
rect 4672 3369 4674 3393
rect 4896 3369 4898 3393
rect 5112 3369 5114 3393
rect 3838 3365 3839 3369
rect 3843 3365 3844 3369
rect 3838 3364 3844 3365
rect 3886 3368 3892 3369
rect 3886 3364 3887 3368
rect 3891 3364 3892 3368
rect 3886 3363 3892 3364
rect 4150 3368 4156 3369
rect 4150 3364 4151 3368
rect 4155 3364 4156 3368
rect 4150 3363 4156 3364
rect 4422 3368 4428 3369
rect 4422 3364 4423 3368
rect 4427 3364 4428 3368
rect 4422 3363 4428 3364
rect 4670 3368 4676 3369
rect 4670 3364 4671 3368
rect 4675 3364 4676 3368
rect 4670 3363 4676 3364
rect 4894 3368 4900 3369
rect 4894 3364 4895 3368
rect 4899 3364 4900 3368
rect 4894 3363 4900 3364
rect 5110 3368 5116 3369
rect 5110 3364 5111 3368
rect 5115 3364 5116 3368
rect 5110 3363 5116 3364
rect 3858 3353 3864 3354
rect 3838 3352 3844 3353
rect 3838 3348 3839 3352
rect 3843 3348 3844 3352
rect 3858 3349 3859 3353
rect 3863 3349 3864 3353
rect 3858 3348 3864 3349
rect 4122 3353 4128 3354
rect 4122 3349 4123 3353
rect 4127 3349 4128 3353
rect 4122 3348 4128 3349
rect 4394 3353 4400 3354
rect 4394 3349 4395 3353
rect 4399 3349 4400 3353
rect 4394 3348 4400 3349
rect 4642 3353 4648 3354
rect 4642 3349 4643 3353
rect 4647 3349 4648 3353
rect 4642 3348 4648 3349
rect 4866 3353 4872 3354
rect 4866 3349 4867 3353
rect 4871 3349 4872 3353
rect 4866 3348 4872 3349
rect 5082 3353 5088 3354
rect 5082 3349 5083 3353
rect 5087 3349 5088 3353
rect 5082 3348 5088 3349
rect 3838 3347 3844 3348
rect 2371 3334 2375 3335
rect 2371 3329 2375 3330
rect 2411 3334 2415 3335
rect 2411 3329 2415 3330
rect 2587 3334 2591 3335
rect 2587 3329 2591 3330
rect 2619 3334 2623 3335
rect 2619 3329 2623 3330
rect 2803 3334 2807 3335
rect 2803 3329 2807 3330
rect 2811 3334 2815 3335
rect 2811 3329 2815 3330
rect 3003 3334 3007 3335
rect 3003 3329 3007 3330
rect 3019 3334 3023 3335
rect 3019 3329 3023 3330
rect 3187 3334 3191 3335
rect 3187 3329 3191 3330
rect 3235 3334 3239 3335
rect 3235 3329 3239 3330
rect 3371 3334 3375 3335
rect 3371 3329 3375 3330
rect 3451 3334 3455 3335
rect 3451 3329 3455 3330
rect 3555 3334 3559 3335
rect 3555 3329 3559 3330
rect 3651 3334 3655 3335
rect 3651 3329 3655 3330
rect 3799 3334 3803 3335
rect 3799 3329 3803 3330
rect 2346 3319 2352 3320
rect 2346 3315 2347 3319
rect 2351 3315 2352 3319
rect 2346 3314 2352 3315
rect 2412 3268 2414 3329
rect 2620 3268 2622 3329
rect 2626 3315 2632 3316
rect 2626 3311 2627 3315
rect 2631 3311 2632 3315
rect 2626 3310 2632 3311
rect 2628 3276 2630 3310
rect 2626 3275 2632 3276
rect 2626 3271 2627 3275
rect 2631 3271 2632 3275
rect 2626 3270 2632 3271
rect 2730 3275 2736 3276
rect 2730 3271 2731 3275
rect 2735 3271 2736 3275
rect 2730 3270 2736 3271
rect 1974 3264 1975 3268
rect 1979 3264 1980 3268
rect 1974 3263 1980 3264
rect 1994 3267 2000 3268
rect 1994 3263 1995 3267
rect 1999 3263 2000 3267
rect 1994 3262 2000 3263
rect 2194 3267 2200 3268
rect 2194 3263 2195 3267
rect 2199 3263 2200 3267
rect 2194 3262 2200 3263
rect 2410 3267 2416 3268
rect 2410 3263 2411 3267
rect 2415 3263 2416 3267
rect 2410 3262 2416 3263
rect 2618 3267 2624 3268
rect 2618 3263 2619 3267
rect 2623 3263 2624 3267
rect 2618 3262 2624 3263
rect 2022 3252 2028 3253
rect 1974 3251 1980 3252
rect 1974 3247 1975 3251
rect 1979 3247 1980 3251
rect 2022 3248 2023 3252
rect 2027 3248 2028 3252
rect 2022 3247 2028 3248
rect 2222 3252 2228 3253
rect 2222 3248 2223 3252
rect 2227 3248 2228 3252
rect 2222 3247 2228 3248
rect 2438 3252 2444 3253
rect 2438 3248 2439 3252
rect 2443 3248 2444 3252
rect 2438 3247 2444 3248
rect 2646 3252 2652 3253
rect 2646 3248 2647 3252
rect 2651 3248 2652 3252
rect 2646 3247 2652 3248
rect 1974 3246 1980 3247
rect 1976 3223 1978 3246
rect 2024 3223 2026 3247
rect 2224 3223 2226 3247
rect 2440 3223 2442 3247
rect 2648 3223 2650 3247
rect 1975 3222 1979 3223
rect 1975 3217 1979 3218
rect 2023 3222 2027 3223
rect 2023 3217 2027 3218
rect 2223 3222 2227 3223
rect 2223 3217 2227 3218
rect 2439 3222 2443 3223
rect 2439 3217 2443 3218
rect 2463 3222 2467 3223
rect 2463 3217 2467 3218
rect 2647 3222 2651 3223
rect 2647 3217 2651 3218
rect 2663 3222 2667 3223
rect 2663 3217 2667 3218
rect 1976 3194 1978 3217
rect 1974 3193 1980 3194
rect 2464 3193 2466 3217
rect 2664 3193 2666 3217
rect 1974 3189 1975 3193
rect 1979 3189 1980 3193
rect 1974 3188 1980 3189
rect 2462 3192 2468 3193
rect 2462 3188 2463 3192
rect 2467 3188 2468 3192
rect 2462 3187 2468 3188
rect 2662 3192 2668 3193
rect 2662 3188 2663 3192
rect 2667 3188 2668 3192
rect 2662 3187 2668 3188
rect 2434 3177 2440 3178
rect 1974 3176 1980 3177
rect 1974 3172 1975 3176
rect 1979 3172 1980 3176
rect 2434 3173 2435 3177
rect 2439 3173 2440 3177
rect 2434 3172 2440 3173
rect 2634 3177 2640 3178
rect 2634 3173 2635 3177
rect 2639 3173 2640 3177
rect 2634 3172 2640 3173
rect 1974 3171 1980 3172
rect 1950 3155 1956 3156
rect 1950 3151 1951 3155
rect 1955 3151 1956 3155
rect 1950 3150 1956 3151
rect 1627 3130 1631 3131
rect 1627 3125 1631 3126
rect 1651 3130 1655 3131
rect 1651 3125 1655 3126
rect 1787 3130 1791 3131
rect 1787 3125 1791 3126
rect 1935 3130 1939 3131
rect 1935 3125 1939 3126
rect 1566 3115 1572 3116
rect 1566 3111 1567 3115
rect 1571 3111 1572 3115
rect 1566 3110 1572 3111
rect 1652 3064 1654 3125
rect 1658 3111 1664 3112
rect 1658 3107 1659 3111
rect 1663 3107 1664 3111
rect 1658 3106 1664 3107
rect 1660 3072 1662 3106
rect 1658 3071 1664 3072
rect 1658 3067 1659 3071
rect 1663 3067 1664 3071
rect 1658 3066 1664 3067
rect 1788 3064 1790 3125
rect 1794 3111 1800 3112
rect 1794 3107 1795 3111
rect 1799 3107 1800 3111
rect 1794 3106 1800 3107
rect 1796 3072 1798 3106
rect 1794 3071 1800 3072
rect 1794 3067 1795 3071
rect 1799 3067 1800 3071
rect 1794 3066 1800 3067
rect 1906 3071 1912 3072
rect 1906 3067 1907 3071
rect 1911 3067 1912 3071
rect 1906 3066 1912 3067
rect 562 3063 568 3064
rect 562 3059 563 3063
rect 567 3059 568 3063
rect 562 3058 568 3059
rect 698 3063 704 3064
rect 698 3059 699 3063
rect 703 3059 704 3063
rect 698 3058 704 3059
rect 834 3063 840 3064
rect 834 3059 835 3063
rect 839 3059 840 3063
rect 834 3058 840 3059
rect 970 3063 976 3064
rect 970 3059 971 3063
rect 975 3059 976 3063
rect 970 3058 976 3059
rect 1106 3063 1112 3064
rect 1106 3059 1107 3063
rect 1111 3059 1112 3063
rect 1106 3058 1112 3059
rect 1242 3063 1248 3064
rect 1242 3059 1243 3063
rect 1247 3059 1248 3063
rect 1242 3058 1248 3059
rect 1378 3063 1384 3064
rect 1378 3059 1379 3063
rect 1383 3059 1384 3063
rect 1378 3058 1384 3059
rect 1514 3063 1520 3064
rect 1514 3059 1515 3063
rect 1519 3059 1520 3063
rect 1514 3058 1520 3059
rect 1650 3063 1656 3064
rect 1650 3059 1651 3063
rect 1655 3059 1656 3063
rect 1650 3058 1656 3059
rect 1786 3063 1792 3064
rect 1786 3059 1787 3063
rect 1791 3059 1792 3063
rect 1786 3058 1792 3059
rect 454 3048 460 3049
rect 454 3044 455 3048
rect 459 3044 460 3048
rect 454 3043 460 3044
rect 590 3048 596 3049
rect 590 3044 591 3048
rect 595 3044 596 3048
rect 590 3043 596 3044
rect 726 3048 732 3049
rect 726 3044 727 3048
rect 731 3044 732 3048
rect 726 3043 732 3044
rect 862 3048 868 3049
rect 862 3044 863 3048
rect 867 3044 868 3048
rect 862 3043 868 3044
rect 998 3048 1004 3049
rect 998 3044 999 3048
rect 1003 3044 1004 3048
rect 998 3043 1004 3044
rect 1134 3048 1140 3049
rect 1134 3044 1135 3048
rect 1139 3044 1140 3048
rect 1134 3043 1140 3044
rect 1270 3048 1276 3049
rect 1270 3044 1271 3048
rect 1275 3044 1276 3048
rect 1270 3043 1276 3044
rect 1406 3048 1412 3049
rect 1406 3044 1407 3048
rect 1411 3044 1412 3048
rect 1406 3043 1412 3044
rect 1542 3048 1548 3049
rect 1542 3044 1543 3048
rect 1547 3044 1548 3048
rect 1542 3043 1548 3044
rect 1678 3048 1684 3049
rect 1678 3044 1679 3048
rect 1683 3044 1684 3048
rect 1678 3043 1684 3044
rect 1814 3048 1820 3049
rect 1814 3044 1815 3048
rect 1819 3044 1820 3048
rect 1814 3043 1820 3044
rect 456 2991 458 3043
rect 592 2991 594 3043
rect 728 2991 730 3043
rect 864 2991 866 3043
rect 1000 2991 1002 3043
rect 1136 2991 1138 3043
rect 1272 2991 1274 3043
rect 1408 2991 1410 3043
rect 1544 2991 1546 3043
rect 1680 2991 1682 3043
rect 1816 2991 1818 3043
rect 455 2990 459 2991
rect 455 2985 459 2986
rect 511 2990 515 2991
rect 511 2985 515 2986
rect 591 2990 595 2991
rect 591 2985 595 2986
rect 727 2990 731 2991
rect 727 2985 731 2986
rect 815 2990 819 2991
rect 815 2985 819 2986
rect 863 2990 867 2991
rect 863 2985 867 2986
rect 999 2990 1003 2991
rect 999 2985 1003 2986
rect 1111 2990 1115 2991
rect 1111 2985 1115 2986
rect 1135 2990 1139 2991
rect 1135 2985 1139 2986
rect 1271 2990 1275 2991
rect 1271 2985 1275 2986
rect 1407 2990 1411 2991
rect 1407 2985 1411 2986
rect 1415 2990 1419 2991
rect 1415 2985 1419 2986
rect 1543 2990 1547 2991
rect 1543 2985 1547 2986
rect 1679 2990 1683 2991
rect 1679 2985 1683 2986
rect 1719 2990 1723 2991
rect 1719 2985 1723 2986
rect 1815 2990 1819 2991
rect 1815 2985 1819 2986
rect 512 2961 514 2985
rect 816 2961 818 2985
rect 1112 2961 1114 2985
rect 1416 2961 1418 2985
rect 1720 2961 1722 2985
rect 510 2960 516 2961
rect 510 2956 511 2960
rect 515 2956 516 2960
rect 510 2955 516 2956
rect 814 2960 820 2961
rect 814 2956 815 2960
rect 819 2956 820 2960
rect 814 2955 820 2956
rect 1110 2960 1116 2961
rect 1110 2956 1111 2960
rect 1115 2956 1116 2960
rect 1110 2955 1116 2956
rect 1414 2960 1420 2961
rect 1414 2956 1415 2960
rect 1419 2956 1420 2960
rect 1414 2955 1420 2956
rect 1718 2960 1724 2961
rect 1718 2956 1719 2960
rect 1723 2956 1724 2960
rect 1718 2955 1724 2956
rect 482 2945 488 2946
rect 482 2941 483 2945
rect 487 2941 488 2945
rect 482 2940 488 2941
rect 786 2945 792 2946
rect 786 2941 787 2945
rect 791 2941 792 2945
rect 786 2940 792 2941
rect 1082 2945 1088 2946
rect 1082 2941 1083 2945
rect 1087 2941 1088 2945
rect 1082 2940 1088 2941
rect 1386 2945 1392 2946
rect 1386 2941 1387 2945
rect 1391 2941 1392 2945
rect 1386 2940 1392 2941
rect 1690 2945 1696 2946
rect 1690 2941 1691 2945
rect 1695 2941 1696 2945
rect 1690 2940 1696 2941
rect 434 2935 440 2936
rect 434 2931 435 2935
rect 439 2931 440 2935
rect 434 2930 440 2931
rect 442 2935 448 2936
rect 442 2931 443 2935
rect 447 2931 448 2935
rect 442 2930 448 2931
rect 444 2896 446 2930
rect 442 2895 448 2896
rect 442 2891 443 2895
rect 447 2891 448 2895
rect 442 2890 448 2891
rect 484 2879 486 2940
rect 722 2935 728 2936
rect 722 2931 723 2935
rect 727 2931 728 2935
rect 722 2930 728 2931
rect 724 2896 726 2930
rect 722 2895 728 2896
rect 722 2891 723 2895
rect 727 2891 728 2895
rect 722 2890 728 2891
rect 788 2879 790 2940
rect 1026 2895 1032 2896
rect 1026 2891 1027 2895
rect 1031 2891 1032 2895
rect 1026 2890 1032 2891
rect 111 2878 115 2879
rect 111 2873 115 2874
rect 131 2878 135 2879
rect 131 2873 135 2874
rect 171 2878 175 2879
rect 171 2873 175 2874
rect 307 2878 311 2879
rect 307 2873 311 2874
rect 483 2878 487 2879
rect 483 2873 487 2874
rect 523 2878 527 2879
rect 523 2873 527 2874
rect 763 2878 767 2879
rect 763 2873 767 2874
rect 787 2878 791 2879
rect 787 2873 791 2874
rect 1011 2878 1015 2879
rect 1011 2873 1015 2874
rect 112 2813 114 2873
rect 110 2812 116 2813
rect 132 2812 134 2873
rect 298 2863 304 2864
rect 298 2859 299 2863
rect 303 2859 304 2863
rect 298 2858 304 2859
rect 110 2808 111 2812
rect 115 2808 116 2812
rect 110 2807 116 2808
rect 130 2811 136 2812
rect 130 2807 131 2811
rect 135 2807 136 2811
rect 130 2806 136 2807
rect 158 2796 164 2797
rect 110 2795 116 2796
rect 110 2791 111 2795
rect 115 2791 116 2795
rect 158 2792 159 2796
rect 163 2792 164 2796
rect 158 2791 164 2792
rect 110 2790 116 2791
rect 112 2763 114 2790
rect 160 2763 162 2791
rect 111 2762 115 2763
rect 111 2757 115 2758
rect 159 2762 163 2763
rect 159 2757 163 2758
rect 279 2762 283 2763
rect 279 2757 283 2758
rect 112 2734 114 2757
rect 110 2733 116 2734
rect 280 2733 282 2757
rect 110 2729 111 2733
rect 115 2729 116 2733
rect 110 2728 116 2729
rect 278 2732 284 2733
rect 278 2728 279 2732
rect 283 2728 284 2732
rect 278 2727 284 2728
rect 250 2717 256 2718
rect 110 2716 116 2717
rect 110 2712 111 2716
rect 115 2712 116 2716
rect 250 2713 251 2717
rect 255 2713 256 2717
rect 250 2712 256 2713
rect 110 2711 116 2712
rect 112 2651 114 2711
rect 252 2651 254 2712
rect 300 2708 302 2858
rect 308 2812 310 2873
rect 314 2859 320 2860
rect 314 2855 315 2859
rect 319 2855 320 2859
rect 314 2854 320 2855
rect 316 2820 318 2854
rect 314 2819 320 2820
rect 314 2815 315 2819
rect 319 2815 320 2819
rect 314 2814 320 2815
rect 524 2812 526 2873
rect 530 2859 536 2860
rect 530 2855 531 2859
rect 535 2855 536 2859
rect 530 2854 536 2855
rect 532 2820 534 2854
rect 530 2819 536 2820
rect 530 2815 531 2819
rect 535 2815 536 2819
rect 530 2814 536 2815
rect 764 2812 766 2873
rect 770 2859 776 2860
rect 770 2855 771 2859
rect 775 2855 776 2859
rect 770 2854 776 2855
rect 772 2820 774 2854
rect 770 2819 776 2820
rect 770 2815 771 2819
rect 775 2815 776 2819
rect 770 2814 776 2815
rect 1012 2812 1014 2873
rect 1018 2859 1024 2860
rect 1018 2855 1019 2859
rect 1023 2855 1024 2859
rect 1018 2854 1024 2855
rect 1020 2820 1022 2854
rect 1028 2820 1030 2890
rect 1084 2879 1086 2940
rect 1210 2935 1216 2936
rect 1210 2931 1211 2935
rect 1215 2931 1216 2935
rect 1210 2930 1216 2931
rect 1083 2878 1087 2879
rect 1083 2873 1087 2874
rect 1212 2864 1214 2930
rect 1388 2879 1390 2940
rect 1670 2935 1676 2936
rect 1670 2931 1671 2935
rect 1675 2931 1676 2935
rect 1670 2930 1676 2931
rect 1672 2896 1674 2930
rect 1670 2895 1676 2896
rect 1670 2891 1671 2895
rect 1675 2891 1676 2895
rect 1670 2890 1676 2891
rect 1692 2879 1694 2940
rect 1908 2896 1910 3066
rect 1936 3065 1938 3125
rect 1976 3099 1978 3171
rect 2426 3167 2432 3168
rect 2426 3163 2427 3167
rect 2431 3163 2432 3167
rect 2426 3162 2432 3163
rect 1975 3098 1979 3099
rect 1975 3093 1979 3094
rect 2331 3098 2335 3099
rect 2331 3093 2335 3094
rect 1934 3064 1940 3065
rect 1934 3060 1935 3064
rect 1939 3060 1940 3064
rect 1934 3059 1940 3060
rect 1934 3047 1940 3048
rect 1934 3043 1935 3047
rect 1939 3043 1940 3047
rect 1934 3042 1940 3043
rect 1936 2991 1938 3042
rect 1976 3033 1978 3093
rect 1974 3032 1980 3033
rect 2332 3032 2334 3093
rect 2428 3084 2430 3162
rect 2436 3099 2438 3172
rect 2636 3099 2638 3172
rect 2732 3128 2734 3270
rect 2812 3268 2814 3329
rect 2906 3315 2912 3316
rect 2906 3311 2907 3315
rect 2911 3311 2912 3315
rect 2906 3310 2912 3311
rect 2810 3267 2816 3268
rect 2810 3263 2811 3267
rect 2815 3263 2816 3267
rect 2810 3262 2816 3263
rect 2838 3252 2844 3253
rect 2838 3248 2839 3252
rect 2843 3248 2844 3252
rect 2838 3247 2844 3248
rect 2840 3223 2842 3247
rect 2839 3222 2843 3223
rect 2839 3217 2843 3218
rect 2863 3222 2867 3223
rect 2863 3217 2867 3218
rect 2864 3193 2866 3217
rect 2862 3192 2868 3193
rect 2862 3188 2863 3192
rect 2867 3188 2868 3192
rect 2862 3187 2868 3188
rect 2834 3177 2840 3178
rect 2834 3173 2835 3177
rect 2839 3173 2840 3177
rect 2834 3172 2840 3173
rect 2730 3127 2736 3128
rect 2730 3123 2731 3127
rect 2735 3123 2736 3127
rect 2730 3122 2736 3123
rect 2836 3099 2838 3172
rect 2908 3168 2910 3310
rect 3004 3268 3006 3329
rect 3010 3315 3016 3316
rect 3010 3311 3011 3315
rect 3015 3311 3016 3315
rect 3010 3310 3016 3311
rect 3012 3276 3014 3310
rect 3010 3275 3016 3276
rect 3010 3271 3011 3275
rect 3015 3271 3016 3275
rect 3010 3270 3016 3271
rect 3188 3268 3190 3329
rect 3194 3315 3200 3316
rect 3194 3311 3195 3315
rect 3199 3311 3200 3315
rect 3194 3310 3200 3311
rect 3196 3276 3198 3310
rect 3194 3275 3200 3276
rect 3194 3271 3195 3275
rect 3199 3271 3200 3275
rect 3194 3270 3200 3271
rect 3372 3268 3374 3329
rect 3378 3315 3384 3316
rect 3378 3311 3379 3315
rect 3383 3311 3384 3315
rect 3378 3310 3384 3311
rect 3380 3276 3382 3310
rect 3378 3275 3384 3276
rect 3378 3271 3379 3275
rect 3383 3271 3384 3275
rect 3378 3270 3384 3271
rect 3556 3268 3558 3329
rect 3562 3315 3568 3316
rect 3562 3311 3563 3315
rect 3567 3311 3568 3315
rect 3562 3310 3568 3311
rect 3564 3276 3566 3310
rect 3562 3275 3568 3276
rect 3562 3271 3563 3275
rect 3567 3271 3568 3275
rect 3562 3270 3568 3271
rect 3678 3275 3684 3276
rect 3678 3271 3679 3275
rect 3683 3271 3684 3275
rect 3678 3270 3684 3271
rect 3002 3267 3008 3268
rect 3002 3263 3003 3267
rect 3007 3263 3008 3267
rect 3002 3262 3008 3263
rect 3186 3267 3192 3268
rect 3186 3263 3187 3267
rect 3191 3263 3192 3267
rect 3186 3262 3192 3263
rect 3370 3267 3376 3268
rect 3370 3263 3371 3267
rect 3375 3263 3376 3267
rect 3370 3262 3376 3263
rect 3554 3267 3560 3268
rect 3554 3263 3555 3267
rect 3559 3263 3560 3267
rect 3554 3262 3560 3263
rect 3030 3252 3036 3253
rect 3030 3248 3031 3252
rect 3035 3248 3036 3252
rect 3030 3247 3036 3248
rect 3214 3252 3220 3253
rect 3214 3248 3215 3252
rect 3219 3248 3220 3252
rect 3214 3247 3220 3248
rect 3398 3252 3404 3253
rect 3398 3248 3399 3252
rect 3403 3248 3404 3252
rect 3398 3247 3404 3248
rect 3582 3252 3588 3253
rect 3582 3248 3583 3252
rect 3587 3248 3588 3252
rect 3582 3247 3588 3248
rect 3032 3223 3034 3247
rect 3216 3223 3218 3247
rect 3400 3223 3402 3247
rect 3584 3223 3586 3247
rect 3031 3222 3035 3223
rect 3031 3217 3035 3218
rect 3055 3222 3059 3223
rect 3055 3217 3059 3218
rect 3215 3222 3219 3223
rect 3215 3217 3219 3218
rect 3239 3222 3243 3223
rect 3239 3217 3243 3218
rect 3399 3222 3403 3223
rect 3399 3217 3403 3218
rect 3431 3222 3435 3223
rect 3431 3217 3435 3218
rect 3583 3222 3587 3223
rect 3583 3217 3587 3218
rect 3623 3222 3627 3223
rect 3623 3217 3627 3218
rect 3056 3193 3058 3217
rect 3240 3193 3242 3217
rect 3432 3193 3434 3217
rect 3624 3193 3626 3217
rect 3054 3192 3060 3193
rect 3054 3188 3055 3192
rect 3059 3188 3060 3192
rect 3054 3187 3060 3188
rect 3238 3192 3244 3193
rect 3238 3188 3239 3192
rect 3243 3188 3244 3192
rect 3238 3187 3244 3188
rect 3430 3192 3436 3193
rect 3430 3188 3431 3192
rect 3435 3188 3436 3192
rect 3430 3187 3436 3188
rect 3622 3192 3628 3193
rect 3622 3188 3623 3192
rect 3627 3188 3628 3192
rect 3622 3187 3628 3188
rect 3026 3177 3032 3178
rect 3026 3173 3027 3177
rect 3031 3173 3032 3177
rect 3026 3172 3032 3173
rect 3210 3177 3216 3178
rect 3210 3173 3211 3177
rect 3215 3173 3216 3177
rect 3210 3172 3216 3173
rect 3402 3177 3408 3178
rect 3402 3173 3403 3177
rect 3407 3173 3408 3177
rect 3402 3172 3408 3173
rect 3594 3177 3600 3178
rect 3594 3173 3595 3177
rect 3599 3173 3600 3177
rect 3594 3172 3600 3173
rect 2906 3167 2912 3168
rect 2906 3163 2907 3167
rect 2911 3163 2912 3167
rect 2906 3162 2912 3163
rect 3028 3099 3030 3172
rect 3122 3127 3128 3128
rect 3122 3123 3123 3127
rect 3127 3123 3128 3127
rect 3122 3122 3128 3123
rect 2435 3098 2439 3099
rect 2435 3093 2439 3094
rect 2555 3098 2559 3099
rect 2555 3093 2559 3094
rect 2635 3098 2639 3099
rect 2635 3093 2639 3094
rect 2779 3098 2783 3099
rect 2779 3093 2783 3094
rect 2835 3098 2839 3099
rect 2835 3093 2839 3094
rect 3003 3098 3007 3099
rect 3003 3093 3007 3094
rect 3027 3098 3031 3099
rect 3027 3093 3031 3094
rect 2426 3083 2432 3084
rect 2426 3079 2427 3083
rect 2431 3079 2432 3083
rect 2426 3078 2432 3079
rect 2556 3032 2558 3093
rect 2562 3079 2568 3080
rect 2562 3075 2563 3079
rect 2567 3075 2568 3079
rect 2562 3074 2568 3075
rect 2564 3040 2566 3074
rect 2562 3039 2568 3040
rect 2562 3035 2563 3039
rect 2567 3035 2568 3039
rect 2562 3034 2568 3035
rect 2610 3039 2616 3040
rect 2610 3035 2611 3039
rect 2615 3035 2616 3039
rect 2610 3034 2616 3035
rect 1974 3028 1975 3032
rect 1979 3028 1980 3032
rect 1974 3027 1980 3028
rect 2330 3031 2336 3032
rect 2330 3027 2331 3031
rect 2335 3027 2336 3031
rect 2330 3026 2336 3027
rect 2554 3031 2560 3032
rect 2554 3027 2555 3031
rect 2559 3027 2560 3031
rect 2554 3026 2560 3027
rect 2358 3016 2364 3017
rect 1974 3015 1980 3016
rect 1974 3011 1975 3015
rect 1979 3011 1980 3015
rect 2358 3012 2359 3016
rect 2363 3012 2364 3016
rect 2358 3011 2364 3012
rect 2582 3016 2588 3017
rect 2582 3012 2583 3016
rect 2587 3012 2588 3016
rect 2582 3011 2588 3012
rect 1974 3010 1980 3011
rect 1935 2990 1939 2991
rect 1935 2985 1939 2986
rect 1936 2962 1938 2985
rect 1976 2975 1978 3010
rect 2360 2975 2362 3011
rect 2584 2975 2586 3011
rect 1975 2974 1979 2975
rect 1975 2969 1979 2970
rect 2143 2974 2147 2975
rect 2143 2969 2147 2970
rect 2343 2974 2347 2975
rect 2343 2969 2347 2970
rect 2359 2974 2363 2975
rect 2359 2969 2363 2970
rect 2543 2974 2547 2975
rect 2543 2969 2547 2970
rect 2583 2974 2587 2975
rect 2583 2969 2587 2970
rect 1934 2961 1940 2962
rect 1934 2957 1935 2961
rect 1939 2957 1940 2961
rect 1934 2956 1940 2957
rect 1976 2946 1978 2969
rect 1974 2945 1980 2946
rect 2144 2945 2146 2969
rect 2344 2945 2346 2969
rect 2544 2945 2546 2969
rect 1934 2944 1940 2945
rect 1934 2940 1935 2944
rect 1939 2940 1940 2944
rect 1974 2941 1975 2945
rect 1979 2941 1980 2945
rect 1974 2940 1980 2941
rect 2142 2944 2148 2945
rect 2142 2940 2143 2944
rect 2147 2940 2148 2944
rect 1934 2939 1940 2940
rect 2142 2939 2148 2940
rect 2342 2944 2348 2945
rect 2342 2940 2343 2944
rect 2347 2940 2348 2944
rect 2342 2939 2348 2940
rect 2542 2944 2548 2945
rect 2542 2940 2543 2944
rect 2547 2940 2548 2944
rect 2542 2939 2548 2940
rect 1906 2895 1912 2896
rect 1906 2891 1907 2895
rect 1911 2891 1912 2895
rect 1906 2890 1912 2891
rect 1936 2879 1938 2939
rect 2114 2929 2120 2930
rect 1974 2928 1980 2929
rect 1974 2924 1975 2928
rect 1979 2924 1980 2928
rect 2114 2925 2115 2929
rect 2119 2925 2120 2929
rect 2114 2924 2120 2925
rect 2314 2929 2320 2930
rect 2314 2925 2315 2929
rect 2319 2925 2320 2929
rect 2314 2924 2320 2925
rect 2514 2929 2520 2930
rect 2514 2925 2515 2929
rect 2519 2925 2520 2929
rect 2514 2924 2520 2925
rect 1974 2923 1980 2924
rect 1275 2878 1279 2879
rect 1275 2873 1279 2874
rect 1387 2878 1391 2879
rect 1387 2873 1391 2874
rect 1539 2878 1543 2879
rect 1539 2873 1543 2874
rect 1691 2878 1695 2879
rect 1691 2873 1695 2874
rect 1935 2878 1939 2879
rect 1935 2873 1939 2874
rect 1210 2863 1216 2864
rect 1210 2859 1211 2863
rect 1215 2859 1216 2863
rect 1210 2858 1216 2859
rect 1018 2819 1024 2820
rect 1018 2815 1019 2819
rect 1023 2815 1024 2819
rect 1018 2814 1024 2815
rect 1026 2819 1032 2820
rect 1026 2815 1027 2819
rect 1031 2815 1032 2819
rect 1026 2814 1032 2815
rect 1276 2812 1278 2873
rect 1540 2812 1542 2873
rect 1546 2859 1552 2860
rect 1546 2855 1547 2859
rect 1551 2855 1552 2859
rect 1546 2854 1552 2855
rect 1548 2820 1550 2854
rect 1546 2819 1552 2820
rect 1546 2815 1547 2819
rect 1551 2815 1552 2819
rect 1546 2814 1552 2815
rect 1618 2819 1624 2820
rect 1618 2815 1619 2819
rect 1623 2815 1624 2819
rect 1618 2814 1624 2815
rect 306 2811 312 2812
rect 306 2807 307 2811
rect 311 2807 312 2811
rect 306 2806 312 2807
rect 522 2811 528 2812
rect 522 2807 523 2811
rect 527 2807 528 2811
rect 522 2806 528 2807
rect 762 2811 768 2812
rect 762 2807 763 2811
rect 767 2807 768 2811
rect 762 2806 768 2807
rect 1010 2811 1016 2812
rect 1010 2807 1011 2811
rect 1015 2807 1016 2811
rect 1010 2806 1016 2807
rect 1274 2811 1280 2812
rect 1274 2807 1275 2811
rect 1279 2807 1280 2811
rect 1274 2806 1280 2807
rect 1538 2811 1544 2812
rect 1538 2807 1539 2811
rect 1543 2807 1544 2811
rect 1538 2806 1544 2807
rect 334 2796 340 2797
rect 334 2792 335 2796
rect 339 2792 340 2796
rect 334 2791 340 2792
rect 550 2796 556 2797
rect 550 2792 551 2796
rect 555 2792 556 2796
rect 550 2791 556 2792
rect 790 2796 796 2797
rect 790 2792 791 2796
rect 795 2792 796 2796
rect 790 2791 796 2792
rect 1038 2796 1044 2797
rect 1038 2792 1039 2796
rect 1043 2792 1044 2796
rect 1038 2791 1044 2792
rect 1302 2796 1308 2797
rect 1302 2792 1303 2796
rect 1307 2792 1308 2796
rect 1302 2791 1308 2792
rect 1566 2796 1572 2797
rect 1566 2792 1567 2796
rect 1571 2792 1572 2796
rect 1566 2791 1572 2792
rect 336 2763 338 2791
rect 552 2763 554 2791
rect 792 2763 794 2791
rect 1040 2763 1042 2791
rect 1304 2763 1306 2791
rect 1568 2763 1570 2791
rect 335 2762 339 2763
rect 335 2757 339 2758
rect 455 2762 459 2763
rect 455 2757 459 2758
rect 551 2762 555 2763
rect 551 2757 555 2758
rect 647 2762 651 2763
rect 647 2757 651 2758
rect 791 2762 795 2763
rect 791 2757 795 2758
rect 855 2762 859 2763
rect 855 2757 859 2758
rect 1039 2762 1043 2763
rect 1039 2757 1043 2758
rect 1079 2762 1083 2763
rect 1079 2757 1083 2758
rect 1303 2762 1307 2763
rect 1303 2757 1307 2758
rect 1311 2762 1315 2763
rect 1311 2757 1315 2758
rect 1551 2762 1555 2763
rect 1551 2757 1555 2758
rect 1567 2762 1571 2763
rect 1567 2757 1571 2758
rect 456 2733 458 2757
rect 648 2733 650 2757
rect 856 2733 858 2757
rect 1080 2733 1082 2757
rect 1312 2733 1314 2757
rect 1552 2733 1554 2757
rect 454 2732 460 2733
rect 454 2728 455 2732
rect 459 2728 460 2732
rect 454 2727 460 2728
rect 646 2732 652 2733
rect 646 2728 647 2732
rect 651 2728 652 2732
rect 646 2727 652 2728
rect 854 2732 860 2733
rect 854 2728 855 2732
rect 859 2728 860 2732
rect 854 2727 860 2728
rect 1078 2732 1084 2733
rect 1078 2728 1079 2732
rect 1083 2728 1084 2732
rect 1078 2727 1084 2728
rect 1310 2732 1316 2733
rect 1310 2728 1311 2732
rect 1315 2728 1316 2732
rect 1310 2727 1316 2728
rect 1550 2732 1556 2733
rect 1550 2728 1551 2732
rect 1555 2728 1556 2732
rect 1550 2727 1556 2728
rect 426 2717 432 2718
rect 426 2713 427 2717
rect 431 2713 432 2717
rect 426 2712 432 2713
rect 618 2717 624 2718
rect 618 2713 619 2717
rect 623 2713 624 2717
rect 618 2712 624 2713
rect 826 2717 832 2718
rect 826 2713 827 2717
rect 831 2713 832 2717
rect 826 2712 832 2713
rect 1050 2717 1056 2718
rect 1050 2713 1051 2717
rect 1055 2713 1056 2717
rect 1050 2712 1056 2713
rect 1282 2717 1288 2718
rect 1282 2713 1283 2717
rect 1287 2713 1288 2717
rect 1282 2712 1288 2713
rect 1522 2717 1528 2718
rect 1522 2713 1523 2717
rect 1527 2713 1528 2717
rect 1522 2712 1528 2713
rect 298 2707 304 2708
rect 298 2703 299 2707
rect 303 2703 304 2707
rect 298 2702 304 2703
rect 406 2707 412 2708
rect 406 2703 407 2707
rect 411 2703 412 2707
rect 406 2702 412 2703
rect 408 2668 410 2702
rect 406 2667 412 2668
rect 406 2663 407 2667
rect 411 2663 412 2667
rect 406 2662 412 2663
rect 428 2651 430 2712
rect 620 2651 622 2712
rect 828 2651 830 2712
rect 1018 2667 1024 2668
rect 1018 2663 1019 2667
rect 1023 2663 1024 2667
rect 1018 2662 1024 2663
rect 111 2650 115 2651
rect 111 2645 115 2646
rect 251 2650 255 2651
rect 251 2645 255 2646
rect 427 2650 431 2651
rect 427 2645 431 2646
rect 571 2650 575 2651
rect 571 2645 575 2646
rect 619 2650 623 2651
rect 619 2645 623 2646
rect 731 2650 735 2651
rect 731 2645 735 2646
rect 827 2650 831 2651
rect 827 2645 831 2646
rect 891 2650 895 2651
rect 891 2645 895 2646
rect 112 2585 114 2645
rect 110 2584 116 2585
rect 572 2584 574 2645
rect 732 2584 734 2645
rect 882 2639 888 2640
rect 882 2635 883 2639
rect 887 2635 888 2639
rect 882 2634 888 2635
rect 738 2631 744 2632
rect 738 2627 739 2631
rect 743 2627 744 2631
rect 738 2626 744 2627
rect 740 2592 742 2626
rect 738 2591 744 2592
rect 738 2587 739 2591
rect 743 2587 744 2591
rect 738 2586 744 2587
rect 110 2580 111 2584
rect 115 2580 116 2584
rect 110 2579 116 2580
rect 570 2583 576 2584
rect 570 2579 571 2583
rect 575 2579 576 2583
rect 570 2578 576 2579
rect 730 2583 736 2584
rect 730 2579 731 2583
rect 735 2579 736 2583
rect 730 2578 736 2579
rect 598 2568 604 2569
rect 110 2567 116 2568
rect 110 2563 111 2567
rect 115 2563 116 2567
rect 598 2564 599 2568
rect 603 2564 604 2568
rect 598 2563 604 2564
rect 758 2568 764 2569
rect 758 2564 759 2568
rect 763 2564 764 2568
rect 758 2563 764 2564
rect 110 2562 116 2563
rect 112 2539 114 2562
rect 600 2539 602 2563
rect 760 2539 762 2563
rect 111 2538 115 2539
rect 111 2533 115 2534
rect 383 2538 387 2539
rect 383 2533 387 2534
rect 599 2538 603 2539
rect 599 2533 603 2534
rect 759 2538 763 2539
rect 759 2533 763 2534
rect 815 2538 819 2539
rect 815 2533 819 2534
rect 112 2510 114 2533
rect 110 2509 116 2510
rect 384 2509 386 2533
rect 600 2509 602 2533
rect 816 2509 818 2533
rect 110 2505 111 2509
rect 115 2505 116 2509
rect 110 2504 116 2505
rect 382 2508 388 2509
rect 382 2504 383 2508
rect 387 2504 388 2508
rect 382 2503 388 2504
rect 598 2508 604 2509
rect 598 2504 599 2508
rect 603 2504 604 2508
rect 598 2503 604 2504
rect 814 2508 820 2509
rect 814 2504 815 2508
rect 819 2504 820 2508
rect 814 2503 820 2504
rect 354 2493 360 2494
rect 110 2492 116 2493
rect 110 2488 111 2492
rect 115 2488 116 2492
rect 354 2489 355 2493
rect 359 2489 360 2493
rect 354 2488 360 2489
rect 570 2493 576 2494
rect 570 2489 571 2493
rect 575 2489 576 2493
rect 570 2488 576 2489
rect 786 2493 792 2494
rect 786 2489 787 2493
rect 791 2489 792 2493
rect 786 2488 792 2489
rect 110 2487 116 2488
rect 112 2423 114 2487
rect 356 2423 358 2488
rect 362 2443 368 2444
rect 362 2439 363 2443
rect 367 2439 368 2443
rect 362 2438 368 2439
rect 111 2422 115 2423
rect 111 2417 115 2418
rect 227 2422 231 2423
rect 227 2417 231 2418
rect 355 2422 359 2423
rect 355 2417 359 2418
rect 112 2357 114 2417
rect 110 2356 116 2357
rect 228 2356 230 2417
rect 364 2364 366 2438
rect 572 2423 574 2488
rect 788 2423 790 2488
rect 884 2484 886 2634
rect 892 2584 894 2645
rect 898 2631 904 2632
rect 898 2627 899 2631
rect 903 2627 904 2631
rect 898 2626 904 2627
rect 900 2592 902 2626
rect 1020 2592 1022 2662
rect 1052 2651 1054 2712
rect 1284 2651 1286 2712
rect 1406 2707 1412 2708
rect 1406 2703 1407 2707
rect 1411 2703 1412 2707
rect 1406 2702 1412 2703
rect 1043 2650 1047 2651
rect 1043 2645 1047 2646
rect 1051 2650 1055 2651
rect 1051 2645 1055 2646
rect 1195 2650 1199 2651
rect 1195 2645 1199 2646
rect 1283 2650 1287 2651
rect 1283 2645 1287 2646
rect 1355 2650 1359 2651
rect 1355 2645 1359 2646
rect 898 2591 904 2592
rect 898 2587 899 2591
rect 903 2587 904 2591
rect 898 2586 904 2587
rect 1018 2591 1024 2592
rect 1018 2587 1019 2591
rect 1023 2587 1024 2591
rect 1018 2586 1024 2587
rect 1044 2584 1046 2645
rect 1186 2635 1192 2636
rect 1186 2631 1187 2635
rect 1191 2631 1192 2635
rect 1186 2630 1192 2631
rect 1188 2592 1190 2630
rect 1090 2591 1096 2592
rect 1090 2587 1091 2591
rect 1095 2587 1096 2591
rect 1090 2586 1096 2587
rect 1186 2591 1192 2592
rect 1186 2587 1187 2591
rect 1191 2587 1192 2591
rect 1186 2586 1192 2587
rect 890 2583 896 2584
rect 890 2579 891 2583
rect 895 2579 896 2583
rect 890 2578 896 2579
rect 1042 2583 1048 2584
rect 1042 2579 1043 2583
rect 1047 2579 1048 2583
rect 1042 2578 1048 2579
rect 918 2568 924 2569
rect 918 2564 919 2568
rect 923 2564 924 2568
rect 918 2563 924 2564
rect 1070 2568 1076 2569
rect 1070 2564 1071 2568
rect 1075 2564 1076 2568
rect 1070 2563 1076 2564
rect 920 2539 922 2563
rect 1072 2539 1074 2563
rect 919 2538 923 2539
rect 919 2533 923 2534
rect 1023 2538 1027 2539
rect 1023 2533 1027 2534
rect 1071 2538 1075 2539
rect 1071 2533 1075 2534
rect 1024 2509 1026 2533
rect 1022 2508 1028 2509
rect 1022 2504 1023 2508
rect 1027 2504 1028 2508
rect 1022 2503 1028 2504
rect 994 2493 1000 2494
rect 994 2489 995 2493
rect 999 2489 1000 2493
rect 994 2488 1000 2489
rect 882 2483 888 2484
rect 882 2479 883 2483
rect 887 2479 888 2483
rect 882 2478 888 2479
rect 996 2423 998 2488
rect 1092 2444 1094 2586
rect 1196 2584 1198 2645
rect 1356 2584 1358 2645
rect 1408 2636 1410 2702
rect 1524 2651 1526 2712
rect 1620 2668 1622 2814
rect 1936 2813 1938 2873
rect 1976 2855 1978 2923
rect 2116 2855 2118 2924
rect 2250 2919 2256 2920
rect 2250 2915 2251 2919
rect 2255 2915 2256 2919
rect 2250 2914 2256 2915
rect 2274 2919 2280 2920
rect 2274 2915 2275 2919
rect 2279 2915 2280 2919
rect 2274 2914 2280 2915
rect 1975 2854 1979 2855
rect 1975 2849 1979 2850
rect 2011 2854 2015 2855
rect 2011 2849 2015 2850
rect 2115 2854 2119 2855
rect 2115 2849 2119 2850
rect 1934 2812 1940 2813
rect 1934 2808 1935 2812
rect 1939 2808 1940 2812
rect 1934 2807 1940 2808
rect 1934 2795 1940 2796
rect 1934 2791 1935 2795
rect 1939 2791 1940 2795
rect 1934 2790 1940 2791
rect 1936 2763 1938 2790
rect 1976 2789 1978 2849
rect 1974 2788 1980 2789
rect 2012 2788 2014 2849
rect 2252 2840 2254 2914
rect 2276 2880 2278 2914
rect 2274 2879 2280 2880
rect 2274 2875 2275 2879
rect 2279 2875 2280 2879
rect 2274 2874 2280 2875
rect 2316 2855 2318 2924
rect 2474 2919 2480 2920
rect 2474 2915 2475 2919
rect 2479 2915 2480 2919
rect 2474 2914 2480 2915
rect 2476 2880 2478 2914
rect 2474 2879 2480 2880
rect 2474 2875 2475 2879
rect 2479 2875 2480 2879
rect 2474 2874 2480 2875
rect 2516 2855 2518 2924
rect 2612 2880 2614 3034
rect 2780 3032 2782 3093
rect 2838 3083 2844 3084
rect 2838 3079 2839 3083
rect 2843 3079 2844 3083
rect 2838 3078 2844 3079
rect 2778 3031 2784 3032
rect 2778 3027 2779 3031
rect 2783 3027 2784 3031
rect 2778 3026 2784 3027
rect 2806 3016 2812 3017
rect 2806 3012 2807 3016
rect 2811 3012 2812 3016
rect 2806 3011 2812 3012
rect 2808 2975 2810 3011
rect 2743 2974 2747 2975
rect 2743 2969 2747 2970
rect 2807 2974 2811 2975
rect 2807 2969 2811 2970
rect 2744 2945 2746 2969
rect 2742 2944 2748 2945
rect 2742 2940 2743 2944
rect 2747 2940 2748 2944
rect 2742 2939 2748 2940
rect 2714 2929 2720 2930
rect 2714 2925 2715 2929
rect 2719 2925 2720 2929
rect 2714 2924 2720 2925
rect 2610 2879 2616 2880
rect 2610 2875 2611 2879
rect 2615 2875 2616 2879
rect 2610 2874 2616 2875
rect 2634 2879 2640 2880
rect 2634 2875 2635 2879
rect 2639 2875 2640 2879
rect 2634 2874 2640 2875
rect 2259 2854 2263 2855
rect 2259 2849 2263 2850
rect 2315 2854 2319 2855
rect 2315 2849 2319 2850
rect 2507 2854 2511 2855
rect 2507 2849 2511 2850
rect 2515 2854 2519 2855
rect 2515 2849 2519 2850
rect 2154 2839 2160 2840
rect 2154 2835 2155 2839
rect 2159 2835 2160 2839
rect 2154 2834 2160 2835
rect 2250 2839 2256 2840
rect 2250 2835 2251 2839
rect 2255 2835 2256 2839
rect 2250 2834 2256 2835
rect 2156 2796 2158 2834
rect 2090 2795 2096 2796
rect 2090 2791 2091 2795
rect 2095 2791 2096 2795
rect 2090 2790 2096 2791
rect 2154 2795 2160 2796
rect 2154 2791 2155 2795
rect 2159 2791 2160 2795
rect 2154 2790 2160 2791
rect 1974 2784 1975 2788
rect 1979 2784 1980 2788
rect 1974 2783 1980 2784
rect 2010 2787 2016 2788
rect 2010 2783 2011 2787
rect 2015 2783 2016 2787
rect 2010 2782 2016 2783
rect 2038 2772 2044 2773
rect 1974 2771 1980 2772
rect 1974 2767 1975 2771
rect 1979 2767 1980 2771
rect 2038 2768 2039 2772
rect 2043 2768 2044 2772
rect 2038 2767 2044 2768
rect 1974 2766 1980 2767
rect 1799 2762 1803 2763
rect 1799 2757 1803 2758
rect 1935 2762 1939 2763
rect 1935 2757 1939 2758
rect 1800 2733 1802 2757
rect 1936 2734 1938 2757
rect 1976 2739 1978 2766
rect 2040 2739 2042 2767
rect 1975 2738 1979 2739
rect 1934 2733 1940 2734
rect 1975 2733 1979 2734
rect 2023 2738 2027 2739
rect 2023 2733 2027 2734
rect 2039 2738 2043 2739
rect 2039 2733 2043 2734
rect 1798 2732 1804 2733
rect 1798 2728 1799 2732
rect 1803 2728 1804 2732
rect 1934 2729 1935 2733
rect 1939 2729 1940 2733
rect 1934 2728 1940 2729
rect 1798 2727 1804 2728
rect 1770 2717 1776 2718
rect 1770 2713 1771 2717
rect 1775 2713 1776 2717
rect 1770 2712 1776 2713
rect 1934 2716 1940 2717
rect 1934 2712 1935 2716
rect 1939 2712 1940 2716
rect 1618 2667 1624 2668
rect 1618 2663 1619 2667
rect 1623 2663 1624 2667
rect 1618 2662 1624 2663
rect 1772 2651 1774 2712
rect 1934 2711 1940 2712
rect 1786 2707 1792 2708
rect 1786 2703 1787 2707
rect 1791 2703 1792 2707
rect 1786 2702 1792 2703
rect 1515 2650 1519 2651
rect 1515 2645 1519 2646
rect 1523 2650 1527 2651
rect 1523 2645 1527 2646
rect 1675 2650 1679 2651
rect 1675 2645 1679 2646
rect 1771 2650 1775 2651
rect 1771 2645 1775 2646
rect 1406 2635 1412 2636
rect 1406 2631 1407 2635
rect 1411 2631 1412 2635
rect 1406 2630 1412 2631
rect 1498 2591 1504 2592
rect 1498 2587 1499 2591
rect 1503 2587 1504 2591
rect 1498 2586 1504 2587
rect 1194 2583 1200 2584
rect 1194 2579 1195 2583
rect 1199 2579 1200 2583
rect 1194 2578 1200 2579
rect 1354 2583 1360 2584
rect 1354 2579 1355 2583
rect 1359 2579 1360 2583
rect 1354 2578 1360 2579
rect 1222 2568 1228 2569
rect 1222 2564 1223 2568
rect 1227 2564 1228 2568
rect 1222 2563 1228 2564
rect 1382 2568 1388 2569
rect 1382 2564 1383 2568
rect 1387 2564 1388 2568
rect 1382 2563 1388 2564
rect 1224 2539 1226 2563
rect 1384 2539 1386 2563
rect 1223 2538 1227 2539
rect 1223 2533 1227 2534
rect 1231 2538 1235 2539
rect 1231 2533 1235 2534
rect 1383 2538 1387 2539
rect 1383 2533 1387 2534
rect 1431 2538 1435 2539
rect 1431 2533 1435 2534
rect 1232 2509 1234 2533
rect 1432 2509 1434 2533
rect 1230 2508 1236 2509
rect 1230 2504 1231 2508
rect 1235 2504 1236 2508
rect 1230 2503 1236 2504
rect 1430 2508 1436 2509
rect 1430 2504 1431 2508
rect 1435 2504 1436 2508
rect 1430 2503 1436 2504
rect 1202 2493 1208 2494
rect 1202 2489 1203 2493
rect 1207 2489 1208 2493
rect 1202 2488 1208 2489
rect 1402 2493 1408 2494
rect 1402 2489 1403 2493
rect 1407 2489 1408 2493
rect 1402 2488 1408 2489
rect 1166 2483 1172 2484
rect 1166 2479 1167 2483
rect 1171 2479 1172 2483
rect 1166 2478 1172 2479
rect 1168 2444 1170 2478
rect 1090 2443 1096 2444
rect 1090 2439 1091 2443
rect 1095 2439 1096 2443
rect 1090 2438 1096 2439
rect 1166 2443 1172 2444
rect 1166 2439 1167 2443
rect 1171 2439 1172 2443
rect 1166 2438 1172 2439
rect 1204 2423 1206 2488
rect 1404 2423 1406 2488
rect 1500 2444 1502 2586
rect 1516 2584 1518 2645
rect 1676 2584 1678 2645
rect 1788 2636 1790 2702
rect 1936 2651 1938 2711
rect 1976 2710 1978 2733
rect 1974 2709 1980 2710
rect 2024 2709 2026 2733
rect 1974 2705 1975 2709
rect 1979 2705 1980 2709
rect 1974 2704 1980 2705
rect 2022 2708 2028 2709
rect 2022 2704 2023 2708
rect 2027 2704 2028 2708
rect 2022 2703 2028 2704
rect 1994 2693 2000 2694
rect 1974 2692 1980 2693
rect 1974 2688 1975 2692
rect 1979 2688 1980 2692
rect 1994 2689 1995 2693
rect 1999 2689 2000 2693
rect 1994 2688 2000 2689
rect 1974 2687 1980 2688
rect 1935 2650 1939 2651
rect 1935 2645 1939 2646
rect 1786 2635 1792 2636
rect 1786 2631 1787 2635
rect 1791 2631 1792 2635
rect 1786 2630 1792 2631
rect 1936 2585 1938 2645
rect 1976 2615 1978 2687
rect 1996 2615 1998 2688
rect 2092 2644 2094 2790
rect 2260 2788 2262 2849
rect 2508 2788 2510 2849
rect 2514 2835 2520 2836
rect 2514 2831 2515 2835
rect 2519 2831 2520 2835
rect 2514 2830 2520 2831
rect 2258 2787 2264 2788
rect 2258 2783 2259 2787
rect 2263 2783 2264 2787
rect 2258 2782 2264 2783
rect 2506 2787 2512 2788
rect 2506 2783 2507 2787
rect 2511 2783 2512 2787
rect 2506 2782 2512 2783
rect 2286 2772 2292 2773
rect 2286 2768 2287 2772
rect 2291 2768 2292 2772
rect 2286 2767 2292 2768
rect 2288 2739 2290 2767
rect 2247 2738 2251 2739
rect 2247 2733 2251 2734
rect 2287 2738 2291 2739
rect 2287 2733 2291 2734
rect 2503 2738 2507 2739
rect 2503 2733 2507 2734
rect 2248 2709 2250 2733
rect 2504 2709 2506 2733
rect 2246 2708 2252 2709
rect 2246 2704 2247 2708
rect 2251 2704 2252 2708
rect 2246 2703 2252 2704
rect 2502 2708 2508 2709
rect 2502 2704 2503 2708
rect 2507 2704 2508 2708
rect 2502 2703 2508 2704
rect 2218 2693 2224 2694
rect 2218 2689 2219 2693
rect 2223 2689 2224 2693
rect 2218 2688 2224 2689
rect 2474 2693 2480 2694
rect 2474 2689 2475 2693
rect 2479 2689 2480 2693
rect 2474 2688 2480 2689
rect 2090 2643 2096 2644
rect 2090 2639 2091 2643
rect 2095 2639 2096 2643
rect 2090 2638 2096 2639
rect 2220 2615 2222 2688
rect 2476 2615 2478 2688
rect 2516 2684 2518 2830
rect 2636 2796 2638 2874
rect 2716 2855 2718 2924
rect 2840 2920 2842 3078
rect 3004 3032 3006 3093
rect 3010 3079 3016 3080
rect 3010 3075 3011 3079
rect 3015 3075 3016 3079
rect 3010 3074 3016 3075
rect 3012 3040 3014 3074
rect 3124 3040 3126 3122
rect 3212 3099 3214 3172
rect 3338 3167 3344 3168
rect 3338 3163 3339 3167
rect 3343 3163 3344 3167
rect 3338 3162 3344 3163
rect 3306 3159 3312 3160
rect 3306 3155 3307 3159
rect 3311 3155 3312 3159
rect 3306 3154 3312 3155
rect 3308 3128 3310 3154
rect 3340 3128 3342 3162
rect 3306 3127 3312 3128
rect 3306 3123 3307 3127
rect 3311 3123 3312 3127
rect 3306 3122 3312 3123
rect 3338 3127 3344 3128
rect 3338 3123 3339 3127
rect 3343 3123 3344 3127
rect 3338 3122 3344 3123
rect 3404 3099 3406 3172
rect 3526 3167 3532 3168
rect 3526 3163 3527 3167
rect 3531 3163 3532 3167
rect 3526 3162 3532 3163
rect 3211 3098 3215 3099
rect 3211 3093 3215 3094
rect 3235 3098 3239 3099
rect 3235 3093 3239 3094
rect 3403 3098 3407 3099
rect 3403 3093 3407 3094
rect 3467 3098 3471 3099
rect 3467 3093 3471 3094
rect 3010 3039 3016 3040
rect 3010 3035 3011 3039
rect 3015 3035 3016 3039
rect 3010 3034 3016 3035
rect 3122 3039 3128 3040
rect 3122 3035 3123 3039
rect 3127 3035 3128 3039
rect 3122 3034 3128 3035
rect 3236 3032 3238 3093
rect 3358 3039 3364 3040
rect 3358 3035 3359 3039
rect 3363 3035 3364 3039
rect 3358 3034 3364 3035
rect 3002 3031 3008 3032
rect 3002 3027 3003 3031
rect 3007 3027 3008 3031
rect 3002 3026 3008 3027
rect 3234 3031 3240 3032
rect 3234 3027 3235 3031
rect 3239 3027 3240 3031
rect 3234 3026 3240 3027
rect 3030 3016 3036 3017
rect 3030 3012 3031 3016
rect 3035 3012 3036 3016
rect 3030 3011 3036 3012
rect 3262 3016 3268 3017
rect 3262 3012 3263 3016
rect 3267 3012 3268 3016
rect 3262 3011 3268 3012
rect 3032 2975 3034 3011
rect 3264 2975 3266 3011
rect 2935 2974 2939 2975
rect 2935 2969 2939 2970
rect 3031 2974 3035 2975
rect 3031 2969 3035 2970
rect 3135 2974 3139 2975
rect 3135 2969 3139 2970
rect 3263 2974 3267 2975
rect 3263 2969 3267 2970
rect 3335 2974 3339 2975
rect 3335 2969 3339 2970
rect 2936 2945 2938 2969
rect 3136 2945 3138 2969
rect 3336 2945 3338 2969
rect 2934 2944 2940 2945
rect 2934 2940 2935 2944
rect 2939 2940 2940 2944
rect 2934 2939 2940 2940
rect 3134 2944 3140 2945
rect 3134 2940 3135 2944
rect 3139 2940 3140 2944
rect 3134 2939 3140 2940
rect 3334 2944 3340 2945
rect 3334 2940 3335 2944
rect 3339 2940 3340 2944
rect 3334 2939 3340 2940
rect 2906 2929 2912 2930
rect 2906 2925 2907 2929
rect 2911 2925 2912 2929
rect 2906 2924 2912 2925
rect 3106 2929 3112 2930
rect 3106 2925 3107 2929
rect 3111 2925 3112 2929
rect 3106 2924 3112 2925
rect 3306 2929 3312 2930
rect 3306 2925 3307 2929
rect 3311 2925 3312 2929
rect 3306 2924 3312 2925
rect 2838 2919 2844 2920
rect 2838 2915 2839 2919
rect 2843 2915 2844 2919
rect 2838 2914 2844 2915
rect 2908 2855 2910 2924
rect 3030 2919 3036 2920
rect 3030 2915 3031 2919
rect 3035 2915 3036 2919
rect 3030 2914 3036 2915
rect 3066 2919 3072 2920
rect 3066 2915 3067 2919
rect 3071 2915 3072 2919
rect 3066 2914 3072 2915
rect 2715 2854 2719 2855
rect 2715 2849 2719 2850
rect 2755 2854 2759 2855
rect 2755 2849 2759 2850
rect 2907 2854 2911 2855
rect 2907 2849 2911 2850
rect 3003 2854 3007 2855
rect 3003 2849 3007 2850
rect 2634 2795 2640 2796
rect 2634 2791 2635 2795
rect 2639 2791 2640 2795
rect 2634 2790 2640 2791
rect 2756 2788 2758 2849
rect 2806 2795 2812 2796
rect 2806 2791 2807 2795
rect 2811 2791 2812 2795
rect 2806 2790 2812 2791
rect 2754 2787 2760 2788
rect 2754 2783 2755 2787
rect 2759 2783 2760 2787
rect 2754 2782 2760 2783
rect 2534 2772 2540 2773
rect 2534 2768 2535 2772
rect 2539 2768 2540 2772
rect 2534 2767 2540 2768
rect 2782 2772 2788 2773
rect 2782 2768 2783 2772
rect 2787 2768 2788 2772
rect 2782 2767 2788 2768
rect 2536 2739 2538 2767
rect 2784 2739 2786 2767
rect 2535 2738 2539 2739
rect 2535 2733 2539 2734
rect 2759 2738 2763 2739
rect 2759 2733 2763 2734
rect 2783 2738 2787 2739
rect 2783 2733 2787 2734
rect 2760 2709 2762 2733
rect 2758 2708 2764 2709
rect 2758 2704 2759 2708
rect 2763 2704 2764 2708
rect 2758 2703 2764 2704
rect 2730 2693 2736 2694
rect 2730 2689 2731 2693
rect 2735 2689 2736 2693
rect 2730 2688 2736 2689
rect 2514 2683 2520 2684
rect 2514 2679 2515 2683
rect 2519 2679 2520 2683
rect 2514 2678 2520 2679
rect 2602 2683 2608 2684
rect 2602 2679 2603 2683
rect 2607 2679 2608 2683
rect 2602 2678 2608 2679
rect 2604 2644 2606 2678
rect 2602 2643 2608 2644
rect 2602 2639 2603 2643
rect 2607 2639 2608 2643
rect 2602 2638 2608 2639
rect 2538 2635 2544 2636
rect 2538 2631 2539 2635
rect 2543 2631 2544 2635
rect 2538 2630 2544 2631
rect 1975 2614 1979 2615
rect 1975 2609 1979 2610
rect 1995 2614 1999 2615
rect 1995 2609 1999 2610
rect 2219 2614 2223 2615
rect 2219 2609 2223 2610
rect 2475 2614 2479 2615
rect 2475 2609 2479 2610
rect 1934 2584 1940 2585
rect 1514 2583 1520 2584
rect 1514 2579 1515 2583
rect 1519 2579 1520 2583
rect 1514 2578 1520 2579
rect 1674 2583 1680 2584
rect 1674 2579 1675 2583
rect 1679 2579 1680 2583
rect 1934 2580 1935 2584
rect 1939 2580 1940 2584
rect 1934 2579 1940 2580
rect 1674 2578 1680 2579
rect 1542 2568 1548 2569
rect 1542 2564 1543 2568
rect 1547 2564 1548 2568
rect 1542 2563 1548 2564
rect 1702 2568 1708 2569
rect 1702 2564 1703 2568
rect 1707 2564 1708 2568
rect 1702 2563 1708 2564
rect 1934 2567 1940 2568
rect 1934 2563 1935 2567
rect 1939 2563 1940 2567
rect 1544 2539 1546 2563
rect 1704 2539 1706 2563
rect 1934 2562 1940 2563
rect 1936 2539 1938 2562
rect 1976 2549 1978 2609
rect 2540 2556 2542 2630
rect 2732 2615 2734 2688
rect 2808 2636 2810 2790
rect 3004 2788 3006 2849
rect 3032 2840 3034 2914
rect 3068 2880 3070 2914
rect 3066 2879 3072 2880
rect 3066 2875 3067 2879
rect 3071 2875 3072 2879
rect 3066 2874 3072 2875
rect 3108 2855 3110 2924
rect 3266 2919 3272 2920
rect 3266 2915 3267 2919
rect 3271 2915 3272 2919
rect 3266 2914 3272 2915
rect 3268 2880 3270 2914
rect 3266 2879 3272 2880
rect 3266 2875 3267 2879
rect 3271 2875 3272 2879
rect 3266 2874 3272 2875
rect 3308 2855 3310 2924
rect 3360 2880 3362 3034
rect 3468 3032 3470 3093
rect 3528 3084 3530 3162
rect 3596 3099 3598 3172
rect 3680 3128 3682 3270
rect 3800 3269 3802 3329
rect 3840 3287 3842 3347
rect 3860 3287 3862 3348
rect 3986 3303 3992 3304
rect 3986 3299 3987 3303
rect 3991 3299 3992 3303
rect 3986 3298 3992 3299
rect 3839 3286 3843 3287
rect 3839 3281 3843 3282
rect 3859 3286 3863 3287
rect 3859 3281 3863 3282
rect 3798 3268 3804 3269
rect 3798 3264 3799 3268
rect 3803 3264 3804 3268
rect 3798 3263 3804 3264
rect 3798 3251 3804 3252
rect 3798 3247 3799 3251
rect 3803 3247 3804 3251
rect 3798 3246 3804 3247
rect 3800 3223 3802 3246
rect 3799 3222 3803 3223
rect 3840 3221 3842 3281
rect 3799 3217 3803 3218
rect 3838 3220 3844 3221
rect 3860 3220 3862 3281
rect 3954 3267 3960 3268
rect 3954 3263 3955 3267
rect 3959 3263 3960 3267
rect 3954 3262 3960 3263
rect 3800 3194 3802 3217
rect 3838 3216 3839 3220
rect 3843 3216 3844 3220
rect 3838 3215 3844 3216
rect 3858 3219 3864 3220
rect 3858 3215 3859 3219
rect 3863 3215 3864 3219
rect 3858 3214 3864 3215
rect 3886 3204 3892 3205
rect 3838 3203 3844 3204
rect 3838 3199 3839 3203
rect 3843 3199 3844 3203
rect 3886 3200 3887 3204
rect 3891 3200 3892 3204
rect 3886 3199 3892 3200
rect 3838 3198 3844 3199
rect 3798 3193 3804 3194
rect 3798 3189 3799 3193
rect 3803 3189 3804 3193
rect 3798 3188 3804 3189
rect 3798 3176 3804 3177
rect 3798 3172 3799 3176
rect 3803 3172 3804 3176
rect 3798 3171 3804 3172
rect 3678 3127 3684 3128
rect 3678 3123 3679 3127
rect 3683 3123 3684 3127
rect 3678 3122 3684 3123
rect 3800 3099 3802 3171
rect 3840 3159 3842 3198
rect 3888 3159 3890 3199
rect 3839 3158 3843 3159
rect 3839 3153 3843 3154
rect 3887 3158 3891 3159
rect 3887 3153 3891 3154
rect 3903 3158 3907 3159
rect 3903 3153 3907 3154
rect 3840 3130 3842 3153
rect 3838 3129 3844 3130
rect 3904 3129 3906 3153
rect 3838 3125 3839 3129
rect 3843 3125 3844 3129
rect 3838 3124 3844 3125
rect 3902 3128 3908 3129
rect 3902 3124 3903 3128
rect 3907 3124 3908 3128
rect 3902 3123 3908 3124
rect 3874 3113 3880 3114
rect 3838 3112 3844 3113
rect 3838 3108 3839 3112
rect 3843 3108 3844 3112
rect 3874 3109 3875 3113
rect 3879 3109 3880 3113
rect 3874 3108 3880 3109
rect 3838 3107 3844 3108
rect 3595 3098 3599 3099
rect 3595 3093 3599 3094
rect 3799 3098 3803 3099
rect 3799 3093 3803 3094
rect 3526 3083 3532 3084
rect 3526 3079 3527 3083
rect 3531 3079 3532 3083
rect 3526 3078 3532 3079
rect 3800 3033 3802 3093
rect 3840 3047 3842 3107
rect 3876 3047 3878 3108
rect 3956 3104 3958 3262
rect 3988 3228 3990 3298
rect 4124 3287 4126 3348
rect 4130 3343 4136 3344
rect 4130 3339 4131 3343
rect 4135 3339 4136 3343
rect 4130 3338 4136 3339
rect 4132 3312 4134 3338
rect 4130 3311 4136 3312
rect 4130 3307 4131 3311
rect 4135 3307 4136 3311
rect 4130 3306 4136 3307
rect 4396 3287 4398 3348
rect 4522 3343 4528 3344
rect 4522 3339 4523 3343
rect 4527 3339 4528 3343
rect 4522 3338 4528 3339
rect 4524 3304 4526 3338
rect 4522 3303 4528 3304
rect 4522 3299 4523 3303
rect 4527 3299 4528 3303
rect 4522 3298 4528 3299
rect 4644 3287 4646 3348
rect 4770 3343 4776 3344
rect 4770 3339 4771 3343
rect 4775 3339 4776 3343
rect 4770 3338 4776 3339
rect 4772 3304 4774 3338
rect 4770 3303 4776 3304
rect 4770 3299 4771 3303
rect 4775 3299 4776 3303
rect 4770 3298 4776 3299
rect 4868 3287 4870 3348
rect 5084 3287 5086 3348
rect 5142 3335 5148 3336
rect 5142 3331 5143 3335
rect 5147 3331 5148 3335
rect 5142 3330 5148 3331
rect 4099 3286 4103 3287
rect 4099 3281 4103 3282
rect 4123 3286 4127 3287
rect 4123 3281 4127 3282
rect 4347 3286 4351 3287
rect 4347 3281 4351 3282
rect 4395 3286 4399 3287
rect 4395 3281 4399 3282
rect 4579 3286 4583 3287
rect 4579 3281 4583 3282
rect 4643 3286 4647 3287
rect 4643 3281 4647 3282
rect 4787 3286 4791 3287
rect 4787 3281 4791 3282
rect 4867 3286 4871 3287
rect 4867 3281 4871 3282
rect 4987 3286 4991 3287
rect 4987 3281 4991 3282
rect 5083 3286 5087 3287
rect 5083 3281 5087 3282
rect 3986 3227 3992 3228
rect 3986 3223 3987 3227
rect 3991 3223 3992 3227
rect 3986 3222 3992 3223
rect 4100 3220 4102 3281
rect 4194 3267 4200 3268
rect 4194 3263 4195 3267
rect 4199 3263 4200 3267
rect 4194 3262 4200 3263
rect 4196 3236 4198 3262
rect 4194 3235 4200 3236
rect 4194 3231 4195 3235
rect 4199 3231 4200 3235
rect 4194 3230 4200 3231
rect 4348 3220 4350 3281
rect 4354 3267 4360 3268
rect 4354 3263 4355 3267
rect 4359 3263 4360 3267
rect 4354 3262 4360 3263
rect 4356 3228 4358 3262
rect 4354 3227 4360 3228
rect 4354 3223 4355 3227
rect 4359 3223 4360 3227
rect 4354 3222 4360 3223
rect 4474 3227 4480 3228
rect 4474 3223 4475 3227
rect 4479 3223 4480 3227
rect 4474 3222 4480 3223
rect 4098 3219 4104 3220
rect 4098 3215 4099 3219
rect 4103 3215 4104 3219
rect 4098 3214 4104 3215
rect 4346 3219 4352 3220
rect 4346 3215 4347 3219
rect 4351 3215 4352 3219
rect 4346 3214 4352 3215
rect 4126 3204 4132 3205
rect 4126 3200 4127 3204
rect 4131 3200 4132 3204
rect 4126 3199 4132 3200
rect 4374 3204 4380 3205
rect 4374 3200 4375 3204
rect 4379 3200 4380 3204
rect 4374 3199 4380 3200
rect 4128 3159 4130 3199
rect 4376 3159 4378 3199
rect 4127 3158 4131 3159
rect 4127 3153 4131 3154
rect 4135 3158 4139 3159
rect 4135 3153 4139 3154
rect 4359 3158 4363 3159
rect 4359 3153 4363 3154
rect 4375 3158 4379 3159
rect 4375 3153 4379 3154
rect 4136 3129 4138 3153
rect 4360 3129 4362 3153
rect 4134 3128 4140 3129
rect 4134 3124 4135 3128
rect 4139 3124 4140 3128
rect 4134 3123 4140 3124
rect 4358 3128 4364 3129
rect 4358 3124 4359 3128
rect 4363 3124 4364 3128
rect 4358 3123 4364 3124
rect 4106 3113 4112 3114
rect 4106 3109 4107 3113
rect 4111 3109 4112 3113
rect 4106 3108 4112 3109
rect 4330 3113 4336 3114
rect 4330 3109 4331 3113
rect 4335 3109 4336 3113
rect 4330 3108 4336 3109
rect 3954 3103 3960 3104
rect 3954 3099 3955 3103
rect 3959 3099 3960 3103
rect 3954 3098 3960 3099
rect 3970 3063 3976 3064
rect 3970 3059 3971 3063
rect 3975 3059 3976 3063
rect 3970 3058 3976 3059
rect 3839 3046 3843 3047
rect 3839 3041 3843 3042
rect 3875 3046 3879 3047
rect 3875 3041 3879 3042
rect 3907 3046 3911 3047
rect 3907 3041 3911 3042
rect 3798 3032 3804 3033
rect 3466 3031 3472 3032
rect 3466 3027 3467 3031
rect 3471 3027 3472 3031
rect 3798 3028 3799 3032
rect 3803 3028 3804 3032
rect 3798 3027 3804 3028
rect 3466 3026 3472 3027
rect 3494 3016 3500 3017
rect 3494 3012 3495 3016
rect 3499 3012 3500 3016
rect 3494 3011 3500 3012
rect 3798 3015 3804 3016
rect 3798 3011 3799 3015
rect 3803 3011 3804 3015
rect 3496 2975 3498 3011
rect 3798 3010 3804 3011
rect 3800 2975 3802 3010
rect 3840 2981 3842 3041
rect 3838 2980 3844 2981
rect 3908 2980 3910 3041
rect 3972 2988 3974 3058
rect 4108 3047 4110 3108
rect 4234 3103 4240 3104
rect 4234 3099 4235 3103
rect 4239 3099 4240 3103
rect 4234 3098 4240 3099
rect 4202 3095 4208 3096
rect 4202 3091 4203 3095
rect 4207 3091 4208 3095
rect 4202 3090 4208 3091
rect 4204 3064 4206 3090
rect 4236 3064 4238 3098
rect 4202 3063 4208 3064
rect 4202 3059 4203 3063
rect 4207 3059 4208 3063
rect 4202 3058 4208 3059
rect 4234 3063 4240 3064
rect 4234 3059 4235 3063
rect 4239 3059 4240 3063
rect 4234 3058 4240 3059
rect 4332 3047 4334 3108
rect 4454 3103 4460 3104
rect 4454 3099 4455 3103
rect 4459 3099 4460 3103
rect 4454 3098 4460 3099
rect 4075 3046 4079 3047
rect 4075 3041 4079 3042
rect 4107 3046 4111 3047
rect 4107 3041 4111 3042
rect 4243 3046 4247 3047
rect 4243 3041 4247 3042
rect 4331 3046 4335 3047
rect 4331 3041 4335 3042
rect 4411 3046 4415 3047
rect 4411 3041 4415 3042
rect 3990 3031 3996 3032
rect 3990 3027 3991 3031
rect 3995 3027 3996 3031
rect 3990 3026 3996 3027
rect 3970 2987 3976 2988
rect 3970 2983 3971 2987
rect 3975 2983 3976 2987
rect 3970 2982 3976 2983
rect 3838 2976 3839 2980
rect 3843 2976 3844 2980
rect 3838 2975 3844 2976
rect 3906 2979 3912 2980
rect 3906 2975 3907 2979
rect 3911 2975 3912 2979
rect 3495 2974 3499 2975
rect 3495 2969 3499 2970
rect 3799 2974 3803 2975
rect 3906 2974 3912 2975
rect 3799 2969 3803 2970
rect 3800 2946 3802 2969
rect 3934 2964 3940 2965
rect 3838 2963 3844 2964
rect 3838 2959 3839 2963
rect 3843 2959 3844 2963
rect 3934 2960 3935 2964
rect 3939 2960 3940 2964
rect 3934 2959 3940 2960
rect 3838 2958 3844 2959
rect 3798 2945 3804 2946
rect 3798 2941 3799 2945
rect 3803 2941 3804 2945
rect 3798 2940 3804 2941
rect 3840 2931 3842 2958
rect 3936 2931 3938 2959
rect 3839 2930 3843 2931
rect 3798 2928 3804 2929
rect 3798 2924 3799 2928
rect 3803 2924 3804 2928
rect 3839 2925 3843 2926
rect 3895 2930 3899 2931
rect 3895 2925 3899 2926
rect 3935 2930 3939 2931
rect 3935 2925 3939 2926
rect 3798 2923 3804 2924
rect 3358 2879 3364 2880
rect 3358 2875 3359 2879
rect 3363 2875 3364 2879
rect 3358 2874 3364 2875
rect 3800 2855 3802 2923
rect 3840 2902 3842 2925
rect 3838 2901 3844 2902
rect 3896 2901 3898 2925
rect 3838 2897 3839 2901
rect 3843 2897 3844 2901
rect 3838 2896 3844 2897
rect 3894 2900 3900 2901
rect 3894 2896 3895 2900
rect 3899 2896 3900 2900
rect 3894 2895 3900 2896
rect 3866 2885 3872 2886
rect 3838 2884 3844 2885
rect 3838 2880 3839 2884
rect 3843 2880 3844 2884
rect 3866 2881 3867 2885
rect 3871 2881 3872 2885
rect 3866 2880 3872 2881
rect 3838 2879 3844 2880
rect 3107 2854 3111 2855
rect 3107 2849 3111 2850
rect 3307 2854 3311 2855
rect 3307 2849 3311 2850
rect 3799 2854 3803 2855
rect 3799 2849 3803 2850
rect 3030 2839 3036 2840
rect 3030 2835 3031 2839
rect 3035 2835 3036 2839
rect 3030 2834 3036 2835
rect 3800 2789 3802 2849
rect 3840 2811 3842 2879
rect 3868 2811 3870 2880
rect 3992 2876 3994 3026
rect 4076 2980 4078 3041
rect 4244 2980 4246 3041
rect 4250 3027 4256 3028
rect 4250 3023 4251 3027
rect 4255 3023 4256 3027
rect 4250 3022 4256 3023
rect 4252 2988 4254 3022
rect 4250 2987 4256 2988
rect 4250 2983 4251 2987
rect 4255 2983 4256 2987
rect 4250 2982 4256 2983
rect 4366 2987 4372 2988
rect 4366 2983 4367 2987
rect 4371 2983 4372 2987
rect 4366 2982 4372 2983
rect 4074 2979 4080 2980
rect 4074 2975 4075 2979
rect 4079 2975 4080 2979
rect 4074 2974 4080 2975
rect 4242 2979 4248 2980
rect 4242 2975 4243 2979
rect 4247 2975 4248 2979
rect 4242 2974 4248 2975
rect 4102 2964 4108 2965
rect 4102 2960 4103 2964
rect 4107 2960 4108 2964
rect 4102 2959 4108 2960
rect 4270 2964 4276 2965
rect 4270 2960 4271 2964
rect 4275 2960 4276 2964
rect 4270 2959 4276 2960
rect 4104 2931 4106 2959
rect 4272 2931 4274 2959
rect 4031 2930 4035 2931
rect 4031 2925 4035 2926
rect 4103 2930 4107 2931
rect 4103 2925 4107 2926
rect 4167 2930 4171 2931
rect 4167 2925 4171 2926
rect 4271 2930 4275 2931
rect 4271 2925 4275 2926
rect 4303 2930 4307 2931
rect 4303 2925 4307 2926
rect 4032 2901 4034 2925
rect 4168 2901 4170 2925
rect 4304 2901 4306 2925
rect 4030 2900 4036 2901
rect 4030 2896 4031 2900
rect 4035 2896 4036 2900
rect 4030 2895 4036 2896
rect 4166 2900 4172 2901
rect 4166 2896 4167 2900
rect 4171 2896 4172 2900
rect 4166 2895 4172 2896
rect 4302 2900 4308 2901
rect 4302 2896 4303 2900
rect 4307 2896 4308 2900
rect 4302 2895 4308 2896
rect 4002 2885 4008 2886
rect 4002 2881 4003 2885
rect 4007 2881 4008 2885
rect 4002 2880 4008 2881
rect 4138 2885 4144 2886
rect 4138 2881 4139 2885
rect 4143 2881 4144 2885
rect 4138 2880 4144 2881
rect 4274 2885 4280 2886
rect 4274 2881 4275 2885
rect 4279 2881 4280 2885
rect 4274 2880 4280 2881
rect 3990 2875 3996 2876
rect 3990 2871 3991 2875
rect 3995 2871 3996 2875
rect 3990 2870 3996 2871
rect 3962 2835 3968 2836
rect 3962 2831 3963 2835
rect 3967 2831 3968 2835
rect 3962 2830 3968 2831
rect 3839 2810 3843 2811
rect 3839 2805 3843 2806
rect 3859 2810 3863 2811
rect 3859 2805 3863 2806
rect 3867 2810 3871 2811
rect 3867 2805 3871 2806
rect 3798 2788 3804 2789
rect 3002 2787 3008 2788
rect 3002 2783 3003 2787
rect 3007 2783 3008 2787
rect 3798 2784 3799 2788
rect 3803 2784 3804 2788
rect 3798 2783 3804 2784
rect 3002 2782 3008 2783
rect 3030 2772 3036 2773
rect 3030 2768 3031 2772
rect 3035 2768 3036 2772
rect 3030 2767 3036 2768
rect 3798 2771 3804 2772
rect 3798 2767 3799 2771
rect 3803 2767 3804 2771
rect 3032 2739 3034 2767
rect 3798 2766 3804 2767
rect 3800 2739 3802 2766
rect 3840 2745 3842 2805
rect 3838 2744 3844 2745
rect 3860 2744 3862 2805
rect 3964 2752 3966 2830
rect 4004 2811 4006 2880
rect 4122 2875 4128 2876
rect 4122 2871 4123 2875
rect 4127 2871 4128 2875
rect 4122 2870 4128 2871
rect 3995 2810 3999 2811
rect 3995 2805 3999 2806
rect 4003 2810 4007 2811
rect 4003 2805 4007 2806
rect 3962 2751 3968 2752
rect 3962 2747 3963 2751
rect 3967 2747 3968 2751
rect 3962 2746 3968 2747
rect 3996 2744 3998 2805
rect 4124 2796 4126 2870
rect 4140 2811 4142 2880
rect 4234 2867 4240 2868
rect 4234 2863 4235 2867
rect 4239 2863 4240 2867
rect 4234 2862 4240 2863
rect 4236 2836 4238 2862
rect 4234 2835 4240 2836
rect 4234 2831 4235 2835
rect 4239 2831 4240 2835
rect 4234 2830 4240 2831
rect 4276 2811 4278 2880
rect 4368 2836 4370 2982
rect 4412 2980 4414 3041
rect 4456 3032 4458 3098
rect 4476 3064 4478 3222
rect 4580 3220 4582 3281
rect 4788 3220 4790 3281
rect 4978 3271 4984 3272
rect 4978 3267 4979 3271
rect 4983 3267 4984 3271
rect 4978 3266 4984 3267
rect 4980 3228 4982 3266
rect 4978 3227 4984 3228
rect 4978 3223 4979 3227
rect 4983 3223 4984 3227
rect 4978 3222 4984 3223
rect 4988 3220 4990 3281
rect 5144 3272 5146 3330
rect 5240 3296 5242 3450
rect 5298 3353 5304 3354
rect 5298 3349 5299 3353
rect 5303 3349 5304 3353
rect 5298 3348 5304 3349
rect 5254 3343 5260 3344
rect 5254 3339 5255 3343
rect 5259 3339 5260 3343
rect 5254 3338 5260 3339
rect 5256 3304 5258 3338
rect 5254 3303 5260 3304
rect 5254 3299 5255 3303
rect 5259 3299 5260 3303
rect 5254 3298 5260 3299
rect 5238 3295 5244 3296
rect 5238 3291 5239 3295
rect 5243 3291 5244 3295
rect 5238 3290 5244 3291
rect 5300 3287 5302 3348
rect 5171 3286 5175 3287
rect 5171 3281 5175 3282
rect 5299 3286 5303 3287
rect 5299 3281 5303 3282
rect 5142 3271 5148 3272
rect 5142 3267 5143 3271
rect 5147 3267 5148 3271
rect 5142 3266 5148 3267
rect 5172 3220 5174 3281
rect 5320 3228 5322 3494
rect 5348 3448 5350 3509
rect 5388 3456 5390 3550
rect 5516 3515 5518 3600
rect 5610 3595 5616 3596
rect 5610 3591 5611 3595
rect 5615 3591 5616 3595
rect 5610 3590 5616 3591
rect 5515 3514 5519 3515
rect 5515 3509 5519 3510
rect 5386 3455 5392 3456
rect 5386 3451 5387 3455
rect 5391 3451 5392 3455
rect 5386 3450 5392 3451
rect 5516 3448 5518 3509
rect 5612 3500 5614 3590
rect 5628 3556 5630 3726
rect 5664 3725 5666 3785
rect 5662 3724 5668 3725
rect 5662 3720 5663 3724
rect 5667 3720 5668 3724
rect 5662 3719 5668 3720
rect 5662 3707 5668 3708
rect 5662 3703 5663 3707
rect 5667 3703 5668 3707
rect 5662 3702 5668 3703
rect 5664 3651 5666 3702
rect 5663 3650 5667 3651
rect 5663 3645 5667 3646
rect 5664 3622 5666 3645
rect 5662 3621 5668 3622
rect 5662 3617 5663 3621
rect 5667 3617 5668 3621
rect 5662 3616 5668 3617
rect 5662 3604 5668 3605
rect 5662 3600 5663 3604
rect 5667 3600 5668 3604
rect 5662 3599 5668 3600
rect 5626 3555 5632 3556
rect 5626 3551 5627 3555
rect 5631 3551 5632 3555
rect 5626 3550 5632 3551
rect 5664 3515 5666 3599
rect 5663 3514 5667 3515
rect 5663 3509 5667 3510
rect 5610 3499 5616 3500
rect 5610 3495 5611 3499
rect 5615 3495 5616 3499
rect 5610 3494 5616 3495
rect 5638 3455 5644 3456
rect 5638 3451 5639 3455
rect 5643 3451 5644 3455
rect 5638 3450 5644 3451
rect 5346 3447 5352 3448
rect 5346 3443 5347 3447
rect 5351 3443 5352 3447
rect 5346 3442 5352 3443
rect 5514 3447 5520 3448
rect 5514 3443 5515 3447
rect 5519 3443 5520 3447
rect 5514 3442 5520 3443
rect 5374 3432 5380 3433
rect 5374 3428 5375 3432
rect 5379 3428 5380 3432
rect 5374 3427 5380 3428
rect 5542 3432 5548 3433
rect 5542 3428 5543 3432
rect 5547 3428 5548 3432
rect 5542 3427 5548 3428
rect 5376 3399 5378 3427
rect 5544 3399 5546 3427
rect 5327 3398 5331 3399
rect 5327 3393 5331 3394
rect 5375 3398 5379 3399
rect 5375 3393 5379 3394
rect 5543 3398 5547 3399
rect 5543 3393 5547 3394
rect 5328 3369 5330 3393
rect 5544 3369 5546 3393
rect 5326 3368 5332 3369
rect 5326 3364 5327 3368
rect 5331 3364 5332 3368
rect 5326 3363 5332 3364
rect 5542 3368 5548 3369
rect 5542 3364 5543 3368
rect 5547 3364 5548 3368
rect 5542 3363 5548 3364
rect 5514 3353 5520 3354
rect 5514 3349 5515 3353
rect 5519 3349 5520 3353
rect 5514 3348 5520 3349
rect 5516 3287 5518 3348
rect 5610 3343 5616 3344
rect 5610 3339 5611 3343
rect 5615 3339 5616 3343
rect 5610 3338 5616 3339
rect 5355 3286 5359 3287
rect 5355 3281 5359 3282
rect 5515 3286 5519 3287
rect 5515 3281 5519 3282
rect 5346 3271 5352 3272
rect 5346 3267 5347 3271
rect 5351 3267 5352 3271
rect 5346 3266 5352 3267
rect 5348 3228 5350 3266
rect 5318 3227 5324 3228
rect 5318 3223 5319 3227
rect 5323 3223 5324 3227
rect 5318 3222 5324 3223
rect 5346 3227 5352 3228
rect 5346 3223 5347 3227
rect 5351 3223 5352 3227
rect 5346 3222 5352 3223
rect 5356 3220 5358 3281
rect 5516 3220 5518 3281
rect 5612 3272 5614 3338
rect 5640 3304 5642 3450
rect 5664 3449 5666 3509
rect 5662 3448 5668 3449
rect 5662 3444 5663 3448
rect 5667 3444 5668 3448
rect 5662 3443 5668 3444
rect 5662 3431 5668 3432
rect 5662 3427 5663 3431
rect 5667 3427 5668 3431
rect 5662 3426 5668 3427
rect 5664 3399 5666 3426
rect 5663 3398 5667 3399
rect 5663 3393 5667 3394
rect 5664 3370 5666 3393
rect 5662 3369 5668 3370
rect 5662 3365 5663 3369
rect 5667 3365 5668 3369
rect 5662 3364 5668 3365
rect 5662 3352 5668 3353
rect 5662 3348 5663 3352
rect 5667 3348 5668 3352
rect 5662 3347 5668 3348
rect 5638 3303 5644 3304
rect 5638 3299 5639 3303
rect 5643 3299 5644 3303
rect 5638 3298 5644 3299
rect 5664 3287 5666 3347
rect 5663 3286 5667 3287
rect 5663 3281 5667 3282
rect 5610 3271 5616 3272
rect 5610 3267 5611 3271
rect 5615 3267 5616 3271
rect 5610 3266 5616 3267
rect 5664 3221 5666 3281
rect 5662 3220 5668 3221
rect 4578 3219 4584 3220
rect 4578 3215 4579 3219
rect 4583 3215 4584 3219
rect 4578 3214 4584 3215
rect 4786 3219 4792 3220
rect 4786 3215 4787 3219
rect 4791 3215 4792 3219
rect 4786 3214 4792 3215
rect 4986 3219 4992 3220
rect 4986 3215 4987 3219
rect 4991 3215 4992 3219
rect 4986 3214 4992 3215
rect 5170 3219 5176 3220
rect 5170 3215 5171 3219
rect 5175 3215 5176 3219
rect 5170 3214 5176 3215
rect 5354 3219 5360 3220
rect 5354 3215 5355 3219
rect 5359 3215 5360 3219
rect 5354 3214 5360 3215
rect 5514 3219 5520 3220
rect 5514 3215 5515 3219
rect 5519 3215 5520 3219
rect 5662 3216 5663 3220
rect 5667 3216 5668 3220
rect 5662 3215 5668 3216
rect 5514 3214 5520 3215
rect 4606 3204 4612 3205
rect 4606 3200 4607 3204
rect 4611 3200 4612 3204
rect 4606 3199 4612 3200
rect 4814 3204 4820 3205
rect 4814 3200 4815 3204
rect 4819 3200 4820 3204
rect 4814 3199 4820 3200
rect 5014 3204 5020 3205
rect 5014 3200 5015 3204
rect 5019 3200 5020 3204
rect 5014 3199 5020 3200
rect 5198 3204 5204 3205
rect 5198 3200 5199 3204
rect 5203 3200 5204 3204
rect 5198 3199 5204 3200
rect 5382 3204 5388 3205
rect 5382 3200 5383 3204
rect 5387 3200 5388 3204
rect 5382 3199 5388 3200
rect 5542 3204 5548 3205
rect 5542 3200 5543 3204
rect 5547 3200 5548 3204
rect 5542 3199 5548 3200
rect 5662 3203 5668 3204
rect 5662 3199 5663 3203
rect 5667 3199 5668 3203
rect 4608 3159 4610 3199
rect 4816 3159 4818 3199
rect 5016 3159 5018 3199
rect 5200 3159 5202 3199
rect 5384 3159 5386 3199
rect 5544 3159 5546 3199
rect 5662 3198 5668 3199
rect 5664 3159 5666 3198
rect 4583 3158 4587 3159
rect 4583 3153 4587 3154
rect 4607 3158 4611 3159
rect 4607 3153 4611 3154
rect 4807 3158 4811 3159
rect 4807 3153 4811 3154
rect 4815 3158 4819 3159
rect 4815 3153 4819 3154
rect 5015 3158 5019 3159
rect 5015 3153 5019 3154
rect 5031 3158 5035 3159
rect 5031 3153 5035 3154
rect 5199 3158 5203 3159
rect 5199 3153 5203 3154
rect 5383 3158 5387 3159
rect 5383 3153 5387 3154
rect 5543 3158 5547 3159
rect 5543 3153 5547 3154
rect 5663 3158 5667 3159
rect 5663 3153 5667 3154
rect 4584 3129 4586 3153
rect 4808 3129 4810 3153
rect 5032 3129 5034 3153
rect 5664 3130 5666 3153
rect 5662 3129 5668 3130
rect 4582 3128 4588 3129
rect 4582 3124 4583 3128
rect 4587 3124 4588 3128
rect 4582 3123 4588 3124
rect 4806 3128 4812 3129
rect 4806 3124 4807 3128
rect 4811 3124 4812 3128
rect 4806 3123 4812 3124
rect 5030 3128 5036 3129
rect 5030 3124 5031 3128
rect 5035 3124 5036 3128
rect 5662 3125 5663 3129
rect 5667 3125 5668 3129
rect 5662 3124 5668 3125
rect 5030 3123 5036 3124
rect 4554 3113 4560 3114
rect 4554 3109 4555 3113
rect 4559 3109 4560 3113
rect 4554 3108 4560 3109
rect 4778 3113 4784 3114
rect 4778 3109 4779 3113
rect 4783 3109 4784 3113
rect 4778 3108 4784 3109
rect 5002 3113 5008 3114
rect 5002 3109 5003 3113
rect 5007 3109 5008 3113
rect 5002 3108 5008 3109
rect 5662 3112 5668 3113
rect 5662 3108 5663 3112
rect 5667 3108 5668 3112
rect 4474 3063 4480 3064
rect 4474 3059 4475 3063
rect 4479 3059 4480 3063
rect 4474 3058 4480 3059
rect 4556 3047 4558 3108
rect 4682 3103 4688 3104
rect 4682 3099 4683 3103
rect 4687 3099 4688 3103
rect 4682 3098 4688 3099
rect 4684 3064 4686 3098
rect 4682 3063 4688 3064
rect 4682 3059 4683 3063
rect 4687 3059 4688 3063
rect 4682 3058 4688 3059
rect 4780 3047 4782 3108
rect 4906 3103 4912 3104
rect 4906 3099 4907 3103
rect 4911 3099 4912 3103
rect 4906 3098 4912 3099
rect 4908 3064 4910 3098
rect 4906 3063 4912 3064
rect 4906 3059 4907 3063
rect 4911 3059 4912 3063
rect 4906 3058 4912 3059
rect 5004 3047 5006 3108
rect 5662 3107 5668 3108
rect 5664 3047 5666 3107
rect 4555 3046 4559 3047
rect 4555 3041 4559 3042
rect 4579 3046 4583 3047
rect 4579 3041 4583 3042
rect 4755 3046 4759 3047
rect 4755 3041 4759 3042
rect 4779 3046 4783 3047
rect 4779 3041 4783 3042
rect 5003 3046 5007 3047
rect 5003 3041 5007 3042
rect 5663 3046 5667 3047
rect 5663 3041 5667 3042
rect 4454 3031 4460 3032
rect 4454 3027 4455 3031
rect 4459 3027 4460 3031
rect 4454 3026 4460 3027
rect 4580 2980 4582 3041
rect 4586 3027 4592 3028
rect 4586 3023 4587 3027
rect 4591 3023 4592 3027
rect 4586 3022 4592 3023
rect 4588 2988 4590 3022
rect 4586 2987 4592 2988
rect 4586 2983 4587 2987
rect 4591 2983 4592 2987
rect 4586 2982 4592 2983
rect 4756 2980 4758 3041
rect 4878 3039 4884 3040
rect 4878 3035 4879 3039
rect 4883 3035 4884 3039
rect 4878 3034 4884 3035
rect 4762 3027 4768 3028
rect 4762 3023 4763 3027
rect 4767 3023 4768 3027
rect 4762 3022 4768 3023
rect 4764 2988 4766 3022
rect 4880 2988 4882 3034
rect 4762 2987 4768 2988
rect 4762 2983 4763 2987
rect 4767 2983 4768 2987
rect 4762 2982 4768 2983
rect 4878 2987 4884 2988
rect 4878 2983 4879 2987
rect 4883 2983 4884 2987
rect 4878 2982 4884 2983
rect 5664 2981 5666 3041
rect 5662 2980 5668 2981
rect 4410 2979 4416 2980
rect 4410 2975 4411 2979
rect 4415 2975 4416 2979
rect 4410 2974 4416 2975
rect 4578 2979 4584 2980
rect 4578 2975 4579 2979
rect 4583 2975 4584 2979
rect 4578 2974 4584 2975
rect 4754 2979 4760 2980
rect 4754 2975 4755 2979
rect 4759 2975 4760 2979
rect 5662 2976 5663 2980
rect 5667 2976 5668 2980
rect 5662 2975 5668 2976
rect 4754 2974 4760 2975
rect 4438 2964 4444 2965
rect 4438 2960 4439 2964
rect 4443 2960 4444 2964
rect 4438 2959 4444 2960
rect 4606 2964 4612 2965
rect 4606 2960 4607 2964
rect 4611 2960 4612 2964
rect 4606 2959 4612 2960
rect 4782 2964 4788 2965
rect 4782 2960 4783 2964
rect 4787 2960 4788 2964
rect 4782 2959 4788 2960
rect 5662 2963 5668 2964
rect 5662 2959 5663 2963
rect 5667 2959 5668 2963
rect 4440 2931 4442 2959
rect 4608 2931 4610 2959
rect 4784 2931 4786 2959
rect 5662 2958 5668 2959
rect 5664 2931 5666 2958
rect 4439 2930 4443 2931
rect 4439 2925 4443 2926
rect 4575 2930 4579 2931
rect 4575 2925 4579 2926
rect 4607 2930 4611 2931
rect 4607 2925 4611 2926
rect 4783 2930 4787 2931
rect 4783 2925 4787 2926
rect 5663 2930 5667 2931
rect 5663 2925 5667 2926
rect 4440 2901 4442 2925
rect 4576 2901 4578 2925
rect 5664 2902 5666 2925
rect 5662 2901 5668 2902
rect 4438 2900 4444 2901
rect 4438 2896 4439 2900
rect 4443 2896 4444 2900
rect 4438 2895 4444 2896
rect 4574 2900 4580 2901
rect 4574 2896 4575 2900
rect 4579 2896 4580 2900
rect 5662 2897 5663 2901
rect 5667 2897 5668 2901
rect 5662 2896 5668 2897
rect 4574 2895 4580 2896
rect 4410 2885 4416 2886
rect 4410 2881 4411 2885
rect 4415 2881 4416 2885
rect 4410 2880 4416 2881
rect 4546 2885 4552 2886
rect 4546 2881 4547 2885
rect 4551 2881 4552 2885
rect 4546 2880 4552 2881
rect 5662 2884 5668 2885
rect 5662 2880 5663 2884
rect 5667 2880 5668 2884
rect 4402 2875 4408 2876
rect 4402 2871 4403 2875
rect 4407 2871 4408 2875
rect 4402 2870 4408 2871
rect 4404 2836 4406 2870
rect 4366 2835 4372 2836
rect 4366 2831 4367 2835
rect 4371 2831 4372 2835
rect 4366 2830 4372 2831
rect 4402 2835 4408 2836
rect 4402 2831 4403 2835
rect 4407 2831 4408 2835
rect 4402 2830 4408 2831
rect 4412 2811 4414 2880
rect 4538 2875 4544 2876
rect 4538 2871 4539 2875
rect 4543 2871 4544 2875
rect 4538 2870 4544 2871
rect 4540 2836 4542 2870
rect 4538 2835 4544 2836
rect 4538 2831 4539 2835
rect 4543 2831 4544 2835
rect 4538 2830 4544 2831
rect 4548 2811 4550 2880
rect 5662 2879 5668 2880
rect 5664 2811 5666 2879
rect 4131 2810 4135 2811
rect 4131 2805 4135 2806
rect 4139 2810 4143 2811
rect 4139 2805 4143 2806
rect 4267 2810 4271 2811
rect 4267 2805 4271 2806
rect 4275 2810 4279 2811
rect 4275 2805 4279 2806
rect 4403 2810 4407 2811
rect 4403 2805 4407 2806
rect 4411 2810 4415 2811
rect 4411 2805 4415 2806
rect 4539 2810 4543 2811
rect 4539 2805 4543 2806
rect 4547 2810 4551 2811
rect 4547 2805 4551 2806
rect 4675 2810 4679 2811
rect 4675 2805 4679 2806
rect 4811 2810 4815 2811
rect 4811 2805 4815 2806
rect 5663 2810 5667 2811
rect 5663 2805 5667 2806
rect 4054 2795 4060 2796
rect 4054 2791 4055 2795
rect 4059 2791 4060 2795
rect 4054 2790 4060 2791
rect 4122 2795 4128 2796
rect 4122 2791 4123 2795
rect 4127 2791 4128 2795
rect 4122 2790 4128 2791
rect 3838 2740 3839 2744
rect 3843 2740 3844 2744
rect 3838 2739 3844 2740
rect 3858 2743 3864 2744
rect 3858 2739 3859 2743
rect 3863 2739 3864 2743
rect 3015 2738 3019 2739
rect 3015 2733 3019 2734
rect 3031 2738 3035 2739
rect 3031 2733 3035 2734
rect 3799 2738 3803 2739
rect 3858 2738 3864 2739
rect 3994 2743 4000 2744
rect 3994 2739 3995 2743
rect 3999 2739 4000 2743
rect 3994 2738 4000 2739
rect 3799 2733 3803 2734
rect 3016 2709 3018 2733
rect 3800 2710 3802 2733
rect 3886 2728 3892 2729
rect 3838 2727 3844 2728
rect 3838 2723 3839 2727
rect 3843 2723 3844 2727
rect 3886 2724 3887 2728
rect 3891 2724 3892 2728
rect 3886 2723 3892 2724
rect 4022 2728 4028 2729
rect 4022 2724 4023 2728
rect 4027 2724 4028 2728
rect 4022 2723 4028 2724
rect 3838 2722 3844 2723
rect 3798 2709 3804 2710
rect 3014 2708 3020 2709
rect 3014 2704 3015 2708
rect 3019 2704 3020 2708
rect 3798 2705 3799 2709
rect 3803 2705 3804 2709
rect 3798 2704 3804 2705
rect 3014 2703 3020 2704
rect 3840 2699 3842 2722
rect 3888 2699 3890 2723
rect 4024 2699 4026 2723
rect 3839 2698 3843 2699
rect 2986 2693 2992 2694
rect 3839 2693 3843 2694
rect 3887 2698 3891 2699
rect 3887 2693 3891 2694
rect 3959 2698 3963 2699
rect 3959 2693 3963 2694
rect 4023 2698 4027 2699
rect 4023 2693 4027 2694
rect 2986 2689 2987 2693
rect 2991 2689 2992 2693
rect 2986 2688 2992 2689
rect 3798 2692 3804 2693
rect 3798 2688 3799 2692
rect 3803 2688 3804 2692
rect 2858 2683 2864 2684
rect 2858 2679 2859 2683
rect 2863 2679 2864 2683
rect 2858 2678 2864 2679
rect 2860 2644 2862 2678
rect 2858 2643 2864 2644
rect 2858 2639 2859 2643
rect 2863 2639 2864 2643
rect 2858 2638 2864 2639
rect 2806 2635 2812 2636
rect 2806 2631 2807 2635
rect 2811 2631 2812 2635
rect 2806 2630 2812 2631
rect 2988 2615 2990 2688
rect 3798 2687 3804 2688
rect 3110 2683 3116 2684
rect 3110 2679 3111 2683
rect 3115 2679 3116 2683
rect 3110 2678 3116 2679
rect 2555 2614 2559 2615
rect 2555 2609 2559 2610
rect 2691 2614 2695 2615
rect 2691 2609 2695 2610
rect 2731 2614 2735 2615
rect 2731 2609 2735 2610
rect 2827 2614 2831 2615
rect 2827 2609 2831 2610
rect 2963 2614 2967 2615
rect 2963 2609 2967 2610
rect 2987 2614 2991 2615
rect 2987 2609 2991 2610
rect 3099 2614 3103 2615
rect 3099 2609 3103 2610
rect 2538 2555 2544 2556
rect 2538 2551 2539 2555
rect 2543 2551 2544 2555
rect 2538 2550 2544 2551
rect 1974 2548 1980 2549
rect 2556 2548 2558 2609
rect 2692 2548 2694 2609
rect 2774 2599 2780 2600
rect 2774 2595 2775 2599
rect 2779 2595 2780 2599
rect 2774 2594 2780 2595
rect 1974 2544 1975 2548
rect 1979 2544 1980 2548
rect 1974 2543 1980 2544
rect 2554 2547 2560 2548
rect 2554 2543 2555 2547
rect 2559 2543 2560 2547
rect 2554 2542 2560 2543
rect 2690 2547 2696 2548
rect 2690 2543 2691 2547
rect 2695 2543 2696 2547
rect 2690 2542 2696 2543
rect 1543 2538 1547 2539
rect 1543 2533 1547 2534
rect 1631 2538 1635 2539
rect 1631 2533 1635 2534
rect 1703 2538 1707 2539
rect 1703 2533 1707 2534
rect 1815 2538 1819 2539
rect 1815 2533 1819 2534
rect 1935 2538 1939 2539
rect 1935 2533 1939 2534
rect 1632 2509 1634 2533
rect 1816 2509 1818 2533
rect 1936 2510 1938 2533
rect 2582 2532 2588 2533
rect 1974 2531 1980 2532
rect 1974 2527 1975 2531
rect 1979 2527 1980 2531
rect 2582 2528 2583 2532
rect 2587 2528 2588 2532
rect 2582 2527 2588 2528
rect 2718 2532 2724 2533
rect 2718 2528 2719 2532
rect 2723 2528 2724 2532
rect 2718 2527 2724 2528
rect 1974 2526 1980 2527
rect 1934 2509 1940 2510
rect 1630 2508 1636 2509
rect 1630 2504 1631 2508
rect 1635 2504 1636 2508
rect 1630 2503 1636 2504
rect 1814 2508 1820 2509
rect 1814 2504 1815 2508
rect 1819 2504 1820 2508
rect 1934 2505 1935 2509
rect 1939 2505 1940 2509
rect 1934 2504 1940 2505
rect 1814 2503 1820 2504
rect 1602 2493 1608 2494
rect 1602 2489 1603 2493
rect 1607 2489 1608 2493
rect 1602 2488 1608 2489
rect 1786 2493 1792 2494
rect 1786 2489 1787 2493
rect 1791 2489 1792 2493
rect 1786 2488 1792 2489
rect 1934 2492 1940 2493
rect 1934 2488 1935 2492
rect 1939 2488 1940 2492
rect 1562 2483 1568 2484
rect 1562 2479 1563 2483
rect 1567 2479 1568 2483
rect 1562 2478 1568 2479
rect 1564 2444 1566 2478
rect 1498 2443 1504 2444
rect 1498 2439 1499 2443
rect 1503 2439 1504 2443
rect 1498 2438 1504 2439
rect 1562 2443 1568 2444
rect 1562 2439 1563 2443
rect 1567 2439 1568 2443
rect 1562 2438 1568 2439
rect 1604 2423 1606 2488
rect 1730 2483 1736 2484
rect 1730 2479 1731 2483
rect 1735 2479 1736 2483
rect 1730 2478 1736 2479
rect 1732 2444 1734 2478
rect 1730 2443 1736 2444
rect 1730 2439 1731 2443
rect 1735 2439 1736 2443
rect 1730 2438 1736 2439
rect 1788 2423 1790 2488
rect 1934 2487 1940 2488
rect 1882 2483 1888 2484
rect 1882 2479 1883 2483
rect 1887 2479 1888 2483
rect 1882 2478 1888 2479
rect 523 2422 527 2423
rect 523 2417 527 2418
rect 571 2422 575 2423
rect 571 2417 575 2418
rect 787 2422 791 2423
rect 787 2417 791 2418
rect 835 2422 839 2423
rect 835 2417 839 2418
rect 995 2422 999 2423
rect 995 2417 999 2418
rect 1155 2422 1159 2423
rect 1155 2417 1159 2418
rect 1203 2422 1207 2423
rect 1203 2417 1207 2418
rect 1403 2422 1407 2423
rect 1403 2417 1407 2418
rect 1483 2422 1487 2423
rect 1483 2417 1487 2418
rect 1603 2422 1607 2423
rect 1603 2417 1607 2418
rect 1787 2422 1791 2423
rect 1787 2417 1791 2418
rect 454 2407 460 2408
rect 454 2403 455 2407
rect 459 2403 460 2407
rect 454 2402 460 2403
rect 456 2364 458 2402
rect 362 2363 368 2364
rect 362 2359 363 2363
rect 367 2359 368 2363
rect 362 2358 368 2359
rect 454 2363 460 2364
rect 454 2359 455 2363
rect 459 2359 460 2363
rect 454 2358 460 2359
rect 524 2356 526 2417
rect 618 2403 624 2404
rect 618 2399 619 2403
rect 623 2399 624 2403
rect 618 2398 624 2399
rect 110 2352 111 2356
rect 115 2352 116 2356
rect 110 2351 116 2352
rect 226 2355 232 2356
rect 226 2351 227 2355
rect 231 2351 232 2355
rect 226 2350 232 2351
rect 522 2355 528 2356
rect 522 2351 523 2355
rect 527 2351 528 2355
rect 522 2350 528 2351
rect 254 2340 260 2341
rect 110 2339 116 2340
rect 110 2335 111 2339
rect 115 2335 116 2339
rect 254 2336 255 2340
rect 259 2336 260 2340
rect 254 2335 260 2336
rect 550 2340 556 2341
rect 550 2336 551 2340
rect 555 2336 556 2340
rect 550 2335 556 2336
rect 110 2334 116 2335
rect 112 2295 114 2334
rect 256 2295 258 2335
rect 552 2295 554 2335
rect 111 2294 115 2295
rect 111 2289 115 2290
rect 159 2294 163 2295
rect 159 2289 163 2290
rect 255 2294 259 2295
rect 255 2289 259 2290
rect 367 2294 371 2295
rect 367 2289 371 2290
rect 551 2294 555 2295
rect 551 2289 555 2290
rect 599 2294 603 2295
rect 599 2289 603 2290
rect 112 2266 114 2289
rect 110 2265 116 2266
rect 160 2265 162 2289
rect 368 2265 370 2289
rect 600 2265 602 2289
rect 110 2261 111 2265
rect 115 2261 116 2265
rect 110 2260 116 2261
rect 158 2264 164 2265
rect 158 2260 159 2264
rect 163 2260 164 2264
rect 158 2259 164 2260
rect 366 2264 372 2265
rect 366 2260 367 2264
rect 371 2260 372 2264
rect 366 2259 372 2260
rect 598 2264 604 2265
rect 598 2260 599 2264
rect 603 2260 604 2264
rect 598 2259 604 2260
rect 130 2249 136 2250
rect 110 2248 116 2249
rect 110 2244 111 2248
rect 115 2244 116 2248
rect 130 2245 131 2249
rect 135 2245 136 2249
rect 130 2244 136 2245
rect 338 2249 344 2250
rect 338 2245 339 2249
rect 343 2245 344 2249
rect 338 2244 344 2245
rect 570 2249 576 2250
rect 570 2245 571 2249
rect 575 2245 576 2249
rect 570 2244 576 2245
rect 110 2243 116 2244
rect 112 2171 114 2243
rect 132 2171 134 2244
rect 278 2239 284 2240
rect 278 2235 279 2239
rect 283 2235 284 2239
rect 278 2234 284 2235
rect 280 2200 282 2234
rect 226 2199 232 2200
rect 226 2195 227 2199
rect 231 2195 232 2199
rect 226 2194 232 2195
rect 278 2199 284 2200
rect 278 2195 279 2199
rect 283 2195 284 2199
rect 278 2194 284 2195
rect 111 2170 115 2171
rect 111 2165 115 2166
rect 131 2170 135 2171
rect 131 2165 135 2166
rect 112 2105 114 2165
rect 110 2104 116 2105
rect 132 2104 134 2165
rect 228 2112 230 2194
rect 340 2171 342 2244
rect 466 2239 472 2240
rect 466 2235 467 2239
rect 471 2235 472 2239
rect 466 2234 472 2235
rect 468 2200 470 2234
rect 466 2199 472 2200
rect 466 2195 467 2199
rect 471 2195 472 2199
rect 466 2194 472 2195
rect 572 2171 574 2244
rect 620 2240 622 2398
rect 836 2356 838 2417
rect 898 2363 904 2364
rect 898 2359 899 2363
rect 903 2359 904 2363
rect 898 2358 904 2359
rect 834 2355 840 2356
rect 834 2351 835 2355
rect 839 2351 840 2355
rect 834 2350 840 2351
rect 862 2340 868 2341
rect 862 2336 863 2340
rect 867 2336 868 2340
rect 862 2335 868 2336
rect 864 2295 866 2335
rect 831 2294 835 2295
rect 831 2289 835 2290
rect 863 2294 867 2295
rect 863 2289 867 2290
rect 832 2265 834 2289
rect 830 2264 836 2265
rect 830 2260 831 2264
rect 835 2260 836 2264
rect 830 2259 836 2260
rect 802 2249 808 2250
rect 802 2245 803 2249
rect 807 2245 808 2249
rect 802 2244 808 2245
rect 618 2239 624 2240
rect 618 2235 619 2239
rect 623 2235 624 2239
rect 618 2234 624 2235
rect 804 2171 806 2244
rect 900 2200 902 2358
rect 1156 2356 1158 2417
rect 1278 2415 1284 2416
rect 1278 2411 1279 2415
rect 1283 2411 1284 2415
rect 1278 2410 1284 2411
rect 1280 2364 1282 2410
rect 1278 2363 1284 2364
rect 1278 2359 1279 2363
rect 1283 2359 1284 2363
rect 1278 2358 1284 2359
rect 1484 2356 1486 2417
rect 1594 2415 1600 2416
rect 1594 2411 1595 2415
rect 1599 2411 1600 2415
rect 1594 2410 1600 2411
rect 1596 2364 1598 2410
rect 1594 2363 1600 2364
rect 1594 2359 1595 2363
rect 1599 2359 1600 2363
rect 1594 2358 1600 2359
rect 1788 2356 1790 2417
rect 1884 2408 1886 2478
rect 1936 2423 1938 2487
rect 1976 2479 1978 2526
rect 2584 2479 2586 2527
rect 2720 2479 2722 2527
rect 1975 2478 1979 2479
rect 1975 2473 1979 2474
rect 2023 2478 2027 2479
rect 2023 2473 2027 2474
rect 2223 2478 2227 2479
rect 2223 2473 2227 2474
rect 2447 2478 2451 2479
rect 2447 2473 2451 2474
rect 2583 2478 2587 2479
rect 2583 2473 2587 2474
rect 2679 2478 2683 2479
rect 2679 2473 2683 2474
rect 2719 2478 2723 2479
rect 2719 2473 2723 2474
rect 1976 2450 1978 2473
rect 1974 2449 1980 2450
rect 2024 2449 2026 2473
rect 2224 2449 2226 2473
rect 2448 2449 2450 2473
rect 2680 2449 2682 2473
rect 1974 2445 1975 2449
rect 1979 2445 1980 2449
rect 1974 2444 1980 2445
rect 2022 2448 2028 2449
rect 2022 2444 2023 2448
rect 2027 2444 2028 2448
rect 2022 2443 2028 2444
rect 2222 2448 2228 2449
rect 2222 2444 2223 2448
rect 2227 2444 2228 2448
rect 2222 2443 2228 2444
rect 2446 2448 2452 2449
rect 2446 2444 2447 2448
rect 2451 2444 2452 2448
rect 2446 2443 2452 2444
rect 2678 2448 2684 2449
rect 2678 2444 2679 2448
rect 2683 2444 2684 2448
rect 2678 2443 2684 2444
rect 1994 2433 2000 2434
rect 1974 2432 1980 2433
rect 1974 2428 1975 2432
rect 1979 2428 1980 2432
rect 1994 2429 1995 2433
rect 1999 2429 2000 2433
rect 1994 2428 2000 2429
rect 2194 2433 2200 2434
rect 2194 2429 2195 2433
rect 2199 2429 2200 2433
rect 2194 2428 2200 2429
rect 2418 2433 2424 2434
rect 2418 2429 2419 2433
rect 2423 2429 2424 2433
rect 2418 2428 2424 2429
rect 2650 2433 2656 2434
rect 2650 2429 2651 2433
rect 2655 2429 2656 2433
rect 2650 2428 2656 2429
rect 1974 2427 1980 2428
rect 1935 2422 1939 2423
rect 1935 2417 1939 2418
rect 1882 2407 1888 2408
rect 1882 2403 1883 2407
rect 1887 2403 1888 2407
rect 1882 2402 1888 2403
rect 1936 2357 1938 2417
rect 1976 2359 1978 2427
rect 1996 2359 1998 2428
rect 2090 2423 2096 2424
rect 2090 2419 2091 2423
rect 2095 2419 2096 2423
rect 2090 2418 2096 2419
rect 1975 2358 1979 2359
rect 1934 2356 1940 2357
rect 1154 2355 1160 2356
rect 1154 2351 1155 2355
rect 1159 2351 1160 2355
rect 1154 2350 1160 2351
rect 1482 2355 1488 2356
rect 1482 2351 1483 2355
rect 1487 2351 1488 2355
rect 1482 2350 1488 2351
rect 1786 2355 1792 2356
rect 1786 2351 1787 2355
rect 1791 2351 1792 2355
rect 1934 2352 1935 2356
rect 1939 2352 1940 2356
rect 1975 2353 1979 2354
rect 1995 2358 1999 2359
rect 1995 2353 1999 2354
rect 1934 2351 1940 2352
rect 1786 2350 1792 2351
rect 1182 2340 1188 2341
rect 1182 2336 1183 2340
rect 1187 2336 1188 2340
rect 1182 2335 1188 2336
rect 1510 2340 1516 2341
rect 1510 2336 1511 2340
rect 1515 2336 1516 2340
rect 1510 2335 1516 2336
rect 1814 2340 1820 2341
rect 1814 2336 1815 2340
rect 1819 2336 1820 2340
rect 1814 2335 1820 2336
rect 1934 2339 1940 2340
rect 1934 2335 1935 2339
rect 1939 2335 1940 2339
rect 1184 2295 1186 2335
rect 1512 2295 1514 2335
rect 1816 2295 1818 2335
rect 1934 2334 1940 2335
rect 1936 2295 1938 2334
rect 1063 2294 1067 2295
rect 1063 2289 1067 2290
rect 1183 2294 1187 2295
rect 1183 2289 1187 2290
rect 1511 2294 1515 2295
rect 1511 2289 1515 2290
rect 1815 2294 1819 2295
rect 1815 2289 1819 2290
rect 1935 2294 1939 2295
rect 1976 2293 1978 2353
rect 1935 2289 1939 2290
rect 1974 2292 1980 2293
rect 1996 2292 1998 2353
rect 2092 2344 2094 2418
rect 2196 2359 2198 2428
rect 2322 2423 2328 2424
rect 2322 2419 2323 2423
rect 2327 2419 2328 2423
rect 2322 2418 2328 2419
rect 2324 2384 2326 2418
rect 2322 2383 2328 2384
rect 2322 2379 2323 2383
rect 2327 2379 2328 2383
rect 2322 2378 2328 2379
rect 2420 2359 2422 2428
rect 2546 2423 2552 2424
rect 2546 2419 2547 2423
rect 2551 2419 2552 2423
rect 2546 2418 2552 2419
rect 2548 2384 2550 2418
rect 2546 2383 2552 2384
rect 2546 2379 2547 2383
rect 2551 2379 2552 2383
rect 2546 2378 2552 2379
rect 2546 2375 2552 2376
rect 2546 2371 2547 2375
rect 2551 2371 2552 2375
rect 2546 2370 2552 2371
rect 2155 2358 2159 2359
rect 2155 2353 2159 2354
rect 2195 2358 2199 2359
rect 2195 2353 2199 2354
rect 2347 2358 2351 2359
rect 2347 2353 2351 2354
rect 2419 2358 2423 2359
rect 2419 2353 2423 2354
rect 2539 2358 2543 2359
rect 2539 2353 2543 2354
rect 2090 2343 2096 2344
rect 2090 2339 2091 2343
rect 2095 2339 2096 2343
rect 2090 2338 2096 2339
rect 2156 2292 2158 2353
rect 2162 2339 2168 2340
rect 2162 2335 2163 2339
rect 2167 2335 2168 2339
rect 2162 2334 2168 2335
rect 2164 2300 2166 2334
rect 2162 2299 2168 2300
rect 2162 2295 2163 2299
rect 2167 2295 2168 2299
rect 2162 2294 2168 2295
rect 2348 2292 2350 2353
rect 2354 2339 2360 2340
rect 2354 2335 2355 2339
rect 2359 2335 2360 2339
rect 2354 2334 2360 2335
rect 2356 2300 2358 2334
rect 2354 2299 2360 2300
rect 2354 2295 2355 2299
rect 2359 2295 2360 2299
rect 2354 2294 2360 2295
rect 2470 2299 2476 2300
rect 2470 2295 2471 2299
rect 2475 2295 2476 2299
rect 2470 2294 2476 2295
rect 1064 2265 1066 2289
rect 1936 2266 1938 2289
rect 1974 2288 1975 2292
rect 1979 2288 1980 2292
rect 1974 2287 1980 2288
rect 1994 2291 2000 2292
rect 1994 2287 1995 2291
rect 1999 2287 2000 2291
rect 1994 2286 2000 2287
rect 2154 2291 2160 2292
rect 2154 2287 2155 2291
rect 2159 2287 2160 2291
rect 2154 2286 2160 2287
rect 2346 2291 2352 2292
rect 2346 2287 2347 2291
rect 2351 2287 2352 2291
rect 2346 2286 2352 2287
rect 2022 2276 2028 2277
rect 1974 2275 1980 2276
rect 1974 2271 1975 2275
rect 1979 2271 1980 2275
rect 2022 2272 2023 2276
rect 2027 2272 2028 2276
rect 2022 2271 2028 2272
rect 2182 2276 2188 2277
rect 2182 2272 2183 2276
rect 2187 2272 2188 2276
rect 2182 2271 2188 2272
rect 2374 2276 2380 2277
rect 2374 2272 2375 2276
rect 2379 2272 2380 2276
rect 2374 2271 2380 2272
rect 1974 2270 1980 2271
rect 1934 2265 1940 2266
rect 1062 2264 1068 2265
rect 1062 2260 1063 2264
rect 1067 2260 1068 2264
rect 1934 2261 1935 2265
rect 1939 2261 1940 2265
rect 1934 2260 1940 2261
rect 1062 2259 1068 2260
rect 1034 2249 1040 2250
rect 1034 2245 1035 2249
rect 1039 2245 1040 2249
rect 1034 2244 1040 2245
rect 1934 2248 1940 2249
rect 1934 2244 1935 2248
rect 1939 2244 1940 2248
rect 930 2239 936 2240
rect 930 2235 931 2239
rect 935 2235 936 2239
rect 930 2234 936 2235
rect 932 2200 934 2234
rect 898 2199 904 2200
rect 898 2195 899 2199
rect 903 2195 904 2199
rect 898 2194 904 2195
rect 930 2199 936 2200
rect 930 2195 931 2199
rect 935 2195 936 2199
rect 930 2194 936 2195
rect 1036 2171 1038 2244
rect 1934 2243 1940 2244
rect 1158 2239 1164 2240
rect 1158 2235 1159 2239
rect 1163 2235 1164 2239
rect 1158 2234 1164 2235
rect 339 2170 343 2171
rect 339 2165 343 2166
rect 347 2170 351 2171
rect 347 2165 351 2166
rect 571 2170 575 2171
rect 571 2165 575 2166
rect 595 2170 599 2171
rect 595 2165 599 2166
rect 803 2170 807 2171
rect 803 2165 807 2166
rect 835 2170 839 2171
rect 835 2165 839 2166
rect 1035 2170 1039 2171
rect 1035 2165 1039 2166
rect 1075 2170 1079 2171
rect 1075 2165 1079 2166
rect 338 2155 344 2156
rect 338 2151 339 2155
rect 343 2151 344 2155
rect 338 2150 344 2151
rect 340 2112 342 2150
rect 226 2111 232 2112
rect 226 2107 227 2111
rect 231 2107 232 2111
rect 226 2106 232 2107
rect 338 2111 344 2112
rect 338 2107 339 2111
rect 343 2107 344 2111
rect 338 2106 344 2107
rect 348 2104 350 2165
rect 596 2104 598 2165
rect 638 2155 644 2156
rect 638 2151 639 2155
rect 643 2151 644 2155
rect 638 2150 644 2151
rect 110 2100 111 2104
rect 115 2100 116 2104
rect 110 2099 116 2100
rect 130 2103 136 2104
rect 130 2099 131 2103
rect 135 2099 136 2103
rect 130 2098 136 2099
rect 346 2103 352 2104
rect 346 2099 347 2103
rect 351 2099 352 2103
rect 346 2098 352 2099
rect 594 2103 600 2104
rect 594 2099 595 2103
rect 599 2099 600 2103
rect 594 2098 600 2099
rect 158 2088 164 2089
rect 110 2087 116 2088
rect 110 2083 111 2087
rect 115 2083 116 2087
rect 158 2084 159 2088
rect 163 2084 164 2088
rect 158 2083 164 2084
rect 374 2088 380 2089
rect 374 2084 375 2088
rect 379 2084 380 2088
rect 374 2083 380 2084
rect 622 2088 628 2089
rect 622 2084 623 2088
rect 627 2084 628 2088
rect 622 2083 628 2084
rect 110 2082 116 2083
rect 112 2055 114 2082
rect 160 2055 162 2083
rect 376 2055 378 2083
rect 624 2055 626 2083
rect 111 2054 115 2055
rect 111 2049 115 2050
rect 159 2054 163 2055
rect 159 2049 163 2050
rect 271 2054 275 2055
rect 271 2049 275 2050
rect 375 2054 379 2055
rect 375 2049 379 2050
rect 407 2054 411 2055
rect 407 2049 411 2050
rect 543 2054 547 2055
rect 543 2049 547 2050
rect 623 2054 627 2055
rect 623 2049 627 2050
rect 112 2026 114 2049
rect 110 2025 116 2026
rect 272 2025 274 2049
rect 408 2025 410 2049
rect 544 2025 546 2049
rect 110 2021 111 2025
rect 115 2021 116 2025
rect 110 2020 116 2021
rect 270 2024 276 2025
rect 270 2020 271 2024
rect 275 2020 276 2024
rect 270 2019 276 2020
rect 406 2024 412 2025
rect 406 2020 407 2024
rect 411 2020 412 2024
rect 406 2019 412 2020
rect 542 2024 548 2025
rect 542 2020 543 2024
rect 547 2020 548 2024
rect 542 2019 548 2020
rect 242 2009 248 2010
rect 110 2008 116 2009
rect 110 2004 111 2008
rect 115 2004 116 2008
rect 242 2005 243 2009
rect 247 2005 248 2009
rect 242 2004 248 2005
rect 378 2009 384 2010
rect 378 2005 379 2009
rect 383 2005 384 2009
rect 378 2004 384 2005
rect 514 2009 520 2010
rect 514 2005 515 2009
rect 519 2005 520 2009
rect 514 2004 520 2005
rect 110 2003 116 2004
rect 112 1939 114 2003
rect 244 1939 246 2004
rect 370 1999 376 2000
rect 370 1995 371 1999
rect 375 1995 376 1999
rect 370 1994 376 1995
rect 372 1960 374 1994
rect 310 1959 316 1960
rect 310 1955 311 1959
rect 315 1955 316 1959
rect 310 1954 316 1955
rect 370 1959 376 1960
rect 370 1955 371 1959
rect 375 1955 376 1959
rect 370 1954 376 1955
rect 111 1938 115 1939
rect 111 1933 115 1934
rect 187 1938 191 1939
rect 187 1933 191 1934
rect 243 1938 247 1939
rect 243 1933 247 1934
rect 112 1873 114 1933
rect 110 1872 116 1873
rect 188 1872 190 1933
rect 312 1880 314 1954
rect 380 1939 382 2004
rect 506 1999 512 2000
rect 506 1995 507 1999
rect 511 1995 512 1999
rect 506 1994 512 1995
rect 508 1960 510 1994
rect 506 1959 512 1960
rect 506 1955 507 1959
rect 511 1955 512 1959
rect 506 1954 512 1955
rect 516 1939 518 2004
rect 640 2000 642 2150
rect 836 2104 838 2165
rect 958 2111 964 2112
rect 958 2107 959 2111
rect 963 2107 964 2111
rect 958 2106 964 2107
rect 834 2103 840 2104
rect 834 2099 835 2103
rect 839 2099 840 2103
rect 834 2098 840 2099
rect 862 2088 868 2089
rect 862 2084 863 2088
rect 867 2084 868 2088
rect 862 2083 868 2084
rect 864 2055 866 2083
rect 687 2054 691 2055
rect 687 2049 691 2050
rect 831 2054 835 2055
rect 831 2049 835 2050
rect 863 2054 867 2055
rect 863 2049 867 2050
rect 688 2025 690 2049
rect 832 2025 834 2049
rect 686 2024 692 2025
rect 686 2020 687 2024
rect 691 2020 692 2024
rect 686 2019 692 2020
rect 830 2024 836 2025
rect 830 2020 831 2024
rect 835 2020 836 2024
rect 830 2019 836 2020
rect 658 2009 664 2010
rect 658 2005 659 2009
rect 663 2005 664 2009
rect 658 2004 664 2005
rect 802 2009 808 2010
rect 802 2005 803 2009
rect 807 2005 808 2009
rect 802 2004 808 2005
rect 946 2009 952 2010
rect 946 2005 947 2009
rect 951 2005 952 2009
rect 946 2004 952 2005
rect 638 1999 644 2000
rect 638 1995 639 1999
rect 643 1995 644 1999
rect 638 1994 644 1995
rect 660 1939 662 2004
rect 682 1999 688 2000
rect 682 1995 683 1999
rect 687 1995 688 1999
rect 682 1994 688 1995
rect 379 1938 383 1939
rect 379 1933 383 1934
rect 515 1938 519 1939
rect 515 1933 519 1934
rect 587 1938 591 1939
rect 587 1933 591 1934
rect 659 1938 663 1939
rect 659 1933 663 1934
rect 310 1879 316 1880
rect 310 1875 311 1879
rect 315 1875 316 1879
rect 310 1874 316 1875
rect 380 1872 382 1933
rect 474 1919 480 1920
rect 474 1915 475 1919
rect 479 1915 480 1919
rect 474 1914 480 1915
rect 110 1868 111 1872
rect 115 1868 116 1872
rect 110 1867 116 1868
rect 186 1871 192 1872
rect 186 1867 187 1871
rect 191 1867 192 1871
rect 186 1866 192 1867
rect 378 1871 384 1872
rect 378 1867 379 1871
rect 383 1867 384 1871
rect 378 1866 384 1867
rect 214 1856 220 1857
rect 110 1855 116 1856
rect 110 1851 111 1855
rect 115 1851 116 1855
rect 214 1852 215 1856
rect 219 1852 220 1856
rect 214 1851 220 1852
rect 406 1856 412 1857
rect 406 1852 407 1856
rect 411 1852 412 1856
rect 406 1851 412 1852
rect 110 1850 116 1851
rect 112 1819 114 1850
rect 216 1819 218 1851
rect 408 1819 410 1851
rect 111 1818 115 1819
rect 111 1813 115 1814
rect 159 1818 163 1819
rect 159 1813 163 1814
rect 215 1818 219 1819
rect 215 1813 219 1814
rect 375 1818 379 1819
rect 375 1813 379 1814
rect 407 1818 411 1819
rect 407 1813 411 1814
rect 112 1790 114 1813
rect 110 1789 116 1790
rect 160 1789 162 1813
rect 376 1789 378 1813
rect 110 1785 111 1789
rect 115 1785 116 1789
rect 110 1784 116 1785
rect 158 1788 164 1789
rect 158 1784 159 1788
rect 163 1784 164 1788
rect 158 1783 164 1784
rect 374 1788 380 1789
rect 374 1784 375 1788
rect 379 1784 380 1788
rect 374 1783 380 1784
rect 130 1773 136 1774
rect 110 1772 116 1773
rect 110 1768 111 1772
rect 115 1768 116 1772
rect 130 1769 131 1773
rect 135 1769 136 1773
rect 130 1768 136 1769
rect 346 1773 352 1774
rect 346 1769 347 1773
rect 351 1769 352 1773
rect 346 1768 352 1769
rect 110 1767 116 1768
rect 112 1683 114 1767
rect 132 1683 134 1768
rect 290 1763 296 1764
rect 290 1759 291 1763
rect 295 1759 296 1763
rect 290 1758 296 1759
rect 292 1724 294 1758
rect 226 1723 232 1724
rect 226 1719 227 1723
rect 231 1719 232 1723
rect 226 1718 232 1719
rect 290 1723 296 1724
rect 290 1719 291 1723
rect 295 1719 296 1723
rect 290 1718 296 1719
rect 111 1682 115 1683
rect 111 1677 115 1678
rect 131 1682 135 1683
rect 131 1677 135 1678
rect 112 1617 114 1677
rect 110 1616 116 1617
rect 132 1616 134 1677
rect 228 1624 230 1718
rect 348 1683 350 1768
rect 476 1764 478 1914
rect 588 1872 590 1933
rect 684 1924 686 1994
rect 804 1939 806 2004
rect 948 1939 950 2004
rect 960 1960 962 2106
rect 1076 2104 1078 2165
rect 1160 2156 1162 2234
rect 1936 2171 1938 2243
rect 1976 2239 1978 2270
rect 2024 2239 2026 2271
rect 2184 2239 2186 2271
rect 2376 2239 2378 2271
rect 1975 2238 1979 2239
rect 1975 2233 1979 2234
rect 2023 2238 2027 2239
rect 2023 2233 2027 2234
rect 2183 2238 2187 2239
rect 2183 2233 2187 2234
rect 2191 2238 2195 2239
rect 2191 2233 2195 2234
rect 2359 2238 2363 2239
rect 2359 2233 2363 2234
rect 2375 2238 2379 2239
rect 2375 2233 2379 2234
rect 1976 2210 1978 2233
rect 1974 2209 1980 2210
rect 2024 2209 2026 2233
rect 2192 2209 2194 2233
rect 2360 2209 2362 2233
rect 1974 2205 1975 2209
rect 1979 2205 1980 2209
rect 1974 2204 1980 2205
rect 2022 2208 2028 2209
rect 2022 2204 2023 2208
rect 2027 2204 2028 2208
rect 2022 2203 2028 2204
rect 2190 2208 2196 2209
rect 2190 2204 2191 2208
rect 2195 2204 2196 2208
rect 2190 2203 2196 2204
rect 2358 2208 2364 2209
rect 2358 2204 2359 2208
rect 2363 2204 2364 2208
rect 2358 2203 2364 2204
rect 1994 2193 2000 2194
rect 1974 2192 1980 2193
rect 1974 2188 1975 2192
rect 1979 2188 1980 2192
rect 1994 2189 1995 2193
rect 1999 2189 2000 2193
rect 1994 2188 2000 2189
rect 2162 2193 2168 2194
rect 2162 2189 2163 2193
rect 2167 2189 2168 2193
rect 2162 2188 2168 2189
rect 2330 2193 2336 2194
rect 2330 2189 2331 2193
rect 2335 2189 2336 2193
rect 2330 2188 2336 2189
rect 1974 2187 1980 2188
rect 1315 2170 1319 2171
rect 1315 2165 1319 2166
rect 1563 2170 1567 2171
rect 1563 2165 1567 2166
rect 1787 2170 1791 2171
rect 1787 2165 1791 2166
rect 1935 2170 1939 2171
rect 1935 2165 1939 2166
rect 1158 2155 1164 2156
rect 1158 2151 1159 2155
rect 1163 2151 1164 2155
rect 1158 2150 1164 2151
rect 1316 2104 1318 2165
rect 1438 2111 1444 2112
rect 1438 2107 1439 2111
rect 1443 2107 1444 2111
rect 1438 2106 1444 2107
rect 1074 2103 1080 2104
rect 1074 2099 1075 2103
rect 1079 2099 1080 2103
rect 1074 2098 1080 2099
rect 1314 2103 1320 2104
rect 1314 2099 1315 2103
rect 1319 2099 1320 2103
rect 1314 2098 1320 2099
rect 1102 2088 1108 2089
rect 1102 2084 1103 2088
rect 1107 2084 1108 2088
rect 1102 2083 1108 2084
rect 1342 2088 1348 2089
rect 1342 2084 1343 2088
rect 1347 2084 1348 2088
rect 1342 2083 1348 2084
rect 1104 2055 1106 2083
rect 1344 2055 1346 2083
rect 975 2054 979 2055
rect 975 2049 979 2050
rect 1103 2054 1107 2055
rect 1103 2049 1107 2050
rect 1119 2054 1123 2055
rect 1119 2049 1123 2050
rect 1263 2054 1267 2055
rect 1263 2049 1267 2050
rect 1343 2054 1347 2055
rect 1343 2049 1347 2050
rect 1407 2054 1411 2055
rect 1407 2049 1411 2050
rect 976 2025 978 2049
rect 1120 2025 1122 2049
rect 1264 2025 1266 2049
rect 1408 2025 1410 2049
rect 974 2024 980 2025
rect 974 2020 975 2024
rect 979 2020 980 2024
rect 974 2019 980 2020
rect 1118 2024 1124 2025
rect 1118 2020 1119 2024
rect 1123 2020 1124 2024
rect 1118 2019 1124 2020
rect 1262 2024 1268 2025
rect 1262 2020 1263 2024
rect 1267 2020 1268 2024
rect 1262 2019 1268 2020
rect 1406 2024 1412 2025
rect 1406 2020 1407 2024
rect 1411 2020 1412 2024
rect 1406 2019 1412 2020
rect 1090 2009 1096 2010
rect 1090 2005 1091 2009
rect 1095 2005 1096 2009
rect 1090 2004 1096 2005
rect 1234 2009 1240 2010
rect 1234 2005 1235 2009
rect 1239 2005 1240 2009
rect 1234 2004 1240 2005
rect 1378 2009 1384 2010
rect 1378 2005 1379 2009
rect 1383 2005 1384 2009
rect 1378 2004 1384 2005
rect 958 1959 964 1960
rect 958 1955 959 1959
rect 963 1955 964 1959
rect 958 1954 964 1955
rect 1092 1939 1094 2004
rect 1218 1999 1224 2000
rect 1218 1995 1219 1999
rect 1223 1995 1224 1999
rect 1218 1994 1224 1995
rect 1186 1991 1192 1992
rect 1186 1987 1187 1991
rect 1191 1987 1192 1991
rect 1186 1986 1192 1987
rect 1188 1960 1190 1986
rect 1220 1960 1222 1994
rect 1186 1959 1192 1960
rect 1186 1955 1187 1959
rect 1191 1955 1192 1959
rect 1186 1954 1192 1955
rect 1218 1959 1224 1960
rect 1218 1955 1219 1959
rect 1223 1955 1224 1959
rect 1218 1954 1224 1955
rect 1236 1939 1238 2004
rect 1358 1999 1364 2000
rect 1358 1995 1359 1999
rect 1363 1995 1364 1999
rect 1358 1994 1364 1995
rect 803 1938 807 1939
rect 803 1933 807 1934
rect 811 1938 815 1939
rect 811 1933 815 1934
rect 947 1938 951 1939
rect 947 1933 951 1934
rect 1051 1938 1055 1939
rect 1051 1933 1055 1934
rect 1091 1938 1095 1939
rect 1091 1933 1095 1934
rect 1235 1938 1239 1939
rect 1235 1933 1239 1934
rect 1299 1938 1303 1939
rect 1299 1933 1303 1934
rect 682 1923 688 1924
rect 682 1919 683 1923
rect 687 1919 688 1923
rect 682 1918 688 1919
rect 812 1872 814 1933
rect 818 1919 824 1920
rect 818 1915 819 1919
rect 823 1915 824 1919
rect 818 1914 824 1915
rect 820 1880 822 1914
rect 818 1879 824 1880
rect 818 1875 819 1879
rect 823 1875 824 1879
rect 818 1874 824 1875
rect 1052 1872 1054 1933
rect 1058 1919 1064 1920
rect 1058 1915 1059 1919
rect 1063 1915 1064 1919
rect 1058 1914 1064 1915
rect 1060 1880 1062 1914
rect 1058 1879 1064 1880
rect 1058 1875 1059 1879
rect 1063 1875 1064 1879
rect 1058 1874 1064 1875
rect 1134 1879 1140 1880
rect 1134 1875 1135 1879
rect 1139 1875 1140 1879
rect 1134 1874 1140 1875
rect 586 1871 592 1872
rect 586 1867 587 1871
rect 591 1867 592 1871
rect 586 1866 592 1867
rect 810 1871 816 1872
rect 810 1867 811 1871
rect 815 1867 816 1871
rect 810 1866 816 1867
rect 1050 1871 1056 1872
rect 1050 1867 1051 1871
rect 1055 1867 1056 1871
rect 1050 1866 1056 1867
rect 614 1856 620 1857
rect 614 1852 615 1856
rect 619 1852 620 1856
rect 614 1851 620 1852
rect 838 1856 844 1857
rect 838 1852 839 1856
rect 843 1852 844 1856
rect 838 1851 844 1852
rect 1078 1856 1084 1857
rect 1078 1852 1079 1856
rect 1083 1852 1084 1856
rect 1078 1851 1084 1852
rect 616 1819 618 1851
rect 840 1819 842 1851
rect 1080 1819 1082 1851
rect 591 1818 595 1819
rect 591 1813 595 1814
rect 615 1818 619 1819
rect 615 1813 619 1814
rect 799 1818 803 1819
rect 799 1813 803 1814
rect 839 1818 843 1819
rect 839 1813 843 1814
rect 999 1818 1003 1819
rect 999 1813 1003 1814
rect 1079 1818 1083 1819
rect 1079 1813 1083 1814
rect 592 1789 594 1813
rect 800 1789 802 1813
rect 1000 1789 1002 1813
rect 590 1788 596 1789
rect 590 1784 591 1788
rect 595 1784 596 1788
rect 590 1783 596 1784
rect 798 1788 804 1789
rect 798 1784 799 1788
rect 803 1784 804 1788
rect 798 1783 804 1784
rect 998 1788 1004 1789
rect 998 1784 999 1788
rect 1003 1784 1004 1788
rect 998 1783 1004 1784
rect 562 1773 568 1774
rect 562 1769 563 1773
rect 567 1769 568 1773
rect 562 1768 568 1769
rect 770 1773 776 1774
rect 770 1769 771 1773
rect 775 1769 776 1773
rect 770 1768 776 1769
rect 970 1773 976 1774
rect 970 1769 971 1773
rect 975 1769 976 1773
rect 970 1768 976 1769
rect 474 1763 480 1764
rect 474 1759 475 1763
rect 479 1759 480 1763
rect 474 1758 480 1759
rect 490 1763 496 1764
rect 490 1759 491 1763
rect 495 1759 496 1763
rect 490 1758 496 1759
rect 347 1682 351 1683
rect 347 1677 351 1678
rect 395 1682 399 1683
rect 395 1677 399 1678
rect 238 1667 244 1668
rect 238 1663 239 1667
rect 243 1663 244 1667
rect 238 1662 244 1663
rect 226 1623 232 1624
rect 226 1619 227 1623
rect 231 1619 232 1623
rect 226 1618 232 1619
rect 110 1612 111 1616
rect 115 1612 116 1616
rect 110 1611 116 1612
rect 130 1615 136 1616
rect 130 1611 131 1615
rect 135 1611 136 1615
rect 130 1610 136 1611
rect 158 1600 164 1601
rect 110 1599 116 1600
rect 110 1595 111 1599
rect 115 1595 116 1599
rect 158 1596 159 1600
rect 163 1596 164 1600
rect 158 1595 164 1596
rect 110 1594 116 1595
rect 112 1559 114 1594
rect 160 1559 162 1595
rect 111 1558 115 1559
rect 111 1553 115 1554
rect 159 1558 163 1559
rect 159 1553 163 1554
rect 112 1530 114 1553
rect 110 1529 116 1530
rect 160 1529 162 1553
rect 110 1525 111 1529
rect 115 1525 116 1529
rect 110 1524 116 1525
rect 158 1528 164 1529
rect 158 1524 159 1528
rect 163 1524 164 1528
rect 158 1523 164 1524
rect 130 1513 136 1514
rect 110 1512 116 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 130 1509 131 1513
rect 135 1509 136 1513
rect 130 1508 136 1509
rect 110 1507 116 1508
rect 112 1435 114 1507
rect 132 1435 134 1508
rect 240 1504 242 1662
rect 396 1616 398 1677
rect 492 1668 494 1758
rect 564 1683 566 1768
rect 772 1683 774 1768
rect 972 1683 974 1768
rect 1106 1763 1112 1764
rect 1106 1759 1107 1763
rect 1111 1759 1112 1763
rect 1106 1758 1112 1759
rect 1066 1755 1072 1756
rect 1066 1751 1067 1755
rect 1071 1751 1072 1755
rect 1066 1750 1072 1751
rect 1068 1724 1070 1750
rect 1108 1724 1110 1758
rect 1066 1723 1072 1724
rect 1066 1719 1067 1723
rect 1071 1719 1072 1723
rect 1066 1718 1072 1719
rect 1106 1723 1112 1724
rect 1106 1719 1107 1723
rect 1111 1719 1112 1723
rect 1106 1718 1112 1719
rect 1136 1716 1138 1874
rect 1300 1872 1302 1933
rect 1360 1924 1362 1994
rect 1380 1939 1382 2004
rect 1440 1960 1442 2106
rect 1564 2104 1566 2165
rect 1788 2104 1790 2165
rect 1794 2151 1800 2152
rect 1794 2147 1795 2151
rect 1799 2147 1800 2151
rect 1794 2146 1800 2147
rect 1562 2103 1568 2104
rect 1562 2099 1563 2103
rect 1567 2099 1568 2103
rect 1562 2098 1568 2099
rect 1786 2103 1792 2104
rect 1786 2099 1787 2103
rect 1791 2099 1792 2103
rect 1786 2098 1792 2099
rect 1590 2088 1596 2089
rect 1590 2084 1591 2088
rect 1595 2084 1596 2088
rect 1590 2083 1596 2084
rect 1592 2055 1594 2083
rect 1543 2054 1547 2055
rect 1543 2049 1547 2050
rect 1591 2054 1595 2055
rect 1591 2049 1595 2050
rect 1679 2054 1683 2055
rect 1679 2049 1683 2050
rect 1544 2025 1546 2049
rect 1680 2025 1682 2049
rect 1542 2024 1548 2025
rect 1542 2020 1543 2024
rect 1547 2020 1548 2024
rect 1542 2019 1548 2020
rect 1678 2024 1684 2025
rect 1678 2020 1679 2024
rect 1683 2020 1684 2024
rect 1678 2019 1684 2020
rect 1514 2009 1520 2010
rect 1514 2005 1515 2009
rect 1519 2005 1520 2009
rect 1514 2004 1520 2005
rect 1650 2009 1656 2010
rect 1650 2005 1651 2009
rect 1655 2005 1656 2009
rect 1650 2004 1656 2005
rect 1786 2009 1792 2010
rect 1786 2005 1787 2009
rect 1791 2005 1792 2009
rect 1786 2004 1792 2005
rect 1506 1999 1512 2000
rect 1506 1995 1507 1999
rect 1511 1995 1512 1999
rect 1506 1994 1512 1995
rect 1508 1960 1510 1994
rect 1438 1959 1444 1960
rect 1438 1955 1439 1959
rect 1443 1955 1444 1959
rect 1438 1954 1444 1955
rect 1506 1959 1512 1960
rect 1506 1955 1507 1959
rect 1511 1955 1512 1959
rect 1506 1954 1512 1955
rect 1516 1939 1518 2004
rect 1652 1939 1654 2004
rect 1746 1991 1752 1992
rect 1746 1987 1747 1991
rect 1751 1987 1752 1991
rect 1746 1986 1752 1987
rect 1748 1960 1750 1986
rect 1746 1959 1752 1960
rect 1746 1955 1747 1959
rect 1751 1955 1752 1959
rect 1746 1954 1752 1955
rect 1788 1939 1790 2004
rect 1796 2000 1798 2146
rect 1936 2105 1938 2165
rect 1976 2111 1978 2187
rect 1996 2111 1998 2188
rect 2122 2183 2128 2184
rect 2122 2179 2123 2183
rect 2127 2179 2128 2183
rect 2122 2178 2128 2179
rect 2124 2144 2126 2178
rect 2122 2143 2128 2144
rect 2122 2139 2123 2143
rect 2127 2139 2128 2143
rect 2122 2138 2128 2139
rect 2164 2111 2166 2188
rect 2290 2183 2296 2184
rect 2290 2179 2291 2183
rect 2295 2179 2296 2183
rect 2290 2178 2296 2179
rect 2292 2144 2294 2178
rect 2290 2143 2296 2144
rect 2290 2139 2291 2143
rect 2295 2139 2296 2143
rect 2290 2138 2296 2139
rect 2332 2111 2334 2188
rect 2458 2183 2464 2184
rect 2458 2179 2459 2183
rect 2463 2179 2464 2183
rect 2458 2178 2464 2179
rect 2460 2144 2462 2178
rect 2458 2143 2464 2144
rect 2458 2139 2459 2143
rect 2463 2139 2464 2143
rect 2458 2138 2464 2139
rect 2472 2136 2474 2294
rect 2540 2292 2542 2353
rect 2548 2300 2550 2370
rect 2652 2359 2654 2428
rect 2776 2424 2778 2594
rect 2828 2548 2830 2609
rect 2950 2555 2956 2556
rect 2950 2551 2951 2555
rect 2955 2551 2956 2555
rect 2950 2550 2956 2551
rect 2826 2547 2832 2548
rect 2826 2543 2827 2547
rect 2831 2543 2832 2547
rect 2826 2542 2832 2543
rect 2854 2532 2860 2533
rect 2854 2528 2855 2532
rect 2859 2528 2860 2532
rect 2854 2527 2860 2528
rect 2856 2479 2858 2527
rect 2855 2478 2859 2479
rect 2855 2473 2859 2474
rect 2927 2478 2931 2479
rect 2927 2473 2931 2474
rect 2928 2449 2930 2473
rect 2926 2448 2932 2449
rect 2926 2444 2927 2448
rect 2931 2444 2932 2448
rect 2926 2443 2932 2444
rect 2898 2433 2904 2434
rect 2898 2429 2899 2433
rect 2903 2429 2904 2433
rect 2898 2428 2904 2429
rect 2774 2423 2780 2424
rect 2774 2419 2775 2423
rect 2779 2419 2780 2423
rect 2774 2418 2780 2419
rect 2900 2359 2902 2428
rect 2952 2384 2954 2550
rect 2964 2548 2966 2609
rect 3100 2548 3102 2609
rect 3112 2600 3114 2678
rect 3800 2615 3802 2687
rect 3840 2670 3842 2693
rect 3838 2669 3844 2670
rect 3960 2669 3962 2693
rect 3838 2665 3839 2669
rect 3843 2665 3844 2669
rect 3838 2664 3844 2665
rect 3958 2668 3964 2669
rect 3958 2664 3959 2668
rect 3963 2664 3964 2668
rect 3958 2663 3964 2664
rect 3930 2653 3936 2654
rect 3838 2652 3844 2653
rect 3838 2648 3839 2652
rect 3843 2648 3844 2652
rect 3930 2649 3931 2653
rect 3935 2649 3936 2653
rect 3930 2648 3936 2649
rect 3838 2647 3844 2648
rect 3799 2614 3803 2615
rect 3799 2609 3803 2610
rect 3110 2599 3116 2600
rect 3110 2595 3111 2599
rect 3115 2595 3116 2599
rect 3110 2594 3116 2595
rect 3800 2549 3802 2609
rect 3840 2587 3842 2647
rect 3932 2587 3934 2648
rect 4056 2644 4058 2790
rect 4132 2744 4134 2805
rect 4268 2744 4270 2805
rect 4274 2791 4280 2792
rect 4274 2787 4275 2791
rect 4279 2787 4280 2791
rect 4274 2786 4280 2787
rect 4276 2752 4278 2786
rect 4274 2751 4280 2752
rect 4274 2747 4275 2751
rect 4279 2747 4280 2751
rect 4274 2746 4280 2747
rect 4404 2744 4406 2805
rect 4410 2791 4416 2792
rect 4410 2787 4411 2791
rect 4415 2787 4416 2791
rect 4410 2786 4416 2787
rect 4412 2752 4414 2786
rect 4410 2751 4416 2752
rect 4410 2747 4411 2751
rect 4415 2747 4416 2751
rect 4410 2746 4416 2747
rect 4540 2744 4542 2805
rect 4546 2791 4552 2792
rect 4546 2787 4547 2791
rect 4551 2787 4552 2791
rect 4546 2786 4552 2787
rect 4548 2752 4550 2786
rect 4546 2751 4552 2752
rect 4546 2747 4547 2751
rect 4551 2747 4552 2751
rect 4546 2746 4552 2747
rect 4676 2744 4678 2805
rect 4682 2791 4688 2792
rect 4682 2787 4683 2791
rect 4687 2787 4688 2791
rect 4682 2786 4688 2787
rect 4684 2752 4686 2786
rect 4682 2751 4688 2752
rect 4682 2747 4683 2751
rect 4687 2747 4688 2751
rect 4682 2746 4688 2747
rect 4812 2744 4814 2805
rect 4818 2791 4824 2792
rect 4818 2787 4819 2791
rect 4823 2787 4824 2791
rect 4818 2786 4824 2787
rect 4820 2752 4822 2786
rect 4818 2751 4824 2752
rect 4818 2747 4819 2751
rect 4823 2747 4824 2751
rect 4818 2746 4824 2747
rect 4830 2751 4836 2752
rect 4830 2747 4831 2751
rect 4835 2747 4836 2751
rect 4830 2746 4836 2747
rect 4130 2743 4136 2744
rect 4130 2739 4131 2743
rect 4135 2739 4136 2743
rect 4130 2738 4136 2739
rect 4266 2743 4272 2744
rect 4266 2739 4267 2743
rect 4271 2739 4272 2743
rect 4266 2738 4272 2739
rect 4402 2743 4408 2744
rect 4402 2739 4403 2743
rect 4407 2739 4408 2743
rect 4402 2738 4408 2739
rect 4538 2743 4544 2744
rect 4538 2739 4539 2743
rect 4543 2739 4544 2743
rect 4538 2738 4544 2739
rect 4674 2743 4680 2744
rect 4674 2739 4675 2743
rect 4679 2739 4680 2743
rect 4674 2738 4680 2739
rect 4810 2743 4816 2744
rect 4810 2739 4811 2743
rect 4815 2739 4816 2743
rect 4810 2738 4816 2739
rect 4158 2728 4164 2729
rect 4158 2724 4159 2728
rect 4163 2724 4164 2728
rect 4158 2723 4164 2724
rect 4294 2728 4300 2729
rect 4294 2724 4295 2728
rect 4299 2724 4300 2728
rect 4294 2723 4300 2724
rect 4430 2728 4436 2729
rect 4430 2724 4431 2728
rect 4435 2724 4436 2728
rect 4430 2723 4436 2724
rect 4566 2728 4572 2729
rect 4566 2724 4567 2728
rect 4571 2724 4572 2728
rect 4566 2723 4572 2724
rect 4702 2728 4708 2729
rect 4702 2724 4703 2728
rect 4707 2724 4708 2728
rect 4702 2723 4708 2724
rect 4160 2699 4162 2723
rect 4296 2699 4298 2723
rect 4432 2699 4434 2723
rect 4568 2699 4570 2723
rect 4704 2699 4706 2723
rect 4159 2698 4163 2699
rect 4159 2693 4163 2694
rect 4255 2698 4259 2699
rect 4255 2693 4259 2694
rect 4295 2698 4299 2699
rect 4295 2693 4299 2694
rect 4431 2698 4435 2699
rect 4431 2693 4435 2694
rect 4543 2698 4547 2699
rect 4543 2693 4547 2694
rect 4567 2698 4571 2699
rect 4567 2693 4571 2694
rect 4703 2698 4707 2699
rect 4703 2693 4707 2694
rect 4823 2698 4827 2699
rect 4823 2693 4827 2694
rect 4256 2669 4258 2693
rect 4544 2669 4546 2693
rect 4824 2669 4826 2693
rect 4254 2668 4260 2669
rect 4254 2664 4255 2668
rect 4259 2664 4260 2668
rect 4254 2663 4260 2664
rect 4542 2668 4548 2669
rect 4542 2664 4543 2668
rect 4547 2664 4548 2668
rect 4542 2663 4548 2664
rect 4822 2668 4828 2669
rect 4822 2664 4823 2668
rect 4827 2664 4828 2668
rect 4822 2663 4828 2664
rect 4226 2653 4232 2654
rect 4226 2649 4227 2653
rect 4231 2649 4232 2653
rect 4226 2648 4232 2649
rect 4514 2653 4520 2654
rect 4514 2649 4515 2653
rect 4519 2649 4520 2653
rect 4514 2648 4520 2649
rect 4794 2653 4800 2654
rect 4794 2649 4795 2653
rect 4799 2649 4800 2653
rect 4794 2648 4800 2649
rect 4054 2643 4060 2644
rect 4054 2639 4055 2643
rect 4059 2639 4060 2643
rect 4054 2638 4060 2639
rect 3982 2603 3988 2604
rect 3982 2599 3983 2603
rect 3987 2599 3988 2603
rect 3982 2598 3988 2599
rect 3839 2586 3843 2587
rect 3839 2581 3843 2582
rect 3859 2586 3863 2587
rect 3859 2581 3863 2582
rect 3931 2586 3935 2587
rect 3931 2581 3935 2582
rect 3798 2548 3804 2549
rect 2962 2547 2968 2548
rect 2962 2543 2963 2547
rect 2967 2543 2968 2547
rect 2962 2542 2968 2543
rect 3098 2547 3104 2548
rect 3098 2543 3099 2547
rect 3103 2543 3104 2547
rect 3798 2544 3799 2548
rect 3803 2544 3804 2548
rect 3798 2543 3804 2544
rect 3098 2542 3104 2543
rect 2990 2532 2996 2533
rect 2990 2528 2991 2532
rect 2995 2528 2996 2532
rect 2990 2527 2996 2528
rect 3126 2532 3132 2533
rect 3126 2528 3127 2532
rect 3131 2528 3132 2532
rect 3126 2527 3132 2528
rect 3798 2531 3804 2532
rect 3798 2527 3799 2531
rect 3803 2527 3804 2531
rect 2992 2479 2994 2527
rect 3128 2479 3130 2527
rect 3798 2526 3804 2527
rect 3800 2479 3802 2526
rect 3840 2521 3842 2581
rect 3838 2520 3844 2521
rect 3860 2520 3862 2581
rect 3984 2528 3986 2598
rect 4228 2587 4230 2648
rect 4442 2643 4448 2644
rect 4442 2639 4443 2643
rect 4447 2639 4448 2643
rect 4442 2638 4448 2639
rect 4322 2627 4328 2628
rect 4322 2623 4323 2627
rect 4327 2623 4328 2627
rect 4322 2622 4328 2623
rect 4324 2604 4326 2622
rect 4444 2604 4446 2638
rect 4322 2603 4328 2604
rect 4322 2599 4323 2603
rect 4327 2599 4328 2603
rect 4322 2598 4328 2599
rect 4442 2603 4448 2604
rect 4442 2599 4443 2603
rect 4447 2599 4448 2603
rect 4442 2598 4448 2599
rect 4516 2587 4518 2648
rect 4638 2643 4644 2644
rect 4638 2639 4639 2643
rect 4643 2639 4644 2643
rect 4638 2638 4644 2639
rect 4083 2586 4087 2587
rect 4083 2581 4087 2582
rect 4227 2586 4231 2587
rect 4227 2581 4231 2582
rect 4331 2586 4335 2587
rect 4331 2581 4335 2582
rect 4515 2586 4519 2587
rect 4515 2581 4519 2582
rect 4579 2586 4583 2587
rect 4579 2581 4583 2582
rect 3982 2527 3988 2528
rect 3982 2523 3983 2527
rect 3987 2523 3988 2527
rect 3982 2522 3988 2523
rect 4084 2520 4086 2581
rect 4178 2567 4184 2568
rect 4178 2563 4179 2567
rect 4183 2563 4184 2567
rect 4178 2562 4184 2563
rect 3838 2516 3839 2520
rect 3843 2516 3844 2520
rect 3838 2515 3844 2516
rect 3858 2519 3864 2520
rect 3858 2515 3859 2519
rect 3863 2515 3864 2519
rect 3858 2514 3864 2515
rect 4082 2519 4088 2520
rect 4082 2515 4083 2519
rect 4087 2515 4088 2519
rect 4082 2514 4088 2515
rect 3886 2504 3892 2505
rect 3838 2503 3844 2504
rect 3838 2499 3839 2503
rect 3843 2499 3844 2503
rect 3886 2500 3887 2504
rect 3891 2500 3892 2504
rect 3886 2499 3892 2500
rect 4110 2504 4116 2505
rect 4110 2500 4111 2504
rect 4115 2500 4116 2504
rect 4110 2499 4116 2500
rect 3838 2498 3844 2499
rect 2991 2478 2995 2479
rect 2991 2473 2995 2474
rect 3127 2478 3131 2479
rect 3127 2473 3131 2474
rect 3183 2478 3187 2479
rect 3183 2473 3187 2474
rect 3439 2478 3443 2479
rect 3439 2473 3443 2474
rect 3679 2478 3683 2479
rect 3679 2473 3683 2474
rect 3799 2478 3803 2479
rect 3799 2473 3803 2474
rect 3184 2449 3186 2473
rect 3440 2449 3442 2473
rect 3680 2449 3682 2473
rect 3800 2450 3802 2473
rect 3840 2471 3842 2498
rect 3888 2471 3890 2499
rect 4112 2471 4114 2499
rect 3839 2470 3843 2471
rect 3839 2465 3843 2466
rect 3887 2470 3891 2471
rect 3887 2465 3891 2466
rect 4087 2470 4091 2471
rect 4087 2465 4091 2466
rect 4111 2470 4115 2471
rect 4111 2465 4115 2466
rect 3798 2449 3804 2450
rect 3182 2448 3188 2449
rect 3182 2444 3183 2448
rect 3187 2444 3188 2448
rect 3182 2443 3188 2444
rect 3438 2448 3444 2449
rect 3438 2444 3439 2448
rect 3443 2444 3444 2448
rect 3438 2443 3444 2444
rect 3678 2448 3684 2449
rect 3678 2444 3679 2448
rect 3683 2444 3684 2448
rect 3798 2445 3799 2449
rect 3803 2445 3804 2449
rect 3798 2444 3804 2445
rect 3678 2443 3684 2444
rect 3840 2442 3842 2465
rect 3838 2441 3844 2442
rect 3888 2441 3890 2465
rect 4088 2441 4090 2465
rect 3838 2437 3839 2441
rect 3843 2437 3844 2441
rect 3838 2436 3844 2437
rect 3886 2440 3892 2441
rect 3886 2436 3887 2440
rect 3891 2436 3892 2440
rect 3886 2435 3892 2436
rect 4086 2440 4092 2441
rect 4086 2436 4087 2440
rect 4091 2436 4092 2440
rect 4086 2435 4092 2436
rect 3154 2433 3160 2434
rect 3154 2429 3155 2433
rect 3159 2429 3160 2433
rect 3154 2428 3160 2429
rect 3410 2433 3416 2434
rect 3410 2429 3411 2433
rect 3415 2429 3416 2433
rect 3410 2428 3416 2429
rect 3650 2433 3656 2434
rect 3650 2429 3651 2433
rect 3655 2429 3656 2433
rect 3650 2428 3656 2429
rect 3798 2432 3804 2433
rect 3798 2428 3799 2432
rect 3803 2428 3804 2432
rect 3026 2423 3032 2424
rect 3026 2419 3027 2423
rect 3031 2419 3032 2423
rect 3026 2418 3032 2419
rect 3028 2384 3030 2418
rect 2950 2383 2956 2384
rect 2950 2379 2951 2383
rect 2955 2379 2956 2383
rect 2950 2378 2956 2379
rect 3026 2383 3032 2384
rect 3026 2379 3027 2383
rect 3031 2379 3032 2383
rect 3026 2378 3032 2379
rect 3156 2359 3158 2428
rect 3282 2423 3288 2424
rect 3282 2419 3283 2423
rect 3287 2419 3288 2423
rect 3282 2418 3288 2419
rect 3284 2384 3286 2418
rect 3282 2383 3288 2384
rect 3282 2379 3283 2383
rect 3287 2379 3288 2383
rect 3282 2378 3288 2379
rect 3412 2359 3414 2428
rect 3534 2423 3540 2424
rect 3534 2419 3535 2423
rect 3539 2419 3540 2423
rect 3534 2418 3540 2419
rect 2651 2358 2655 2359
rect 2651 2353 2655 2354
rect 2731 2358 2735 2359
rect 2731 2353 2735 2354
rect 2899 2358 2903 2359
rect 2899 2353 2903 2354
rect 2923 2358 2927 2359
rect 2923 2353 2927 2354
rect 3115 2358 3119 2359
rect 3115 2353 3119 2354
rect 3155 2358 3159 2359
rect 3155 2353 3159 2354
rect 3299 2358 3303 2359
rect 3299 2353 3303 2354
rect 3411 2358 3415 2359
rect 3411 2353 3415 2354
rect 3483 2358 3487 2359
rect 3483 2353 3487 2354
rect 2546 2299 2552 2300
rect 2546 2295 2547 2299
rect 2551 2295 2552 2299
rect 2546 2294 2552 2295
rect 2732 2292 2734 2353
rect 2806 2343 2812 2344
rect 2806 2339 2807 2343
rect 2811 2339 2812 2343
rect 2806 2338 2812 2339
rect 2538 2291 2544 2292
rect 2538 2287 2539 2291
rect 2543 2287 2544 2291
rect 2538 2286 2544 2287
rect 2730 2291 2736 2292
rect 2730 2287 2731 2291
rect 2735 2287 2736 2291
rect 2730 2286 2736 2287
rect 2566 2276 2572 2277
rect 2566 2272 2567 2276
rect 2571 2272 2572 2276
rect 2566 2271 2572 2272
rect 2758 2276 2764 2277
rect 2758 2272 2759 2276
rect 2763 2272 2764 2276
rect 2758 2271 2764 2272
rect 2568 2239 2570 2271
rect 2760 2239 2762 2271
rect 2535 2238 2539 2239
rect 2535 2233 2539 2234
rect 2567 2238 2571 2239
rect 2567 2233 2571 2234
rect 2711 2238 2715 2239
rect 2711 2233 2715 2234
rect 2759 2238 2763 2239
rect 2759 2233 2763 2234
rect 2536 2209 2538 2233
rect 2712 2209 2714 2233
rect 2534 2208 2540 2209
rect 2534 2204 2535 2208
rect 2539 2204 2540 2208
rect 2534 2203 2540 2204
rect 2710 2208 2716 2209
rect 2710 2204 2711 2208
rect 2715 2204 2716 2208
rect 2710 2203 2716 2204
rect 2506 2193 2512 2194
rect 2506 2189 2507 2193
rect 2511 2189 2512 2193
rect 2506 2188 2512 2189
rect 2682 2193 2688 2194
rect 2682 2189 2683 2193
rect 2687 2189 2688 2193
rect 2682 2188 2688 2189
rect 2470 2135 2476 2136
rect 2470 2131 2471 2135
rect 2475 2131 2476 2135
rect 2470 2130 2476 2131
rect 2508 2111 2510 2188
rect 2634 2183 2640 2184
rect 2634 2179 2635 2183
rect 2639 2179 2640 2183
rect 2634 2178 2640 2179
rect 2636 2144 2638 2178
rect 2634 2143 2640 2144
rect 2634 2139 2635 2143
rect 2639 2139 2640 2143
rect 2634 2138 2640 2139
rect 2684 2111 2686 2188
rect 2808 2184 2810 2338
rect 2924 2292 2926 2353
rect 3018 2339 3024 2340
rect 3018 2335 3019 2339
rect 3023 2335 3024 2339
rect 3018 2334 3024 2335
rect 3020 2308 3022 2334
rect 3018 2307 3024 2308
rect 3018 2303 3019 2307
rect 3023 2303 3024 2307
rect 3018 2302 3024 2303
rect 3116 2292 3118 2353
rect 3122 2339 3128 2340
rect 3122 2335 3123 2339
rect 3127 2335 3128 2339
rect 3122 2334 3128 2335
rect 3124 2300 3126 2334
rect 3122 2299 3128 2300
rect 3122 2295 3123 2299
rect 3127 2295 3128 2299
rect 3122 2294 3128 2295
rect 3238 2299 3244 2300
rect 3238 2295 3239 2299
rect 3243 2295 3244 2299
rect 3238 2294 3244 2295
rect 2922 2291 2928 2292
rect 2922 2287 2923 2291
rect 2927 2287 2928 2291
rect 2922 2286 2928 2287
rect 3114 2291 3120 2292
rect 3114 2287 3115 2291
rect 3119 2287 3120 2291
rect 3114 2286 3120 2287
rect 2950 2276 2956 2277
rect 2950 2272 2951 2276
rect 2955 2272 2956 2276
rect 2950 2271 2956 2272
rect 3142 2276 3148 2277
rect 3142 2272 3143 2276
rect 3147 2272 3148 2276
rect 3142 2271 3148 2272
rect 2952 2239 2954 2271
rect 3144 2239 3146 2271
rect 2879 2238 2883 2239
rect 2879 2233 2883 2234
rect 2951 2238 2955 2239
rect 2951 2233 2955 2234
rect 3047 2238 3051 2239
rect 3047 2233 3051 2234
rect 3143 2238 3147 2239
rect 3143 2233 3147 2234
rect 3207 2238 3211 2239
rect 3207 2233 3211 2234
rect 2880 2209 2882 2233
rect 3048 2209 3050 2233
rect 3208 2209 3210 2233
rect 2878 2208 2884 2209
rect 2878 2204 2879 2208
rect 2883 2204 2884 2208
rect 2878 2203 2884 2204
rect 3046 2208 3052 2209
rect 3046 2204 3047 2208
rect 3051 2204 3052 2208
rect 3046 2203 3052 2204
rect 3206 2208 3212 2209
rect 3206 2204 3207 2208
rect 3211 2204 3212 2208
rect 3206 2203 3212 2204
rect 2850 2193 2856 2194
rect 2850 2189 2851 2193
rect 2855 2189 2856 2193
rect 2850 2188 2856 2189
rect 3018 2193 3024 2194
rect 3018 2189 3019 2193
rect 3023 2189 3024 2193
rect 3018 2188 3024 2189
rect 3178 2193 3184 2194
rect 3178 2189 3179 2193
rect 3183 2189 3184 2193
rect 3178 2188 3184 2189
rect 2806 2183 2812 2184
rect 2806 2179 2807 2183
rect 2811 2179 2812 2183
rect 2806 2178 2812 2179
rect 2852 2111 2854 2188
rect 2978 2183 2984 2184
rect 2978 2179 2979 2183
rect 2983 2179 2984 2183
rect 2978 2178 2984 2179
rect 2946 2175 2952 2176
rect 2946 2171 2947 2175
rect 2951 2171 2952 2175
rect 2946 2170 2952 2171
rect 2948 2144 2950 2170
rect 2980 2144 2982 2178
rect 2946 2143 2952 2144
rect 2946 2139 2947 2143
rect 2951 2139 2952 2143
rect 2946 2138 2952 2139
rect 2978 2143 2984 2144
rect 2978 2139 2979 2143
rect 2983 2139 2984 2143
rect 2978 2138 2984 2139
rect 3020 2111 3022 2188
rect 3142 2183 3148 2184
rect 3142 2179 3143 2183
rect 3147 2179 3148 2183
rect 3142 2178 3148 2179
rect 1975 2110 1979 2111
rect 1975 2105 1979 2106
rect 1995 2110 1999 2111
rect 1995 2105 1999 2106
rect 2163 2110 2167 2111
rect 2163 2105 2167 2106
rect 2331 2110 2335 2111
rect 2331 2105 2335 2106
rect 2507 2110 2511 2111
rect 2507 2105 2511 2106
rect 2683 2110 2687 2111
rect 2683 2105 2687 2106
rect 2851 2110 2855 2111
rect 2851 2105 2855 2106
rect 3019 2110 3023 2111
rect 3019 2105 3023 2106
rect 3107 2110 3111 2111
rect 3107 2105 3111 2106
rect 1934 2104 1940 2105
rect 1934 2100 1935 2104
rect 1939 2100 1940 2104
rect 1934 2099 1940 2100
rect 1814 2088 1820 2089
rect 1814 2084 1815 2088
rect 1819 2084 1820 2088
rect 1814 2083 1820 2084
rect 1934 2087 1940 2088
rect 1934 2083 1935 2087
rect 1939 2083 1940 2087
rect 1816 2055 1818 2083
rect 1934 2082 1940 2083
rect 1936 2055 1938 2082
rect 1815 2054 1819 2055
rect 1815 2049 1819 2050
rect 1935 2054 1939 2055
rect 1935 2049 1939 2050
rect 1816 2025 1818 2049
rect 1936 2026 1938 2049
rect 1976 2045 1978 2105
rect 1974 2044 1980 2045
rect 3108 2044 3110 2105
rect 3144 2096 3146 2178
rect 3180 2111 3182 2188
rect 3240 2144 3242 2294
rect 3300 2292 3302 2353
rect 3394 2339 3400 2340
rect 3394 2335 3395 2339
rect 3399 2335 3400 2339
rect 3394 2334 3400 2335
rect 3298 2291 3304 2292
rect 3298 2287 3299 2291
rect 3303 2287 3304 2291
rect 3298 2286 3304 2287
rect 3326 2276 3332 2277
rect 3326 2272 3327 2276
rect 3331 2272 3332 2276
rect 3326 2271 3332 2272
rect 3328 2239 3330 2271
rect 3327 2238 3331 2239
rect 3327 2233 3331 2234
rect 3367 2238 3371 2239
rect 3367 2233 3371 2234
rect 3368 2209 3370 2233
rect 3366 2208 3372 2209
rect 3366 2204 3367 2208
rect 3371 2204 3372 2208
rect 3366 2203 3372 2204
rect 3338 2193 3344 2194
rect 3338 2189 3339 2193
rect 3343 2189 3344 2193
rect 3338 2188 3344 2189
rect 3238 2143 3244 2144
rect 3238 2139 3239 2143
rect 3243 2139 3244 2143
rect 3238 2138 3244 2139
rect 3340 2111 3342 2188
rect 3396 2184 3398 2334
rect 3484 2292 3486 2353
rect 3536 2344 3538 2418
rect 3652 2359 3654 2428
rect 3798 2427 3804 2428
rect 3746 2383 3752 2384
rect 3746 2379 3747 2383
rect 3751 2379 3752 2383
rect 3746 2378 3752 2379
rect 3651 2358 3655 2359
rect 3651 2353 3655 2354
rect 3534 2343 3540 2344
rect 3534 2339 3535 2343
rect 3539 2339 3540 2343
rect 3534 2338 3540 2339
rect 3652 2292 3654 2353
rect 3658 2339 3664 2340
rect 3658 2335 3659 2339
rect 3663 2335 3664 2339
rect 3658 2334 3664 2335
rect 3660 2300 3662 2334
rect 3748 2300 3750 2378
rect 3800 2359 3802 2427
rect 3858 2425 3864 2426
rect 3838 2424 3844 2425
rect 3822 2423 3828 2424
rect 3822 2419 3823 2423
rect 3827 2419 3828 2423
rect 3838 2420 3839 2424
rect 3843 2420 3844 2424
rect 3858 2421 3859 2425
rect 3863 2421 3864 2425
rect 3858 2420 3864 2421
rect 4058 2425 4064 2426
rect 4058 2421 4059 2425
rect 4063 2421 4064 2425
rect 4058 2420 4064 2421
rect 3838 2419 3844 2420
rect 3822 2418 3828 2419
rect 3824 2376 3826 2418
rect 3822 2375 3828 2376
rect 3822 2371 3823 2375
rect 3827 2371 3828 2375
rect 3822 2370 3828 2371
rect 3799 2358 3803 2359
rect 3799 2353 3803 2354
rect 3658 2299 3664 2300
rect 3658 2295 3659 2299
rect 3663 2295 3664 2299
rect 3658 2294 3664 2295
rect 3746 2299 3752 2300
rect 3746 2295 3747 2299
rect 3751 2295 3752 2299
rect 3746 2294 3752 2295
rect 3800 2293 3802 2353
rect 3840 2347 3842 2419
rect 3860 2347 3862 2420
rect 4022 2415 4028 2416
rect 4022 2411 4023 2415
rect 4027 2411 4028 2415
rect 4022 2410 4028 2411
rect 4024 2376 4026 2410
rect 4022 2375 4028 2376
rect 4022 2371 4023 2375
rect 4027 2371 4028 2375
rect 4022 2370 4028 2371
rect 4060 2347 4062 2420
rect 4180 2416 4182 2562
rect 4332 2520 4334 2581
rect 4394 2527 4400 2528
rect 4394 2523 4395 2527
rect 4399 2523 4400 2527
rect 4394 2522 4400 2523
rect 4330 2519 4336 2520
rect 4330 2515 4331 2519
rect 4335 2515 4336 2519
rect 4330 2514 4336 2515
rect 4358 2504 4364 2505
rect 4358 2500 4359 2504
rect 4363 2500 4364 2504
rect 4358 2499 4364 2500
rect 4360 2471 4362 2499
rect 4327 2470 4331 2471
rect 4327 2465 4331 2466
rect 4359 2470 4363 2471
rect 4359 2465 4363 2466
rect 4328 2441 4330 2465
rect 4326 2440 4332 2441
rect 4326 2436 4327 2440
rect 4331 2436 4332 2440
rect 4326 2435 4332 2436
rect 4298 2425 4304 2426
rect 4298 2421 4299 2425
rect 4303 2421 4304 2425
rect 4298 2420 4304 2421
rect 4178 2415 4184 2416
rect 4178 2411 4179 2415
rect 4183 2411 4184 2415
rect 4178 2410 4184 2411
rect 4300 2347 4302 2420
rect 4396 2376 4398 2522
rect 4580 2520 4582 2581
rect 4640 2572 4642 2638
rect 4796 2587 4798 2648
rect 4832 2628 4834 2746
rect 5664 2745 5666 2805
rect 5662 2744 5668 2745
rect 5662 2740 5663 2744
rect 5667 2740 5668 2744
rect 5662 2739 5668 2740
rect 4838 2728 4844 2729
rect 4838 2724 4839 2728
rect 4843 2724 4844 2728
rect 4838 2723 4844 2724
rect 5662 2727 5668 2728
rect 5662 2723 5663 2727
rect 5667 2723 5668 2727
rect 4840 2699 4842 2723
rect 5662 2722 5668 2723
rect 5664 2699 5666 2722
rect 4839 2698 4843 2699
rect 4839 2693 4843 2694
rect 5111 2698 5115 2699
rect 5111 2693 5115 2694
rect 5399 2698 5403 2699
rect 5399 2693 5403 2694
rect 5663 2698 5667 2699
rect 5663 2693 5667 2694
rect 5112 2669 5114 2693
rect 5400 2669 5402 2693
rect 5664 2670 5666 2693
rect 5662 2669 5668 2670
rect 5110 2668 5116 2669
rect 5110 2664 5111 2668
rect 5115 2664 5116 2668
rect 5110 2663 5116 2664
rect 5398 2668 5404 2669
rect 5398 2664 5399 2668
rect 5403 2664 5404 2668
rect 5662 2665 5663 2669
rect 5667 2665 5668 2669
rect 5662 2664 5668 2665
rect 5398 2663 5404 2664
rect 5082 2653 5088 2654
rect 5082 2649 5083 2653
rect 5087 2649 5088 2653
rect 5082 2648 5088 2649
rect 5370 2653 5376 2654
rect 5370 2649 5371 2653
rect 5375 2649 5376 2653
rect 5370 2648 5376 2649
rect 5662 2652 5668 2653
rect 5662 2648 5663 2652
rect 5667 2648 5668 2652
rect 4974 2643 4980 2644
rect 4974 2639 4975 2643
rect 4979 2639 4980 2643
rect 4974 2638 4980 2639
rect 4830 2627 4836 2628
rect 4830 2623 4831 2627
rect 4835 2623 4836 2627
rect 4830 2622 4836 2623
rect 4976 2604 4978 2638
rect 4890 2603 4896 2604
rect 4890 2599 4891 2603
rect 4895 2599 4896 2603
rect 4890 2598 4896 2599
rect 4974 2603 4980 2604
rect 4974 2599 4975 2603
rect 4979 2599 4980 2603
rect 4974 2598 4980 2599
rect 4795 2586 4799 2587
rect 4795 2581 4799 2582
rect 4827 2586 4831 2587
rect 4827 2581 4831 2582
rect 4638 2571 4644 2572
rect 4638 2567 4639 2571
rect 4643 2567 4644 2571
rect 4638 2566 4644 2567
rect 4828 2520 4830 2581
rect 4892 2528 4894 2598
rect 5084 2587 5086 2648
rect 5266 2643 5272 2644
rect 5266 2639 5267 2643
rect 5271 2639 5272 2643
rect 5266 2638 5272 2639
rect 5268 2604 5270 2638
rect 5266 2603 5272 2604
rect 5266 2599 5267 2603
rect 5271 2599 5272 2603
rect 5266 2598 5272 2599
rect 5372 2587 5374 2648
rect 5662 2647 5668 2648
rect 5418 2643 5424 2644
rect 5418 2639 5419 2643
rect 5423 2639 5424 2643
rect 5418 2638 5424 2639
rect 5075 2586 5079 2587
rect 5075 2581 5079 2582
rect 5083 2586 5087 2587
rect 5083 2581 5087 2582
rect 5323 2586 5327 2587
rect 5323 2581 5327 2582
rect 5371 2586 5375 2587
rect 5371 2581 5375 2582
rect 4890 2527 4896 2528
rect 4890 2523 4891 2527
rect 4895 2523 4896 2527
rect 4890 2522 4896 2523
rect 5076 2520 5078 2581
rect 5170 2567 5176 2568
rect 5170 2563 5171 2567
rect 5175 2563 5176 2567
rect 5170 2562 5176 2563
rect 4578 2519 4584 2520
rect 4578 2515 4579 2519
rect 4583 2515 4584 2519
rect 4578 2514 4584 2515
rect 4826 2519 4832 2520
rect 4826 2515 4827 2519
rect 4831 2515 4832 2519
rect 4826 2514 4832 2515
rect 5074 2519 5080 2520
rect 5074 2515 5075 2519
rect 5079 2515 5080 2519
rect 5074 2514 5080 2515
rect 4606 2504 4612 2505
rect 4606 2500 4607 2504
rect 4611 2500 4612 2504
rect 4606 2499 4612 2500
rect 4854 2504 4860 2505
rect 4854 2500 4855 2504
rect 4859 2500 4860 2504
rect 4854 2499 4860 2500
rect 5102 2504 5108 2505
rect 5102 2500 5103 2504
rect 5107 2500 5108 2504
rect 5102 2499 5108 2500
rect 4608 2471 4610 2499
rect 4856 2471 4858 2499
rect 5104 2471 5106 2499
rect 4583 2470 4587 2471
rect 4583 2465 4587 2466
rect 4607 2470 4611 2471
rect 4607 2465 4611 2466
rect 4847 2470 4851 2471
rect 4847 2465 4851 2466
rect 4855 2470 4859 2471
rect 4855 2465 4859 2466
rect 5103 2470 5107 2471
rect 5103 2465 5107 2466
rect 5119 2470 5123 2471
rect 5119 2465 5123 2466
rect 4584 2441 4586 2465
rect 4848 2441 4850 2465
rect 5120 2441 5122 2465
rect 4582 2440 4588 2441
rect 4582 2436 4583 2440
rect 4587 2436 4588 2440
rect 4582 2435 4588 2436
rect 4846 2440 4852 2441
rect 4846 2436 4847 2440
rect 4851 2436 4852 2440
rect 4846 2435 4852 2436
rect 5118 2440 5124 2441
rect 5118 2436 5119 2440
rect 5123 2436 5124 2440
rect 5118 2435 5124 2436
rect 4554 2425 4560 2426
rect 4554 2421 4555 2425
rect 4559 2421 4560 2425
rect 4554 2420 4560 2421
rect 4818 2425 4824 2426
rect 4818 2421 4819 2425
rect 4823 2421 4824 2425
rect 4818 2420 4824 2421
rect 5090 2425 5096 2426
rect 5090 2421 5091 2425
rect 5095 2421 5096 2425
rect 5090 2420 5096 2421
rect 4394 2375 4400 2376
rect 4394 2371 4395 2375
rect 4399 2371 4400 2375
rect 4394 2370 4400 2371
rect 4556 2347 4558 2420
rect 4682 2415 4688 2416
rect 4682 2411 4683 2415
rect 4687 2411 4688 2415
rect 4682 2410 4688 2411
rect 4684 2376 4686 2410
rect 4682 2375 4688 2376
rect 4682 2371 4683 2375
rect 4687 2371 4688 2375
rect 4682 2370 4688 2371
rect 4820 2347 4822 2420
rect 4890 2415 4896 2416
rect 4890 2411 4891 2415
rect 4895 2411 4896 2415
rect 4890 2410 4896 2411
rect 3839 2346 3843 2347
rect 3839 2341 3843 2342
rect 3859 2346 3863 2347
rect 3859 2341 3863 2342
rect 4059 2346 4063 2347
rect 4059 2341 4063 2342
rect 4299 2346 4303 2347
rect 4299 2341 4303 2342
rect 4443 2346 4447 2347
rect 4443 2341 4447 2342
rect 4555 2346 4559 2347
rect 4555 2341 4559 2342
rect 4611 2346 4615 2347
rect 4611 2341 4615 2342
rect 4787 2346 4791 2347
rect 4787 2341 4791 2342
rect 4819 2346 4823 2347
rect 4819 2341 4823 2342
rect 3798 2292 3804 2293
rect 3482 2291 3488 2292
rect 3482 2287 3483 2291
rect 3487 2287 3488 2291
rect 3482 2286 3488 2287
rect 3650 2291 3656 2292
rect 3650 2287 3651 2291
rect 3655 2287 3656 2291
rect 3798 2288 3799 2292
rect 3803 2288 3804 2292
rect 3798 2287 3804 2288
rect 3650 2286 3656 2287
rect 3840 2281 3842 2341
rect 3838 2280 3844 2281
rect 4444 2280 4446 2341
rect 4612 2280 4614 2341
rect 4618 2327 4624 2328
rect 4618 2323 4619 2327
rect 4623 2323 4624 2327
rect 4618 2322 4624 2323
rect 4620 2288 4622 2322
rect 4618 2287 4624 2288
rect 4618 2283 4619 2287
rect 4623 2283 4624 2287
rect 4618 2282 4624 2283
rect 4788 2280 4790 2341
rect 4892 2336 4894 2410
rect 5092 2347 5094 2420
rect 5172 2416 5174 2562
rect 5324 2520 5326 2581
rect 5420 2572 5422 2638
rect 5664 2587 5666 2647
rect 5663 2586 5667 2587
rect 5663 2581 5667 2582
rect 5418 2571 5424 2572
rect 5418 2567 5419 2571
rect 5423 2567 5424 2571
rect 5418 2566 5424 2567
rect 5446 2527 5452 2528
rect 5446 2523 5447 2527
rect 5451 2523 5452 2527
rect 5446 2522 5452 2523
rect 5322 2519 5328 2520
rect 5322 2515 5323 2519
rect 5327 2515 5328 2519
rect 5322 2514 5328 2515
rect 5350 2504 5356 2505
rect 5350 2500 5351 2504
rect 5355 2500 5356 2504
rect 5350 2499 5356 2500
rect 5352 2471 5354 2499
rect 5351 2470 5355 2471
rect 5351 2465 5355 2466
rect 5399 2470 5403 2471
rect 5399 2465 5403 2466
rect 5400 2441 5402 2465
rect 5398 2440 5404 2441
rect 5398 2436 5399 2440
rect 5403 2436 5404 2440
rect 5398 2435 5404 2436
rect 5370 2425 5376 2426
rect 5370 2421 5371 2425
rect 5375 2421 5376 2425
rect 5370 2420 5376 2421
rect 5170 2415 5176 2416
rect 5170 2411 5171 2415
rect 5175 2411 5176 2415
rect 5170 2410 5176 2411
rect 5098 2375 5104 2376
rect 5098 2371 5099 2375
rect 5103 2371 5104 2375
rect 5098 2370 5104 2371
rect 4963 2346 4967 2347
rect 4963 2341 4967 2342
rect 5091 2346 5095 2347
rect 5091 2341 5095 2342
rect 4890 2335 4896 2336
rect 4890 2331 4891 2335
rect 4895 2331 4896 2335
rect 4890 2330 4896 2331
rect 4794 2327 4800 2328
rect 4794 2323 4795 2327
rect 4799 2323 4800 2327
rect 4794 2322 4800 2323
rect 4796 2288 4798 2322
rect 4794 2287 4800 2288
rect 4794 2283 4795 2287
rect 4799 2283 4800 2287
rect 4794 2282 4800 2283
rect 4902 2287 4908 2288
rect 4902 2283 4903 2287
rect 4907 2283 4908 2287
rect 4902 2282 4908 2283
rect 3510 2276 3516 2277
rect 3510 2272 3511 2276
rect 3515 2272 3516 2276
rect 3510 2271 3516 2272
rect 3678 2276 3684 2277
rect 3838 2276 3839 2280
rect 3843 2276 3844 2280
rect 3678 2272 3679 2276
rect 3683 2272 3684 2276
rect 3678 2271 3684 2272
rect 3798 2275 3804 2276
rect 3838 2275 3844 2276
rect 4442 2279 4448 2280
rect 4442 2275 4443 2279
rect 4447 2275 4448 2279
rect 3798 2271 3799 2275
rect 3803 2271 3804 2275
rect 4442 2274 4448 2275
rect 4610 2279 4616 2280
rect 4610 2275 4611 2279
rect 4615 2275 4616 2279
rect 4610 2274 4616 2275
rect 4786 2279 4792 2280
rect 4786 2275 4787 2279
rect 4791 2275 4792 2279
rect 4786 2274 4792 2275
rect 3512 2239 3514 2271
rect 3680 2239 3682 2271
rect 3798 2270 3804 2271
rect 3800 2239 3802 2270
rect 4470 2264 4476 2265
rect 3838 2263 3844 2264
rect 3838 2259 3839 2263
rect 3843 2259 3844 2263
rect 4470 2260 4471 2264
rect 4475 2260 4476 2264
rect 4470 2259 4476 2260
rect 4638 2264 4644 2265
rect 4638 2260 4639 2264
rect 4643 2260 4644 2264
rect 4638 2259 4644 2260
rect 4814 2264 4820 2265
rect 4814 2260 4815 2264
rect 4819 2260 4820 2264
rect 4814 2259 4820 2260
rect 3838 2258 3844 2259
rect 3511 2238 3515 2239
rect 3511 2233 3515 2234
rect 3535 2238 3539 2239
rect 3535 2233 3539 2234
rect 3679 2238 3683 2239
rect 3679 2233 3683 2234
rect 3799 2238 3803 2239
rect 3799 2233 3803 2234
rect 3536 2209 3538 2233
rect 3680 2209 3682 2233
rect 3800 2210 3802 2233
rect 3840 2223 3842 2258
rect 4472 2223 4474 2259
rect 4640 2223 4642 2259
rect 4816 2223 4818 2259
rect 3839 2222 3843 2223
rect 3839 2217 3843 2218
rect 4471 2222 4475 2223
rect 4471 2217 4475 2218
rect 4543 2222 4547 2223
rect 4543 2217 4547 2218
rect 4639 2222 4643 2223
rect 4639 2217 4643 2218
rect 4719 2222 4723 2223
rect 4719 2217 4723 2218
rect 4815 2222 4819 2223
rect 4815 2217 4819 2218
rect 3798 2209 3804 2210
rect 3534 2208 3540 2209
rect 3534 2204 3535 2208
rect 3539 2204 3540 2208
rect 3534 2203 3540 2204
rect 3678 2208 3684 2209
rect 3678 2204 3679 2208
rect 3683 2204 3684 2208
rect 3798 2205 3799 2209
rect 3803 2205 3804 2209
rect 3798 2204 3804 2205
rect 3678 2203 3684 2204
rect 3840 2194 3842 2217
rect 3506 2193 3512 2194
rect 3506 2189 3507 2193
rect 3511 2189 3512 2193
rect 3506 2188 3512 2189
rect 3650 2193 3656 2194
rect 3838 2193 3844 2194
rect 4544 2193 4546 2217
rect 4720 2193 4722 2217
rect 3650 2189 3651 2193
rect 3655 2189 3656 2193
rect 3650 2188 3656 2189
rect 3798 2192 3804 2193
rect 3798 2188 3799 2192
rect 3803 2188 3804 2192
rect 3838 2189 3839 2193
rect 3843 2189 3844 2193
rect 3838 2188 3844 2189
rect 4542 2192 4548 2193
rect 4542 2188 4543 2192
rect 4547 2188 4548 2192
rect 3394 2183 3400 2184
rect 3394 2179 3395 2183
rect 3399 2179 3400 2183
rect 3394 2178 3400 2179
rect 3478 2183 3484 2184
rect 3478 2179 3479 2183
rect 3483 2179 3484 2183
rect 3478 2178 3484 2179
rect 3480 2144 3482 2178
rect 3478 2143 3484 2144
rect 3478 2139 3479 2143
rect 3483 2139 3484 2143
rect 3478 2138 3484 2139
rect 3508 2111 3510 2188
rect 3652 2111 3654 2188
rect 3798 2187 3804 2188
rect 4542 2187 4548 2188
rect 4718 2192 4724 2193
rect 4718 2188 4719 2192
rect 4723 2188 4724 2192
rect 4718 2187 4724 2188
rect 3746 2143 3752 2144
rect 3746 2139 3747 2143
rect 3751 2139 3752 2143
rect 3746 2138 3752 2139
rect 3179 2110 3183 2111
rect 3179 2105 3183 2106
rect 3243 2110 3247 2111
rect 3243 2105 3247 2106
rect 3339 2110 3343 2111
rect 3339 2105 3343 2106
rect 3379 2110 3383 2111
rect 3379 2105 3383 2106
rect 3507 2110 3511 2111
rect 3507 2105 3511 2106
rect 3515 2110 3519 2111
rect 3515 2105 3519 2106
rect 3651 2110 3655 2111
rect 3651 2105 3655 2106
rect 3142 2095 3148 2096
rect 3142 2091 3143 2095
rect 3147 2091 3148 2095
rect 3142 2090 3148 2091
rect 3244 2044 3246 2105
rect 3250 2091 3256 2092
rect 3250 2087 3251 2091
rect 3255 2087 3256 2091
rect 3250 2086 3256 2087
rect 3252 2052 3254 2086
rect 3250 2051 3256 2052
rect 3250 2047 3251 2051
rect 3255 2047 3256 2051
rect 3250 2046 3256 2047
rect 3380 2044 3382 2105
rect 3386 2091 3392 2092
rect 3386 2087 3387 2091
rect 3391 2087 3392 2091
rect 3386 2086 3392 2087
rect 3388 2052 3390 2086
rect 3386 2051 3392 2052
rect 3386 2047 3387 2051
rect 3391 2047 3392 2051
rect 3386 2046 3392 2047
rect 3466 2051 3472 2052
rect 3466 2047 3467 2051
rect 3471 2047 3472 2051
rect 3466 2046 3472 2047
rect 1974 2040 1975 2044
rect 1979 2040 1980 2044
rect 1974 2039 1980 2040
rect 3106 2043 3112 2044
rect 3106 2039 3107 2043
rect 3111 2039 3112 2043
rect 3106 2038 3112 2039
rect 3242 2043 3248 2044
rect 3242 2039 3243 2043
rect 3247 2039 3248 2043
rect 3242 2038 3248 2039
rect 3378 2043 3384 2044
rect 3378 2039 3379 2043
rect 3383 2039 3384 2043
rect 3378 2038 3384 2039
rect 3134 2028 3140 2029
rect 1974 2027 1980 2028
rect 1934 2025 1940 2026
rect 1814 2024 1820 2025
rect 1814 2020 1815 2024
rect 1819 2020 1820 2024
rect 1934 2021 1935 2025
rect 1939 2021 1940 2025
rect 1974 2023 1975 2027
rect 1979 2023 1980 2027
rect 3134 2024 3135 2028
rect 3139 2024 3140 2028
rect 3134 2023 3140 2024
rect 3270 2028 3276 2029
rect 3270 2024 3271 2028
rect 3275 2024 3276 2028
rect 3270 2023 3276 2024
rect 3406 2028 3412 2029
rect 3406 2024 3407 2028
rect 3411 2024 3412 2028
rect 3406 2023 3412 2024
rect 1974 2022 1980 2023
rect 1934 2020 1940 2021
rect 1814 2019 1820 2020
rect 1934 2008 1940 2009
rect 1934 2004 1935 2008
rect 1939 2004 1940 2008
rect 1934 2003 1940 2004
rect 1794 1999 1800 2000
rect 1794 1995 1795 1999
rect 1799 1995 1800 1999
rect 1794 1994 1800 1995
rect 1882 1959 1888 1960
rect 1882 1955 1883 1959
rect 1887 1955 1888 1959
rect 1882 1954 1888 1955
rect 1379 1938 1383 1939
rect 1379 1933 1383 1934
rect 1515 1938 1519 1939
rect 1515 1933 1519 1934
rect 1555 1938 1559 1939
rect 1555 1933 1559 1934
rect 1651 1938 1655 1939
rect 1651 1933 1655 1934
rect 1787 1938 1791 1939
rect 1787 1933 1791 1934
rect 1358 1923 1364 1924
rect 1358 1919 1359 1923
rect 1363 1919 1364 1923
rect 1358 1918 1364 1919
rect 1556 1872 1558 1933
rect 1562 1919 1568 1920
rect 1562 1915 1563 1919
rect 1567 1915 1568 1919
rect 1562 1914 1568 1915
rect 1564 1880 1566 1914
rect 1562 1879 1568 1880
rect 1562 1875 1563 1879
rect 1567 1875 1568 1879
rect 1562 1874 1568 1875
rect 1642 1879 1648 1880
rect 1642 1875 1643 1879
rect 1647 1875 1648 1879
rect 1642 1874 1648 1875
rect 1298 1871 1304 1872
rect 1298 1867 1299 1871
rect 1303 1867 1304 1871
rect 1298 1866 1304 1867
rect 1554 1871 1560 1872
rect 1554 1867 1555 1871
rect 1559 1867 1560 1871
rect 1554 1866 1560 1867
rect 1326 1856 1332 1857
rect 1326 1852 1327 1856
rect 1331 1852 1332 1856
rect 1326 1851 1332 1852
rect 1582 1856 1588 1857
rect 1582 1852 1583 1856
rect 1587 1852 1588 1856
rect 1582 1851 1588 1852
rect 1328 1819 1330 1851
rect 1584 1819 1586 1851
rect 1191 1818 1195 1819
rect 1191 1813 1195 1814
rect 1327 1818 1331 1819
rect 1327 1813 1331 1814
rect 1383 1818 1387 1819
rect 1383 1813 1387 1814
rect 1575 1818 1579 1819
rect 1575 1813 1579 1814
rect 1583 1818 1587 1819
rect 1583 1813 1587 1814
rect 1192 1789 1194 1813
rect 1384 1789 1386 1813
rect 1576 1789 1578 1813
rect 1190 1788 1196 1789
rect 1190 1784 1191 1788
rect 1195 1784 1196 1788
rect 1190 1783 1196 1784
rect 1382 1788 1388 1789
rect 1382 1784 1383 1788
rect 1387 1784 1388 1788
rect 1382 1783 1388 1784
rect 1574 1788 1580 1789
rect 1574 1784 1575 1788
rect 1579 1784 1580 1788
rect 1574 1783 1580 1784
rect 1162 1773 1168 1774
rect 1162 1769 1163 1773
rect 1167 1769 1168 1773
rect 1162 1768 1168 1769
rect 1354 1773 1360 1774
rect 1354 1769 1355 1773
rect 1359 1769 1360 1773
rect 1354 1768 1360 1769
rect 1546 1773 1552 1774
rect 1546 1769 1547 1773
rect 1551 1769 1552 1773
rect 1546 1768 1552 1769
rect 1134 1715 1140 1716
rect 1134 1711 1135 1715
rect 1139 1711 1140 1715
rect 1134 1710 1140 1711
rect 1164 1683 1166 1768
rect 1286 1763 1292 1764
rect 1286 1759 1287 1763
rect 1291 1759 1292 1763
rect 1286 1758 1292 1759
rect 563 1682 567 1683
rect 563 1677 567 1678
rect 683 1682 687 1683
rect 683 1677 687 1678
rect 771 1682 775 1683
rect 771 1677 775 1678
rect 971 1682 975 1683
rect 971 1677 975 1678
rect 979 1682 983 1683
rect 979 1677 983 1678
rect 1163 1682 1167 1683
rect 1163 1677 1167 1678
rect 1275 1682 1279 1683
rect 1275 1677 1279 1678
rect 490 1667 496 1668
rect 490 1663 491 1667
rect 495 1663 496 1667
rect 490 1662 496 1663
rect 684 1616 686 1677
rect 690 1663 696 1664
rect 690 1659 691 1663
rect 695 1659 696 1663
rect 690 1658 696 1659
rect 692 1624 694 1658
rect 690 1623 696 1624
rect 690 1619 691 1623
rect 695 1619 696 1623
rect 690 1618 696 1619
rect 980 1616 982 1677
rect 1074 1663 1080 1664
rect 1074 1659 1075 1663
rect 1079 1659 1080 1663
rect 1074 1658 1080 1659
rect 1076 1636 1078 1658
rect 1074 1635 1080 1636
rect 1074 1631 1075 1635
rect 1079 1631 1080 1635
rect 1074 1630 1080 1631
rect 986 1623 992 1624
rect 986 1619 987 1623
rect 991 1619 992 1623
rect 986 1618 992 1619
rect 994 1623 1000 1624
rect 994 1619 995 1623
rect 999 1619 1000 1623
rect 994 1618 1000 1619
rect 394 1615 400 1616
rect 394 1611 395 1615
rect 399 1611 400 1615
rect 394 1610 400 1611
rect 682 1615 688 1616
rect 682 1611 683 1615
rect 687 1611 688 1615
rect 682 1610 688 1611
rect 978 1615 984 1616
rect 978 1611 979 1615
rect 983 1611 984 1615
rect 978 1610 984 1611
rect 422 1600 428 1601
rect 422 1596 423 1600
rect 427 1596 428 1600
rect 422 1595 428 1596
rect 710 1600 716 1601
rect 710 1596 711 1600
rect 715 1596 716 1600
rect 710 1595 716 1596
rect 424 1559 426 1595
rect 712 1559 714 1595
rect 375 1558 379 1559
rect 375 1553 379 1554
rect 423 1558 427 1559
rect 423 1553 427 1554
rect 607 1558 611 1559
rect 607 1553 611 1554
rect 711 1558 715 1559
rect 711 1553 715 1554
rect 839 1558 843 1559
rect 839 1553 843 1554
rect 376 1529 378 1553
rect 608 1529 610 1553
rect 840 1529 842 1553
rect 374 1528 380 1529
rect 374 1524 375 1528
rect 379 1524 380 1528
rect 374 1523 380 1524
rect 606 1528 612 1529
rect 606 1524 607 1528
rect 611 1524 612 1528
rect 606 1523 612 1524
rect 838 1528 844 1529
rect 838 1524 839 1528
rect 843 1524 844 1528
rect 838 1523 844 1524
rect 346 1513 352 1514
rect 346 1509 347 1513
rect 351 1509 352 1513
rect 346 1508 352 1509
rect 578 1513 584 1514
rect 578 1509 579 1513
rect 583 1509 584 1513
rect 578 1508 584 1509
rect 810 1513 816 1514
rect 810 1509 811 1513
rect 815 1509 816 1513
rect 810 1508 816 1509
rect 238 1503 244 1504
rect 238 1499 239 1503
rect 243 1499 244 1503
rect 238 1498 244 1499
rect 348 1435 350 1508
rect 354 1503 360 1504
rect 354 1499 355 1503
rect 359 1499 360 1503
rect 354 1498 360 1499
rect 356 1472 358 1498
rect 354 1471 360 1472
rect 354 1467 355 1471
rect 359 1467 360 1471
rect 354 1466 360 1467
rect 580 1435 582 1508
rect 718 1503 724 1504
rect 718 1499 719 1503
rect 723 1499 724 1503
rect 718 1498 724 1499
rect 802 1503 808 1504
rect 802 1499 803 1503
rect 807 1499 808 1503
rect 802 1498 808 1499
rect 111 1434 115 1435
rect 111 1429 115 1430
rect 131 1434 135 1435
rect 131 1429 135 1430
rect 347 1434 351 1435
rect 347 1429 351 1430
rect 411 1434 415 1435
rect 411 1429 415 1430
rect 579 1434 583 1435
rect 579 1429 583 1430
rect 112 1369 114 1429
rect 110 1368 116 1369
rect 132 1368 134 1429
rect 226 1415 232 1416
rect 226 1411 227 1415
rect 231 1411 232 1415
rect 226 1410 232 1411
rect 110 1364 111 1368
rect 115 1364 116 1368
rect 110 1363 116 1364
rect 130 1367 136 1368
rect 130 1363 131 1367
rect 135 1363 136 1367
rect 130 1362 136 1363
rect 158 1352 164 1353
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 158 1348 159 1352
rect 163 1348 164 1352
rect 158 1347 164 1348
rect 110 1346 116 1347
rect 112 1323 114 1346
rect 160 1323 162 1347
rect 111 1322 115 1323
rect 111 1317 115 1318
rect 159 1322 163 1323
rect 159 1317 163 1318
rect 112 1294 114 1317
rect 110 1293 116 1294
rect 160 1293 162 1317
rect 110 1289 111 1293
rect 115 1289 116 1293
rect 110 1288 116 1289
rect 158 1292 164 1293
rect 158 1288 159 1292
rect 163 1288 164 1292
rect 158 1287 164 1288
rect 130 1277 136 1278
rect 110 1276 116 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 130 1273 131 1277
rect 135 1273 136 1277
rect 130 1272 136 1273
rect 110 1271 116 1272
rect 112 1199 114 1271
rect 132 1199 134 1272
rect 228 1268 230 1410
rect 412 1368 414 1429
rect 720 1420 722 1498
rect 804 1464 806 1498
rect 802 1463 808 1464
rect 802 1459 803 1463
rect 807 1459 808 1463
rect 802 1458 808 1459
rect 812 1435 814 1508
rect 988 1464 990 1618
rect 996 1472 998 1618
rect 1276 1616 1278 1677
rect 1288 1668 1290 1758
rect 1356 1683 1358 1768
rect 1548 1683 1550 1768
rect 1644 1724 1646 1874
rect 1788 1872 1790 1933
rect 1884 1880 1886 1954
rect 1936 1939 1938 2003
rect 1976 1999 1978 2022
rect 3136 1999 3138 2023
rect 3272 1999 3274 2023
rect 3408 1999 3410 2023
rect 1975 1998 1979 1999
rect 1975 1993 1979 1994
rect 3127 1998 3131 1999
rect 3127 1993 3131 1994
rect 3135 1998 3139 1999
rect 3135 1993 3139 1994
rect 3263 1998 3267 1999
rect 3263 1993 3267 1994
rect 3271 1998 3275 1999
rect 3271 1993 3275 1994
rect 3399 1998 3403 1999
rect 3399 1993 3403 1994
rect 3407 1998 3411 1999
rect 3407 1993 3411 1994
rect 1976 1970 1978 1993
rect 1974 1969 1980 1970
rect 3128 1969 3130 1993
rect 3264 1969 3266 1993
rect 3400 1969 3402 1993
rect 1974 1965 1975 1969
rect 1979 1965 1980 1969
rect 1974 1964 1980 1965
rect 3126 1968 3132 1969
rect 3126 1964 3127 1968
rect 3131 1964 3132 1968
rect 3126 1963 3132 1964
rect 3262 1968 3268 1969
rect 3262 1964 3263 1968
rect 3267 1964 3268 1968
rect 3262 1963 3268 1964
rect 3398 1968 3404 1969
rect 3398 1964 3399 1968
rect 3403 1964 3404 1968
rect 3398 1963 3404 1964
rect 3098 1953 3104 1954
rect 1974 1952 1980 1953
rect 1974 1948 1975 1952
rect 1979 1948 1980 1952
rect 3098 1949 3099 1953
rect 3103 1949 3104 1953
rect 3098 1948 3104 1949
rect 3234 1953 3240 1954
rect 3234 1949 3235 1953
rect 3239 1949 3240 1953
rect 3234 1948 3240 1949
rect 3370 1953 3376 1954
rect 3370 1949 3371 1953
rect 3375 1949 3376 1953
rect 3370 1948 3376 1949
rect 1974 1947 1980 1948
rect 1935 1938 1939 1939
rect 1935 1933 1939 1934
rect 1882 1879 1888 1880
rect 1882 1875 1883 1879
rect 1887 1875 1888 1879
rect 1882 1874 1888 1875
rect 1936 1873 1938 1933
rect 1976 1875 1978 1947
rect 2118 1923 2124 1924
rect 2118 1919 2119 1923
rect 2123 1919 2124 1923
rect 2118 1918 2124 1919
rect 1975 1874 1979 1875
rect 1934 1872 1940 1873
rect 1786 1871 1792 1872
rect 1786 1867 1787 1871
rect 1791 1867 1792 1871
rect 1934 1868 1935 1872
rect 1939 1868 1940 1872
rect 1975 1869 1979 1870
rect 1995 1874 1999 1875
rect 1995 1869 1999 1870
rect 1934 1867 1940 1868
rect 1786 1866 1792 1867
rect 1814 1856 1820 1857
rect 1814 1852 1815 1856
rect 1819 1852 1820 1856
rect 1814 1851 1820 1852
rect 1934 1855 1940 1856
rect 1934 1851 1935 1855
rect 1939 1851 1940 1855
rect 1816 1819 1818 1851
rect 1934 1850 1940 1851
rect 1936 1819 1938 1850
rect 1815 1818 1819 1819
rect 1815 1813 1819 1814
rect 1935 1818 1939 1819
rect 1935 1813 1939 1814
rect 1936 1790 1938 1813
rect 1976 1809 1978 1869
rect 1974 1808 1980 1809
rect 1996 1808 1998 1869
rect 2120 1816 2122 1918
rect 3100 1875 3102 1948
rect 3202 1943 3208 1944
rect 3202 1939 3203 1943
rect 3207 1939 3208 1943
rect 3202 1938 3208 1939
rect 2227 1874 2231 1875
rect 2227 1869 2231 1870
rect 2467 1874 2471 1875
rect 2467 1869 2471 1870
rect 2691 1874 2695 1875
rect 2691 1869 2695 1870
rect 2907 1874 2911 1875
rect 2907 1869 2911 1870
rect 3099 1874 3103 1875
rect 3099 1869 3103 1870
rect 3107 1874 3111 1875
rect 3107 1869 3111 1870
rect 2218 1859 2224 1860
rect 2218 1855 2219 1859
rect 2223 1855 2224 1859
rect 2218 1854 2224 1855
rect 2220 1816 2222 1854
rect 2118 1815 2124 1816
rect 2118 1811 2119 1815
rect 2123 1811 2124 1815
rect 2118 1810 2124 1811
rect 2218 1815 2224 1816
rect 2218 1811 2219 1815
rect 2223 1811 2224 1815
rect 2218 1810 2224 1811
rect 2228 1808 2230 1869
rect 2402 1859 2408 1860
rect 2402 1855 2403 1859
rect 2407 1855 2408 1859
rect 2402 1854 2408 1855
rect 2410 1859 2416 1860
rect 2410 1855 2411 1859
rect 2415 1855 2416 1859
rect 2410 1854 2416 1855
rect 2404 1816 2406 1854
rect 2402 1815 2408 1816
rect 2402 1811 2403 1815
rect 2407 1811 2408 1815
rect 2402 1810 2408 1811
rect 1974 1804 1975 1808
rect 1979 1804 1980 1808
rect 1974 1803 1980 1804
rect 1994 1807 2000 1808
rect 1994 1803 1995 1807
rect 1999 1803 2000 1807
rect 1994 1802 2000 1803
rect 2226 1807 2232 1808
rect 2226 1803 2227 1807
rect 2231 1803 2232 1807
rect 2226 1802 2232 1803
rect 2022 1792 2028 1793
rect 1974 1791 1980 1792
rect 1934 1789 1940 1790
rect 1934 1785 1935 1789
rect 1939 1785 1940 1789
rect 1974 1787 1975 1791
rect 1979 1787 1980 1791
rect 2022 1788 2023 1792
rect 2027 1788 2028 1792
rect 2022 1787 2028 1788
rect 2254 1792 2260 1793
rect 2254 1788 2255 1792
rect 2259 1788 2260 1792
rect 2254 1787 2260 1788
rect 1974 1786 1980 1787
rect 1934 1784 1940 1785
rect 1934 1772 1940 1773
rect 1934 1768 1935 1772
rect 1939 1768 1940 1772
rect 1934 1767 1940 1768
rect 1642 1723 1648 1724
rect 1642 1719 1643 1723
rect 1647 1719 1648 1723
rect 1642 1718 1648 1719
rect 1936 1683 1938 1767
rect 1976 1755 1978 1786
rect 2024 1755 2026 1787
rect 2256 1755 2258 1787
rect 1975 1754 1979 1755
rect 1975 1749 1979 1750
rect 2023 1754 2027 1755
rect 2023 1749 2027 1750
rect 2159 1754 2163 1755
rect 2159 1749 2163 1750
rect 2255 1754 2259 1755
rect 2255 1749 2259 1750
rect 2311 1754 2315 1755
rect 2311 1749 2315 1750
rect 1976 1726 1978 1749
rect 1974 1725 1980 1726
rect 2024 1725 2026 1749
rect 2160 1725 2162 1749
rect 2312 1725 2314 1749
rect 1974 1721 1975 1725
rect 1979 1721 1980 1725
rect 1974 1720 1980 1721
rect 2022 1724 2028 1725
rect 2022 1720 2023 1724
rect 2027 1720 2028 1724
rect 2022 1719 2028 1720
rect 2158 1724 2164 1725
rect 2158 1720 2159 1724
rect 2163 1720 2164 1724
rect 2158 1719 2164 1720
rect 2310 1724 2316 1725
rect 2310 1720 2311 1724
rect 2315 1720 2316 1724
rect 2310 1719 2316 1720
rect 1994 1709 2000 1710
rect 1974 1708 1980 1709
rect 1974 1704 1975 1708
rect 1979 1704 1980 1708
rect 1994 1705 1995 1709
rect 1999 1705 2000 1709
rect 1994 1704 2000 1705
rect 2130 1709 2136 1710
rect 2130 1705 2131 1709
rect 2135 1705 2136 1709
rect 2130 1704 2136 1705
rect 2282 1709 2288 1710
rect 2282 1705 2283 1709
rect 2287 1705 2288 1709
rect 2282 1704 2288 1705
rect 1974 1703 1980 1704
rect 1355 1682 1359 1683
rect 1355 1677 1359 1678
rect 1547 1682 1551 1683
rect 1547 1677 1551 1678
rect 1935 1682 1939 1683
rect 1935 1677 1939 1678
rect 1286 1667 1292 1668
rect 1286 1663 1287 1667
rect 1291 1663 1292 1667
rect 1286 1662 1292 1663
rect 1936 1617 1938 1677
rect 1976 1635 1978 1703
rect 1996 1635 1998 1704
rect 2122 1699 2128 1700
rect 2122 1695 2123 1699
rect 2127 1695 2128 1699
rect 2122 1694 2128 1695
rect 2090 1691 2096 1692
rect 2090 1687 2091 1691
rect 2095 1687 2096 1691
rect 2090 1686 2096 1687
rect 2092 1660 2094 1686
rect 2124 1660 2126 1694
rect 2090 1659 2096 1660
rect 2090 1655 2091 1659
rect 2095 1655 2096 1659
rect 2090 1654 2096 1655
rect 2122 1659 2128 1660
rect 2122 1655 2123 1659
rect 2127 1655 2128 1659
rect 2122 1654 2128 1655
rect 2132 1635 2134 1704
rect 2258 1699 2264 1700
rect 2258 1695 2259 1699
rect 2263 1695 2264 1699
rect 2258 1694 2264 1695
rect 2260 1660 2262 1694
rect 2258 1659 2264 1660
rect 2258 1655 2259 1659
rect 2263 1655 2264 1659
rect 2258 1654 2264 1655
rect 2284 1635 2286 1704
rect 2412 1700 2414 1854
rect 2468 1808 2470 1869
rect 2692 1808 2694 1869
rect 2786 1855 2792 1856
rect 2786 1851 2787 1855
rect 2791 1851 2792 1855
rect 2786 1850 2792 1851
rect 2788 1824 2790 1850
rect 2786 1823 2792 1824
rect 2786 1819 2787 1823
rect 2791 1819 2792 1823
rect 2786 1818 2792 1819
rect 2908 1808 2910 1869
rect 2914 1855 2920 1856
rect 2914 1851 2915 1855
rect 2919 1851 2920 1855
rect 2914 1850 2920 1851
rect 2916 1816 2918 1850
rect 2914 1815 2920 1816
rect 2914 1811 2915 1815
rect 2919 1811 2920 1815
rect 2914 1810 2920 1811
rect 3030 1815 3036 1816
rect 3030 1811 3031 1815
rect 3035 1811 3036 1815
rect 3030 1810 3036 1811
rect 2466 1807 2472 1808
rect 2466 1803 2467 1807
rect 2471 1803 2472 1807
rect 2466 1802 2472 1803
rect 2690 1807 2696 1808
rect 2690 1803 2691 1807
rect 2695 1803 2696 1807
rect 2690 1802 2696 1803
rect 2906 1807 2912 1808
rect 2906 1803 2907 1807
rect 2911 1803 2912 1807
rect 2906 1802 2912 1803
rect 2494 1792 2500 1793
rect 2494 1788 2495 1792
rect 2499 1788 2500 1792
rect 2494 1787 2500 1788
rect 2718 1792 2724 1793
rect 2718 1788 2719 1792
rect 2723 1788 2724 1792
rect 2718 1787 2724 1788
rect 2934 1792 2940 1793
rect 2934 1788 2935 1792
rect 2939 1788 2940 1792
rect 2934 1787 2940 1788
rect 2496 1755 2498 1787
rect 2720 1755 2722 1787
rect 2936 1755 2938 1787
rect 2471 1754 2475 1755
rect 2471 1749 2475 1750
rect 2495 1754 2499 1755
rect 2495 1749 2499 1750
rect 2639 1754 2643 1755
rect 2639 1749 2643 1750
rect 2719 1754 2723 1755
rect 2719 1749 2723 1750
rect 2807 1754 2811 1755
rect 2807 1749 2811 1750
rect 2935 1754 2939 1755
rect 2935 1749 2939 1750
rect 2975 1754 2979 1755
rect 2975 1749 2979 1750
rect 2472 1725 2474 1749
rect 2640 1725 2642 1749
rect 2808 1725 2810 1749
rect 2976 1725 2978 1749
rect 2470 1724 2476 1725
rect 2470 1720 2471 1724
rect 2475 1720 2476 1724
rect 2470 1719 2476 1720
rect 2638 1724 2644 1725
rect 2638 1720 2639 1724
rect 2643 1720 2644 1724
rect 2638 1719 2644 1720
rect 2806 1724 2812 1725
rect 2806 1720 2807 1724
rect 2811 1720 2812 1724
rect 2806 1719 2812 1720
rect 2974 1724 2980 1725
rect 2974 1720 2975 1724
rect 2979 1720 2980 1724
rect 2974 1719 2980 1720
rect 2442 1709 2448 1710
rect 2442 1705 2443 1709
rect 2447 1705 2448 1709
rect 2442 1704 2448 1705
rect 2610 1709 2616 1710
rect 2610 1705 2611 1709
rect 2615 1705 2616 1709
rect 2610 1704 2616 1705
rect 2778 1709 2784 1710
rect 2778 1705 2779 1709
rect 2783 1705 2784 1709
rect 2778 1704 2784 1705
rect 2946 1709 2952 1710
rect 2946 1705 2947 1709
rect 2951 1705 2952 1709
rect 2946 1704 2952 1705
rect 2410 1699 2416 1700
rect 2410 1695 2411 1699
rect 2415 1695 2416 1699
rect 2410 1694 2416 1695
rect 2444 1635 2446 1704
rect 2602 1699 2608 1700
rect 2602 1695 2603 1699
rect 2607 1695 2608 1699
rect 2602 1694 2608 1695
rect 2604 1660 2606 1694
rect 2602 1659 2608 1660
rect 2602 1655 2603 1659
rect 2607 1655 2608 1659
rect 2602 1654 2608 1655
rect 2612 1635 2614 1704
rect 2706 1659 2712 1660
rect 2706 1655 2707 1659
rect 2711 1655 2712 1659
rect 2706 1654 2712 1655
rect 1975 1634 1979 1635
rect 1975 1629 1979 1630
rect 1995 1634 1999 1635
rect 1995 1629 1999 1630
rect 2091 1634 2095 1635
rect 2091 1629 2095 1630
rect 2131 1634 2135 1635
rect 2131 1629 2135 1630
rect 2227 1634 2231 1635
rect 2227 1629 2231 1630
rect 2283 1634 2287 1635
rect 2283 1629 2287 1630
rect 2363 1634 2367 1635
rect 2363 1629 2367 1630
rect 2443 1634 2447 1635
rect 2443 1629 2447 1630
rect 2499 1634 2503 1635
rect 2499 1629 2503 1630
rect 2611 1634 2615 1635
rect 2611 1629 2615 1630
rect 2635 1634 2639 1635
rect 2635 1629 2639 1630
rect 1934 1616 1940 1617
rect 1274 1615 1280 1616
rect 1274 1611 1275 1615
rect 1279 1611 1280 1615
rect 1934 1612 1935 1616
rect 1939 1612 1940 1616
rect 1934 1611 1940 1612
rect 1274 1610 1280 1611
rect 1006 1600 1012 1601
rect 1006 1596 1007 1600
rect 1011 1596 1012 1600
rect 1006 1595 1012 1596
rect 1302 1600 1308 1601
rect 1302 1596 1303 1600
rect 1307 1596 1308 1600
rect 1302 1595 1308 1596
rect 1934 1599 1940 1600
rect 1934 1595 1935 1599
rect 1939 1595 1940 1599
rect 1008 1559 1010 1595
rect 1304 1559 1306 1595
rect 1934 1594 1940 1595
rect 1936 1559 1938 1594
rect 1976 1569 1978 1629
rect 1974 1568 1980 1569
rect 2092 1568 2094 1629
rect 2186 1615 2192 1616
rect 2186 1611 2187 1615
rect 2191 1611 2192 1615
rect 2186 1610 2192 1611
rect 1974 1564 1975 1568
rect 1979 1564 1980 1568
rect 1974 1563 1980 1564
rect 2090 1567 2096 1568
rect 2090 1563 2091 1567
rect 2095 1563 2096 1567
rect 2090 1562 2096 1563
rect 1007 1558 1011 1559
rect 1007 1553 1011 1554
rect 1071 1558 1075 1559
rect 1071 1553 1075 1554
rect 1303 1558 1307 1559
rect 1303 1553 1307 1554
rect 1935 1558 1939 1559
rect 1935 1553 1939 1554
rect 1072 1529 1074 1553
rect 1304 1529 1306 1553
rect 1936 1530 1938 1553
rect 2118 1552 2124 1553
rect 1974 1551 1980 1552
rect 1974 1547 1975 1551
rect 1979 1547 1980 1551
rect 2118 1548 2119 1552
rect 2123 1548 2124 1552
rect 2118 1547 2124 1548
rect 1974 1546 1980 1547
rect 1934 1529 1940 1530
rect 1070 1528 1076 1529
rect 1070 1524 1071 1528
rect 1075 1524 1076 1528
rect 1070 1523 1076 1524
rect 1302 1528 1308 1529
rect 1302 1524 1303 1528
rect 1307 1524 1308 1528
rect 1934 1525 1935 1529
rect 1939 1525 1940 1529
rect 1934 1524 1940 1525
rect 1302 1523 1308 1524
rect 1042 1513 1048 1514
rect 1042 1509 1043 1513
rect 1047 1509 1048 1513
rect 1042 1508 1048 1509
rect 1274 1513 1280 1514
rect 1274 1509 1275 1513
rect 1279 1509 1280 1513
rect 1274 1508 1280 1509
rect 1934 1512 1940 1513
rect 1934 1508 1935 1512
rect 1939 1508 1940 1512
rect 994 1471 1000 1472
rect 994 1467 995 1471
rect 999 1467 1000 1471
rect 994 1466 1000 1467
rect 986 1463 992 1464
rect 986 1459 987 1463
rect 991 1459 992 1463
rect 986 1458 992 1459
rect 1044 1435 1046 1508
rect 1170 1503 1176 1504
rect 1170 1499 1171 1503
rect 1175 1499 1176 1503
rect 1170 1498 1176 1499
rect 1172 1464 1174 1498
rect 1170 1463 1176 1464
rect 1170 1459 1171 1463
rect 1175 1459 1176 1463
rect 1170 1458 1176 1459
rect 1276 1435 1278 1508
rect 1934 1507 1940 1508
rect 1402 1503 1408 1504
rect 1402 1499 1403 1503
rect 1407 1499 1408 1503
rect 1402 1498 1408 1499
rect 739 1434 743 1435
rect 739 1429 743 1430
rect 811 1434 815 1435
rect 811 1429 815 1430
rect 1043 1434 1047 1435
rect 1043 1429 1047 1430
rect 1091 1434 1095 1435
rect 1091 1429 1095 1430
rect 1275 1434 1279 1435
rect 1275 1429 1279 1430
rect 718 1419 724 1420
rect 506 1415 512 1416
rect 506 1411 507 1415
rect 511 1411 512 1415
rect 718 1415 719 1419
rect 723 1415 724 1419
rect 718 1414 724 1415
rect 506 1410 512 1411
rect 508 1396 510 1410
rect 506 1395 512 1396
rect 506 1391 507 1395
rect 511 1391 512 1395
rect 506 1390 512 1391
rect 740 1368 742 1429
rect 862 1395 868 1396
rect 862 1391 863 1395
rect 867 1391 868 1395
rect 862 1390 868 1391
rect 864 1376 866 1390
rect 862 1375 868 1376
rect 862 1371 863 1375
rect 867 1371 868 1375
rect 862 1370 868 1371
rect 1034 1375 1040 1376
rect 1034 1371 1035 1375
rect 1039 1371 1040 1375
rect 1034 1370 1040 1371
rect 410 1367 416 1368
rect 410 1363 411 1367
rect 415 1363 416 1367
rect 410 1362 416 1363
rect 738 1367 744 1368
rect 738 1363 739 1367
rect 743 1363 744 1367
rect 738 1362 744 1363
rect 438 1352 444 1353
rect 438 1348 439 1352
rect 443 1348 444 1352
rect 438 1347 444 1348
rect 766 1352 772 1353
rect 766 1348 767 1352
rect 771 1348 772 1352
rect 766 1347 772 1348
rect 440 1323 442 1347
rect 768 1323 770 1347
rect 359 1322 363 1323
rect 359 1317 363 1318
rect 439 1322 443 1323
rect 439 1317 443 1318
rect 575 1322 579 1323
rect 575 1317 579 1318
rect 767 1322 771 1323
rect 767 1317 771 1318
rect 775 1322 779 1323
rect 775 1317 779 1318
rect 967 1322 971 1323
rect 967 1317 971 1318
rect 360 1293 362 1317
rect 576 1293 578 1317
rect 776 1293 778 1317
rect 968 1293 970 1317
rect 358 1292 364 1293
rect 358 1288 359 1292
rect 363 1288 364 1292
rect 358 1287 364 1288
rect 574 1292 580 1293
rect 574 1288 575 1292
rect 579 1288 580 1292
rect 574 1287 580 1288
rect 774 1292 780 1293
rect 774 1288 775 1292
rect 779 1288 780 1292
rect 774 1287 780 1288
rect 966 1292 972 1293
rect 966 1288 967 1292
rect 971 1288 972 1292
rect 966 1287 972 1288
rect 330 1277 336 1278
rect 330 1273 331 1277
rect 335 1273 336 1277
rect 330 1272 336 1273
rect 546 1277 552 1278
rect 546 1273 547 1277
rect 551 1273 552 1277
rect 546 1272 552 1273
rect 746 1277 752 1278
rect 746 1273 747 1277
rect 751 1273 752 1277
rect 746 1272 752 1273
rect 938 1277 944 1278
rect 938 1273 939 1277
rect 943 1273 944 1277
rect 938 1272 944 1273
rect 226 1267 232 1268
rect 226 1263 227 1267
rect 231 1263 232 1267
rect 226 1262 232 1263
rect 226 1227 232 1228
rect 226 1223 227 1227
rect 231 1223 232 1227
rect 226 1222 232 1223
rect 111 1198 115 1199
rect 111 1193 115 1194
rect 131 1198 135 1199
rect 131 1193 135 1194
rect 112 1133 114 1193
rect 110 1132 116 1133
rect 132 1132 134 1193
rect 228 1140 230 1222
rect 332 1199 334 1272
rect 386 1267 392 1268
rect 386 1263 387 1267
rect 391 1263 392 1267
rect 386 1262 392 1263
rect 291 1198 295 1199
rect 291 1193 295 1194
rect 331 1198 335 1199
rect 331 1193 335 1194
rect 270 1183 276 1184
rect 270 1179 271 1183
rect 275 1179 276 1183
rect 270 1178 276 1179
rect 226 1139 232 1140
rect 226 1135 227 1139
rect 231 1135 232 1139
rect 226 1134 232 1135
rect 110 1128 111 1132
rect 115 1128 116 1132
rect 110 1127 116 1128
rect 130 1131 136 1132
rect 130 1127 131 1131
rect 135 1127 136 1131
rect 130 1126 136 1127
rect 158 1116 164 1117
rect 110 1115 116 1116
rect 110 1111 111 1115
rect 115 1111 116 1115
rect 158 1112 159 1116
rect 163 1112 164 1116
rect 158 1111 164 1112
rect 110 1110 116 1111
rect 112 1075 114 1110
rect 160 1075 162 1111
rect 111 1074 115 1075
rect 111 1069 115 1070
rect 159 1074 163 1075
rect 159 1069 163 1070
rect 175 1074 179 1075
rect 175 1069 179 1070
rect 112 1046 114 1069
rect 110 1045 116 1046
rect 176 1045 178 1069
rect 110 1041 111 1045
rect 115 1041 116 1045
rect 110 1040 116 1041
rect 174 1044 180 1045
rect 174 1040 175 1044
rect 179 1040 180 1044
rect 174 1039 180 1040
rect 146 1029 152 1030
rect 110 1028 116 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 146 1025 147 1029
rect 151 1025 152 1029
rect 146 1024 152 1025
rect 110 1023 116 1024
rect 112 951 114 1023
rect 148 951 150 1024
rect 272 1020 274 1178
rect 292 1132 294 1193
rect 388 1184 390 1262
rect 548 1199 550 1272
rect 748 1199 750 1272
rect 870 1267 876 1268
rect 870 1263 871 1267
rect 875 1263 876 1267
rect 870 1262 876 1263
rect 475 1198 479 1199
rect 475 1193 479 1194
rect 547 1198 551 1199
rect 547 1193 551 1194
rect 659 1198 663 1199
rect 659 1193 663 1194
rect 747 1198 751 1199
rect 747 1193 751 1194
rect 835 1198 839 1199
rect 835 1193 839 1194
rect 386 1183 392 1184
rect 386 1179 387 1183
rect 391 1179 392 1183
rect 386 1178 392 1179
rect 476 1132 478 1193
rect 482 1179 488 1180
rect 482 1175 483 1179
rect 487 1175 488 1179
rect 482 1174 488 1175
rect 484 1140 486 1174
rect 482 1139 488 1140
rect 482 1135 483 1139
rect 487 1135 488 1139
rect 482 1134 488 1135
rect 660 1132 662 1193
rect 666 1179 672 1180
rect 666 1175 667 1179
rect 671 1175 672 1179
rect 666 1174 672 1175
rect 668 1140 670 1174
rect 666 1139 672 1140
rect 666 1135 667 1139
rect 671 1135 672 1139
rect 666 1134 672 1135
rect 754 1139 760 1140
rect 754 1135 755 1139
rect 759 1135 760 1139
rect 754 1134 760 1135
rect 290 1131 296 1132
rect 290 1127 291 1131
rect 295 1127 296 1131
rect 290 1126 296 1127
rect 474 1131 480 1132
rect 474 1127 475 1131
rect 479 1127 480 1131
rect 474 1126 480 1127
rect 658 1131 664 1132
rect 658 1127 659 1131
rect 663 1127 664 1131
rect 658 1126 664 1127
rect 318 1116 324 1117
rect 318 1112 319 1116
rect 323 1112 324 1116
rect 318 1111 324 1112
rect 502 1116 508 1117
rect 502 1112 503 1116
rect 507 1112 508 1116
rect 502 1111 508 1112
rect 686 1116 692 1117
rect 686 1112 687 1116
rect 691 1112 692 1116
rect 686 1111 692 1112
rect 320 1075 322 1111
rect 504 1075 506 1111
rect 688 1075 690 1111
rect 319 1074 323 1075
rect 319 1069 323 1070
rect 431 1074 435 1075
rect 431 1069 435 1070
rect 503 1074 507 1075
rect 503 1069 507 1070
rect 687 1074 691 1075
rect 687 1069 691 1070
rect 432 1045 434 1069
rect 688 1045 690 1069
rect 430 1044 436 1045
rect 430 1040 431 1044
rect 435 1040 436 1044
rect 430 1039 436 1040
rect 686 1044 692 1045
rect 686 1040 687 1044
rect 691 1040 692 1044
rect 686 1039 692 1040
rect 402 1029 408 1030
rect 402 1025 403 1029
rect 407 1025 408 1029
rect 402 1024 408 1025
rect 658 1029 664 1030
rect 658 1025 659 1029
rect 663 1025 664 1029
rect 658 1024 664 1025
rect 270 1019 276 1020
rect 270 1015 271 1019
rect 275 1015 276 1019
rect 270 1014 276 1015
rect 354 1019 360 1020
rect 354 1015 355 1019
rect 359 1015 360 1019
rect 354 1014 360 1015
rect 356 980 358 1014
rect 354 979 360 980
rect 354 975 355 979
rect 359 975 360 979
rect 354 974 360 975
rect 362 979 368 980
rect 362 975 363 979
rect 367 975 368 979
rect 362 974 368 975
rect 111 950 115 951
rect 111 945 115 946
rect 147 950 151 951
rect 147 945 151 946
rect 235 950 239 951
rect 235 945 239 946
rect 112 885 114 945
rect 110 884 116 885
rect 236 884 238 945
rect 270 935 276 936
rect 270 931 271 935
rect 275 931 276 935
rect 270 930 276 931
rect 110 880 111 884
rect 115 880 116 884
rect 110 879 116 880
rect 234 883 240 884
rect 234 879 235 883
rect 239 879 240 883
rect 234 878 240 879
rect 262 868 268 869
rect 110 867 116 868
rect 110 863 111 867
rect 115 863 116 867
rect 262 864 263 868
rect 267 864 268 868
rect 262 863 268 864
rect 110 862 116 863
rect 112 823 114 862
rect 264 823 266 863
rect 111 822 115 823
rect 111 817 115 818
rect 175 822 179 823
rect 175 817 179 818
rect 263 822 267 823
rect 263 817 267 818
rect 112 794 114 817
rect 110 793 116 794
rect 176 793 178 817
rect 110 789 111 793
rect 115 789 116 793
rect 110 788 116 789
rect 174 792 180 793
rect 174 788 175 792
rect 179 788 180 792
rect 174 787 180 788
rect 146 777 152 778
rect 110 776 116 777
rect 110 772 111 776
rect 115 772 116 776
rect 146 773 147 777
rect 151 773 152 777
rect 146 772 152 773
rect 110 771 116 772
rect 112 711 114 771
rect 148 711 150 772
rect 272 768 274 930
rect 364 892 366 974
rect 404 951 406 1024
rect 660 951 662 1024
rect 756 980 758 1134
rect 836 1132 838 1193
rect 872 1184 874 1262
rect 940 1199 942 1272
rect 1036 1228 1038 1370
rect 1092 1368 1094 1429
rect 1404 1420 1406 1498
rect 1936 1435 1938 1507
rect 1976 1503 1978 1546
rect 2120 1503 2122 1547
rect 2188 1512 2190 1610
rect 2228 1568 2230 1629
rect 2234 1615 2240 1616
rect 2234 1611 2235 1615
rect 2239 1611 2240 1615
rect 2234 1610 2240 1611
rect 2236 1576 2238 1610
rect 2234 1575 2240 1576
rect 2234 1571 2235 1575
rect 2239 1571 2240 1575
rect 2234 1570 2240 1571
rect 2364 1568 2366 1629
rect 2370 1615 2376 1616
rect 2370 1611 2371 1615
rect 2375 1611 2376 1615
rect 2370 1610 2376 1611
rect 2372 1576 2374 1610
rect 2370 1575 2376 1576
rect 2370 1571 2371 1575
rect 2375 1571 2376 1575
rect 2370 1570 2376 1571
rect 2500 1568 2502 1629
rect 2506 1615 2512 1616
rect 2506 1611 2507 1615
rect 2511 1611 2512 1615
rect 2506 1610 2512 1611
rect 2508 1576 2510 1610
rect 2506 1575 2512 1576
rect 2506 1571 2507 1575
rect 2511 1571 2512 1575
rect 2506 1570 2512 1571
rect 2636 1568 2638 1629
rect 2642 1615 2648 1616
rect 2642 1611 2643 1615
rect 2647 1611 2648 1615
rect 2642 1610 2648 1611
rect 2644 1576 2646 1610
rect 2708 1584 2710 1654
rect 2780 1635 2782 1704
rect 2914 1699 2920 1700
rect 2914 1695 2915 1699
rect 2919 1695 2920 1699
rect 2914 1694 2920 1695
rect 2874 1691 2880 1692
rect 2874 1687 2875 1691
rect 2879 1687 2880 1691
rect 2874 1686 2880 1687
rect 2876 1660 2878 1686
rect 2874 1659 2880 1660
rect 2874 1655 2875 1659
rect 2879 1655 2880 1659
rect 2874 1654 2880 1655
rect 2771 1634 2775 1635
rect 2771 1629 2775 1630
rect 2779 1634 2783 1635
rect 2779 1629 2783 1630
rect 2907 1634 2911 1635
rect 2907 1629 2911 1630
rect 2706 1583 2712 1584
rect 2706 1579 2707 1583
rect 2711 1579 2712 1583
rect 2706 1578 2712 1579
rect 2642 1575 2648 1576
rect 2642 1571 2643 1575
rect 2647 1571 2648 1575
rect 2642 1570 2648 1571
rect 2772 1568 2774 1629
rect 2778 1615 2784 1616
rect 2778 1611 2779 1615
rect 2783 1611 2784 1615
rect 2778 1610 2784 1611
rect 2780 1576 2782 1610
rect 2778 1575 2784 1576
rect 2778 1571 2779 1575
rect 2783 1571 2784 1575
rect 2778 1570 2784 1571
rect 2908 1568 2910 1629
rect 2916 1620 2918 1694
rect 2948 1635 2950 1704
rect 3032 1660 3034 1810
rect 3108 1808 3110 1869
rect 3204 1860 3206 1938
rect 3236 1875 3238 1948
rect 3372 1875 3374 1948
rect 3468 1904 3470 2046
rect 3516 2044 3518 2105
rect 3652 2044 3654 2105
rect 3658 2091 3664 2092
rect 3658 2087 3659 2091
rect 3663 2087 3664 2091
rect 3658 2086 3664 2087
rect 3660 2052 3662 2086
rect 3748 2052 3750 2138
rect 3800 2111 3802 2187
rect 4514 2177 4520 2178
rect 3838 2176 3844 2177
rect 3838 2172 3839 2176
rect 3843 2172 3844 2176
rect 4514 2173 4515 2177
rect 4519 2173 4520 2177
rect 4514 2172 4520 2173
rect 4690 2177 4696 2178
rect 4690 2173 4691 2177
rect 4695 2173 4696 2177
rect 4690 2172 4696 2173
rect 4882 2177 4888 2178
rect 4882 2173 4883 2177
rect 4887 2173 4888 2177
rect 4882 2172 4888 2173
rect 3838 2171 3844 2172
rect 3840 2111 3842 2171
rect 4516 2111 4518 2172
rect 4642 2167 4648 2168
rect 4642 2163 4643 2167
rect 4647 2163 4648 2167
rect 4642 2162 4648 2163
rect 4670 2167 4676 2168
rect 4670 2163 4671 2167
rect 4675 2163 4676 2167
rect 4670 2162 4676 2163
rect 3799 2110 3803 2111
rect 3799 2105 3803 2106
rect 3839 2110 3843 2111
rect 3839 2105 3843 2106
rect 4515 2110 4519 2111
rect 4515 2105 4519 2106
rect 4635 2110 4639 2111
rect 4635 2105 4639 2106
rect 3766 2099 3772 2100
rect 3766 2095 3767 2099
rect 3771 2095 3772 2099
rect 3766 2094 3772 2095
rect 3658 2051 3664 2052
rect 3658 2047 3659 2051
rect 3663 2047 3664 2051
rect 3658 2046 3664 2047
rect 3746 2051 3752 2052
rect 3746 2047 3747 2051
rect 3751 2047 3752 2051
rect 3746 2046 3752 2047
rect 3514 2043 3520 2044
rect 3514 2039 3515 2043
rect 3519 2039 3520 2043
rect 3514 2038 3520 2039
rect 3650 2043 3656 2044
rect 3650 2039 3651 2043
rect 3655 2039 3656 2043
rect 3650 2038 3656 2039
rect 3542 2028 3548 2029
rect 3542 2024 3543 2028
rect 3547 2024 3548 2028
rect 3542 2023 3548 2024
rect 3678 2028 3684 2029
rect 3678 2024 3679 2028
rect 3683 2024 3684 2028
rect 3678 2023 3684 2024
rect 3544 1999 3546 2023
rect 3680 1999 3682 2023
rect 3535 1998 3539 1999
rect 3535 1993 3539 1994
rect 3543 1998 3547 1999
rect 3543 1993 3547 1994
rect 3671 1998 3675 1999
rect 3671 1993 3675 1994
rect 3679 1998 3683 1999
rect 3679 1993 3683 1994
rect 3536 1969 3538 1993
rect 3672 1969 3674 1993
rect 3534 1968 3540 1969
rect 3534 1964 3535 1968
rect 3539 1964 3540 1968
rect 3534 1963 3540 1964
rect 3670 1968 3676 1969
rect 3670 1964 3671 1968
rect 3675 1964 3676 1968
rect 3670 1963 3676 1964
rect 3506 1953 3512 1954
rect 3506 1949 3507 1953
rect 3511 1949 3512 1953
rect 3506 1948 3512 1949
rect 3642 1953 3648 1954
rect 3642 1949 3643 1953
rect 3647 1949 3648 1953
rect 3642 1948 3648 1949
rect 3466 1903 3472 1904
rect 3466 1899 3467 1903
rect 3471 1899 3472 1903
rect 3466 1898 3472 1899
rect 3508 1875 3510 1948
rect 3634 1943 3640 1944
rect 3634 1939 3635 1943
rect 3639 1939 3640 1943
rect 3634 1938 3640 1939
rect 3636 1904 3638 1938
rect 3602 1903 3608 1904
rect 3602 1899 3603 1903
rect 3607 1899 3608 1903
rect 3602 1898 3608 1899
rect 3634 1903 3640 1904
rect 3634 1899 3635 1903
rect 3639 1899 3640 1903
rect 3634 1898 3640 1899
rect 3235 1874 3239 1875
rect 3235 1869 3239 1870
rect 3299 1874 3303 1875
rect 3299 1869 3303 1870
rect 3371 1874 3375 1875
rect 3371 1869 3375 1870
rect 3483 1874 3487 1875
rect 3483 1869 3487 1870
rect 3507 1874 3511 1875
rect 3507 1869 3511 1870
rect 3202 1859 3208 1860
rect 3202 1855 3203 1859
rect 3207 1855 3208 1859
rect 3202 1854 3208 1855
rect 3300 1808 3302 1869
rect 3394 1855 3400 1856
rect 3394 1851 3395 1855
rect 3399 1851 3400 1855
rect 3394 1850 3400 1851
rect 3396 1824 3398 1850
rect 3394 1823 3400 1824
rect 3394 1819 3395 1823
rect 3399 1819 3400 1823
rect 3394 1818 3400 1819
rect 3484 1808 3486 1869
rect 3490 1855 3496 1856
rect 3490 1851 3491 1855
rect 3495 1851 3496 1855
rect 3490 1850 3496 1851
rect 3492 1816 3494 1850
rect 3604 1816 3606 1898
rect 3644 1875 3646 1948
rect 3768 1944 3770 2094
rect 3800 2045 3802 2105
rect 3840 2045 3842 2105
rect 3798 2044 3804 2045
rect 3798 2040 3799 2044
rect 3803 2040 3804 2044
rect 3798 2039 3804 2040
rect 3838 2044 3844 2045
rect 4636 2044 4638 2105
rect 4644 2096 4646 2162
rect 4672 2128 4674 2162
rect 4670 2127 4676 2128
rect 4670 2123 4671 2127
rect 4675 2123 4676 2127
rect 4670 2122 4676 2123
rect 4692 2111 4694 2172
rect 4884 2111 4886 2172
rect 4904 2128 4906 2282
rect 4964 2280 4966 2341
rect 5100 2288 5102 2370
rect 5372 2347 5374 2420
rect 5434 2415 5440 2416
rect 5434 2411 5435 2415
rect 5439 2411 5440 2415
rect 5434 2410 5440 2411
rect 5147 2346 5151 2347
rect 5147 2341 5151 2342
rect 5339 2346 5343 2347
rect 5339 2341 5343 2342
rect 5371 2346 5375 2347
rect 5371 2341 5375 2342
rect 5098 2287 5104 2288
rect 5098 2283 5099 2287
rect 5103 2283 5104 2287
rect 5098 2282 5104 2283
rect 5148 2280 5150 2341
rect 5326 2331 5332 2332
rect 5326 2327 5327 2331
rect 5331 2327 5332 2331
rect 5326 2326 5332 2327
rect 4962 2279 4968 2280
rect 4962 2275 4963 2279
rect 4967 2275 4968 2279
rect 4962 2274 4968 2275
rect 5146 2279 5152 2280
rect 5146 2275 5147 2279
rect 5151 2275 5152 2279
rect 5146 2274 5152 2275
rect 4990 2264 4996 2265
rect 4990 2260 4991 2264
rect 4995 2260 4996 2264
rect 4990 2259 4996 2260
rect 5174 2264 5180 2265
rect 5174 2260 5175 2264
rect 5179 2260 5180 2264
rect 5174 2259 5180 2260
rect 4992 2223 4994 2259
rect 5176 2223 5178 2259
rect 4911 2222 4915 2223
rect 4911 2217 4915 2218
rect 4991 2222 4995 2223
rect 4991 2217 4995 2218
rect 5119 2222 5123 2223
rect 5119 2217 5123 2218
rect 5175 2222 5179 2223
rect 5175 2217 5179 2218
rect 4912 2193 4914 2217
rect 5120 2193 5122 2217
rect 4910 2192 4916 2193
rect 4910 2188 4911 2192
rect 4915 2188 4916 2192
rect 4910 2187 4916 2188
rect 5118 2192 5124 2193
rect 5118 2188 5119 2192
rect 5123 2188 5124 2192
rect 5118 2187 5124 2188
rect 5090 2177 5096 2178
rect 5090 2173 5091 2177
rect 5095 2173 5096 2177
rect 5090 2172 5096 2173
rect 5306 2177 5312 2178
rect 5306 2173 5307 2177
rect 5311 2173 5312 2177
rect 5306 2172 5312 2173
rect 4902 2127 4908 2128
rect 4902 2123 4903 2127
rect 4907 2123 4908 2127
rect 4902 2122 4908 2123
rect 5092 2111 5094 2172
rect 5278 2167 5284 2168
rect 5278 2163 5279 2167
rect 5283 2163 5284 2167
rect 5278 2162 5284 2163
rect 5280 2128 5282 2162
rect 5166 2127 5172 2128
rect 5166 2123 5167 2127
rect 5171 2123 5172 2127
rect 5166 2122 5172 2123
rect 5278 2127 5284 2128
rect 5278 2123 5279 2127
rect 5283 2123 5284 2127
rect 5278 2122 5284 2123
rect 4691 2110 4695 2111
rect 4691 2105 4695 2106
rect 4771 2110 4775 2111
rect 4771 2105 4775 2106
rect 4883 2110 4887 2111
rect 4883 2105 4887 2106
rect 4907 2110 4911 2111
rect 4907 2105 4911 2106
rect 5043 2110 5047 2111
rect 5043 2105 5047 2106
rect 5091 2110 5095 2111
rect 5091 2105 5095 2106
rect 4642 2095 4648 2096
rect 4642 2091 4643 2095
rect 4647 2091 4648 2095
rect 4642 2090 4648 2091
rect 4772 2044 4774 2105
rect 4778 2091 4784 2092
rect 4778 2087 4779 2091
rect 4783 2087 4784 2091
rect 4778 2086 4784 2087
rect 4780 2052 4782 2086
rect 4778 2051 4784 2052
rect 4778 2047 4779 2051
rect 4783 2047 4784 2051
rect 4778 2046 4784 2047
rect 4908 2044 4910 2105
rect 4914 2091 4920 2092
rect 4914 2087 4915 2091
rect 4919 2087 4920 2091
rect 4914 2086 4920 2087
rect 4916 2052 4918 2086
rect 4914 2051 4920 2052
rect 4914 2047 4915 2051
rect 4919 2047 4920 2051
rect 4914 2046 4920 2047
rect 5044 2044 5046 2105
rect 5050 2091 5056 2092
rect 5050 2087 5051 2091
rect 5055 2087 5056 2091
rect 5050 2086 5056 2087
rect 5052 2052 5054 2086
rect 5168 2052 5170 2122
rect 5308 2111 5310 2172
rect 5328 2168 5330 2326
rect 5340 2280 5342 2341
rect 5436 2332 5438 2410
rect 5448 2376 5450 2522
rect 5664 2521 5666 2581
rect 5662 2520 5668 2521
rect 5662 2516 5663 2520
rect 5667 2516 5668 2520
rect 5662 2515 5668 2516
rect 5662 2503 5668 2504
rect 5662 2499 5663 2503
rect 5667 2499 5668 2503
rect 5662 2498 5668 2499
rect 5664 2471 5666 2498
rect 5663 2470 5667 2471
rect 5663 2465 5667 2466
rect 5664 2442 5666 2465
rect 5662 2441 5668 2442
rect 5662 2437 5663 2441
rect 5667 2437 5668 2441
rect 5662 2436 5668 2437
rect 5662 2424 5668 2425
rect 5662 2420 5663 2424
rect 5667 2420 5668 2424
rect 5662 2419 5668 2420
rect 5446 2375 5452 2376
rect 5446 2371 5447 2375
rect 5451 2371 5452 2375
rect 5446 2370 5452 2371
rect 5664 2347 5666 2419
rect 5515 2346 5519 2347
rect 5515 2341 5519 2342
rect 5663 2346 5667 2347
rect 5663 2341 5667 2342
rect 5434 2331 5440 2332
rect 5434 2327 5435 2331
rect 5439 2327 5440 2331
rect 5434 2326 5440 2327
rect 5516 2280 5518 2341
rect 5522 2327 5528 2328
rect 5522 2323 5523 2327
rect 5527 2323 5528 2327
rect 5522 2322 5528 2323
rect 5524 2288 5526 2322
rect 5522 2287 5528 2288
rect 5522 2283 5523 2287
rect 5527 2283 5528 2287
rect 5522 2282 5528 2283
rect 5610 2287 5616 2288
rect 5610 2283 5611 2287
rect 5615 2283 5616 2287
rect 5610 2282 5616 2283
rect 5338 2279 5344 2280
rect 5338 2275 5339 2279
rect 5343 2275 5344 2279
rect 5338 2274 5344 2275
rect 5514 2279 5520 2280
rect 5514 2275 5515 2279
rect 5519 2275 5520 2279
rect 5514 2274 5520 2275
rect 5366 2264 5372 2265
rect 5366 2260 5367 2264
rect 5371 2260 5372 2264
rect 5366 2259 5372 2260
rect 5542 2264 5548 2265
rect 5542 2260 5543 2264
rect 5547 2260 5548 2264
rect 5542 2259 5548 2260
rect 5368 2223 5370 2259
rect 5544 2223 5546 2259
rect 5335 2222 5339 2223
rect 5335 2217 5339 2218
rect 5367 2222 5371 2223
rect 5367 2217 5371 2218
rect 5543 2222 5547 2223
rect 5543 2217 5547 2218
rect 5336 2193 5338 2217
rect 5544 2193 5546 2217
rect 5334 2192 5340 2193
rect 5334 2188 5335 2192
rect 5339 2188 5340 2192
rect 5334 2187 5340 2188
rect 5542 2192 5548 2193
rect 5542 2188 5543 2192
rect 5547 2188 5548 2192
rect 5542 2187 5548 2188
rect 5514 2177 5520 2178
rect 5514 2173 5515 2177
rect 5519 2173 5520 2177
rect 5514 2172 5520 2173
rect 5326 2167 5332 2168
rect 5326 2163 5327 2167
rect 5331 2163 5332 2167
rect 5326 2162 5332 2163
rect 5516 2111 5518 2172
rect 5612 2128 5614 2282
rect 5664 2281 5666 2341
rect 5662 2280 5668 2281
rect 5662 2276 5663 2280
rect 5667 2276 5668 2280
rect 5662 2275 5668 2276
rect 5662 2263 5668 2264
rect 5662 2259 5663 2263
rect 5667 2259 5668 2263
rect 5662 2258 5668 2259
rect 5664 2223 5666 2258
rect 5663 2222 5667 2223
rect 5663 2217 5667 2218
rect 5664 2194 5666 2217
rect 5662 2193 5668 2194
rect 5662 2189 5663 2193
rect 5667 2189 5668 2193
rect 5662 2188 5668 2189
rect 5662 2176 5668 2177
rect 5662 2172 5663 2176
rect 5667 2172 5668 2176
rect 5662 2171 5668 2172
rect 5638 2167 5644 2168
rect 5638 2163 5639 2167
rect 5643 2163 5644 2167
rect 5638 2162 5644 2163
rect 5610 2127 5616 2128
rect 5610 2123 5611 2127
rect 5615 2123 5616 2127
rect 5610 2122 5616 2123
rect 5179 2110 5183 2111
rect 5179 2105 5183 2106
rect 5307 2110 5311 2111
rect 5307 2105 5311 2106
rect 5515 2110 5519 2111
rect 5515 2105 5519 2106
rect 5050 2051 5056 2052
rect 5050 2047 5051 2051
rect 5055 2047 5056 2051
rect 5050 2046 5056 2047
rect 5166 2051 5172 2052
rect 5166 2047 5167 2051
rect 5171 2047 5172 2051
rect 5166 2046 5172 2047
rect 5180 2044 5182 2105
rect 5366 2095 5372 2096
rect 5366 2091 5367 2095
rect 5371 2091 5372 2095
rect 5366 2090 5372 2091
rect 5218 2051 5224 2052
rect 5218 2047 5219 2051
rect 5223 2047 5224 2051
rect 5218 2046 5224 2047
rect 3838 2040 3839 2044
rect 3843 2040 3844 2044
rect 3838 2039 3844 2040
rect 4634 2043 4640 2044
rect 4634 2039 4635 2043
rect 4639 2039 4640 2043
rect 4634 2038 4640 2039
rect 4770 2043 4776 2044
rect 4770 2039 4771 2043
rect 4775 2039 4776 2043
rect 4770 2038 4776 2039
rect 4906 2043 4912 2044
rect 4906 2039 4907 2043
rect 4911 2039 4912 2043
rect 4906 2038 4912 2039
rect 5042 2043 5048 2044
rect 5042 2039 5043 2043
rect 5047 2039 5048 2043
rect 5042 2038 5048 2039
rect 5178 2043 5184 2044
rect 5178 2039 5179 2043
rect 5183 2039 5184 2043
rect 5178 2038 5184 2039
rect 4662 2028 4668 2029
rect 3798 2027 3804 2028
rect 3798 2023 3799 2027
rect 3803 2023 3804 2027
rect 3798 2022 3804 2023
rect 3838 2027 3844 2028
rect 3838 2023 3839 2027
rect 3843 2023 3844 2027
rect 4662 2024 4663 2028
rect 4667 2024 4668 2028
rect 4662 2023 4668 2024
rect 4798 2028 4804 2029
rect 4798 2024 4799 2028
rect 4803 2024 4804 2028
rect 4798 2023 4804 2024
rect 4934 2028 4940 2029
rect 4934 2024 4935 2028
rect 4939 2024 4940 2028
rect 4934 2023 4940 2024
rect 5070 2028 5076 2029
rect 5070 2024 5071 2028
rect 5075 2024 5076 2028
rect 5070 2023 5076 2024
rect 5206 2028 5212 2029
rect 5206 2024 5207 2028
rect 5211 2024 5212 2028
rect 5206 2023 5212 2024
rect 3838 2022 3844 2023
rect 3800 1999 3802 2022
rect 3840 1999 3842 2022
rect 4664 1999 4666 2023
rect 4800 1999 4802 2023
rect 4936 1999 4938 2023
rect 5072 1999 5074 2023
rect 5208 1999 5210 2023
rect 3799 1998 3803 1999
rect 3799 1993 3803 1994
rect 3839 1998 3843 1999
rect 3839 1993 3843 1994
rect 4663 1998 4667 1999
rect 4663 1993 4667 1994
rect 4799 1998 4803 1999
rect 4799 1993 4803 1994
rect 4863 1998 4867 1999
rect 4863 1993 4867 1994
rect 4935 1998 4939 1999
rect 4935 1993 4939 1994
rect 4999 1998 5003 1999
rect 4999 1993 5003 1994
rect 5071 1998 5075 1999
rect 5071 1993 5075 1994
rect 5135 1998 5139 1999
rect 5135 1993 5139 1994
rect 5207 1998 5211 1999
rect 5207 1993 5211 1994
rect 3800 1970 3802 1993
rect 3840 1970 3842 1993
rect 3798 1969 3804 1970
rect 3798 1965 3799 1969
rect 3803 1965 3804 1969
rect 3798 1964 3804 1965
rect 3838 1969 3844 1970
rect 4864 1969 4866 1993
rect 5000 1969 5002 1993
rect 5136 1969 5138 1993
rect 3838 1965 3839 1969
rect 3843 1965 3844 1969
rect 3838 1964 3844 1965
rect 4862 1968 4868 1969
rect 4862 1964 4863 1968
rect 4867 1964 4868 1968
rect 4862 1963 4868 1964
rect 4998 1968 5004 1969
rect 4998 1964 4999 1968
rect 5003 1964 5004 1968
rect 4998 1963 5004 1964
rect 5134 1968 5140 1969
rect 5134 1964 5135 1968
rect 5139 1964 5140 1968
rect 5134 1963 5140 1964
rect 4834 1953 4840 1954
rect 3798 1952 3804 1953
rect 3798 1948 3799 1952
rect 3803 1948 3804 1952
rect 3798 1947 3804 1948
rect 3838 1952 3844 1953
rect 3838 1948 3839 1952
rect 3843 1948 3844 1952
rect 4834 1949 4835 1953
rect 4839 1949 4840 1953
rect 4834 1948 4840 1949
rect 4970 1953 4976 1954
rect 4970 1949 4971 1953
rect 4975 1949 4976 1953
rect 4970 1948 4976 1949
rect 5106 1953 5112 1954
rect 5106 1949 5107 1953
rect 5111 1949 5112 1953
rect 5106 1948 5112 1949
rect 3838 1947 3844 1948
rect 3766 1943 3772 1944
rect 3766 1939 3767 1943
rect 3771 1939 3772 1943
rect 3766 1938 3772 1939
rect 3800 1875 3802 1947
rect 3840 1875 3842 1947
rect 4770 1943 4776 1944
rect 4770 1939 4771 1943
rect 4775 1939 4776 1943
rect 4770 1938 4776 1939
rect 3643 1874 3647 1875
rect 3643 1869 3647 1870
rect 3651 1874 3655 1875
rect 3651 1869 3655 1870
rect 3799 1874 3803 1875
rect 3799 1869 3803 1870
rect 3839 1874 3843 1875
rect 3839 1869 3843 1870
rect 4675 1874 4679 1875
rect 4675 1869 4679 1870
rect 3490 1815 3496 1816
rect 3490 1811 3491 1815
rect 3495 1811 3496 1815
rect 3490 1810 3496 1811
rect 3602 1815 3608 1816
rect 3602 1811 3603 1815
rect 3607 1811 3608 1815
rect 3602 1810 3608 1811
rect 3652 1808 3654 1869
rect 3800 1809 3802 1869
rect 3840 1809 3842 1869
rect 3982 1859 3988 1860
rect 3982 1855 3983 1859
rect 3987 1855 3988 1859
rect 3982 1854 3988 1855
rect 3798 1808 3804 1809
rect 3106 1807 3112 1808
rect 3106 1803 3107 1807
rect 3111 1803 3112 1807
rect 3106 1802 3112 1803
rect 3298 1807 3304 1808
rect 3298 1803 3299 1807
rect 3303 1803 3304 1807
rect 3298 1802 3304 1803
rect 3482 1807 3488 1808
rect 3482 1803 3483 1807
rect 3487 1803 3488 1807
rect 3482 1802 3488 1803
rect 3650 1807 3656 1808
rect 3650 1803 3651 1807
rect 3655 1803 3656 1807
rect 3798 1804 3799 1808
rect 3803 1804 3804 1808
rect 3798 1803 3804 1804
rect 3838 1808 3844 1809
rect 3838 1804 3839 1808
rect 3843 1804 3844 1808
rect 3838 1803 3844 1804
rect 3650 1802 3656 1803
rect 3134 1792 3140 1793
rect 3134 1788 3135 1792
rect 3139 1788 3140 1792
rect 3134 1787 3140 1788
rect 3326 1792 3332 1793
rect 3326 1788 3327 1792
rect 3331 1788 3332 1792
rect 3326 1787 3332 1788
rect 3510 1792 3516 1793
rect 3510 1788 3511 1792
rect 3515 1788 3516 1792
rect 3510 1787 3516 1788
rect 3678 1792 3684 1793
rect 3678 1788 3679 1792
rect 3683 1788 3684 1792
rect 3678 1787 3684 1788
rect 3798 1791 3804 1792
rect 3798 1787 3799 1791
rect 3803 1787 3804 1791
rect 3136 1755 3138 1787
rect 3328 1755 3330 1787
rect 3512 1755 3514 1787
rect 3680 1755 3682 1787
rect 3798 1786 3804 1787
rect 3838 1791 3844 1792
rect 3838 1787 3839 1791
rect 3843 1787 3844 1791
rect 3838 1786 3844 1787
rect 3800 1755 3802 1786
rect 3135 1754 3139 1755
rect 3135 1749 3139 1750
rect 3151 1754 3155 1755
rect 3151 1749 3155 1750
rect 3327 1754 3331 1755
rect 3327 1749 3331 1750
rect 3511 1754 3515 1755
rect 3511 1749 3515 1750
rect 3679 1754 3683 1755
rect 3679 1749 3683 1750
rect 3799 1754 3803 1755
rect 3799 1749 3803 1750
rect 3152 1725 3154 1749
rect 3800 1726 3802 1749
rect 3840 1747 3842 1786
rect 3839 1746 3843 1747
rect 3839 1741 3843 1742
rect 3887 1746 3891 1747
rect 3887 1741 3891 1742
rect 3798 1725 3804 1726
rect 3150 1724 3156 1725
rect 3150 1720 3151 1724
rect 3155 1720 3156 1724
rect 3798 1721 3799 1725
rect 3803 1721 3804 1725
rect 3798 1720 3804 1721
rect 3150 1719 3156 1720
rect 3840 1718 3842 1741
rect 3838 1717 3844 1718
rect 3888 1717 3890 1741
rect 3838 1713 3839 1717
rect 3843 1713 3844 1717
rect 3838 1712 3844 1713
rect 3886 1716 3892 1717
rect 3886 1712 3887 1716
rect 3891 1712 3892 1716
rect 3886 1711 3892 1712
rect 3122 1709 3128 1710
rect 3122 1705 3123 1709
rect 3127 1705 3128 1709
rect 3122 1704 3128 1705
rect 3798 1708 3804 1709
rect 3798 1704 3799 1708
rect 3803 1704 3804 1708
rect 3074 1699 3080 1700
rect 3074 1695 3075 1699
rect 3079 1695 3080 1699
rect 3074 1694 3080 1695
rect 3076 1660 3078 1694
rect 3030 1659 3036 1660
rect 3030 1655 3031 1659
rect 3035 1655 3036 1659
rect 3030 1654 3036 1655
rect 3074 1659 3080 1660
rect 3074 1655 3075 1659
rect 3079 1655 3080 1659
rect 3074 1654 3080 1655
rect 3124 1635 3126 1704
rect 3798 1703 3804 1704
rect 3800 1635 3802 1703
rect 3858 1701 3864 1702
rect 3838 1700 3844 1701
rect 3838 1696 3839 1700
rect 3843 1696 3844 1700
rect 3858 1697 3859 1701
rect 3863 1697 3864 1701
rect 3858 1696 3864 1697
rect 3838 1695 3844 1696
rect 3840 1635 3842 1695
rect 3860 1635 3862 1696
rect 3984 1692 3986 1854
rect 4676 1808 4678 1869
rect 4772 1860 4774 1938
rect 4836 1875 4838 1948
rect 4972 1875 4974 1948
rect 5108 1875 5110 1948
rect 5220 1904 5222 2046
rect 5271 1998 5275 1999
rect 5271 1993 5275 1994
rect 5272 1969 5274 1993
rect 5270 1968 5276 1969
rect 5270 1964 5271 1968
rect 5275 1964 5276 1968
rect 5270 1963 5276 1964
rect 5242 1953 5248 1954
rect 5242 1949 5243 1953
rect 5247 1949 5248 1953
rect 5242 1948 5248 1949
rect 5218 1903 5224 1904
rect 5218 1899 5219 1903
rect 5223 1899 5224 1903
rect 5218 1898 5224 1899
rect 5244 1875 5246 1948
rect 5368 1944 5370 2090
rect 5407 1998 5411 1999
rect 5407 1993 5411 1994
rect 5543 1998 5547 1999
rect 5543 1993 5547 1994
rect 5408 1969 5410 1993
rect 5544 1969 5546 1993
rect 5406 1968 5412 1969
rect 5406 1964 5407 1968
rect 5411 1964 5412 1968
rect 5406 1963 5412 1964
rect 5542 1968 5548 1969
rect 5542 1964 5543 1968
rect 5547 1964 5548 1968
rect 5542 1963 5548 1964
rect 5378 1953 5384 1954
rect 5378 1949 5379 1953
rect 5383 1949 5384 1953
rect 5378 1948 5384 1949
rect 5514 1953 5520 1954
rect 5514 1949 5515 1953
rect 5519 1949 5520 1953
rect 5514 1948 5520 1949
rect 5366 1943 5372 1944
rect 5366 1939 5367 1943
rect 5371 1939 5372 1943
rect 5366 1938 5372 1939
rect 5380 1875 5382 1948
rect 5386 1943 5392 1944
rect 5386 1939 5387 1943
rect 5391 1939 5392 1943
rect 5386 1938 5392 1939
rect 5388 1912 5390 1938
rect 5386 1911 5392 1912
rect 5386 1907 5387 1911
rect 5391 1907 5392 1911
rect 5386 1906 5392 1907
rect 5516 1875 5518 1948
rect 5610 1943 5616 1944
rect 5610 1939 5611 1943
rect 5615 1939 5616 1943
rect 5610 1938 5616 1939
rect 4819 1874 4823 1875
rect 4819 1869 4823 1870
rect 4835 1874 4839 1875
rect 4835 1869 4839 1870
rect 4963 1874 4967 1875
rect 4963 1869 4967 1870
rect 4971 1874 4975 1875
rect 4971 1869 4975 1870
rect 5107 1874 5111 1875
rect 5107 1869 5111 1870
rect 5243 1874 5247 1875
rect 5243 1869 5247 1870
rect 5379 1874 5383 1875
rect 5379 1869 5383 1870
rect 5515 1874 5519 1875
rect 5515 1869 5519 1870
rect 4770 1859 4776 1860
rect 4770 1855 4771 1859
rect 4775 1855 4776 1859
rect 4770 1854 4776 1855
rect 4820 1808 4822 1869
rect 4826 1855 4832 1856
rect 4826 1851 4827 1855
rect 4831 1851 4832 1855
rect 4826 1850 4832 1851
rect 4828 1816 4830 1850
rect 4826 1815 4832 1816
rect 4826 1811 4827 1815
rect 4831 1811 4832 1815
rect 4826 1810 4832 1811
rect 4964 1808 4966 1869
rect 4970 1855 4976 1856
rect 4970 1851 4971 1855
rect 4975 1851 4976 1855
rect 4970 1850 4976 1851
rect 4972 1816 4974 1850
rect 4970 1815 4976 1816
rect 4970 1811 4971 1815
rect 4975 1811 4976 1815
rect 4970 1810 4976 1811
rect 5086 1815 5092 1816
rect 5086 1811 5087 1815
rect 5091 1811 5092 1815
rect 5086 1810 5092 1811
rect 4674 1807 4680 1808
rect 4674 1803 4675 1807
rect 4679 1803 4680 1807
rect 4674 1802 4680 1803
rect 4818 1807 4824 1808
rect 4818 1803 4819 1807
rect 4823 1803 4824 1807
rect 4818 1802 4824 1803
rect 4962 1807 4968 1808
rect 4962 1803 4963 1807
rect 4967 1803 4968 1807
rect 4962 1802 4968 1803
rect 4702 1792 4708 1793
rect 4702 1788 4703 1792
rect 4707 1788 4708 1792
rect 4702 1787 4708 1788
rect 4846 1792 4852 1793
rect 4846 1788 4847 1792
rect 4851 1788 4852 1792
rect 4846 1787 4852 1788
rect 4990 1792 4996 1793
rect 4990 1788 4991 1792
rect 4995 1788 4996 1792
rect 4990 1787 4996 1788
rect 4704 1747 4706 1787
rect 4848 1747 4850 1787
rect 4992 1747 4994 1787
rect 4079 1746 4083 1747
rect 4079 1741 4083 1742
rect 4303 1746 4307 1747
rect 4303 1741 4307 1742
rect 4535 1746 4539 1747
rect 4535 1741 4539 1742
rect 4703 1746 4707 1747
rect 4703 1741 4707 1742
rect 4775 1746 4779 1747
rect 4775 1741 4779 1742
rect 4847 1746 4851 1747
rect 4847 1741 4851 1742
rect 4991 1746 4995 1747
rect 4991 1741 4995 1742
rect 5023 1746 5027 1747
rect 5023 1741 5027 1742
rect 4080 1717 4082 1741
rect 4304 1717 4306 1741
rect 4536 1717 4538 1741
rect 4776 1717 4778 1741
rect 5024 1717 5026 1741
rect 4078 1716 4084 1717
rect 4078 1712 4079 1716
rect 4083 1712 4084 1716
rect 4078 1711 4084 1712
rect 4302 1716 4308 1717
rect 4302 1712 4303 1716
rect 4307 1712 4308 1716
rect 4302 1711 4308 1712
rect 4534 1716 4540 1717
rect 4534 1712 4535 1716
rect 4539 1712 4540 1716
rect 4534 1711 4540 1712
rect 4774 1716 4780 1717
rect 4774 1712 4775 1716
rect 4779 1712 4780 1716
rect 4774 1711 4780 1712
rect 5022 1716 5028 1717
rect 5022 1712 5023 1716
rect 5027 1712 5028 1716
rect 5022 1711 5028 1712
rect 4050 1701 4056 1702
rect 4050 1697 4051 1701
rect 4055 1697 4056 1701
rect 4050 1696 4056 1697
rect 4274 1701 4280 1702
rect 4274 1697 4275 1701
rect 4279 1697 4280 1701
rect 4274 1696 4280 1697
rect 4506 1701 4512 1702
rect 4506 1697 4507 1701
rect 4511 1697 4512 1701
rect 4506 1696 4512 1697
rect 4746 1701 4752 1702
rect 4746 1697 4747 1701
rect 4751 1697 4752 1701
rect 4746 1696 4752 1697
rect 4994 1701 5000 1702
rect 4994 1697 4995 1701
rect 4999 1697 5000 1701
rect 4994 1696 5000 1697
rect 3982 1691 3988 1692
rect 3982 1687 3983 1691
rect 3987 1687 3988 1691
rect 3982 1686 3988 1687
rect 4052 1635 4054 1696
rect 4146 1651 4152 1652
rect 4146 1647 4147 1651
rect 4151 1647 4152 1651
rect 4146 1646 4152 1647
rect 2947 1634 2951 1635
rect 2947 1629 2951 1630
rect 3043 1634 3047 1635
rect 3043 1629 3047 1630
rect 3123 1634 3127 1635
rect 3123 1629 3127 1630
rect 3179 1634 3183 1635
rect 3179 1629 3183 1630
rect 3799 1634 3803 1635
rect 3799 1629 3803 1630
rect 3839 1634 3843 1635
rect 3839 1629 3843 1630
rect 3859 1634 3863 1635
rect 3859 1629 3863 1630
rect 3995 1634 3999 1635
rect 3995 1629 3999 1630
rect 4051 1634 4055 1635
rect 4051 1629 4055 1630
rect 2914 1619 2920 1620
rect 2914 1615 2915 1619
rect 2919 1615 2920 1619
rect 2914 1614 2920 1615
rect 3044 1568 3046 1629
rect 3050 1615 3056 1616
rect 3050 1611 3051 1615
rect 3055 1611 3056 1615
rect 3050 1610 3056 1611
rect 3052 1576 3054 1610
rect 3050 1575 3056 1576
rect 3050 1571 3051 1575
rect 3055 1571 3056 1575
rect 3050 1570 3056 1571
rect 3180 1568 3182 1629
rect 3186 1615 3192 1616
rect 3186 1611 3187 1615
rect 3191 1611 3192 1615
rect 3186 1610 3192 1611
rect 3188 1576 3190 1610
rect 3186 1575 3192 1576
rect 3186 1571 3187 1575
rect 3191 1571 3192 1575
rect 3186 1570 3192 1571
rect 3298 1575 3304 1576
rect 3298 1571 3299 1575
rect 3303 1571 3304 1575
rect 3298 1570 3304 1571
rect 2226 1567 2232 1568
rect 2226 1563 2227 1567
rect 2231 1563 2232 1567
rect 2226 1562 2232 1563
rect 2362 1567 2368 1568
rect 2362 1563 2363 1567
rect 2367 1563 2368 1567
rect 2362 1562 2368 1563
rect 2498 1567 2504 1568
rect 2498 1563 2499 1567
rect 2503 1563 2504 1567
rect 2498 1562 2504 1563
rect 2634 1567 2640 1568
rect 2634 1563 2635 1567
rect 2639 1563 2640 1567
rect 2634 1562 2640 1563
rect 2770 1567 2776 1568
rect 2770 1563 2771 1567
rect 2775 1563 2776 1567
rect 2770 1562 2776 1563
rect 2906 1567 2912 1568
rect 2906 1563 2907 1567
rect 2911 1563 2912 1567
rect 2906 1562 2912 1563
rect 3042 1567 3048 1568
rect 3042 1563 3043 1567
rect 3047 1563 3048 1567
rect 3042 1562 3048 1563
rect 3178 1567 3184 1568
rect 3178 1563 3179 1567
rect 3183 1563 3184 1567
rect 3178 1562 3184 1563
rect 2254 1552 2260 1553
rect 2254 1548 2255 1552
rect 2259 1548 2260 1552
rect 2254 1547 2260 1548
rect 2390 1552 2396 1553
rect 2390 1548 2391 1552
rect 2395 1548 2396 1552
rect 2390 1547 2396 1548
rect 2526 1552 2532 1553
rect 2526 1548 2527 1552
rect 2531 1548 2532 1552
rect 2526 1547 2532 1548
rect 2662 1552 2668 1553
rect 2662 1548 2663 1552
rect 2667 1548 2668 1552
rect 2662 1547 2668 1548
rect 2798 1552 2804 1553
rect 2798 1548 2799 1552
rect 2803 1548 2804 1552
rect 2798 1547 2804 1548
rect 2934 1552 2940 1553
rect 2934 1548 2935 1552
rect 2939 1548 2940 1552
rect 2934 1547 2940 1548
rect 3070 1552 3076 1553
rect 3070 1548 3071 1552
rect 3075 1548 3076 1552
rect 3070 1547 3076 1548
rect 3206 1552 3212 1553
rect 3206 1548 3207 1552
rect 3211 1548 3212 1552
rect 3206 1547 3212 1548
rect 2186 1511 2192 1512
rect 2186 1507 2187 1511
rect 2191 1507 2192 1511
rect 2186 1506 2192 1507
rect 2256 1503 2258 1547
rect 2392 1503 2394 1547
rect 2528 1503 2530 1547
rect 2654 1511 2660 1512
rect 2654 1507 2655 1511
rect 2659 1507 2660 1511
rect 2654 1506 2660 1507
rect 1975 1502 1979 1503
rect 1975 1497 1979 1498
rect 2023 1502 2027 1503
rect 2023 1497 2027 1498
rect 2119 1502 2123 1503
rect 2119 1497 2123 1498
rect 2159 1502 2163 1503
rect 2159 1497 2163 1498
rect 2255 1502 2259 1503
rect 2255 1497 2259 1498
rect 2295 1502 2299 1503
rect 2295 1497 2299 1498
rect 2391 1502 2395 1503
rect 2391 1497 2395 1498
rect 2431 1502 2435 1503
rect 2431 1497 2435 1498
rect 2527 1502 2531 1503
rect 2527 1497 2531 1498
rect 2567 1502 2571 1503
rect 2567 1497 2571 1498
rect 1976 1474 1978 1497
rect 1974 1473 1980 1474
rect 2024 1473 2026 1497
rect 2160 1473 2162 1497
rect 2296 1473 2298 1497
rect 2432 1473 2434 1497
rect 2568 1473 2570 1497
rect 1974 1469 1975 1473
rect 1979 1469 1980 1473
rect 1974 1468 1980 1469
rect 2022 1472 2028 1473
rect 2022 1468 2023 1472
rect 2027 1468 2028 1472
rect 2022 1467 2028 1468
rect 2158 1472 2164 1473
rect 2158 1468 2159 1472
rect 2163 1468 2164 1472
rect 2158 1467 2164 1468
rect 2294 1472 2300 1473
rect 2294 1468 2295 1472
rect 2299 1468 2300 1472
rect 2294 1467 2300 1468
rect 2430 1472 2436 1473
rect 2430 1468 2431 1472
rect 2435 1468 2436 1472
rect 2430 1467 2436 1468
rect 2566 1472 2572 1473
rect 2566 1468 2567 1472
rect 2571 1468 2572 1472
rect 2566 1467 2572 1468
rect 1994 1457 2000 1458
rect 1974 1456 1980 1457
rect 1974 1452 1975 1456
rect 1979 1452 1980 1456
rect 1994 1453 1995 1457
rect 1999 1453 2000 1457
rect 1994 1452 2000 1453
rect 2130 1457 2136 1458
rect 2130 1453 2131 1457
rect 2135 1453 2136 1457
rect 2130 1452 2136 1453
rect 2266 1457 2272 1458
rect 2266 1453 2267 1457
rect 2271 1453 2272 1457
rect 2266 1452 2272 1453
rect 2402 1457 2408 1458
rect 2402 1453 2403 1457
rect 2407 1453 2408 1457
rect 2402 1452 2408 1453
rect 2538 1457 2544 1458
rect 2538 1453 2539 1457
rect 2543 1453 2544 1457
rect 2538 1452 2544 1453
rect 1974 1451 1980 1452
rect 1451 1434 1455 1435
rect 1451 1429 1455 1430
rect 1787 1434 1791 1435
rect 1787 1429 1791 1430
rect 1935 1434 1939 1435
rect 1935 1429 1939 1430
rect 1402 1419 1408 1420
rect 1186 1415 1192 1416
rect 1186 1411 1187 1415
rect 1191 1411 1192 1415
rect 1402 1415 1403 1419
rect 1407 1415 1408 1419
rect 1402 1414 1408 1415
rect 1186 1410 1192 1411
rect 1188 1396 1190 1410
rect 1186 1395 1192 1396
rect 1186 1391 1187 1395
rect 1191 1391 1192 1395
rect 1186 1390 1192 1391
rect 1452 1368 1454 1429
rect 1574 1395 1580 1396
rect 1574 1391 1575 1395
rect 1579 1391 1580 1395
rect 1574 1390 1580 1391
rect 1576 1376 1578 1390
rect 1574 1375 1580 1376
rect 1574 1371 1575 1375
rect 1579 1371 1580 1375
rect 1574 1370 1580 1371
rect 1788 1368 1790 1429
rect 1882 1415 1888 1416
rect 1882 1411 1883 1415
rect 1887 1411 1888 1415
rect 1882 1410 1888 1411
rect 1090 1367 1096 1368
rect 1090 1363 1091 1367
rect 1095 1363 1096 1367
rect 1090 1362 1096 1363
rect 1450 1367 1456 1368
rect 1450 1363 1451 1367
rect 1455 1363 1456 1367
rect 1450 1362 1456 1363
rect 1786 1367 1792 1368
rect 1786 1363 1787 1367
rect 1791 1363 1792 1367
rect 1786 1362 1792 1363
rect 1118 1352 1124 1353
rect 1118 1348 1119 1352
rect 1123 1348 1124 1352
rect 1118 1347 1124 1348
rect 1478 1352 1484 1353
rect 1478 1348 1479 1352
rect 1483 1348 1484 1352
rect 1478 1347 1484 1348
rect 1814 1352 1820 1353
rect 1814 1348 1815 1352
rect 1819 1348 1820 1352
rect 1814 1347 1820 1348
rect 1120 1323 1122 1347
rect 1480 1323 1482 1347
rect 1816 1323 1818 1347
rect 1119 1322 1123 1323
rect 1119 1317 1123 1318
rect 1151 1322 1155 1323
rect 1151 1317 1155 1318
rect 1327 1322 1331 1323
rect 1327 1317 1331 1318
rect 1479 1322 1483 1323
rect 1479 1317 1483 1318
rect 1495 1322 1499 1323
rect 1495 1317 1499 1318
rect 1663 1322 1667 1323
rect 1663 1317 1667 1318
rect 1815 1322 1819 1323
rect 1815 1317 1819 1318
rect 1152 1293 1154 1317
rect 1328 1293 1330 1317
rect 1496 1293 1498 1317
rect 1664 1293 1666 1317
rect 1816 1293 1818 1317
rect 1150 1292 1156 1293
rect 1150 1288 1151 1292
rect 1155 1288 1156 1292
rect 1150 1287 1156 1288
rect 1326 1292 1332 1293
rect 1326 1288 1327 1292
rect 1331 1288 1332 1292
rect 1326 1287 1332 1288
rect 1494 1292 1500 1293
rect 1494 1288 1495 1292
rect 1499 1288 1500 1292
rect 1494 1287 1500 1288
rect 1662 1292 1668 1293
rect 1662 1288 1663 1292
rect 1667 1288 1668 1292
rect 1662 1287 1668 1288
rect 1814 1292 1820 1293
rect 1814 1288 1815 1292
rect 1819 1288 1820 1292
rect 1814 1287 1820 1288
rect 1122 1277 1128 1278
rect 1122 1273 1123 1277
rect 1127 1273 1128 1277
rect 1122 1272 1128 1273
rect 1298 1277 1304 1278
rect 1298 1273 1299 1277
rect 1303 1273 1304 1277
rect 1298 1272 1304 1273
rect 1466 1277 1472 1278
rect 1466 1273 1467 1277
rect 1471 1273 1472 1277
rect 1466 1272 1472 1273
rect 1634 1277 1640 1278
rect 1634 1273 1635 1277
rect 1639 1273 1640 1277
rect 1634 1272 1640 1273
rect 1786 1277 1792 1278
rect 1786 1273 1787 1277
rect 1791 1273 1792 1277
rect 1786 1272 1792 1273
rect 1034 1227 1040 1228
rect 1034 1223 1035 1227
rect 1039 1223 1040 1227
rect 1034 1222 1040 1223
rect 1124 1199 1126 1272
rect 1250 1267 1256 1268
rect 1250 1263 1251 1267
rect 1255 1263 1256 1267
rect 1250 1262 1256 1263
rect 1252 1228 1254 1262
rect 1218 1227 1224 1228
rect 1218 1223 1219 1227
rect 1223 1223 1224 1227
rect 1218 1222 1224 1223
rect 1250 1227 1256 1228
rect 1250 1223 1251 1227
rect 1255 1223 1256 1227
rect 1250 1222 1256 1223
rect 939 1198 943 1199
rect 939 1193 943 1194
rect 1003 1198 1007 1199
rect 1003 1193 1007 1194
rect 1123 1198 1127 1199
rect 1123 1193 1127 1194
rect 1171 1198 1175 1199
rect 1171 1193 1175 1194
rect 870 1183 876 1184
rect 870 1179 871 1183
rect 875 1179 876 1183
rect 870 1178 876 1179
rect 1004 1132 1006 1193
rect 1010 1179 1016 1180
rect 1010 1175 1011 1179
rect 1015 1175 1016 1179
rect 1010 1174 1016 1175
rect 1012 1140 1014 1174
rect 1010 1139 1016 1140
rect 1010 1135 1011 1139
rect 1015 1135 1016 1139
rect 1010 1134 1016 1135
rect 1142 1139 1148 1140
rect 1142 1135 1143 1139
rect 1147 1135 1148 1139
rect 1142 1134 1148 1135
rect 834 1131 840 1132
rect 834 1127 835 1131
rect 839 1127 840 1131
rect 834 1126 840 1127
rect 1002 1131 1008 1132
rect 1002 1127 1003 1131
rect 1007 1127 1008 1131
rect 1002 1126 1008 1127
rect 862 1116 868 1117
rect 862 1112 863 1116
rect 867 1112 868 1116
rect 862 1111 868 1112
rect 1030 1116 1036 1117
rect 1030 1112 1031 1116
rect 1035 1112 1036 1116
rect 1030 1111 1036 1112
rect 864 1075 866 1111
rect 1032 1075 1034 1111
rect 863 1074 867 1075
rect 863 1069 867 1070
rect 951 1074 955 1075
rect 951 1069 955 1070
rect 1031 1074 1035 1075
rect 1031 1069 1035 1070
rect 952 1045 954 1069
rect 950 1044 956 1045
rect 950 1040 951 1044
rect 955 1040 956 1044
rect 950 1039 956 1040
rect 922 1029 928 1030
rect 922 1025 923 1029
rect 927 1025 928 1029
rect 922 1024 928 1025
rect 778 1019 784 1020
rect 778 1015 779 1019
rect 783 1015 784 1019
rect 778 1014 784 1015
rect 754 979 760 980
rect 754 975 755 979
rect 759 975 760 979
rect 754 974 760 975
rect 403 950 407 951
rect 403 945 407 946
rect 459 950 463 951
rect 459 945 463 946
rect 659 950 663 951
rect 659 945 663 946
rect 683 950 687 951
rect 683 945 687 946
rect 362 891 368 892
rect 362 887 363 891
rect 367 887 368 891
rect 362 886 368 887
rect 460 884 462 945
rect 498 891 504 892
rect 498 887 499 891
rect 503 887 504 891
rect 498 886 504 887
rect 458 883 464 884
rect 458 879 459 883
rect 463 879 464 883
rect 458 878 464 879
rect 486 868 492 869
rect 486 864 487 868
rect 491 864 492 868
rect 486 863 492 864
rect 488 823 490 863
rect 431 822 435 823
rect 431 817 435 818
rect 487 822 491 823
rect 487 817 491 818
rect 432 793 434 817
rect 430 792 436 793
rect 430 788 431 792
rect 435 788 436 792
rect 430 787 436 788
rect 402 777 408 778
rect 402 773 403 777
rect 407 773 408 777
rect 402 772 408 773
rect 270 767 276 768
rect 270 763 271 767
rect 275 763 276 767
rect 270 762 276 763
rect 242 727 248 728
rect 242 723 243 727
rect 247 723 248 727
rect 242 722 248 723
rect 111 710 115 711
rect 111 705 115 706
rect 131 710 135 711
rect 131 705 135 706
rect 147 710 151 711
rect 147 705 151 706
rect 112 645 114 705
rect 110 644 116 645
rect 132 644 134 705
rect 244 652 246 722
rect 404 711 406 772
rect 500 728 502 886
rect 684 884 686 945
rect 780 936 782 1014
rect 924 951 926 1024
rect 1002 1019 1008 1020
rect 1002 1015 1003 1019
rect 1007 1015 1008 1019
rect 1002 1014 1008 1015
rect 1134 1019 1140 1020
rect 1134 1015 1135 1019
rect 1139 1015 1140 1019
rect 1134 1014 1140 1015
rect 907 950 911 951
rect 907 945 911 946
rect 923 950 927 951
rect 923 945 927 946
rect 778 935 784 936
rect 778 931 779 935
rect 783 931 784 935
rect 778 930 784 931
rect 908 884 910 945
rect 1004 936 1006 1014
rect 1136 980 1138 1014
rect 1144 980 1146 1134
rect 1172 1132 1174 1193
rect 1220 1140 1222 1222
rect 1300 1199 1302 1272
rect 1426 1267 1432 1268
rect 1426 1263 1427 1267
rect 1431 1263 1432 1267
rect 1426 1262 1432 1263
rect 1428 1228 1430 1262
rect 1426 1227 1432 1228
rect 1426 1223 1427 1227
rect 1431 1223 1432 1227
rect 1426 1222 1432 1223
rect 1468 1199 1470 1272
rect 1594 1267 1600 1268
rect 1594 1263 1595 1267
rect 1599 1263 1600 1267
rect 1594 1262 1600 1263
rect 1596 1228 1598 1262
rect 1594 1227 1600 1228
rect 1594 1223 1595 1227
rect 1599 1223 1600 1227
rect 1594 1222 1600 1223
rect 1636 1199 1638 1272
rect 1762 1267 1768 1268
rect 1762 1263 1763 1267
rect 1767 1263 1768 1267
rect 1762 1262 1768 1263
rect 1764 1228 1766 1262
rect 1762 1227 1768 1228
rect 1762 1223 1763 1227
rect 1767 1223 1768 1227
rect 1762 1222 1768 1223
rect 1788 1199 1790 1272
rect 1884 1268 1886 1410
rect 1936 1369 1938 1429
rect 1976 1383 1978 1451
rect 1996 1383 1998 1452
rect 2122 1447 2128 1448
rect 2122 1443 2123 1447
rect 2127 1443 2128 1447
rect 2122 1442 2128 1443
rect 2124 1408 2126 1442
rect 2122 1407 2128 1408
rect 2122 1403 2123 1407
rect 2127 1403 2128 1407
rect 2122 1402 2128 1403
rect 2132 1383 2134 1452
rect 2258 1447 2264 1448
rect 2258 1443 2259 1447
rect 2263 1443 2264 1447
rect 2258 1442 2264 1443
rect 2260 1408 2262 1442
rect 2258 1407 2264 1408
rect 2258 1403 2259 1407
rect 2263 1403 2264 1407
rect 2258 1402 2264 1403
rect 2268 1383 2270 1452
rect 2394 1447 2400 1448
rect 2394 1443 2395 1447
rect 2399 1443 2400 1447
rect 2394 1442 2400 1443
rect 2396 1408 2398 1442
rect 2394 1407 2400 1408
rect 2394 1403 2395 1407
rect 2399 1403 2400 1407
rect 2394 1402 2400 1403
rect 2298 1399 2304 1400
rect 2298 1395 2299 1399
rect 2303 1395 2304 1399
rect 2298 1394 2304 1395
rect 1975 1382 1979 1383
rect 1975 1377 1979 1378
rect 1995 1382 1999 1383
rect 1995 1377 1999 1378
rect 2131 1382 2135 1383
rect 2131 1377 2135 1378
rect 2267 1382 2271 1383
rect 2267 1377 2271 1378
rect 2275 1382 2279 1383
rect 2275 1377 2279 1378
rect 1934 1368 1940 1369
rect 1934 1364 1935 1368
rect 1939 1364 1940 1368
rect 1934 1363 1940 1364
rect 1934 1351 1940 1352
rect 1934 1347 1935 1351
rect 1939 1347 1940 1351
rect 1934 1346 1940 1347
rect 1936 1323 1938 1346
rect 1935 1322 1939 1323
rect 1935 1317 1939 1318
rect 1976 1317 1978 1377
rect 1936 1294 1938 1317
rect 1974 1316 1980 1317
rect 1996 1316 1998 1377
rect 2276 1316 2278 1377
rect 2282 1363 2288 1364
rect 2282 1359 2283 1363
rect 2287 1359 2288 1363
rect 2282 1358 2288 1359
rect 2284 1324 2286 1358
rect 2300 1324 2302 1394
rect 2404 1383 2406 1452
rect 2530 1447 2536 1448
rect 2530 1443 2531 1447
rect 2535 1443 2536 1447
rect 2530 1442 2536 1443
rect 2532 1408 2534 1442
rect 2530 1407 2536 1408
rect 2530 1403 2531 1407
rect 2535 1403 2536 1407
rect 2530 1402 2536 1403
rect 2540 1383 2542 1452
rect 2656 1448 2658 1506
rect 2664 1503 2666 1547
rect 2800 1503 2802 1547
rect 2936 1503 2938 1547
rect 3072 1503 3074 1547
rect 3208 1503 3210 1547
rect 2663 1502 2667 1503
rect 2663 1497 2667 1498
rect 2703 1502 2707 1503
rect 2703 1497 2707 1498
rect 2799 1502 2803 1503
rect 2799 1497 2803 1498
rect 2839 1502 2843 1503
rect 2839 1497 2843 1498
rect 2935 1502 2939 1503
rect 2935 1497 2939 1498
rect 2975 1502 2979 1503
rect 2975 1497 2979 1498
rect 3071 1502 3075 1503
rect 3071 1497 3075 1498
rect 3207 1502 3211 1503
rect 3207 1497 3211 1498
rect 2704 1473 2706 1497
rect 2840 1473 2842 1497
rect 2976 1473 2978 1497
rect 2702 1472 2708 1473
rect 2702 1468 2703 1472
rect 2707 1468 2708 1472
rect 2702 1467 2708 1468
rect 2838 1472 2844 1473
rect 2838 1468 2839 1472
rect 2843 1468 2844 1472
rect 2838 1467 2844 1468
rect 2974 1472 2980 1473
rect 2974 1468 2975 1472
rect 2979 1468 2980 1472
rect 2974 1467 2980 1468
rect 2674 1457 2680 1458
rect 2674 1453 2675 1457
rect 2679 1453 2680 1457
rect 2674 1452 2680 1453
rect 2810 1457 2816 1458
rect 2810 1453 2811 1457
rect 2815 1453 2816 1457
rect 2810 1452 2816 1453
rect 2946 1457 2952 1458
rect 2946 1453 2947 1457
rect 2951 1453 2952 1457
rect 2946 1452 2952 1453
rect 2654 1447 2660 1448
rect 2654 1443 2655 1447
rect 2659 1443 2660 1447
rect 2654 1442 2660 1443
rect 2676 1383 2678 1452
rect 2802 1447 2808 1448
rect 2802 1443 2803 1447
rect 2807 1443 2808 1447
rect 2802 1442 2808 1443
rect 2770 1439 2776 1440
rect 2770 1435 2771 1439
rect 2775 1435 2776 1439
rect 2770 1434 2776 1435
rect 2772 1408 2774 1434
rect 2804 1408 2806 1442
rect 2770 1407 2776 1408
rect 2770 1403 2771 1407
rect 2775 1403 2776 1407
rect 2770 1402 2776 1403
rect 2802 1407 2808 1408
rect 2802 1403 2803 1407
rect 2807 1403 2808 1407
rect 2802 1402 2808 1403
rect 2812 1383 2814 1452
rect 2934 1447 2940 1448
rect 2934 1443 2935 1447
rect 2939 1443 2940 1447
rect 2934 1442 2940 1443
rect 2403 1382 2407 1383
rect 2403 1377 2407 1378
rect 2539 1382 2543 1383
rect 2539 1377 2543 1378
rect 2563 1382 2567 1383
rect 2563 1377 2567 1378
rect 2675 1382 2679 1383
rect 2675 1377 2679 1378
rect 2811 1382 2815 1383
rect 2811 1377 2815 1378
rect 2843 1382 2847 1383
rect 2843 1377 2847 1378
rect 2282 1323 2288 1324
rect 2282 1319 2283 1323
rect 2287 1319 2288 1323
rect 2282 1318 2288 1319
rect 2298 1323 2304 1324
rect 2298 1319 2299 1323
rect 2303 1319 2304 1323
rect 2298 1318 2304 1319
rect 2564 1316 2566 1377
rect 2686 1323 2692 1324
rect 2686 1319 2687 1323
rect 2691 1319 2692 1323
rect 2686 1318 2692 1319
rect 1974 1312 1975 1316
rect 1979 1312 1980 1316
rect 1974 1311 1980 1312
rect 1994 1315 2000 1316
rect 1994 1311 1995 1315
rect 1999 1311 2000 1315
rect 1994 1310 2000 1311
rect 2274 1315 2280 1316
rect 2274 1311 2275 1315
rect 2279 1311 2280 1315
rect 2274 1310 2280 1311
rect 2562 1315 2568 1316
rect 2562 1311 2563 1315
rect 2567 1311 2568 1315
rect 2562 1310 2568 1311
rect 2022 1300 2028 1301
rect 1974 1299 1980 1300
rect 1974 1295 1975 1299
rect 1979 1295 1980 1299
rect 2022 1296 2023 1300
rect 2027 1296 2028 1300
rect 2022 1295 2028 1296
rect 2302 1300 2308 1301
rect 2302 1296 2303 1300
rect 2307 1296 2308 1300
rect 2302 1295 2308 1296
rect 2590 1300 2596 1301
rect 2590 1296 2591 1300
rect 2595 1296 2596 1300
rect 2590 1295 2596 1296
rect 1974 1294 1980 1295
rect 1934 1293 1940 1294
rect 1934 1289 1935 1293
rect 1939 1289 1940 1293
rect 1934 1288 1940 1289
rect 1934 1276 1940 1277
rect 1934 1272 1935 1276
rect 1939 1272 1940 1276
rect 1934 1271 1940 1272
rect 1882 1267 1888 1268
rect 1882 1263 1883 1267
rect 1887 1263 1888 1267
rect 1882 1262 1888 1263
rect 1936 1199 1938 1271
rect 1976 1247 1978 1294
rect 2024 1247 2026 1295
rect 2304 1247 2306 1295
rect 2592 1247 2594 1295
rect 1975 1246 1979 1247
rect 1975 1241 1979 1242
rect 2023 1246 2027 1247
rect 2023 1241 2027 1242
rect 2303 1246 2307 1247
rect 2303 1241 2307 1242
rect 2591 1246 2595 1247
rect 2591 1241 2595 1242
rect 2655 1246 2659 1247
rect 2655 1241 2659 1242
rect 1976 1218 1978 1241
rect 1974 1217 1980 1218
rect 2656 1217 2658 1241
rect 1974 1213 1975 1217
rect 1979 1213 1980 1217
rect 1974 1212 1980 1213
rect 2654 1216 2660 1217
rect 2654 1212 2655 1216
rect 2659 1212 2660 1216
rect 2654 1211 2660 1212
rect 2626 1201 2632 1202
rect 1974 1200 1980 1201
rect 1299 1198 1303 1199
rect 1299 1193 1303 1194
rect 1331 1198 1335 1199
rect 1331 1193 1335 1194
rect 1467 1198 1471 1199
rect 1467 1193 1471 1194
rect 1491 1198 1495 1199
rect 1491 1193 1495 1194
rect 1635 1198 1639 1199
rect 1635 1193 1639 1194
rect 1651 1198 1655 1199
rect 1651 1193 1655 1194
rect 1787 1198 1791 1199
rect 1787 1193 1791 1194
rect 1935 1198 1939 1199
rect 1974 1196 1975 1200
rect 1979 1196 1980 1200
rect 2626 1197 2627 1201
rect 2631 1197 2632 1201
rect 2626 1196 2632 1197
rect 1974 1195 1980 1196
rect 1935 1193 1939 1194
rect 1218 1139 1224 1140
rect 1218 1135 1219 1139
rect 1223 1135 1224 1139
rect 1218 1134 1224 1135
rect 1332 1132 1334 1193
rect 1482 1183 1488 1184
rect 1482 1179 1483 1183
rect 1487 1179 1488 1183
rect 1482 1178 1488 1179
rect 1484 1140 1486 1178
rect 1482 1139 1488 1140
rect 1482 1135 1483 1139
rect 1487 1135 1488 1139
rect 1482 1134 1488 1135
rect 1492 1132 1494 1193
rect 1652 1132 1654 1193
rect 1746 1179 1752 1180
rect 1746 1175 1747 1179
rect 1751 1175 1752 1179
rect 1746 1174 1752 1175
rect 1748 1148 1750 1174
rect 1746 1147 1752 1148
rect 1746 1143 1747 1147
rect 1751 1143 1752 1147
rect 1746 1142 1752 1143
rect 1788 1132 1790 1193
rect 1936 1133 1938 1193
rect 1934 1132 1940 1133
rect 1170 1131 1176 1132
rect 1170 1127 1171 1131
rect 1175 1127 1176 1131
rect 1170 1126 1176 1127
rect 1330 1131 1336 1132
rect 1330 1127 1331 1131
rect 1335 1127 1336 1131
rect 1330 1126 1336 1127
rect 1490 1131 1496 1132
rect 1490 1127 1491 1131
rect 1495 1127 1496 1131
rect 1490 1126 1496 1127
rect 1650 1131 1656 1132
rect 1650 1127 1651 1131
rect 1655 1127 1656 1131
rect 1650 1126 1656 1127
rect 1786 1131 1792 1132
rect 1786 1127 1787 1131
rect 1791 1127 1792 1131
rect 1934 1128 1935 1132
rect 1939 1128 1940 1132
rect 1934 1127 1940 1128
rect 1786 1126 1792 1127
rect 1976 1119 1978 1195
rect 2118 1183 2124 1184
rect 2118 1179 2119 1183
rect 2123 1179 2124 1183
rect 2118 1178 2124 1179
rect 2266 1183 2272 1184
rect 2266 1179 2267 1183
rect 2271 1179 2272 1183
rect 2266 1178 2272 1179
rect 1975 1118 1979 1119
rect 1198 1116 1204 1117
rect 1198 1112 1199 1116
rect 1203 1112 1204 1116
rect 1198 1111 1204 1112
rect 1358 1116 1364 1117
rect 1358 1112 1359 1116
rect 1363 1112 1364 1116
rect 1358 1111 1364 1112
rect 1518 1116 1524 1117
rect 1518 1112 1519 1116
rect 1523 1112 1524 1116
rect 1518 1111 1524 1112
rect 1678 1116 1684 1117
rect 1678 1112 1679 1116
rect 1683 1112 1684 1116
rect 1678 1111 1684 1112
rect 1814 1116 1820 1117
rect 1814 1112 1815 1116
rect 1819 1112 1820 1116
rect 1814 1111 1820 1112
rect 1934 1115 1940 1116
rect 1934 1111 1935 1115
rect 1939 1111 1940 1115
rect 1975 1113 1979 1114
rect 1995 1118 1999 1119
rect 1995 1113 1999 1114
rect 1200 1075 1202 1111
rect 1360 1075 1362 1111
rect 1520 1075 1522 1111
rect 1680 1075 1682 1111
rect 1816 1075 1818 1111
rect 1934 1110 1940 1111
rect 1936 1075 1938 1110
rect 1199 1074 1203 1075
rect 1199 1069 1203 1070
rect 1215 1074 1219 1075
rect 1215 1069 1219 1070
rect 1359 1074 1363 1075
rect 1359 1069 1363 1070
rect 1519 1074 1523 1075
rect 1519 1069 1523 1070
rect 1679 1074 1683 1075
rect 1679 1069 1683 1070
rect 1815 1074 1819 1075
rect 1815 1069 1819 1070
rect 1935 1074 1939 1075
rect 1935 1069 1939 1070
rect 1216 1045 1218 1069
rect 1936 1046 1938 1069
rect 1976 1053 1978 1113
rect 1974 1052 1980 1053
rect 1996 1052 1998 1113
rect 2090 1099 2096 1100
rect 2090 1095 2091 1099
rect 2095 1095 2096 1099
rect 2090 1094 2096 1095
rect 1974 1048 1975 1052
rect 1979 1048 1980 1052
rect 1974 1047 1980 1048
rect 1994 1051 2000 1052
rect 1994 1047 1995 1051
rect 1999 1047 2000 1051
rect 1994 1046 2000 1047
rect 1934 1045 1940 1046
rect 1214 1044 1220 1045
rect 1214 1040 1215 1044
rect 1219 1040 1220 1044
rect 1934 1041 1935 1045
rect 1939 1041 1940 1045
rect 1934 1040 1940 1041
rect 1214 1039 1220 1040
rect 2022 1036 2028 1037
rect 1974 1035 1980 1036
rect 1974 1031 1975 1035
rect 1979 1031 1980 1035
rect 2022 1032 2023 1036
rect 2027 1032 2028 1036
rect 2022 1031 2028 1032
rect 1974 1030 1980 1031
rect 1186 1029 1192 1030
rect 1186 1025 1187 1029
rect 1191 1025 1192 1029
rect 1186 1024 1192 1025
rect 1934 1028 1940 1029
rect 1934 1024 1935 1028
rect 1939 1024 1940 1028
rect 1134 979 1140 980
rect 1134 975 1135 979
rect 1139 975 1140 979
rect 1134 974 1140 975
rect 1142 979 1148 980
rect 1142 975 1143 979
rect 1147 975 1148 979
rect 1142 974 1148 975
rect 1188 951 1190 1024
rect 1934 1023 1940 1024
rect 1936 951 1938 1023
rect 1976 1007 1978 1030
rect 2024 1007 2026 1031
rect 1975 1006 1979 1007
rect 1975 1001 1979 1002
rect 2023 1006 2027 1007
rect 2023 1001 2027 1002
rect 1976 978 1978 1001
rect 1974 977 1980 978
rect 2024 977 2026 1001
rect 1974 973 1975 977
rect 1979 973 1980 977
rect 1974 972 1980 973
rect 2022 976 2028 977
rect 2022 972 2023 976
rect 2027 972 2028 976
rect 2022 971 2028 972
rect 1994 961 2000 962
rect 1974 960 1980 961
rect 1974 956 1975 960
rect 1979 956 1980 960
rect 1994 957 1995 961
rect 1999 957 2000 961
rect 1994 956 2000 957
rect 1974 955 1980 956
rect 1131 950 1135 951
rect 1131 945 1135 946
rect 1187 950 1191 951
rect 1187 945 1191 946
rect 1363 950 1367 951
rect 1363 945 1367 946
rect 1935 950 1939 951
rect 1935 945 1939 946
rect 1002 935 1008 936
rect 1002 931 1003 935
rect 1007 931 1008 935
rect 1002 930 1008 931
rect 1132 884 1134 945
rect 1138 931 1144 932
rect 1138 927 1139 931
rect 1143 927 1144 931
rect 1138 926 1144 927
rect 1140 892 1142 926
rect 1138 891 1144 892
rect 1138 887 1139 891
rect 1143 887 1144 891
rect 1138 886 1144 887
rect 1364 884 1366 945
rect 1370 931 1376 932
rect 1370 927 1371 931
rect 1375 927 1376 931
rect 1370 926 1376 927
rect 1372 892 1374 926
rect 1370 891 1376 892
rect 1370 887 1371 891
rect 1375 887 1376 891
rect 1370 886 1376 887
rect 1490 891 1496 892
rect 1490 887 1491 891
rect 1495 887 1496 891
rect 1490 886 1496 887
rect 682 883 688 884
rect 682 879 683 883
rect 687 879 688 883
rect 682 878 688 879
rect 906 883 912 884
rect 906 879 907 883
rect 911 879 912 883
rect 906 878 912 879
rect 1130 883 1136 884
rect 1130 879 1131 883
rect 1135 879 1136 883
rect 1130 878 1136 879
rect 1362 883 1368 884
rect 1362 879 1363 883
rect 1367 879 1368 883
rect 1362 878 1368 879
rect 710 868 716 869
rect 710 864 711 868
rect 715 864 716 868
rect 710 863 716 864
rect 934 868 940 869
rect 934 864 935 868
rect 939 864 940 868
rect 934 863 940 864
rect 1158 868 1164 869
rect 1158 864 1159 868
rect 1163 864 1164 868
rect 1158 863 1164 864
rect 1390 868 1396 869
rect 1390 864 1391 868
rect 1395 864 1396 868
rect 1390 863 1396 864
rect 712 823 714 863
rect 936 823 938 863
rect 1160 823 1162 863
rect 1392 823 1394 863
rect 671 822 675 823
rect 671 817 675 818
rect 711 822 715 823
rect 711 817 715 818
rect 903 822 907 823
rect 903 817 907 818
rect 935 822 939 823
rect 935 817 939 818
rect 1127 822 1131 823
rect 1127 817 1131 818
rect 1159 822 1163 823
rect 1159 817 1163 818
rect 1351 822 1355 823
rect 1351 817 1355 818
rect 1391 822 1395 823
rect 1391 817 1395 818
rect 672 793 674 817
rect 904 793 906 817
rect 1128 793 1130 817
rect 1352 793 1354 817
rect 670 792 676 793
rect 670 788 671 792
rect 675 788 676 792
rect 670 787 676 788
rect 902 792 908 793
rect 902 788 903 792
rect 907 788 908 792
rect 902 787 908 788
rect 1126 792 1132 793
rect 1126 788 1127 792
rect 1131 788 1132 792
rect 1126 787 1132 788
rect 1350 792 1356 793
rect 1350 788 1351 792
rect 1355 788 1356 792
rect 1350 787 1356 788
rect 642 777 648 778
rect 642 773 643 777
rect 647 773 648 777
rect 642 772 648 773
rect 874 777 880 778
rect 874 773 875 777
rect 879 773 880 777
rect 874 772 880 773
rect 1098 777 1104 778
rect 1098 773 1099 777
rect 1103 773 1104 777
rect 1098 772 1104 773
rect 1322 777 1328 778
rect 1322 773 1323 777
rect 1327 773 1328 777
rect 1322 772 1328 773
rect 530 767 536 768
rect 530 763 531 767
rect 535 763 536 767
rect 530 762 536 763
rect 532 728 534 762
rect 498 727 504 728
rect 498 723 499 727
rect 503 723 504 727
rect 498 722 504 723
rect 530 727 536 728
rect 530 723 531 727
rect 535 723 536 727
rect 530 722 536 723
rect 644 711 646 772
rect 766 767 772 768
rect 766 763 767 767
rect 771 763 772 767
rect 766 762 772 763
rect 315 710 319 711
rect 315 705 319 706
rect 403 710 407 711
rect 403 705 407 706
rect 523 710 527 711
rect 523 705 527 706
rect 643 710 647 711
rect 643 705 647 706
rect 723 710 727 711
rect 723 705 727 706
rect 306 695 312 696
rect 306 691 307 695
rect 311 691 312 695
rect 306 690 312 691
rect 308 652 310 690
rect 242 651 248 652
rect 242 647 243 651
rect 247 647 248 651
rect 242 646 248 647
rect 306 651 312 652
rect 306 647 307 651
rect 311 647 312 651
rect 306 646 312 647
rect 316 644 318 705
rect 410 691 416 692
rect 410 687 411 691
rect 415 687 416 691
rect 410 686 416 687
rect 110 640 111 644
rect 115 640 116 644
rect 110 639 116 640
rect 130 643 136 644
rect 130 639 131 643
rect 135 639 136 643
rect 130 638 136 639
rect 314 643 320 644
rect 314 639 315 643
rect 319 639 320 643
rect 314 638 320 639
rect 158 628 164 629
rect 110 627 116 628
rect 110 623 111 627
rect 115 623 116 627
rect 158 624 159 628
rect 163 624 164 628
rect 158 623 164 624
rect 342 628 348 629
rect 342 624 343 628
rect 347 624 348 628
rect 342 623 348 624
rect 110 622 116 623
rect 112 599 114 622
rect 160 599 162 623
rect 344 599 346 623
rect 111 598 115 599
rect 111 593 115 594
rect 159 598 163 599
rect 159 593 163 594
rect 343 598 347 599
rect 343 593 347 594
rect 375 598 379 599
rect 375 593 379 594
rect 112 570 114 593
rect 110 569 116 570
rect 160 569 162 593
rect 376 569 378 593
rect 110 565 111 569
rect 115 565 116 569
rect 110 564 116 565
rect 158 568 164 569
rect 158 564 159 568
rect 163 564 164 568
rect 158 563 164 564
rect 374 568 380 569
rect 374 564 375 568
rect 379 564 380 568
rect 374 563 380 564
rect 130 553 136 554
rect 110 552 116 553
rect 110 548 111 552
rect 115 548 116 552
rect 130 549 131 553
rect 135 549 136 553
rect 130 548 136 549
rect 346 553 352 554
rect 346 549 347 553
rect 351 549 352 553
rect 346 548 352 549
rect 110 547 116 548
rect 112 487 114 547
rect 132 487 134 548
rect 254 543 260 544
rect 254 539 255 543
rect 259 539 260 543
rect 254 538 260 539
rect 256 504 258 538
rect 226 503 232 504
rect 226 499 227 503
rect 231 499 232 503
rect 226 498 232 499
rect 254 503 260 504
rect 254 499 255 503
rect 259 499 260 503
rect 254 498 260 499
rect 111 486 115 487
rect 111 481 115 482
rect 131 486 135 487
rect 131 481 135 482
rect 155 486 159 487
rect 155 481 159 482
rect 112 421 114 481
rect 110 420 116 421
rect 156 420 158 481
rect 228 428 230 498
rect 348 487 350 548
rect 412 544 414 686
rect 524 644 526 705
rect 618 691 624 692
rect 618 687 619 691
rect 623 687 624 691
rect 618 686 624 687
rect 620 660 622 686
rect 618 659 624 660
rect 618 655 619 659
rect 623 655 624 659
rect 618 654 624 655
rect 646 651 652 652
rect 646 647 647 651
rect 651 647 652 651
rect 646 646 652 647
rect 522 643 528 644
rect 522 639 523 643
rect 527 639 528 643
rect 522 638 528 639
rect 550 628 556 629
rect 550 624 551 628
rect 555 624 556 628
rect 550 623 556 624
rect 552 599 554 623
rect 551 598 555 599
rect 551 593 555 594
rect 599 598 603 599
rect 599 593 603 594
rect 600 569 602 593
rect 598 568 604 569
rect 598 564 599 568
rect 603 564 604 568
rect 598 563 604 564
rect 570 553 576 554
rect 570 549 571 553
rect 575 549 576 553
rect 570 548 576 549
rect 410 543 416 544
rect 410 539 411 543
rect 415 539 416 543
rect 410 538 416 539
rect 572 487 574 548
rect 648 504 650 646
rect 724 644 726 705
rect 768 696 770 762
rect 876 711 878 772
rect 1062 767 1068 768
rect 1062 763 1063 767
rect 1067 763 1068 767
rect 1062 762 1068 763
rect 1064 728 1066 762
rect 1062 727 1068 728
rect 1062 723 1063 727
rect 1067 723 1068 727
rect 1062 722 1068 723
rect 1100 711 1102 772
rect 1324 711 1326 772
rect 1482 767 1488 768
rect 1482 763 1483 767
rect 1487 763 1488 767
rect 1482 762 1488 763
rect 1484 728 1486 762
rect 1492 728 1494 886
rect 1936 885 1938 945
rect 1976 891 1978 955
rect 1996 891 1998 956
rect 2092 952 2094 1094
rect 2120 1060 2122 1178
rect 2171 1118 2175 1119
rect 2171 1113 2175 1114
rect 2118 1059 2124 1060
rect 2118 1055 2119 1059
rect 2123 1055 2124 1059
rect 2118 1054 2124 1055
rect 2172 1052 2174 1113
rect 2268 1104 2270 1178
rect 2628 1119 2630 1196
rect 2688 1152 2690 1318
rect 2844 1316 2846 1377
rect 2936 1368 2938 1442
rect 2948 1383 2950 1452
rect 3300 1408 3302 1570
rect 3800 1569 3802 1629
rect 3840 1569 3842 1629
rect 3798 1568 3804 1569
rect 3798 1564 3799 1568
rect 3803 1564 3804 1568
rect 3798 1563 3804 1564
rect 3838 1568 3844 1569
rect 3860 1568 3862 1629
rect 3954 1615 3960 1616
rect 3954 1611 3955 1615
rect 3959 1611 3960 1615
rect 3954 1610 3960 1611
rect 3956 1584 3958 1610
rect 3954 1583 3960 1584
rect 3954 1579 3955 1583
rect 3959 1579 3960 1583
rect 3954 1578 3960 1579
rect 3996 1568 3998 1629
rect 4002 1615 4008 1616
rect 4002 1611 4003 1615
rect 4007 1611 4008 1615
rect 4002 1610 4008 1611
rect 4004 1576 4006 1610
rect 4148 1576 4150 1646
rect 4276 1635 4278 1696
rect 4434 1691 4440 1692
rect 4434 1687 4435 1691
rect 4439 1687 4440 1691
rect 4434 1686 4440 1687
rect 4370 1683 4376 1684
rect 4370 1679 4371 1683
rect 4375 1679 4376 1683
rect 4370 1678 4376 1679
rect 4372 1652 4374 1678
rect 4436 1652 4438 1686
rect 4370 1651 4376 1652
rect 4370 1647 4371 1651
rect 4375 1647 4376 1651
rect 4370 1646 4376 1647
rect 4434 1651 4440 1652
rect 4434 1647 4435 1651
rect 4439 1647 4440 1651
rect 4434 1646 4440 1647
rect 4508 1635 4510 1696
rect 4634 1691 4640 1692
rect 4634 1687 4635 1691
rect 4639 1687 4640 1691
rect 4634 1686 4640 1687
rect 4636 1652 4638 1686
rect 4634 1651 4640 1652
rect 4634 1647 4635 1651
rect 4639 1647 4640 1651
rect 4634 1646 4640 1647
rect 4748 1635 4750 1696
rect 4870 1691 4876 1692
rect 4870 1687 4871 1691
rect 4875 1687 4876 1691
rect 4870 1686 4876 1687
rect 4155 1634 4159 1635
rect 4155 1629 4159 1630
rect 4275 1634 4279 1635
rect 4275 1629 4279 1630
rect 4355 1634 4359 1635
rect 4355 1629 4359 1630
rect 4507 1634 4511 1635
rect 4507 1629 4511 1630
rect 4587 1634 4591 1635
rect 4587 1629 4591 1630
rect 4747 1634 4751 1635
rect 4747 1629 4751 1630
rect 4851 1634 4855 1635
rect 4851 1629 4855 1630
rect 4002 1575 4008 1576
rect 4002 1571 4003 1575
rect 4007 1571 4008 1575
rect 4002 1570 4008 1571
rect 4122 1575 4128 1576
rect 4122 1571 4123 1575
rect 4127 1571 4128 1575
rect 4122 1570 4128 1571
rect 4146 1575 4152 1576
rect 4146 1571 4147 1575
rect 4151 1571 4152 1575
rect 4146 1570 4152 1571
rect 3838 1564 3839 1568
rect 3843 1564 3844 1568
rect 3838 1563 3844 1564
rect 3858 1567 3864 1568
rect 3858 1563 3859 1567
rect 3863 1563 3864 1567
rect 3858 1562 3864 1563
rect 3994 1567 4000 1568
rect 3994 1563 3995 1567
rect 3999 1563 4000 1567
rect 3994 1562 4000 1563
rect 3886 1552 3892 1553
rect 3798 1551 3804 1552
rect 3798 1547 3799 1551
rect 3803 1547 3804 1551
rect 3798 1546 3804 1547
rect 3838 1551 3844 1552
rect 3838 1547 3839 1551
rect 3843 1547 3844 1551
rect 3886 1548 3887 1552
rect 3891 1548 3892 1552
rect 3886 1547 3892 1548
rect 4022 1552 4028 1553
rect 4022 1548 4023 1552
rect 4027 1548 4028 1552
rect 4022 1547 4028 1548
rect 3838 1546 3844 1547
rect 3800 1503 3802 1546
rect 3840 1523 3842 1546
rect 3888 1523 3890 1547
rect 4024 1523 4026 1547
rect 3839 1522 3843 1523
rect 3839 1517 3843 1518
rect 3887 1522 3891 1523
rect 3887 1517 3891 1518
rect 4023 1522 4027 1523
rect 4023 1517 4027 1518
rect 3799 1502 3803 1503
rect 3799 1497 3803 1498
rect 3800 1474 3802 1497
rect 3840 1494 3842 1517
rect 3838 1493 3844 1494
rect 3888 1493 3890 1517
rect 4024 1493 4026 1517
rect 4124 1508 4126 1570
rect 4156 1568 4158 1629
rect 4250 1615 4256 1616
rect 4250 1611 4251 1615
rect 4255 1611 4256 1615
rect 4250 1610 4256 1611
rect 4154 1567 4160 1568
rect 4154 1563 4155 1567
rect 4159 1563 4160 1567
rect 4154 1562 4160 1563
rect 4182 1552 4188 1553
rect 4182 1548 4183 1552
rect 4187 1548 4188 1552
rect 4182 1547 4188 1548
rect 4184 1523 4186 1547
rect 4159 1522 4163 1523
rect 4159 1517 4163 1518
rect 4183 1522 4187 1523
rect 4183 1517 4187 1518
rect 4122 1507 4128 1508
rect 4122 1503 4123 1507
rect 4127 1503 4128 1507
rect 4122 1502 4128 1503
rect 4160 1493 4162 1517
rect 3838 1489 3839 1493
rect 3843 1489 3844 1493
rect 3838 1488 3844 1489
rect 3886 1492 3892 1493
rect 3886 1488 3887 1492
rect 3891 1488 3892 1492
rect 3886 1487 3892 1488
rect 4022 1492 4028 1493
rect 4022 1488 4023 1492
rect 4027 1488 4028 1492
rect 4022 1487 4028 1488
rect 4158 1492 4164 1493
rect 4158 1488 4159 1492
rect 4163 1488 4164 1492
rect 4158 1487 4164 1488
rect 3858 1477 3864 1478
rect 3838 1476 3844 1477
rect 3798 1473 3804 1474
rect 3798 1469 3799 1473
rect 3803 1469 3804 1473
rect 3838 1472 3839 1476
rect 3843 1472 3844 1476
rect 3858 1473 3859 1477
rect 3863 1473 3864 1477
rect 3858 1472 3864 1473
rect 3994 1477 4000 1478
rect 3994 1473 3995 1477
rect 3999 1473 4000 1477
rect 3994 1472 4000 1473
rect 4130 1477 4136 1478
rect 4130 1473 4131 1477
rect 4135 1473 4136 1477
rect 4130 1472 4136 1473
rect 3838 1471 3844 1472
rect 3798 1468 3804 1469
rect 3798 1456 3804 1457
rect 3798 1452 3799 1456
rect 3803 1452 3804 1456
rect 3798 1451 3804 1452
rect 3298 1407 3304 1408
rect 3298 1403 3299 1407
rect 3303 1403 3304 1407
rect 3298 1402 3304 1403
rect 3778 1391 3784 1392
rect 3778 1387 3779 1391
rect 3783 1387 3784 1391
rect 3778 1386 3784 1387
rect 2947 1382 2951 1383
rect 2947 1377 2951 1378
rect 3123 1382 3127 1383
rect 3123 1377 3127 1378
rect 3395 1382 3399 1383
rect 3395 1377 3399 1378
rect 3651 1382 3655 1383
rect 3651 1377 3655 1378
rect 2934 1367 2940 1368
rect 2934 1363 2935 1367
rect 2939 1363 2940 1367
rect 2934 1362 2940 1363
rect 3124 1316 3126 1377
rect 3370 1367 3376 1368
rect 3370 1363 3371 1367
rect 3375 1363 3376 1367
rect 3370 1362 3376 1363
rect 2842 1315 2848 1316
rect 2842 1311 2843 1315
rect 2847 1311 2848 1315
rect 2842 1310 2848 1311
rect 3122 1315 3128 1316
rect 3122 1311 3123 1315
rect 3127 1311 3128 1315
rect 3122 1310 3128 1311
rect 2870 1300 2876 1301
rect 2870 1296 2871 1300
rect 2875 1296 2876 1300
rect 2870 1295 2876 1296
rect 3150 1300 3156 1301
rect 3150 1296 3151 1300
rect 3155 1296 3156 1300
rect 3150 1295 3156 1296
rect 2872 1247 2874 1295
rect 3152 1247 3154 1295
rect 2831 1246 2835 1247
rect 2831 1241 2835 1242
rect 2871 1246 2875 1247
rect 2871 1241 2875 1242
rect 3007 1246 3011 1247
rect 3007 1241 3011 1242
rect 3151 1246 3155 1247
rect 3151 1241 3155 1242
rect 3183 1246 3187 1247
rect 3183 1241 3187 1242
rect 3359 1246 3363 1247
rect 3359 1241 3363 1242
rect 2832 1217 2834 1241
rect 3008 1217 3010 1241
rect 3184 1217 3186 1241
rect 3360 1217 3362 1241
rect 2830 1216 2836 1217
rect 2830 1212 2831 1216
rect 2835 1212 2836 1216
rect 2830 1211 2836 1212
rect 3006 1216 3012 1217
rect 3006 1212 3007 1216
rect 3011 1212 3012 1216
rect 3006 1211 3012 1212
rect 3182 1216 3188 1217
rect 3182 1212 3183 1216
rect 3187 1212 3188 1216
rect 3182 1211 3188 1212
rect 3358 1216 3364 1217
rect 3358 1212 3359 1216
rect 3363 1212 3364 1216
rect 3358 1211 3364 1212
rect 2802 1201 2808 1202
rect 2802 1197 2803 1201
rect 2807 1197 2808 1201
rect 2802 1196 2808 1197
rect 2978 1201 2984 1202
rect 2978 1197 2979 1201
rect 2983 1197 2984 1201
rect 2978 1196 2984 1197
rect 3154 1201 3160 1202
rect 3154 1197 3155 1201
rect 3159 1197 3160 1201
rect 3154 1196 3160 1197
rect 3330 1201 3336 1202
rect 3330 1197 3331 1201
rect 3335 1197 3336 1201
rect 3330 1196 3336 1197
rect 2754 1191 2760 1192
rect 2754 1187 2755 1191
rect 2759 1187 2760 1191
rect 2754 1186 2760 1187
rect 2756 1152 2758 1186
rect 2686 1151 2692 1152
rect 2686 1147 2687 1151
rect 2691 1147 2692 1151
rect 2686 1146 2692 1147
rect 2754 1151 2760 1152
rect 2754 1147 2755 1151
rect 2759 1147 2760 1151
rect 2754 1146 2760 1147
rect 2804 1119 2806 1196
rect 2980 1119 2982 1196
rect 3156 1119 3158 1196
rect 3282 1191 3288 1192
rect 3282 1187 3283 1191
rect 3287 1187 3288 1191
rect 3282 1186 3288 1187
rect 3284 1152 3286 1186
rect 3282 1151 3288 1152
rect 3282 1147 3283 1151
rect 3287 1147 3288 1151
rect 3282 1146 3288 1147
rect 3234 1143 3240 1144
rect 3234 1139 3235 1143
rect 3239 1139 3240 1143
rect 3234 1138 3240 1139
rect 2363 1118 2367 1119
rect 2363 1113 2367 1114
rect 2547 1118 2551 1119
rect 2547 1113 2551 1114
rect 2627 1118 2631 1119
rect 2627 1113 2631 1114
rect 2723 1118 2727 1119
rect 2723 1113 2727 1114
rect 2803 1118 2807 1119
rect 2803 1113 2807 1114
rect 2891 1118 2895 1119
rect 2891 1113 2895 1114
rect 2979 1118 2983 1119
rect 2979 1113 2983 1114
rect 3059 1118 3063 1119
rect 3059 1113 3063 1114
rect 3155 1118 3159 1119
rect 3155 1113 3159 1114
rect 3219 1118 3223 1119
rect 3219 1113 3223 1114
rect 2266 1103 2272 1104
rect 2266 1099 2267 1103
rect 2271 1099 2272 1103
rect 2266 1098 2272 1099
rect 2364 1052 2366 1113
rect 2370 1099 2376 1100
rect 2370 1095 2371 1099
rect 2375 1095 2376 1099
rect 2370 1094 2376 1095
rect 2372 1060 2374 1094
rect 2370 1059 2376 1060
rect 2370 1055 2371 1059
rect 2375 1055 2376 1059
rect 2370 1054 2376 1055
rect 2490 1059 2496 1060
rect 2490 1055 2491 1059
rect 2495 1055 2496 1059
rect 2490 1054 2496 1055
rect 2170 1051 2176 1052
rect 2170 1047 2171 1051
rect 2175 1047 2176 1051
rect 2170 1046 2176 1047
rect 2362 1051 2368 1052
rect 2362 1047 2363 1051
rect 2367 1047 2368 1051
rect 2362 1046 2368 1047
rect 2198 1036 2204 1037
rect 2198 1032 2199 1036
rect 2203 1032 2204 1036
rect 2198 1031 2204 1032
rect 2390 1036 2396 1037
rect 2390 1032 2391 1036
rect 2395 1032 2396 1036
rect 2390 1031 2396 1032
rect 2200 1007 2202 1031
rect 2392 1007 2394 1031
rect 2191 1006 2195 1007
rect 2191 1001 2195 1002
rect 2199 1006 2203 1007
rect 2199 1001 2203 1002
rect 2375 1006 2379 1007
rect 2375 1001 2379 1002
rect 2391 1006 2395 1007
rect 2391 1001 2395 1002
rect 2192 977 2194 1001
rect 2376 977 2378 1001
rect 2190 976 2196 977
rect 2190 972 2191 976
rect 2195 972 2196 976
rect 2190 971 2196 972
rect 2374 976 2380 977
rect 2374 972 2375 976
rect 2379 972 2380 976
rect 2374 971 2380 972
rect 2162 961 2168 962
rect 2162 957 2163 961
rect 2167 957 2168 961
rect 2162 956 2168 957
rect 2346 961 2352 962
rect 2346 957 2347 961
rect 2351 957 2352 961
rect 2346 956 2352 957
rect 2090 951 2096 952
rect 2090 947 2091 951
rect 2095 947 2096 951
rect 2090 946 2096 947
rect 2154 951 2160 952
rect 2154 947 2155 951
rect 2159 947 2160 951
rect 2154 946 2160 947
rect 2156 912 2158 946
rect 2154 911 2160 912
rect 2154 907 2155 911
rect 2159 907 2160 911
rect 2154 906 2160 907
rect 2164 891 2166 956
rect 2348 891 2350 956
rect 2492 912 2494 1054
rect 2548 1052 2550 1113
rect 2642 1099 2648 1100
rect 2642 1095 2643 1099
rect 2647 1095 2648 1099
rect 2642 1094 2648 1095
rect 2644 1068 2646 1094
rect 2642 1067 2648 1068
rect 2642 1063 2643 1067
rect 2647 1063 2648 1067
rect 2642 1062 2648 1063
rect 2724 1052 2726 1113
rect 2730 1099 2736 1100
rect 2730 1095 2731 1099
rect 2735 1095 2736 1099
rect 2730 1094 2736 1095
rect 2732 1060 2734 1094
rect 2730 1059 2736 1060
rect 2730 1055 2731 1059
rect 2735 1055 2736 1059
rect 2730 1054 2736 1055
rect 2892 1052 2894 1113
rect 2898 1099 2904 1100
rect 2898 1095 2899 1099
rect 2903 1095 2904 1099
rect 2898 1094 2904 1095
rect 2900 1060 2902 1094
rect 2898 1059 2904 1060
rect 2898 1055 2899 1059
rect 2903 1055 2904 1059
rect 2898 1054 2904 1055
rect 3060 1052 3062 1113
rect 3066 1099 3072 1100
rect 3066 1095 3067 1099
rect 3071 1095 3072 1099
rect 3066 1094 3072 1095
rect 3068 1060 3070 1094
rect 3066 1059 3072 1060
rect 3066 1055 3067 1059
rect 3071 1055 3072 1059
rect 3066 1054 3072 1055
rect 3220 1052 3222 1113
rect 3226 1099 3232 1100
rect 3226 1095 3227 1099
rect 3231 1095 3232 1099
rect 3226 1094 3232 1095
rect 3228 1060 3230 1094
rect 3236 1060 3238 1138
rect 3332 1119 3334 1196
rect 3372 1184 3374 1362
rect 3396 1316 3398 1377
rect 3402 1363 3408 1364
rect 3402 1359 3403 1363
rect 3407 1359 3408 1363
rect 3402 1358 3408 1359
rect 3404 1324 3406 1358
rect 3402 1323 3408 1324
rect 3402 1319 3403 1323
rect 3407 1319 3408 1323
rect 3402 1318 3408 1319
rect 3652 1316 3654 1377
rect 3658 1363 3664 1364
rect 3658 1359 3659 1363
rect 3663 1359 3664 1363
rect 3658 1358 3664 1359
rect 3660 1324 3662 1358
rect 3780 1324 3782 1386
rect 3800 1383 3802 1451
rect 3840 1407 3842 1471
rect 3860 1407 3862 1472
rect 3986 1467 3992 1468
rect 3986 1463 3987 1467
rect 3991 1463 3992 1467
rect 3986 1462 3992 1463
rect 3988 1428 3990 1462
rect 3954 1427 3960 1428
rect 3954 1423 3955 1427
rect 3959 1423 3960 1427
rect 3954 1422 3960 1423
rect 3986 1427 3992 1428
rect 3986 1423 3987 1427
rect 3991 1423 3992 1427
rect 3986 1422 3992 1423
rect 3839 1406 3843 1407
rect 3839 1401 3843 1402
rect 3859 1406 3863 1407
rect 3859 1401 3863 1402
rect 3799 1382 3803 1383
rect 3799 1377 3803 1378
rect 3658 1323 3664 1324
rect 3658 1319 3659 1323
rect 3663 1319 3664 1323
rect 3658 1318 3664 1319
rect 3778 1323 3784 1324
rect 3778 1319 3779 1323
rect 3783 1319 3784 1323
rect 3778 1318 3784 1319
rect 3800 1317 3802 1377
rect 3840 1341 3842 1401
rect 3838 1340 3844 1341
rect 3860 1340 3862 1401
rect 3956 1348 3958 1422
rect 3996 1407 3998 1472
rect 4122 1467 4128 1468
rect 4122 1463 4123 1467
rect 4127 1463 4128 1467
rect 4122 1462 4128 1463
rect 4124 1428 4126 1462
rect 4122 1427 4128 1428
rect 4122 1423 4123 1427
rect 4127 1423 4128 1427
rect 4122 1422 4128 1423
rect 4132 1407 4134 1472
rect 4252 1468 4254 1610
rect 4356 1568 4358 1629
rect 4398 1619 4404 1620
rect 4398 1615 4399 1619
rect 4403 1615 4404 1619
rect 4398 1614 4404 1615
rect 4354 1567 4360 1568
rect 4354 1563 4355 1567
rect 4359 1563 4360 1567
rect 4354 1562 4360 1563
rect 4382 1552 4388 1553
rect 4382 1548 4383 1552
rect 4387 1548 4388 1552
rect 4382 1547 4388 1548
rect 4384 1523 4386 1547
rect 4303 1522 4307 1523
rect 4303 1517 4307 1518
rect 4383 1522 4387 1523
rect 4383 1517 4387 1518
rect 4258 1507 4264 1508
rect 4258 1503 4259 1507
rect 4263 1503 4264 1507
rect 4258 1502 4264 1503
rect 4250 1467 4256 1468
rect 4250 1463 4251 1467
rect 4255 1463 4256 1467
rect 4250 1462 4256 1463
rect 4154 1459 4160 1460
rect 4154 1455 4155 1459
rect 4159 1455 4160 1459
rect 4154 1454 4160 1455
rect 3995 1406 3999 1407
rect 3995 1401 3999 1402
rect 4059 1406 4063 1407
rect 4059 1401 4063 1402
rect 4131 1406 4135 1407
rect 4131 1401 4135 1402
rect 3954 1347 3960 1348
rect 3954 1343 3955 1347
rect 3959 1343 3960 1347
rect 3954 1342 3960 1343
rect 4060 1340 4062 1401
rect 4156 1392 4158 1454
rect 4260 1428 4262 1502
rect 4304 1493 4306 1517
rect 4302 1492 4308 1493
rect 4302 1488 4303 1492
rect 4307 1488 4308 1492
rect 4302 1487 4308 1488
rect 4274 1477 4280 1478
rect 4274 1473 4275 1477
rect 4279 1473 4280 1477
rect 4274 1472 4280 1473
rect 4258 1427 4264 1428
rect 4258 1423 4259 1427
rect 4263 1423 4264 1427
rect 4258 1422 4264 1423
rect 4276 1407 4278 1472
rect 4400 1468 4402 1614
rect 4478 1575 4484 1576
rect 4478 1571 4479 1575
rect 4483 1571 4484 1575
rect 4478 1570 4484 1571
rect 4466 1477 4472 1478
rect 4466 1473 4467 1477
rect 4471 1473 4472 1477
rect 4466 1472 4472 1473
rect 4398 1467 4404 1468
rect 4398 1463 4399 1467
rect 4403 1463 4404 1467
rect 4398 1462 4404 1463
rect 4468 1407 4470 1472
rect 4480 1428 4482 1570
rect 4588 1568 4590 1629
rect 4682 1615 4688 1616
rect 4682 1611 4683 1615
rect 4687 1611 4688 1615
rect 4682 1610 4688 1611
rect 4684 1584 4686 1610
rect 4682 1583 4688 1584
rect 4682 1579 4683 1583
rect 4687 1579 4688 1583
rect 4682 1578 4688 1579
rect 4852 1568 4854 1629
rect 4872 1620 4874 1686
rect 4996 1635 4998 1696
rect 5088 1652 5090 1810
rect 5108 1808 5110 1869
rect 5244 1808 5246 1869
rect 5250 1855 5256 1856
rect 5250 1851 5251 1855
rect 5255 1851 5256 1855
rect 5250 1850 5256 1851
rect 5252 1816 5254 1850
rect 5250 1815 5256 1816
rect 5250 1811 5251 1815
rect 5255 1811 5256 1815
rect 5250 1810 5256 1811
rect 5380 1808 5382 1869
rect 5498 1815 5504 1816
rect 5498 1811 5499 1815
rect 5503 1811 5504 1815
rect 5498 1810 5504 1811
rect 5106 1807 5112 1808
rect 5106 1803 5107 1807
rect 5111 1803 5112 1807
rect 5106 1802 5112 1803
rect 5242 1807 5248 1808
rect 5242 1803 5243 1807
rect 5247 1803 5248 1807
rect 5242 1802 5248 1803
rect 5378 1807 5384 1808
rect 5378 1803 5379 1807
rect 5383 1803 5384 1807
rect 5378 1802 5384 1803
rect 5134 1792 5140 1793
rect 5134 1788 5135 1792
rect 5139 1788 5140 1792
rect 5134 1787 5140 1788
rect 5270 1792 5276 1793
rect 5270 1788 5271 1792
rect 5275 1788 5276 1792
rect 5270 1787 5276 1788
rect 5406 1792 5412 1793
rect 5406 1788 5407 1792
rect 5411 1788 5412 1792
rect 5406 1787 5412 1788
rect 5136 1747 5138 1787
rect 5272 1747 5274 1787
rect 5408 1747 5410 1787
rect 5135 1746 5139 1747
rect 5135 1741 5139 1742
rect 5271 1746 5275 1747
rect 5271 1741 5275 1742
rect 5279 1746 5283 1747
rect 5279 1741 5283 1742
rect 5407 1746 5411 1747
rect 5407 1741 5411 1742
rect 5280 1717 5282 1741
rect 5278 1716 5284 1717
rect 5278 1712 5279 1716
rect 5283 1712 5284 1716
rect 5278 1711 5284 1712
rect 5250 1701 5256 1702
rect 5250 1697 5251 1701
rect 5255 1697 5256 1701
rect 5250 1696 5256 1697
rect 5086 1651 5092 1652
rect 5086 1647 5087 1651
rect 5091 1647 5092 1651
rect 5086 1646 5092 1647
rect 5252 1635 5254 1696
rect 5500 1652 5502 1810
rect 5516 1808 5518 1869
rect 5612 1860 5614 1938
rect 5640 1904 5642 2162
rect 5664 2111 5666 2171
rect 5663 2110 5667 2111
rect 5663 2105 5667 2106
rect 5664 2045 5666 2105
rect 5662 2044 5668 2045
rect 5662 2040 5663 2044
rect 5667 2040 5668 2044
rect 5662 2039 5668 2040
rect 5662 2027 5668 2028
rect 5662 2023 5663 2027
rect 5667 2023 5668 2027
rect 5662 2022 5668 2023
rect 5664 1999 5666 2022
rect 5663 1998 5667 1999
rect 5663 1993 5667 1994
rect 5664 1970 5666 1993
rect 5662 1969 5668 1970
rect 5662 1965 5663 1969
rect 5667 1965 5668 1969
rect 5662 1964 5668 1965
rect 5662 1952 5668 1953
rect 5662 1948 5663 1952
rect 5667 1948 5668 1952
rect 5662 1947 5668 1948
rect 5638 1903 5644 1904
rect 5638 1899 5639 1903
rect 5643 1899 5644 1903
rect 5638 1898 5644 1899
rect 5664 1875 5666 1947
rect 5663 1874 5667 1875
rect 5663 1869 5667 1870
rect 5610 1859 5616 1860
rect 5610 1855 5611 1859
rect 5615 1855 5616 1859
rect 5610 1854 5616 1855
rect 5664 1809 5666 1869
rect 5662 1808 5668 1809
rect 5514 1807 5520 1808
rect 5514 1803 5515 1807
rect 5519 1803 5520 1807
rect 5662 1804 5663 1808
rect 5667 1804 5668 1808
rect 5662 1803 5668 1804
rect 5514 1802 5520 1803
rect 5542 1792 5548 1793
rect 5542 1788 5543 1792
rect 5547 1788 5548 1792
rect 5542 1787 5548 1788
rect 5662 1791 5668 1792
rect 5662 1787 5663 1791
rect 5667 1787 5668 1791
rect 5544 1747 5546 1787
rect 5662 1786 5668 1787
rect 5664 1747 5666 1786
rect 5535 1746 5539 1747
rect 5535 1741 5539 1742
rect 5543 1746 5547 1747
rect 5543 1741 5547 1742
rect 5663 1746 5667 1747
rect 5663 1741 5667 1742
rect 5536 1717 5538 1741
rect 5664 1718 5666 1741
rect 5662 1717 5668 1718
rect 5534 1716 5540 1717
rect 5534 1712 5535 1716
rect 5539 1712 5540 1716
rect 5662 1713 5663 1717
rect 5667 1713 5668 1717
rect 5662 1712 5668 1713
rect 5534 1711 5540 1712
rect 5506 1701 5512 1702
rect 5506 1697 5507 1701
rect 5511 1697 5512 1701
rect 5506 1696 5512 1697
rect 5662 1700 5668 1701
rect 5662 1696 5663 1700
rect 5667 1696 5668 1700
rect 5346 1651 5352 1652
rect 5346 1647 5347 1651
rect 5351 1647 5352 1651
rect 5346 1646 5352 1647
rect 5498 1651 5504 1652
rect 5498 1647 5499 1651
rect 5503 1647 5504 1651
rect 5498 1646 5504 1647
rect 4995 1634 4999 1635
rect 4995 1629 4999 1630
rect 5131 1634 5135 1635
rect 5131 1629 5135 1630
rect 5251 1634 5255 1635
rect 5251 1629 5255 1630
rect 4870 1619 4876 1620
rect 4870 1615 4871 1619
rect 4875 1615 4876 1619
rect 4870 1614 4876 1615
rect 5132 1568 5134 1629
rect 5138 1615 5144 1616
rect 5138 1611 5139 1615
rect 5143 1611 5144 1615
rect 5138 1610 5144 1611
rect 5140 1576 5142 1610
rect 5348 1576 5350 1646
rect 5508 1635 5510 1696
rect 5662 1695 5668 1696
rect 5554 1691 5560 1692
rect 5554 1687 5555 1691
rect 5559 1687 5560 1691
rect 5554 1686 5560 1687
rect 5419 1634 5423 1635
rect 5419 1629 5423 1630
rect 5507 1634 5511 1635
rect 5507 1629 5511 1630
rect 5138 1575 5144 1576
rect 5138 1571 5139 1575
rect 5143 1571 5144 1575
rect 5138 1570 5144 1571
rect 5346 1575 5352 1576
rect 5346 1571 5347 1575
rect 5351 1571 5352 1575
rect 5346 1570 5352 1571
rect 5420 1568 5422 1629
rect 5466 1619 5472 1620
rect 5466 1615 5467 1619
rect 5471 1615 5472 1619
rect 5466 1614 5472 1615
rect 4586 1567 4592 1568
rect 4586 1563 4587 1567
rect 4591 1563 4592 1567
rect 4586 1562 4592 1563
rect 4850 1567 4856 1568
rect 4850 1563 4851 1567
rect 4855 1563 4856 1567
rect 4850 1562 4856 1563
rect 5130 1567 5136 1568
rect 5130 1563 5131 1567
rect 5135 1563 5136 1567
rect 5130 1562 5136 1563
rect 5418 1567 5424 1568
rect 5418 1563 5419 1567
rect 5423 1563 5424 1567
rect 5418 1562 5424 1563
rect 4614 1552 4620 1553
rect 4614 1548 4615 1552
rect 4619 1548 4620 1552
rect 4614 1547 4620 1548
rect 4878 1552 4884 1553
rect 4878 1548 4879 1552
rect 4883 1548 4884 1552
rect 4878 1547 4884 1548
rect 5158 1552 5164 1553
rect 5158 1548 5159 1552
rect 5163 1548 5164 1552
rect 5158 1547 5164 1548
rect 5446 1552 5452 1553
rect 5446 1548 5447 1552
rect 5451 1548 5452 1552
rect 5446 1547 5452 1548
rect 4616 1523 4618 1547
rect 4880 1523 4882 1547
rect 5160 1523 5162 1547
rect 5448 1523 5450 1547
rect 4495 1522 4499 1523
rect 4495 1517 4499 1518
rect 4615 1522 4619 1523
rect 4615 1517 4619 1518
rect 4719 1522 4723 1523
rect 4719 1517 4723 1518
rect 4879 1522 4883 1523
rect 4879 1517 4883 1518
rect 4967 1522 4971 1523
rect 4967 1517 4971 1518
rect 5159 1522 5163 1523
rect 5159 1517 5163 1518
rect 5223 1522 5227 1523
rect 5223 1517 5227 1518
rect 5447 1522 5451 1523
rect 5447 1517 5451 1518
rect 4496 1493 4498 1517
rect 4720 1493 4722 1517
rect 4968 1493 4970 1517
rect 5224 1493 5226 1517
rect 4494 1492 4500 1493
rect 4494 1488 4495 1492
rect 4499 1488 4500 1492
rect 4494 1487 4500 1488
rect 4718 1492 4724 1493
rect 4718 1488 4719 1492
rect 4723 1488 4724 1492
rect 4718 1487 4724 1488
rect 4966 1492 4972 1493
rect 4966 1488 4967 1492
rect 4971 1488 4972 1492
rect 4966 1487 4972 1488
rect 5222 1492 5228 1493
rect 5222 1488 5223 1492
rect 5227 1488 5228 1492
rect 5222 1487 5228 1488
rect 4690 1477 4696 1478
rect 4690 1473 4691 1477
rect 4695 1473 4696 1477
rect 4690 1472 4696 1473
rect 4938 1477 4944 1478
rect 4938 1473 4939 1477
rect 4943 1473 4944 1477
rect 4938 1472 4944 1473
rect 5194 1477 5200 1478
rect 5194 1473 5195 1477
rect 5199 1473 5200 1477
rect 5194 1472 5200 1473
rect 5458 1477 5464 1478
rect 5458 1473 5459 1477
rect 5463 1473 5464 1477
rect 5458 1472 5464 1473
rect 4594 1467 4600 1468
rect 4594 1463 4595 1467
rect 4599 1463 4600 1467
rect 4594 1462 4600 1463
rect 4596 1428 4598 1462
rect 4478 1427 4484 1428
rect 4478 1423 4479 1427
rect 4483 1423 4484 1427
rect 4478 1422 4484 1423
rect 4594 1427 4600 1428
rect 4594 1423 4595 1427
rect 4599 1423 4600 1427
rect 4594 1422 4600 1423
rect 4692 1407 4694 1472
rect 4818 1467 4824 1468
rect 4818 1463 4819 1467
rect 4823 1463 4824 1467
rect 4818 1462 4824 1463
rect 4820 1428 4822 1462
rect 4818 1427 4824 1428
rect 4818 1423 4819 1427
rect 4823 1423 4824 1427
rect 4818 1422 4824 1423
rect 4940 1407 4942 1472
rect 5066 1467 5072 1468
rect 5066 1463 5067 1467
rect 5071 1463 5072 1467
rect 5066 1462 5072 1463
rect 5068 1428 5070 1462
rect 5066 1427 5072 1428
rect 5066 1423 5067 1427
rect 5071 1423 5072 1427
rect 5066 1422 5072 1423
rect 5196 1407 5198 1472
rect 5460 1407 5462 1472
rect 4275 1406 4279 1407
rect 4275 1401 4279 1402
rect 4307 1406 4311 1407
rect 4307 1401 4311 1402
rect 4467 1406 4471 1407
rect 4467 1401 4471 1402
rect 4579 1406 4583 1407
rect 4579 1401 4583 1402
rect 4691 1406 4695 1407
rect 4691 1401 4695 1402
rect 4875 1406 4879 1407
rect 4875 1401 4879 1402
rect 4939 1406 4943 1407
rect 4939 1401 4943 1402
rect 5187 1406 5191 1407
rect 5187 1401 5191 1402
rect 5195 1406 5199 1407
rect 5195 1401 5199 1402
rect 5459 1406 5463 1407
rect 5459 1401 5463 1402
rect 4154 1391 4160 1392
rect 4154 1387 4155 1391
rect 4159 1387 4160 1391
rect 4154 1386 4160 1387
rect 4308 1340 4310 1401
rect 4314 1387 4320 1388
rect 4314 1383 4315 1387
rect 4319 1383 4320 1387
rect 4314 1382 4320 1383
rect 4316 1348 4318 1382
rect 4314 1347 4320 1348
rect 4314 1343 4315 1347
rect 4319 1343 4320 1347
rect 4314 1342 4320 1343
rect 4580 1340 4582 1401
rect 4586 1387 4592 1388
rect 4586 1383 4587 1387
rect 4591 1383 4592 1387
rect 4586 1382 4592 1383
rect 4588 1348 4590 1382
rect 4682 1355 4688 1356
rect 4682 1351 4683 1355
rect 4687 1351 4688 1355
rect 4682 1350 4688 1351
rect 4586 1347 4592 1348
rect 4586 1343 4587 1347
rect 4591 1343 4592 1347
rect 4586 1342 4592 1343
rect 3838 1336 3839 1340
rect 3843 1336 3844 1340
rect 3838 1335 3844 1336
rect 3858 1339 3864 1340
rect 3858 1335 3859 1339
rect 3863 1335 3864 1339
rect 3858 1334 3864 1335
rect 4058 1339 4064 1340
rect 4058 1335 4059 1339
rect 4063 1335 4064 1339
rect 4058 1334 4064 1335
rect 4306 1339 4312 1340
rect 4306 1335 4307 1339
rect 4311 1335 4312 1339
rect 4306 1334 4312 1335
rect 4578 1339 4584 1340
rect 4578 1335 4579 1339
rect 4583 1335 4584 1339
rect 4578 1334 4584 1335
rect 3886 1324 3892 1325
rect 3838 1323 3844 1324
rect 3838 1319 3839 1323
rect 3843 1319 3844 1323
rect 3886 1320 3887 1324
rect 3891 1320 3892 1324
rect 3886 1319 3892 1320
rect 4086 1324 4092 1325
rect 4086 1320 4087 1324
rect 4091 1320 4092 1324
rect 4086 1319 4092 1320
rect 4334 1324 4340 1325
rect 4334 1320 4335 1324
rect 4339 1320 4340 1324
rect 4334 1319 4340 1320
rect 4606 1324 4612 1325
rect 4606 1320 4607 1324
rect 4611 1320 4612 1324
rect 4606 1319 4612 1320
rect 3838 1318 3844 1319
rect 3798 1316 3804 1317
rect 3394 1315 3400 1316
rect 3394 1311 3395 1315
rect 3399 1311 3400 1315
rect 3394 1310 3400 1311
rect 3650 1315 3656 1316
rect 3650 1311 3651 1315
rect 3655 1311 3656 1315
rect 3798 1312 3799 1316
rect 3803 1312 3804 1316
rect 3798 1311 3804 1312
rect 3650 1310 3656 1311
rect 3422 1300 3428 1301
rect 3422 1296 3423 1300
rect 3427 1296 3428 1300
rect 3422 1295 3428 1296
rect 3678 1300 3684 1301
rect 3678 1296 3679 1300
rect 3683 1296 3684 1300
rect 3678 1295 3684 1296
rect 3798 1299 3804 1300
rect 3798 1295 3799 1299
rect 3803 1295 3804 1299
rect 3424 1247 3426 1295
rect 3680 1247 3682 1295
rect 3798 1294 3804 1295
rect 3800 1247 3802 1294
rect 3840 1287 3842 1318
rect 3888 1287 3890 1319
rect 4088 1287 4090 1319
rect 4336 1287 4338 1319
rect 4608 1287 4610 1319
rect 3839 1286 3843 1287
rect 3839 1281 3843 1282
rect 3887 1286 3891 1287
rect 3887 1281 3891 1282
rect 4087 1286 4091 1287
rect 4087 1281 4091 1282
rect 4335 1286 4339 1287
rect 4335 1281 4339 1282
rect 4607 1286 4611 1287
rect 4607 1281 4611 1282
rect 4615 1286 4619 1287
rect 4615 1281 4619 1282
rect 3840 1258 3842 1281
rect 3838 1257 3844 1258
rect 4616 1257 4618 1281
rect 3838 1253 3839 1257
rect 3843 1253 3844 1257
rect 3838 1252 3844 1253
rect 4614 1256 4620 1257
rect 4614 1252 4615 1256
rect 4619 1252 4620 1256
rect 4614 1251 4620 1252
rect 3423 1246 3427 1247
rect 3423 1241 3427 1242
rect 3543 1246 3547 1247
rect 3543 1241 3547 1242
rect 3679 1246 3683 1247
rect 3679 1241 3683 1242
rect 3799 1246 3803 1247
rect 3799 1241 3803 1242
rect 4586 1241 4592 1242
rect 3544 1217 3546 1241
rect 3800 1218 3802 1241
rect 3838 1240 3844 1241
rect 3838 1236 3839 1240
rect 3843 1236 3844 1240
rect 4586 1237 4587 1241
rect 4591 1237 4592 1241
rect 4586 1236 4592 1237
rect 3838 1235 3844 1236
rect 3798 1217 3804 1218
rect 3542 1216 3548 1217
rect 3542 1212 3543 1216
rect 3547 1212 3548 1216
rect 3798 1213 3799 1217
rect 3803 1213 3804 1217
rect 3798 1212 3804 1213
rect 3542 1211 3548 1212
rect 3514 1201 3520 1202
rect 3514 1197 3515 1201
rect 3519 1197 3520 1201
rect 3514 1196 3520 1197
rect 3798 1200 3804 1201
rect 3798 1196 3799 1200
rect 3803 1196 3804 1200
rect 3458 1191 3464 1192
rect 3458 1187 3459 1191
rect 3463 1187 3464 1191
rect 3458 1186 3464 1187
rect 3370 1183 3376 1184
rect 3370 1179 3371 1183
rect 3375 1179 3376 1183
rect 3370 1178 3376 1179
rect 3460 1152 3462 1186
rect 3458 1151 3464 1152
rect 3458 1147 3459 1151
rect 3463 1147 3464 1151
rect 3458 1146 3464 1147
rect 3516 1119 3518 1196
rect 3798 1195 3804 1196
rect 3800 1119 3802 1195
rect 3840 1171 3842 1235
rect 4588 1171 4590 1236
rect 4684 1192 4686 1350
rect 4876 1340 4878 1401
rect 4882 1387 4888 1388
rect 4882 1383 4883 1387
rect 4887 1383 4888 1387
rect 4882 1382 4888 1383
rect 4884 1348 4886 1382
rect 4882 1347 4888 1348
rect 4882 1343 4883 1347
rect 4887 1343 4888 1347
rect 4882 1342 4888 1343
rect 5188 1340 5190 1401
rect 5194 1387 5200 1388
rect 5194 1383 5195 1387
rect 5199 1383 5200 1387
rect 5194 1382 5200 1383
rect 5196 1348 5198 1382
rect 5194 1347 5200 1348
rect 5194 1343 5195 1347
rect 5199 1343 5200 1347
rect 5194 1342 5200 1343
rect 4874 1339 4880 1340
rect 4874 1335 4875 1339
rect 4879 1335 4880 1339
rect 4874 1334 4880 1335
rect 5186 1339 5192 1340
rect 5186 1335 5187 1339
rect 5191 1335 5192 1339
rect 5186 1334 5192 1335
rect 4902 1324 4908 1325
rect 4902 1320 4903 1324
rect 4907 1320 4908 1324
rect 4902 1319 4908 1320
rect 5214 1324 5220 1325
rect 5214 1320 5215 1324
rect 5219 1320 5220 1324
rect 5214 1319 5220 1320
rect 4904 1287 4906 1319
rect 5216 1287 5218 1319
rect 4791 1286 4795 1287
rect 4791 1281 4795 1282
rect 4903 1286 4907 1287
rect 4903 1281 4907 1282
rect 4975 1286 4979 1287
rect 4975 1281 4979 1282
rect 5167 1286 5171 1287
rect 5167 1281 5171 1282
rect 5215 1286 5219 1287
rect 5215 1281 5219 1282
rect 5367 1286 5371 1287
rect 5367 1281 5371 1282
rect 4792 1257 4794 1281
rect 4976 1257 4978 1281
rect 5168 1257 5170 1281
rect 5368 1257 5370 1281
rect 4790 1256 4796 1257
rect 4790 1252 4791 1256
rect 4795 1252 4796 1256
rect 4790 1251 4796 1252
rect 4974 1256 4980 1257
rect 4974 1252 4975 1256
rect 4979 1252 4980 1256
rect 4974 1251 4980 1252
rect 5166 1256 5172 1257
rect 5166 1252 5167 1256
rect 5171 1252 5172 1256
rect 5166 1251 5172 1252
rect 5366 1256 5372 1257
rect 5366 1252 5367 1256
rect 5371 1252 5372 1256
rect 5366 1251 5372 1252
rect 4762 1241 4768 1242
rect 4762 1237 4763 1241
rect 4767 1237 4768 1241
rect 4762 1236 4768 1237
rect 4946 1241 4952 1242
rect 4946 1237 4947 1241
rect 4951 1237 4952 1241
rect 4946 1236 4952 1237
rect 5138 1241 5144 1242
rect 5138 1237 5139 1241
rect 5143 1237 5144 1241
rect 5138 1236 5144 1237
rect 5338 1241 5344 1242
rect 5338 1237 5339 1241
rect 5343 1237 5344 1241
rect 5338 1236 5344 1237
rect 4714 1231 4720 1232
rect 4714 1227 4715 1231
rect 4719 1227 4720 1231
rect 4714 1226 4720 1227
rect 4716 1192 4718 1226
rect 4682 1191 4688 1192
rect 4682 1187 4683 1191
rect 4687 1187 4688 1191
rect 4682 1186 4688 1187
rect 4714 1191 4720 1192
rect 4714 1187 4715 1191
rect 4719 1187 4720 1191
rect 4714 1186 4720 1187
rect 4764 1171 4766 1236
rect 4890 1231 4896 1232
rect 4890 1227 4891 1231
rect 4895 1227 4896 1231
rect 4890 1226 4896 1227
rect 4892 1192 4894 1226
rect 4890 1191 4896 1192
rect 4890 1187 4891 1191
rect 4895 1187 4896 1191
rect 4890 1186 4896 1187
rect 4948 1171 4950 1236
rect 5074 1231 5080 1232
rect 5074 1227 5075 1231
rect 5079 1227 5080 1231
rect 5074 1226 5080 1227
rect 5082 1231 5088 1232
rect 5082 1227 5083 1231
rect 5087 1227 5088 1231
rect 5082 1226 5088 1227
rect 5076 1192 5078 1226
rect 5074 1191 5080 1192
rect 5074 1187 5075 1191
rect 5079 1187 5080 1191
rect 5074 1186 5080 1187
rect 3839 1170 3843 1171
rect 3839 1165 3843 1166
rect 4587 1170 4591 1171
rect 4587 1165 4591 1166
rect 4763 1170 4767 1171
rect 4763 1165 4767 1166
rect 4835 1170 4839 1171
rect 4835 1165 4839 1166
rect 4947 1170 4951 1171
rect 4947 1165 4951 1166
rect 4971 1170 4975 1171
rect 4971 1165 4975 1166
rect 3331 1118 3335 1119
rect 3331 1113 3335 1114
rect 3387 1118 3391 1119
rect 3387 1113 3391 1114
rect 3515 1118 3519 1119
rect 3515 1113 3519 1114
rect 3799 1118 3803 1119
rect 3799 1113 3803 1114
rect 3226 1059 3232 1060
rect 3226 1055 3227 1059
rect 3231 1055 3232 1059
rect 3226 1054 3232 1055
rect 3234 1059 3240 1060
rect 3234 1055 3235 1059
rect 3239 1055 3240 1059
rect 3234 1054 3240 1055
rect 3388 1052 3390 1113
rect 3406 1103 3412 1104
rect 3406 1099 3407 1103
rect 3411 1099 3412 1103
rect 3406 1098 3412 1099
rect 2546 1051 2552 1052
rect 2546 1047 2547 1051
rect 2551 1047 2552 1051
rect 2546 1046 2552 1047
rect 2722 1051 2728 1052
rect 2722 1047 2723 1051
rect 2727 1047 2728 1051
rect 2722 1046 2728 1047
rect 2890 1051 2896 1052
rect 2890 1047 2891 1051
rect 2895 1047 2896 1051
rect 2890 1046 2896 1047
rect 3058 1051 3064 1052
rect 3058 1047 3059 1051
rect 3063 1047 3064 1051
rect 3058 1046 3064 1047
rect 3218 1051 3224 1052
rect 3218 1047 3219 1051
rect 3223 1047 3224 1051
rect 3218 1046 3224 1047
rect 3386 1051 3392 1052
rect 3386 1047 3387 1051
rect 3391 1047 3392 1051
rect 3386 1046 3392 1047
rect 2574 1036 2580 1037
rect 2574 1032 2575 1036
rect 2579 1032 2580 1036
rect 2574 1031 2580 1032
rect 2750 1036 2756 1037
rect 2750 1032 2751 1036
rect 2755 1032 2756 1036
rect 2750 1031 2756 1032
rect 2918 1036 2924 1037
rect 2918 1032 2919 1036
rect 2923 1032 2924 1036
rect 2918 1031 2924 1032
rect 3086 1036 3092 1037
rect 3086 1032 3087 1036
rect 3091 1032 3092 1036
rect 3086 1031 3092 1032
rect 3246 1036 3252 1037
rect 3246 1032 3247 1036
rect 3251 1032 3252 1036
rect 3246 1031 3252 1032
rect 2576 1007 2578 1031
rect 2752 1007 2754 1031
rect 2920 1007 2922 1031
rect 3088 1007 3090 1031
rect 3248 1007 3250 1031
rect 2567 1006 2571 1007
rect 2567 1001 2571 1002
rect 2575 1006 2579 1007
rect 2575 1001 2579 1002
rect 2751 1006 2755 1007
rect 2751 1001 2755 1002
rect 2759 1006 2763 1007
rect 2759 1001 2763 1002
rect 2919 1006 2923 1007
rect 2919 1001 2923 1002
rect 2943 1006 2947 1007
rect 2943 1001 2947 1002
rect 3087 1006 3091 1007
rect 3087 1001 3091 1002
rect 3127 1006 3131 1007
rect 3127 1001 3131 1002
rect 3247 1006 3251 1007
rect 3247 1001 3251 1002
rect 3311 1006 3315 1007
rect 3311 1001 3315 1002
rect 2568 977 2570 1001
rect 2760 977 2762 1001
rect 2944 977 2946 1001
rect 3128 977 3130 1001
rect 3312 977 3314 1001
rect 2566 976 2572 977
rect 2566 972 2567 976
rect 2571 972 2572 976
rect 2566 971 2572 972
rect 2758 976 2764 977
rect 2758 972 2759 976
rect 2763 972 2764 976
rect 2758 971 2764 972
rect 2942 976 2948 977
rect 2942 972 2943 976
rect 2947 972 2948 976
rect 2942 971 2948 972
rect 3126 976 3132 977
rect 3126 972 3127 976
rect 3131 972 3132 976
rect 3126 971 3132 972
rect 3310 976 3316 977
rect 3310 972 3311 976
rect 3315 972 3316 976
rect 3310 971 3316 972
rect 2538 961 2544 962
rect 2538 957 2539 961
rect 2543 957 2544 961
rect 2538 956 2544 957
rect 2730 961 2736 962
rect 2730 957 2731 961
rect 2735 957 2736 961
rect 2730 956 2736 957
rect 2914 961 2920 962
rect 2914 957 2915 961
rect 2919 957 2920 961
rect 2914 956 2920 957
rect 3098 961 3104 962
rect 3098 957 3099 961
rect 3103 957 3104 961
rect 3098 956 3104 957
rect 3282 961 3288 962
rect 3282 957 3283 961
rect 3287 957 3288 961
rect 3282 956 3288 957
rect 2490 911 2496 912
rect 2490 907 2491 911
rect 2495 907 2496 911
rect 2490 906 2496 907
rect 2540 891 2542 956
rect 2666 951 2672 952
rect 2666 947 2667 951
rect 2671 947 2672 951
rect 2666 946 2672 947
rect 2668 912 2670 946
rect 2666 911 2672 912
rect 2666 907 2667 911
rect 2671 907 2672 911
rect 2666 906 2672 907
rect 2732 891 2734 956
rect 2894 951 2900 952
rect 2894 947 2895 951
rect 2899 947 2900 951
rect 2894 946 2900 947
rect 1975 890 1979 891
rect 1975 885 1979 886
rect 1995 890 1999 891
rect 1995 885 1999 886
rect 2163 890 2167 891
rect 2163 885 2167 886
rect 2179 890 2183 891
rect 2179 885 2183 886
rect 2347 890 2351 891
rect 2347 885 2351 886
rect 2403 890 2407 891
rect 2403 885 2407 886
rect 2539 890 2543 891
rect 2539 885 2543 886
rect 2675 890 2679 891
rect 2675 885 2679 886
rect 2731 890 2735 891
rect 2731 885 2735 886
rect 1934 884 1940 885
rect 1934 880 1935 884
rect 1939 880 1940 884
rect 1934 879 1940 880
rect 1934 867 1940 868
rect 1934 863 1935 867
rect 1939 863 1940 867
rect 1934 862 1940 863
rect 1936 823 1938 862
rect 1976 825 1978 885
rect 1974 824 1980 825
rect 1996 824 1998 885
rect 2180 824 2182 885
rect 2186 871 2192 872
rect 2186 867 2187 871
rect 2191 867 2192 871
rect 2186 866 2192 867
rect 2188 832 2190 866
rect 2186 831 2192 832
rect 2186 827 2187 831
rect 2191 827 2192 831
rect 2186 826 2192 827
rect 2404 824 2406 885
rect 2526 883 2532 884
rect 2526 879 2527 883
rect 2531 879 2532 883
rect 2526 878 2532 879
rect 2528 832 2530 878
rect 2526 831 2532 832
rect 2526 827 2527 831
rect 2531 827 2532 831
rect 2526 826 2532 827
rect 2676 824 2678 885
rect 2896 876 2898 946
rect 2916 891 2918 956
rect 3042 951 3048 952
rect 3042 947 3043 951
rect 3047 947 3048 951
rect 3042 946 3048 947
rect 3010 943 3016 944
rect 3010 939 3011 943
rect 3015 939 3016 943
rect 3010 938 3016 939
rect 3012 912 3014 938
rect 3044 912 3046 946
rect 3010 911 3016 912
rect 3010 907 3011 911
rect 3015 907 3016 911
rect 3010 906 3016 907
rect 3042 911 3048 912
rect 3042 907 3043 911
rect 3047 907 3048 911
rect 3042 906 3048 907
rect 3100 891 3102 956
rect 3226 951 3232 952
rect 3226 947 3227 951
rect 3231 947 3232 951
rect 3226 946 3232 947
rect 3228 912 3230 946
rect 3226 911 3232 912
rect 3226 907 3227 911
rect 3231 907 3232 911
rect 3226 906 3232 907
rect 3284 891 3286 956
rect 3408 952 3410 1098
rect 3800 1053 3802 1113
rect 3840 1105 3842 1165
rect 3838 1104 3844 1105
rect 4836 1104 4838 1165
rect 4972 1104 4974 1165
rect 5084 1160 5086 1226
rect 5140 1171 5142 1236
rect 5340 1171 5342 1236
rect 5468 1232 5470 1614
rect 5487 1522 5491 1523
rect 5487 1517 5491 1518
rect 5488 1493 5490 1517
rect 5486 1492 5492 1493
rect 5486 1488 5487 1492
rect 5491 1488 5492 1492
rect 5486 1487 5492 1488
rect 5556 1428 5558 1686
rect 5664 1635 5666 1695
rect 5663 1634 5667 1635
rect 5663 1629 5667 1630
rect 5664 1569 5666 1629
rect 5662 1568 5668 1569
rect 5662 1564 5663 1568
rect 5667 1564 5668 1568
rect 5662 1563 5668 1564
rect 5662 1551 5668 1552
rect 5662 1547 5663 1551
rect 5667 1547 5668 1551
rect 5662 1546 5668 1547
rect 5664 1523 5666 1546
rect 5663 1522 5667 1523
rect 5663 1517 5667 1518
rect 5664 1494 5666 1517
rect 5662 1493 5668 1494
rect 5662 1489 5663 1493
rect 5667 1489 5668 1493
rect 5662 1488 5668 1489
rect 5662 1476 5668 1477
rect 5662 1472 5663 1476
rect 5667 1472 5668 1476
rect 5662 1471 5668 1472
rect 5582 1467 5588 1468
rect 5582 1463 5583 1467
rect 5587 1463 5588 1467
rect 5582 1462 5588 1463
rect 5554 1427 5560 1428
rect 5554 1423 5555 1427
rect 5559 1423 5560 1427
rect 5554 1422 5560 1423
rect 5499 1406 5503 1407
rect 5499 1401 5503 1402
rect 5500 1340 5502 1401
rect 5584 1392 5586 1462
rect 5664 1407 5666 1471
rect 5663 1406 5667 1407
rect 5663 1401 5667 1402
rect 5582 1391 5588 1392
rect 5582 1387 5583 1391
rect 5587 1387 5588 1391
rect 5582 1386 5588 1387
rect 5610 1347 5616 1348
rect 5610 1343 5611 1347
rect 5615 1343 5616 1347
rect 5610 1342 5616 1343
rect 5498 1339 5504 1340
rect 5498 1335 5499 1339
rect 5503 1335 5504 1339
rect 5498 1334 5504 1335
rect 5526 1324 5532 1325
rect 5526 1320 5527 1324
rect 5531 1320 5532 1324
rect 5526 1319 5532 1320
rect 5528 1287 5530 1319
rect 5527 1286 5531 1287
rect 5527 1281 5531 1282
rect 5543 1286 5547 1287
rect 5543 1281 5547 1282
rect 5544 1257 5546 1281
rect 5542 1256 5548 1257
rect 5542 1252 5543 1256
rect 5547 1252 5548 1256
rect 5542 1251 5548 1252
rect 5514 1241 5520 1242
rect 5514 1237 5515 1241
rect 5519 1237 5520 1241
rect 5514 1236 5520 1237
rect 5466 1231 5472 1232
rect 5466 1227 5467 1231
rect 5471 1227 5472 1231
rect 5466 1226 5472 1227
rect 5478 1191 5484 1192
rect 5478 1187 5479 1191
rect 5483 1187 5484 1191
rect 5478 1186 5484 1187
rect 5107 1170 5111 1171
rect 5107 1165 5111 1166
rect 5139 1170 5143 1171
rect 5139 1165 5143 1166
rect 5243 1170 5247 1171
rect 5243 1165 5247 1166
rect 5339 1170 5343 1171
rect 5339 1165 5343 1166
rect 5379 1170 5383 1171
rect 5379 1165 5383 1166
rect 5082 1159 5088 1160
rect 5082 1155 5083 1159
rect 5087 1155 5088 1159
rect 5082 1154 5088 1155
rect 4978 1151 4984 1152
rect 4978 1147 4979 1151
rect 4983 1147 4984 1151
rect 4978 1146 4984 1147
rect 4980 1112 4982 1146
rect 4978 1111 4984 1112
rect 4978 1107 4979 1111
rect 4983 1107 4984 1111
rect 4978 1106 4984 1107
rect 5108 1104 5110 1165
rect 5114 1151 5120 1152
rect 5114 1147 5115 1151
rect 5119 1147 5120 1151
rect 5114 1146 5120 1147
rect 5116 1112 5118 1146
rect 5114 1111 5120 1112
rect 5114 1107 5115 1111
rect 5119 1107 5120 1111
rect 5114 1106 5120 1107
rect 5244 1104 5246 1165
rect 5250 1151 5256 1152
rect 5250 1147 5251 1151
rect 5255 1147 5256 1151
rect 5250 1146 5256 1147
rect 5252 1112 5254 1146
rect 5250 1111 5256 1112
rect 5250 1107 5251 1111
rect 5255 1107 5256 1111
rect 5250 1106 5256 1107
rect 5380 1104 5382 1165
rect 5386 1151 5392 1152
rect 5386 1147 5387 1151
rect 5391 1147 5392 1151
rect 5386 1146 5392 1147
rect 5388 1112 5390 1146
rect 5386 1111 5392 1112
rect 5386 1107 5387 1111
rect 5391 1107 5392 1111
rect 5386 1106 5392 1107
rect 5418 1111 5424 1112
rect 5418 1107 5419 1111
rect 5423 1107 5424 1111
rect 5418 1106 5424 1107
rect 3838 1100 3839 1104
rect 3843 1100 3844 1104
rect 3838 1099 3844 1100
rect 4834 1103 4840 1104
rect 4834 1099 4835 1103
rect 4839 1099 4840 1103
rect 4834 1098 4840 1099
rect 4970 1103 4976 1104
rect 4970 1099 4971 1103
rect 4975 1099 4976 1103
rect 4970 1098 4976 1099
rect 5106 1103 5112 1104
rect 5106 1099 5107 1103
rect 5111 1099 5112 1103
rect 5106 1098 5112 1099
rect 5242 1103 5248 1104
rect 5242 1099 5243 1103
rect 5247 1099 5248 1103
rect 5242 1098 5248 1099
rect 5378 1103 5384 1104
rect 5378 1099 5379 1103
rect 5383 1099 5384 1103
rect 5378 1098 5384 1099
rect 4862 1088 4868 1089
rect 3838 1087 3844 1088
rect 3838 1083 3839 1087
rect 3843 1083 3844 1087
rect 4862 1084 4863 1088
rect 4867 1084 4868 1088
rect 4862 1083 4868 1084
rect 4998 1088 5004 1089
rect 4998 1084 4999 1088
rect 5003 1084 5004 1088
rect 4998 1083 5004 1084
rect 5134 1088 5140 1089
rect 5134 1084 5135 1088
rect 5139 1084 5140 1088
rect 5134 1083 5140 1084
rect 5270 1088 5276 1089
rect 5270 1084 5271 1088
rect 5275 1084 5276 1088
rect 5270 1083 5276 1084
rect 5406 1088 5412 1089
rect 5406 1084 5407 1088
rect 5411 1084 5412 1088
rect 5406 1083 5412 1084
rect 3838 1082 3844 1083
rect 3840 1055 3842 1082
rect 4864 1055 4866 1083
rect 5000 1055 5002 1083
rect 5136 1055 5138 1083
rect 5272 1055 5274 1083
rect 5408 1055 5410 1083
rect 3839 1054 3843 1055
rect 3798 1052 3804 1053
rect 3798 1048 3799 1052
rect 3803 1048 3804 1052
rect 3839 1049 3843 1050
rect 4807 1054 4811 1055
rect 4807 1049 4811 1050
rect 4863 1054 4867 1055
rect 4863 1049 4867 1050
rect 4943 1054 4947 1055
rect 4943 1049 4947 1050
rect 4999 1054 5003 1055
rect 4999 1049 5003 1050
rect 5079 1054 5083 1055
rect 5079 1049 5083 1050
rect 5135 1054 5139 1055
rect 5135 1049 5139 1050
rect 5215 1054 5219 1055
rect 5215 1049 5219 1050
rect 5271 1054 5275 1055
rect 5271 1049 5275 1050
rect 5351 1054 5355 1055
rect 5351 1049 5355 1050
rect 5407 1054 5411 1055
rect 5407 1049 5411 1050
rect 3798 1047 3804 1048
rect 3414 1036 3420 1037
rect 3414 1032 3415 1036
rect 3419 1032 3420 1036
rect 3414 1031 3420 1032
rect 3798 1035 3804 1036
rect 3798 1031 3799 1035
rect 3803 1031 3804 1035
rect 3416 1007 3418 1031
rect 3798 1030 3804 1031
rect 3800 1007 3802 1030
rect 3840 1026 3842 1049
rect 3838 1025 3844 1026
rect 4808 1025 4810 1049
rect 4944 1025 4946 1049
rect 5080 1025 5082 1049
rect 5216 1025 5218 1049
rect 5352 1025 5354 1049
rect 3838 1021 3839 1025
rect 3843 1021 3844 1025
rect 3838 1020 3844 1021
rect 4806 1024 4812 1025
rect 4806 1020 4807 1024
rect 4811 1020 4812 1024
rect 4806 1019 4812 1020
rect 4942 1024 4948 1025
rect 4942 1020 4943 1024
rect 4947 1020 4948 1024
rect 4942 1019 4948 1020
rect 5078 1024 5084 1025
rect 5078 1020 5079 1024
rect 5083 1020 5084 1024
rect 5078 1019 5084 1020
rect 5214 1024 5220 1025
rect 5214 1020 5215 1024
rect 5219 1020 5220 1024
rect 5214 1019 5220 1020
rect 5350 1024 5356 1025
rect 5350 1020 5351 1024
rect 5355 1020 5356 1024
rect 5350 1019 5356 1020
rect 4778 1009 4784 1010
rect 3838 1008 3844 1009
rect 3415 1006 3419 1007
rect 3415 1001 3419 1002
rect 3495 1006 3499 1007
rect 3495 1001 3499 1002
rect 3679 1006 3683 1007
rect 3679 1001 3683 1002
rect 3799 1006 3803 1007
rect 3838 1004 3839 1008
rect 3843 1004 3844 1008
rect 4778 1005 4779 1009
rect 4783 1005 4784 1009
rect 4778 1004 4784 1005
rect 4914 1009 4920 1010
rect 4914 1005 4915 1009
rect 4919 1005 4920 1009
rect 4914 1004 4920 1005
rect 5050 1009 5056 1010
rect 5050 1005 5051 1009
rect 5055 1005 5056 1009
rect 5050 1004 5056 1005
rect 5186 1009 5192 1010
rect 5186 1005 5187 1009
rect 5191 1005 5192 1009
rect 5186 1004 5192 1005
rect 5322 1009 5328 1010
rect 5322 1005 5323 1009
rect 5327 1005 5328 1009
rect 5322 1004 5328 1005
rect 3838 1003 3844 1004
rect 3799 1001 3803 1002
rect 3496 977 3498 1001
rect 3680 977 3682 1001
rect 3800 978 3802 1001
rect 3798 977 3804 978
rect 3494 976 3500 977
rect 3494 972 3495 976
rect 3499 972 3500 976
rect 3494 971 3500 972
rect 3678 976 3684 977
rect 3678 972 3679 976
rect 3683 972 3684 976
rect 3798 973 3799 977
rect 3803 973 3804 977
rect 3798 972 3804 973
rect 3678 971 3684 972
rect 3466 961 3472 962
rect 3466 957 3467 961
rect 3471 957 3472 961
rect 3466 956 3472 957
rect 3650 961 3656 962
rect 3650 957 3651 961
rect 3655 957 3656 961
rect 3650 956 3656 957
rect 3798 960 3804 961
rect 3798 956 3799 960
rect 3803 956 3804 960
rect 3406 951 3412 952
rect 3406 947 3407 951
rect 3411 947 3412 951
rect 3406 946 3412 947
rect 3468 891 3470 956
rect 3642 951 3648 952
rect 3642 947 3643 951
rect 3647 947 3648 951
rect 3642 946 3648 947
rect 3644 912 3646 946
rect 3642 911 3648 912
rect 3642 907 3643 911
rect 3647 907 3648 911
rect 3642 906 3648 907
rect 3652 891 3654 956
rect 3798 955 3804 956
rect 3746 911 3752 912
rect 3746 907 3747 911
rect 3751 907 3752 911
rect 3746 906 3752 907
rect 2915 890 2919 891
rect 2915 885 2919 886
rect 2987 890 2991 891
rect 2987 885 2991 886
rect 3099 890 3103 891
rect 3099 885 3103 886
rect 3283 890 3287 891
rect 3283 885 3287 886
rect 3323 890 3327 891
rect 3323 885 3327 886
rect 3467 890 3471 891
rect 3467 885 3471 886
rect 3651 890 3655 891
rect 3651 885 3655 886
rect 2894 875 2900 876
rect 2770 871 2776 872
rect 2770 867 2771 871
rect 2775 867 2776 871
rect 2894 871 2895 875
rect 2899 871 2900 875
rect 2894 870 2900 871
rect 2770 866 2776 867
rect 2772 840 2774 866
rect 2770 839 2776 840
rect 2770 835 2771 839
rect 2775 835 2776 839
rect 2770 834 2776 835
rect 2988 824 2990 885
rect 3324 824 3326 885
rect 3330 871 3336 872
rect 3330 867 3331 871
rect 3335 867 3336 871
rect 3330 866 3336 867
rect 3332 832 3334 866
rect 3330 831 3336 832
rect 3330 827 3331 831
rect 3335 827 3336 831
rect 3330 826 3336 827
rect 3652 824 3654 885
rect 3748 832 3750 906
rect 3800 891 3802 955
rect 3840 939 3842 1003
rect 4780 939 4782 1004
rect 4906 999 4912 1000
rect 4906 995 4907 999
rect 4911 995 4912 999
rect 4906 994 4912 995
rect 4874 991 4880 992
rect 4874 987 4875 991
rect 4879 987 4880 991
rect 4874 986 4880 987
rect 4876 960 4878 986
rect 4908 960 4910 994
rect 4874 959 4880 960
rect 4874 955 4875 959
rect 4879 955 4880 959
rect 4874 954 4880 955
rect 4906 959 4912 960
rect 4906 955 4907 959
rect 4911 955 4912 959
rect 4906 954 4912 955
rect 4916 939 4918 1004
rect 5042 999 5048 1000
rect 5042 995 5043 999
rect 5047 995 5048 999
rect 5042 994 5048 995
rect 5044 960 5046 994
rect 5042 959 5048 960
rect 5042 955 5043 959
rect 5047 955 5048 959
rect 5042 954 5048 955
rect 5052 939 5054 1004
rect 5178 999 5184 1000
rect 5178 995 5179 999
rect 5183 995 5184 999
rect 5178 994 5184 995
rect 3839 938 3843 939
rect 3839 933 3843 934
rect 3859 938 3863 939
rect 3859 933 3863 934
rect 3995 938 3999 939
rect 3995 933 3999 934
rect 4171 938 4175 939
rect 4171 933 4175 934
rect 4387 938 4391 939
rect 4387 933 4391 934
rect 4643 938 4647 939
rect 4643 933 4647 934
rect 4779 938 4783 939
rect 4779 933 4783 934
rect 4915 938 4919 939
rect 4915 933 4919 934
rect 4931 938 4935 939
rect 4931 933 4935 934
rect 5051 938 5055 939
rect 5051 933 5055 934
rect 3799 890 3803 891
rect 3799 885 3803 886
rect 3746 831 3752 832
rect 3746 827 3747 831
rect 3751 827 3752 831
rect 3746 826 3752 827
rect 3800 825 3802 885
rect 3840 873 3842 933
rect 3838 872 3844 873
rect 3860 872 3862 933
rect 3954 919 3960 920
rect 3954 915 3955 919
rect 3959 915 3960 919
rect 3954 914 3960 915
rect 3838 868 3839 872
rect 3843 868 3844 872
rect 3838 867 3844 868
rect 3858 871 3864 872
rect 3858 867 3859 871
rect 3863 867 3864 871
rect 3858 866 3864 867
rect 3886 856 3892 857
rect 3838 855 3844 856
rect 3838 851 3839 855
rect 3843 851 3844 855
rect 3886 852 3887 856
rect 3891 852 3892 856
rect 3886 851 3892 852
rect 3838 850 3844 851
rect 3840 827 3842 850
rect 3888 827 3890 851
rect 3839 826 3843 827
rect 3798 824 3804 825
rect 1575 822 1579 823
rect 1575 817 1579 818
rect 1935 822 1939 823
rect 1974 820 1975 824
rect 1979 820 1980 824
rect 1974 819 1980 820
rect 1994 823 2000 824
rect 1994 819 1995 823
rect 1999 819 2000 823
rect 1994 818 2000 819
rect 2178 823 2184 824
rect 2178 819 2179 823
rect 2183 819 2184 823
rect 2178 818 2184 819
rect 2402 823 2408 824
rect 2402 819 2403 823
rect 2407 819 2408 823
rect 2402 818 2408 819
rect 2674 823 2680 824
rect 2674 819 2675 823
rect 2679 819 2680 823
rect 2674 818 2680 819
rect 2986 823 2992 824
rect 2986 819 2987 823
rect 2991 819 2992 823
rect 2986 818 2992 819
rect 3322 823 3328 824
rect 3322 819 3323 823
rect 3327 819 3328 823
rect 3322 818 3328 819
rect 3650 823 3656 824
rect 3650 819 3651 823
rect 3655 819 3656 823
rect 3798 820 3799 824
rect 3803 820 3804 824
rect 3839 821 3843 822
rect 3887 826 3891 827
rect 3887 821 3891 822
rect 3798 819 3804 820
rect 3650 818 3656 819
rect 1935 817 1939 818
rect 1576 793 1578 817
rect 1936 794 1938 817
rect 2022 808 2028 809
rect 1974 807 1980 808
rect 1974 803 1975 807
rect 1979 803 1980 807
rect 2022 804 2023 808
rect 2027 804 2028 808
rect 2022 803 2028 804
rect 2206 808 2212 809
rect 2206 804 2207 808
rect 2211 804 2212 808
rect 2206 803 2212 804
rect 2430 808 2436 809
rect 2430 804 2431 808
rect 2435 804 2436 808
rect 2430 803 2436 804
rect 2702 808 2708 809
rect 2702 804 2703 808
rect 2707 804 2708 808
rect 2702 803 2708 804
rect 3014 808 3020 809
rect 3014 804 3015 808
rect 3019 804 3020 808
rect 3014 803 3020 804
rect 3350 808 3356 809
rect 3350 804 3351 808
rect 3355 804 3356 808
rect 3350 803 3356 804
rect 3678 808 3684 809
rect 3678 804 3679 808
rect 3683 804 3684 808
rect 3678 803 3684 804
rect 3798 807 3804 808
rect 3798 803 3799 807
rect 3803 803 3804 807
rect 1974 802 1980 803
rect 1934 793 1940 794
rect 1574 792 1580 793
rect 1574 788 1575 792
rect 1579 788 1580 792
rect 1934 789 1935 793
rect 1939 789 1940 793
rect 1934 788 1940 789
rect 1574 787 1580 788
rect 1546 777 1552 778
rect 1546 773 1547 777
rect 1551 773 1552 777
rect 1546 772 1552 773
rect 1934 776 1940 777
rect 1934 772 1935 776
rect 1939 772 1940 776
rect 1482 727 1488 728
rect 1482 723 1483 727
rect 1487 723 1488 727
rect 1482 722 1488 723
rect 1490 727 1496 728
rect 1490 723 1491 727
rect 1495 723 1496 727
rect 1490 722 1496 723
rect 1548 711 1550 772
rect 1934 771 1940 772
rect 1936 711 1938 771
rect 875 710 879 711
rect 875 705 879 706
rect 907 710 911 711
rect 907 705 911 706
rect 1083 710 1087 711
rect 1083 705 1087 706
rect 1099 710 1103 711
rect 1099 705 1103 706
rect 1259 710 1263 711
rect 1259 705 1263 706
rect 1323 710 1327 711
rect 1323 705 1327 706
rect 1427 710 1431 711
rect 1427 705 1431 706
rect 1547 710 1551 711
rect 1547 705 1551 706
rect 1595 710 1599 711
rect 1595 705 1599 706
rect 1771 710 1775 711
rect 1771 705 1775 706
rect 1935 710 1939 711
rect 1935 705 1939 706
rect 766 695 772 696
rect 766 691 767 695
rect 771 691 772 695
rect 766 690 772 691
rect 908 644 910 705
rect 914 691 920 692
rect 914 687 915 691
rect 919 687 920 691
rect 914 686 920 687
rect 916 652 918 686
rect 914 651 920 652
rect 914 647 915 651
rect 919 647 920 651
rect 914 646 920 647
rect 1084 644 1086 705
rect 1260 644 1262 705
rect 1266 691 1272 692
rect 1266 687 1267 691
rect 1271 687 1272 691
rect 1266 686 1272 687
rect 1268 652 1270 686
rect 1266 651 1272 652
rect 1266 647 1267 651
rect 1271 647 1272 651
rect 1266 646 1272 647
rect 1428 644 1430 705
rect 1434 691 1440 692
rect 1434 687 1435 691
rect 1439 687 1440 691
rect 1434 686 1440 687
rect 1436 652 1438 686
rect 1434 651 1440 652
rect 1434 647 1435 651
rect 1439 647 1440 651
rect 1434 646 1440 647
rect 1596 644 1598 705
rect 1602 691 1608 692
rect 1602 687 1603 691
rect 1607 687 1608 691
rect 1602 686 1608 687
rect 1604 652 1606 686
rect 1602 651 1608 652
rect 1602 647 1603 651
rect 1607 647 1608 651
rect 1602 646 1608 647
rect 1772 644 1774 705
rect 1778 691 1784 692
rect 1778 687 1779 691
rect 1783 687 1784 691
rect 1778 686 1784 687
rect 1780 652 1782 686
rect 1778 651 1784 652
rect 1778 647 1779 651
rect 1783 647 1784 651
rect 1778 646 1784 647
rect 1894 651 1900 652
rect 1894 647 1895 651
rect 1899 647 1900 651
rect 1894 646 1900 647
rect 722 643 728 644
rect 722 639 723 643
rect 727 639 728 643
rect 722 638 728 639
rect 906 643 912 644
rect 906 639 907 643
rect 911 639 912 643
rect 906 638 912 639
rect 1082 643 1088 644
rect 1082 639 1083 643
rect 1087 639 1088 643
rect 1082 638 1088 639
rect 1258 643 1264 644
rect 1258 639 1259 643
rect 1263 639 1264 643
rect 1258 638 1264 639
rect 1426 643 1432 644
rect 1426 639 1427 643
rect 1431 639 1432 643
rect 1426 638 1432 639
rect 1594 643 1600 644
rect 1594 639 1595 643
rect 1599 639 1600 643
rect 1594 638 1600 639
rect 1770 643 1776 644
rect 1770 639 1771 643
rect 1775 639 1776 643
rect 1770 638 1776 639
rect 750 628 756 629
rect 750 624 751 628
rect 755 624 756 628
rect 750 623 756 624
rect 934 628 940 629
rect 934 624 935 628
rect 939 624 940 628
rect 934 623 940 624
rect 1110 628 1116 629
rect 1110 624 1111 628
rect 1115 624 1116 628
rect 1110 623 1116 624
rect 1286 628 1292 629
rect 1286 624 1287 628
rect 1291 624 1292 628
rect 1286 623 1292 624
rect 1454 628 1460 629
rect 1454 624 1455 628
rect 1459 624 1460 628
rect 1454 623 1460 624
rect 1622 628 1628 629
rect 1622 624 1623 628
rect 1627 624 1628 628
rect 1622 623 1628 624
rect 1798 628 1804 629
rect 1798 624 1799 628
rect 1803 624 1804 628
rect 1798 623 1804 624
rect 752 599 754 623
rect 936 599 938 623
rect 1112 599 1114 623
rect 1288 599 1290 623
rect 1456 599 1458 623
rect 1624 599 1626 623
rect 1800 599 1802 623
rect 751 598 755 599
rect 751 593 755 594
rect 807 598 811 599
rect 807 593 811 594
rect 935 598 939 599
rect 935 593 939 594
rect 999 598 1003 599
rect 999 593 1003 594
rect 1111 598 1115 599
rect 1111 593 1115 594
rect 1175 598 1179 599
rect 1175 593 1179 594
rect 1287 598 1291 599
rect 1287 593 1291 594
rect 1343 598 1347 599
rect 1343 593 1347 594
rect 1455 598 1459 599
rect 1455 593 1459 594
rect 1511 598 1515 599
rect 1511 593 1515 594
rect 1623 598 1627 599
rect 1623 593 1627 594
rect 1671 598 1675 599
rect 1671 593 1675 594
rect 1799 598 1803 599
rect 1799 593 1803 594
rect 1815 598 1819 599
rect 1815 593 1819 594
rect 808 569 810 593
rect 1000 569 1002 593
rect 1176 569 1178 593
rect 1344 569 1346 593
rect 1512 569 1514 593
rect 1672 569 1674 593
rect 1816 569 1818 593
rect 806 568 812 569
rect 806 564 807 568
rect 811 564 812 568
rect 806 563 812 564
rect 998 568 1004 569
rect 998 564 999 568
rect 1003 564 1004 568
rect 998 563 1004 564
rect 1174 568 1180 569
rect 1174 564 1175 568
rect 1179 564 1180 568
rect 1174 563 1180 564
rect 1342 568 1348 569
rect 1342 564 1343 568
rect 1347 564 1348 568
rect 1342 563 1348 564
rect 1510 568 1516 569
rect 1510 564 1511 568
rect 1515 564 1516 568
rect 1510 563 1516 564
rect 1670 568 1676 569
rect 1670 564 1671 568
rect 1675 564 1676 568
rect 1670 563 1676 564
rect 1814 568 1820 569
rect 1814 564 1815 568
rect 1819 564 1820 568
rect 1814 563 1820 564
rect 778 553 784 554
rect 778 549 779 553
rect 783 549 784 553
rect 778 548 784 549
rect 970 553 976 554
rect 970 549 971 553
rect 975 549 976 553
rect 970 548 976 549
rect 1146 553 1152 554
rect 1146 549 1147 553
rect 1151 549 1152 553
rect 1146 548 1152 549
rect 1314 553 1320 554
rect 1314 549 1315 553
rect 1319 549 1320 553
rect 1314 548 1320 549
rect 1482 553 1488 554
rect 1482 549 1483 553
rect 1487 549 1488 553
rect 1482 548 1488 549
rect 1642 553 1648 554
rect 1642 549 1643 553
rect 1647 549 1648 553
rect 1642 548 1648 549
rect 1786 553 1792 554
rect 1786 549 1787 553
rect 1791 549 1792 553
rect 1786 548 1792 549
rect 742 543 748 544
rect 742 539 743 543
rect 747 539 748 543
rect 742 538 748 539
rect 744 504 746 538
rect 646 503 652 504
rect 646 499 647 503
rect 651 499 652 503
rect 646 498 652 499
rect 742 503 748 504
rect 742 499 743 503
rect 747 499 748 503
rect 742 498 748 499
rect 780 487 782 548
rect 906 543 912 544
rect 906 539 907 543
rect 911 539 912 543
rect 906 538 912 539
rect 908 504 910 538
rect 906 503 912 504
rect 906 499 907 503
rect 911 499 912 503
rect 906 498 912 499
rect 972 487 974 548
rect 1148 487 1150 548
rect 1274 543 1280 544
rect 1274 539 1275 543
rect 1279 539 1280 543
rect 1274 538 1280 539
rect 1276 504 1278 538
rect 1274 503 1280 504
rect 1274 499 1275 503
rect 1279 499 1280 503
rect 1274 498 1280 499
rect 1316 487 1318 548
rect 1442 543 1448 544
rect 1442 539 1443 543
rect 1447 539 1448 543
rect 1442 538 1448 539
rect 1444 504 1446 538
rect 1442 503 1448 504
rect 1442 499 1443 503
rect 1447 499 1448 503
rect 1442 498 1448 499
rect 1484 487 1486 548
rect 1630 543 1636 544
rect 1630 539 1631 543
rect 1635 539 1636 543
rect 1630 538 1636 539
rect 1632 504 1634 538
rect 1630 503 1636 504
rect 1630 499 1631 503
rect 1635 499 1636 503
rect 1630 498 1636 499
rect 1644 487 1646 548
rect 1770 543 1776 544
rect 1770 539 1771 543
rect 1775 539 1776 543
rect 1770 538 1776 539
rect 1772 504 1774 538
rect 1770 503 1776 504
rect 1770 499 1771 503
rect 1775 499 1776 503
rect 1770 498 1776 499
rect 1788 487 1790 548
rect 1882 543 1888 544
rect 1882 539 1883 543
rect 1887 539 1888 543
rect 1882 538 1888 539
rect 347 486 351 487
rect 347 481 351 482
rect 483 486 487 487
rect 483 481 487 482
rect 571 486 575 487
rect 571 481 575 482
rect 779 486 783 487
rect 779 481 783 482
rect 811 486 815 487
rect 811 481 815 482
rect 971 486 975 487
rect 971 481 975 482
rect 1139 486 1143 487
rect 1139 481 1143 482
rect 1147 486 1151 487
rect 1147 481 1151 482
rect 1315 486 1319 487
rect 1315 481 1319 482
rect 1475 486 1479 487
rect 1475 481 1479 482
rect 1483 486 1487 487
rect 1483 481 1487 482
rect 1643 486 1647 487
rect 1643 481 1647 482
rect 1787 486 1791 487
rect 1787 481 1791 482
rect 250 467 256 468
rect 250 463 251 467
rect 255 463 256 467
rect 250 462 256 463
rect 252 436 254 462
rect 250 435 256 436
rect 250 431 251 435
rect 255 431 256 435
rect 250 430 256 431
rect 226 427 232 428
rect 226 423 227 427
rect 231 423 232 427
rect 226 422 232 423
rect 484 420 486 481
rect 578 467 584 468
rect 578 463 579 467
rect 583 463 584 467
rect 578 462 584 463
rect 110 416 111 420
rect 115 416 116 420
rect 110 415 116 416
rect 154 419 160 420
rect 154 415 155 419
rect 159 415 160 419
rect 154 414 160 415
rect 482 419 488 420
rect 482 415 483 419
rect 487 415 488 419
rect 482 414 488 415
rect 182 404 188 405
rect 110 403 116 404
rect 110 399 111 403
rect 115 399 116 403
rect 182 400 183 404
rect 187 400 188 404
rect 182 399 188 400
rect 510 404 516 405
rect 510 400 511 404
rect 515 400 516 404
rect 510 399 516 400
rect 110 398 116 399
rect 112 363 114 398
rect 184 363 186 399
rect 512 363 514 399
rect 111 362 115 363
rect 111 357 115 358
rect 183 362 187 363
rect 183 357 187 358
rect 279 362 283 363
rect 279 357 283 358
rect 487 362 491 363
rect 487 357 491 358
rect 511 362 515 363
rect 511 357 515 358
rect 112 334 114 357
rect 110 333 116 334
rect 280 333 282 357
rect 488 333 490 357
rect 110 329 111 333
rect 115 329 116 333
rect 110 328 116 329
rect 278 332 284 333
rect 278 328 279 332
rect 283 328 284 332
rect 278 327 284 328
rect 486 332 492 333
rect 486 328 487 332
rect 491 328 492 332
rect 486 327 492 328
rect 250 317 256 318
rect 110 316 116 317
rect 110 312 111 316
rect 115 312 116 316
rect 250 313 251 317
rect 255 313 256 317
rect 250 312 256 313
rect 458 317 464 318
rect 458 313 459 317
rect 463 313 464 317
rect 458 312 464 313
rect 110 311 116 312
rect 112 211 114 311
rect 252 211 254 312
rect 346 267 352 268
rect 346 263 347 267
rect 351 263 352 267
rect 346 262 352 263
rect 111 210 115 211
rect 111 205 115 206
rect 131 210 135 211
rect 131 205 135 206
rect 251 210 255 211
rect 251 205 255 206
rect 267 210 271 211
rect 267 205 271 206
rect 112 145 114 205
rect 110 144 116 145
rect 132 144 134 205
rect 226 191 232 192
rect 226 187 227 191
rect 231 187 232 191
rect 226 186 232 187
rect 228 160 230 186
rect 226 159 232 160
rect 226 155 227 159
rect 231 155 232 159
rect 226 154 232 155
rect 268 144 270 205
rect 274 191 280 192
rect 274 187 275 191
rect 279 187 280 191
rect 274 186 280 187
rect 276 152 278 186
rect 348 152 350 262
rect 460 211 462 312
rect 580 308 582 462
rect 812 420 814 481
rect 906 467 912 468
rect 906 463 907 467
rect 911 463 912 467
rect 906 462 912 463
rect 908 436 910 462
rect 906 435 912 436
rect 906 431 907 435
rect 911 431 912 435
rect 906 430 912 431
rect 934 427 940 428
rect 934 423 935 427
rect 939 423 940 427
rect 934 422 940 423
rect 810 419 816 420
rect 810 415 811 419
rect 815 415 816 419
rect 810 414 816 415
rect 838 404 844 405
rect 838 400 839 404
rect 843 400 844 404
rect 838 399 844 400
rect 840 363 842 399
rect 703 362 707 363
rect 703 357 707 358
rect 839 362 843 363
rect 839 357 843 358
rect 919 362 923 363
rect 919 357 923 358
rect 704 333 706 357
rect 920 333 922 357
rect 702 332 708 333
rect 702 328 703 332
rect 707 328 708 332
rect 702 327 708 328
rect 918 332 924 333
rect 918 328 919 332
rect 923 328 924 332
rect 918 327 924 328
rect 674 317 680 318
rect 674 313 675 317
rect 679 313 680 317
rect 674 312 680 313
rect 890 317 896 318
rect 890 313 891 317
rect 895 313 896 317
rect 890 312 896 313
rect 578 307 584 308
rect 578 303 579 307
rect 583 303 584 307
rect 578 302 584 303
rect 676 211 678 312
rect 770 299 776 300
rect 770 295 771 299
rect 775 295 776 299
rect 770 294 776 295
rect 772 268 774 294
rect 770 267 776 268
rect 770 263 771 267
rect 775 263 776 267
rect 770 262 776 263
rect 892 211 894 312
rect 936 268 938 422
rect 1140 420 1142 481
rect 1476 420 1478 481
rect 1482 467 1488 468
rect 1482 463 1483 467
rect 1487 463 1488 467
rect 1482 462 1488 463
rect 1484 428 1486 462
rect 1482 427 1488 428
rect 1482 423 1483 427
rect 1487 423 1488 427
rect 1482 422 1488 423
rect 1788 420 1790 481
rect 1884 472 1886 538
rect 1896 496 1898 646
rect 1936 645 1938 705
rect 1934 644 1940 645
rect 1934 640 1935 644
rect 1939 640 1940 644
rect 1934 639 1940 640
rect 1934 627 1940 628
rect 1934 623 1935 627
rect 1939 623 1940 627
rect 1934 622 1940 623
rect 1936 599 1938 622
rect 1935 598 1939 599
rect 1935 593 1939 594
rect 1936 570 1938 593
rect 1976 579 1978 802
rect 2024 579 2026 803
rect 2208 579 2210 803
rect 2432 579 2434 803
rect 2704 579 2706 803
rect 3016 579 3018 803
rect 3352 579 3354 803
rect 3680 579 3682 803
rect 3798 802 3804 803
rect 3800 579 3802 802
rect 3840 798 3842 821
rect 3838 797 3844 798
rect 3888 797 3890 821
rect 3838 793 3839 797
rect 3843 793 3844 797
rect 3838 792 3844 793
rect 3886 796 3892 797
rect 3886 792 3887 796
rect 3891 792 3892 796
rect 3886 791 3892 792
rect 3858 781 3864 782
rect 3838 780 3844 781
rect 3838 776 3839 780
rect 3843 776 3844 780
rect 3858 777 3859 781
rect 3863 777 3864 781
rect 3858 776 3864 777
rect 3838 775 3844 776
rect 3840 711 3842 775
rect 3860 711 3862 776
rect 3956 772 3958 914
rect 3996 872 3998 933
rect 4162 923 4168 924
rect 4162 919 4163 923
rect 4167 919 4168 923
rect 4162 918 4168 919
rect 4164 880 4166 918
rect 4090 879 4096 880
rect 4090 875 4091 879
rect 4095 875 4096 879
rect 4090 874 4096 875
rect 4162 879 4168 880
rect 4162 875 4163 879
rect 4167 875 4168 879
rect 4162 874 4168 875
rect 3994 871 4000 872
rect 3994 867 3995 871
rect 3999 867 4000 871
rect 3994 866 4000 867
rect 4022 856 4028 857
rect 4022 852 4023 856
rect 4027 852 4028 856
rect 4022 851 4028 852
rect 4024 827 4026 851
rect 4023 826 4027 827
rect 4023 821 4027 822
rect 4024 797 4026 821
rect 4022 796 4028 797
rect 4022 792 4023 796
rect 4027 792 4028 796
rect 4022 791 4028 792
rect 3994 781 4000 782
rect 3994 777 3995 781
rect 3999 777 4000 781
rect 3994 776 4000 777
rect 3954 771 3960 772
rect 3954 767 3955 771
rect 3959 767 3960 771
rect 3954 766 3960 767
rect 3954 731 3960 732
rect 3954 727 3955 731
rect 3959 727 3960 731
rect 3954 726 3960 727
rect 3839 710 3843 711
rect 3839 705 3843 706
rect 3859 710 3863 711
rect 3859 705 3863 706
rect 3840 645 3842 705
rect 3838 644 3844 645
rect 3860 644 3862 705
rect 3956 652 3958 726
rect 3996 711 3998 776
rect 4092 732 4094 874
rect 4172 872 4174 933
rect 4274 923 4280 924
rect 4274 919 4275 923
rect 4279 919 4280 923
rect 4274 918 4280 919
rect 4170 871 4176 872
rect 4170 867 4171 871
rect 4175 867 4176 871
rect 4170 866 4176 867
rect 4198 856 4204 857
rect 4198 852 4199 856
rect 4203 852 4204 856
rect 4198 851 4204 852
rect 4200 827 4202 851
rect 4159 826 4163 827
rect 4159 821 4163 822
rect 4199 826 4203 827
rect 4199 821 4203 822
rect 4160 797 4162 821
rect 4158 796 4164 797
rect 4158 792 4159 796
rect 4163 792 4164 796
rect 4158 791 4164 792
rect 4130 781 4136 782
rect 4130 777 4131 781
rect 4135 777 4136 781
rect 4130 776 4136 777
rect 4266 781 4272 782
rect 4266 777 4267 781
rect 4271 777 4272 781
rect 4266 776 4272 777
rect 4122 771 4128 772
rect 4122 767 4123 771
rect 4127 767 4128 771
rect 4122 766 4128 767
rect 4124 732 4126 766
rect 4090 731 4096 732
rect 4090 727 4091 731
rect 4095 727 4096 731
rect 4090 726 4096 727
rect 4122 731 4128 732
rect 4122 727 4123 731
rect 4127 727 4128 731
rect 4122 726 4128 727
rect 4132 711 4134 776
rect 4258 771 4264 772
rect 4258 767 4259 771
rect 4263 767 4264 771
rect 4258 766 4264 767
rect 4260 732 4262 766
rect 4258 731 4264 732
rect 4258 727 4259 731
rect 4263 727 4264 731
rect 4258 726 4264 727
rect 4268 711 4270 776
rect 4276 764 4278 918
rect 4388 872 4390 933
rect 4482 919 4488 920
rect 4482 915 4483 919
rect 4487 915 4488 919
rect 4482 914 4488 915
rect 4484 888 4486 914
rect 4482 887 4488 888
rect 4482 883 4483 887
rect 4487 883 4488 887
rect 4482 882 4488 883
rect 4644 872 4646 933
rect 4650 919 4656 920
rect 4650 915 4651 919
rect 4655 915 4656 919
rect 4650 914 4656 915
rect 4652 880 4654 914
rect 4650 879 4656 880
rect 4650 875 4651 879
rect 4655 875 4656 879
rect 4650 874 4656 875
rect 4932 872 4934 933
rect 5180 924 5182 994
rect 5188 939 5190 1004
rect 5324 939 5326 1004
rect 5330 999 5336 1000
rect 5330 995 5331 999
rect 5335 995 5336 999
rect 5330 994 5336 995
rect 5332 968 5334 994
rect 5330 967 5336 968
rect 5330 963 5331 967
rect 5335 963 5336 967
rect 5330 962 5336 963
rect 5420 960 5422 1106
rect 5458 1009 5464 1010
rect 5458 1005 5459 1009
rect 5463 1005 5464 1009
rect 5458 1004 5464 1005
rect 5418 959 5424 960
rect 5418 955 5419 959
rect 5423 955 5424 959
rect 5418 954 5424 955
rect 5460 939 5462 1004
rect 5480 1000 5482 1186
rect 5516 1171 5518 1236
rect 5612 1192 5614 1342
rect 5664 1341 5666 1401
rect 5662 1340 5668 1341
rect 5662 1336 5663 1340
rect 5667 1336 5668 1340
rect 5662 1335 5668 1336
rect 5662 1323 5668 1324
rect 5662 1319 5663 1323
rect 5667 1319 5668 1323
rect 5662 1318 5668 1319
rect 5664 1287 5666 1318
rect 5663 1286 5667 1287
rect 5663 1281 5667 1282
rect 5664 1258 5666 1281
rect 5662 1257 5668 1258
rect 5662 1253 5663 1257
rect 5667 1253 5668 1257
rect 5662 1252 5668 1253
rect 5662 1240 5668 1241
rect 5662 1236 5663 1240
rect 5667 1236 5668 1240
rect 5662 1235 5668 1236
rect 5618 1231 5624 1232
rect 5618 1227 5619 1231
rect 5623 1227 5624 1231
rect 5618 1226 5624 1227
rect 5610 1191 5616 1192
rect 5610 1187 5611 1191
rect 5615 1187 5616 1191
rect 5610 1186 5616 1187
rect 5515 1170 5519 1171
rect 5515 1165 5519 1166
rect 5516 1104 5518 1165
rect 5620 1156 5622 1226
rect 5664 1171 5666 1235
rect 5663 1170 5667 1171
rect 5663 1165 5667 1166
rect 5618 1155 5624 1156
rect 5618 1151 5619 1155
rect 5623 1151 5624 1155
rect 5618 1150 5624 1151
rect 5610 1111 5616 1112
rect 5610 1107 5611 1111
rect 5615 1107 5616 1111
rect 5610 1106 5616 1107
rect 5514 1103 5520 1104
rect 5514 1099 5515 1103
rect 5519 1099 5520 1103
rect 5514 1098 5520 1099
rect 5542 1088 5548 1089
rect 5542 1084 5543 1088
rect 5547 1084 5548 1088
rect 5542 1083 5548 1084
rect 5544 1055 5546 1083
rect 5487 1054 5491 1055
rect 5487 1049 5491 1050
rect 5543 1054 5547 1055
rect 5543 1049 5547 1050
rect 5488 1025 5490 1049
rect 5486 1024 5492 1025
rect 5486 1020 5487 1024
rect 5491 1020 5492 1024
rect 5486 1019 5492 1020
rect 5478 999 5484 1000
rect 5478 995 5479 999
rect 5483 995 5484 999
rect 5478 994 5484 995
rect 5554 959 5560 960
rect 5554 955 5555 959
rect 5559 955 5560 959
rect 5554 954 5560 955
rect 5187 938 5191 939
rect 5187 933 5191 934
rect 5235 938 5239 939
rect 5235 933 5239 934
rect 5323 938 5327 939
rect 5323 933 5327 934
rect 5459 938 5463 939
rect 5459 933 5463 934
rect 5515 938 5519 939
rect 5515 933 5519 934
rect 5178 923 5184 924
rect 4938 919 4944 920
rect 4938 915 4939 919
rect 4943 915 4944 919
rect 5178 919 5179 923
rect 5183 919 5184 923
rect 5178 918 5184 919
rect 4938 914 4944 915
rect 4940 880 4942 914
rect 4938 879 4944 880
rect 4938 875 4939 879
rect 4943 875 4944 879
rect 4938 874 4944 875
rect 5066 879 5072 880
rect 5066 875 5067 879
rect 5071 875 5072 879
rect 5066 874 5072 875
rect 4386 871 4392 872
rect 4386 867 4387 871
rect 4391 867 4392 871
rect 4386 866 4392 867
rect 4642 871 4648 872
rect 4642 867 4643 871
rect 4647 867 4648 871
rect 4642 866 4648 867
rect 4930 871 4936 872
rect 4930 867 4931 871
rect 4935 867 4936 871
rect 4930 866 4936 867
rect 4414 856 4420 857
rect 4414 852 4415 856
rect 4419 852 4420 856
rect 4414 851 4420 852
rect 4670 856 4676 857
rect 4670 852 4671 856
rect 4675 852 4676 856
rect 4670 851 4676 852
rect 4958 856 4964 857
rect 4958 852 4959 856
rect 4963 852 4964 856
rect 4958 851 4964 852
rect 4416 827 4418 851
rect 4672 827 4674 851
rect 4960 827 4962 851
rect 4295 826 4299 827
rect 4295 821 4299 822
rect 4415 826 4419 827
rect 4415 821 4419 822
rect 4431 826 4435 827
rect 4431 821 4435 822
rect 4567 826 4571 827
rect 4567 821 4571 822
rect 4671 826 4675 827
rect 4671 821 4675 822
rect 4719 826 4723 827
rect 4719 821 4723 822
rect 4895 826 4899 827
rect 4895 821 4899 822
rect 4959 826 4963 827
rect 4959 821 4963 822
rect 4296 797 4298 821
rect 4432 797 4434 821
rect 4568 797 4570 821
rect 4720 797 4722 821
rect 4896 797 4898 821
rect 4294 796 4300 797
rect 4294 792 4295 796
rect 4299 792 4300 796
rect 4294 791 4300 792
rect 4430 796 4436 797
rect 4430 792 4431 796
rect 4435 792 4436 796
rect 4430 791 4436 792
rect 4566 796 4572 797
rect 4566 792 4567 796
rect 4571 792 4572 796
rect 4566 791 4572 792
rect 4718 796 4724 797
rect 4718 792 4719 796
rect 4723 792 4724 796
rect 4718 791 4724 792
rect 4894 796 4900 797
rect 4894 792 4895 796
rect 4899 792 4900 796
rect 4894 791 4900 792
rect 4402 781 4408 782
rect 4402 777 4403 781
rect 4407 777 4408 781
rect 4402 776 4408 777
rect 4538 781 4544 782
rect 4538 777 4539 781
rect 4543 777 4544 781
rect 4538 776 4544 777
rect 4690 781 4696 782
rect 4690 777 4691 781
rect 4695 777 4696 781
rect 4690 776 4696 777
rect 4866 781 4872 782
rect 4866 777 4867 781
rect 4871 777 4872 781
rect 4866 776 4872 777
rect 5058 781 5064 782
rect 5058 777 5059 781
rect 5063 777 5064 781
rect 5058 776 5064 777
rect 4394 771 4400 772
rect 4394 767 4395 771
rect 4399 767 4400 771
rect 4394 766 4400 767
rect 4274 763 4280 764
rect 4274 759 4275 763
rect 4279 759 4280 763
rect 4274 758 4280 759
rect 4396 732 4398 766
rect 4394 731 4400 732
rect 4394 727 4395 731
rect 4399 727 4400 731
rect 4394 726 4400 727
rect 4404 711 4406 776
rect 4530 771 4536 772
rect 4530 767 4531 771
rect 4535 767 4536 771
rect 4530 766 4536 767
rect 4532 732 4534 766
rect 4530 731 4536 732
rect 4530 727 4531 731
rect 4535 727 4536 731
rect 4530 726 4536 727
rect 4540 711 4542 776
rect 4634 771 4640 772
rect 4634 767 4635 771
rect 4639 767 4640 771
rect 4634 766 4640 767
rect 3995 710 3999 711
rect 3995 705 3999 706
rect 4131 710 4135 711
rect 4131 705 4135 706
rect 4267 710 4271 711
rect 4267 705 4271 706
rect 4403 710 4407 711
rect 4403 705 4407 706
rect 4539 710 4543 711
rect 4539 705 4543 706
rect 3954 651 3960 652
rect 3954 647 3955 651
rect 3959 647 3960 651
rect 3954 646 3960 647
rect 3996 644 3998 705
rect 4002 691 4008 692
rect 4002 687 4003 691
rect 4007 687 4008 691
rect 4002 686 4008 687
rect 3838 640 3839 644
rect 3843 640 3844 644
rect 3838 639 3844 640
rect 3858 643 3864 644
rect 3858 639 3859 643
rect 3863 639 3864 643
rect 3858 638 3864 639
rect 3994 643 4000 644
rect 3994 639 3995 643
rect 3999 639 4000 643
rect 3994 638 4000 639
rect 3886 628 3892 629
rect 3838 627 3844 628
rect 3838 623 3839 627
rect 3843 623 3844 627
rect 3886 624 3887 628
rect 3891 624 3892 628
rect 3886 623 3892 624
rect 3838 622 3844 623
rect 3840 599 3842 622
rect 3888 599 3890 623
rect 3839 598 3843 599
rect 3839 593 3843 594
rect 3887 598 3891 599
rect 3887 593 3891 594
rect 1975 578 1979 579
rect 1975 573 1979 574
rect 2023 578 2027 579
rect 2023 573 2027 574
rect 2207 578 2211 579
rect 2207 573 2211 574
rect 2431 578 2435 579
rect 2431 573 2435 574
rect 2703 578 2707 579
rect 2703 573 2707 574
rect 3015 578 3019 579
rect 3015 573 3019 574
rect 3135 578 3139 579
rect 3135 573 3139 574
rect 3271 578 3275 579
rect 3271 573 3275 574
rect 3351 578 3355 579
rect 3351 573 3355 574
rect 3407 578 3411 579
rect 3407 573 3411 574
rect 3543 578 3547 579
rect 3543 573 3547 574
rect 3679 578 3683 579
rect 3679 573 3683 574
rect 3799 578 3803 579
rect 3799 573 3803 574
rect 1934 569 1940 570
rect 1934 565 1935 569
rect 1939 565 1940 569
rect 1934 564 1940 565
rect 1934 552 1940 553
rect 1934 548 1935 552
rect 1939 548 1940 552
rect 1976 550 1978 573
rect 1934 547 1940 548
rect 1974 549 1980 550
rect 3136 549 3138 573
rect 3272 549 3274 573
rect 3408 549 3410 573
rect 3544 549 3546 573
rect 3680 549 3682 573
rect 3800 550 3802 573
rect 3840 570 3842 593
rect 3838 569 3844 570
rect 3888 569 3890 593
rect 3838 565 3839 569
rect 3843 565 3844 569
rect 3838 564 3844 565
rect 3886 568 3892 569
rect 3886 564 3887 568
rect 3891 564 3892 568
rect 3886 563 3892 564
rect 3858 553 3864 554
rect 3838 552 3844 553
rect 3798 549 3804 550
rect 1894 495 1900 496
rect 1894 491 1895 495
rect 1899 491 1900 495
rect 1894 490 1900 491
rect 1936 487 1938 547
rect 1974 545 1975 549
rect 1979 545 1980 549
rect 1974 544 1980 545
rect 3134 548 3140 549
rect 3134 544 3135 548
rect 3139 544 3140 548
rect 3134 543 3140 544
rect 3270 548 3276 549
rect 3270 544 3271 548
rect 3275 544 3276 548
rect 3270 543 3276 544
rect 3406 548 3412 549
rect 3406 544 3407 548
rect 3411 544 3412 548
rect 3406 543 3412 544
rect 3542 548 3548 549
rect 3542 544 3543 548
rect 3547 544 3548 548
rect 3542 543 3548 544
rect 3678 548 3684 549
rect 3678 544 3679 548
rect 3683 544 3684 548
rect 3798 545 3799 549
rect 3803 545 3804 549
rect 3838 548 3839 552
rect 3843 548 3844 552
rect 3858 549 3859 553
rect 3863 549 3864 553
rect 3858 548 3864 549
rect 3838 547 3844 548
rect 3798 544 3804 545
rect 3678 543 3684 544
rect 3106 533 3112 534
rect 1974 532 1980 533
rect 1974 528 1975 532
rect 1979 528 1980 532
rect 3106 529 3107 533
rect 3111 529 3112 533
rect 3106 528 3112 529
rect 3242 533 3248 534
rect 3242 529 3243 533
rect 3247 529 3248 533
rect 3242 528 3248 529
rect 3378 533 3384 534
rect 3378 529 3379 533
rect 3383 529 3384 533
rect 3378 528 3384 529
rect 3514 533 3520 534
rect 3514 529 3515 533
rect 3519 529 3520 533
rect 3514 528 3520 529
rect 3650 533 3656 534
rect 3650 529 3651 533
rect 3655 529 3656 533
rect 3650 528 3656 529
rect 3798 532 3804 533
rect 3798 528 3799 532
rect 3803 528 3804 532
rect 1974 527 1980 528
rect 1935 486 1939 487
rect 1935 481 1939 482
rect 1882 471 1888 472
rect 1882 467 1883 471
rect 1887 467 1888 471
rect 1882 466 1888 467
rect 1914 451 1920 452
rect 1914 447 1915 451
rect 1919 447 1920 451
rect 1914 446 1920 447
rect 1916 428 1918 446
rect 1914 427 1920 428
rect 1914 423 1915 427
rect 1919 423 1920 427
rect 1914 422 1920 423
rect 1936 421 1938 481
rect 1976 467 1978 527
rect 3108 467 3110 528
rect 3234 523 3240 524
rect 3234 519 3235 523
rect 3239 519 3240 523
rect 3234 518 3240 519
rect 3236 484 3238 518
rect 3202 483 3208 484
rect 3202 479 3203 483
rect 3207 479 3208 483
rect 3202 478 3208 479
rect 3234 483 3240 484
rect 3234 479 3235 483
rect 3239 479 3240 483
rect 3234 478 3240 479
rect 1975 466 1979 467
rect 1975 461 1979 462
rect 1995 466 1999 467
rect 1995 461 1999 462
rect 2203 466 2207 467
rect 2203 461 2207 462
rect 2427 466 2431 467
rect 2427 461 2431 462
rect 2651 466 2655 467
rect 2651 461 2655 462
rect 2859 466 2863 467
rect 2859 461 2863 462
rect 3067 466 3071 467
rect 3067 461 3071 462
rect 3107 466 3111 467
rect 3107 461 3111 462
rect 1934 420 1940 421
rect 1138 419 1144 420
rect 1138 415 1139 419
rect 1143 415 1144 419
rect 1138 414 1144 415
rect 1474 419 1480 420
rect 1474 415 1475 419
rect 1479 415 1480 419
rect 1474 414 1480 415
rect 1786 419 1792 420
rect 1786 415 1787 419
rect 1791 415 1792 419
rect 1934 416 1935 420
rect 1939 416 1940 420
rect 1934 415 1940 416
rect 1786 414 1792 415
rect 1166 404 1172 405
rect 1166 400 1167 404
rect 1171 400 1172 404
rect 1166 399 1172 400
rect 1502 404 1508 405
rect 1502 400 1503 404
rect 1507 400 1508 404
rect 1502 399 1508 400
rect 1814 404 1820 405
rect 1814 400 1815 404
rect 1819 400 1820 404
rect 1814 399 1820 400
rect 1934 403 1940 404
rect 1934 399 1935 403
rect 1939 399 1940 403
rect 1976 401 1978 461
rect 1168 363 1170 399
rect 1504 363 1506 399
rect 1816 363 1818 399
rect 1934 398 1940 399
rect 1974 400 1980 401
rect 1996 400 1998 461
rect 2204 400 2206 461
rect 2210 447 2216 448
rect 2210 443 2211 447
rect 2215 443 2216 447
rect 2210 442 2216 443
rect 2212 408 2214 442
rect 2210 407 2216 408
rect 2210 403 2211 407
rect 2215 403 2216 407
rect 2210 402 2216 403
rect 2428 400 2430 461
rect 2434 447 2440 448
rect 2434 443 2435 447
rect 2439 443 2440 447
rect 2434 442 2440 443
rect 2436 408 2438 442
rect 2434 407 2440 408
rect 2434 403 2435 407
rect 2439 403 2440 407
rect 2434 402 2440 403
rect 2652 400 2654 461
rect 2658 447 2664 448
rect 2658 443 2659 447
rect 2663 443 2664 447
rect 2658 442 2664 443
rect 2660 408 2662 442
rect 2658 407 2664 408
rect 2658 403 2659 407
rect 2663 403 2664 407
rect 2658 402 2664 403
rect 2686 407 2692 408
rect 2686 403 2687 407
rect 2691 403 2692 407
rect 2686 402 2692 403
rect 1936 363 1938 398
rect 1974 396 1975 400
rect 1979 396 1980 400
rect 1974 395 1980 396
rect 1994 399 2000 400
rect 1994 395 1995 399
rect 1999 395 2000 399
rect 1994 394 2000 395
rect 2202 399 2208 400
rect 2202 395 2203 399
rect 2207 395 2208 399
rect 2202 394 2208 395
rect 2426 399 2432 400
rect 2426 395 2427 399
rect 2431 395 2432 399
rect 2426 394 2432 395
rect 2650 399 2656 400
rect 2650 395 2651 399
rect 2655 395 2656 399
rect 2650 394 2656 395
rect 2022 384 2028 385
rect 1974 383 1980 384
rect 1974 379 1975 383
rect 1979 379 1980 383
rect 2022 380 2023 384
rect 2027 380 2028 384
rect 2022 379 2028 380
rect 2230 384 2236 385
rect 2230 380 2231 384
rect 2235 380 2236 384
rect 2230 379 2236 380
rect 2454 384 2460 385
rect 2454 380 2455 384
rect 2459 380 2460 384
rect 2454 379 2460 380
rect 2678 384 2684 385
rect 2678 380 2679 384
rect 2683 380 2684 384
rect 2678 379 2684 380
rect 1974 378 1980 379
rect 1135 362 1139 363
rect 1135 357 1139 358
rect 1167 362 1171 363
rect 1167 357 1171 358
rect 1503 362 1507 363
rect 1503 357 1507 358
rect 1815 362 1819 363
rect 1815 357 1819 358
rect 1935 362 1939 363
rect 1935 357 1939 358
rect 1136 333 1138 357
rect 1936 334 1938 357
rect 1976 339 1978 378
rect 2024 339 2026 379
rect 2232 339 2234 379
rect 2456 339 2458 379
rect 2680 339 2682 379
rect 1975 338 1979 339
rect 1934 333 1940 334
rect 1975 333 1979 334
rect 2023 338 2027 339
rect 2023 333 2027 334
rect 2159 338 2163 339
rect 2159 333 2163 334
rect 2231 338 2235 339
rect 2231 333 2235 334
rect 2295 338 2299 339
rect 2295 333 2299 334
rect 2431 338 2435 339
rect 2431 333 2435 334
rect 2455 338 2459 339
rect 2455 333 2459 334
rect 2567 338 2571 339
rect 2567 333 2571 334
rect 2679 338 2683 339
rect 2679 333 2683 334
rect 1134 332 1140 333
rect 1134 328 1135 332
rect 1139 328 1140 332
rect 1934 329 1935 333
rect 1939 329 1940 333
rect 1934 328 1940 329
rect 1134 327 1140 328
rect 1106 317 1112 318
rect 1106 313 1107 317
rect 1111 313 1112 317
rect 1106 312 1112 313
rect 1934 316 1940 317
rect 1934 312 1935 316
rect 1939 312 1940 316
rect 1062 307 1068 308
rect 1062 303 1063 307
rect 1067 303 1068 307
rect 1062 302 1068 303
rect 1064 268 1066 302
rect 934 267 940 268
rect 934 263 935 267
rect 939 263 940 267
rect 934 262 940 263
rect 1062 267 1068 268
rect 1062 263 1063 267
rect 1067 263 1068 267
rect 1062 262 1068 263
rect 1108 211 1110 312
rect 1934 311 1940 312
rect 1936 211 1938 311
rect 1976 310 1978 333
rect 1974 309 1980 310
rect 2024 309 2026 333
rect 2160 309 2162 333
rect 2296 309 2298 333
rect 2432 309 2434 333
rect 2568 309 2570 333
rect 1974 305 1975 309
rect 1979 305 1980 309
rect 1974 304 1980 305
rect 2022 308 2028 309
rect 2022 304 2023 308
rect 2027 304 2028 308
rect 2022 303 2028 304
rect 2158 308 2164 309
rect 2158 304 2159 308
rect 2163 304 2164 308
rect 2158 303 2164 304
rect 2294 308 2300 309
rect 2294 304 2295 308
rect 2299 304 2300 308
rect 2294 303 2300 304
rect 2430 308 2436 309
rect 2430 304 2431 308
rect 2435 304 2436 308
rect 2430 303 2436 304
rect 2566 308 2572 309
rect 2566 304 2567 308
rect 2571 304 2572 308
rect 2566 303 2572 304
rect 1994 293 2000 294
rect 1974 292 1980 293
rect 1974 288 1975 292
rect 1979 288 1980 292
rect 1994 289 1995 293
rect 1999 289 2000 293
rect 1994 288 2000 289
rect 2130 293 2136 294
rect 2130 289 2131 293
rect 2135 289 2136 293
rect 2130 288 2136 289
rect 2266 293 2272 294
rect 2266 289 2267 293
rect 2271 289 2272 293
rect 2266 288 2272 289
rect 2402 293 2408 294
rect 2402 289 2403 293
rect 2407 289 2408 293
rect 2402 288 2408 289
rect 2538 293 2544 294
rect 2538 289 2539 293
rect 2543 289 2544 293
rect 2538 288 2544 289
rect 2674 293 2680 294
rect 2674 289 2675 293
rect 2679 289 2680 293
rect 2674 288 2680 289
rect 1974 287 1980 288
rect 403 210 407 211
rect 403 205 407 206
rect 459 210 463 211
rect 459 205 463 206
rect 539 210 543 211
rect 539 205 543 206
rect 675 210 679 211
rect 675 205 679 206
rect 811 210 815 211
rect 811 205 815 206
rect 891 210 895 211
rect 891 205 895 206
rect 947 210 951 211
rect 947 205 951 206
rect 1083 210 1087 211
rect 1083 205 1087 206
rect 1107 210 1111 211
rect 1107 205 1111 206
rect 1935 210 1939 211
rect 1935 205 1939 206
rect 274 151 280 152
rect 274 147 275 151
rect 279 147 280 151
rect 274 146 280 147
rect 346 151 352 152
rect 346 147 347 151
rect 351 147 352 151
rect 346 146 352 147
rect 404 144 406 205
rect 540 144 542 205
rect 634 191 640 192
rect 634 187 635 191
rect 639 187 640 191
rect 634 186 640 187
rect 636 160 638 186
rect 634 159 640 160
rect 634 155 635 159
rect 639 155 640 159
rect 634 154 640 155
rect 676 144 678 205
rect 812 144 814 205
rect 948 144 950 205
rect 954 191 960 192
rect 954 187 955 191
rect 959 187 960 191
rect 954 186 960 187
rect 956 152 958 186
rect 954 151 960 152
rect 954 147 955 151
rect 959 147 960 151
rect 954 146 960 147
rect 1084 144 1086 205
rect 1206 203 1212 204
rect 1206 199 1207 203
rect 1211 199 1212 203
rect 1206 198 1212 199
rect 1090 191 1096 192
rect 1090 187 1091 191
rect 1095 187 1096 191
rect 1090 186 1096 187
rect 1092 152 1094 186
rect 1208 152 1210 198
rect 1090 151 1096 152
rect 1090 147 1091 151
rect 1095 147 1096 151
rect 1090 146 1096 147
rect 1206 151 1212 152
rect 1206 147 1207 151
rect 1211 147 1212 151
rect 1206 146 1212 147
rect 1936 145 1938 205
rect 1976 191 1978 287
rect 1996 191 1998 288
rect 2122 283 2128 284
rect 2122 279 2123 283
rect 2127 279 2128 283
rect 2122 278 2128 279
rect 2090 275 2096 276
rect 2090 271 2091 275
rect 2095 271 2096 275
rect 2090 270 2096 271
rect 2092 244 2094 270
rect 2124 244 2126 278
rect 2090 243 2096 244
rect 2090 239 2091 243
rect 2095 239 2096 243
rect 2090 238 2096 239
rect 2122 243 2128 244
rect 2122 239 2123 243
rect 2127 239 2128 243
rect 2122 238 2128 239
rect 2090 235 2096 236
rect 2090 231 2091 235
rect 2095 231 2096 235
rect 2090 230 2096 231
rect 1975 190 1979 191
rect 1975 185 1979 186
rect 1995 190 1999 191
rect 1995 185 1999 186
rect 1934 144 1940 145
rect 110 140 111 144
rect 115 140 116 144
rect 110 139 116 140
rect 130 143 136 144
rect 130 139 131 143
rect 135 139 136 143
rect 130 138 136 139
rect 266 143 272 144
rect 266 139 267 143
rect 271 139 272 143
rect 266 138 272 139
rect 402 143 408 144
rect 402 139 403 143
rect 407 139 408 143
rect 402 138 408 139
rect 538 143 544 144
rect 538 139 539 143
rect 543 139 544 143
rect 538 138 544 139
rect 674 143 680 144
rect 674 139 675 143
rect 679 139 680 143
rect 674 138 680 139
rect 810 143 816 144
rect 810 139 811 143
rect 815 139 816 143
rect 810 138 816 139
rect 946 143 952 144
rect 946 139 947 143
rect 951 139 952 143
rect 946 138 952 139
rect 1082 143 1088 144
rect 1082 139 1083 143
rect 1087 139 1088 143
rect 1934 140 1935 144
rect 1939 140 1940 144
rect 1934 139 1940 140
rect 1082 138 1088 139
rect 158 128 164 129
rect 110 127 116 128
rect 110 123 111 127
rect 115 123 116 127
rect 158 124 159 128
rect 163 124 164 128
rect 158 123 164 124
rect 294 128 300 129
rect 294 124 295 128
rect 299 124 300 128
rect 294 123 300 124
rect 430 128 436 129
rect 430 124 431 128
rect 435 124 436 128
rect 430 123 436 124
rect 566 128 572 129
rect 566 124 567 128
rect 571 124 572 128
rect 566 123 572 124
rect 702 128 708 129
rect 702 124 703 128
rect 707 124 708 128
rect 702 123 708 124
rect 838 128 844 129
rect 838 124 839 128
rect 843 124 844 128
rect 838 123 844 124
rect 974 128 980 129
rect 974 124 975 128
rect 979 124 980 128
rect 974 123 980 124
rect 1110 128 1116 129
rect 1110 124 1111 128
rect 1115 124 1116 128
rect 1110 123 1116 124
rect 1934 127 1940 128
rect 1934 123 1935 127
rect 1939 123 1940 127
rect 1976 125 1978 185
rect 110 122 116 123
rect 112 99 114 122
rect 160 99 162 123
rect 296 99 298 123
rect 432 99 434 123
rect 568 99 570 123
rect 704 99 706 123
rect 840 99 842 123
rect 976 99 978 123
rect 1112 99 1114 123
rect 1934 122 1940 123
rect 1974 124 1980 125
rect 1996 124 1998 185
rect 2092 176 2094 230
rect 2132 191 2134 288
rect 2258 283 2264 284
rect 2258 279 2259 283
rect 2263 279 2264 283
rect 2258 278 2264 279
rect 2260 244 2262 278
rect 2258 243 2264 244
rect 2258 239 2259 243
rect 2263 239 2264 243
rect 2258 238 2264 239
rect 2268 191 2270 288
rect 2394 283 2400 284
rect 2394 279 2395 283
rect 2399 279 2400 283
rect 2394 278 2400 279
rect 2396 244 2398 278
rect 2394 243 2400 244
rect 2394 239 2395 243
rect 2399 239 2400 243
rect 2394 238 2400 239
rect 2404 191 2406 288
rect 2530 283 2536 284
rect 2530 279 2531 283
rect 2535 279 2536 283
rect 2530 278 2536 279
rect 2532 244 2534 278
rect 2530 243 2536 244
rect 2530 239 2531 243
rect 2535 239 2536 243
rect 2530 238 2536 239
rect 2540 191 2542 288
rect 2666 283 2672 284
rect 2666 279 2667 283
rect 2671 279 2672 283
rect 2666 278 2672 279
rect 2668 244 2670 278
rect 2666 243 2672 244
rect 2666 239 2667 243
rect 2671 239 2672 243
rect 2666 238 2672 239
rect 2676 191 2678 288
rect 2688 276 2690 402
rect 2860 400 2862 461
rect 2954 447 2960 448
rect 2954 443 2955 447
rect 2959 443 2960 447
rect 2954 442 2960 443
rect 2858 399 2864 400
rect 2858 395 2859 399
rect 2863 395 2864 399
rect 2858 394 2864 395
rect 2886 384 2892 385
rect 2886 380 2887 384
rect 2891 380 2892 384
rect 2886 379 2892 380
rect 2888 339 2890 379
rect 2703 338 2707 339
rect 2703 333 2707 334
rect 2839 338 2843 339
rect 2839 333 2843 334
rect 2887 338 2891 339
rect 2887 333 2891 334
rect 2704 309 2706 333
rect 2840 309 2842 333
rect 2702 308 2708 309
rect 2702 304 2703 308
rect 2707 304 2708 308
rect 2702 303 2708 304
rect 2838 308 2844 309
rect 2838 304 2839 308
rect 2843 304 2844 308
rect 2838 303 2844 304
rect 2810 293 2816 294
rect 2810 289 2811 293
rect 2815 289 2816 293
rect 2810 288 2816 289
rect 2946 293 2952 294
rect 2946 289 2947 293
rect 2951 289 2952 293
rect 2946 288 2952 289
rect 2802 283 2808 284
rect 2802 279 2803 283
rect 2807 279 2808 283
rect 2802 278 2808 279
rect 2686 275 2692 276
rect 2686 271 2687 275
rect 2691 271 2692 275
rect 2686 270 2692 271
rect 2804 244 2806 278
rect 2802 243 2808 244
rect 2802 239 2803 243
rect 2807 239 2808 243
rect 2802 238 2808 239
rect 2812 191 2814 288
rect 2854 283 2860 284
rect 2854 279 2855 283
rect 2859 279 2860 283
rect 2854 278 2860 279
rect 2856 236 2858 278
rect 2854 235 2860 236
rect 2854 231 2855 235
rect 2859 231 2860 235
rect 2854 230 2860 231
rect 2948 191 2950 288
rect 2956 268 2958 442
rect 3068 400 3070 461
rect 3074 447 3080 448
rect 3074 443 3075 447
rect 3079 443 3080 447
rect 3074 442 3080 443
rect 3076 408 3078 442
rect 3204 416 3206 478
rect 3244 467 3246 528
rect 3370 523 3376 524
rect 3370 519 3371 523
rect 3375 519 3376 523
rect 3370 518 3376 519
rect 3372 484 3374 518
rect 3370 483 3376 484
rect 3370 479 3371 483
rect 3375 479 3376 483
rect 3370 478 3376 479
rect 3380 467 3382 528
rect 3506 523 3512 524
rect 3506 519 3507 523
rect 3511 519 3512 523
rect 3506 518 3512 519
rect 3508 484 3510 518
rect 3506 483 3512 484
rect 3506 479 3507 483
rect 3511 479 3512 483
rect 3506 478 3512 479
rect 3516 467 3518 528
rect 3642 523 3648 524
rect 3642 519 3643 523
rect 3647 519 3648 523
rect 3642 518 3648 519
rect 3644 484 3646 518
rect 3642 483 3648 484
rect 3642 479 3643 483
rect 3647 479 3648 483
rect 3642 478 3648 479
rect 3652 467 3654 528
rect 3798 527 3804 528
rect 3778 523 3784 524
rect 3778 519 3779 523
rect 3783 519 3784 523
rect 3778 518 3784 519
rect 3780 504 3782 518
rect 3778 503 3784 504
rect 3778 499 3779 503
rect 3783 499 3784 503
rect 3778 498 3784 499
rect 3800 467 3802 527
rect 3840 475 3842 547
rect 3860 475 3862 548
rect 4004 544 4006 686
rect 4132 644 4134 705
rect 4138 691 4144 692
rect 4138 687 4139 691
rect 4143 687 4144 691
rect 4138 686 4144 687
rect 4140 652 4142 686
rect 4138 651 4144 652
rect 4138 647 4139 651
rect 4143 647 4144 651
rect 4138 646 4144 647
rect 4268 644 4270 705
rect 4274 691 4280 692
rect 4274 687 4275 691
rect 4279 687 4280 691
rect 4274 686 4280 687
rect 4276 652 4278 686
rect 4274 651 4280 652
rect 4274 647 4275 651
rect 4279 647 4280 651
rect 4274 646 4280 647
rect 4404 644 4406 705
rect 4410 691 4416 692
rect 4410 687 4411 691
rect 4415 687 4416 691
rect 4410 686 4416 687
rect 4412 652 4414 686
rect 4410 651 4416 652
rect 4410 647 4411 651
rect 4415 647 4416 651
rect 4410 646 4416 647
rect 4540 644 4542 705
rect 4636 696 4638 766
rect 4692 711 4694 776
rect 4842 771 4848 772
rect 4842 767 4843 771
rect 4847 767 4848 771
rect 4842 766 4848 767
rect 4844 732 4846 766
rect 4842 731 4848 732
rect 4842 727 4843 731
rect 4847 727 4848 731
rect 4842 726 4848 727
rect 4868 711 4870 776
rect 4962 763 4968 764
rect 4962 759 4963 763
rect 4967 759 4968 763
rect 4962 758 4968 759
rect 4964 732 4966 758
rect 4962 731 4968 732
rect 4962 727 4963 731
rect 4967 727 4968 731
rect 4962 726 4968 727
rect 5060 711 5062 776
rect 5068 732 5070 874
rect 5236 872 5238 933
rect 5516 872 5518 933
rect 5234 871 5240 872
rect 5234 867 5235 871
rect 5239 867 5240 871
rect 5234 866 5240 867
rect 5514 871 5520 872
rect 5514 867 5515 871
rect 5519 867 5520 871
rect 5514 866 5520 867
rect 5262 856 5268 857
rect 5262 852 5263 856
rect 5267 852 5268 856
rect 5262 851 5268 852
rect 5542 856 5548 857
rect 5542 852 5543 856
rect 5547 852 5548 856
rect 5542 851 5548 852
rect 5264 827 5266 851
rect 5544 827 5546 851
rect 5087 826 5091 827
rect 5087 821 5091 822
rect 5263 826 5267 827
rect 5263 821 5267 822
rect 5287 826 5291 827
rect 5287 821 5291 822
rect 5487 826 5491 827
rect 5487 821 5491 822
rect 5543 826 5547 827
rect 5543 821 5547 822
rect 5088 797 5090 821
rect 5288 797 5290 821
rect 5488 797 5490 821
rect 5086 796 5092 797
rect 5086 792 5087 796
rect 5091 792 5092 796
rect 5086 791 5092 792
rect 5286 796 5292 797
rect 5286 792 5287 796
rect 5291 792 5292 796
rect 5286 791 5292 792
rect 5486 796 5492 797
rect 5486 792 5487 796
rect 5491 792 5492 796
rect 5486 791 5492 792
rect 5258 781 5264 782
rect 5258 777 5259 781
rect 5263 777 5264 781
rect 5258 776 5264 777
rect 5458 781 5464 782
rect 5458 777 5459 781
rect 5463 777 5464 781
rect 5458 776 5464 777
rect 5218 771 5224 772
rect 5218 767 5219 771
rect 5223 767 5224 771
rect 5218 766 5224 767
rect 5220 732 5222 766
rect 5066 731 5072 732
rect 5066 727 5067 731
rect 5071 727 5072 731
rect 5066 726 5072 727
rect 5218 731 5224 732
rect 5218 727 5219 731
rect 5223 727 5224 731
rect 5218 726 5224 727
rect 5260 711 5262 776
rect 5460 711 5462 776
rect 5556 772 5558 954
rect 5612 924 5614 1106
rect 5664 1105 5666 1165
rect 5662 1104 5668 1105
rect 5662 1100 5663 1104
rect 5667 1100 5668 1104
rect 5662 1099 5668 1100
rect 5662 1087 5668 1088
rect 5662 1083 5663 1087
rect 5667 1083 5668 1087
rect 5662 1082 5668 1083
rect 5664 1055 5666 1082
rect 5663 1054 5667 1055
rect 5663 1049 5667 1050
rect 5664 1026 5666 1049
rect 5662 1025 5668 1026
rect 5662 1021 5663 1025
rect 5667 1021 5668 1025
rect 5662 1020 5668 1021
rect 5662 1008 5668 1009
rect 5662 1004 5663 1008
rect 5667 1004 5668 1008
rect 5662 1003 5668 1004
rect 5664 939 5666 1003
rect 5663 938 5667 939
rect 5663 933 5667 934
rect 5610 923 5616 924
rect 5610 919 5611 923
rect 5615 919 5616 923
rect 5610 918 5616 919
rect 5610 879 5616 880
rect 5610 875 5611 879
rect 5615 875 5616 879
rect 5610 874 5616 875
rect 5554 771 5560 772
rect 5554 767 5555 771
rect 5559 767 5560 771
rect 5554 766 5560 767
rect 5554 731 5560 732
rect 5554 727 5555 731
rect 5559 727 5560 731
rect 5554 726 5560 727
rect 4691 710 4695 711
rect 4691 705 4695 706
rect 4699 710 4703 711
rect 4699 705 4703 706
rect 4867 710 4871 711
rect 4867 705 4871 706
rect 4891 710 4895 711
rect 4891 705 4895 706
rect 5059 710 5063 711
rect 5059 705 5063 706
rect 5099 710 5103 711
rect 5099 705 5103 706
rect 5259 710 5263 711
rect 5259 705 5263 706
rect 5315 710 5319 711
rect 5315 705 5319 706
rect 5459 710 5463 711
rect 5459 705 5463 706
rect 5515 710 5519 711
rect 5515 705 5519 706
rect 4634 695 4640 696
rect 4634 691 4635 695
rect 4639 691 4640 695
rect 4634 690 4640 691
rect 4700 644 4702 705
rect 4706 691 4712 692
rect 4706 687 4707 691
rect 4711 687 4712 691
rect 4706 686 4712 687
rect 4708 652 4710 686
rect 4706 651 4712 652
rect 4706 647 4707 651
rect 4711 647 4712 651
rect 4706 646 4712 647
rect 4892 644 4894 705
rect 4898 691 4904 692
rect 4898 687 4899 691
rect 4903 687 4904 691
rect 4898 686 4904 687
rect 4900 652 4902 686
rect 4898 651 4904 652
rect 4898 647 4899 651
rect 4903 647 4904 651
rect 4898 646 4904 647
rect 5100 644 5102 705
rect 5106 691 5112 692
rect 5106 687 5107 691
rect 5111 687 5112 691
rect 5106 686 5112 687
rect 5108 652 5110 686
rect 5106 651 5112 652
rect 5106 647 5107 651
rect 5111 647 5112 651
rect 5106 646 5112 647
rect 5316 644 5318 705
rect 5322 691 5328 692
rect 5322 687 5323 691
rect 5327 687 5328 691
rect 5322 686 5328 687
rect 5324 652 5326 686
rect 5322 651 5328 652
rect 5322 647 5323 651
rect 5327 647 5328 651
rect 5322 646 5328 647
rect 5366 651 5372 652
rect 5366 647 5367 651
rect 5371 647 5372 651
rect 5366 646 5372 647
rect 4130 643 4136 644
rect 4130 639 4131 643
rect 4135 639 4136 643
rect 4130 638 4136 639
rect 4266 643 4272 644
rect 4266 639 4267 643
rect 4271 639 4272 643
rect 4266 638 4272 639
rect 4402 643 4408 644
rect 4402 639 4403 643
rect 4407 639 4408 643
rect 4402 638 4408 639
rect 4538 643 4544 644
rect 4538 639 4539 643
rect 4543 639 4544 643
rect 4538 638 4544 639
rect 4698 643 4704 644
rect 4698 639 4699 643
rect 4703 639 4704 643
rect 4698 638 4704 639
rect 4890 643 4896 644
rect 4890 639 4891 643
rect 4895 639 4896 643
rect 4890 638 4896 639
rect 5098 643 5104 644
rect 5098 639 5099 643
rect 5103 639 5104 643
rect 5098 638 5104 639
rect 5314 643 5320 644
rect 5314 639 5315 643
rect 5319 639 5320 643
rect 5314 638 5320 639
rect 4022 628 4028 629
rect 4022 624 4023 628
rect 4027 624 4028 628
rect 4022 623 4028 624
rect 4158 628 4164 629
rect 4158 624 4159 628
rect 4163 624 4164 628
rect 4158 623 4164 624
rect 4294 628 4300 629
rect 4294 624 4295 628
rect 4299 624 4300 628
rect 4294 623 4300 624
rect 4430 628 4436 629
rect 4430 624 4431 628
rect 4435 624 4436 628
rect 4430 623 4436 624
rect 4566 628 4572 629
rect 4566 624 4567 628
rect 4571 624 4572 628
rect 4566 623 4572 624
rect 4726 628 4732 629
rect 4726 624 4727 628
rect 4731 624 4732 628
rect 4726 623 4732 624
rect 4918 628 4924 629
rect 4918 624 4919 628
rect 4923 624 4924 628
rect 4918 623 4924 624
rect 5126 628 5132 629
rect 5126 624 5127 628
rect 5131 624 5132 628
rect 5126 623 5132 624
rect 5342 628 5348 629
rect 5342 624 5343 628
rect 5347 624 5348 628
rect 5342 623 5348 624
rect 4024 599 4026 623
rect 4160 599 4162 623
rect 4296 599 4298 623
rect 4432 599 4434 623
rect 4568 599 4570 623
rect 4728 599 4730 623
rect 4920 599 4922 623
rect 5128 599 5130 623
rect 5344 599 5346 623
rect 4023 598 4027 599
rect 4023 593 4027 594
rect 4071 598 4075 599
rect 4071 593 4075 594
rect 4159 598 4163 599
rect 4159 593 4163 594
rect 4295 598 4299 599
rect 4295 593 4299 594
rect 4311 598 4315 599
rect 4311 593 4315 594
rect 4431 598 4435 599
rect 4431 593 4435 594
rect 4567 598 4571 599
rect 4567 593 4571 594
rect 4575 598 4579 599
rect 4575 593 4579 594
rect 4727 598 4731 599
rect 4727 593 4731 594
rect 4855 598 4859 599
rect 4855 593 4859 594
rect 4919 598 4923 599
rect 4919 593 4923 594
rect 5127 598 5131 599
rect 5127 593 5131 594
rect 5151 598 5155 599
rect 5151 593 5155 594
rect 5343 598 5347 599
rect 5343 593 5347 594
rect 4072 569 4074 593
rect 4312 569 4314 593
rect 4576 569 4578 593
rect 4856 569 4858 593
rect 5152 569 5154 593
rect 4070 568 4076 569
rect 4070 564 4071 568
rect 4075 564 4076 568
rect 4070 563 4076 564
rect 4310 568 4316 569
rect 4310 564 4311 568
rect 4315 564 4316 568
rect 4310 563 4316 564
rect 4574 568 4580 569
rect 4574 564 4575 568
rect 4579 564 4580 568
rect 4574 563 4580 564
rect 4854 568 4860 569
rect 4854 564 4855 568
rect 4859 564 4860 568
rect 4854 563 4860 564
rect 5150 568 5156 569
rect 5150 564 5151 568
rect 5155 564 5156 568
rect 5150 563 5156 564
rect 4042 553 4048 554
rect 4042 549 4043 553
rect 4047 549 4048 553
rect 4042 548 4048 549
rect 4282 553 4288 554
rect 4282 549 4283 553
rect 4287 549 4288 553
rect 4282 548 4288 549
rect 4546 553 4552 554
rect 4546 549 4547 553
rect 4551 549 4552 553
rect 4546 548 4552 549
rect 4826 553 4832 554
rect 4826 549 4827 553
rect 4831 549 4832 553
rect 4826 548 4832 549
rect 5122 553 5128 554
rect 5122 549 5123 553
rect 5127 549 5128 553
rect 5122 548 5128 549
rect 4002 543 4008 544
rect 4002 539 4003 543
rect 4007 539 4008 543
rect 4002 538 4008 539
rect 4044 475 4046 548
rect 4170 543 4176 544
rect 4170 539 4171 543
rect 4175 539 4176 543
rect 4170 538 4176 539
rect 4172 504 4174 538
rect 4170 503 4176 504
rect 4170 499 4171 503
rect 4175 499 4176 503
rect 4170 498 4176 499
rect 4284 475 4286 548
rect 4548 475 4550 548
rect 4674 543 4680 544
rect 4674 539 4675 543
rect 4679 539 4680 543
rect 4674 538 4680 539
rect 4634 535 4640 536
rect 4634 531 4635 535
rect 4639 531 4640 535
rect 4634 530 4640 531
rect 3839 474 3843 475
rect 3839 469 3843 470
rect 3859 474 3863 475
rect 3859 469 3863 470
rect 4043 474 4047 475
rect 4043 469 4047 470
rect 4283 474 4287 475
rect 4283 469 4287 470
rect 4451 474 4455 475
rect 4451 469 4455 470
rect 4547 474 4551 475
rect 4547 469 4551 470
rect 3243 466 3247 467
rect 3243 461 3247 462
rect 3267 466 3271 467
rect 3267 461 3271 462
rect 3379 466 3383 467
rect 3379 461 3383 462
rect 3467 466 3471 467
rect 3467 461 3471 462
rect 3515 466 3519 467
rect 3515 461 3519 462
rect 3651 466 3655 467
rect 3651 461 3655 462
rect 3799 466 3803 467
rect 3799 461 3803 462
rect 3202 415 3208 416
rect 3202 411 3203 415
rect 3207 411 3208 415
rect 3202 410 3208 411
rect 3074 407 3080 408
rect 3074 403 3075 407
rect 3079 403 3080 407
rect 3074 402 3080 403
rect 3268 400 3270 461
rect 3274 447 3280 448
rect 3274 443 3275 447
rect 3279 443 3280 447
rect 3274 442 3280 443
rect 3276 408 3278 442
rect 3274 407 3280 408
rect 3274 403 3275 407
rect 3279 403 3280 407
rect 3274 402 3280 403
rect 3468 400 3470 461
rect 3634 451 3640 452
rect 3474 447 3480 448
rect 3474 443 3475 447
rect 3479 443 3480 447
rect 3634 447 3635 451
rect 3639 447 3640 451
rect 3634 446 3640 447
rect 3474 442 3480 443
rect 3476 408 3478 442
rect 3474 407 3480 408
rect 3474 403 3475 407
rect 3479 403 3480 407
rect 3636 404 3638 446
rect 3474 402 3480 403
rect 3634 403 3640 404
rect 3066 399 3072 400
rect 3066 395 3067 399
rect 3071 395 3072 399
rect 3066 394 3072 395
rect 3266 399 3272 400
rect 3266 395 3267 399
rect 3271 395 3272 399
rect 3266 394 3272 395
rect 3466 399 3472 400
rect 3466 395 3467 399
rect 3471 395 3472 399
rect 3634 399 3635 403
rect 3639 399 3640 403
rect 3652 400 3654 461
rect 3800 401 3802 461
rect 3840 409 3842 469
rect 3838 408 3844 409
rect 4452 408 4454 469
rect 4636 460 4638 530
rect 4676 504 4678 538
rect 4674 503 4680 504
rect 4674 499 4675 503
rect 4679 499 4680 503
rect 4674 498 4680 499
rect 4828 475 4830 548
rect 5124 475 5126 548
rect 5368 488 5370 646
rect 5516 644 5518 705
rect 5556 652 5558 726
rect 5612 696 5614 874
rect 5664 873 5666 933
rect 5662 872 5668 873
rect 5662 868 5663 872
rect 5667 868 5668 872
rect 5662 867 5668 868
rect 5662 855 5668 856
rect 5662 851 5663 855
rect 5667 851 5668 855
rect 5662 850 5668 851
rect 5664 827 5666 850
rect 5663 826 5667 827
rect 5663 821 5667 822
rect 5664 798 5666 821
rect 5662 797 5668 798
rect 5662 793 5663 797
rect 5667 793 5668 797
rect 5662 792 5668 793
rect 5662 780 5668 781
rect 5662 776 5663 780
rect 5667 776 5668 780
rect 5662 775 5668 776
rect 5664 711 5666 775
rect 5663 710 5667 711
rect 5663 705 5667 706
rect 5610 695 5616 696
rect 5610 691 5611 695
rect 5615 691 5616 695
rect 5610 690 5616 691
rect 5554 651 5560 652
rect 5554 647 5555 651
rect 5559 647 5560 651
rect 5554 646 5560 647
rect 5664 645 5666 705
rect 5662 644 5668 645
rect 5514 643 5520 644
rect 5514 639 5515 643
rect 5519 639 5520 643
rect 5662 640 5663 644
rect 5667 640 5668 644
rect 5662 639 5668 640
rect 5514 638 5520 639
rect 5542 628 5548 629
rect 5542 624 5543 628
rect 5547 624 5548 628
rect 5542 623 5548 624
rect 5662 627 5668 628
rect 5662 623 5663 627
rect 5667 623 5668 627
rect 5544 599 5546 623
rect 5662 622 5668 623
rect 5664 599 5666 622
rect 5447 598 5451 599
rect 5447 593 5451 594
rect 5543 598 5547 599
rect 5543 593 5547 594
rect 5663 598 5667 599
rect 5663 593 5667 594
rect 5448 569 5450 593
rect 5664 570 5666 593
rect 5662 569 5668 570
rect 5446 568 5452 569
rect 5446 564 5447 568
rect 5451 564 5452 568
rect 5662 565 5663 569
rect 5667 565 5668 569
rect 5662 564 5668 565
rect 5446 563 5452 564
rect 5418 553 5424 554
rect 5418 549 5419 553
rect 5423 549 5424 553
rect 5418 548 5424 549
rect 5662 552 5668 553
rect 5662 548 5663 552
rect 5667 548 5668 552
rect 5394 503 5400 504
rect 5394 499 5395 503
rect 5399 499 5400 503
rect 5394 498 5400 499
rect 5366 487 5372 488
rect 5366 483 5367 487
rect 5371 483 5372 487
rect 5366 482 5372 483
rect 4643 474 4647 475
rect 4643 469 4647 470
rect 4827 474 4831 475
rect 4827 469 4831 470
rect 4843 474 4847 475
rect 4843 469 4847 470
rect 5051 474 5055 475
rect 5051 469 5055 470
rect 5123 474 5127 475
rect 5123 469 5127 470
rect 5267 474 5271 475
rect 5267 469 5271 470
rect 4634 459 4640 460
rect 4634 455 4635 459
rect 4639 455 4640 459
rect 4634 454 4640 455
rect 4644 408 4646 469
rect 4650 455 4656 456
rect 4650 451 4651 455
rect 4655 451 4656 455
rect 4650 450 4656 451
rect 4652 416 4654 450
rect 4650 415 4656 416
rect 4650 411 4651 415
rect 4655 411 4656 415
rect 4650 410 4656 411
rect 4844 408 4846 469
rect 4850 455 4856 456
rect 4850 451 4851 455
rect 4855 451 4856 455
rect 4850 450 4856 451
rect 4852 416 4854 450
rect 4850 415 4856 416
rect 4850 411 4851 415
rect 4855 411 4856 415
rect 4850 410 4856 411
rect 5052 408 5054 469
rect 5058 455 5064 456
rect 5058 451 5059 455
rect 5063 451 5064 455
rect 5058 450 5064 451
rect 5060 416 5062 450
rect 5058 415 5064 416
rect 5058 411 5059 415
rect 5063 411 5064 415
rect 5058 410 5064 411
rect 5118 415 5124 416
rect 5118 411 5119 415
rect 5123 411 5124 415
rect 5118 410 5124 411
rect 3838 404 3839 408
rect 3843 404 3844 408
rect 3838 403 3844 404
rect 4450 407 4456 408
rect 4450 403 4451 407
rect 4455 403 4456 407
rect 4450 402 4456 403
rect 4642 407 4648 408
rect 4642 403 4643 407
rect 4647 403 4648 407
rect 4642 402 4648 403
rect 4842 407 4848 408
rect 4842 403 4843 407
rect 4847 403 4848 407
rect 4842 402 4848 403
rect 5050 407 5056 408
rect 5050 403 5051 407
rect 5055 403 5056 407
rect 5050 402 5056 403
rect 3798 400 3804 401
rect 3634 398 3640 399
rect 3650 399 3656 400
rect 3466 394 3472 395
rect 3650 395 3651 399
rect 3655 395 3656 399
rect 3798 396 3799 400
rect 3803 396 3804 400
rect 3798 395 3804 396
rect 3650 394 3656 395
rect 4478 392 4484 393
rect 3838 391 3844 392
rect 3838 387 3839 391
rect 3843 387 3844 391
rect 4478 388 4479 392
rect 4483 388 4484 392
rect 4478 387 4484 388
rect 4670 392 4676 393
rect 4670 388 4671 392
rect 4675 388 4676 392
rect 4670 387 4676 388
rect 4870 392 4876 393
rect 4870 388 4871 392
rect 4875 388 4876 392
rect 4870 387 4876 388
rect 5078 392 5084 393
rect 5078 388 5079 392
rect 5083 388 5084 392
rect 5078 387 5084 388
rect 3838 386 3844 387
rect 3094 384 3100 385
rect 3094 380 3095 384
rect 3099 380 3100 384
rect 3094 379 3100 380
rect 3294 384 3300 385
rect 3294 380 3295 384
rect 3299 380 3300 384
rect 3294 379 3300 380
rect 3494 384 3500 385
rect 3494 380 3495 384
rect 3499 380 3500 384
rect 3494 379 3500 380
rect 3678 384 3684 385
rect 3678 380 3679 384
rect 3683 380 3684 384
rect 3678 379 3684 380
rect 3798 383 3804 384
rect 3798 379 3799 383
rect 3803 379 3804 383
rect 3096 339 3098 379
rect 3296 339 3298 379
rect 3496 339 3498 379
rect 3680 339 3682 379
rect 3798 378 3804 379
rect 3800 339 3802 378
rect 3840 359 3842 386
rect 4480 359 4482 387
rect 4672 359 4674 387
rect 4872 359 4874 387
rect 5080 359 5082 387
rect 3839 358 3843 359
rect 3839 353 3843 354
rect 4479 358 4483 359
rect 4479 353 4483 354
rect 4615 358 4619 359
rect 4615 353 4619 354
rect 4671 358 4675 359
rect 4671 353 4675 354
rect 4775 358 4779 359
rect 4775 353 4779 354
rect 4871 358 4875 359
rect 4871 353 4875 354
rect 4951 358 4955 359
rect 4951 353 4955 354
rect 5079 358 5083 359
rect 5079 353 5083 354
rect 2975 338 2979 339
rect 2975 333 2979 334
rect 3095 338 3099 339
rect 3095 333 3099 334
rect 3111 338 3115 339
rect 3111 333 3115 334
rect 3247 338 3251 339
rect 3247 333 3251 334
rect 3295 338 3299 339
rect 3295 333 3299 334
rect 3383 338 3387 339
rect 3383 333 3387 334
rect 3495 338 3499 339
rect 3495 333 3499 334
rect 3519 338 3523 339
rect 3519 333 3523 334
rect 3655 338 3659 339
rect 3655 333 3659 334
rect 3679 338 3683 339
rect 3679 333 3683 334
rect 3799 338 3803 339
rect 3799 333 3803 334
rect 2976 309 2978 333
rect 3112 309 3114 333
rect 3248 309 3250 333
rect 3384 309 3386 333
rect 3520 309 3522 333
rect 3656 309 3658 333
rect 3800 310 3802 333
rect 3840 330 3842 353
rect 3838 329 3844 330
rect 4616 329 4618 353
rect 4776 329 4778 353
rect 4952 329 4954 353
rect 3838 325 3839 329
rect 3843 325 3844 329
rect 3838 324 3844 325
rect 4614 328 4620 329
rect 4614 324 4615 328
rect 4619 324 4620 328
rect 4614 323 4620 324
rect 4774 328 4780 329
rect 4774 324 4775 328
rect 4779 324 4780 328
rect 4774 323 4780 324
rect 4950 328 4956 329
rect 4950 324 4951 328
rect 4955 324 4956 328
rect 4950 323 4956 324
rect 4586 313 4592 314
rect 3838 312 3844 313
rect 3798 309 3804 310
rect 2974 308 2980 309
rect 2974 304 2975 308
rect 2979 304 2980 308
rect 2974 303 2980 304
rect 3110 308 3116 309
rect 3110 304 3111 308
rect 3115 304 3116 308
rect 3110 303 3116 304
rect 3246 308 3252 309
rect 3246 304 3247 308
rect 3251 304 3252 308
rect 3246 303 3252 304
rect 3382 308 3388 309
rect 3382 304 3383 308
rect 3387 304 3388 308
rect 3382 303 3388 304
rect 3518 308 3524 309
rect 3518 304 3519 308
rect 3523 304 3524 308
rect 3518 303 3524 304
rect 3654 308 3660 309
rect 3654 304 3655 308
rect 3659 304 3660 308
rect 3798 305 3799 309
rect 3803 305 3804 309
rect 3838 308 3839 312
rect 3843 308 3844 312
rect 4586 309 4587 313
rect 4591 309 4592 313
rect 4586 308 4592 309
rect 4746 313 4752 314
rect 4746 309 4747 313
rect 4751 309 4752 313
rect 4746 308 4752 309
rect 4922 313 4928 314
rect 4922 309 4923 313
rect 4927 309 4928 313
rect 4922 308 4928 309
rect 5106 313 5112 314
rect 5106 309 5107 313
rect 5111 309 5112 313
rect 5106 308 5112 309
rect 3838 307 3844 308
rect 3798 304 3804 305
rect 3654 303 3660 304
rect 3082 293 3088 294
rect 3082 289 3083 293
rect 3087 289 3088 293
rect 3082 288 3088 289
rect 3218 293 3224 294
rect 3218 289 3219 293
rect 3223 289 3224 293
rect 3218 288 3224 289
rect 3354 293 3360 294
rect 3354 289 3355 293
rect 3359 289 3360 293
rect 3354 288 3360 289
rect 3490 293 3496 294
rect 3490 289 3491 293
rect 3495 289 3496 293
rect 3490 288 3496 289
rect 3626 293 3632 294
rect 3626 289 3627 293
rect 3631 289 3632 293
rect 3626 288 3632 289
rect 3798 292 3804 293
rect 3798 288 3799 292
rect 3803 288 3804 292
rect 3074 283 3080 284
rect 3074 279 3075 283
rect 3079 279 3080 283
rect 3074 278 3080 279
rect 2954 267 2960 268
rect 2954 263 2955 267
rect 2959 263 2960 267
rect 2954 262 2960 263
rect 3076 244 3078 278
rect 3042 243 3048 244
rect 3042 239 3043 243
rect 3047 239 3048 243
rect 3042 238 3048 239
rect 3074 243 3080 244
rect 3074 239 3075 243
rect 3079 239 3080 243
rect 3074 238 3080 239
rect 2131 190 2135 191
rect 2131 185 2135 186
rect 2267 190 2271 191
rect 2267 185 2271 186
rect 2403 190 2407 191
rect 2403 185 2407 186
rect 2539 190 2543 191
rect 2539 185 2543 186
rect 2675 190 2679 191
rect 2675 185 2679 186
rect 2811 190 2815 191
rect 2811 185 2815 186
rect 2947 190 2951 191
rect 2947 185 2951 186
rect 2090 175 2096 176
rect 2090 171 2091 175
rect 2095 171 2096 175
rect 2090 170 2096 171
rect 2132 124 2134 185
rect 2138 171 2144 172
rect 2138 167 2139 171
rect 2143 167 2144 171
rect 2138 166 2144 167
rect 2140 132 2142 166
rect 2138 131 2144 132
rect 2138 127 2139 131
rect 2143 127 2144 131
rect 2138 126 2144 127
rect 2268 124 2270 185
rect 2274 171 2280 172
rect 2274 167 2275 171
rect 2279 167 2280 171
rect 2274 166 2280 167
rect 2276 132 2278 166
rect 2274 131 2280 132
rect 2274 127 2275 131
rect 2279 127 2280 131
rect 2274 126 2280 127
rect 2404 124 2406 185
rect 2410 171 2416 172
rect 2410 167 2411 171
rect 2415 167 2416 171
rect 2410 166 2416 167
rect 2412 132 2414 166
rect 2410 131 2416 132
rect 2410 127 2411 131
rect 2415 127 2416 131
rect 2410 126 2416 127
rect 2540 124 2542 185
rect 2546 171 2552 172
rect 2546 167 2547 171
rect 2551 167 2552 171
rect 2546 166 2552 167
rect 2548 132 2550 166
rect 2546 131 2552 132
rect 2546 127 2547 131
rect 2551 127 2552 131
rect 2546 126 2552 127
rect 2676 124 2678 185
rect 2682 171 2688 172
rect 2682 167 2683 171
rect 2687 167 2688 171
rect 2682 166 2688 167
rect 2684 132 2686 166
rect 2682 131 2688 132
rect 2682 127 2683 131
rect 2687 127 2688 131
rect 2682 126 2688 127
rect 2812 124 2814 185
rect 2818 171 2824 172
rect 2818 167 2819 171
rect 2823 167 2824 171
rect 2818 166 2824 167
rect 2820 132 2822 166
rect 2818 131 2824 132
rect 2818 127 2819 131
rect 2823 127 2824 131
rect 2818 126 2824 127
rect 2948 124 2950 185
rect 2954 171 2960 172
rect 2954 167 2955 171
rect 2959 167 2960 171
rect 2954 166 2960 167
rect 2956 132 2958 166
rect 3044 133 3046 238
rect 3084 191 3086 288
rect 3210 283 3216 284
rect 3210 279 3211 283
rect 3215 279 3216 283
rect 3210 278 3216 279
rect 3212 244 3214 278
rect 3210 243 3216 244
rect 3210 239 3211 243
rect 3215 239 3216 243
rect 3210 238 3216 239
rect 3220 191 3222 288
rect 3346 283 3352 284
rect 3346 279 3347 283
rect 3351 279 3352 283
rect 3346 278 3352 279
rect 3348 244 3350 278
rect 3346 243 3352 244
rect 3346 239 3347 243
rect 3351 239 3352 243
rect 3346 238 3352 239
rect 3356 191 3358 288
rect 3482 283 3488 284
rect 3482 279 3483 283
rect 3487 279 3488 283
rect 3482 278 3488 279
rect 3484 244 3486 278
rect 3482 243 3488 244
rect 3482 239 3483 243
rect 3487 239 3488 243
rect 3482 238 3488 239
rect 3492 191 3494 288
rect 3628 191 3630 288
rect 3798 287 3804 288
rect 3800 191 3802 287
rect 3840 207 3842 307
rect 4386 255 4392 256
rect 4386 251 4387 255
rect 4391 251 4392 255
rect 4386 250 4392 251
rect 3839 206 3843 207
rect 3839 201 3843 202
rect 4291 206 4295 207
rect 4291 201 4295 202
rect 3083 190 3087 191
rect 3083 185 3087 186
rect 3219 190 3223 191
rect 3219 185 3223 186
rect 3355 190 3359 191
rect 3355 185 3359 186
rect 3491 190 3495 191
rect 3491 185 3495 186
rect 3627 190 3631 191
rect 3627 185 3631 186
rect 3799 190 3803 191
rect 3799 185 3803 186
rect 3043 132 3047 133
rect 2954 131 2960 132
rect 2954 127 2955 131
rect 2959 127 2960 131
rect 3043 127 3047 128
rect 2954 126 2960 127
rect 3084 124 3086 185
rect 3090 171 3096 172
rect 3090 167 3091 171
rect 3095 167 3096 171
rect 3090 166 3096 167
rect 3092 132 3094 166
rect 3090 131 3096 132
rect 3090 127 3091 131
rect 3095 127 3096 131
rect 3090 126 3096 127
rect 3220 124 3222 185
rect 3226 171 3232 172
rect 3226 167 3227 171
rect 3231 167 3232 171
rect 3226 166 3232 167
rect 3228 132 3230 166
rect 3226 131 3232 132
rect 3226 127 3227 131
rect 3231 127 3232 131
rect 3226 126 3232 127
rect 3356 124 3358 185
rect 3362 171 3368 172
rect 3362 167 3363 171
rect 3367 167 3368 171
rect 3362 166 3368 167
rect 3364 132 3366 166
rect 3362 131 3368 132
rect 3362 127 3363 131
rect 3367 127 3368 131
rect 3362 126 3368 127
rect 3492 124 3494 185
rect 3498 171 3504 172
rect 3498 167 3499 171
rect 3503 167 3504 171
rect 3498 166 3504 167
rect 3500 132 3502 166
rect 3498 131 3504 132
rect 3498 127 3499 131
rect 3503 127 3504 131
rect 3498 126 3504 127
rect 3628 124 3630 185
rect 3634 171 3640 172
rect 3634 167 3635 171
rect 3639 167 3640 171
rect 3634 166 3640 167
rect 3636 132 3638 166
rect 3647 132 3651 133
rect 3634 131 3640 132
rect 3634 127 3635 131
rect 3639 127 3640 131
rect 3634 126 3640 127
rect 3646 127 3647 132
rect 3651 127 3652 132
rect 3646 126 3652 127
rect 3800 125 3802 185
rect 3840 141 3842 201
rect 3838 140 3844 141
rect 4292 140 4294 201
rect 4388 192 4390 250
rect 4588 207 4590 308
rect 4734 303 4740 304
rect 4734 299 4735 303
rect 4739 299 4740 303
rect 4734 298 4740 299
rect 4674 295 4680 296
rect 4674 291 4675 295
rect 4679 291 4680 295
rect 4674 290 4680 291
rect 4676 256 4678 290
rect 4736 264 4738 298
rect 4734 263 4740 264
rect 4734 259 4735 263
rect 4739 259 4740 263
rect 4734 258 4740 259
rect 4674 255 4680 256
rect 4674 251 4675 255
rect 4679 251 4680 255
rect 4674 250 4680 251
rect 4748 207 4750 308
rect 4874 303 4880 304
rect 4874 299 4875 303
rect 4879 299 4880 303
rect 4874 298 4880 299
rect 4876 264 4878 298
rect 4874 263 4880 264
rect 4874 259 4875 263
rect 4879 259 4880 263
rect 4874 258 4880 259
rect 4924 207 4926 308
rect 5050 303 5056 304
rect 5050 299 5051 303
rect 5055 299 5056 303
rect 5050 298 5056 299
rect 5052 264 5054 298
rect 5050 263 5056 264
rect 5050 259 5051 263
rect 5055 259 5056 263
rect 5050 258 5056 259
rect 5108 207 5110 308
rect 5120 256 5122 410
rect 5268 408 5270 469
rect 5362 455 5368 456
rect 5362 451 5363 455
rect 5367 451 5368 455
rect 5362 450 5368 451
rect 5266 407 5272 408
rect 5266 403 5267 407
rect 5271 403 5272 407
rect 5266 402 5272 403
rect 5294 392 5300 393
rect 5294 388 5295 392
rect 5299 388 5300 392
rect 5294 387 5300 388
rect 5296 359 5298 387
rect 5135 358 5139 359
rect 5135 353 5139 354
rect 5295 358 5299 359
rect 5295 353 5299 354
rect 5327 358 5331 359
rect 5327 353 5331 354
rect 5136 329 5138 353
rect 5328 329 5330 353
rect 5134 328 5140 329
rect 5134 324 5135 328
rect 5139 324 5140 328
rect 5134 323 5140 324
rect 5326 328 5332 329
rect 5326 324 5327 328
rect 5331 324 5332 328
rect 5326 323 5332 324
rect 5298 313 5304 314
rect 5298 309 5299 313
rect 5303 309 5304 313
rect 5298 308 5304 309
rect 5118 255 5124 256
rect 5118 251 5119 255
rect 5123 251 5124 255
rect 5118 250 5124 251
rect 5300 207 5302 308
rect 4427 206 4431 207
rect 4427 201 4431 202
rect 4563 206 4567 207
rect 4563 201 4567 202
rect 4587 206 4591 207
rect 4587 201 4591 202
rect 4699 206 4703 207
rect 4699 201 4703 202
rect 4747 206 4751 207
rect 4747 201 4751 202
rect 4835 206 4839 207
rect 4835 201 4839 202
rect 4923 206 4927 207
rect 4923 201 4927 202
rect 4971 206 4975 207
rect 4971 201 4975 202
rect 5107 206 5111 207
rect 5107 201 5111 202
rect 5243 206 5247 207
rect 5243 201 5247 202
rect 5299 206 5303 207
rect 5299 201 5303 202
rect 4386 191 4392 192
rect 4386 187 4387 191
rect 4391 187 4392 191
rect 4386 186 4392 187
rect 4428 140 4430 201
rect 4434 187 4440 188
rect 4434 183 4435 187
rect 4439 183 4440 187
rect 4434 182 4440 183
rect 4436 148 4438 182
rect 4434 147 4440 148
rect 4434 143 4435 147
rect 4439 143 4440 147
rect 4434 142 4440 143
rect 4564 140 4566 201
rect 4570 187 4576 188
rect 4570 183 4571 187
rect 4575 183 4576 187
rect 4570 182 4576 183
rect 4572 148 4574 182
rect 4570 147 4576 148
rect 4570 143 4571 147
rect 4575 143 4576 147
rect 4570 142 4576 143
rect 4700 140 4702 201
rect 4706 187 4712 188
rect 4706 183 4707 187
rect 4711 183 4712 187
rect 4706 182 4712 183
rect 4708 148 4710 182
rect 4706 147 4712 148
rect 4706 143 4707 147
rect 4711 143 4712 147
rect 4706 142 4712 143
rect 4836 140 4838 201
rect 4842 187 4848 188
rect 4842 183 4843 187
rect 4847 183 4848 187
rect 4842 182 4848 183
rect 4844 148 4846 182
rect 4842 147 4848 148
rect 4842 143 4843 147
rect 4847 143 4848 147
rect 4842 142 4848 143
rect 4972 140 4974 201
rect 4978 187 4984 188
rect 4978 183 4979 187
rect 4983 183 4984 187
rect 4978 182 4984 183
rect 4980 148 4982 182
rect 4978 147 4984 148
rect 4978 143 4979 147
rect 4983 143 4984 147
rect 4978 142 4984 143
rect 5108 140 5110 201
rect 5114 187 5120 188
rect 5114 183 5115 187
rect 5119 183 5120 187
rect 5114 182 5120 183
rect 5116 148 5118 182
rect 5114 147 5120 148
rect 5114 143 5115 147
rect 5119 143 5120 147
rect 5114 142 5120 143
rect 5244 140 5246 201
rect 5250 187 5256 188
rect 5250 183 5251 187
rect 5255 183 5256 187
rect 5250 182 5256 183
rect 5252 148 5254 182
rect 5364 148 5366 450
rect 5396 416 5398 498
rect 5420 475 5422 548
rect 5662 547 5668 548
rect 5542 543 5548 544
rect 5542 539 5543 543
rect 5547 539 5548 543
rect 5542 538 5548 539
rect 5419 474 5423 475
rect 5419 469 5423 470
rect 5483 474 5487 475
rect 5483 469 5487 470
rect 5394 415 5400 416
rect 5394 411 5395 415
rect 5399 411 5400 415
rect 5394 410 5400 411
rect 5484 408 5486 469
rect 5544 460 5546 538
rect 5664 475 5666 547
rect 5663 474 5667 475
rect 5663 469 5667 470
rect 5542 459 5548 460
rect 5542 455 5543 459
rect 5547 455 5548 459
rect 5542 454 5548 455
rect 5594 415 5600 416
rect 5594 411 5595 415
rect 5599 411 5600 415
rect 5594 410 5600 411
rect 5482 407 5488 408
rect 5482 403 5483 407
rect 5487 403 5488 407
rect 5482 402 5488 403
rect 5510 392 5516 393
rect 5510 388 5511 392
rect 5515 388 5516 392
rect 5510 387 5516 388
rect 5512 359 5514 387
rect 5511 358 5515 359
rect 5511 353 5515 354
rect 5527 358 5531 359
rect 5527 353 5531 354
rect 5528 329 5530 353
rect 5526 328 5532 329
rect 5526 324 5527 328
rect 5531 324 5532 328
rect 5526 323 5532 324
rect 5498 313 5504 314
rect 5498 309 5499 313
rect 5503 309 5504 313
rect 5498 308 5504 309
rect 5500 207 5502 308
rect 5596 264 5598 410
rect 5664 409 5666 469
rect 5662 408 5668 409
rect 5662 404 5663 408
rect 5667 404 5668 408
rect 5662 403 5668 404
rect 5662 391 5668 392
rect 5662 387 5663 391
rect 5667 387 5668 391
rect 5662 386 5668 387
rect 5664 359 5666 386
rect 5663 358 5667 359
rect 5663 353 5667 354
rect 5664 330 5666 353
rect 5662 329 5668 330
rect 5662 325 5663 329
rect 5667 325 5668 329
rect 5662 324 5668 325
rect 5662 312 5668 313
rect 5662 308 5663 312
rect 5667 308 5668 312
rect 5662 307 5668 308
rect 5610 303 5616 304
rect 5610 299 5611 303
rect 5615 299 5616 303
rect 5610 298 5616 299
rect 5594 263 5600 264
rect 5594 259 5595 263
rect 5599 259 5600 263
rect 5594 258 5600 259
rect 5379 206 5383 207
rect 5379 201 5383 202
rect 5499 206 5503 207
rect 5499 201 5503 202
rect 5515 206 5519 207
rect 5515 201 5519 202
rect 5250 147 5256 148
rect 5250 143 5251 147
rect 5255 143 5256 147
rect 5250 142 5256 143
rect 5362 147 5368 148
rect 5362 143 5363 147
rect 5367 143 5368 147
rect 5362 142 5368 143
rect 5380 140 5382 201
rect 5474 187 5480 188
rect 5474 183 5475 187
rect 5479 183 5480 187
rect 5474 182 5480 183
rect 5476 148 5478 182
rect 5474 147 5480 148
rect 5474 143 5475 147
rect 5479 143 5480 147
rect 5474 142 5480 143
rect 5516 140 5518 201
rect 5612 192 5614 298
rect 5664 207 5666 307
rect 5663 206 5667 207
rect 5663 201 5667 202
rect 5610 191 5616 192
rect 5610 187 5611 191
rect 5615 187 5616 191
rect 5610 186 5616 187
rect 5664 141 5666 201
rect 5662 140 5668 141
rect 3838 136 3839 140
rect 3843 136 3844 140
rect 3838 135 3844 136
rect 4290 139 4296 140
rect 4290 135 4291 139
rect 4295 135 4296 139
rect 4290 134 4296 135
rect 4426 139 4432 140
rect 4426 135 4427 139
rect 4431 135 4432 139
rect 4426 134 4432 135
rect 4562 139 4568 140
rect 4562 135 4563 139
rect 4567 135 4568 139
rect 4562 134 4568 135
rect 4698 139 4704 140
rect 4698 135 4699 139
rect 4703 135 4704 139
rect 4698 134 4704 135
rect 4834 139 4840 140
rect 4834 135 4835 139
rect 4839 135 4840 139
rect 4834 134 4840 135
rect 4970 139 4976 140
rect 4970 135 4971 139
rect 4975 135 4976 139
rect 4970 134 4976 135
rect 5106 139 5112 140
rect 5106 135 5107 139
rect 5111 135 5112 139
rect 5106 134 5112 135
rect 5242 139 5248 140
rect 5242 135 5243 139
rect 5247 135 5248 139
rect 5242 134 5248 135
rect 5378 139 5384 140
rect 5378 135 5379 139
rect 5383 135 5384 139
rect 5378 134 5384 135
rect 5514 139 5520 140
rect 5514 135 5515 139
rect 5519 135 5520 139
rect 5662 136 5663 140
rect 5667 136 5668 140
rect 5662 135 5668 136
rect 5514 134 5520 135
rect 3798 124 3804 125
rect 4318 124 4324 125
rect 1936 99 1938 122
rect 1974 120 1975 124
rect 1979 120 1980 124
rect 1974 119 1980 120
rect 1994 123 2000 124
rect 1994 119 1995 123
rect 1999 119 2000 123
rect 1994 118 2000 119
rect 2130 123 2136 124
rect 2130 119 2131 123
rect 2135 119 2136 123
rect 2130 118 2136 119
rect 2266 123 2272 124
rect 2266 119 2267 123
rect 2271 119 2272 123
rect 2266 118 2272 119
rect 2402 123 2408 124
rect 2402 119 2403 123
rect 2407 119 2408 123
rect 2402 118 2408 119
rect 2538 123 2544 124
rect 2538 119 2539 123
rect 2543 119 2544 123
rect 2538 118 2544 119
rect 2674 123 2680 124
rect 2674 119 2675 123
rect 2679 119 2680 123
rect 2674 118 2680 119
rect 2810 123 2816 124
rect 2810 119 2811 123
rect 2815 119 2816 123
rect 2810 118 2816 119
rect 2946 123 2952 124
rect 2946 119 2947 123
rect 2951 119 2952 123
rect 2946 118 2952 119
rect 3082 123 3088 124
rect 3082 119 3083 123
rect 3087 119 3088 123
rect 3082 118 3088 119
rect 3218 123 3224 124
rect 3218 119 3219 123
rect 3223 119 3224 123
rect 3218 118 3224 119
rect 3354 123 3360 124
rect 3354 119 3355 123
rect 3359 119 3360 123
rect 3354 118 3360 119
rect 3490 123 3496 124
rect 3490 119 3491 123
rect 3495 119 3496 123
rect 3490 118 3496 119
rect 3626 123 3632 124
rect 3626 119 3627 123
rect 3631 119 3632 123
rect 3798 120 3799 124
rect 3803 120 3804 124
rect 3798 119 3804 120
rect 3838 123 3844 124
rect 3838 119 3839 123
rect 3843 119 3844 123
rect 4318 120 4319 124
rect 4323 120 4324 124
rect 4318 119 4324 120
rect 4454 124 4460 125
rect 4454 120 4455 124
rect 4459 120 4460 124
rect 4454 119 4460 120
rect 4590 124 4596 125
rect 4590 120 4591 124
rect 4595 120 4596 124
rect 4590 119 4596 120
rect 4726 124 4732 125
rect 4726 120 4727 124
rect 4731 120 4732 124
rect 4726 119 4732 120
rect 4862 124 4868 125
rect 4862 120 4863 124
rect 4867 120 4868 124
rect 4862 119 4868 120
rect 4998 124 5004 125
rect 4998 120 4999 124
rect 5003 120 5004 124
rect 4998 119 5004 120
rect 5134 124 5140 125
rect 5134 120 5135 124
rect 5139 120 5140 124
rect 5134 119 5140 120
rect 5270 124 5276 125
rect 5270 120 5271 124
rect 5275 120 5276 124
rect 5270 119 5276 120
rect 5406 124 5412 125
rect 5406 120 5407 124
rect 5411 120 5412 124
rect 5406 119 5412 120
rect 5542 124 5548 125
rect 5542 120 5543 124
rect 5547 120 5548 124
rect 5542 119 5548 120
rect 5662 123 5668 124
rect 5662 119 5663 123
rect 5667 119 5668 123
rect 3626 118 3632 119
rect 3838 118 3844 119
rect 2022 108 2028 109
rect 1974 107 1980 108
rect 1974 103 1975 107
rect 1979 103 1980 107
rect 2022 104 2023 108
rect 2027 104 2028 108
rect 2022 103 2028 104
rect 2158 108 2164 109
rect 2158 104 2159 108
rect 2163 104 2164 108
rect 2158 103 2164 104
rect 2294 108 2300 109
rect 2294 104 2295 108
rect 2299 104 2300 108
rect 2294 103 2300 104
rect 2430 108 2436 109
rect 2430 104 2431 108
rect 2435 104 2436 108
rect 2430 103 2436 104
rect 2566 108 2572 109
rect 2566 104 2567 108
rect 2571 104 2572 108
rect 2566 103 2572 104
rect 2702 108 2708 109
rect 2702 104 2703 108
rect 2707 104 2708 108
rect 2702 103 2708 104
rect 2838 108 2844 109
rect 2838 104 2839 108
rect 2843 104 2844 108
rect 2838 103 2844 104
rect 2974 108 2980 109
rect 2974 104 2975 108
rect 2979 104 2980 108
rect 2974 103 2980 104
rect 3110 108 3116 109
rect 3110 104 3111 108
rect 3115 104 3116 108
rect 3110 103 3116 104
rect 3246 108 3252 109
rect 3246 104 3247 108
rect 3251 104 3252 108
rect 3246 103 3252 104
rect 3382 108 3388 109
rect 3382 104 3383 108
rect 3387 104 3388 108
rect 3382 103 3388 104
rect 3518 108 3524 109
rect 3518 104 3519 108
rect 3523 104 3524 108
rect 3518 103 3524 104
rect 3654 108 3660 109
rect 3654 104 3655 108
rect 3659 104 3660 108
rect 3654 103 3660 104
rect 3798 107 3804 108
rect 3798 103 3799 107
rect 3803 103 3804 107
rect 1974 102 1980 103
rect 111 98 115 99
rect 111 93 115 94
rect 159 98 163 99
rect 159 93 163 94
rect 295 98 299 99
rect 295 93 299 94
rect 431 98 435 99
rect 431 93 435 94
rect 567 98 571 99
rect 567 93 571 94
rect 703 98 707 99
rect 703 93 707 94
rect 839 98 843 99
rect 839 93 843 94
rect 975 98 979 99
rect 975 93 979 94
rect 1111 98 1115 99
rect 1111 93 1115 94
rect 1935 98 1939 99
rect 1935 93 1939 94
rect 1976 79 1978 102
rect 2024 79 2026 103
rect 2160 79 2162 103
rect 2296 79 2298 103
rect 2432 79 2434 103
rect 2568 79 2570 103
rect 2704 79 2706 103
rect 2840 79 2842 103
rect 2976 79 2978 103
rect 3112 79 3114 103
rect 3248 79 3250 103
rect 3384 79 3386 103
rect 3520 79 3522 103
rect 3656 79 3658 103
rect 3798 102 3804 103
rect 3800 79 3802 102
rect 3840 95 3842 118
rect 4320 95 4322 119
rect 4456 95 4458 119
rect 4592 95 4594 119
rect 4728 95 4730 119
rect 4864 95 4866 119
rect 5000 95 5002 119
rect 5136 95 5138 119
rect 5272 95 5274 119
rect 5408 95 5410 119
rect 5544 95 5546 119
rect 5662 118 5668 119
rect 5664 95 5666 118
rect 3839 94 3843 95
rect 3839 89 3843 90
rect 4319 94 4323 95
rect 4319 89 4323 90
rect 4455 94 4459 95
rect 4455 89 4459 90
rect 4591 94 4595 95
rect 4591 89 4595 90
rect 4727 94 4731 95
rect 4727 89 4731 90
rect 4863 94 4867 95
rect 4863 89 4867 90
rect 4999 94 5003 95
rect 4999 89 5003 90
rect 5135 94 5139 95
rect 5135 89 5139 90
rect 5271 94 5275 95
rect 5271 89 5275 90
rect 5407 94 5411 95
rect 5407 89 5411 90
rect 5543 94 5547 95
rect 5543 89 5547 90
rect 5663 94 5667 95
rect 5663 89 5667 90
rect 1975 78 1979 79
rect 1975 73 1979 74
rect 2023 78 2027 79
rect 2023 73 2027 74
rect 2159 78 2163 79
rect 2159 73 2163 74
rect 2295 78 2299 79
rect 2295 73 2299 74
rect 2431 78 2435 79
rect 2431 73 2435 74
rect 2567 78 2571 79
rect 2567 73 2571 74
rect 2703 78 2707 79
rect 2703 73 2707 74
rect 2839 78 2843 79
rect 2839 73 2843 74
rect 2975 78 2979 79
rect 2975 73 2979 74
rect 3111 78 3115 79
rect 3111 73 3115 74
rect 3247 78 3251 79
rect 3247 73 3251 74
rect 3383 78 3387 79
rect 3383 73 3387 74
rect 3519 78 3523 79
rect 3519 73 3523 74
rect 3655 78 3659 79
rect 3655 73 3659 74
rect 3799 78 3803 79
rect 3799 73 3803 74
<< m4c >>
rect 111 5754 115 5758
rect 159 5754 163 5758
rect 295 5754 299 5758
rect 1935 5754 1939 5758
rect 111 5642 115 5646
rect 131 5642 135 5646
rect 267 5642 271 5646
rect 275 5642 279 5646
rect 1975 5654 1979 5658
rect 2023 5654 2027 5658
rect 2183 5654 2187 5658
rect 2367 5654 2371 5658
rect 2551 5654 2555 5658
rect 2727 5654 2731 5658
rect 2895 5654 2899 5658
rect 3063 5654 3067 5658
rect 3223 5654 3227 5658
rect 3383 5654 3387 5658
rect 3543 5654 3547 5658
rect 3679 5654 3683 5658
rect 3799 5654 3803 5658
rect 475 5642 479 5646
rect 699 5642 703 5646
rect 955 5642 959 5646
rect 1227 5642 1231 5646
rect 1515 5642 1519 5646
rect 1787 5642 1791 5646
rect 1935 5642 1939 5646
rect 111 5530 115 5534
rect 159 5530 163 5534
rect 279 5530 283 5534
rect 303 5530 307 5534
rect 503 5530 507 5534
rect 519 5530 523 5534
rect 727 5530 731 5534
rect 767 5530 771 5534
rect 983 5530 987 5534
rect 1015 5530 1019 5534
rect 1255 5530 1259 5534
rect 1263 5530 1267 5534
rect 111 5418 115 5422
rect 251 5418 255 5422
rect 411 5418 415 5422
rect 491 5418 495 5422
rect 1511 5530 1515 5534
rect 1543 5530 1547 5534
rect 1767 5530 1771 5534
rect 611 5418 615 5422
rect 739 5418 743 5422
rect 819 5418 823 5422
rect 987 5418 991 5422
rect 1035 5418 1039 5422
rect 1235 5418 1239 5422
rect 1259 5418 1263 5422
rect 111 5306 115 5310
rect 439 5306 443 5310
rect 591 5306 595 5310
rect 639 5306 643 5310
rect 3839 5650 3843 5654
rect 4335 5650 4339 5654
rect 4471 5650 4475 5654
rect 4607 5650 4611 5654
rect 4743 5650 4747 5654
rect 4879 5650 4883 5654
rect 5015 5650 5019 5654
rect 5663 5650 5667 5654
rect 1975 5542 1979 5546
rect 1995 5542 1999 5546
rect 2139 5542 2143 5546
rect 2155 5542 2159 5546
rect 2339 5542 2343 5546
rect 2355 5542 2359 5546
rect 2523 5542 2527 5546
rect 2563 5542 2567 5546
rect 1815 5530 1819 5534
rect 1935 5530 1939 5534
rect 1483 5418 1487 5422
rect 1491 5418 1495 5422
rect 1739 5418 1743 5422
rect 1935 5418 1939 5422
rect 1975 5422 1979 5426
rect 2167 5422 2171 5426
rect 727 5306 731 5310
rect 847 5306 851 5310
rect 863 5306 867 5310
rect 999 5306 1003 5310
rect 1063 5306 1067 5310
rect 1135 5306 1139 5310
rect 1271 5306 1275 5310
rect 1287 5306 1291 5310
rect 1407 5306 1411 5310
rect 1519 5306 1523 5310
rect 1543 5306 1547 5310
rect 2699 5542 2703 5546
rect 2755 5542 2759 5546
rect 2867 5542 2871 5546
rect 2939 5542 2943 5546
rect 3035 5542 3039 5546
rect 3115 5542 3119 5546
rect 3195 5542 3199 5546
rect 3291 5542 3295 5546
rect 3355 5542 3359 5546
rect 3467 5542 3471 5546
rect 3515 5542 3519 5546
rect 3643 5542 3647 5546
rect 3651 5542 3655 5546
rect 2311 5422 2315 5426
rect 2383 5422 2387 5426
rect 2511 5422 2515 5426
rect 2591 5422 2595 5426
rect 2703 5422 2707 5426
rect 2783 5422 2787 5426
rect 2887 5422 2891 5426
rect 2967 5422 2971 5426
rect 3071 5422 3075 5426
rect 3143 5422 3147 5426
rect 1935 5306 1939 5310
rect 1975 5310 1979 5314
rect 2195 5310 2199 5314
rect 2283 5310 2287 5314
rect 2339 5310 2343 5314
rect 2483 5310 2487 5314
rect 2491 5310 2495 5314
rect 2651 5310 2655 5314
rect 2675 5310 2679 5314
rect 1975 5198 1979 5202
rect 2023 5198 2027 5202
rect 2159 5198 2163 5202
rect 2223 5198 2227 5202
rect 111 5090 115 5094
rect 347 5090 351 5094
rect 483 5090 487 5094
rect 563 5090 567 5094
rect 619 5090 623 5094
rect 699 5090 703 5094
rect 755 5090 759 5094
rect 835 5090 839 5094
rect 891 5090 895 5094
rect 971 5090 975 5094
rect 1035 5090 1039 5094
rect 1107 5090 1111 5094
rect 1187 5090 1191 5094
rect 1243 5090 1247 5094
rect 1339 5090 1343 5094
rect 1379 5090 1383 5094
rect 1491 5090 1495 5094
rect 1515 5090 1519 5094
rect 1651 5090 1655 5094
rect 1787 5090 1791 5094
rect 1935 5090 1939 5094
rect 111 4978 115 4982
rect 159 4978 163 4982
rect 343 4978 347 4982
rect 375 4978 379 4982
rect 511 4978 515 4982
rect 551 4978 555 4982
rect 111 4858 115 4862
rect 131 4858 135 4862
rect 647 4978 651 4982
rect 751 4978 755 4982
rect 783 4978 787 4982
rect 919 4978 923 4982
rect 943 4978 947 4982
rect 1063 4978 1067 4982
rect 1127 4978 1131 4982
rect 1215 4978 1219 4982
rect 1311 4978 1315 4982
rect 1367 4978 1371 4982
rect 1487 4978 1491 4982
rect 1519 4978 1523 4982
rect 1663 4978 1667 4982
rect 1679 4978 1683 4982
rect 1975 5086 1979 5090
rect 1995 5086 1999 5090
rect 2819 5310 2823 5314
rect 2859 5310 2863 5314
rect 3247 5422 3251 5426
rect 3319 5422 3323 5426
rect 3799 5542 3803 5546
rect 3839 5538 3843 5542
rect 4251 5538 4255 5542
rect 4307 5538 4311 5542
rect 4403 5538 4407 5542
rect 4443 5538 4447 5542
rect 4555 5538 4559 5542
rect 4579 5538 4583 5542
rect 4707 5538 4711 5542
rect 4715 5538 4719 5542
rect 4851 5538 4855 5542
rect 4859 5538 4863 5542
rect 4987 5538 4991 5542
rect 5019 5538 5023 5542
rect 3423 5422 3427 5426
rect 3495 5422 3499 5426
rect 3607 5422 3611 5426
rect 3671 5422 3675 5426
rect 3799 5422 3803 5426
rect 3839 5406 3843 5410
rect 4279 5406 4283 5410
rect 4431 5406 4435 5410
rect 4487 5406 4491 5410
rect 3003 5310 3007 5314
rect 3043 5310 3047 5314
rect 3187 5310 3191 5314
rect 3219 5310 3223 5314
rect 3379 5310 3383 5314
rect 3395 5310 3399 5314
rect 3579 5310 3583 5314
rect 2327 5198 2331 5202
rect 2367 5198 2371 5202
rect 2511 5198 2515 5202
rect 2519 5198 2523 5202
rect 2679 5198 2683 5202
rect 2695 5198 2699 5202
rect 2847 5198 2851 5202
rect 2887 5198 2891 5202
rect 3031 5198 3035 5202
rect 3087 5198 3091 5202
rect 3215 5198 3219 5202
rect 3287 5198 3291 5202
rect 3799 5310 3803 5314
rect 3839 5278 3843 5282
rect 4251 5278 4255 5282
rect 4583 5406 4587 5410
rect 4695 5406 4699 5410
rect 4735 5406 4739 5410
rect 5663 5538 5667 5542
rect 4887 5406 4891 5410
rect 4911 5406 4915 5410
rect 5047 5406 5051 5410
rect 5127 5406 5131 5410
rect 5663 5406 5667 5410
rect 4459 5278 4463 5282
rect 4483 5278 4487 5282
rect 4667 5278 4671 5282
rect 4715 5278 4719 5282
rect 4883 5278 4887 5282
rect 4947 5278 4951 5282
rect 5099 5278 5103 5282
rect 5187 5278 5191 5282
rect 3407 5198 3411 5202
rect 3495 5198 3499 5202
rect 3607 5198 3611 5202
rect 3679 5198 3683 5202
rect 3799 5198 3803 5202
rect 2131 5086 2135 5090
rect 2299 5086 2303 5090
rect 2483 5086 2487 5090
rect 2531 5086 2535 5090
rect 2667 5086 2671 5090
rect 2859 5086 2863 5090
rect 3059 5086 3063 5090
rect 3099 5086 3103 5090
rect 3259 5086 3263 5090
rect 3467 5086 3471 5090
rect 3651 5086 3655 5090
rect 1815 4978 1819 4982
rect 1935 4978 1939 4982
rect 1975 4942 1979 4946
rect 2023 4942 2027 4946
rect 2559 4942 2563 4946
rect 2871 4942 2875 4946
rect 3007 4942 3011 4946
rect 267 4858 271 4862
rect 315 4858 319 4862
rect 403 4858 407 4862
rect 523 4858 527 4862
rect 539 4858 543 4862
rect 675 4858 679 4862
rect 723 4858 727 4862
rect 915 4858 919 4862
rect 1099 4858 1103 4862
rect 1283 4858 1287 4862
rect 1459 4858 1463 4862
rect 1635 4858 1639 4862
rect 1787 4858 1791 4862
rect 1935 4858 1939 4862
rect 3839 5138 3843 5142
rect 3887 5138 3891 5142
rect 4135 5138 4139 5142
rect 4279 5138 4283 5142
rect 4407 5138 4411 5142
rect 3799 5086 3803 5090
rect 3839 5014 3843 5018
rect 3859 5014 3863 5018
rect 4511 5138 4515 5142
rect 4679 5138 4683 5142
rect 4743 5138 4747 5142
rect 5663 5278 5667 5282
rect 4959 5138 4963 5142
rect 4975 5138 4979 5142
rect 5215 5138 5219 5142
rect 5239 5138 5243 5142
rect 5663 5138 5667 5142
rect 4019 5014 4023 5018
rect 4107 5014 4111 5018
rect 4211 5014 4215 5018
rect 4379 5014 4383 5018
rect 4411 5014 4415 5018
rect 4627 5014 4631 5018
rect 4651 5014 4655 5018
rect 3127 4942 3131 4946
rect 3679 4942 3683 4946
rect 3799 4942 3803 4946
rect 1975 4806 1979 4810
rect 1995 4806 1999 4810
rect 2155 4806 2159 4810
rect 2347 4806 2351 4810
rect 2539 4806 2543 4810
rect 2731 4806 2735 4810
rect 2843 4806 2847 4810
rect 2931 4806 2935 4810
rect 2979 4806 2983 4810
rect 3131 4806 3135 4810
rect 111 4738 115 4742
rect 159 4738 163 4742
rect 295 4738 299 4742
rect 343 4738 347 4742
rect 431 4738 435 4742
rect 567 4738 571 4742
rect 703 4738 707 4742
rect 807 4738 811 4742
rect 1055 4738 1059 4742
rect 1311 4738 1315 4742
rect 1575 4738 1579 4742
rect 1815 4738 1819 4742
rect 1935 4738 1939 4742
rect 111 4610 115 4614
rect 131 4610 135 4614
rect 171 4610 175 4614
rect 315 4610 319 4614
rect 395 4610 399 4614
rect 539 4610 543 4614
rect 643 4610 647 4614
rect 779 4610 783 4614
rect 907 4610 911 4614
rect 1027 4610 1031 4614
rect 1195 4610 1199 4614
rect 1283 4610 1287 4614
rect 1491 4610 1495 4614
rect 111 4494 115 4498
rect 199 4494 203 4498
rect 423 4494 427 4498
rect 447 4494 451 4498
rect 655 4494 659 4498
rect 671 4494 675 4498
rect 887 4494 891 4498
rect 935 4494 939 4498
rect 1143 4494 1147 4498
rect 1223 4494 1227 4498
rect 1975 4690 1979 4694
rect 2023 4690 2027 4694
rect 2183 4690 2187 4694
rect 2239 4690 2243 4694
rect 2375 4690 2379 4694
rect 2471 4690 2475 4694
rect 2567 4690 2571 4694
rect 1547 4610 1551 4614
rect 1787 4610 1791 4614
rect 1935 4610 1939 4614
rect 1407 4494 1411 4498
rect 1519 4494 1523 4498
rect 1679 4494 1683 4498
rect 111 4378 115 4382
rect 419 4378 423 4382
rect 627 4378 631 4382
rect 667 4378 671 4382
rect 811 4378 815 4382
rect 859 4378 863 4382
rect 963 4378 967 4382
rect 1115 4378 1119 4382
rect 1123 4378 1127 4382
rect 2695 4690 2699 4694
rect 2759 4690 2763 4694
rect 3839 4882 3843 4886
rect 3887 4882 3891 4886
rect 4047 4882 4051 4886
rect 4071 4882 4075 4886
rect 4239 4882 4243 4886
rect 4287 4882 4291 4886
rect 3799 4806 3803 4810
rect 3839 4766 3843 4770
rect 3859 4766 3863 4770
rect 3915 4766 3919 4770
rect 4843 5014 4847 5018
rect 4931 5014 4935 5018
rect 5067 5014 5071 5018
rect 5211 5014 5215 5018
rect 5299 5014 5303 5018
rect 4439 4882 4443 4886
rect 4511 4882 4515 4886
rect 4655 4882 4659 4886
rect 4735 4882 4739 4886
rect 4871 4882 4875 4886
rect 4959 4882 4963 4886
rect 5095 4882 5099 4886
rect 5183 4882 5187 4886
rect 4043 4766 4047 4770
rect 4187 4766 4191 4770
rect 4259 4766 4263 4770
rect 4467 4766 4471 4770
rect 4483 4766 4487 4770
rect 4707 4766 4711 4770
rect 4763 4766 4767 4770
rect 4931 4766 4935 4770
rect 5067 4766 5071 4770
rect 2919 4690 2923 4694
rect 2959 4690 2963 4694
rect 3143 4690 3147 4694
rect 3159 4690 3163 4694
rect 3367 4690 3371 4694
rect 3799 4690 3803 4694
rect 3839 4654 3843 4658
rect 3943 4654 3947 4658
rect 4063 4654 4067 4658
rect 4215 4654 4219 4658
rect 4327 4654 4331 4658
rect 4495 4654 4499 4658
rect 1975 4574 1979 4578
rect 1995 4574 1999 4578
rect 2099 4574 2103 4578
rect 2211 4574 2215 4578
rect 2347 4574 2351 4578
rect 2443 4574 2447 4578
rect 2579 4574 2583 4578
rect 2667 4574 2671 4578
rect 2795 4574 2799 4578
rect 2891 4574 2895 4578
rect 3003 4574 3007 4578
rect 3115 4574 3119 4578
rect 1815 4494 1819 4498
rect 1935 4494 1939 4498
rect 1975 4454 1979 4458
rect 2127 4454 2131 4458
rect 1291 4378 1295 4382
rect 1379 4378 1383 4382
rect 1467 4378 1471 4382
rect 1651 4378 1655 4382
rect 111 4250 115 4254
rect 695 4250 699 4254
rect 815 4250 819 4254
rect 839 4250 843 4254
rect 951 4250 955 4254
rect 991 4250 995 4254
rect 1087 4250 1091 4254
rect 1151 4250 1155 4254
rect 1223 4250 1227 4254
rect 1319 4250 1323 4254
rect 1359 4250 1363 4254
rect 1495 4250 1499 4254
rect 111 4134 115 4138
rect 731 4134 735 4138
rect 787 4134 791 4138
rect 867 4134 871 4138
rect 923 4134 927 4138
rect 1003 4134 1007 4138
rect 1059 4134 1063 4138
rect 1139 4134 1143 4138
rect 1195 4134 1199 4138
rect 1275 4134 1279 4138
rect 1331 4134 1335 4138
rect 111 3998 115 4002
rect 511 3998 515 4002
rect 663 3998 667 4002
rect 759 3998 763 4002
rect 823 3998 827 4002
rect 111 3858 115 3862
rect 131 3858 135 3862
rect 307 3858 311 3862
rect 483 3858 487 3862
rect 515 3858 519 3862
rect 635 3858 639 3862
rect 723 3858 727 3862
rect 111 3746 115 3750
rect 159 3746 163 3750
rect 335 3746 339 3750
rect 111 3622 115 3626
rect 131 3622 135 3626
rect 147 3622 151 3626
rect 1935 4378 1939 4382
rect 3203 4574 3207 4578
rect 3339 4574 3343 4578
rect 3403 4574 3407 4578
rect 3611 4574 3615 4578
rect 3799 4574 3803 4578
rect 2231 4454 2235 4458
rect 2375 4454 2379 4458
rect 2447 4454 2451 4458
rect 2607 4454 2611 4458
rect 2663 4454 2667 4458
rect 2823 4454 2827 4458
rect 2871 4454 2875 4458
rect 3031 4454 3035 4458
rect 3079 4454 3083 4458
rect 3231 4454 3235 4458
rect 3287 4454 3291 4458
rect 3431 4454 3435 4458
rect 3495 4454 3499 4458
rect 3639 4454 3643 4458
rect 3679 4454 3683 4458
rect 1975 4334 1979 4338
rect 2203 4334 2207 4338
rect 2307 4334 2311 4338
rect 2419 4334 2423 4338
rect 2459 4334 2463 4338
rect 2627 4334 2631 4338
rect 2635 4334 2639 4338
rect 2811 4334 2815 4338
rect 2843 4334 2847 4338
rect 3011 4334 3015 4338
rect 3051 4334 3055 4338
rect 3227 4334 3231 4338
rect 3259 4334 3263 4338
rect 3839 4542 3843 4546
rect 4035 4542 4039 4546
rect 4599 4654 4603 4658
rect 4791 4654 4795 4658
rect 5663 5014 5667 5018
rect 5327 4882 5331 4886
rect 5407 4882 5411 4886
rect 5663 4882 5667 4886
rect 5155 4766 5159 4770
rect 5371 4766 5375 4770
rect 5379 4766 5383 4770
rect 5663 4766 5667 4770
rect 4871 4654 4875 4658
rect 5095 4654 5099 4658
rect 5151 4654 5155 4658
rect 5399 4654 5403 4658
rect 5439 4654 5443 4658
rect 4179 4542 4183 4546
rect 4299 4542 4303 4546
rect 4411 4542 4415 4546
rect 4571 4542 4575 4546
rect 4659 4542 4663 4546
rect 4843 4542 4847 4546
rect 4915 4542 4919 4546
rect 5123 4542 5127 4546
rect 5179 4542 5183 4546
rect 3799 4454 3803 4458
rect 3839 4422 3843 4426
rect 4207 4422 4211 4426
rect 4359 4422 4363 4426
rect 4439 4422 4443 4426
rect 4519 4422 4523 4426
rect 4687 4422 4691 4426
rect 3451 4334 3455 4338
rect 3467 4334 3471 4338
rect 3651 4334 3655 4338
rect 3799 4334 3803 4338
rect 1631 4250 1635 4254
rect 1679 4250 1683 4254
rect 1767 4250 1771 4254
rect 1935 4250 1939 4254
rect 1975 4214 1979 4218
rect 2335 4214 2339 4218
rect 2487 4214 2491 4218
rect 2567 4214 2571 4218
rect 2655 4214 2659 4218
rect 2703 4214 2707 4218
rect 2839 4214 2843 4218
rect 2975 4214 2979 4218
rect 3039 4214 3043 4218
rect 3255 4214 3259 4218
rect 1411 4134 1415 4138
rect 1467 4134 1471 4138
rect 1547 4134 1551 4138
rect 1603 4134 1607 4138
rect 895 3998 899 4002
rect 983 3998 987 4002
rect 1031 3998 1035 4002
rect 1151 3998 1155 4002
rect 1167 3998 1171 4002
rect 1303 3998 1307 4002
rect 1319 3998 1323 4002
rect 795 3858 799 3862
rect 939 3858 943 3862
rect 955 3858 959 3862
rect 1123 3858 1127 3862
rect 1163 3858 1167 3862
rect 527 3746 531 3750
rect 543 3746 547 3750
rect 711 3746 715 3750
rect 751 3746 755 3750
rect 887 3746 891 3750
rect 967 3746 971 3750
rect 1055 3746 1059 3750
rect 1739 4134 1743 4138
rect 1935 4134 1939 4138
rect 1975 4082 1979 4086
rect 2291 4082 2295 4086
rect 2427 4082 2431 4086
rect 2539 4082 2543 4086
rect 2563 4082 2567 4086
rect 2387 4048 2391 4052
rect 1439 3998 1443 4002
rect 1575 3998 1579 4002
rect 1935 3998 1939 4002
rect 1975 3966 1979 3970
rect 2119 3966 2123 3970
rect 2319 3966 2323 3970
rect 2327 3966 2331 3970
rect 2455 3966 2459 3970
rect 2535 3966 2539 3970
rect 1291 3858 1295 3862
rect 1935 3858 1939 3862
rect 1975 3842 1979 3846
rect 2091 3842 2095 3846
rect 2139 3842 2143 3846
rect 3839 4310 3843 4314
rect 3859 4310 3863 4314
rect 4043 4310 4047 4314
rect 4251 4310 4255 4314
rect 4331 4310 4335 4314
rect 3479 4214 3483 4218
rect 3679 4214 3683 4218
rect 3799 4214 3803 4218
rect 3839 4162 3843 4166
rect 3887 4162 3891 4166
rect 2675 4082 2679 4086
rect 2699 4082 2703 4086
rect 2811 4082 2815 4086
rect 2835 4082 2839 4086
rect 2947 4082 2951 4086
rect 3799 4082 3803 4086
rect 2959 4048 2963 4052
rect 4879 4422 4883 4426
rect 4943 4422 4947 4426
rect 5663 4654 5667 4658
rect 5411 4542 5415 4546
rect 5443 4542 5447 4546
rect 5663 4542 5667 4546
rect 5079 4422 5083 4426
rect 5207 4422 5211 4426
rect 5287 4422 5291 4426
rect 5471 4422 5475 4426
rect 5503 4422 5507 4426
rect 4475 4310 4479 4314
rect 4491 4310 4495 4314
rect 4659 4310 4663 4314
rect 4715 4310 4719 4314
rect 4851 4310 4855 4314
rect 4971 4310 4975 4314
rect 5051 4310 5055 4314
rect 5235 4310 5239 4314
rect 5259 4310 5263 4314
rect 5663 4422 5667 4426
rect 5475 4310 5479 4314
rect 5499 4310 5503 4314
rect 5663 4310 5667 4314
rect 4071 4162 4075 4166
rect 4279 4162 4283 4166
rect 4415 4162 4419 4166
rect 4503 4162 4507 4166
rect 4743 4162 4747 4166
rect 4975 4162 4979 4166
rect 4999 4162 5003 4166
rect 5263 4162 5267 4166
rect 5527 4162 5531 4166
rect 5543 4162 5547 4166
rect 5663 4162 5667 4166
rect 3839 4050 3843 4054
rect 3859 4050 3863 4054
rect 4003 4050 4007 4054
rect 4171 4050 4175 4054
rect 4339 4050 4343 4054
rect 4387 4050 4391 4054
rect 4499 4050 4503 4054
rect 4651 4050 4655 4054
rect 4803 4050 4807 4054
rect 4947 4050 4951 4054
rect 5091 4050 5095 4054
rect 5235 4050 5239 4054
rect 5379 4050 5383 4054
rect 5515 4050 5519 4054
rect 2591 3966 2595 3970
rect 2727 3966 2731 3970
rect 2743 3966 2747 3970
rect 2863 3966 2867 3970
rect 2943 3966 2947 3970
rect 3135 3966 3139 3970
rect 3319 3966 3323 3970
rect 3511 3966 3515 3970
rect 3679 3966 3683 3970
rect 3799 3966 3803 3970
rect 2299 3842 2303 3846
rect 2371 3842 2375 3846
rect 2507 3842 2511 3846
rect 2587 3842 2591 3846
rect 2715 3842 2719 3846
rect 2795 3842 2799 3846
rect 2915 3842 2919 3846
rect 2995 3842 2999 3846
rect 1191 3746 1195 3750
rect 1215 3746 1219 3750
rect 1367 3746 1371 3750
rect 1519 3746 1523 3750
rect 1679 3746 1683 3750
rect 1815 3746 1819 3750
rect 1935 3746 1939 3750
rect 1975 3726 1979 3730
rect 2167 3726 2171 3730
rect 2279 3726 2283 3730
rect 307 3622 311 3626
rect 355 3622 359 3626
rect 499 3622 503 3626
rect 571 3622 575 3626
rect 683 3622 687 3626
rect 803 3622 807 3626
rect 859 3622 863 3626
rect 1027 3622 1031 3626
rect 1043 3622 1047 3626
rect 111 3486 115 3490
rect 175 3486 179 3490
rect 303 3486 307 3490
rect 383 3486 387 3490
rect 447 3486 451 3490
rect 599 3486 603 3490
rect 759 3486 763 3490
rect 831 3486 835 3490
rect 111 3358 115 3362
rect 275 3358 279 3362
rect 419 3358 423 3362
rect 467 3358 471 3362
rect 571 3358 575 3362
rect 667 3358 671 3362
rect 731 3358 735 3362
rect 111 3246 115 3250
rect 495 3246 499 3250
rect 535 3246 539 3250
rect 1187 3622 1191 3626
rect 1291 3622 1295 3626
rect 1339 3622 1343 3626
rect 935 3486 939 3490
rect 1071 3486 1075 3490
rect 1111 3486 1115 3490
rect 1491 3622 1495 3626
rect 1547 3622 1551 3626
rect 1651 3622 1655 3626
rect 1787 3622 1791 3626
rect 1295 3486 1299 3490
rect 1319 3486 1323 3490
rect 1487 3486 1491 3490
rect 1575 3486 1579 3490
rect 875 3358 879 3362
rect 907 3358 911 3362
rect 1083 3358 1087 3362
rect 1091 3358 1095 3362
rect 1267 3358 1271 3362
rect 1315 3358 1319 3362
rect 695 3246 699 3250
rect 727 3246 731 3250
rect 903 3246 907 3250
rect 919 3246 923 3250
rect 1111 3246 1115 3250
rect 1119 3246 1123 3250
rect 111 3126 115 3130
rect 427 3126 431 3130
rect 507 3126 511 3130
rect 111 2986 115 2990
rect 199 2986 203 2990
rect 563 3126 567 3130
rect 1935 3622 1939 3626
rect 1975 3602 1979 3606
rect 1995 3602 1999 3606
rect 2251 3602 2255 3606
rect 1815 3486 1819 3490
rect 1935 3486 1939 3490
rect 1975 3482 1979 3486
rect 2023 3482 2027 3486
rect 1459 3358 1463 3362
rect 1935 3358 1939 3362
rect 1295 3246 1299 3250
rect 1343 3246 1347 3250
rect 2399 3726 2403 3730
rect 2479 3726 2483 3730
rect 3839 3914 3843 3918
rect 3887 3914 3891 3918
rect 4031 3914 4035 3918
rect 4199 3914 4203 3918
rect 4367 3914 4371 3918
rect 4383 3914 4387 3918
rect 3107 3842 3111 3846
rect 3195 3842 3199 3846
rect 3291 3842 3295 3846
rect 3403 3842 3407 3846
rect 3483 3842 3487 3846
rect 3651 3842 3655 3846
rect 3799 3842 3803 3846
rect 3011 3824 3015 3828
rect 3419 3824 3423 3828
rect 4527 3914 4531 3918
rect 4599 3914 4603 3918
rect 4679 3914 4683 3918
rect 4823 3914 4827 3918
rect 4831 3914 4835 3918
rect 4975 3914 4979 3918
rect 5063 3914 5067 3918
rect 5119 3914 5123 3918
rect 5263 3914 5267 3918
rect 5311 3914 5315 3918
rect 3839 3786 3843 3790
rect 3995 3786 3999 3790
rect 4203 3786 4207 3790
rect 4355 3786 4359 3790
rect 4435 3786 4439 3790
rect 4571 3786 4575 3790
rect 4691 3786 4695 3790
rect 4795 3786 4799 3790
rect 4963 3786 4967 3790
rect 5035 3786 5039 3790
rect 2615 3726 2619 3730
rect 2679 3726 2683 3730
rect 2823 3726 2827 3730
rect 2879 3726 2883 3730
rect 3023 3726 3027 3730
rect 3079 3726 3083 3730
rect 3223 3726 3227 3730
rect 3279 3726 3283 3730
rect 3431 3726 3435 3730
rect 3799 3726 3803 3730
rect 4091 3728 4095 3732
rect 4939 3731 4943 3732
rect 4939 3728 4943 3731
rect 2451 3602 2455 3606
rect 2515 3602 2519 3606
rect 2651 3602 2655 3606
rect 2755 3602 2759 3606
rect 2851 3602 2855 3606
rect 2979 3602 2983 3606
rect 3051 3602 3055 3606
rect 2191 3482 2195 3486
rect 2279 3482 2283 3486
rect 2399 3482 2403 3486
rect 2543 3482 2547 3486
rect 2615 3482 2619 3486
rect 1975 3330 1979 3334
rect 1995 3330 1999 3334
rect 2163 3330 2167 3334
rect 2195 3330 2199 3334
rect 1471 3246 1475 3250
rect 1655 3246 1659 3250
rect 1815 3246 1819 3250
rect 1935 3246 1939 3250
rect 699 3126 703 3130
rect 835 3126 839 3130
rect 891 3126 895 3130
rect 971 3126 975 3130
rect 1083 3126 1087 3130
rect 1107 3126 1111 3130
rect 1243 3126 1247 3130
rect 1267 3126 1271 3130
rect 1379 3126 1383 3130
rect 1443 3126 1447 3130
rect 1515 3126 1519 3130
rect 3839 3646 3843 3650
rect 4023 3646 4027 3650
rect 4215 3646 4219 3650
rect 4231 3646 4235 3650
rect 4399 3646 4403 3650
rect 4463 3646 4467 3650
rect 4607 3646 4611 3650
rect 4719 3646 4723 3650
rect 3195 3602 3199 3606
rect 3251 3602 3255 3606
rect 3411 3602 3415 3606
rect 3627 3602 3631 3606
rect 3799 3602 3803 3606
rect 2783 3482 2787 3486
rect 2831 3482 2835 3486
rect 3007 3482 3011 3486
rect 3047 3482 3051 3486
rect 3223 3482 3227 3486
rect 3263 3482 3267 3486
rect 3439 3482 3443 3486
rect 3479 3482 3483 3486
rect 3839 3510 3843 3514
rect 4187 3510 4191 3514
rect 4371 3510 4375 3514
rect 4531 3510 4535 3514
rect 4579 3510 4583 3514
rect 3655 3482 3659 3486
rect 3679 3482 3683 3486
rect 3799 3482 3803 3486
rect 5663 4050 5667 4054
rect 5407 3914 5411 3918
rect 5543 3914 5547 3918
rect 5251 3786 5255 3790
rect 5283 3786 5287 3790
rect 4831 3646 4835 3650
rect 4991 3646 4995 3650
rect 5071 3646 5075 3650
rect 5279 3646 5283 3650
rect 5319 3646 5323 3650
rect 5515 3786 5519 3790
rect 5663 3914 5667 3918
rect 5663 3786 5667 3790
rect 5543 3646 5547 3650
rect 4683 3510 4687 3514
rect 4803 3510 4807 3514
rect 4843 3510 4847 3514
rect 5003 3510 5007 3514
rect 5043 3510 5047 3514
rect 5171 3510 5175 3514
rect 5291 3510 5295 3514
rect 5347 3510 5351 3514
rect 3839 3394 3843 3398
rect 3887 3394 3891 3398
rect 4151 3394 4155 3398
rect 4423 3394 4427 3398
rect 4559 3394 4563 3398
rect 4671 3394 4675 3398
rect 4711 3394 4715 3398
rect 4871 3394 4875 3398
rect 4895 3394 4899 3398
rect 5031 3394 5035 3398
rect 5111 3394 5115 3398
rect 5199 3394 5203 3398
rect 2371 3330 2375 3334
rect 2411 3330 2415 3334
rect 2587 3330 2591 3334
rect 2619 3330 2623 3334
rect 2803 3330 2807 3334
rect 2811 3330 2815 3334
rect 3003 3330 3007 3334
rect 3019 3330 3023 3334
rect 3187 3330 3191 3334
rect 3235 3330 3239 3334
rect 3371 3330 3375 3334
rect 3451 3330 3455 3334
rect 3555 3330 3559 3334
rect 3651 3330 3655 3334
rect 3799 3330 3803 3334
rect 1975 3218 1979 3222
rect 2023 3218 2027 3222
rect 2223 3218 2227 3222
rect 2439 3218 2443 3222
rect 2463 3218 2467 3222
rect 2647 3218 2651 3222
rect 2663 3218 2667 3222
rect 1627 3126 1631 3130
rect 1651 3126 1655 3130
rect 1787 3126 1791 3130
rect 1935 3126 1939 3130
rect 455 2986 459 2990
rect 511 2986 515 2990
rect 591 2986 595 2990
rect 727 2986 731 2990
rect 815 2986 819 2990
rect 863 2986 867 2990
rect 999 2986 1003 2990
rect 1111 2986 1115 2990
rect 1135 2986 1139 2990
rect 1271 2986 1275 2990
rect 1407 2986 1411 2990
rect 1415 2986 1419 2990
rect 1543 2986 1547 2990
rect 1679 2986 1683 2990
rect 1719 2986 1723 2990
rect 1815 2986 1819 2990
rect 111 2874 115 2878
rect 131 2874 135 2878
rect 171 2874 175 2878
rect 307 2874 311 2878
rect 483 2874 487 2878
rect 523 2874 527 2878
rect 763 2874 767 2878
rect 787 2874 791 2878
rect 1011 2874 1015 2878
rect 111 2758 115 2762
rect 159 2758 163 2762
rect 279 2758 283 2762
rect 1083 2874 1087 2878
rect 1975 3094 1979 3098
rect 2331 3094 2335 3098
rect 2839 3218 2843 3222
rect 2863 3218 2867 3222
rect 3031 3218 3035 3222
rect 3055 3218 3059 3222
rect 3215 3218 3219 3222
rect 3239 3218 3243 3222
rect 3399 3218 3403 3222
rect 3431 3218 3435 3222
rect 3583 3218 3587 3222
rect 3623 3218 3627 3222
rect 2435 3094 2439 3098
rect 2555 3094 2559 3098
rect 2635 3094 2639 3098
rect 2779 3094 2783 3098
rect 2835 3094 2839 3098
rect 3003 3094 3007 3098
rect 3027 3094 3031 3098
rect 1935 2986 1939 2990
rect 1975 2970 1979 2974
rect 2143 2970 2147 2974
rect 2343 2970 2347 2974
rect 2359 2970 2363 2974
rect 2543 2970 2547 2974
rect 2583 2970 2587 2974
rect 1275 2874 1279 2878
rect 1387 2874 1391 2878
rect 1539 2874 1543 2878
rect 1691 2874 1695 2878
rect 1935 2874 1939 2878
rect 335 2758 339 2762
rect 455 2758 459 2762
rect 551 2758 555 2762
rect 647 2758 651 2762
rect 791 2758 795 2762
rect 855 2758 859 2762
rect 1039 2758 1043 2762
rect 1079 2758 1083 2762
rect 1303 2758 1307 2762
rect 1311 2758 1315 2762
rect 1551 2758 1555 2762
rect 1567 2758 1571 2762
rect 111 2646 115 2650
rect 251 2646 255 2650
rect 427 2646 431 2650
rect 571 2646 575 2650
rect 619 2646 623 2650
rect 731 2646 735 2650
rect 827 2646 831 2650
rect 891 2646 895 2650
rect 111 2534 115 2538
rect 383 2534 387 2538
rect 599 2534 603 2538
rect 759 2534 763 2538
rect 815 2534 819 2538
rect 111 2418 115 2422
rect 227 2418 231 2422
rect 355 2418 359 2422
rect 1043 2646 1047 2650
rect 1051 2646 1055 2650
rect 1195 2646 1199 2650
rect 1283 2646 1287 2650
rect 1355 2646 1359 2650
rect 919 2534 923 2538
rect 1023 2534 1027 2538
rect 1071 2534 1075 2538
rect 1975 2850 1979 2854
rect 2011 2850 2015 2854
rect 2115 2850 2119 2854
rect 2743 2970 2747 2974
rect 2807 2970 2811 2974
rect 2259 2850 2263 2854
rect 2315 2850 2319 2854
rect 2507 2850 2511 2854
rect 2515 2850 2519 2854
rect 1799 2758 1803 2762
rect 1935 2758 1939 2762
rect 1975 2734 1979 2738
rect 2023 2734 2027 2738
rect 2039 2734 2043 2738
rect 1515 2646 1519 2650
rect 1523 2646 1527 2650
rect 1675 2646 1679 2650
rect 1771 2646 1775 2650
rect 1223 2534 1227 2538
rect 1231 2534 1235 2538
rect 1383 2534 1387 2538
rect 1431 2534 1435 2538
rect 1935 2646 1939 2650
rect 2247 2734 2251 2738
rect 2287 2734 2291 2738
rect 2503 2734 2507 2738
rect 3211 3094 3215 3098
rect 3235 3094 3239 3098
rect 3403 3094 3407 3098
rect 3467 3094 3471 3098
rect 2935 2970 2939 2974
rect 3031 2970 3035 2974
rect 3135 2970 3139 2974
rect 3263 2970 3267 2974
rect 3335 2970 3339 2974
rect 2715 2850 2719 2854
rect 2755 2850 2759 2854
rect 2907 2850 2911 2854
rect 3003 2850 3007 2854
rect 2535 2734 2539 2738
rect 2759 2734 2763 2738
rect 2783 2734 2787 2738
rect 1975 2610 1979 2614
rect 1995 2610 1999 2614
rect 2219 2610 2223 2614
rect 2475 2610 2479 2614
rect 3839 3282 3843 3286
rect 3859 3282 3863 3286
rect 3799 3218 3803 3222
rect 3839 3154 3843 3158
rect 3887 3154 3891 3158
rect 3903 3154 3907 3158
rect 3595 3094 3599 3098
rect 3799 3094 3803 3098
rect 4099 3282 4103 3286
rect 4123 3282 4127 3286
rect 4347 3282 4351 3286
rect 4395 3282 4399 3286
rect 4579 3282 4583 3286
rect 4643 3282 4647 3286
rect 4787 3282 4791 3286
rect 4867 3282 4871 3286
rect 4987 3282 4991 3286
rect 5083 3282 5087 3286
rect 4127 3154 4131 3158
rect 4135 3154 4139 3158
rect 4359 3154 4363 3158
rect 4375 3154 4379 3158
rect 3839 3042 3843 3046
rect 3875 3042 3879 3046
rect 3907 3042 3911 3046
rect 4075 3042 4079 3046
rect 4107 3042 4111 3046
rect 4243 3042 4247 3046
rect 4331 3042 4335 3046
rect 4411 3042 4415 3046
rect 3495 2970 3499 2974
rect 3799 2970 3803 2974
rect 3839 2926 3843 2930
rect 3895 2926 3899 2930
rect 3935 2926 3939 2930
rect 3107 2850 3111 2854
rect 3307 2850 3311 2854
rect 3799 2850 3803 2854
rect 4031 2926 4035 2930
rect 4103 2926 4107 2930
rect 4167 2926 4171 2930
rect 4271 2926 4275 2930
rect 4303 2926 4307 2930
rect 3839 2806 3843 2810
rect 3859 2806 3863 2810
rect 3867 2806 3871 2810
rect 3995 2806 3999 2810
rect 4003 2806 4007 2810
rect 5171 3282 5175 3286
rect 5299 3282 5303 3286
rect 5515 3510 5519 3514
rect 5663 3646 5667 3650
rect 5663 3510 5667 3514
rect 5327 3394 5331 3398
rect 5375 3394 5379 3398
rect 5543 3394 5547 3398
rect 5355 3282 5359 3286
rect 5515 3282 5519 3286
rect 5663 3394 5667 3398
rect 5663 3282 5667 3286
rect 4583 3154 4587 3158
rect 4607 3154 4611 3158
rect 4807 3154 4811 3158
rect 4815 3154 4819 3158
rect 5015 3154 5019 3158
rect 5031 3154 5035 3158
rect 5199 3154 5203 3158
rect 5383 3154 5387 3158
rect 5543 3154 5547 3158
rect 5663 3154 5667 3158
rect 4555 3042 4559 3046
rect 4579 3042 4583 3046
rect 4755 3042 4759 3046
rect 4779 3042 4783 3046
rect 5003 3042 5007 3046
rect 5663 3042 5667 3046
rect 4439 2926 4443 2930
rect 4575 2926 4579 2930
rect 4607 2926 4611 2930
rect 4783 2926 4787 2930
rect 5663 2926 5667 2930
rect 4131 2806 4135 2810
rect 4139 2806 4143 2810
rect 4267 2806 4271 2810
rect 4275 2806 4279 2810
rect 4403 2806 4407 2810
rect 4411 2806 4415 2810
rect 4539 2806 4543 2810
rect 4547 2806 4551 2810
rect 4675 2806 4679 2810
rect 4811 2806 4815 2810
rect 5663 2806 5667 2810
rect 3015 2734 3019 2738
rect 3031 2734 3035 2738
rect 3799 2734 3803 2738
rect 3839 2694 3843 2698
rect 3887 2694 3891 2698
rect 3959 2694 3963 2698
rect 4023 2694 4027 2698
rect 2555 2610 2559 2614
rect 2691 2610 2695 2614
rect 2731 2610 2735 2614
rect 2827 2610 2831 2614
rect 2963 2610 2967 2614
rect 2987 2610 2991 2614
rect 3099 2610 3103 2614
rect 1543 2534 1547 2538
rect 1631 2534 1635 2538
rect 1703 2534 1707 2538
rect 1815 2534 1819 2538
rect 1935 2534 1939 2538
rect 523 2418 527 2422
rect 571 2418 575 2422
rect 787 2418 791 2422
rect 835 2418 839 2422
rect 995 2418 999 2422
rect 1155 2418 1159 2422
rect 1203 2418 1207 2422
rect 1403 2418 1407 2422
rect 1483 2418 1487 2422
rect 1603 2418 1607 2422
rect 1787 2418 1791 2422
rect 111 2290 115 2294
rect 159 2290 163 2294
rect 255 2290 259 2294
rect 367 2290 371 2294
rect 551 2290 555 2294
rect 599 2290 603 2294
rect 111 2166 115 2170
rect 131 2166 135 2170
rect 831 2290 835 2294
rect 863 2290 867 2294
rect 1975 2474 1979 2478
rect 2023 2474 2027 2478
rect 2223 2474 2227 2478
rect 2447 2474 2451 2478
rect 2583 2474 2587 2478
rect 2679 2474 2683 2478
rect 2719 2474 2723 2478
rect 1935 2418 1939 2422
rect 1975 2354 1979 2358
rect 1995 2354 1999 2358
rect 1063 2290 1067 2294
rect 1183 2290 1187 2294
rect 1511 2290 1515 2294
rect 1815 2290 1819 2294
rect 1935 2290 1939 2294
rect 2155 2354 2159 2358
rect 2195 2354 2199 2358
rect 2347 2354 2351 2358
rect 2419 2354 2423 2358
rect 2539 2354 2543 2358
rect 339 2166 343 2170
rect 347 2166 351 2170
rect 571 2166 575 2170
rect 595 2166 599 2170
rect 803 2166 807 2170
rect 835 2166 839 2170
rect 1035 2166 1039 2170
rect 1075 2166 1079 2170
rect 111 2050 115 2054
rect 159 2050 163 2054
rect 271 2050 275 2054
rect 375 2050 379 2054
rect 407 2050 411 2054
rect 543 2050 547 2054
rect 623 2050 627 2054
rect 111 1934 115 1938
rect 187 1934 191 1938
rect 243 1934 247 1938
rect 687 2050 691 2054
rect 831 2050 835 2054
rect 863 2050 867 2054
rect 379 1934 383 1938
rect 515 1934 519 1938
rect 587 1934 591 1938
rect 659 1934 663 1938
rect 111 1814 115 1818
rect 159 1814 163 1818
rect 215 1814 219 1818
rect 375 1814 379 1818
rect 407 1814 411 1818
rect 111 1678 115 1682
rect 131 1678 135 1682
rect 1975 2234 1979 2238
rect 2023 2234 2027 2238
rect 2183 2234 2187 2238
rect 2191 2234 2195 2238
rect 2359 2234 2363 2238
rect 2375 2234 2379 2238
rect 1315 2166 1319 2170
rect 1563 2166 1567 2170
rect 1787 2166 1791 2170
rect 1935 2166 1939 2170
rect 975 2050 979 2054
rect 1103 2050 1107 2054
rect 1119 2050 1123 2054
rect 1263 2050 1267 2054
rect 1343 2050 1347 2054
rect 1407 2050 1411 2054
rect 803 1934 807 1938
rect 811 1934 815 1938
rect 947 1934 951 1938
rect 1051 1934 1055 1938
rect 1091 1934 1095 1938
rect 1235 1934 1239 1938
rect 1299 1934 1303 1938
rect 591 1814 595 1818
rect 615 1814 619 1818
rect 799 1814 803 1818
rect 839 1814 843 1818
rect 999 1814 1003 1818
rect 1079 1814 1083 1818
rect 347 1678 351 1682
rect 395 1678 399 1682
rect 111 1554 115 1558
rect 159 1554 163 1558
rect 1543 2050 1547 2054
rect 1591 2050 1595 2054
rect 1679 2050 1683 2054
rect 2855 2474 2859 2478
rect 2927 2474 2931 2478
rect 3799 2610 3803 2614
rect 4159 2694 4163 2698
rect 4255 2694 4259 2698
rect 4295 2694 4299 2698
rect 4431 2694 4435 2698
rect 4543 2694 4547 2698
rect 4567 2694 4571 2698
rect 4703 2694 4707 2698
rect 4823 2694 4827 2698
rect 3839 2582 3843 2586
rect 3859 2582 3863 2586
rect 3931 2582 3935 2586
rect 4083 2582 4087 2586
rect 4227 2582 4231 2586
rect 4331 2582 4335 2586
rect 4515 2582 4519 2586
rect 4579 2582 4583 2586
rect 2991 2474 2995 2478
rect 3127 2474 3131 2478
rect 3183 2474 3187 2478
rect 3439 2474 3443 2478
rect 3679 2474 3683 2478
rect 3799 2474 3803 2478
rect 3839 2466 3843 2470
rect 3887 2466 3891 2470
rect 4087 2466 4091 2470
rect 4111 2466 4115 2470
rect 2651 2354 2655 2358
rect 2731 2354 2735 2358
rect 2899 2354 2903 2358
rect 2923 2354 2927 2358
rect 3115 2354 3119 2358
rect 3155 2354 3159 2358
rect 3299 2354 3303 2358
rect 3411 2354 3415 2358
rect 3483 2354 3487 2358
rect 2535 2234 2539 2238
rect 2567 2234 2571 2238
rect 2711 2234 2715 2238
rect 2759 2234 2763 2238
rect 2879 2234 2883 2238
rect 2951 2234 2955 2238
rect 3047 2234 3051 2238
rect 3143 2234 3147 2238
rect 3207 2234 3211 2238
rect 1975 2106 1979 2110
rect 1995 2106 1999 2110
rect 2163 2106 2167 2110
rect 2331 2106 2335 2110
rect 2507 2106 2511 2110
rect 2683 2106 2687 2110
rect 2851 2106 2855 2110
rect 3019 2106 3023 2110
rect 3107 2106 3111 2110
rect 1815 2050 1819 2054
rect 1935 2050 1939 2054
rect 3327 2234 3331 2238
rect 3367 2234 3371 2238
rect 3651 2354 3655 2358
rect 3799 2354 3803 2358
rect 4327 2466 4331 2470
rect 4359 2466 4363 2470
rect 4839 2694 4843 2698
rect 5111 2694 5115 2698
rect 5399 2694 5403 2698
rect 5663 2694 5667 2698
rect 4795 2582 4799 2586
rect 4827 2582 4831 2586
rect 5075 2582 5079 2586
rect 5083 2582 5087 2586
rect 5323 2582 5327 2586
rect 5371 2582 5375 2586
rect 4583 2466 4587 2470
rect 4607 2466 4611 2470
rect 4847 2466 4851 2470
rect 4855 2466 4859 2470
rect 5103 2466 5107 2470
rect 5119 2466 5123 2470
rect 3839 2342 3843 2346
rect 3859 2342 3863 2346
rect 4059 2342 4063 2346
rect 4299 2342 4303 2346
rect 4443 2342 4447 2346
rect 4555 2342 4559 2346
rect 4611 2342 4615 2346
rect 4787 2342 4791 2346
rect 4819 2342 4823 2346
rect 5663 2582 5667 2586
rect 5351 2466 5355 2470
rect 5399 2466 5403 2470
rect 4963 2342 4967 2346
rect 5091 2342 5095 2346
rect 3511 2234 3515 2238
rect 3535 2234 3539 2238
rect 3679 2234 3683 2238
rect 3799 2234 3803 2238
rect 3839 2218 3843 2222
rect 4471 2218 4475 2222
rect 4543 2218 4547 2222
rect 4639 2218 4643 2222
rect 4719 2218 4723 2222
rect 4815 2218 4819 2222
rect 3179 2106 3183 2110
rect 3243 2106 3247 2110
rect 3339 2106 3343 2110
rect 3379 2106 3383 2110
rect 3507 2106 3511 2110
rect 3515 2106 3519 2110
rect 3651 2106 3655 2110
rect 1379 1934 1383 1938
rect 1515 1934 1519 1938
rect 1555 1934 1559 1938
rect 1651 1934 1655 1938
rect 1787 1934 1791 1938
rect 1191 1814 1195 1818
rect 1327 1814 1331 1818
rect 1383 1814 1387 1818
rect 1575 1814 1579 1818
rect 1583 1814 1587 1818
rect 563 1678 567 1682
rect 683 1678 687 1682
rect 771 1678 775 1682
rect 971 1678 975 1682
rect 979 1678 983 1682
rect 1163 1678 1167 1682
rect 1275 1678 1279 1682
rect 375 1554 379 1558
rect 423 1554 427 1558
rect 607 1554 611 1558
rect 711 1554 715 1558
rect 839 1554 843 1558
rect 111 1430 115 1434
rect 131 1430 135 1434
rect 347 1430 351 1434
rect 411 1430 415 1434
rect 579 1430 583 1434
rect 111 1318 115 1322
rect 159 1318 163 1322
rect 1975 1994 1979 1998
rect 3127 1994 3131 1998
rect 3135 1994 3139 1998
rect 3263 1994 3267 1998
rect 3271 1994 3275 1998
rect 3399 1994 3403 1998
rect 3407 1994 3411 1998
rect 1935 1934 1939 1938
rect 1975 1870 1979 1874
rect 1995 1870 1999 1874
rect 1815 1814 1819 1818
rect 1935 1814 1939 1818
rect 2227 1870 2231 1874
rect 2467 1870 2471 1874
rect 2691 1870 2695 1874
rect 2907 1870 2911 1874
rect 3099 1870 3103 1874
rect 3107 1870 3111 1874
rect 1975 1750 1979 1754
rect 2023 1750 2027 1754
rect 2159 1750 2163 1754
rect 2255 1750 2259 1754
rect 2311 1750 2315 1754
rect 1355 1678 1359 1682
rect 1547 1678 1551 1682
rect 1935 1678 1939 1682
rect 2471 1750 2475 1754
rect 2495 1750 2499 1754
rect 2639 1750 2643 1754
rect 2719 1750 2723 1754
rect 2807 1750 2811 1754
rect 2935 1750 2939 1754
rect 2975 1750 2979 1754
rect 1975 1630 1979 1634
rect 1995 1630 1999 1634
rect 2091 1630 2095 1634
rect 2131 1630 2135 1634
rect 2227 1630 2231 1634
rect 2283 1630 2287 1634
rect 2363 1630 2367 1634
rect 2443 1630 2447 1634
rect 2499 1630 2503 1634
rect 2611 1630 2615 1634
rect 2635 1630 2639 1634
rect 1007 1554 1011 1558
rect 1071 1554 1075 1558
rect 1303 1554 1307 1558
rect 1935 1554 1939 1558
rect 739 1430 743 1434
rect 811 1430 815 1434
rect 1043 1430 1047 1434
rect 1091 1430 1095 1434
rect 1275 1430 1279 1434
rect 359 1318 363 1322
rect 439 1318 443 1322
rect 575 1318 579 1322
rect 767 1318 771 1322
rect 775 1318 779 1322
rect 967 1318 971 1322
rect 111 1194 115 1198
rect 131 1194 135 1198
rect 291 1194 295 1198
rect 331 1194 335 1198
rect 111 1070 115 1074
rect 159 1070 163 1074
rect 175 1070 179 1074
rect 475 1194 479 1198
rect 547 1194 551 1198
rect 659 1194 663 1198
rect 747 1194 751 1198
rect 835 1194 839 1198
rect 319 1070 323 1074
rect 431 1070 435 1074
rect 503 1070 507 1074
rect 687 1070 691 1074
rect 111 946 115 950
rect 147 946 151 950
rect 235 946 239 950
rect 111 818 115 822
rect 175 818 179 822
rect 263 818 267 822
rect 2771 1630 2775 1634
rect 2779 1630 2783 1634
rect 2907 1630 2911 1634
rect 3799 2106 3803 2110
rect 3839 2106 3843 2110
rect 4515 2106 4519 2110
rect 4635 2106 4639 2110
rect 3535 1994 3539 1998
rect 3543 1994 3547 1998
rect 3671 1994 3675 1998
rect 3679 1994 3683 1998
rect 3235 1870 3239 1874
rect 3299 1870 3303 1874
rect 3371 1870 3375 1874
rect 3483 1870 3487 1874
rect 3507 1870 3511 1874
rect 5147 2342 5151 2346
rect 5339 2342 5343 2346
rect 5371 2342 5375 2346
rect 4911 2218 4915 2222
rect 4991 2218 4995 2222
rect 5119 2218 5123 2222
rect 5175 2218 5179 2222
rect 4691 2106 4695 2110
rect 4771 2106 4775 2110
rect 4883 2106 4887 2110
rect 4907 2106 4911 2110
rect 5043 2106 5047 2110
rect 5091 2106 5095 2110
rect 5663 2466 5667 2470
rect 5515 2342 5519 2346
rect 5663 2342 5667 2346
rect 5335 2218 5339 2222
rect 5367 2218 5371 2222
rect 5543 2218 5547 2222
rect 5663 2218 5667 2222
rect 5179 2106 5183 2110
rect 5307 2106 5311 2110
rect 5515 2106 5519 2110
rect 3799 1994 3803 1998
rect 3839 1994 3843 1998
rect 4663 1994 4667 1998
rect 4799 1994 4803 1998
rect 4863 1994 4867 1998
rect 4935 1994 4939 1998
rect 4999 1994 5003 1998
rect 5071 1994 5075 1998
rect 5135 1994 5139 1998
rect 5207 1994 5211 1998
rect 3643 1870 3647 1874
rect 3651 1870 3655 1874
rect 3799 1870 3803 1874
rect 3839 1870 3843 1874
rect 4675 1870 4679 1874
rect 3135 1750 3139 1754
rect 3151 1750 3155 1754
rect 3327 1750 3331 1754
rect 3511 1750 3515 1754
rect 3679 1750 3683 1754
rect 3799 1750 3803 1754
rect 3839 1742 3843 1746
rect 3887 1742 3891 1746
rect 5271 1994 5275 1998
rect 5407 1994 5411 1998
rect 5543 1994 5547 1998
rect 4819 1870 4823 1874
rect 4835 1870 4839 1874
rect 4963 1870 4967 1874
rect 4971 1870 4975 1874
rect 5107 1870 5111 1874
rect 5243 1870 5247 1874
rect 5379 1870 5383 1874
rect 5515 1870 5519 1874
rect 4079 1742 4083 1746
rect 4303 1742 4307 1746
rect 4535 1742 4539 1746
rect 4703 1742 4707 1746
rect 4775 1742 4779 1746
rect 4847 1742 4851 1746
rect 4991 1742 4995 1746
rect 5023 1742 5027 1746
rect 2947 1630 2951 1634
rect 3043 1630 3047 1634
rect 3123 1630 3127 1634
rect 3179 1630 3183 1634
rect 3799 1630 3803 1634
rect 3839 1630 3843 1634
rect 3859 1630 3863 1634
rect 3995 1630 3999 1634
rect 4051 1630 4055 1634
rect 1975 1498 1979 1502
rect 2023 1498 2027 1502
rect 2119 1498 2123 1502
rect 2159 1498 2163 1502
rect 2255 1498 2259 1502
rect 2295 1498 2299 1502
rect 2391 1498 2395 1502
rect 2431 1498 2435 1502
rect 2527 1498 2531 1502
rect 2567 1498 2571 1502
rect 1451 1430 1455 1434
rect 1787 1430 1791 1434
rect 1935 1430 1939 1434
rect 1119 1318 1123 1322
rect 1151 1318 1155 1322
rect 1327 1318 1331 1322
rect 1479 1318 1483 1322
rect 1495 1318 1499 1322
rect 1663 1318 1667 1322
rect 1815 1318 1819 1322
rect 939 1194 943 1198
rect 1003 1194 1007 1198
rect 1123 1194 1127 1198
rect 1171 1194 1175 1198
rect 863 1070 867 1074
rect 951 1070 955 1074
rect 1031 1070 1035 1074
rect 403 946 407 950
rect 459 946 463 950
rect 659 946 663 950
rect 683 946 687 950
rect 431 818 435 822
rect 487 818 491 822
rect 111 706 115 710
rect 131 706 135 710
rect 147 706 151 710
rect 907 946 911 950
rect 923 946 927 950
rect 1975 1378 1979 1382
rect 1995 1378 1999 1382
rect 2131 1378 2135 1382
rect 2267 1378 2271 1382
rect 2275 1378 2279 1382
rect 1935 1318 1939 1322
rect 2663 1498 2667 1502
rect 2703 1498 2707 1502
rect 2799 1498 2803 1502
rect 2839 1498 2843 1502
rect 2935 1498 2939 1502
rect 2975 1498 2979 1502
rect 3071 1498 3075 1502
rect 3207 1498 3211 1502
rect 2403 1378 2407 1382
rect 2539 1378 2543 1382
rect 2563 1378 2567 1382
rect 2675 1378 2679 1382
rect 2811 1378 2815 1382
rect 2843 1378 2847 1382
rect 1975 1242 1979 1246
rect 2023 1242 2027 1246
rect 2303 1242 2307 1246
rect 2591 1242 2595 1246
rect 2655 1242 2659 1246
rect 1299 1194 1303 1198
rect 1331 1194 1335 1198
rect 1467 1194 1471 1198
rect 1491 1194 1495 1198
rect 1635 1194 1639 1198
rect 1651 1194 1655 1198
rect 1787 1194 1791 1198
rect 1935 1194 1939 1198
rect 1975 1114 1979 1118
rect 1995 1114 1999 1118
rect 1199 1070 1203 1074
rect 1215 1070 1219 1074
rect 1359 1070 1363 1074
rect 1519 1070 1523 1074
rect 1679 1070 1683 1074
rect 1815 1070 1819 1074
rect 1935 1070 1939 1074
rect 1975 1002 1979 1006
rect 2023 1002 2027 1006
rect 1131 946 1135 950
rect 1187 946 1191 950
rect 1363 946 1367 950
rect 1935 946 1939 950
rect 671 818 675 822
rect 711 818 715 822
rect 903 818 907 822
rect 935 818 939 822
rect 1127 818 1131 822
rect 1159 818 1163 822
rect 1351 818 1355 822
rect 1391 818 1395 822
rect 315 706 319 710
rect 403 706 407 710
rect 523 706 527 710
rect 643 706 647 710
rect 723 706 727 710
rect 111 594 115 598
rect 159 594 163 598
rect 343 594 347 598
rect 375 594 379 598
rect 111 482 115 486
rect 131 482 135 486
rect 155 482 159 486
rect 551 594 555 598
rect 599 594 603 598
rect 2171 1114 2175 1118
rect 4155 1630 4159 1634
rect 4275 1630 4279 1634
rect 4355 1630 4359 1634
rect 4507 1630 4511 1634
rect 4587 1630 4591 1634
rect 4747 1630 4751 1634
rect 4851 1630 4855 1634
rect 3839 1518 3843 1522
rect 3887 1518 3891 1522
rect 4023 1518 4027 1522
rect 3799 1498 3803 1502
rect 4159 1518 4163 1522
rect 4183 1518 4187 1522
rect 2947 1378 2951 1382
rect 3123 1378 3127 1382
rect 3395 1378 3399 1382
rect 3651 1378 3655 1382
rect 2831 1242 2835 1246
rect 2871 1242 2875 1246
rect 3007 1242 3011 1246
rect 3151 1242 3155 1246
rect 3183 1242 3187 1246
rect 3359 1242 3363 1246
rect 2363 1114 2367 1118
rect 2547 1114 2551 1118
rect 2627 1114 2631 1118
rect 2723 1114 2727 1118
rect 2803 1114 2807 1118
rect 2891 1114 2895 1118
rect 2979 1114 2983 1118
rect 3059 1114 3063 1118
rect 3155 1114 3159 1118
rect 3219 1114 3223 1118
rect 2191 1002 2195 1006
rect 2199 1002 2203 1006
rect 2375 1002 2379 1006
rect 2391 1002 2395 1006
rect 3839 1402 3843 1406
rect 3859 1402 3863 1406
rect 3799 1378 3803 1382
rect 4303 1518 4307 1522
rect 4383 1518 4387 1522
rect 3995 1402 3999 1406
rect 4059 1402 4063 1406
rect 4131 1402 4135 1406
rect 5135 1742 5139 1746
rect 5271 1742 5275 1746
rect 5279 1742 5283 1746
rect 5407 1742 5411 1746
rect 5663 2106 5667 2110
rect 5663 1994 5667 1998
rect 5663 1870 5667 1874
rect 5535 1742 5539 1746
rect 5543 1742 5547 1746
rect 5663 1742 5667 1746
rect 4995 1630 4999 1634
rect 5131 1630 5135 1634
rect 5251 1630 5255 1634
rect 5419 1630 5423 1634
rect 5507 1630 5511 1634
rect 4495 1518 4499 1522
rect 4615 1518 4619 1522
rect 4719 1518 4723 1522
rect 4879 1518 4883 1522
rect 4967 1518 4971 1522
rect 5159 1518 5163 1522
rect 5223 1518 5227 1522
rect 5447 1518 5451 1522
rect 4275 1402 4279 1406
rect 4307 1402 4311 1406
rect 4467 1402 4471 1406
rect 4579 1402 4583 1406
rect 4691 1402 4695 1406
rect 4875 1402 4879 1406
rect 4939 1402 4943 1406
rect 5187 1402 5191 1406
rect 5195 1402 5199 1406
rect 5459 1402 5463 1406
rect 3839 1282 3843 1286
rect 3887 1282 3891 1286
rect 4087 1282 4091 1286
rect 4335 1282 4339 1286
rect 4607 1282 4611 1286
rect 4615 1282 4619 1286
rect 3423 1242 3427 1246
rect 3543 1242 3547 1246
rect 3679 1242 3683 1246
rect 3799 1242 3803 1246
rect 4791 1282 4795 1286
rect 4903 1282 4907 1286
rect 4975 1282 4979 1286
rect 5167 1282 5171 1286
rect 5215 1282 5219 1286
rect 5367 1282 5371 1286
rect 3839 1166 3843 1170
rect 4587 1166 4591 1170
rect 4763 1166 4767 1170
rect 4835 1166 4839 1170
rect 4947 1166 4951 1170
rect 4971 1166 4975 1170
rect 3331 1114 3335 1118
rect 3387 1114 3391 1118
rect 3515 1114 3519 1118
rect 3799 1114 3803 1118
rect 2567 1002 2571 1006
rect 2575 1002 2579 1006
rect 2751 1002 2755 1006
rect 2759 1002 2763 1006
rect 2919 1002 2923 1006
rect 2943 1002 2947 1006
rect 3087 1002 3091 1006
rect 3127 1002 3131 1006
rect 3247 1002 3251 1006
rect 3311 1002 3315 1006
rect 1975 886 1979 890
rect 1995 886 1999 890
rect 2163 886 2167 890
rect 2179 886 2183 890
rect 2347 886 2351 890
rect 2403 886 2407 890
rect 2539 886 2543 890
rect 2675 886 2679 890
rect 2731 886 2735 890
rect 5487 1518 5491 1522
rect 5663 1630 5667 1634
rect 5663 1518 5667 1522
rect 5499 1402 5503 1406
rect 5663 1402 5667 1406
rect 5527 1282 5531 1286
rect 5543 1282 5547 1286
rect 5107 1166 5111 1170
rect 5139 1166 5143 1170
rect 5243 1166 5247 1170
rect 5339 1166 5343 1170
rect 5379 1166 5383 1170
rect 3839 1050 3843 1054
rect 4807 1050 4811 1054
rect 4863 1050 4867 1054
rect 4943 1050 4947 1054
rect 4999 1050 5003 1054
rect 5079 1050 5083 1054
rect 5135 1050 5139 1054
rect 5215 1050 5219 1054
rect 5271 1050 5275 1054
rect 5351 1050 5355 1054
rect 5407 1050 5411 1054
rect 3415 1002 3419 1006
rect 3495 1002 3499 1006
rect 3679 1002 3683 1006
rect 3799 1002 3803 1006
rect 2915 886 2919 890
rect 2987 886 2991 890
rect 3099 886 3103 890
rect 3283 886 3287 890
rect 3323 886 3327 890
rect 3467 886 3471 890
rect 3651 886 3655 890
rect 3839 934 3843 938
rect 3859 934 3863 938
rect 3995 934 3999 938
rect 4171 934 4175 938
rect 4387 934 4391 938
rect 4643 934 4647 938
rect 4779 934 4783 938
rect 4915 934 4919 938
rect 4931 934 4935 938
rect 5051 934 5055 938
rect 3799 886 3803 890
rect 1575 818 1579 822
rect 1935 818 1939 822
rect 3839 822 3843 826
rect 3887 822 3891 826
rect 875 706 879 710
rect 907 706 911 710
rect 1083 706 1087 710
rect 1099 706 1103 710
rect 1259 706 1263 710
rect 1323 706 1327 710
rect 1427 706 1431 710
rect 1547 706 1551 710
rect 1595 706 1599 710
rect 1771 706 1775 710
rect 1935 706 1939 710
rect 751 594 755 598
rect 807 594 811 598
rect 935 594 939 598
rect 999 594 1003 598
rect 1111 594 1115 598
rect 1175 594 1179 598
rect 1287 594 1291 598
rect 1343 594 1347 598
rect 1455 594 1459 598
rect 1511 594 1515 598
rect 1623 594 1627 598
rect 1671 594 1675 598
rect 1799 594 1803 598
rect 1815 594 1819 598
rect 347 482 351 486
rect 483 482 487 486
rect 571 482 575 486
rect 779 482 783 486
rect 811 482 815 486
rect 971 482 975 486
rect 1139 482 1143 486
rect 1147 482 1151 486
rect 1315 482 1319 486
rect 1475 482 1479 486
rect 1483 482 1487 486
rect 1643 482 1647 486
rect 1787 482 1791 486
rect 111 358 115 362
rect 183 358 187 362
rect 279 358 283 362
rect 487 358 491 362
rect 511 358 515 362
rect 111 206 115 210
rect 131 206 135 210
rect 251 206 255 210
rect 267 206 271 210
rect 703 358 707 362
rect 839 358 843 362
rect 919 358 923 362
rect 1935 594 1939 598
rect 4023 822 4027 826
rect 3839 706 3843 710
rect 3859 706 3863 710
rect 4159 822 4163 826
rect 4199 822 4203 826
rect 5663 1282 5667 1286
rect 5515 1166 5519 1170
rect 5663 1166 5667 1170
rect 5487 1050 5491 1054
rect 5543 1050 5547 1054
rect 5187 934 5191 938
rect 5235 934 5239 938
rect 5323 934 5327 938
rect 5459 934 5463 938
rect 5515 934 5519 938
rect 4295 822 4299 826
rect 4415 822 4419 826
rect 4431 822 4435 826
rect 4567 822 4571 826
rect 4671 822 4675 826
rect 4719 822 4723 826
rect 4895 822 4899 826
rect 4959 822 4963 826
rect 3995 706 3999 710
rect 4131 706 4135 710
rect 4267 706 4271 710
rect 4403 706 4407 710
rect 4539 706 4543 710
rect 3839 594 3843 598
rect 3887 594 3891 598
rect 1975 574 1979 578
rect 2023 574 2027 578
rect 2207 574 2211 578
rect 2431 574 2435 578
rect 2703 574 2707 578
rect 3015 574 3019 578
rect 3135 574 3139 578
rect 3271 574 3275 578
rect 3351 574 3355 578
rect 3407 574 3411 578
rect 3543 574 3547 578
rect 3679 574 3683 578
rect 3799 574 3803 578
rect 1935 482 1939 486
rect 1975 462 1979 466
rect 1995 462 1999 466
rect 2203 462 2207 466
rect 2427 462 2431 466
rect 2651 462 2655 466
rect 2859 462 2863 466
rect 3067 462 3071 466
rect 3107 462 3111 466
rect 1135 358 1139 362
rect 1167 358 1171 362
rect 1503 358 1507 362
rect 1815 358 1819 362
rect 1935 358 1939 362
rect 1975 334 1979 338
rect 2023 334 2027 338
rect 2159 334 2163 338
rect 2231 334 2235 338
rect 2295 334 2299 338
rect 2431 334 2435 338
rect 2455 334 2459 338
rect 2567 334 2571 338
rect 2679 334 2683 338
rect 403 206 407 210
rect 459 206 463 210
rect 539 206 543 210
rect 675 206 679 210
rect 811 206 815 210
rect 891 206 895 210
rect 947 206 951 210
rect 1083 206 1087 210
rect 1107 206 1111 210
rect 1935 206 1939 210
rect 1975 186 1979 190
rect 1995 186 1999 190
rect 2703 334 2707 338
rect 2839 334 2843 338
rect 2887 334 2891 338
rect 5087 822 5091 826
rect 5263 822 5267 826
rect 5287 822 5291 826
rect 5487 822 5491 826
rect 5543 822 5547 826
rect 5663 1050 5667 1054
rect 5663 934 5667 938
rect 4691 706 4695 710
rect 4699 706 4703 710
rect 4867 706 4871 710
rect 4891 706 4895 710
rect 5059 706 5063 710
rect 5099 706 5103 710
rect 5259 706 5263 710
rect 5315 706 5319 710
rect 5459 706 5463 710
rect 5515 706 5519 710
rect 4023 594 4027 598
rect 4071 594 4075 598
rect 4159 594 4163 598
rect 4295 594 4299 598
rect 4311 594 4315 598
rect 4431 594 4435 598
rect 4567 594 4571 598
rect 4575 594 4579 598
rect 4727 594 4731 598
rect 4855 594 4859 598
rect 4919 594 4923 598
rect 5127 594 5131 598
rect 5151 594 5155 598
rect 5343 594 5347 598
rect 3839 470 3843 474
rect 3859 470 3863 474
rect 4043 470 4047 474
rect 4283 470 4287 474
rect 4451 470 4455 474
rect 4547 470 4551 474
rect 3243 462 3247 466
rect 3267 462 3271 466
rect 3379 462 3383 466
rect 3467 462 3471 466
rect 3515 462 3519 466
rect 3651 462 3655 466
rect 3799 462 3803 466
rect 5663 822 5667 826
rect 5663 706 5667 710
rect 5447 594 5451 598
rect 5543 594 5547 598
rect 5663 594 5667 598
rect 4643 470 4647 474
rect 4827 470 4831 474
rect 4843 470 4847 474
rect 5051 470 5055 474
rect 5123 470 5127 474
rect 5267 470 5271 474
rect 3839 354 3843 358
rect 4479 354 4483 358
rect 4615 354 4619 358
rect 4671 354 4675 358
rect 4775 354 4779 358
rect 4871 354 4875 358
rect 4951 354 4955 358
rect 5079 354 5083 358
rect 2975 334 2979 338
rect 3095 334 3099 338
rect 3111 334 3115 338
rect 3247 334 3251 338
rect 3295 334 3299 338
rect 3383 334 3387 338
rect 3495 334 3499 338
rect 3519 334 3523 338
rect 3655 334 3659 338
rect 3679 334 3683 338
rect 3799 334 3803 338
rect 2131 186 2135 190
rect 2267 186 2271 190
rect 2403 186 2407 190
rect 2539 186 2543 190
rect 2675 186 2679 190
rect 2811 186 2815 190
rect 2947 186 2951 190
rect 3839 202 3843 206
rect 4291 202 4295 206
rect 3083 186 3087 190
rect 3219 186 3223 190
rect 3355 186 3359 190
rect 3491 186 3495 190
rect 3627 186 3631 190
rect 3799 186 3803 190
rect 3043 128 3047 132
rect 3647 131 3651 132
rect 3647 128 3651 131
rect 5135 354 5139 358
rect 5295 354 5299 358
rect 5327 354 5331 358
rect 4427 202 4431 206
rect 4563 202 4567 206
rect 4587 202 4591 206
rect 4699 202 4703 206
rect 4747 202 4751 206
rect 4835 202 4839 206
rect 4923 202 4927 206
rect 4971 202 4975 206
rect 5107 202 5111 206
rect 5243 202 5247 206
rect 5299 202 5303 206
rect 5419 470 5423 474
rect 5483 470 5487 474
rect 5663 470 5667 474
rect 5511 354 5515 358
rect 5527 354 5531 358
rect 5663 354 5667 358
rect 5379 202 5383 206
rect 5499 202 5503 206
rect 5515 202 5519 206
rect 5663 202 5667 206
rect 111 94 115 98
rect 159 94 163 98
rect 295 94 299 98
rect 431 94 435 98
rect 567 94 571 98
rect 703 94 707 98
rect 839 94 843 98
rect 975 94 979 98
rect 1111 94 1115 98
rect 1935 94 1939 98
rect 3839 90 3843 94
rect 4319 90 4323 94
rect 4455 90 4459 94
rect 4591 90 4595 94
rect 4727 90 4731 94
rect 4863 90 4867 94
rect 4999 90 5003 94
rect 5135 90 5139 94
rect 5271 90 5275 94
rect 5407 90 5411 94
rect 5543 90 5547 94
rect 5663 90 5667 94
rect 1975 74 1979 78
rect 2023 74 2027 78
rect 2159 74 2163 78
rect 2295 74 2299 78
rect 2431 74 2435 78
rect 2567 74 2571 78
rect 2703 74 2707 78
rect 2839 74 2843 78
rect 2975 74 2979 78
rect 3111 74 3115 78
rect 3247 74 3251 78
rect 3383 74 3387 78
rect 3519 74 3523 78
rect 3655 74 3659 78
rect 3799 74 3803 78
<< m4 >>
rect 84 5753 85 5759
rect 91 5758 1947 5759
rect 91 5754 111 5758
rect 115 5754 159 5758
rect 163 5754 295 5758
rect 299 5754 1935 5758
rect 1939 5754 1947 5758
rect 91 5753 1947 5754
rect 1953 5753 1954 5759
rect 1946 5653 1947 5659
rect 1953 5658 3811 5659
rect 1953 5654 1975 5658
rect 1979 5654 2023 5658
rect 2027 5654 2183 5658
rect 2187 5654 2367 5658
rect 2371 5654 2551 5658
rect 2555 5654 2727 5658
rect 2731 5654 2895 5658
rect 2899 5654 3063 5658
rect 3067 5654 3223 5658
rect 3227 5654 3383 5658
rect 3387 5654 3543 5658
rect 3547 5654 3679 5658
rect 3683 5654 3799 5658
rect 3803 5654 3811 5658
rect 1953 5653 3811 5654
rect 3817 5655 3818 5659
rect 3817 5654 5702 5655
rect 3817 5653 3839 5654
rect 3810 5650 3839 5653
rect 3843 5650 4335 5654
rect 4339 5650 4471 5654
rect 4475 5650 4607 5654
rect 4611 5650 4743 5654
rect 4747 5650 4879 5654
rect 4883 5650 5015 5654
rect 5019 5650 5663 5654
rect 5667 5650 5702 5654
rect 3810 5649 5702 5650
rect 96 5641 97 5647
rect 103 5646 1959 5647
rect 103 5642 111 5646
rect 115 5642 131 5646
rect 135 5642 267 5646
rect 271 5642 275 5646
rect 279 5642 475 5646
rect 479 5642 699 5646
rect 703 5642 955 5646
rect 959 5642 1227 5646
rect 1231 5642 1515 5646
rect 1519 5642 1787 5646
rect 1791 5642 1935 5646
rect 1939 5642 1959 5646
rect 103 5641 1959 5642
rect 1965 5641 1966 5647
rect 1958 5541 1959 5547
rect 1965 5546 3823 5547
rect 1965 5542 1975 5546
rect 1979 5542 1995 5546
rect 1999 5542 2139 5546
rect 2143 5542 2155 5546
rect 2159 5542 2339 5546
rect 2343 5542 2355 5546
rect 2359 5542 2523 5546
rect 2527 5542 2563 5546
rect 2567 5542 2699 5546
rect 2703 5542 2755 5546
rect 2759 5542 2867 5546
rect 2871 5542 2939 5546
rect 2943 5542 3035 5546
rect 3039 5542 3115 5546
rect 3119 5542 3195 5546
rect 3199 5542 3291 5546
rect 3295 5542 3355 5546
rect 3359 5542 3467 5546
rect 3471 5542 3515 5546
rect 3519 5542 3643 5546
rect 3647 5542 3651 5546
rect 3655 5542 3799 5546
rect 3803 5542 3823 5546
rect 1965 5541 3823 5542
rect 3829 5543 3830 5547
rect 3829 5542 5714 5543
rect 3829 5541 3839 5542
rect 3822 5538 3839 5541
rect 3843 5538 4251 5542
rect 4255 5538 4307 5542
rect 4311 5538 4403 5542
rect 4407 5538 4443 5542
rect 4447 5538 4555 5542
rect 4559 5538 4579 5542
rect 4583 5538 4707 5542
rect 4711 5538 4715 5542
rect 4719 5538 4851 5542
rect 4855 5538 4859 5542
rect 4863 5538 4987 5542
rect 4991 5538 5019 5542
rect 5023 5538 5663 5542
rect 5667 5538 5714 5542
rect 3822 5537 5714 5538
rect 84 5529 85 5535
rect 91 5534 1947 5535
rect 91 5530 111 5534
rect 115 5530 159 5534
rect 163 5530 279 5534
rect 283 5530 303 5534
rect 307 5530 503 5534
rect 507 5530 519 5534
rect 523 5530 727 5534
rect 731 5530 767 5534
rect 771 5530 983 5534
rect 987 5530 1015 5534
rect 1019 5530 1255 5534
rect 1259 5530 1263 5534
rect 1267 5530 1511 5534
rect 1515 5530 1543 5534
rect 1547 5530 1767 5534
rect 1771 5530 1815 5534
rect 1819 5530 1935 5534
rect 1939 5530 1947 5534
rect 91 5529 1947 5530
rect 1953 5529 1954 5535
rect 1946 5427 1947 5433
rect 1953 5427 1978 5433
rect 1972 5426 3811 5427
rect 96 5417 97 5423
rect 103 5422 1959 5423
rect 103 5418 111 5422
rect 115 5418 251 5422
rect 255 5418 411 5422
rect 415 5418 491 5422
rect 495 5418 611 5422
rect 615 5418 739 5422
rect 743 5418 819 5422
rect 823 5418 987 5422
rect 991 5418 1035 5422
rect 1039 5418 1235 5422
rect 1239 5418 1259 5422
rect 1263 5418 1483 5422
rect 1487 5418 1491 5422
rect 1495 5418 1739 5422
rect 1743 5418 1935 5422
rect 1939 5418 1959 5422
rect 103 5417 1959 5418
rect 1965 5417 1966 5423
rect 1972 5422 1975 5426
rect 1979 5422 2167 5426
rect 2171 5422 2311 5426
rect 2315 5422 2383 5426
rect 2387 5422 2511 5426
rect 2515 5422 2591 5426
rect 2595 5422 2703 5426
rect 2707 5422 2783 5426
rect 2787 5422 2887 5426
rect 2891 5422 2967 5426
rect 2971 5422 3071 5426
rect 3075 5422 3143 5426
rect 3147 5422 3247 5426
rect 3251 5422 3319 5426
rect 3323 5422 3423 5426
rect 3427 5422 3495 5426
rect 3499 5422 3607 5426
rect 3611 5422 3671 5426
rect 3675 5422 3799 5426
rect 3803 5422 3811 5426
rect 1972 5421 3811 5422
rect 3817 5421 3818 5427
rect 3810 5405 3811 5411
rect 3817 5410 5695 5411
rect 3817 5406 3839 5410
rect 3843 5406 4279 5410
rect 4283 5406 4431 5410
rect 4435 5406 4487 5410
rect 4491 5406 4583 5410
rect 4587 5406 4695 5410
rect 4699 5406 4735 5410
rect 4739 5406 4887 5410
rect 4891 5406 4911 5410
rect 4915 5406 5047 5410
rect 5051 5406 5127 5410
rect 5131 5406 5663 5410
rect 5667 5406 5695 5410
rect 3817 5405 5695 5406
rect 5701 5405 5702 5411
rect 84 5305 85 5311
rect 91 5310 1947 5311
rect 91 5306 111 5310
rect 115 5306 439 5310
rect 443 5306 591 5310
rect 595 5306 639 5310
rect 643 5306 727 5310
rect 731 5306 847 5310
rect 851 5306 863 5310
rect 867 5306 999 5310
rect 1003 5306 1063 5310
rect 1067 5306 1135 5310
rect 1139 5306 1271 5310
rect 1275 5306 1287 5310
rect 1291 5306 1407 5310
rect 1411 5306 1519 5310
rect 1523 5306 1543 5310
rect 1547 5306 1935 5310
rect 1939 5306 1947 5310
rect 91 5305 1947 5306
rect 1953 5305 1954 5311
rect 1958 5309 1959 5315
rect 1965 5314 3823 5315
rect 1965 5310 1975 5314
rect 1979 5310 2195 5314
rect 2199 5310 2283 5314
rect 2287 5310 2339 5314
rect 2343 5310 2483 5314
rect 2487 5310 2491 5314
rect 2495 5310 2651 5314
rect 2655 5310 2675 5314
rect 2679 5310 2819 5314
rect 2823 5310 2859 5314
rect 2863 5310 3003 5314
rect 3007 5310 3043 5314
rect 3047 5310 3187 5314
rect 3191 5310 3219 5314
rect 3223 5310 3379 5314
rect 3383 5310 3395 5314
rect 3399 5310 3579 5314
rect 3583 5310 3799 5314
rect 3803 5310 3823 5314
rect 1965 5309 3823 5310
rect 3829 5309 3830 5315
rect 3822 5277 3823 5283
rect 3829 5282 5707 5283
rect 3829 5278 3839 5282
rect 3843 5278 4251 5282
rect 4255 5278 4459 5282
rect 4463 5278 4483 5282
rect 4487 5278 4667 5282
rect 4671 5278 4715 5282
rect 4719 5278 4883 5282
rect 4887 5278 4947 5282
rect 4951 5278 5099 5282
rect 5103 5278 5187 5282
rect 5191 5278 5663 5282
rect 5667 5278 5707 5282
rect 3829 5277 5707 5278
rect 5713 5277 5714 5283
rect 1946 5197 1947 5203
rect 1953 5202 3811 5203
rect 1953 5198 1975 5202
rect 1979 5198 2023 5202
rect 2027 5198 2159 5202
rect 2163 5198 2223 5202
rect 2227 5198 2327 5202
rect 2331 5198 2367 5202
rect 2371 5198 2511 5202
rect 2515 5198 2519 5202
rect 2523 5198 2679 5202
rect 2683 5198 2695 5202
rect 2699 5198 2847 5202
rect 2851 5198 2887 5202
rect 2891 5198 3031 5202
rect 3035 5198 3087 5202
rect 3091 5198 3215 5202
rect 3219 5198 3287 5202
rect 3291 5198 3407 5202
rect 3411 5198 3495 5202
rect 3499 5198 3607 5202
rect 3611 5198 3679 5202
rect 3683 5198 3799 5202
rect 3803 5198 3811 5202
rect 1953 5197 3811 5198
rect 3817 5197 3818 5203
rect 3810 5137 3811 5143
rect 3817 5142 5695 5143
rect 3817 5138 3839 5142
rect 3843 5138 3887 5142
rect 3891 5138 4135 5142
rect 4139 5138 4279 5142
rect 4283 5138 4407 5142
rect 4411 5138 4511 5142
rect 4515 5138 4679 5142
rect 4683 5138 4743 5142
rect 4747 5138 4959 5142
rect 4963 5138 4975 5142
rect 4979 5138 5215 5142
rect 5219 5138 5239 5142
rect 5243 5138 5663 5142
rect 5667 5138 5695 5142
rect 3817 5137 5695 5138
rect 5701 5137 5702 5143
rect 96 5089 97 5095
rect 103 5094 1959 5095
rect 103 5090 111 5094
rect 115 5090 347 5094
rect 351 5090 483 5094
rect 487 5090 563 5094
rect 567 5090 619 5094
rect 623 5090 699 5094
rect 703 5090 755 5094
rect 759 5090 835 5094
rect 839 5090 891 5094
rect 895 5090 971 5094
rect 975 5090 1035 5094
rect 1039 5090 1107 5094
rect 1111 5090 1187 5094
rect 1191 5090 1243 5094
rect 1247 5090 1339 5094
rect 1343 5090 1379 5094
rect 1383 5090 1491 5094
rect 1495 5090 1515 5094
rect 1519 5090 1651 5094
rect 1655 5090 1787 5094
rect 1791 5090 1935 5094
rect 1939 5090 1959 5094
rect 103 5089 1959 5090
rect 1965 5091 1966 5095
rect 1965 5090 3830 5091
rect 1965 5089 1975 5090
rect 1958 5086 1975 5089
rect 1979 5086 1995 5090
rect 1999 5086 2131 5090
rect 2135 5086 2299 5090
rect 2303 5086 2483 5090
rect 2487 5086 2531 5090
rect 2535 5086 2667 5090
rect 2671 5086 2859 5090
rect 2863 5086 3059 5090
rect 3063 5086 3099 5090
rect 3103 5086 3259 5090
rect 3263 5086 3467 5090
rect 3471 5086 3651 5090
rect 3655 5086 3799 5090
rect 3803 5086 3830 5090
rect 1958 5085 3830 5086
rect 3822 5013 3823 5019
rect 3829 5018 5707 5019
rect 3829 5014 3839 5018
rect 3843 5014 3859 5018
rect 3863 5014 4019 5018
rect 4023 5014 4107 5018
rect 4111 5014 4211 5018
rect 4215 5014 4379 5018
rect 4383 5014 4411 5018
rect 4415 5014 4627 5018
rect 4631 5014 4651 5018
rect 4655 5014 4843 5018
rect 4847 5014 4931 5018
rect 4935 5014 5067 5018
rect 5071 5014 5211 5018
rect 5215 5014 5299 5018
rect 5303 5014 5663 5018
rect 5667 5014 5707 5018
rect 3829 5013 5707 5014
rect 5713 5013 5714 5019
rect 84 4977 85 4983
rect 91 4982 1947 4983
rect 91 4978 111 4982
rect 115 4978 159 4982
rect 163 4978 343 4982
rect 347 4978 375 4982
rect 379 4978 511 4982
rect 515 4978 551 4982
rect 555 4978 647 4982
rect 651 4978 751 4982
rect 755 4978 783 4982
rect 787 4978 919 4982
rect 923 4978 943 4982
rect 947 4978 1063 4982
rect 1067 4978 1127 4982
rect 1131 4978 1215 4982
rect 1219 4978 1311 4982
rect 1315 4978 1367 4982
rect 1371 4978 1487 4982
rect 1491 4978 1519 4982
rect 1523 4978 1663 4982
rect 1667 4978 1679 4982
rect 1683 4978 1815 4982
rect 1819 4978 1935 4982
rect 1939 4978 1947 4982
rect 91 4977 1947 4978
rect 1953 4977 1954 4983
rect 1946 4941 1947 4947
rect 1953 4946 3811 4947
rect 1953 4942 1975 4946
rect 1979 4942 2023 4946
rect 2027 4942 2559 4946
rect 2563 4942 2871 4946
rect 2875 4942 3007 4946
rect 3011 4942 3127 4946
rect 3131 4942 3679 4946
rect 3683 4942 3799 4946
rect 3803 4942 3811 4946
rect 1953 4941 3811 4942
rect 3817 4941 3818 4947
rect 3810 4881 3811 4887
rect 3817 4886 5695 4887
rect 3817 4882 3839 4886
rect 3843 4882 3887 4886
rect 3891 4882 4047 4886
rect 4051 4882 4071 4886
rect 4075 4882 4239 4886
rect 4243 4882 4287 4886
rect 4291 4882 4439 4886
rect 4443 4882 4511 4886
rect 4515 4882 4655 4886
rect 4659 4882 4735 4886
rect 4739 4882 4871 4886
rect 4875 4882 4959 4886
rect 4963 4882 5095 4886
rect 5099 4882 5183 4886
rect 5187 4882 5327 4886
rect 5331 4882 5407 4886
rect 5411 4882 5663 4886
rect 5667 4882 5695 4886
rect 3817 4881 5695 4882
rect 5701 4881 5702 4887
rect 96 4857 97 4863
rect 103 4862 1959 4863
rect 103 4858 111 4862
rect 115 4858 131 4862
rect 135 4858 267 4862
rect 271 4858 315 4862
rect 319 4858 403 4862
rect 407 4858 523 4862
rect 527 4858 539 4862
rect 543 4858 675 4862
rect 679 4858 723 4862
rect 727 4858 915 4862
rect 919 4858 1099 4862
rect 1103 4858 1283 4862
rect 1287 4858 1459 4862
rect 1463 4858 1635 4862
rect 1639 4858 1787 4862
rect 1791 4858 1935 4862
rect 1939 4858 1959 4862
rect 103 4857 1959 4858
rect 1965 4857 1966 4863
rect 1958 4805 1959 4811
rect 1965 4810 3823 4811
rect 1965 4806 1975 4810
rect 1979 4806 1995 4810
rect 1999 4806 2155 4810
rect 2159 4806 2347 4810
rect 2351 4806 2539 4810
rect 2543 4806 2731 4810
rect 2735 4806 2843 4810
rect 2847 4806 2931 4810
rect 2935 4806 2979 4810
rect 2983 4806 3131 4810
rect 3135 4806 3799 4810
rect 3803 4806 3823 4810
rect 1965 4805 3823 4806
rect 3829 4805 3830 4811
rect 3822 4765 3823 4771
rect 3829 4770 5707 4771
rect 3829 4766 3839 4770
rect 3843 4766 3859 4770
rect 3863 4766 3915 4770
rect 3919 4766 4043 4770
rect 4047 4766 4187 4770
rect 4191 4766 4259 4770
rect 4263 4766 4467 4770
rect 4471 4766 4483 4770
rect 4487 4766 4707 4770
rect 4711 4766 4763 4770
rect 4767 4766 4931 4770
rect 4935 4766 5067 4770
rect 5071 4766 5155 4770
rect 5159 4766 5371 4770
rect 5375 4766 5379 4770
rect 5383 4766 5663 4770
rect 5667 4766 5707 4770
rect 3829 4765 5707 4766
rect 5713 4765 5714 4771
rect 84 4737 85 4743
rect 91 4742 1947 4743
rect 91 4738 111 4742
rect 115 4738 159 4742
rect 163 4738 295 4742
rect 299 4738 343 4742
rect 347 4738 431 4742
rect 435 4738 567 4742
rect 571 4738 703 4742
rect 707 4738 807 4742
rect 811 4738 1055 4742
rect 1059 4738 1311 4742
rect 1315 4738 1575 4742
rect 1579 4738 1815 4742
rect 1819 4738 1935 4742
rect 1939 4738 1947 4742
rect 91 4737 1947 4738
rect 1953 4737 1954 4743
rect 1946 4689 1947 4695
rect 1953 4694 3811 4695
rect 1953 4690 1975 4694
rect 1979 4690 2023 4694
rect 2027 4690 2183 4694
rect 2187 4690 2239 4694
rect 2243 4690 2375 4694
rect 2379 4690 2471 4694
rect 2475 4690 2567 4694
rect 2571 4690 2695 4694
rect 2699 4690 2759 4694
rect 2763 4690 2919 4694
rect 2923 4690 2959 4694
rect 2963 4690 3143 4694
rect 3147 4690 3159 4694
rect 3163 4690 3367 4694
rect 3371 4690 3799 4694
rect 3803 4690 3811 4694
rect 1953 4689 3811 4690
rect 3817 4689 3818 4695
rect 3810 4653 3811 4659
rect 3817 4658 5695 4659
rect 3817 4654 3839 4658
rect 3843 4654 3943 4658
rect 3947 4654 4063 4658
rect 4067 4654 4215 4658
rect 4219 4654 4327 4658
rect 4331 4654 4495 4658
rect 4499 4654 4599 4658
rect 4603 4654 4791 4658
rect 4795 4654 4871 4658
rect 4875 4654 5095 4658
rect 5099 4654 5151 4658
rect 5155 4654 5399 4658
rect 5403 4654 5439 4658
rect 5443 4654 5663 4658
rect 5667 4654 5695 4658
rect 3817 4653 5695 4654
rect 5701 4653 5702 4659
rect 96 4609 97 4615
rect 103 4614 1959 4615
rect 103 4610 111 4614
rect 115 4610 131 4614
rect 135 4610 171 4614
rect 175 4610 315 4614
rect 319 4610 395 4614
rect 399 4610 539 4614
rect 543 4610 643 4614
rect 647 4610 779 4614
rect 783 4610 907 4614
rect 911 4610 1027 4614
rect 1031 4610 1195 4614
rect 1199 4610 1283 4614
rect 1287 4610 1491 4614
rect 1495 4610 1547 4614
rect 1551 4610 1787 4614
rect 1791 4610 1935 4614
rect 1939 4610 1959 4614
rect 103 4609 1959 4610
rect 1965 4609 1966 4615
rect 1958 4573 1959 4579
rect 1965 4578 3823 4579
rect 1965 4574 1975 4578
rect 1979 4574 1995 4578
rect 1999 4574 2099 4578
rect 2103 4574 2211 4578
rect 2215 4574 2347 4578
rect 2351 4574 2443 4578
rect 2447 4574 2579 4578
rect 2583 4574 2667 4578
rect 2671 4574 2795 4578
rect 2799 4574 2891 4578
rect 2895 4574 3003 4578
rect 3007 4574 3115 4578
rect 3119 4574 3203 4578
rect 3207 4574 3339 4578
rect 3343 4574 3403 4578
rect 3407 4574 3611 4578
rect 3615 4574 3799 4578
rect 3803 4574 3823 4578
rect 1965 4573 3823 4574
rect 3829 4573 3830 4579
rect 3822 4541 3823 4547
rect 3829 4546 5707 4547
rect 3829 4542 3839 4546
rect 3843 4542 4035 4546
rect 4039 4542 4179 4546
rect 4183 4542 4299 4546
rect 4303 4542 4411 4546
rect 4415 4542 4571 4546
rect 4575 4542 4659 4546
rect 4663 4542 4843 4546
rect 4847 4542 4915 4546
rect 4919 4542 5123 4546
rect 5127 4542 5179 4546
rect 5183 4542 5411 4546
rect 5415 4542 5443 4546
rect 5447 4542 5663 4546
rect 5667 4542 5707 4546
rect 3829 4541 5707 4542
rect 5713 4541 5714 4547
rect 84 4493 85 4499
rect 91 4498 1947 4499
rect 91 4494 111 4498
rect 115 4494 199 4498
rect 203 4494 423 4498
rect 427 4494 447 4498
rect 451 4494 655 4498
rect 659 4494 671 4498
rect 675 4494 887 4498
rect 891 4494 935 4498
rect 939 4494 1143 4498
rect 1147 4494 1223 4498
rect 1227 4494 1407 4498
rect 1411 4494 1519 4498
rect 1523 4494 1679 4498
rect 1683 4494 1815 4498
rect 1819 4494 1935 4498
rect 1939 4494 1947 4498
rect 91 4493 1947 4494
rect 1953 4493 1954 4499
rect 1946 4453 1947 4459
rect 1953 4458 3811 4459
rect 1953 4454 1975 4458
rect 1979 4454 2127 4458
rect 2131 4454 2231 4458
rect 2235 4454 2375 4458
rect 2379 4454 2447 4458
rect 2451 4454 2607 4458
rect 2611 4454 2663 4458
rect 2667 4454 2823 4458
rect 2827 4454 2871 4458
rect 2875 4454 3031 4458
rect 3035 4454 3079 4458
rect 3083 4454 3231 4458
rect 3235 4454 3287 4458
rect 3291 4454 3431 4458
rect 3435 4454 3495 4458
rect 3499 4454 3639 4458
rect 3643 4454 3679 4458
rect 3683 4454 3799 4458
rect 3803 4454 3811 4458
rect 1953 4453 3811 4454
rect 3817 4453 3818 4459
rect 3810 4421 3811 4427
rect 3817 4426 5695 4427
rect 3817 4422 3839 4426
rect 3843 4422 4207 4426
rect 4211 4422 4359 4426
rect 4363 4422 4439 4426
rect 4443 4422 4519 4426
rect 4523 4422 4687 4426
rect 4691 4422 4879 4426
rect 4883 4422 4943 4426
rect 4947 4422 5079 4426
rect 5083 4422 5207 4426
rect 5211 4422 5287 4426
rect 5291 4422 5471 4426
rect 5475 4422 5503 4426
rect 5507 4422 5663 4426
rect 5667 4422 5695 4426
rect 3817 4421 5695 4422
rect 5701 4421 5702 4427
rect 96 4377 97 4383
rect 103 4382 1959 4383
rect 103 4378 111 4382
rect 115 4378 419 4382
rect 423 4378 627 4382
rect 631 4378 667 4382
rect 671 4378 811 4382
rect 815 4378 859 4382
rect 863 4378 963 4382
rect 967 4378 1115 4382
rect 1119 4378 1123 4382
rect 1127 4378 1291 4382
rect 1295 4378 1379 4382
rect 1383 4378 1467 4382
rect 1471 4378 1651 4382
rect 1655 4378 1935 4382
rect 1939 4378 1959 4382
rect 103 4377 1959 4378
rect 1965 4377 1966 4383
rect 1958 4333 1959 4339
rect 1965 4338 3823 4339
rect 1965 4334 1975 4338
rect 1979 4334 2203 4338
rect 2207 4334 2307 4338
rect 2311 4334 2419 4338
rect 2423 4334 2459 4338
rect 2463 4334 2627 4338
rect 2631 4334 2635 4338
rect 2639 4334 2811 4338
rect 2815 4334 2843 4338
rect 2847 4334 3011 4338
rect 3015 4334 3051 4338
rect 3055 4334 3227 4338
rect 3231 4334 3259 4338
rect 3263 4334 3451 4338
rect 3455 4334 3467 4338
rect 3471 4334 3651 4338
rect 3655 4334 3799 4338
rect 3803 4334 3823 4338
rect 1965 4333 3823 4334
rect 3829 4333 3830 4339
rect 3822 4309 3823 4315
rect 3829 4314 5707 4315
rect 3829 4310 3839 4314
rect 3843 4310 3859 4314
rect 3863 4310 4043 4314
rect 4047 4310 4251 4314
rect 4255 4310 4331 4314
rect 4335 4310 4475 4314
rect 4479 4310 4491 4314
rect 4495 4310 4659 4314
rect 4663 4310 4715 4314
rect 4719 4310 4851 4314
rect 4855 4310 4971 4314
rect 4975 4310 5051 4314
rect 5055 4310 5235 4314
rect 5239 4310 5259 4314
rect 5263 4310 5475 4314
rect 5479 4310 5499 4314
rect 5503 4310 5663 4314
rect 5667 4310 5707 4314
rect 3829 4309 5707 4310
rect 5713 4309 5714 4315
rect 84 4249 85 4255
rect 91 4254 1947 4255
rect 91 4250 111 4254
rect 115 4250 695 4254
rect 699 4250 815 4254
rect 819 4250 839 4254
rect 843 4250 951 4254
rect 955 4250 991 4254
rect 995 4250 1087 4254
rect 1091 4250 1151 4254
rect 1155 4250 1223 4254
rect 1227 4250 1319 4254
rect 1323 4250 1359 4254
rect 1363 4250 1495 4254
rect 1499 4250 1631 4254
rect 1635 4250 1679 4254
rect 1683 4250 1767 4254
rect 1771 4250 1935 4254
rect 1939 4250 1947 4254
rect 91 4249 1947 4250
rect 1953 4249 1954 4255
rect 1946 4213 1947 4219
rect 1953 4218 3811 4219
rect 1953 4214 1975 4218
rect 1979 4214 2335 4218
rect 2339 4214 2487 4218
rect 2491 4214 2567 4218
rect 2571 4214 2655 4218
rect 2659 4214 2703 4218
rect 2707 4214 2839 4218
rect 2843 4214 2975 4218
rect 2979 4214 3039 4218
rect 3043 4214 3255 4218
rect 3259 4214 3479 4218
rect 3483 4214 3679 4218
rect 3683 4214 3799 4218
rect 3803 4214 3811 4218
rect 1953 4213 3811 4214
rect 3817 4213 3818 4219
rect 3810 4161 3811 4167
rect 3817 4166 5695 4167
rect 3817 4162 3839 4166
rect 3843 4162 3887 4166
rect 3891 4162 4071 4166
rect 4075 4162 4279 4166
rect 4283 4162 4415 4166
rect 4419 4162 4503 4166
rect 4507 4162 4743 4166
rect 4747 4162 4975 4166
rect 4979 4162 4999 4166
rect 5003 4162 5263 4166
rect 5267 4162 5527 4166
rect 5531 4162 5543 4166
rect 5547 4162 5663 4166
rect 5667 4162 5695 4166
rect 3817 4161 5695 4162
rect 5701 4161 5702 4167
rect 96 4133 97 4139
rect 103 4138 1959 4139
rect 103 4134 111 4138
rect 115 4134 731 4138
rect 735 4134 787 4138
rect 791 4134 867 4138
rect 871 4134 923 4138
rect 927 4134 1003 4138
rect 1007 4134 1059 4138
rect 1063 4134 1139 4138
rect 1143 4134 1195 4138
rect 1199 4134 1275 4138
rect 1279 4134 1331 4138
rect 1335 4134 1411 4138
rect 1415 4134 1467 4138
rect 1471 4134 1547 4138
rect 1551 4134 1603 4138
rect 1607 4134 1739 4138
rect 1743 4134 1935 4138
rect 1939 4134 1959 4138
rect 103 4133 1959 4134
rect 1965 4133 1966 4139
rect 1958 4081 1959 4087
rect 1965 4086 3823 4087
rect 1965 4082 1975 4086
rect 1979 4082 2291 4086
rect 2295 4082 2427 4086
rect 2431 4082 2539 4086
rect 2543 4082 2563 4086
rect 2567 4082 2675 4086
rect 2679 4082 2699 4086
rect 2703 4082 2811 4086
rect 2815 4082 2835 4086
rect 2839 4082 2947 4086
rect 2951 4082 3799 4086
rect 3803 4082 3823 4086
rect 1965 4081 3823 4082
rect 3829 4081 3830 4087
rect 2386 4052 2392 4053
rect 2958 4052 2964 4053
rect 2386 4048 2387 4052
rect 2391 4048 2959 4052
rect 2963 4048 2964 4052
rect 3822 4049 3823 4055
rect 3829 4054 5707 4055
rect 3829 4050 3839 4054
rect 3843 4050 3859 4054
rect 3863 4050 4003 4054
rect 4007 4050 4171 4054
rect 4175 4050 4339 4054
rect 4343 4050 4387 4054
rect 4391 4050 4499 4054
rect 4503 4050 4651 4054
rect 4655 4050 4803 4054
rect 4807 4050 4947 4054
rect 4951 4050 5091 4054
rect 5095 4050 5235 4054
rect 5239 4050 5379 4054
rect 5383 4050 5515 4054
rect 5519 4050 5663 4054
rect 5667 4050 5707 4054
rect 3829 4049 5707 4050
rect 5713 4049 5714 4055
rect 2386 4047 2392 4048
rect 2958 4047 2964 4048
rect 84 3997 85 4003
rect 91 4002 1947 4003
rect 91 3998 111 4002
rect 115 3998 511 4002
rect 515 3998 663 4002
rect 667 3998 759 4002
rect 763 3998 823 4002
rect 827 3998 895 4002
rect 899 3998 983 4002
rect 987 3998 1031 4002
rect 1035 3998 1151 4002
rect 1155 3998 1167 4002
rect 1171 3998 1303 4002
rect 1307 3998 1319 4002
rect 1323 3998 1439 4002
rect 1443 3998 1575 4002
rect 1579 3998 1935 4002
rect 1939 3998 1947 4002
rect 91 3997 1947 3998
rect 1953 3997 1954 4003
rect 1946 3965 1947 3971
rect 1953 3970 3811 3971
rect 1953 3966 1975 3970
rect 1979 3966 2119 3970
rect 2123 3966 2319 3970
rect 2323 3966 2327 3970
rect 2331 3966 2455 3970
rect 2459 3966 2535 3970
rect 2539 3966 2591 3970
rect 2595 3966 2727 3970
rect 2731 3966 2743 3970
rect 2747 3966 2863 3970
rect 2867 3966 2943 3970
rect 2947 3966 3135 3970
rect 3139 3966 3319 3970
rect 3323 3966 3511 3970
rect 3515 3966 3679 3970
rect 3683 3966 3799 3970
rect 3803 3966 3811 3970
rect 1953 3965 3811 3966
rect 3817 3965 3818 3971
rect 3810 3913 3811 3919
rect 3817 3918 5695 3919
rect 3817 3914 3839 3918
rect 3843 3914 3887 3918
rect 3891 3914 4031 3918
rect 4035 3914 4199 3918
rect 4203 3914 4367 3918
rect 4371 3914 4383 3918
rect 4387 3914 4527 3918
rect 4531 3914 4599 3918
rect 4603 3914 4679 3918
rect 4683 3914 4823 3918
rect 4827 3914 4831 3918
rect 4835 3914 4975 3918
rect 4979 3914 5063 3918
rect 5067 3914 5119 3918
rect 5123 3914 5263 3918
rect 5267 3914 5311 3918
rect 5315 3914 5407 3918
rect 5411 3914 5543 3918
rect 5547 3914 5663 3918
rect 5667 3914 5695 3918
rect 3817 3913 5695 3914
rect 5701 3913 5702 3919
rect 96 3857 97 3863
rect 103 3862 1959 3863
rect 103 3858 111 3862
rect 115 3858 131 3862
rect 135 3858 307 3862
rect 311 3858 483 3862
rect 487 3858 515 3862
rect 519 3858 635 3862
rect 639 3858 723 3862
rect 727 3858 795 3862
rect 799 3858 939 3862
rect 943 3858 955 3862
rect 959 3858 1123 3862
rect 1127 3858 1163 3862
rect 1167 3858 1291 3862
rect 1295 3858 1935 3862
rect 1939 3858 1959 3862
rect 103 3857 1959 3858
rect 1965 3857 1966 3863
rect 1958 3841 1959 3847
rect 1965 3846 3823 3847
rect 1965 3842 1975 3846
rect 1979 3842 2091 3846
rect 2095 3842 2139 3846
rect 2143 3842 2299 3846
rect 2303 3842 2371 3846
rect 2375 3842 2507 3846
rect 2511 3842 2587 3846
rect 2591 3842 2715 3846
rect 2719 3842 2795 3846
rect 2799 3842 2915 3846
rect 2919 3842 2995 3846
rect 2999 3842 3107 3846
rect 3111 3842 3195 3846
rect 3199 3842 3291 3846
rect 3295 3842 3403 3846
rect 3407 3842 3483 3846
rect 3487 3842 3651 3846
rect 3655 3842 3799 3846
rect 3803 3842 3823 3846
rect 1965 3841 3823 3842
rect 3829 3841 3830 3847
rect 3010 3828 3016 3829
rect 3418 3828 3424 3829
rect 3010 3824 3011 3828
rect 3015 3824 3419 3828
rect 3423 3824 3424 3828
rect 3010 3823 3016 3824
rect 3418 3823 3424 3824
rect 3822 3785 3823 3791
rect 3829 3790 5707 3791
rect 3829 3786 3839 3790
rect 3843 3786 3995 3790
rect 3999 3786 4203 3790
rect 4207 3786 4355 3790
rect 4359 3786 4435 3790
rect 4439 3786 4571 3790
rect 4575 3786 4691 3790
rect 4695 3786 4795 3790
rect 4799 3786 4963 3790
rect 4967 3786 5035 3790
rect 5039 3786 5251 3790
rect 5255 3786 5283 3790
rect 5287 3786 5515 3790
rect 5519 3786 5663 3790
rect 5667 3786 5707 3790
rect 3829 3785 5707 3786
rect 5713 3785 5714 3791
rect 84 3745 85 3751
rect 91 3750 1947 3751
rect 91 3746 111 3750
rect 115 3746 159 3750
rect 163 3746 335 3750
rect 339 3746 527 3750
rect 531 3746 543 3750
rect 547 3746 711 3750
rect 715 3746 751 3750
rect 755 3746 887 3750
rect 891 3746 967 3750
rect 971 3746 1055 3750
rect 1059 3746 1191 3750
rect 1195 3746 1215 3750
rect 1219 3746 1367 3750
rect 1371 3746 1519 3750
rect 1523 3746 1679 3750
rect 1683 3746 1815 3750
rect 1819 3746 1935 3750
rect 1939 3746 1947 3750
rect 91 3745 1947 3746
rect 1953 3745 1954 3751
rect 4090 3732 4096 3733
rect 4938 3732 4944 3733
rect 1946 3725 1947 3731
rect 1953 3730 3811 3731
rect 1953 3726 1975 3730
rect 1979 3726 2167 3730
rect 2171 3726 2279 3730
rect 2283 3726 2399 3730
rect 2403 3726 2479 3730
rect 2483 3726 2615 3730
rect 2619 3726 2679 3730
rect 2683 3726 2823 3730
rect 2827 3726 2879 3730
rect 2883 3726 3023 3730
rect 3027 3726 3079 3730
rect 3083 3726 3223 3730
rect 3227 3726 3279 3730
rect 3283 3726 3431 3730
rect 3435 3726 3799 3730
rect 3803 3726 3811 3730
rect 1953 3725 3811 3726
rect 3817 3725 3818 3731
rect 4090 3728 4091 3732
rect 4095 3728 4939 3732
rect 4943 3728 4944 3732
rect 4090 3727 4096 3728
rect 4938 3727 4944 3728
rect 3810 3645 3811 3651
rect 3817 3650 5695 3651
rect 3817 3646 3839 3650
rect 3843 3646 4023 3650
rect 4027 3646 4215 3650
rect 4219 3646 4231 3650
rect 4235 3646 4399 3650
rect 4403 3646 4463 3650
rect 4467 3646 4607 3650
rect 4611 3646 4719 3650
rect 4723 3646 4831 3650
rect 4835 3646 4991 3650
rect 4995 3646 5071 3650
rect 5075 3646 5279 3650
rect 5283 3646 5319 3650
rect 5323 3646 5543 3650
rect 5547 3646 5663 3650
rect 5667 3646 5695 3650
rect 3817 3645 5695 3646
rect 5701 3645 5702 3651
rect 96 3621 97 3627
rect 103 3626 1959 3627
rect 103 3622 111 3626
rect 115 3622 131 3626
rect 135 3622 147 3626
rect 151 3622 307 3626
rect 311 3622 355 3626
rect 359 3622 499 3626
rect 503 3622 571 3626
rect 575 3622 683 3626
rect 687 3622 803 3626
rect 807 3622 859 3626
rect 863 3622 1027 3626
rect 1031 3622 1043 3626
rect 1047 3622 1187 3626
rect 1191 3622 1291 3626
rect 1295 3622 1339 3626
rect 1343 3622 1491 3626
rect 1495 3622 1547 3626
rect 1551 3622 1651 3626
rect 1655 3622 1787 3626
rect 1791 3622 1935 3626
rect 1939 3622 1959 3626
rect 103 3621 1959 3622
rect 1965 3621 1966 3627
rect 1958 3601 1959 3607
rect 1965 3606 3823 3607
rect 1965 3602 1975 3606
rect 1979 3602 1995 3606
rect 1999 3602 2251 3606
rect 2255 3602 2451 3606
rect 2455 3602 2515 3606
rect 2519 3602 2651 3606
rect 2655 3602 2755 3606
rect 2759 3602 2851 3606
rect 2855 3602 2979 3606
rect 2983 3602 3051 3606
rect 3055 3602 3195 3606
rect 3199 3602 3251 3606
rect 3255 3602 3411 3606
rect 3415 3602 3627 3606
rect 3631 3602 3799 3606
rect 3803 3602 3823 3606
rect 1965 3601 3823 3602
rect 3829 3601 3830 3607
rect 3822 3509 3823 3515
rect 3829 3514 5707 3515
rect 3829 3510 3839 3514
rect 3843 3510 4187 3514
rect 4191 3510 4371 3514
rect 4375 3510 4531 3514
rect 4535 3510 4579 3514
rect 4583 3510 4683 3514
rect 4687 3510 4803 3514
rect 4807 3510 4843 3514
rect 4847 3510 5003 3514
rect 5007 3510 5043 3514
rect 5047 3510 5171 3514
rect 5175 3510 5291 3514
rect 5295 3510 5347 3514
rect 5351 3510 5515 3514
rect 5519 3510 5663 3514
rect 5667 3510 5707 3514
rect 3829 3509 5707 3510
rect 5713 3509 5714 3515
rect 84 3485 85 3491
rect 91 3490 1947 3491
rect 91 3486 111 3490
rect 115 3486 175 3490
rect 179 3486 303 3490
rect 307 3486 383 3490
rect 387 3486 447 3490
rect 451 3486 599 3490
rect 603 3486 759 3490
rect 763 3486 831 3490
rect 835 3486 935 3490
rect 939 3486 1071 3490
rect 1075 3486 1111 3490
rect 1115 3486 1295 3490
rect 1299 3486 1319 3490
rect 1323 3486 1487 3490
rect 1491 3486 1575 3490
rect 1579 3486 1815 3490
rect 1819 3486 1935 3490
rect 1939 3486 1947 3490
rect 91 3485 1947 3486
rect 1953 3487 1954 3491
rect 1953 3486 3818 3487
rect 1953 3485 1975 3486
rect 1946 3482 1975 3485
rect 1979 3482 2023 3486
rect 2027 3482 2191 3486
rect 2195 3482 2279 3486
rect 2283 3482 2399 3486
rect 2403 3482 2543 3486
rect 2547 3482 2615 3486
rect 2619 3482 2783 3486
rect 2787 3482 2831 3486
rect 2835 3482 3007 3486
rect 3011 3482 3047 3486
rect 3051 3482 3223 3486
rect 3227 3482 3263 3486
rect 3267 3482 3439 3486
rect 3443 3482 3479 3486
rect 3483 3482 3655 3486
rect 3659 3482 3679 3486
rect 3683 3482 3799 3486
rect 3803 3482 3818 3486
rect 1946 3481 3818 3482
rect 3810 3393 3811 3399
rect 3817 3398 5695 3399
rect 3817 3394 3839 3398
rect 3843 3394 3887 3398
rect 3891 3394 4151 3398
rect 4155 3394 4423 3398
rect 4427 3394 4559 3398
rect 4563 3394 4671 3398
rect 4675 3394 4711 3398
rect 4715 3394 4871 3398
rect 4875 3394 4895 3398
rect 4899 3394 5031 3398
rect 5035 3394 5111 3398
rect 5115 3394 5199 3398
rect 5203 3394 5327 3398
rect 5331 3394 5375 3398
rect 5379 3394 5543 3398
rect 5547 3394 5663 3398
rect 5667 3394 5695 3398
rect 3817 3393 5695 3394
rect 5701 3393 5702 3399
rect 96 3357 97 3363
rect 103 3362 1959 3363
rect 103 3358 111 3362
rect 115 3358 275 3362
rect 279 3358 419 3362
rect 423 3358 467 3362
rect 471 3358 571 3362
rect 575 3358 667 3362
rect 671 3358 731 3362
rect 735 3358 875 3362
rect 879 3358 907 3362
rect 911 3358 1083 3362
rect 1087 3358 1091 3362
rect 1095 3358 1267 3362
rect 1271 3358 1315 3362
rect 1319 3358 1459 3362
rect 1463 3358 1935 3362
rect 1939 3358 1959 3362
rect 103 3357 1959 3358
rect 1965 3357 1966 3363
rect 1958 3329 1959 3335
rect 1965 3334 3823 3335
rect 1965 3330 1975 3334
rect 1979 3330 1995 3334
rect 1999 3330 2163 3334
rect 2167 3330 2195 3334
rect 2199 3330 2371 3334
rect 2375 3330 2411 3334
rect 2415 3330 2587 3334
rect 2591 3330 2619 3334
rect 2623 3330 2803 3334
rect 2807 3330 2811 3334
rect 2815 3330 3003 3334
rect 3007 3330 3019 3334
rect 3023 3330 3187 3334
rect 3191 3330 3235 3334
rect 3239 3330 3371 3334
rect 3375 3330 3451 3334
rect 3455 3330 3555 3334
rect 3559 3330 3651 3334
rect 3655 3330 3799 3334
rect 3803 3330 3823 3334
rect 1965 3329 3823 3330
rect 3829 3329 3830 3335
rect 3822 3281 3823 3287
rect 3829 3286 5707 3287
rect 3829 3282 3839 3286
rect 3843 3282 3859 3286
rect 3863 3282 4099 3286
rect 4103 3282 4123 3286
rect 4127 3282 4347 3286
rect 4351 3282 4395 3286
rect 4399 3282 4579 3286
rect 4583 3282 4643 3286
rect 4647 3282 4787 3286
rect 4791 3282 4867 3286
rect 4871 3282 4987 3286
rect 4991 3282 5083 3286
rect 5087 3282 5171 3286
rect 5175 3282 5299 3286
rect 5303 3282 5355 3286
rect 5359 3282 5515 3286
rect 5519 3282 5663 3286
rect 5667 3282 5707 3286
rect 3829 3281 5707 3282
rect 5713 3281 5714 3287
rect 84 3245 85 3251
rect 91 3250 1947 3251
rect 91 3246 111 3250
rect 115 3246 495 3250
rect 499 3246 535 3250
rect 539 3246 695 3250
rect 699 3246 727 3250
rect 731 3246 903 3250
rect 907 3246 919 3250
rect 923 3246 1111 3250
rect 1115 3246 1119 3250
rect 1123 3246 1295 3250
rect 1299 3246 1343 3250
rect 1347 3246 1471 3250
rect 1475 3246 1655 3250
rect 1659 3246 1815 3250
rect 1819 3246 1935 3250
rect 1939 3246 1947 3250
rect 91 3245 1947 3246
rect 1953 3245 1954 3251
rect 1946 3217 1947 3223
rect 1953 3222 3811 3223
rect 1953 3218 1975 3222
rect 1979 3218 2023 3222
rect 2027 3218 2223 3222
rect 2227 3218 2439 3222
rect 2443 3218 2463 3222
rect 2467 3218 2647 3222
rect 2651 3218 2663 3222
rect 2667 3218 2839 3222
rect 2843 3218 2863 3222
rect 2867 3218 3031 3222
rect 3035 3218 3055 3222
rect 3059 3218 3215 3222
rect 3219 3218 3239 3222
rect 3243 3218 3399 3222
rect 3403 3218 3431 3222
rect 3435 3218 3583 3222
rect 3587 3218 3623 3222
rect 3627 3218 3799 3222
rect 3803 3218 3811 3222
rect 1953 3217 3811 3218
rect 3817 3217 3818 3223
rect 3810 3153 3811 3159
rect 3817 3158 5695 3159
rect 3817 3154 3839 3158
rect 3843 3154 3887 3158
rect 3891 3154 3903 3158
rect 3907 3154 4127 3158
rect 4131 3154 4135 3158
rect 4139 3154 4359 3158
rect 4363 3154 4375 3158
rect 4379 3154 4583 3158
rect 4587 3154 4607 3158
rect 4611 3154 4807 3158
rect 4811 3154 4815 3158
rect 4819 3154 5015 3158
rect 5019 3154 5031 3158
rect 5035 3154 5199 3158
rect 5203 3154 5383 3158
rect 5387 3154 5543 3158
rect 5547 3154 5663 3158
rect 5667 3154 5695 3158
rect 3817 3153 5695 3154
rect 5701 3153 5702 3159
rect 96 3125 97 3131
rect 103 3130 1959 3131
rect 103 3126 111 3130
rect 115 3126 427 3130
rect 431 3126 507 3130
rect 511 3126 563 3130
rect 567 3126 699 3130
rect 703 3126 835 3130
rect 839 3126 891 3130
rect 895 3126 971 3130
rect 975 3126 1083 3130
rect 1087 3126 1107 3130
rect 1111 3126 1243 3130
rect 1247 3126 1267 3130
rect 1271 3126 1379 3130
rect 1383 3126 1443 3130
rect 1447 3126 1515 3130
rect 1519 3126 1627 3130
rect 1631 3126 1651 3130
rect 1655 3126 1787 3130
rect 1791 3126 1935 3130
rect 1939 3126 1959 3130
rect 103 3125 1959 3126
rect 1965 3125 1966 3131
rect 1958 3093 1959 3099
rect 1965 3098 3823 3099
rect 1965 3094 1975 3098
rect 1979 3094 2331 3098
rect 2335 3094 2435 3098
rect 2439 3094 2555 3098
rect 2559 3094 2635 3098
rect 2639 3094 2779 3098
rect 2783 3094 2835 3098
rect 2839 3094 3003 3098
rect 3007 3094 3027 3098
rect 3031 3094 3211 3098
rect 3215 3094 3235 3098
rect 3239 3094 3403 3098
rect 3407 3094 3467 3098
rect 3471 3094 3595 3098
rect 3599 3094 3799 3098
rect 3803 3094 3823 3098
rect 1965 3093 3823 3094
rect 3829 3093 3830 3099
rect 3822 3041 3823 3047
rect 3829 3046 5707 3047
rect 3829 3042 3839 3046
rect 3843 3042 3875 3046
rect 3879 3042 3907 3046
rect 3911 3042 4075 3046
rect 4079 3042 4107 3046
rect 4111 3042 4243 3046
rect 4247 3042 4331 3046
rect 4335 3042 4411 3046
rect 4415 3042 4555 3046
rect 4559 3042 4579 3046
rect 4583 3042 4755 3046
rect 4759 3042 4779 3046
rect 4783 3042 5003 3046
rect 5007 3042 5663 3046
rect 5667 3042 5707 3046
rect 3829 3041 5707 3042
rect 5713 3041 5714 3047
rect 84 2985 85 2991
rect 91 2990 1947 2991
rect 91 2986 111 2990
rect 115 2986 199 2990
rect 203 2986 455 2990
rect 459 2986 511 2990
rect 515 2986 591 2990
rect 595 2986 727 2990
rect 731 2986 815 2990
rect 819 2986 863 2990
rect 867 2986 999 2990
rect 1003 2986 1111 2990
rect 1115 2986 1135 2990
rect 1139 2986 1271 2990
rect 1275 2986 1407 2990
rect 1411 2986 1415 2990
rect 1419 2986 1543 2990
rect 1547 2986 1679 2990
rect 1683 2986 1719 2990
rect 1723 2986 1815 2990
rect 1819 2986 1935 2990
rect 1939 2986 1947 2990
rect 91 2985 1947 2986
rect 1953 2985 1954 2991
rect 1946 2969 1947 2975
rect 1953 2974 3811 2975
rect 1953 2970 1975 2974
rect 1979 2970 2143 2974
rect 2147 2970 2343 2974
rect 2347 2970 2359 2974
rect 2363 2970 2543 2974
rect 2547 2970 2583 2974
rect 2587 2970 2743 2974
rect 2747 2970 2807 2974
rect 2811 2970 2935 2974
rect 2939 2970 3031 2974
rect 3035 2970 3135 2974
rect 3139 2970 3263 2974
rect 3267 2970 3335 2974
rect 3339 2970 3495 2974
rect 3499 2970 3799 2974
rect 3803 2970 3811 2974
rect 1953 2969 3811 2970
rect 3817 2969 3818 2975
rect 3810 2925 3811 2931
rect 3817 2930 5695 2931
rect 3817 2926 3839 2930
rect 3843 2926 3895 2930
rect 3899 2926 3935 2930
rect 3939 2926 4031 2930
rect 4035 2926 4103 2930
rect 4107 2926 4167 2930
rect 4171 2926 4271 2930
rect 4275 2926 4303 2930
rect 4307 2926 4439 2930
rect 4443 2926 4575 2930
rect 4579 2926 4607 2930
rect 4611 2926 4783 2930
rect 4787 2926 5663 2930
rect 5667 2926 5695 2930
rect 3817 2925 5695 2926
rect 5701 2925 5702 2931
rect 96 2873 97 2879
rect 103 2878 1959 2879
rect 103 2874 111 2878
rect 115 2874 131 2878
rect 135 2874 171 2878
rect 175 2874 307 2878
rect 311 2874 483 2878
rect 487 2874 523 2878
rect 527 2874 763 2878
rect 767 2874 787 2878
rect 791 2874 1011 2878
rect 1015 2874 1083 2878
rect 1087 2874 1275 2878
rect 1279 2874 1387 2878
rect 1391 2874 1539 2878
rect 1543 2874 1691 2878
rect 1695 2874 1935 2878
rect 1939 2874 1959 2878
rect 103 2873 1959 2874
rect 1965 2873 1966 2879
rect 1958 2849 1959 2855
rect 1965 2854 3823 2855
rect 1965 2850 1975 2854
rect 1979 2850 2011 2854
rect 2015 2850 2115 2854
rect 2119 2850 2259 2854
rect 2263 2850 2315 2854
rect 2319 2850 2507 2854
rect 2511 2850 2515 2854
rect 2519 2850 2715 2854
rect 2719 2850 2755 2854
rect 2759 2850 2907 2854
rect 2911 2850 3003 2854
rect 3007 2850 3107 2854
rect 3111 2850 3307 2854
rect 3311 2850 3799 2854
rect 3803 2850 3823 2854
rect 1965 2849 3823 2850
rect 3829 2849 3830 2855
rect 3822 2805 3823 2811
rect 3829 2810 5707 2811
rect 3829 2806 3839 2810
rect 3843 2806 3859 2810
rect 3863 2806 3867 2810
rect 3871 2806 3995 2810
rect 3999 2806 4003 2810
rect 4007 2806 4131 2810
rect 4135 2806 4139 2810
rect 4143 2806 4267 2810
rect 4271 2806 4275 2810
rect 4279 2806 4403 2810
rect 4407 2806 4411 2810
rect 4415 2806 4539 2810
rect 4543 2806 4547 2810
rect 4551 2806 4675 2810
rect 4679 2806 4811 2810
rect 4815 2806 5663 2810
rect 5667 2806 5707 2810
rect 3829 2805 5707 2806
rect 5713 2805 5714 2811
rect 84 2757 85 2763
rect 91 2762 1947 2763
rect 91 2758 111 2762
rect 115 2758 159 2762
rect 163 2758 279 2762
rect 283 2758 335 2762
rect 339 2758 455 2762
rect 459 2758 551 2762
rect 555 2758 647 2762
rect 651 2758 791 2762
rect 795 2758 855 2762
rect 859 2758 1039 2762
rect 1043 2758 1079 2762
rect 1083 2758 1303 2762
rect 1307 2758 1311 2762
rect 1315 2758 1551 2762
rect 1555 2758 1567 2762
rect 1571 2758 1799 2762
rect 1803 2758 1935 2762
rect 1939 2758 1947 2762
rect 91 2757 1947 2758
rect 1953 2757 1954 2763
rect 1946 2733 1947 2739
rect 1953 2738 3811 2739
rect 1953 2734 1975 2738
rect 1979 2734 2023 2738
rect 2027 2734 2039 2738
rect 2043 2734 2247 2738
rect 2251 2734 2287 2738
rect 2291 2734 2503 2738
rect 2507 2734 2535 2738
rect 2539 2734 2759 2738
rect 2763 2734 2783 2738
rect 2787 2734 3015 2738
rect 3019 2734 3031 2738
rect 3035 2734 3799 2738
rect 3803 2734 3811 2738
rect 1953 2733 3811 2734
rect 3817 2733 3818 2739
rect 3810 2693 3811 2699
rect 3817 2698 5695 2699
rect 3817 2694 3839 2698
rect 3843 2694 3887 2698
rect 3891 2694 3959 2698
rect 3963 2694 4023 2698
rect 4027 2694 4159 2698
rect 4163 2694 4255 2698
rect 4259 2694 4295 2698
rect 4299 2694 4431 2698
rect 4435 2694 4543 2698
rect 4547 2694 4567 2698
rect 4571 2694 4703 2698
rect 4707 2694 4823 2698
rect 4827 2694 4839 2698
rect 4843 2694 5111 2698
rect 5115 2694 5399 2698
rect 5403 2694 5663 2698
rect 5667 2694 5695 2698
rect 3817 2693 5695 2694
rect 5701 2693 5702 2699
rect 96 2645 97 2651
rect 103 2650 1959 2651
rect 103 2646 111 2650
rect 115 2646 251 2650
rect 255 2646 427 2650
rect 431 2646 571 2650
rect 575 2646 619 2650
rect 623 2646 731 2650
rect 735 2646 827 2650
rect 831 2646 891 2650
rect 895 2646 1043 2650
rect 1047 2646 1051 2650
rect 1055 2646 1195 2650
rect 1199 2646 1283 2650
rect 1287 2646 1355 2650
rect 1359 2646 1515 2650
rect 1519 2646 1523 2650
rect 1527 2646 1675 2650
rect 1679 2646 1771 2650
rect 1775 2646 1935 2650
rect 1939 2646 1959 2650
rect 103 2645 1959 2646
rect 1965 2645 1966 2651
rect 1958 2609 1959 2615
rect 1965 2614 3823 2615
rect 1965 2610 1975 2614
rect 1979 2610 1995 2614
rect 1999 2610 2219 2614
rect 2223 2610 2475 2614
rect 2479 2610 2555 2614
rect 2559 2610 2691 2614
rect 2695 2610 2731 2614
rect 2735 2610 2827 2614
rect 2831 2610 2963 2614
rect 2967 2610 2987 2614
rect 2991 2610 3099 2614
rect 3103 2610 3799 2614
rect 3803 2610 3823 2614
rect 1965 2609 3823 2610
rect 3829 2609 3830 2615
rect 3822 2581 3823 2587
rect 3829 2586 5707 2587
rect 3829 2582 3839 2586
rect 3843 2582 3859 2586
rect 3863 2582 3931 2586
rect 3935 2582 4083 2586
rect 4087 2582 4227 2586
rect 4231 2582 4331 2586
rect 4335 2582 4515 2586
rect 4519 2582 4579 2586
rect 4583 2582 4795 2586
rect 4799 2582 4827 2586
rect 4831 2582 5075 2586
rect 5079 2582 5083 2586
rect 5087 2582 5323 2586
rect 5327 2582 5371 2586
rect 5375 2582 5663 2586
rect 5667 2582 5707 2586
rect 3829 2581 5707 2582
rect 5713 2581 5714 2587
rect 84 2533 85 2539
rect 91 2538 1947 2539
rect 91 2534 111 2538
rect 115 2534 383 2538
rect 387 2534 599 2538
rect 603 2534 759 2538
rect 763 2534 815 2538
rect 819 2534 919 2538
rect 923 2534 1023 2538
rect 1027 2534 1071 2538
rect 1075 2534 1223 2538
rect 1227 2534 1231 2538
rect 1235 2534 1383 2538
rect 1387 2534 1431 2538
rect 1435 2534 1543 2538
rect 1547 2534 1631 2538
rect 1635 2534 1703 2538
rect 1707 2534 1815 2538
rect 1819 2534 1935 2538
rect 1939 2534 1947 2538
rect 91 2533 1947 2534
rect 1953 2533 1954 2539
rect 1946 2473 1947 2479
rect 1953 2478 3811 2479
rect 1953 2474 1975 2478
rect 1979 2474 2023 2478
rect 2027 2474 2223 2478
rect 2227 2474 2447 2478
rect 2451 2474 2583 2478
rect 2587 2474 2679 2478
rect 2683 2474 2719 2478
rect 2723 2474 2855 2478
rect 2859 2474 2927 2478
rect 2931 2474 2991 2478
rect 2995 2474 3127 2478
rect 3131 2474 3183 2478
rect 3187 2474 3439 2478
rect 3443 2474 3679 2478
rect 3683 2474 3799 2478
rect 3803 2474 3811 2478
rect 1953 2473 3811 2474
rect 3817 2473 3818 2479
rect 3810 2471 3818 2473
rect 3810 2465 3811 2471
rect 3817 2470 5695 2471
rect 3817 2466 3839 2470
rect 3843 2466 3887 2470
rect 3891 2466 4087 2470
rect 4091 2466 4111 2470
rect 4115 2466 4327 2470
rect 4331 2466 4359 2470
rect 4363 2466 4583 2470
rect 4587 2466 4607 2470
rect 4611 2466 4847 2470
rect 4851 2466 4855 2470
rect 4859 2466 5103 2470
rect 5107 2466 5119 2470
rect 5123 2466 5351 2470
rect 5355 2466 5399 2470
rect 5403 2466 5663 2470
rect 5667 2466 5695 2470
rect 3817 2465 5695 2466
rect 5701 2465 5702 2471
rect 96 2417 97 2423
rect 103 2422 1959 2423
rect 103 2418 111 2422
rect 115 2418 227 2422
rect 231 2418 355 2422
rect 359 2418 523 2422
rect 527 2418 571 2422
rect 575 2418 787 2422
rect 791 2418 835 2422
rect 839 2418 995 2422
rect 999 2418 1155 2422
rect 1159 2418 1203 2422
rect 1207 2418 1403 2422
rect 1407 2418 1483 2422
rect 1487 2418 1603 2422
rect 1607 2418 1787 2422
rect 1791 2418 1935 2422
rect 1939 2418 1959 2422
rect 103 2417 1959 2418
rect 1965 2417 1966 2423
rect 1958 2353 1959 2359
rect 1965 2358 3823 2359
rect 1965 2354 1975 2358
rect 1979 2354 1995 2358
rect 1999 2354 2155 2358
rect 2159 2354 2195 2358
rect 2199 2354 2347 2358
rect 2351 2354 2419 2358
rect 2423 2354 2539 2358
rect 2543 2354 2651 2358
rect 2655 2354 2731 2358
rect 2735 2354 2899 2358
rect 2903 2354 2923 2358
rect 2927 2354 3115 2358
rect 3119 2354 3155 2358
rect 3159 2354 3299 2358
rect 3303 2354 3411 2358
rect 3415 2354 3483 2358
rect 3487 2354 3651 2358
rect 3655 2354 3799 2358
rect 3803 2354 3823 2358
rect 1965 2353 3823 2354
rect 3829 2353 3830 2359
rect 3822 2341 3823 2347
rect 3829 2346 5707 2347
rect 3829 2342 3839 2346
rect 3843 2342 3859 2346
rect 3863 2342 4059 2346
rect 4063 2342 4299 2346
rect 4303 2342 4443 2346
rect 4447 2342 4555 2346
rect 4559 2342 4611 2346
rect 4615 2342 4787 2346
rect 4791 2342 4819 2346
rect 4823 2342 4963 2346
rect 4967 2342 5091 2346
rect 5095 2342 5147 2346
rect 5151 2342 5339 2346
rect 5343 2342 5371 2346
rect 5375 2342 5515 2346
rect 5519 2342 5663 2346
rect 5667 2342 5707 2346
rect 3829 2341 5707 2342
rect 5713 2341 5714 2347
rect 84 2289 85 2295
rect 91 2294 1947 2295
rect 91 2290 111 2294
rect 115 2290 159 2294
rect 163 2290 255 2294
rect 259 2290 367 2294
rect 371 2290 551 2294
rect 555 2290 599 2294
rect 603 2290 831 2294
rect 835 2290 863 2294
rect 867 2290 1063 2294
rect 1067 2290 1183 2294
rect 1187 2290 1511 2294
rect 1515 2290 1815 2294
rect 1819 2290 1935 2294
rect 1939 2290 1947 2294
rect 91 2289 1947 2290
rect 1953 2289 1954 2295
rect 1946 2233 1947 2239
rect 1953 2238 3811 2239
rect 1953 2234 1975 2238
rect 1979 2234 2023 2238
rect 2027 2234 2183 2238
rect 2187 2234 2191 2238
rect 2195 2234 2359 2238
rect 2363 2234 2375 2238
rect 2379 2234 2535 2238
rect 2539 2234 2567 2238
rect 2571 2234 2711 2238
rect 2715 2234 2759 2238
rect 2763 2234 2879 2238
rect 2883 2234 2951 2238
rect 2955 2234 3047 2238
rect 3051 2234 3143 2238
rect 3147 2234 3207 2238
rect 3211 2234 3327 2238
rect 3331 2234 3367 2238
rect 3371 2234 3511 2238
rect 3515 2234 3535 2238
rect 3539 2234 3679 2238
rect 3683 2234 3799 2238
rect 3803 2234 3811 2238
rect 1953 2233 3811 2234
rect 3817 2233 3818 2239
rect 3810 2217 3811 2223
rect 3817 2222 5695 2223
rect 3817 2218 3839 2222
rect 3843 2218 4471 2222
rect 4475 2218 4543 2222
rect 4547 2218 4639 2222
rect 4643 2218 4719 2222
rect 4723 2218 4815 2222
rect 4819 2218 4911 2222
rect 4915 2218 4991 2222
rect 4995 2218 5119 2222
rect 5123 2218 5175 2222
rect 5179 2218 5335 2222
rect 5339 2218 5367 2222
rect 5371 2218 5543 2222
rect 5547 2218 5663 2222
rect 5667 2218 5695 2222
rect 3817 2217 5695 2218
rect 5701 2217 5702 2223
rect 96 2165 97 2171
rect 103 2170 1959 2171
rect 103 2166 111 2170
rect 115 2166 131 2170
rect 135 2166 339 2170
rect 343 2166 347 2170
rect 351 2166 571 2170
rect 575 2166 595 2170
rect 599 2166 803 2170
rect 807 2166 835 2170
rect 839 2166 1035 2170
rect 1039 2166 1075 2170
rect 1079 2166 1315 2170
rect 1319 2166 1563 2170
rect 1567 2166 1787 2170
rect 1791 2166 1935 2170
rect 1939 2166 1959 2170
rect 103 2165 1959 2166
rect 1965 2165 1966 2171
rect 1958 2105 1959 2111
rect 1965 2110 3823 2111
rect 1965 2106 1975 2110
rect 1979 2106 1995 2110
rect 1999 2106 2163 2110
rect 2167 2106 2331 2110
rect 2335 2106 2507 2110
rect 2511 2106 2683 2110
rect 2687 2106 2851 2110
rect 2855 2106 3019 2110
rect 3023 2106 3107 2110
rect 3111 2106 3179 2110
rect 3183 2106 3243 2110
rect 3247 2106 3339 2110
rect 3343 2106 3379 2110
rect 3383 2106 3507 2110
rect 3511 2106 3515 2110
rect 3519 2106 3651 2110
rect 3655 2106 3799 2110
rect 3803 2106 3823 2110
rect 1965 2105 3823 2106
rect 3829 2110 5714 2111
rect 3829 2106 3839 2110
rect 3843 2106 4515 2110
rect 4519 2106 4635 2110
rect 4639 2106 4691 2110
rect 4695 2106 4771 2110
rect 4775 2106 4883 2110
rect 4887 2106 4907 2110
rect 4911 2106 5043 2110
rect 5047 2106 5091 2110
rect 5095 2106 5179 2110
rect 5183 2106 5307 2110
rect 5311 2106 5515 2110
rect 5519 2106 5663 2110
rect 5667 2106 5714 2110
rect 3829 2105 5714 2106
rect 84 2049 85 2055
rect 91 2054 1947 2055
rect 91 2050 111 2054
rect 115 2050 159 2054
rect 163 2050 271 2054
rect 275 2050 375 2054
rect 379 2050 407 2054
rect 411 2050 543 2054
rect 547 2050 623 2054
rect 627 2050 687 2054
rect 691 2050 831 2054
rect 835 2050 863 2054
rect 867 2050 975 2054
rect 979 2050 1103 2054
rect 1107 2050 1119 2054
rect 1123 2050 1263 2054
rect 1267 2050 1343 2054
rect 1347 2050 1407 2054
rect 1411 2050 1543 2054
rect 1547 2050 1591 2054
rect 1595 2050 1679 2054
rect 1683 2050 1815 2054
rect 1819 2050 1935 2054
rect 1939 2050 1947 2054
rect 91 2049 1947 2050
rect 1953 2049 1954 2055
rect 1946 1993 1947 1999
rect 1953 1998 3811 1999
rect 1953 1994 1975 1998
rect 1979 1994 3127 1998
rect 3131 1994 3135 1998
rect 3139 1994 3263 1998
rect 3267 1994 3271 1998
rect 3275 1994 3399 1998
rect 3403 1994 3407 1998
rect 3411 1994 3535 1998
rect 3539 1994 3543 1998
rect 3547 1994 3671 1998
rect 3675 1994 3679 1998
rect 3683 1994 3799 1998
rect 3803 1994 3811 1998
rect 1953 1993 3811 1994
rect 3817 1998 5702 1999
rect 3817 1994 3839 1998
rect 3843 1994 4663 1998
rect 4667 1994 4799 1998
rect 4803 1994 4863 1998
rect 4867 1994 4935 1998
rect 4939 1994 4999 1998
rect 5003 1994 5071 1998
rect 5075 1994 5135 1998
rect 5139 1994 5207 1998
rect 5211 1994 5271 1998
rect 5275 1994 5407 1998
rect 5411 1994 5543 1998
rect 5547 1994 5663 1998
rect 5667 1994 5702 1998
rect 3817 1993 5702 1994
rect 96 1933 97 1939
rect 103 1938 1959 1939
rect 103 1934 111 1938
rect 115 1934 187 1938
rect 191 1934 243 1938
rect 247 1934 379 1938
rect 383 1934 515 1938
rect 519 1934 587 1938
rect 591 1934 659 1938
rect 663 1934 803 1938
rect 807 1934 811 1938
rect 815 1934 947 1938
rect 951 1934 1051 1938
rect 1055 1934 1091 1938
rect 1095 1934 1235 1938
rect 1239 1934 1299 1938
rect 1303 1934 1379 1938
rect 1383 1934 1515 1938
rect 1519 1934 1555 1938
rect 1559 1934 1651 1938
rect 1655 1934 1787 1938
rect 1791 1934 1935 1938
rect 1939 1934 1959 1938
rect 103 1933 1959 1934
rect 1965 1933 1966 1939
rect 1958 1869 1959 1875
rect 1965 1874 3823 1875
rect 1965 1870 1975 1874
rect 1979 1870 1995 1874
rect 1999 1870 2227 1874
rect 2231 1870 2467 1874
rect 2471 1870 2691 1874
rect 2695 1870 2907 1874
rect 2911 1870 3099 1874
rect 3103 1870 3107 1874
rect 3111 1870 3235 1874
rect 3239 1870 3299 1874
rect 3303 1870 3371 1874
rect 3375 1870 3483 1874
rect 3487 1870 3507 1874
rect 3511 1870 3643 1874
rect 3647 1870 3651 1874
rect 3655 1870 3799 1874
rect 3803 1870 3823 1874
rect 1965 1869 3823 1870
rect 3829 1874 5714 1875
rect 3829 1870 3839 1874
rect 3843 1870 4675 1874
rect 4679 1870 4819 1874
rect 4823 1870 4835 1874
rect 4839 1870 4963 1874
rect 4967 1870 4971 1874
rect 4975 1870 5107 1874
rect 5111 1870 5243 1874
rect 5247 1870 5379 1874
rect 5383 1870 5515 1874
rect 5519 1870 5663 1874
rect 5667 1870 5714 1874
rect 3829 1869 5714 1870
rect 84 1813 85 1819
rect 91 1818 1947 1819
rect 91 1814 111 1818
rect 115 1814 159 1818
rect 163 1814 215 1818
rect 219 1814 375 1818
rect 379 1814 407 1818
rect 411 1814 591 1818
rect 595 1814 615 1818
rect 619 1814 799 1818
rect 803 1814 839 1818
rect 843 1814 999 1818
rect 1003 1814 1079 1818
rect 1083 1814 1191 1818
rect 1195 1814 1327 1818
rect 1331 1814 1383 1818
rect 1387 1814 1575 1818
rect 1579 1814 1583 1818
rect 1587 1814 1815 1818
rect 1819 1814 1935 1818
rect 1939 1814 1947 1818
rect 91 1813 1947 1814
rect 1953 1813 1954 1819
rect 1946 1749 1947 1755
rect 1953 1754 3811 1755
rect 1953 1750 1975 1754
rect 1979 1750 2023 1754
rect 2027 1750 2159 1754
rect 2163 1750 2255 1754
rect 2259 1750 2311 1754
rect 2315 1750 2471 1754
rect 2475 1750 2495 1754
rect 2499 1750 2639 1754
rect 2643 1750 2719 1754
rect 2723 1750 2807 1754
rect 2811 1750 2935 1754
rect 2939 1750 2975 1754
rect 2979 1750 3135 1754
rect 3139 1750 3151 1754
rect 3155 1750 3327 1754
rect 3331 1750 3511 1754
rect 3515 1750 3679 1754
rect 3683 1750 3799 1754
rect 3803 1750 3811 1754
rect 1953 1749 3811 1750
rect 3817 1749 3818 1755
rect 3810 1747 3818 1749
rect 3810 1741 3811 1747
rect 3817 1746 5695 1747
rect 3817 1742 3839 1746
rect 3843 1742 3887 1746
rect 3891 1742 4079 1746
rect 4083 1742 4303 1746
rect 4307 1742 4535 1746
rect 4539 1742 4703 1746
rect 4707 1742 4775 1746
rect 4779 1742 4847 1746
rect 4851 1742 4991 1746
rect 4995 1742 5023 1746
rect 5027 1742 5135 1746
rect 5139 1742 5271 1746
rect 5275 1742 5279 1746
rect 5283 1742 5407 1746
rect 5411 1742 5535 1746
rect 5539 1742 5543 1746
rect 5547 1742 5663 1746
rect 5667 1742 5695 1746
rect 3817 1741 5695 1742
rect 5701 1741 5702 1747
rect 96 1677 97 1683
rect 103 1682 1959 1683
rect 103 1678 111 1682
rect 115 1678 131 1682
rect 135 1678 347 1682
rect 351 1678 395 1682
rect 399 1678 563 1682
rect 567 1678 683 1682
rect 687 1678 771 1682
rect 775 1678 971 1682
rect 975 1678 979 1682
rect 983 1678 1163 1682
rect 1167 1678 1275 1682
rect 1279 1678 1355 1682
rect 1359 1678 1547 1682
rect 1551 1678 1935 1682
rect 1939 1678 1959 1682
rect 103 1677 1959 1678
rect 1965 1677 1966 1683
rect 1958 1629 1959 1635
rect 1965 1634 3823 1635
rect 1965 1630 1975 1634
rect 1979 1630 1995 1634
rect 1999 1630 2091 1634
rect 2095 1630 2131 1634
rect 2135 1630 2227 1634
rect 2231 1630 2283 1634
rect 2287 1630 2363 1634
rect 2367 1630 2443 1634
rect 2447 1630 2499 1634
rect 2503 1630 2611 1634
rect 2615 1630 2635 1634
rect 2639 1630 2771 1634
rect 2775 1630 2779 1634
rect 2783 1630 2907 1634
rect 2911 1630 2947 1634
rect 2951 1630 3043 1634
rect 3047 1630 3123 1634
rect 3127 1630 3179 1634
rect 3183 1630 3799 1634
rect 3803 1630 3823 1634
rect 1965 1629 3823 1630
rect 3829 1634 5714 1635
rect 3829 1630 3839 1634
rect 3843 1630 3859 1634
rect 3863 1630 3995 1634
rect 3999 1630 4051 1634
rect 4055 1630 4155 1634
rect 4159 1630 4275 1634
rect 4279 1630 4355 1634
rect 4359 1630 4507 1634
rect 4511 1630 4587 1634
rect 4591 1630 4747 1634
rect 4751 1630 4851 1634
rect 4855 1630 4995 1634
rect 4999 1630 5131 1634
rect 5135 1630 5251 1634
rect 5255 1630 5419 1634
rect 5423 1630 5507 1634
rect 5511 1630 5663 1634
rect 5667 1630 5714 1634
rect 3829 1629 5714 1630
rect 84 1553 85 1559
rect 91 1558 1947 1559
rect 91 1554 111 1558
rect 115 1554 159 1558
rect 163 1554 375 1558
rect 379 1554 423 1558
rect 427 1554 607 1558
rect 611 1554 711 1558
rect 715 1554 839 1558
rect 843 1554 1007 1558
rect 1011 1554 1071 1558
rect 1075 1554 1303 1558
rect 1307 1554 1935 1558
rect 1939 1554 1947 1558
rect 91 1553 1947 1554
rect 1953 1553 1954 1559
rect 3810 1517 3811 1523
rect 3817 1522 5695 1523
rect 3817 1518 3839 1522
rect 3843 1518 3887 1522
rect 3891 1518 4023 1522
rect 4027 1518 4159 1522
rect 4163 1518 4183 1522
rect 4187 1518 4303 1522
rect 4307 1518 4383 1522
rect 4387 1518 4495 1522
rect 4499 1518 4615 1522
rect 4619 1518 4719 1522
rect 4723 1518 4879 1522
rect 4883 1518 4967 1522
rect 4971 1518 5159 1522
rect 5163 1518 5223 1522
rect 5227 1518 5447 1522
rect 5451 1518 5487 1522
rect 5491 1518 5663 1522
rect 5667 1518 5695 1522
rect 3817 1517 5695 1518
rect 5701 1517 5702 1523
rect 1946 1497 1947 1503
rect 1953 1502 3811 1503
rect 1953 1498 1975 1502
rect 1979 1498 2023 1502
rect 2027 1498 2119 1502
rect 2123 1498 2159 1502
rect 2163 1498 2255 1502
rect 2259 1498 2295 1502
rect 2299 1498 2391 1502
rect 2395 1498 2431 1502
rect 2435 1498 2527 1502
rect 2531 1498 2567 1502
rect 2571 1498 2663 1502
rect 2667 1498 2703 1502
rect 2707 1498 2799 1502
rect 2803 1498 2839 1502
rect 2843 1498 2935 1502
rect 2939 1498 2975 1502
rect 2979 1498 3071 1502
rect 3075 1498 3207 1502
rect 3211 1498 3799 1502
rect 3803 1498 3811 1502
rect 1953 1497 3811 1498
rect 3817 1497 3818 1503
rect 96 1429 97 1435
rect 103 1434 1959 1435
rect 103 1430 111 1434
rect 115 1430 131 1434
rect 135 1430 347 1434
rect 351 1430 411 1434
rect 415 1430 579 1434
rect 583 1430 739 1434
rect 743 1430 811 1434
rect 815 1430 1043 1434
rect 1047 1430 1091 1434
rect 1095 1430 1275 1434
rect 1279 1430 1451 1434
rect 1455 1430 1787 1434
rect 1791 1430 1935 1434
rect 1939 1430 1959 1434
rect 103 1429 1959 1430
rect 1965 1429 1966 1435
rect 3822 1401 3823 1407
rect 3829 1406 5707 1407
rect 3829 1402 3839 1406
rect 3843 1402 3859 1406
rect 3863 1402 3995 1406
rect 3999 1402 4059 1406
rect 4063 1402 4131 1406
rect 4135 1402 4275 1406
rect 4279 1402 4307 1406
rect 4311 1402 4467 1406
rect 4471 1402 4579 1406
rect 4583 1402 4691 1406
rect 4695 1402 4875 1406
rect 4879 1402 4939 1406
rect 4943 1402 5187 1406
rect 5191 1402 5195 1406
rect 5199 1402 5459 1406
rect 5463 1402 5499 1406
rect 5503 1402 5663 1406
rect 5667 1402 5707 1406
rect 3829 1401 5707 1402
rect 5713 1401 5714 1407
rect 1958 1377 1959 1383
rect 1965 1382 3823 1383
rect 1965 1378 1975 1382
rect 1979 1378 1995 1382
rect 1999 1378 2131 1382
rect 2135 1378 2267 1382
rect 2271 1378 2275 1382
rect 2279 1378 2403 1382
rect 2407 1378 2539 1382
rect 2543 1378 2563 1382
rect 2567 1378 2675 1382
rect 2679 1378 2811 1382
rect 2815 1378 2843 1382
rect 2847 1378 2947 1382
rect 2951 1378 3123 1382
rect 3127 1378 3395 1382
rect 3399 1378 3651 1382
rect 3655 1378 3799 1382
rect 3803 1378 3823 1382
rect 1965 1377 3823 1378
rect 3829 1377 3830 1383
rect 84 1317 85 1323
rect 91 1322 1947 1323
rect 91 1318 111 1322
rect 115 1318 159 1322
rect 163 1318 359 1322
rect 363 1318 439 1322
rect 443 1318 575 1322
rect 579 1318 767 1322
rect 771 1318 775 1322
rect 779 1318 967 1322
rect 971 1318 1119 1322
rect 1123 1318 1151 1322
rect 1155 1318 1327 1322
rect 1331 1318 1479 1322
rect 1483 1318 1495 1322
rect 1499 1318 1663 1322
rect 1667 1318 1815 1322
rect 1819 1318 1935 1322
rect 1939 1318 1947 1322
rect 91 1317 1947 1318
rect 1953 1317 1954 1323
rect 3810 1281 3811 1287
rect 3817 1286 5695 1287
rect 3817 1282 3839 1286
rect 3843 1282 3887 1286
rect 3891 1282 4087 1286
rect 4091 1282 4335 1286
rect 4339 1282 4607 1286
rect 4611 1282 4615 1286
rect 4619 1282 4791 1286
rect 4795 1282 4903 1286
rect 4907 1282 4975 1286
rect 4979 1282 5167 1286
rect 5171 1282 5215 1286
rect 5219 1282 5367 1286
rect 5371 1282 5527 1286
rect 5531 1282 5543 1286
rect 5547 1282 5663 1286
rect 5667 1282 5695 1286
rect 3817 1281 5695 1282
rect 5701 1281 5702 1287
rect 1946 1241 1947 1247
rect 1953 1246 3811 1247
rect 1953 1242 1975 1246
rect 1979 1242 2023 1246
rect 2027 1242 2303 1246
rect 2307 1242 2591 1246
rect 2595 1242 2655 1246
rect 2659 1242 2831 1246
rect 2835 1242 2871 1246
rect 2875 1242 3007 1246
rect 3011 1242 3151 1246
rect 3155 1242 3183 1246
rect 3187 1242 3359 1246
rect 3363 1242 3423 1246
rect 3427 1242 3543 1246
rect 3547 1242 3679 1246
rect 3683 1242 3799 1246
rect 3803 1242 3811 1246
rect 1953 1241 3811 1242
rect 3817 1241 3818 1247
rect 96 1193 97 1199
rect 103 1198 1959 1199
rect 103 1194 111 1198
rect 115 1194 131 1198
rect 135 1194 291 1198
rect 295 1194 331 1198
rect 335 1194 475 1198
rect 479 1194 547 1198
rect 551 1194 659 1198
rect 663 1194 747 1198
rect 751 1194 835 1198
rect 839 1194 939 1198
rect 943 1194 1003 1198
rect 1007 1194 1123 1198
rect 1127 1194 1171 1198
rect 1175 1194 1299 1198
rect 1303 1194 1331 1198
rect 1335 1194 1467 1198
rect 1471 1194 1491 1198
rect 1495 1194 1635 1198
rect 1639 1194 1651 1198
rect 1655 1194 1787 1198
rect 1791 1194 1935 1198
rect 1939 1194 1959 1198
rect 103 1193 1959 1194
rect 1965 1193 1966 1199
rect 3822 1165 3823 1171
rect 3829 1170 5707 1171
rect 3829 1166 3839 1170
rect 3843 1166 4587 1170
rect 4591 1166 4763 1170
rect 4767 1166 4835 1170
rect 4839 1166 4947 1170
rect 4951 1166 4971 1170
rect 4975 1166 5107 1170
rect 5111 1166 5139 1170
rect 5143 1166 5243 1170
rect 5247 1166 5339 1170
rect 5343 1166 5379 1170
rect 5383 1166 5515 1170
rect 5519 1166 5663 1170
rect 5667 1166 5707 1170
rect 3829 1165 5707 1166
rect 5713 1165 5714 1171
rect 1958 1113 1959 1119
rect 1965 1118 3823 1119
rect 1965 1114 1975 1118
rect 1979 1114 1995 1118
rect 1999 1114 2171 1118
rect 2175 1114 2363 1118
rect 2367 1114 2547 1118
rect 2551 1114 2627 1118
rect 2631 1114 2723 1118
rect 2727 1114 2803 1118
rect 2807 1114 2891 1118
rect 2895 1114 2979 1118
rect 2983 1114 3059 1118
rect 3063 1114 3155 1118
rect 3159 1114 3219 1118
rect 3223 1114 3331 1118
rect 3335 1114 3387 1118
rect 3391 1114 3515 1118
rect 3519 1114 3799 1118
rect 3803 1114 3823 1118
rect 1965 1113 3823 1114
rect 3829 1113 3830 1119
rect 84 1069 85 1075
rect 91 1074 1947 1075
rect 91 1070 111 1074
rect 115 1070 159 1074
rect 163 1070 175 1074
rect 179 1070 319 1074
rect 323 1070 431 1074
rect 435 1070 503 1074
rect 507 1070 687 1074
rect 691 1070 863 1074
rect 867 1070 951 1074
rect 955 1070 1031 1074
rect 1035 1070 1199 1074
rect 1203 1070 1215 1074
rect 1219 1070 1359 1074
rect 1363 1070 1519 1074
rect 1523 1070 1679 1074
rect 1683 1070 1815 1074
rect 1819 1070 1935 1074
rect 1939 1070 1947 1074
rect 91 1069 1947 1070
rect 1953 1069 1954 1075
rect 3810 1049 3811 1055
rect 3817 1054 5695 1055
rect 3817 1050 3839 1054
rect 3843 1050 4807 1054
rect 4811 1050 4863 1054
rect 4867 1050 4943 1054
rect 4947 1050 4999 1054
rect 5003 1050 5079 1054
rect 5083 1050 5135 1054
rect 5139 1050 5215 1054
rect 5219 1050 5271 1054
rect 5275 1050 5351 1054
rect 5355 1050 5407 1054
rect 5411 1050 5487 1054
rect 5491 1050 5543 1054
rect 5547 1050 5663 1054
rect 5667 1050 5695 1054
rect 3817 1049 5695 1050
rect 5701 1049 5702 1055
rect 1946 1001 1947 1007
rect 1953 1006 3811 1007
rect 1953 1002 1975 1006
rect 1979 1002 2023 1006
rect 2027 1002 2191 1006
rect 2195 1002 2199 1006
rect 2203 1002 2375 1006
rect 2379 1002 2391 1006
rect 2395 1002 2567 1006
rect 2571 1002 2575 1006
rect 2579 1002 2751 1006
rect 2755 1002 2759 1006
rect 2763 1002 2919 1006
rect 2923 1002 2943 1006
rect 2947 1002 3087 1006
rect 3091 1002 3127 1006
rect 3131 1002 3247 1006
rect 3251 1002 3311 1006
rect 3315 1002 3415 1006
rect 3419 1002 3495 1006
rect 3499 1002 3679 1006
rect 3683 1002 3799 1006
rect 3803 1002 3811 1006
rect 1953 1001 3811 1002
rect 3817 1001 3818 1007
rect 96 945 97 951
rect 103 950 1959 951
rect 103 946 111 950
rect 115 946 147 950
rect 151 946 235 950
rect 239 946 403 950
rect 407 946 459 950
rect 463 946 659 950
rect 663 946 683 950
rect 687 946 907 950
rect 911 946 923 950
rect 927 946 1131 950
rect 1135 946 1187 950
rect 1191 946 1363 950
rect 1367 946 1935 950
rect 1939 946 1959 950
rect 103 945 1959 946
rect 1965 945 1966 951
rect 3822 933 3823 939
rect 3829 938 5707 939
rect 3829 934 3839 938
rect 3843 934 3859 938
rect 3863 934 3995 938
rect 3999 934 4171 938
rect 4175 934 4387 938
rect 4391 934 4643 938
rect 4647 934 4779 938
rect 4783 934 4915 938
rect 4919 934 4931 938
rect 4935 934 5051 938
rect 5055 934 5187 938
rect 5191 934 5235 938
rect 5239 934 5323 938
rect 5327 934 5459 938
rect 5463 934 5515 938
rect 5519 934 5663 938
rect 5667 934 5707 938
rect 3829 933 5707 934
rect 5713 933 5714 939
rect 1958 885 1959 891
rect 1965 890 3823 891
rect 1965 886 1975 890
rect 1979 886 1995 890
rect 1999 886 2163 890
rect 2167 886 2179 890
rect 2183 886 2347 890
rect 2351 886 2403 890
rect 2407 886 2539 890
rect 2543 886 2675 890
rect 2679 886 2731 890
rect 2735 886 2915 890
rect 2919 886 2987 890
rect 2991 886 3099 890
rect 3103 886 3283 890
rect 3287 886 3323 890
rect 3327 886 3467 890
rect 3471 886 3651 890
rect 3655 886 3799 890
rect 3803 886 3823 890
rect 1965 885 3823 886
rect 3829 885 3830 891
rect 84 817 85 823
rect 91 822 1947 823
rect 91 818 111 822
rect 115 818 175 822
rect 179 818 263 822
rect 267 818 431 822
rect 435 818 487 822
rect 491 818 671 822
rect 675 818 711 822
rect 715 818 903 822
rect 907 818 935 822
rect 939 818 1127 822
rect 1131 818 1159 822
rect 1163 818 1351 822
rect 1355 818 1391 822
rect 1395 818 1575 822
rect 1579 818 1935 822
rect 1939 818 1947 822
rect 91 817 1947 818
rect 1953 817 1954 823
rect 3810 821 3811 827
rect 3817 826 5695 827
rect 3817 822 3839 826
rect 3843 822 3887 826
rect 3891 822 4023 826
rect 4027 822 4159 826
rect 4163 822 4199 826
rect 4203 822 4295 826
rect 4299 822 4415 826
rect 4419 822 4431 826
rect 4435 822 4567 826
rect 4571 822 4671 826
rect 4675 822 4719 826
rect 4723 822 4895 826
rect 4899 822 4959 826
rect 4963 822 5087 826
rect 5091 822 5263 826
rect 5267 822 5287 826
rect 5291 822 5487 826
rect 5491 822 5543 826
rect 5547 822 5663 826
rect 5667 822 5695 826
rect 3817 821 5695 822
rect 5701 821 5702 827
rect 96 705 97 711
rect 103 710 1959 711
rect 103 706 111 710
rect 115 706 131 710
rect 135 706 147 710
rect 151 706 315 710
rect 319 706 403 710
rect 407 706 523 710
rect 527 706 643 710
rect 647 706 723 710
rect 727 706 875 710
rect 879 706 907 710
rect 911 706 1083 710
rect 1087 706 1099 710
rect 1103 706 1259 710
rect 1263 706 1323 710
rect 1327 706 1427 710
rect 1431 706 1547 710
rect 1551 706 1595 710
rect 1599 706 1771 710
rect 1775 706 1935 710
rect 1939 706 1959 710
rect 103 705 1959 706
rect 1965 705 1966 711
rect 3822 705 3823 711
rect 3829 710 5707 711
rect 3829 706 3839 710
rect 3843 706 3859 710
rect 3863 706 3995 710
rect 3999 706 4131 710
rect 4135 706 4267 710
rect 4271 706 4403 710
rect 4407 706 4539 710
rect 4543 706 4691 710
rect 4695 706 4699 710
rect 4703 706 4867 710
rect 4871 706 4891 710
rect 4895 706 5059 710
rect 5063 706 5099 710
rect 5103 706 5259 710
rect 5263 706 5315 710
rect 5319 706 5459 710
rect 5463 706 5515 710
rect 5519 706 5663 710
rect 5667 706 5707 710
rect 3829 705 5707 706
rect 5713 705 5714 711
rect 84 593 85 599
rect 91 598 1947 599
rect 91 594 111 598
rect 115 594 159 598
rect 163 594 343 598
rect 347 594 375 598
rect 379 594 551 598
rect 555 594 599 598
rect 603 594 751 598
rect 755 594 807 598
rect 811 594 935 598
rect 939 594 999 598
rect 1003 594 1111 598
rect 1115 594 1175 598
rect 1179 594 1287 598
rect 1291 594 1343 598
rect 1347 594 1455 598
rect 1459 594 1511 598
rect 1515 594 1623 598
rect 1627 594 1671 598
rect 1675 594 1799 598
rect 1803 594 1815 598
rect 1819 594 1935 598
rect 1939 594 1947 598
rect 91 593 1947 594
rect 1953 593 1954 599
rect 3810 593 3811 599
rect 3817 598 5695 599
rect 3817 594 3839 598
rect 3843 594 3887 598
rect 3891 594 4023 598
rect 4027 594 4071 598
rect 4075 594 4159 598
rect 4163 594 4295 598
rect 4299 594 4311 598
rect 4315 594 4431 598
rect 4435 594 4567 598
rect 4571 594 4575 598
rect 4579 594 4727 598
rect 4731 594 4855 598
rect 4859 594 4919 598
rect 4923 594 5127 598
rect 5131 594 5151 598
rect 5155 594 5343 598
rect 5347 594 5447 598
rect 5451 594 5543 598
rect 5547 594 5663 598
rect 5667 594 5695 598
rect 3817 593 5695 594
rect 5701 593 5702 599
rect 1946 573 1947 579
rect 1953 578 3811 579
rect 1953 574 1975 578
rect 1979 574 2023 578
rect 2027 574 2207 578
rect 2211 574 2431 578
rect 2435 574 2703 578
rect 2707 574 3015 578
rect 3019 574 3135 578
rect 3139 574 3271 578
rect 3275 574 3351 578
rect 3355 574 3407 578
rect 3411 574 3543 578
rect 3547 574 3679 578
rect 3683 574 3799 578
rect 3803 574 3811 578
rect 1953 573 3811 574
rect 3817 573 3818 579
rect 96 481 97 487
rect 103 486 1959 487
rect 103 482 111 486
rect 115 482 131 486
rect 135 482 155 486
rect 159 482 347 486
rect 351 482 483 486
rect 487 482 571 486
rect 575 482 779 486
rect 783 482 811 486
rect 815 482 971 486
rect 975 482 1139 486
rect 1143 482 1147 486
rect 1151 482 1315 486
rect 1319 482 1475 486
rect 1479 482 1483 486
rect 1487 482 1643 486
rect 1647 482 1787 486
rect 1791 482 1935 486
rect 1939 482 1959 486
rect 103 481 1959 482
rect 1965 481 1966 487
rect 3822 469 3823 475
rect 3829 474 5707 475
rect 3829 470 3839 474
rect 3843 470 3859 474
rect 3863 470 4043 474
rect 4047 470 4283 474
rect 4287 470 4451 474
rect 4455 470 4547 474
rect 4551 470 4643 474
rect 4647 470 4827 474
rect 4831 470 4843 474
rect 4847 470 5051 474
rect 5055 470 5123 474
rect 5127 470 5267 474
rect 5271 470 5419 474
rect 5423 470 5483 474
rect 5487 470 5663 474
rect 5667 470 5707 474
rect 3829 469 5707 470
rect 5713 469 5714 475
rect 3822 467 3830 469
rect 1958 461 1959 467
rect 1965 466 3823 467
rect 1965 462 1975 466
rect 1979 462 1995 466
rect 1999 462 2203 466
rect 2207 462 2427 466
rect 2431 462 2651 466
rect 2655 462 2859 466
rect 2863 462 3067 466
rect 3071 462 3107 466
rect 3111 462 3243 466
rect 3247 462 3267 466
rect 3271 462 3379 466
rect 3383 462 3467 466
rect 3471 462 3515 466
rect 3519 462 3651 466
rect 3655 462 3799 466
rect 3803 462 3823 466
rect 1965 461 3823 462
rect 3829 461 3830 467
rect 84 357 85 363
rect 91 362 1947 363
rect 91 358 111 362
rect 115 358 183 362
rect 187 358 279 362
rect 283 358 487 362
rect 491 358 511 362
rect 515 358 703 362
rect 707 358 839 362
rect 843 358 919 362
rect 923 358 1135 362
rect 1139 358 1167 362
rect 1171 358 1503 362
rect 1507 358 1815 362
rect 1819 358 1935 362
rect 1939 358 1947 362
rect 91 357 1947 358
rect 1953 357 1954 363
rect 3810 353 3811 359
rect 3817 358 5695 359
rect 3817 354 3839 358
rect 3843 354 4479 358
rect 4483 354 4615 358
rect 4619 354 4671 358
rect 4675 354 4775 358
rect 4779 354 4871 358
rect 4875 354 4951 358
rect 4955 354 5079 358
rect 5083 354 5135 358
rect 5139 354 5295 358
rect 5299 354 5327 358
rect 5331 354 5511 358
rect 5515 354 5527 358
rect 5531 354 5663 358
rect 5667 354 5695 358
rect 3817 353 5695 354
rect 5701 353 5702 359
rect 1946 333 1947 339
rect 1953 338 3811 339
rect 1953 334 1975 338
rect 1979 334 2023 338
rect 2027 334 2159 338
rect 2163 334 2231 338
rect 2235 334 2295 338
rect 2299 334 2431 338
rect 2435 334 2455 338
rect 2459 334 2567 338
rect 2571 334 2679 338
rect 2683 334 2703 338
rect 2707 334 2839 338
rect 2843 334 2887 338
rect 2891 334 2975 338
rect 2979 334 3095 338
rect 3099 334 3111 338
rect 3115 334 3247 338
rect 3251 334 3295 338
rect 3299 334 3383 338
rect 3387 334 3495 338
rect 3499 334 3519 338
rect 3523 334 3655 338
rect 3659 334 3679 338
rect 3683 334 3799 338
rect 3803 334 3811 338
rect 1953 333 3811 334
rect 3817 333 3818 339
rect 96 205 97 211
rect 103 210 1959 211
rect 103 206 111 210
rect 115 206 131 210
rect 135 206 251 210
rect 255 206 267 210
rect 271 206 403 210
rect 407 206 459 210
rect 463 206 539 210
rect 543 206 675 210
rect 679 206 811 210
rect 815 206 891 210
rect 895 206 947 210
rect 951 206 1083 210
rect 1087 206 1107 210
rect 1111 206 1935 210
rect 1939 206 1959 210
rect 103 205 1959 206
rect 1965 205 1966 211
rect 3822 201 3823 207
rect 3829 206 5707 207
rect 3829 202 3839 206
rect 3843 202 4291 206
rect 4295 202 4427 206
rect 4431 202 4563 206
rect 4567 202 4587 206
rect 4591 202 4699 206
rect 4703 202 4747 206
rect 4751 202 4835 206
rect 4839 202 4923 206
rect 4927 202 4971 206
rect 4975 202 5107 206
rect 5111 202 5243 206
rect 5247 202 5299 206
rect 5303 202 5379 206
rect 5383 202 5499 206
rect 5503 202 5515 206
rect 5519 202 5663 206
rect 5667 202 5707 206
rect 3829 201 5707 202
rect 5713 201 5714 207
rect 1958 185 1959 191
rect 1965 190 3823 191
rect 1965 186 1975 190
rect 1979 186 1995 190
rect 1999 186 2131 190
rect 2135 186 2267 190
rect 2271 186 2403 190
rect 2407 186 2539 190
rect 2543 186 2675 190
rect 2679 186 2811 190
rect 2815 186 2947 190
rect 2951 186 3083 190
rect 3087 186 3219 190
rect 3223 186 3355 190
rect 3359 186 3491 190
rect 3495 186 3627 190
rect 3631 186 3799 190
rect 3803 186 3823 190
rect 1965 185 3823 186
rect 3829 185 3830 191
rect 3042 132 3048 133
rect 3646 132 3652 133
rect 3042 128 3043 132
rect 3047 128 3647 132
rect 3651 128 3652 132
rect 3042 127 3048 128
rect 3646 127 3652 128
rect 84 93 85 99
rect 91 98 1947 99
rect 91 94 111 98
rect 115 94 159 98
rect 163 94 295 98
rect 299 94 431 98
rect 435 94 567 98
rect 571 94 703 98
rect 707 94 839 98
rect 843 94 975 98
rect 979 94 1111 98
rect 1115 94 1935 98
rect 1939 94 1947 98
rect 91 93 1947 94
rect 1953 93 1954 99
rect 3810 89 3811 95
rect 3817 94 5695 95
rect 3817 90 3839 94
rect 3843 90 4319 94
rect 4323 90 4455 94
rect 4459 90 4591 94
rect 4595 90 4727 94
rect 4731 90 4863 94
rect 4867 90 4999 94
rect 5003 90 5135 94
rect 5139 90 5271 94
rect 5275 90 5407 94
rect 5411 90 5543 94
rect 5547 90 5663 94
rect 5667 90 5695 94
rect 3817 89 5695 90
rect 5701 89 5702 95
rect 1946 73 1947 79
rect 1953 78 3811 79
rect 1953 74 1975 78
rect 1979 74 2023 78
rect 2027 74 2159 78
rect 2163 74 2295 78
rect 2299 74 2431 78
rect 2435 74 2567 78
rect 2571 74 2703 78
rect 2707 74 2839 78
rect 2843 74 2975 78
rect 2979 74 3111 78
rect 3115 74 3247 78
rect 3251 74 3383 78
rect 3387 74 3519 78
rect 3523 74 3655 78
rect 3659 74 3799 78
rect 3803 74 3811 78
rect 1953 73 3811 74
rect 3817 73 3818 79
<< m5c >>
rect 85 5753 91 5759
rect 1947 5753 1953 5759
rect 1947 5653 1953 5659
rect 3811 5653 3817 5659
rect 97 5641 103 5647
rect 1959 5641 1965 5647
rect 1959 5541 1965 5547
rect 3823 5541 3829 5547
rect 85 5529 91 5535
rect 1947 5529 1953 5535
rect 1947 5427 1953 5433
rect 97 5417 103 5423
rect 1959 5417 1965 5423
rect 3811 5421 3817 5427
rect 3811 5405 3817 5411
rect 5695 5405 5701 5411
rect 85 5305 91 5311
rect 1947 5305 1953 5311
rect 1959 5309 1965 5315
rect 3823 5309 3829 5315
rect 3823 5277 3829 5283
rect 5707 5277 5713 5283
rect 1947 5197 1953 5203
rect 3811 5197 3817 5203
rect 3811 5137 3817 5143
rect 5695 5137 5701 5143
rect 97 5089 103 5095
rect 1959 5089 1965 5095
rect 3823 5013 3829 5019
rect 5707 5013 5713 5019
rect 85 4977 91 4983
rect 1947 4977 1953 4983
rect 1947 4941 1953 4947
rect 3811 4941 3817 4947
rect 3811 4881 3817 4887
rect 5695 4881 5701 4887
rect 97 4857 103 4863
rect 1959 4857 1965 4863
rect 1959 4805 1965 4811
rect 3823 4805 3829 4811
rect 3823 4765 3829 4771
rect 5707 4765 5713 4771
rect 85 4737 91 4743
rect 1947 4737 1953 4743
rect 1947 4689 1953 4695
rect 3811 4689 3817 4695
rect 3811 4653 3817 4659
rect 5695 4653 5701 4659
rect 97 4609 103 4615
rect 1959 4609 1965 4615
rect 1959 4573 1965 4579
rect 3823 4573 3829 4579
rect 3823 4541 3829 4547
rect 5707 4541 5713 4547
rect 85 4493 91 4499
rect 1947 4493 1953 4499
rect 1947 4453 1953 4459
rect 3811 4453 3817 4459
rect 3811 4421 3817 4427
rect 5695 4421 5701 4427
rect 97 4377 103 4383
rect 1959 4377 1965 4383
rect 1959 4333 1965 4339
rect 3823 4333 3829 4339
rect 3823 4309 3829 4315
rect 5707 4309 5713 4315
rect 85 4249 91 4255
rect 1947 4249 1953 4255
rect 1947 4213 1953 4219
rect 3811 4213 3817 4219
rect 3811 4161 3817 4167
rect 5695 4161 5701 4167
rect 97 4133 103 4139
rect 1959 4133 1965 4139
rect 1959 4081 1965 4087
rect 3823 4081 3829 4087
rect 3823 4049 3829 4055
rect 5707 4049 5713 4055
rect 85 3997 91 4003
rect 1947 3997 1953 4003
rect 1947 3965 1953 3971
rect 3811 3965 3817 3971
rect 3811 3913 3817 3919
rect 5695 3913 5701 3919
rect 97 3857 103 3863
rect 1959 3857 1965 3863
rect 1959 3841 1965 3847
rect 3823 3841 3829 3847
rect 3823 3785 3829 3791
rect 5707 3785 5713 3791
rect 85 3745 91 3751
rect 1947 3745 1953 3751
rect 1947 3725 1953 3731
rect 3811 3725 3817 3731
rect 3811 3645 3817 3651
rect 5695 3645 5701 3651
rect 97 3621 103 3627
rect 1959 3621 1965 3627
rect 1959 3601 1965 3607
rect 3823 3601 3829 3607
rect 3823 3509 3829 3515
rect 5707 3509 5713 3515
rect 85 3485 91 3491
rect 1947 3485 1953 3491
rect 3811 3393 3817 3399
rect 5695 3393 5701 3399
rect 97 3357 103 3363
rect 1959 3357 1965 3363
rect 1959 3329 1965 3335
rect 3823 3329 3829 3335
rect 3823 3281 3829 3287
rect 5707 3281 5713 3287
rect 85 3245 91 3251
rect 1947 3245 1953 3251
rect 1947 3217 1953 3223
rect 3811 3217 3817 3223
rect 3811 3153 3817 3159
rect 5695 3153 5701 3159
rect 97 3125 103 3131
rect 1959 3125 1965 3131
rect 1959 3093 1965 3099
rect 3823 3093 3829 3099
rect 3823 3041 3829 3047
rect 5707 3041 5713 3047
rect 85 2985 91 2991
rect 1947 2985 1953 2991
rect 1947 2969 1953 2975
rect 3811 2969 3817 2975
rect 3811 2925 3817 2931
rect 5695 2925 5701 2931
rect 97 2873 103 2879
rect 1959 2873 1965 2879
rect 1959 2849 1965 2855
rect 3823 2849 3829 2855
rect 3823 2805 3829 2811
rect 5707 2805 5713 2811
rect 85 2757 91 2763
rect 1947 2757 1953 2763
rect 1947 2733 1953 2739
rect 3811 2733 3817 2739
rect 3811 2693 3817 2699
rect 5695 2693 5701 2699
rect 97 2645 103 2651
rect 1959 2645 1965 2651
rect 1959 2609 1965 2615
rect 3823 2609 3829 2615
rect 3823 2581 3829 2587
rect 5707 2581 5713 2587
rect 85 2533 91 2539
rect 1947 2533 1953 2539
rect 1947 2473 1953 2479
rect 3811 2473 3817 2479
rect 3811 2465 3817 2471
rect 5695 2465 5701 2471
rect 97 2417 103 2423
rect 1959 2417 1965 2423
rect 1959 2353 1965 2359
rect 3823 2353 3829 2359
rect 3823 2341 3829 2347
rect 5707 2341 5713 2347
rect 85 2289 91 2295
rect 1947 2289 1953 2295
rect 1947 2233 1953 2239
rect 3811 2233 3817 2239
rect 3811 2217 3817 2223
rect 5695 2217 5701 2223
rect 97 2165 103 2171
rect 1959 2165 1965 2171
rect 1959 2105 1965 2111
rect 3823 2105 3829 2111
rect 85 2049 91 2055
rect 1947 2049 1953 2055
rect 1947 1993 1953 1999
rect 3811 1993 3817 1999
rect 97 1933 103 1939
rect 1959 1933 1965 1939
rect 1959 1869 1965 1875
rect 3823 1869 3829 1875
rect 85 1813 91 1819
rect 1947 1813 1953 1819
rect 1947 1749 1953 1755
rect 3811 1749 3817 1755
rect 3811 1741 3817 1747
rect 5695 1741 5701 1747
rect 97 1677 103 1683
rect 1959 1677 1965 1683
rect 1959 1629 1965 1635
rect 3823 1629 3829 1635
rect 85 1553 91 1559
rect 1947 1553 1953 1559
rect 3811 1517 3817 1523
rect 5695 1517 5701 1523
rect 1947 1497 1953 1503
rect 3811 1497 3817 1503
rect 97 1429 103 1435
rect 1959 1429 1965 1435
rect 3823 1401 3829 1407
rect 5707 1401 5713 1407
rect 1959 1377 1965 1383
rect 3823 1377 3829 1383
rect 85 1317 91 1323
rect 1947 1317 1953 1323
rect 3811 1281 3817 1287
rect 5695 1281 5701 1287
rect 1947 1241 1953 1247
rect 3811 1241 3817 1247
rect 97 1193 103 1199
rect 1959 1193 1965 1199
rect 3823 1165 3829 1171
rect 5707 1165 5713 1171
rect 1959 1113 1965 1119
rect 3823 1113 3829 1119
rect 85 1069 91 1075
rect 1947 1069 1953 1075
rect 3811 1049 3817 1055
rect 5695 1049 5701 1055
rect 1947 1001 1953 1007
rect 3811 1001 3817 1007
rect 97 945 103 951
rect 1959 945 1965 951
rect 3823 933 3829 939
rect 5707 933 5713 939
rect 1959 885 1965 891
rect 3823 885 3829 891
rect 85 817 91 823
rect 1947 817 1953 823
rect 3811 821 3817 827
rect 5695 821 5701 827
rect 97 705 103 711
rect 1959 705 1965 711
rect 3823 705 3829 711
rect 5707 705 5713 711
rect 85 593 91 599
rect 1947 593 1953 599
rect 3811 593 3817 599
rect 5695 593 5701 599
rect 1947 573 1953 579
rect 3811 573 3817 579
rect 97 481 103 487
rect 1959 481 1965 487
rect 3823 469 3829 475
rect 5707 469 5713 475
rect 1959 461 1965 467
rect 3823 461 3829 467
rect 85 357 91 363
rect 1947 357 1953 363
rect 3811 353 3817 359
rect 5695 353 5701 359
rect 1947 333 1953 339
rect 3811 333 3817 339
rect 97 205 103 211
rect 1959 205 1965 211
rect 3823 201 3829 207
rect 5707 201 5713 207
rect 1959 185 1965 191
rect 3823 185 3829 191
rect 85 93 91 99
rect 1947 93 1953 99
rect 3811 89 3817 95
rect 5695 89 5701 95
rect 1947 73 1953 79
rect 3811 73 3817 79
<< m5 >>
rect 84 5759 92 5760
rect 84 5753 85 5759
rect 91 5753 92 5759
rect 84 5535 92 5753
rect 84 5529 85 5535
rect 91 5529 92 5535
rect 84 5311 92 5529
rect 84 5305 85 5311
rect 91 5305 92 5311
rect 84 4983 92 5305
rect 84 4977 85 4983
rect 91 4977 92 4983
rect 84 4743 92 4977
rect 84 4737 85 4743
rect 91 4737 92 4743
rect 84 4499 92 4737
rect 84 4493 85 4499
rect 91 4493 92 4499
rect 84 4255 92 4493
rect 84 4249 85 4255
rect 91 4249 92 4255
rect 84 4003 92 4249
rect 84 3997 85 4003
rect 91 3997 92 4003
rect 84 3751 92 3997
rect 84 3745 85 3751
rect 91 3745 92 3751
rect 84 3491 92 3745
rect 84 3485 85 3491
rect 91 3485 92 3491
rect 84 3251 92 3485
rect 84 3245 85 3251
rect 91 3245 92 3251
rect 84 2991 92 3245
rect 84 2985 85 2991
rect 91 2985 92 2991
rect 84 2763 92 2985
rect 84 2757 85 2763
rect 91 2757 92 2763
rect 84 2539 92 2757
rect 84 2533 85 2539
rect 91 2533 92 2539
rect 84 2295 92 2533
rect 84 2289 85 2295
rect 91 2289 92 2295
rect 84 2055 92 2289
rect 84 2049 85 2055
rect 91 2049 92 2055
rect 84 1819 92 2049
rect 84 1813 85 1819
rect 91 1813 92 1819
rect 84 1559 92 1813
rect 84 1553 85 1559
rect 91 1553 92 1559
rect 84 1323 92 1553
rect 84 1317 85 1323
rect 91 1317 92 1323
rect 84 1075 92 1317
rect 84 1069 85 1075
rect 91 1069 92 1075
rect 84 823 92 1069
rect 84 817 85 823
rect 91 817 92 823
rect 84 599 92 817
rect 84 593 85 599
rect 91 593 92 599
rect 84 363 92 593
rect 84 357 85 363
rect 91 357 92 363
rect 84 99 92 357
rect 84 93 85 99
rect 91 93 92 99
rect 84 72 92 93
rect 96 5647 104 5760
rect 96 5641 97 5647
rect 103 5641 104 5647
rect 96 5423 104 5641
rect 96 5417 97 5423
rect 103 5417 104 5423
rect 96 5095 104 5417
rect 96 5089 97 5095
rect 103 5089 104 5095
rect 96 4863 104 5089
rect 96 4857 97 4863
rect 103 4857 104 4863
rect 96 4615 104 4857
rect 96 4609 97 4615
rect 103 4609 104 4615
rect 96 4383 104 4609
rect 96 4377 97 4383
rect 103 4377 104 4383
rect 96 4139 104 4377
rect 96 4133 97 4139
rect 103 4133 104 4139
rect 96 3863 104 4133
rect 96 3857 97 3863
rect 103 3857 104 3863
rect 96 3627 104 3857
rect 96 3621 97 3627
rect 103 3621 104 3627
rect 96 3363 104 3621
rect 96 3357 97 3363
rect 103 3357 104 3363
rect 96 3131 104 3357
rect 96 3125 97 3131
rect 103 3125 104 3131
rect 96 2879 104 3125
rect 96 2873 97 2879
rect 103 2873 104 2879
rect 96 2651 104 2873
rect 96 2645 97 2651
rect 103 2645 104 2651
rect 96 2423 104 2645
rect 96 2417 97 2423
rect 103 2417 104 2423
rect 96 2171 104 2417
rect 96 2165 97 2171
rect 103 2165 104 2171
rect 96 1939 104 2165
rect 96 1933 97 1939
rect 103 1933 104 1939
rect 96 1683 104 1933
rect 96 1677 97 1683
rect 103 1677 104 1683
rect 96 1435 104 1677
rect 96 1429 97 1435
rect 103 1429 104 1435
rect 96 1199 104 1429
rect 96 1193 97 1199
rect 103 1193 104 1199
rect 96 951 104 1193
rect 96 945 97 951
rect 103 945 104 951
rect 96 711 104 945
rect 96 705 97 711
rect 103 705 104 711
rect 96 487 104 705
rect 96 481 97 487
rect 103 481 104 487
rect 96 211 104 481
rect 96 205 97 211
rect 103 205 104 211
rect 96 72 104 205
rect 1946 5759 1954 5760
rect 1946 5753 1947 5759
rect 1953 5753 1954 5759
rect 1946 5659 1954 5753
rect 1946 5653 1947 5659
rect 1953 5653 1954 5659
rect 1946 5535 1954 5653
rect 1946 5529 1947 5535
rect 1953 5529 1954 5535
rect 1946 5433 1954 5529
rect 1946 5427 1947 5433
rect 1953 5427 1954 5433
rect 1946 5311 1954 5427
rect 1946 5305 1947 5311
rect 1953 5305 1954 5311
rect 1946 5203 1954 5305
rect 1946 5197 1947 5203
rect 1953 5197 1954 5203
rect 1946 4983 1954 5197
rect 1946 4977 1947 4983
rect 1953 4977 1954 4983
rect 1946 4947 1954 4977
rect 1946 4941 1947 4947
rect 1953 4941 1954 4947
rect 1946 4743 1954 4941
rect 1946 4737 1947 4743
rect 1953 4737 1954 4743
rect 1946 4695 1954 4737
rect 1946 4689 1947 4695
rect 1953 4689 1954 4695
rect 1946 4499 1954 4689
rect 1946 4493 1947 4499
rect 1953 4493 1954 4499
rect 1946 4459 1954 4493
rect 1946 4453 1947 4459
rect 1953 4453 1954 4459
rect 1946 4255 1954 4453
rect 1946 4249 1947 4255
rect 1953 4249 1954 4255
rect 1946 4219 1954 4249
rect 1946 4213 1947 4219
rect 1953 4213 1954 4219
rect 1946 4003 1954 4213
rect 1946 3997 1947 4003
rect 1953 3997 1954 4003
rect 1946 3971 1954 3997
rect 1946 3965 1947 3971
rect 1953 3965 1954 3971
rect 1946 3751 1954 3965
rect 1946 3745 1947 3751
rect 1953 3745 1954 3751
rect 1946 3731 1954 3745
rect 1946 3725 1947 3731
rect 1953 3725 1954 3731
rect 1946 3491 1954 3725
rect 1946 3485 1947 3491
rect 1953 3485 1954 3491
rect 1946 3251 1954 3485
rect 1946 3245 1947 3251
rect 1953 3245 1954 3251
rect 1946 3223 1954 3245
rect 1946 3217 1947 3223
rect 1953 3217 1954 3223
rect 1946 2991 1954 3217
rect 1946 2985 1947 2991
rect 1953 2985 1954 2991
rect 1946 2975 1954 2985
rect 1946 2969 1947 2975
rect 1953 2969 1954 2975
rect 1946 2763 1954 2969
rect 1946 2757 1947 2763
rect 1953 2757 1954 2763
rect 1946 2739 1954 2757
rect 1946 2733 1947 2739
rect 1953 2733 1954 2739
rect 1946 2539 1954 2733
rect 1946 2533 1947 2539
rect 1953 2533 1954 2539
rect 1946 2479 1954 2533
rect 1946 2473 1947 2479
rect 1953 2473 1954 2479
rect 1946 2295 1954 2473
rect 1946 2289 1947 2295
rect 1953 2289 1954 2295
rect 1946 2239 1954 2289
rect 1946 2233 1947 2239
rect 1953 2233 1954 2239
rect 1946 2055 1954 2233
rect 1946 2049 1947 2055
rect 1953 2049 1954 2055
rect 1946 1999 1954 2049
rect 1946 1993 1947 1999
rect 1953 1993 1954 1999
rect 1946 1819 1954 1993
rect 1946 1813 1947 1819
rect 1953 1813 1954 1819
rect 1946 1755 1954 1813
rect 1946 1749 1947 1755
rect 1953 1749 1954 1755
rect 1946 1559 1954 1749
rect 1946 1553 1947 1559
rect 1953 1553 1954 1559
rect 1946 1503 1954 1553
rect 1946 1497 1947 1503
rect 1953 1497 1954 1503
rect 1946 1323 1954 1497
rect 1946 1317 1947 1323
rect 1953 1317 1954 1323
rect 1946 1247 1954 1317
rect 1946 1241 1947 1247
rect 1953 1241 1954 1247
rect 1946 1075 1954 1241
rect 1946 1069 1947 1075
rect 1953 1069 1954 1075
rect 1946 1007 1954 1069
rect 1946 1001 1947 1007
rect 1953 1001 1954 1007
rect 1946 823 1954 1001
rect 1946 817 1947 823
rect 1953 817 1954 823
rect 1946 599 1954 817
rect 1946 593 1947 599
rect 1953 593 1954 599
rect 1946 579 1954 593
rect 1946 573 1947 579
rect 1953 573 1954 579
rect 1946 363 1954 573
rect 1946 357 1947 363
rect 1953 357 1954 363
rect 1946 339 1954 357
rect 1946 333 1947 339
rect 1953 333 1954 339
rect 1946 99 1954 333
rect 1946 93 1947 99
rect 1953 93 1954 99
rect 1946 79 1954 93
rect 1946 73 1947 79
rect 1953 73 1954 79
rect 1946 72 1954 73
rect 1958 5647 1966 5760
rect 1958 5641 1959 5647
rect 1965 5641 1966 5647
rect 1958 5547 1966 5641
rect 1958 5541 1959 5547
rect 1965 5541 1966 5547
rect 1958 5423 1966 5541
rect 1958 5417 1959 5423
rect 1965 5417 1966 5423
rect 1958 5315 1966 5417
rect 1958 5309 1959 5315
rect 1965 5309 1966 5315
rect 1958 5095 1966 5309
rect 1958 5089 1959 5095
rect 1965 5089 1966 5095
rect 1958 4863 1966 5089
rect 1958 4857 1959 4863
rect 1965 4857 1966 4863
rect 1958 4811 1966 4857
rect 1958 4805 1959 4811
rect 1965 4805 1966 4811
rect 1958 4615 1966 4805
rect 1958 4609 1959 4615
rect 1965 4609 1966 4615
rect 1958 4579 1966 4609
rect 1958 4573 1959 4579
rect 1965 4573 1966 4579
rect 1958 4383 1966 4573
rect 1958 4377 1959 4383
rect 1965 4377 1966 4383
rect 1958 4339 1966 4377
rect 1958 4333 1959 4339
rect 1965 4333 1966 4339
rect 1958 4139 1966 4333
rect 1958 4133 1959 4139
rect 1965 4133 1966 4139
rect 1958 4087 1966 4133
rect 1958 4081 1959 4087
rect 1965 4081 1966 4087
rect 1958 3863 1966 4081
rect 1958 3857 1959 3863
rect 1965 3857 1966 3863
rect 1958 3847 1966 3857
rect 1958 3841 1959 3847
rect 1965 3841 1966 3847
rect 1958 3627 1966 3841
rect 1958 3621 1959 3627
rect 1965 3621 1966 3627
rect 1958 3607 1966 3621
rect 1958 3601 1959 3607
rect 1965 3601 1966 3607
rect 1958 3363 1966 3601
rect 1958 3357 1959 3363
rect 1965 3357 1966 3363
rect 1958 3335 1966 3357
rect 1958 3329 1959 3335
rect 1965 3329 1966 3335
rect 1958 3131 1966 3329
rect 1958 3125 1959 3131
rect 1965 3125 1966 3131
rect 1958 3099 1966 3125
rect 1958 3093 1959 3099
rect 1965 3093 1966 3099
rect 1958 2879 1966 3093
rect 1958 2873 1959 2879
rect 1965 2873 1966 2879
rect 1958 2855 1966 2873
rect 1958 2849 1959 2855
rect 1965 2849 1966 2855
rect 1958 2651 1966 2849
rect 1958 2645 1959 2651
rect 1965 2645 1966 2651
rect 1958 2615 1966 2645
rect 1958 2609 1959 2615
rect 1965 2609 1966 2615
rect 1958 2423 1966 2609
rect 1958 2417 1959 2423
rect 1965 2417 1966 2423
rect 1958 2359 1966 2417
rect 1958 2353 1959 2359
rect 1965 2353 1966 2359
rect 1958 2171 1966 2353
rect 1958 2165 1959 2171
rect 1965 2165 1966 2171
rect 1958 2111 1966 2165
rect 1958 2105 1959 2111
rect 1965 2105 1966 2111
rect 1958 1939 1966 2105
rect 1958 1933 1959 1939
rect 1965 1933 1966 1939
rect 1958 1875 1966 1933
rect 1958 1869 1959 1875
rect 1965 1869 1966 1875
rect 1958 1683 1966 1869
rect 1958 1677 1959 1683
rect 1965 1677 1966 1683
rect 1958 1635 1966 1677
rect 1958 1629 1959 1635
rect 1965 1629 1966 1635
rect 1958 1435 1966 1629
rect 1958 1429 1959 1435
rect 1965 1429 1966 1435
rect 1958 1383 1966 1429
rect 1958 1377 1959 1383
rect 1965 1377 1966 1383
rect 1958 1199 1966 1377
rect 1958 1193 1959 1199
rect 1965 1193 1966 1199
rect 1958 1119 1966 1193
rect 1958 1113 1959 1119
rect 1965 1113 1966 1119
rect 1958 951 1966 1113
rect 1958 945 1959 951
rect 1965 945 1966 951
rect 1958 891 1966 945
rect 1958 885 1959 891
rect 1965 885 1966 891
rect 1958 711 1966 885
rect 1958 705 1959 711
rect 1965 705 1966 711
rect 1958 487 1966 705
rect 1958 481 1959 487
rect 1965 481 1966 487
rect 1958 467 1966 481
rect 1958 461 1959 467
rect 1965 461 1966 467
rect 1958 211 1966 461
rect 1958 205 1959 211
rect 1965 205 1966 211
rect 1958 191 1966 205
rect 1958 185 1959 191
rect 1965 185 1966 191
rect 1958 72 1966 185
rect 3810 5659 3818 5760
rect 3810 5653 3811 5659
rect 3817 5653 3818 5659
rect 3810 5427 3818 5653
rect 3810 5421 3811 5427
rect 3817 5421 3818 5427
rect 3810 5411 3818 5421
rect 3810 5405 3811 5411
rect 3817 5405 3818 5411
rect 3810 5203 3818 5405
rect 3810 5197 3811 5203
rect 3817 5197 3818 5203
rect 3810 5143 3818 5197
rect 3810 5137 3811 5143
rect 3817 5137 3818 5143
rect 3810 4947 3818 5137
rect 3810 4941 3811 4947
rect 3817 4941 3818 4947
rect 3810 4887 3818 4941
rect 3810 4881 3811 4887
rect 3817 4881 3818 4887
rect 3810 4695 3818 4881
rect 3810 4689 3811 4695
rect 3817 4689 3818 4695
rect 3810 4659 3818 4689
rect 3810 4653 3811 4659
rect 3817 4653 3818 4659
rect 3810 4459 3818 4653
rect 3810 4453 3811 4459
rect 3817 4453 3818 4459
rect 3810 4427 3818 4453
rect 3810 4421 3811 4427
rect 3817 4421 3818 4427
rect 3810 4219 3818 4421
rect 3810 4213 3811 4219
rect 3817 4213 3818 4219
rect 3810 4167 3818 4213
rect 3810 4161 3811 4167
rect 3817 4161 3818 4167
rect 3810 3971 3818 4161
rect 3810 3965 3811 3971
rect 3817 3965 3818 3971
rect 3810 3919 3818 3965
rect 3810 3913 3811 3919
rect 3817 3913 3818 3919
rect 3810 3731 3818 3913
rect 3810 3725 3811 3731
rect 3817 3725 3818 3731
rect 3810 3651 3818 3725
rect 3810 3645 3811 3651
rect 3817 3645 3818 3651
rect 3810 3399 3818 3645
rect 3810 3393 3811 3399
rect 3817 3393 3818 3399
rect 3810 3223 3818 3393
rect 3810 3217 3811 3223
rect 3817 3217 3818 3223
rect 3810 3159 3818 3217
rect 3810 3153 3811 3159
rect 3817 3153 3818 3159
rect 3810 2975 3818 3153
rect 3810 2969 3811 2975
rect 3817 2969 3818 2975
rect 3810 2931 3818 2969
rect 3810 2925 3811 2931
rect 3817 2925 3818 2931
rect 3810 2739 3818 2925
rect 3810 2733 3811 2739
rect 3817 2733 3818 2739
rect 3810 2699 3818 2733
rect 3810 2693 3811 2699
rect 3817 2693 3818 2699
rect 3810 2479 3818 2693
rect 3810 2473 3811 2479
rect 3817 2473 3818 2479
rect 3810 2471 3818 2473
rect 3810 2465 3811 2471
rect 3817 2465 3818 2471
rect 3810 2239 3818 2465
rect 3810 2233 3811 2239
rect 3817 2233 3818 2239
rect 3810 2223 3818 2233
rect 3810 2217 3811 2223
rect 3817 2217 3818 2223
rect 3810 1999 3818 2217
rect 3810 1993 3811 1999
rect 3817 1993 3818 1999
rect 3810 1755 3818 1993
rect 3810 1749 3811 1755
rect 3817 1749 3818 1755
rect 3810 1747 3818 1749
rect 3810 1741 3811 1747
rect 3817 1741 3818 1747
rect 3810 1523 3818 1741
rect 3810 1517 3811 1523
rect 3817 1517 3818 1523
rect 3810 1503 3818 1517
rect 3810 1497 3811 1503
rect 3817 1497 3818 1503
rect 3810 1287 3818 1497
rect 3810 1281 3811 1287
rect 3817 1281 3818 1287
rect 3810 1247 3818 1281
rect 3810 1241 3811 1247
rect 3817 1241 3818 1247
rect 3810 1055 3818 1241
rect 3810 1049 3811 1055
rect 3817 1049 3818 1055
rect 3810 1007 3818 1049
rect 3810 1001 3811 1007
rect 3817 1001 3818 1007
rect 3810 827 3818 1001
rect 3810 821 3811 827
rect 3817 821 3818 827
rect 3810 599 3818 821
rect 3810 593 3811 599
rect 3817 593 3818 599
rect 3810 579 3818 593
rect 3810 573 3811 579
rect 3817 573 3818 579
rect 3810 359 3818 573
rect 3810 353 3811 359
rect 3817 353 3818 359
rect 3810 339 3818 353
rect 3810 333 3811 339
rect 3817 333 3818 339
rect 3810 95 3818 333
rect 3810 89 3811 95
rect 3817 89 3818 95
rect 3810 79 3818 89
rect 3810 73 3811 79
rect 3817 73 3818 79
rect 3810 72 3818 73
rect 3822 5547 3830 5760
rect 3822 5541 3823 5547
rect 3829 5541 3830 5547
rect 3822 5315 3830 5541
rect 3822 5309 3823 5315
rect 3829 5309 3830 5315
rect 3822 5283 3830 5309
rect 3822 5277 3823 5283
rect 3829 5277 3830 5283
rect 3822 5019 3830 5277
rect 3822 5013 3823 5019
rect 3829 5013 3830 5019
rect 3822 4811 3830 5013
rect 3822 4805 3823 4811
rect 3829 4805 3830 4811
rect 3822 4771 3830 4805
rect 3822 4765 3823 4771
rect 3829 4765 3830 4771
rect 3822 4579 3830 4765
rect 3822 4573 3823 4579
rect 3829 4573 3830 4579
rect 3822 4547 3830 4573
rect 3822 4541 3823 4547
rect 3829 4541 3830 4547
rect 3822 4339 3830 4541
rect 3822 4333 3823 4339
rect 3829 4333 3830 4339
rect 3822 4315 3830 4333
rect 3822 4309 3823 4315
rect 3829 4309 3830 4315
rect 3822 4087 3830 4309
rect 3822 4081 3823 4087
rect 3829 4081 3830 4087
rect 3822 4055 3830 4081
rect 3822 4049 3823 4055
rect 3829 4049 3830 4055
rect 3822 3847 3830 4049
rect 3822 3841 3823 3847
rect 3829 3841 3830 3847
rect 3822 3791 3830 3841
rect 3822 3785 3823 3791
rect 3829 3785 3830 3791
rect 3822 3607 3830 3785
rect 3822 3601 3823 3607
rect 3829 3601 3830 3607
rect 3822 3515 3830 3601
rect 3822 3509 3823 3515
rect 3829 3509 3830 3515
rect 3822 3335 3830 3509
rect 3822 3329 3823 3335
rect 3829 3329 3830 3335
rect 3822 3287 3830 3329
rect 3822 3281 3823 3287
rect 3829 3281 3830 3287
rect 3822 3099 3830 3281
rect 3822 3093 3823 3099
rect 3829 3093 3830 3099
rect 3822 3047 3830 3093
rect 3822 3041 3823 3047
rect 3829 3041 3830 3047
rect 3822 2855 3830 3041
rect 3822 2849 3823 2855
rect 3829 2849 3830 2855
rect 3822 2811 3830 2849
rect 3822 2805 3823 2811
rect 3829 2805 3830 2811
rect 3822 2615 3830 2805
rect 3822 2609 3823 2615
rect 3829 2609 3830 2615
rect 3822 2587 3830 2609
rect 3822 2581 3823 2587
rect 3829 2581 3830 2587
rect 3822 2359 3830 2581
rect 3822 2353 3823 2359
rect 3829 2353 3830 2359
rect 3822 2347 3830 2353
rect 3822 2341 3823 2347
rect 3829 2341 3830 2347
rect 3822 2111 3830 2341
rect 3822 2105 3823 2111
rect 3829 2105 3830 2111
rect 3822 1875 3830 2105
rect 3822 1869 3823 1875
rect 3829 1869 3830 1875
rect 3822 1635 3830 1869
rect 3822 1629 3823 1635
rect 3829 1629 3830 1635
rect 3822 1407 3830 1629
rect 3822 1401 3823 1407
rect 3829 1401 3830 1407
rect 3822 1383 3830 1401
rect 3822 1377 3823 1383
rect 3829 1377 3830 1383
rect 3822 1171 3830 1377
rect 3822 1165 3823 1171
rect 3829 1165 3830 1171
rect 3822 1119 3830 1165
rect 3822 1113 3823 1119
rect 3829 1113 3830 1119
rect 3822 939 3830 1113
rect 3822 933 3823 939
rect 3829 933 3830 939
rect 3822 891 3830 933
rect 3822 885 3823 891
rect 3829 885 3830 891
rect 3822 711 3830 885
rect 3822 705 3823 711
rect 3829 705 3830 711
rect 3822 475 3830 705
rect 3822 469 3823 475
rect 3829 469 3830 475
rect 3822 467 3830 469
rect 3822 461 3823 467
rect 3829 461 3830 467
rect 3822 207 3830 461
rect 3822 201 3823 207
rect 3829 201 3830 207
rect 3822 191 3830 201
rect 3822 185 3823 191
rect 3829 185 3830 191
rect 3822 72 3830 185
rect 5694 5411 5702 5760
rect 5694 5405 5695 5411
rect 5701 5405 5702 5411
rect 5694 5143 5702 5405
rect 5694 5137 5695 5143
rect 5701 5137 5702 5143
rect 5694 4887 5702 5137
rect 5694 4881 5695 4887
rect 5701 4881 5702 4887
rect 5694 4659 5702 4881
rect 5694 4653 5695 4659
rect 5701 4653 5702 4659
rect 5694 4427 5702 4653
rect 5694 4421 5695 4427
rect 5701 4421 5702 4427
rect 5694 4167 5702 4421
rect 5694 4161 5695 4167
rect 5701 4161 5702 4167
rect 5694 3919 5702 4161
rect 5694 3913 5695 3919
rect 5701 3913 5702 3919
rect 5694 3651 5702 3913
rect 5694 3645 5695 3651
rect 5701 3645 5702 3651
rect 5694 3399 5702 3645
rect 5694 3393 5695 3399
rect 5701 3393 5702 3399
rect 5694 3159 5702 3393
rect 5694 3153 5695 3159
rect 5701 3153 5702 3159
rect 5694 2931 5702 3153
rect 5694 2925 5695 2931
rect 5701 2925 5702 2931
rect 5694 2699 5702 2925
rect 5694 2693 5695 2699
rect 5701 2693 5702 2699
rect 5694 2471 5702 2693
rect 5694 2465 5695 2471
rect 5701 2465 5702 2471
rect 5694 2223 5702 2465
rect 5694 2217 5695 2223
rect 5701 2217 5702 2223
rect 5694 1747 5702 2217
rect 5694 1741 5695 1747
rect 5701 1741 5702 1747
rect 5694 1523 5702 1741
rect 5694 1517 5695 1523
rect 5701 1517 5702 1523
rect 5694 1287 5702 1517
rect 5694 1281 5695 1287
rect 5701 1281 5702 1287
rect 5694 1055 5702 1281
rect 5694 1049 5695 1055
rect 5701 1049 5702 1055
rect 5694 827 5702 1049
rect 5694 821 5695 827
rect 5701 821 5702 827
rect 5694 599 5702 821
rect 5694 593 5695 599
rect 5701 593 5702 599
rect 5694 359 5702 593
rect 5694 353 5695 359
rect 5701 353 5702 359
rect 5694 95 5702 353
rect 5694 89 5695 95
rect 5701 89 5702 95
rect 5694 72 5702 89
rect 5706 5283 5714 5760
rect 5706 5277 5707 5283
rect 5713 5277 5714 5283
rect 5706 5019 5714 5277
rect 5706 5013 5707 5019
rect 5713 5013 5714 5019
rect 5706 4771 5714 5013
rect 5706 4765 5707 4771
rect 5713 4765 5714 4771
rect 5706 4547 5714 4765
rect 5706 4541 5707 4547
rect 5713 4541 5714 4547
rect 5706 4315 5714 4541
rect 5706 4309 5707 4315
rect 5713 4309 5714 4315
rect 5706 4055 5714 4309
rect 5706 4049 5707 4055
rect 5713 4049 5714 4055
rect 5706 3791 5714 4049
rect 5706 3785 5707 3791
rect 5713 3785 5714 3791
rect 5706 3515 5714 3785
rect 5706 3509 5707 3515
rect 5713 3509 5714 3515
rect 5706 3287 5714 3509
rect 5706 3281 5707 3287
rect 5713 3281 5714 3287
rect 5706 3047 5714 3281
rect 5706 3041 5707 3047
rect 5713 3041 5714 3047
rect 5706 2811 5714 3041
rect 5706 2805 5707 2811
rect 5713 2805 5714 2811
rect 5706 2587 5714 2805
rect 5706 2581 5707 2587
rect 5713 2581 5714 2587
rect 5706 2347 5714 2581
rect 5706 2341 5707 2347
rect 5713 2341 5714 2347
rect 5706 1407 5714 2341
rect 5706 1401 5707 1407
rect 5713 1401 5714 1407
rect 5706 1171 5714 1401
rect 5706 1165 5707 1171
rect 5713 1165 5714 1171
rect 5706 939 5714 1165
rect 5706 933 5707 939
rect 5713 933 5714 939
rect 5706 711 5714 933
rect 5706 705 5707 711
rect 5713 705 5714 711
rect 5706 475 5714 705
rect 5706 469 5707 475
rect 5713 469 5714 475
rect 5706 207 5714 469
rect 5706 201 5707 207
rect 5713 201 5714 207
rect 5706 72 5714 201
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__271
timestamp 1731220469
transform 1 0 5656 0 -1 5628
box 7 3 12 24
use welltap_svt  __well_tap__270
timestamp 1731220469
transform 1 0 3832 0 -1 5628
box 7 3 12 24
use welltap_svt  __well_tap__269
timestamp 1731220469
transform 1 0 5656 0 1 5452
box 7 3 12 24
use welltap_svt  __well_tap__268
timestamp 1731220469
transform 1 0 3832 0 1 5452
box 7 3 12 24
use welltap_svt  __well_tap__267
timestamp 1731220469
transform 1 0 5656 0 -1 5384
box 7 3 12 24
use welltap_svt  __well_tap__266
timestamp 1731220469
transform 1 0 3832 0 -1 5384
box 7 3 12 24
use welltap_svt  __well_tap__265
timestamp 1731220469
transform 1 0 5656 0 1 5192
box 7 3 12 24
use welltap_svt  __well_tap__264
timestamp 1731220469
transform 1 0 3832 0 1 5192
box 7 3 12 24
use welltap_svt  __well_tap__263
timestamp 1731220469
transform 1 0 5656 0 -1 5116
box 7 3 12 24
use welltap_svt  __well_tap__262
timestamp 1731220469
transform 1 0 3832 0 -1 5116
box 7 3 12 24
use welltap_svt  __well_tap__261
timestamp 1731220469
transform 1 0 5656 0 1 4928
box 7 3 12 24
use welltap_svt  __well_tap__260
timestamp 1731220469
transform 1 0 3832 0 1 4928
box 7 3 12 24
use welltap_svt  __well_tap__259
timestamp 1731220469
transform 1 0 5656 0 -1 4860
box 7 3 12 24
use welltap_svt  __well_tap__258
timestamp 1731220469
transform 1 0 3832 0 -1 4860
box 7 3 12 24
use welltap_svt  __well_tap__257
timestamp 1731220469
transform 1 0 5656 0 1 4680
box 7 3 12 24
use welltap_svt  __well_tap__256
timestamp 1731220469
transform 1 0 3832 0 1 4680
box 7 3 12 24
use welltap_svt  __well_tap__255
timestamp 1731220469
transform 1 0 5656 0 -1 4632
box 7 3 12 24
use welltap_svt  __well_tap__254
timestamp 1731220469
transform 1 0 3832 0 -1 4632
box 7 3 12 24
use welltap_svt  __well_tap__253
timestamp 1731220469
transform 1 0 5656 0 1 4456
box 7 3 12 24
use welltap_svt  __well_tap__252
timestamp 1731220469
transform 1 0 3832 0 1 4456
box 7 3 12 24
use welltap_svt  __well_tap__251
timestamp 1731220469
transform 1 0 5656 0 -1 4400
box 7 3 12 24
use welltap_svt  __well_tap__250
timestamp 1731220469
transform 1 0 3832 0 -1 4400
box 7 3 12 24
use welltap_svt  __well_tap__249
timestamp 1731220469
transform 1 0 5656 0 1 4224
box 7 3 12 24
use welltap_svt  __well_tap__248
timestamp 1731220469
transform 1 0 3832 0 1 4224
box 7 3 12 24
use welltap_svt  __well_tap__247
timestamp 1731220469
transform 1 0 5656 0 -1 4140
box 7 3 12 24
use welltap_svt  __well_tap__246
timestamp 1731220469
transform 1 0 3832 0 -1 4140
box 7 3 12 24
use welltap_svt  __well_tap__245
timestamp 1731220469
transform 1 0 5656 0 1 3964
box 7 3 12 24
use welltap_svt  __well_tap__244
timestamp 1731220469
transform 1 0 3832 0 1 3964
box 7 3 12 24
use welltap_svt  __well_tap__243
timestamp 1731220469
transform 1 0 5656 0 -1 3892
box 7 3 12 24
use welltap_svt  __well_tap__242
timestamp 1731220469
transform 1 0 3832 0 -1 3892
box 7 3 12 24
use welltap_svt  __well_tap__241
timestamp 1731220469
transform 1 0 5656 0 1 3700
box 7 3 12 24
use welltap_svt  __well_tap__240
timestamp 1731220469
transform 1 0 3832 0 1 3700
box 7 3 12 24
use welltap_svt  __well_tap__239
timestamp 1731220469
transform 1 0 5656 0 -1 3624
box 7 3 12 24
use welltap_svt  __well_tap__238
timestamp 1731220469
transform 1 0 3832 0 -1 3624
box 7 3 12 24
use welltap_svt  __well_tap__237
timestamp 1731220469
transform 1 0 5656 0 1 3424
box 7 3 12 24
use welltap_svt  __well_tap__236
timestamp 1731220469
transform 1 0 3832 0 1 3424
box 7 3 12 24
use welltap_svt  __well_tap__235
timestamp 1731220469
transform 1 0 5656 0 -1 3372
box 7 3 12 24
use welltap_svt  __well_tap__234
timestamp 1731220469
transform 1 0 3832 0 -1 3372
box 7 3 12 24
use welltap_svt  __well_tap__233
timestamp 1731220469
transform 1 0 5656 0 1 3196
box 7 3 12 24
use welltap_svt  __well_tap__232
timestamp 1731220469
transform 1 0 3832 0 1 3196
box 7 3 12 24
use welltap_svt  __well_tap__231
timestamp 1731220469
transform 1 0 5656 0 -1 3132
box 7 3 12 24
use welltap_svt  __well_tap__230
timestamp 1731220469
transform 1 0 3832 0 -1 3132
box 7 3 12 24
use welltap_svt  __well_tap__229
timestamp 1731220469
transform 1 0 5656 0 1 2956
box 7 3 12 24
use welltap_svt  __well_tap__228
timestamp 1731220469
transform 1 0 3832 0 1 2956
box 7 3 12 24
use welltap_svt  __well_tap__227
timestamp 1731220469
transform 1 0 5656 0 -1 2904
box 7 3 12 24
use welltap_svt  __well_tap__226
timestamp 1731220469
transform 1 0 3832 0 -1 2904
box 7 3 12 24
use welltap_svt  __well_tap__225
timestamp 1731220469
transform 1 0 5656 0 1 2720
box 7 3 12 24
use welltap_svt  __well_tap__224
timestamp 1731220469
transform 1 0 3832 0 1 2720
box 7 3 12 24
use welltap_svt  __well_tap__223
timestamp 1731220469
transform 1 0 5656 0 -1 2672
box 7 3 12 24
use welltap_svt  __well_tap__222
timestamp 1731220469
transform 1 0 3832 0 -1 2672
box 7 3 12 24
use welltap_svt  __well_tap__221
timestamp 1731220469
transform 1 0 5656 0 1 2496
box 7 3 12 24
use welltap_svt  __well_tap__220
timestamp 1731220469
transform 1 0 3832 0 1 2496
box 7 3 12 24
use welltap_svt  __well_tap__219
timestamp 1731220469
transform 1 0 5656 0 -1 2444
box 7 3 12 24
use welltap_svt  __well_tap__218
timestamp 1731220469
transform 1 0 3832 0 -1 2444
box 7 3 12 24
use welltap_svt  __well_tap__217
timestamp 1731220469
transform 1 0 5656 0 1 2256
box 7 3 12 24
use welltap_svt  __well_tap__216
timestamp 1731220469
transform 1 0 3832 0 1 2256
box 7 3 12 24
use welltap_svt  __well_tap__215
timestamp 1731220469
transform 1 0 5656 0 -1 2196
box 7 3 12 24
use welltap_svt  __well_tap__214
timestamp 1731220469
transform 1 0 3832 0 -1 2196
box 7 3 12 24
use welltap_svt  __well_tap__213
timestamp 1731220469
transform 1 0 5656 0 1 2020
box 7 3 12 24
use welltap_svt  __well_tap__212
timestamp 1731220469
transform 1 0 3832 0 1 2020
box 7 3 12 24
use welltap_svt  __well_tap__211
timestamp 1731220469
transform 1 0 5656 0 -1 1972
box 7 3 12 24
use welltap_svt  __well_tap__210
timestamp 1731220469
transform 1 0 3832 0 -1 1972
box 7 3 12 24
use welltap_svt  __well_tap__209
timestamp 1731220469
transform 1 0 5656 0 1 1784
box 7 3 12 24
use welltap_svt  __well_tap__208
timestamp 1731220469
transform 1 0 3832 0 1 1784
box 7 3 12 24
use welltap_svt  __well_tap__207
timestamp 1731220469
transform 1 0 5656 0 -1 1720
box 7 3 12 24
use welltap_svt  __well_tap__206
timestamp 1731220469
transform 1 0 3832 0 -1 1720
box 7 3 12 24
use welltap_svt  __well_tap__205
timestamp 1731220469
transform 1 0 5656 0 1 1544
box 7 3 12 24
use welltap_svt  __well_tap__204
timestamp 1731220469
transform 1 0 3832 0 1 1544
box 7 3 12 24
use welltap_svt  __well_tap__203
timestamp 1731220469
transform 1 0 5656 0 -1 1496
box 7 3 12 24
use welltap_svt  __well_tap__202
timestamp 1731220469
transform 1 0 3832 0 -1 1496
box 7 3 12 24
use welltap_svt  __well_tap__201
timestamp 1731220469
transform 1 0 5656 0 1 1316
box 7 3 12 24
use welltap_svt  __well_tap__200
timestamp 1731220469
transform 1 0 3832 0 1 1316
box 7 3 12 24
use welltap_svt  __well_tap__199
timestamp 1731220469
transform 1 0 5656 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__198
timestamp 1731220469
transform 1 0 3832 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__197
timestamp 1731220469
transform 1 0 5656 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__196
timestamp 1731220469
transform 1 0 3832 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__195
timestamp 1731220469
transform 1 0 5656 0 -1 1028
box 7 3 12 24
use welltap_svt  __well_tap__194
timestamp 1731220469
transform 1 0 3832 0 -1 1028
box 7 3 12 24
use welltap_svt  __well_tap__193
timestamp 1731220469
transform 1 0 5656 0 1 848
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220469
transform 1 0 3832 0 1 848
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220469
transform 1 0 5656 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220469
transform 1 0 3832 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220469
transform 1 0 5656 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220469
transform 1 0 3832 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220469
transform 1 0 5656 0 -1 572
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220469
transform 1 0 3832 0 -1 572
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220469
transform 1 0 5656 0 1 384
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220469
transform 1 0 3832 0 1 384
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220469
transform 1 0 5656 0 -1 332
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220469
transform 1 0 3832 0 -1 332
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220469
transform 1 0 5656 0 1 116
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220469
transform 1 0 3832 0 1 116
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220469
transform 1 0 3792 0 -1 5632
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220469
transform 1 0 1968 0 -1 5632
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220469
transform 1 0 3792 0 1 5456
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220469
transform 1 0 1968 0 1 5456
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220469
transform 1 0 3792 0 -1 5400
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220469
transform 1 0 1968 0 -1 5400
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220469
transform 1 0 3792 0 1 5224
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220469
transform 1 0 1968 0 1 5224
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220469
transform 1 0 3792 0 -1 5176
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220469
transform 1 0 1968 0 -1 5176
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220469
transform 1 0 3792 0 1 5000
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220469
transform 1 0 1968 0 1 5000
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220469
transform 1 0 3792 0 -1 4920
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220469
transform 1 0 1968 0 -1 4920
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220469
transform 1 0 3792 0 1 4720
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220469
transform 1 0 1968 0 1 4720
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220469
transform 1 0 3792 0 -1 4668
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220469
transform 1 0 1968 0 -1 4668
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220469
transform 1 0 3792 0 1 4488
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220469
transform 1 0 1968 0 1 4488
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220469
transform 1 0 3792 0 -1 4432
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220469
transform 1 0 1968 0 -1 4432
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220469
transform 1 0 3792 0 1 4248
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220469
transform 1 0 1968 0 1 4248
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220469
transform 1 0 3792 0 -1 4192
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220469
transform 1 0 1968 0 -1 4192
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220469
transform 1 0 3792 0 1 3996
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220469
transform 1 0 1968 0 1 3996
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220469
transform 1 0 3792 0 -1 3944
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220469
transform 1 0 1968 0 -1 3944
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220469
transform 1 0 3792 0 1 3756
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220469
transform 1 0 1968 0 1 3756
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220469
transform 1 0 3792 0 -1 3704
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220469
transform 1 0 1968 0 -1 3704
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220469
transform 1 0 3792 0 1 3516
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220469
transform 1 0 1968 0 1 3516
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220469
transform 1 0 3792 0 -1 3460
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220469
transform 1 0 1968 0 -1 3460
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220469
transform 1 0 3792 0 1 3244
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220469
transform 1 0 1968 0 1 3244
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220469
transform 1 0 3792 0 -1 3196
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220469
transform 1 0 1968 0 -1 3196
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220469
transform 1 0 3792 0 1 3008
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220469
transform 1 0 1968 0 1 3008
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220469
transform 1 0 3792 0 -1 2948
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220469
transform 1 0 1968 0 -1 2948
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220469
transform 1 0 3792 0 1 2764
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220469
transform 1 0 1968 0 1 2764
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220469
transform 1 0 3792 0 -1 2712
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220469
transform 1 0 1968 0 -1 2712
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220469
transform 1 0 3792 0 1 2524
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220469
transform 1 0 1968 0 1 2524
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220469
transform 1 0 3792 0 -1 2452
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220469
transform 1 0 1968 0 -1 2452
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220469
transform 1 0 3792 0 1 2268
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220469
transform 1 0 1968 0 1 2268
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220469
transform 1 0 3792 0 -1 2212
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220469
transform 1 0 1968 0 -1 2212
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220469
transform 1 0 3792 0 1 2020
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220469
transform 1 0 1968 0 1 2020
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220469
transform 1 0 3792 0 -1 1972
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220469
transform 1 0 1968 0 -1 1972
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220469
transform 1 0 3792 0 1 1784
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220469
transform 1 0 1968 0 1 1784
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220469
transform 1 0 3792 0 -1 1728
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220469
transform 1 0 1968 0 -1 1728
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220469
transform 1 0 3792 0 1 1544
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220469
transform 1 0 1968 0 1 1544
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220469
transform 1 0 3792 0 -1 1476
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220469
transform 1 0 1968 0 -1 1476
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220469
transform 1 0 3792 0 1 1292
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220469
transform 1 0 1968 0 1 1292
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220469
transform 1 0 3792 0 -1 1220
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220469
transform 1 0 1968 0 -1 1220
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220469
transform 1 0 3792 0 1 1028
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220469
transform 1 0 1968 0 1 1028
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220469
transform 1 0 3792 0 -1 980
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220469
transform 1 0 1968 0 -1 980
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220469
transform 1 0 3792 0 1 800
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220469
transform 1 0 1968 0 1 800
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220469
transform 1 0 3792 0 -1 552
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220469
transform 1 0 1968 0 -1 552
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220469
transform 1 0 3792 0 1 376
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220469
transform 1 0 1968 0 1 376
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220469
transform 1 0 3792 0 -1 312
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220469
transform 1 0 1968 0 -1 312
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220469
transform 1 0 3792 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220469
transform 1 0 1968 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220469
transform 1 0 1928 0 -1 5732
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220469
transform 1 0 104 0 -1 5732
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220469
transform 1 0 1928 0 1 5556
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220469
transform 1 0 104 0 1 5556
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220469
transform 1 0 1928 0 -1 5508
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220469
transform 1 0 104 0 -1 5508
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220469
transform 1 0 1928 0 1 5332
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220469
transform 1 0 104 0 1 5332
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220469
transform 1 0 1928 0 -1 5284
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220469
transform 1 0 104 0 -1 5284
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220469
transform 1 0 1928 0 1 5004
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220469
transform 1 0 104 0 1 5004
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220469
transform 1 0 1928 0 -1 4956
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220469
transform 1 0 104 0 -1 4956
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220469
transform 1 0 1928 0 1 4772
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220469
transform 1 0 104 0 1 4772
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220469
transform 1 0 1928 0 -1 4716
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220469
transform 1 0 104 0 -1 4716
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220469
transform 1 0 1928 0 1 4524
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220469
transform 1 0 104 0 1 4524
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220469
transform 1 0 1928 0 -1 4472
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220469
transform 1 0 104 0 -1 4472
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220469
transform 1 0 1928 0 1 4292
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220469
transform 1 0 104 0 1 4292
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220469
transform 1 0 1928 0 -1 4228
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220469
transform 1 0 104 0 -1 4228
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220469
transform 1 0 1928 0 1 4048
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220469
transform 1 0 104 0 1 4048
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220469
transform 1 0 1928 0 -1 3976
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220469
transform 1 0 104 0 -1 3976
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220469
transform 1 0 1928 0 1 3772
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220469
transform 1 0 104 0 1 3772
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220469
transform 1 0 1928 0 -1 3724
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220469
transform 1 0 104 0 -1 3724
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220469
transform 1 0 1928 0 1 3536
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220469
transform 1 0 104 0 1 3536
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220469
transform 1 0 1928 0 -1 3464
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220469
transform 1 0 104 0 -1 3464
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220469
transform 1 0 1928 0 1 3272
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220469
transform 1 0 104 0 1 3272
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220469
transform 1 0 1928 0 -1 3224
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220469
transform 1 0 104 0 -1 3224
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220469
transform 1 0 1928 0 1 3040
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220469
transform 1 0 104 0 1 3040
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220469
transform 1 0 1928 0 -1 2964
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220469
transform 1 0 104 0 -1 2964
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220469
transform 1 0 1928 0 1 2788
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220469
transform 1 0 104 0 1 2788
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220469
transform 1 0 1928 0 -1 2736
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220469
transform 1 0 104 0 -1 2736
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220469
transform 1 0 1928 0 1 2560
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220469
transform 1 0 104 0 1 2560
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220469
transform 1 0 1928 0 -1 2512
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220469
transform 1 0 104 0 -1 2512
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220469
transform 1 0 1928 0 1 2332
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220469
transform 1 0 104 0 1 2332
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220469
transform 1 0 1928 0 -1 2268
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220469
transform 1 0 104 0 -1 2268
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220469
transform 1 0 1928 0 1 2080
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220469
transform 1 0 104 0 1 2080
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220469
transform 1 0 1928 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220469
transform 1 0 104 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220469
transform 1 0 1928 0 1 1848
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220469
transform 1 0 104 0 1 1848
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220469
transform 1 0 1928 0 -1 1792
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220469
transform 1 0 104 0 -1 1792
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220469
transform 1 0 1928 0 1 1592
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220469
transform 1 0 104 0 1 1592
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220469
transform 1 0 1928 0 -1 1532
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220469
transform 1 0 104 0 -1 1532
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220469
transform 1 0 1928 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220469
transform 1 0 104 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220469
transform 1 0 1928 0 -1 1296
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220469
transform 1 0 104 0 -1 1296
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220469
transform 1 0 1928 0 1 1108
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220469
transform 1 0 104 0 1 1108
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220469
transform 1 0 1928 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220469
transform 1 0 104 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220469
transform 1 0 1928 0 1 860
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220469
transform 1 0 104 0 1 860
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220469
transform 1 0 1928 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220469
transform 1 0 104 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220469
transform 1 0 1928 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220469
transform 1 0 104 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220469
transform 1 0 1928 0 -1 572
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220469
transform 1 0 104 0 -1 572
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220469
transform 1 0 1928 0 1 396
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220469
transform 1 0 104 0 1 396
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220469
transform 1 0 1928 0 -1 336
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220469
transform 1 0 104 0 -1 336
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220469
transform 1 0 1928 0 1 120
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220469
transform 1 0 104 0 1 120
box 7 3 12 24
use _0_0std_0_0cells_0_0FAX1  tst_5999_6
timestamp 1731220469
transform 1 0 5376 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5998_6
timestamp 1731220469
transform 1 0 5512 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5997_6
timestamp 1731220469
transform 1 0 5496 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5996_6
timestamp 1731220469
transform 1 0 5480 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5995_6
timestamp 1731220469
transform 1 0 5416 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5994_6
timestamp 1731220469
transform 1 0 5264 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5993_6
timestamp 1731220469
transform 1 0 5240 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5992_6
timestamp 1731220469
transform 1 0 5104 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5991_6
timestamp 1731220469
transform 1 0 4968 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5990_6
timestamp 1731220469
transform 1 0 4832 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5989_6
timestamp 1731220469
transform 1 0 4696 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5988_6
timestamp 1731220469
transform 1 0 4560 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5987_6
timestamp 1731220469
transform 1 0 4424 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5986_6
timestamp 1731220469
transform 1 0 4288 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5985_6
timestamp 1731220469
transform 1 0 5296 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5984_6
timestamp 1731220469
transform 1 0 5104 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5983_6
timestamp 1731220469
transform 1 0 4920 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5982_6
timestamp 1731220469
transform 1 0 4744 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5981_6
timestamp 1731220469
transform 1 0 4584 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5980_6
timestamp 1731220469
transform 1 0 5048 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5979_6
timestamp 1731220469
transform 1 0 4840 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5978_6
timestamp 1731220469
transform 1 0 4640 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5977_6
timestamp 1731220469
transform 1 0 4448 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5976_6
timestamp 1731220469
transform 1 0 5120 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5975_6
timestamp 1731220469
transform 1 0 4824 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5974_6
timestamp 1731220469
transform 1 0 4544 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5973_6
timestamp 1731220469
transform 1 0 4280 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5972_6
timestamp 1731220469
transform 1 0 4040 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5971_6
timestamp 1731220469
transform 1 0 5312 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5970_6
timestamp 1731220469
transform 1 0 5096 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5969_6
timestamp 1731220469
transform 1 0 4888 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5968_6
timestamp 1731220469
transform 1 0 4696 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5967_6
timestamp 1731220469
transform 1 0 4536 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5966_6
timestamp 1731220469
transform 1 0 4536 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5965_6
timestamp 1731220469
transform 1 0 4400 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5964_6
timestamp 1731220469
transform 1 0 4264 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5963_6
timestamp 1731220469
transform 1 0 4128 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5962_6
timestamp 1731220469
transform 1 0 3992 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5961_6
timestamp 1731220469
transform 1 0 3992 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5960_6
timestamp 1731220469
transform 1 0 4168 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5959_6
timestamp 1731220469
transform 1 0 4688 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5958_6
timestamp 1731220469
transform 1 0 4864 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5957_6
timestamp 1731220469
transform 1 0 5256 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5956_6
timestamp 1731220469
transform 1 0 5056 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5955_6
timestamp 1731220469
transform 1 0 4928 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5954_6
timestamp 1731220469
transform 1 0 4640 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5953_6
timestamp 1731220469
transform 1 0 4384 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5952_6
timestamp 1731220469
transform 1 0 5232 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5951_6
timestamp 1731220469
transform 1 0 5048 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5950_6
timestamp 1731220469
transform 1 0 4912 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5949_6
timestamp 1731220469
transform 1 0 4776 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5948_6
timestamp 1731220469
transform 1 0 5184 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5947_6
timestamp 1731220469
transform 1 0 5320 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5946_6
timestamp 1731220469
transform 1 0 5376 0 1 1056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5945_6
timestamp 1731220469
transform 1 0 5240 0 1 1056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5944_6
timestamp 1731220469
transform 1 0 5104 0 1 1056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5943_6
timestamp 1731220469
transform 1 0 4968 0 1 1056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5942_6
timestamp 1731220469
transform 1 0 4832 0 1 1056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5941_6
timestamp 1731220469
transform 1 0 5136 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5940_6
timestamp 1731220469
transform 1 0 4944 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5939_6
timestamp 1731220469
transform 1 0 4760 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5938_6
timestamp 1731220469
transform 1 0 4584 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5937_6
timestamp 1731220469
transform 1 0 5184 0 1 1292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5936_6
timestamp 1731220469
transform 1 0 4872 0 1 1292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5935_6
timestamp 1731220469
transform 1 0 4576 0 1 1292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5934_6
timestamp 1731220469
transform 1 0 4304 0 1 1292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5933_6
timestamp 1731220469
transform 1 0 4056 0 1 1292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5932_6
timestamp 1731220469
transform 1 0 5192 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5931_6
timestamp 1731220469
transform 1 0 4936 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5930_6
timestamp 1731220469
transform 1 0 4688 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5929_6
timestamp 1731220469
transform 1 0 4464 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5928_6
timestamp 1731220469
transform 1 0 4352 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5927_6
timestamp 1731220469
transform 1 0 4272 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5926_6
timestamp 1731220469
transform 1 0 3992 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5925_6
timestamp 1731220469
transform 1 0 3856 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5924_6
timestamp 1731220469
transform 1 0 4584 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5923_6
timestamp 1731220469
transform 1 0 5128 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5922_6
timestamp 1731220469
transform 1 0 4848 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5921_6
timestamp 1731220469
transform 1 0 4744 0 -1 1744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5920_6
timestamp 1731220469
transform 1 0 4504 0 -1 1744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5919_6
timestamp 1731220469
transform 1 0 4272 0 -1 1744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5918_6
timestamp 1731220469
transform 1 0 4992 0 -1 1744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5917_6
timestamp 1731220469
transform 1 0 4960 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5916_6
timestamp 1731220469
transform 1 0 4816 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5915_6
timestamp 1731220469
transform 1 0 4672 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5914_6
timestamp 1731220469
transform 1 0 4832 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5913_6
timestamp 1731220469
transform 1 0 4968 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5912_6
timestamp 1731220469
transform 1 0 5104 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5911_6
timestamp 1731220469
transform 1 0 5176 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5910_6
timestamp 1731220469
transform 1 0 5240 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5909_6
timestamp 1731220469
transform 1 0 5376 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5908_6
timestamp 1731220469
transform 1 0 5240 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5907_6
timestamp 1731220469
transform 1 0 5104 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5906_6
timestamp 1731220469
transform 1 0 5248 0 -1 1744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5905_6
timestamp 1731220469
transform 1 0 5416 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5904_6
timestamp 1731220469
transform 1 0 5336 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5903_6
timestamp 1731220469
transform 1 0 5456 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5902_6
timestamp 1731220469
transform 1 0 5456 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5901_6
timestamp 1731220469
transform 1 0 5512 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5900_6
timestamp 1731220469
transform 1 0 5512 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5899_6
timestamp 1731220469
transform 1 0 5512 0 1 1056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5898_6
timestamp 1731220469
transform 1 0 5512 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5897_6
timestamp 1731220469
transform 1 0 5496 0 1 1292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5896_6
timestamp 1731220469
transform 1 0 5456 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5895_6
timestamp 1731220469
transform 1 0 5504 0 -1 1744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5894_6
timestamp 1731220469
transform 1 0 5376 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5893_6
timestamp 1731220469
transform 1 0 5512 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5892_6
timestamp 1731220469
transform 1 0 5512 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5891_6
timestamp 1731220469
transform 1 0 5512 0 -1 2220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5890_6
timestamp 1731220469
transform 1 0 5512 0 1 2232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5889_6
timestamp 1731220469
transform 1 0 5336 0 1 2232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5888_6
timestamp 1731220469
transform 1 0 5368 0 -1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5887_6
timestamp 1731220469
transform 1 0 5320 0 1 2472
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5886_6
timestamp 1731220469
transform 1 0 5368 0 -1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5885_6
timestamp 1731220469
transform 1 0 5080 0 -1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5884_6
timestamp 1731220469
transform 1 0 4792 0 -1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5883_6
timestamp 1731220469
transform 1 0 4824 0 1 2472
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5882_6
timestamp 1731220469
transform 1 0 5072 0 1 2472
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5881_6
timestamp 1731220469
transform 1 0 5088 0 -1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5880_6
timestamp 1731220469
transform 1 0 4960 0 1 2232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5879_6
timestamp 1731220469
transform 1 0 5144 0 1 2232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5878_6
timestamp 1731220469
transform 1 0 5304 0 -1 2220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5877_6
timestamp 1731220469
transform 1 0 5088 0 -1 2220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5876_6
timestamp 1731220469
transform 1 0 5040 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5875_6
timestamp 1731220469
transform 1 0 4904 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5874_6
timestamp 1731220469
transform 1 0 4768 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5873_6
timestamp 1731220469
transform 1 0 4632 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5872_6
timestamp 1731220469
transform 1 0 4512 0 -1 2220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5871_6
timestamp 1731220469
transform 1 0 4688 0 -1 2220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5870_6
timestamp 1731220469
transform 1 0 4880 0 -1 2220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5869_6
timestamp 1731220469
transform 1 0 4784 0 1 2232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5868_6
timestamp 1731220469
transform 1 0 4608 0 1 2232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5867_6
timestamp 1731220469
transform 1 0 4440 0 1 2232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5866_6
timestamp 1731220469
transform 1 0 4816 0 -1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5865_6
timestamp 1731220469
transform 1 0 4552 0 -1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5864_6
timestamp 1731220469
transform 1 0 4296 0 -1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5863_6
timestamp 1731220469
transform 1 0 4328 0 1 2472
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5862_6
timestamp 1731220469
transform 1 0 4576 0 1 2472
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5861_6
timestamp 1731220469
transform 1 0 4512 0 -1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5860_6
timestamp 1731220469
transform 1 0 4224 0 -1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5859_6
timestamp 1731220469
transform 1 0 4808 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5858_6
timestamp 1731220469
transform 1 0 4672 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5857_6
timestamp 1731220469
transform 1 0 4536 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5856_6
timestamp 1731220469
transform 1 0 4400 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5855_6
timestamp 1731220469
transform 1 0 4264 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5854_6
timestamp 1731220469
transform 1 0 4128 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5853_6
timestamp 1731220469
transform 1 0 4000 0 -1 2928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5852_6
timestamp 1731220469
transform 1 0 4136 0 -1 2928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5851_6
timestamp 1731220469
transform 1 0 4544 0 -1 2928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5850_6
timestamp 1731220469
transform 1 0 4408 0 -1 2928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5849_6
timestamp 1731220469
transform 1 0 4272 0 -1 2928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5848_6
timestamp 1731220469
transform 1 0 4240 0 1 2932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5847_6
timestamp 1731220469
transform 1 0 4072 0 1 2932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5846_6
timestamp 1731220469
transform 1 0 4752 0 1 2932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5845_6
timestamp 1731220469
transform 1 0 4576 0 1 2932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5844_6
timestamp 1731220469
transform 1 0 4408 0 1 2932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5843_6
timestamp 1731220469
transform 1 0 4328 0 -1 3156
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5842_6
timestamp 1731220469
transform 1 0 4104 0 -1 3156
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5841_6
timestamp 1731220469
transform 1 0 5000 0 -1 3156
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5840_6
timestamp 1731220469
transform 1 0 4776 0 -1 3156
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5839_6
timestamp 1731220469
transform 1 0 4552 0 -1 3156
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5838_6
timestamp 1731220469
transform 1 0 4344 0 1 3172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5837_6
timestamp 1731220469
transform 1 0 4096 0 1 3172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5836_6
timestamp 1731220469
transform 1 0 4576 0 1 3172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5835_6
timestamp 1731220469
transform 1 0 4784 0 1 3172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5834_6
timestamp 1731220469
transform 1 0 4984 0 1 3172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5833_6
timestamp 1731220469
transform 1 0 5296 0 -1 3396
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5832_6
timestamp 1731220469
transform 1 0 5080 0 -1 3396
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5831_6
timestamp 1731220469
transform 1 0 4864 0 -1 3396
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5830_6
timestamp 1731220469
transform 1 0 4640 0 -1 3396
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5829_6
timestamp 1731220469
transform 1 0 4392 0 -1 3396
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5828_6
timestamp 1731220469
transform 1 0 5168 0 1 3400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5827_6
timestamp 1731220469
transform 1 0 5000 0 1 3400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5826_6
timestamp 1731220469
transform 1 0 4840 0 1 3400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5825_6
timestamp 1731220469
transform 1 0 4680 0 1 3400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5824_6
timestamp 1731220469
transform 1 0 4528 0 1 3400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5823_6
timestamp 1731220469
transform 1 0 5040 0 -1 3648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5822_6
timestamp 1731220469
transform 1 0 4800 0 -1 3648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5821_6
timestamp 1731220469
transform 1 0 4576 0 -1 3648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5820_6
timestamp 1731220469
transform 1 0 4368 0 -1 3648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5819_6
timestamp 1731220469
transform 1 0 4184 0 -1 3648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5818_6
timestamp 1731220469
transform 1 0 4688 0 1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5817_6
timestamp 1731220469
transform 1 0 4432 0 1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5816_6
timestamp 1731220469
transform 1 0 4200 0 1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5815_6
timestamp 1731220469
transform 1 0 3992 0 1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5814_6
timestamp 1731220469
transform 1 0 4960 0 1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5813_6
timestamp 1731220469
transform 1 0 5032 0 -1 3916
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5812_6
timestamp 1731220469
transform 1 0 4792 0 -1 3916
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5811_6
timestamp 1731220469
transform 1 0 4568 0 -1 3916
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5810_6
timestamp 1731220469
transform 1 0 4352 0 -1 3916
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5809_6
timestamp 1731220469
transform 1 0 4336 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5808_6
timestamp 1731220469
transform 1 0 4496 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5807_6
timestamp 1731220469
transform 1 0 4648 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5806_6
timestamp 1731220469
transform 1 0 4800 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5805_6
timestamp 1731220469
transform 1 0 4944 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5804_6
timestamp 1731220469
transform 1 0 5088 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5803_6
timestamp 1731220469
transform 1 0 5232 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5802_6
timestamp 1731220469
transform 1 0 5376 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5801_6
timestamp 1731220469
transform 1 0 5280 0 -1 3916
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5800_6
timestamp 1731220469
transform 1 0 5248 0 1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5799_6
timestamp 1731220469
transform 1 0 5288 0 -1 3648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5798_6
timestamp 1731220469
transform 1 0 5344 0 1 3400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5797_6
timestamp 1731220469
transform 1 0 5168 0 1 3172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5796_6
timestamp 1731220469
transform 1 0 5352 0 1 3172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5795_6
timestamp 1731220469
transform 1 0 5512 0 1 3172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5794_6
timestamp 1731220469
transform 1 0 5512 0 -1 3396
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5793_6
timestamp 1731220469
transform 1 0 5512 0 1 3400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5792_6
timestamp 1731220469
transform 1 0 5512 0 -1 3648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5791_6
timestamp 1731220469
transform 1 0 5512 0 1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5790_6
timestamp 1731220469
transform 1 0 5512 0 -1 3916
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5789_6
timestamp 1731220469
transform 1 0 5512 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5788_6
timestamp 1731220469
transform 1 0 5512 0 -1 4164
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5787_6
timestamp 1731220469
transform 1 0 5496 0 1 4200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5786_6
timestamp 1731220469
transform 1 0 5472 0 -1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5785_6
timestamp 1731220469
transform 1 0 5440 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5784_6
timestamp 1731220469
transform 1 0 5408 0 -1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5783_6
timestamp 1731220469
transform 1 0 5368 0 1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5782_6
timestamp 1731220469
transform 1 0 5376 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5781_6
timestamp 1731220469
transform 1 0 5152 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5780_6
timestamp 1731220469
transform 1 0 5064 0 1 4904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5779_6
timestamp 1731220469
transform 1 0 5296 0 1 4904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5778_6
timestamp 1731220469
transform 1 0 5208 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5777_6
timestamp 1731220469
transform 1 0 4928 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5776_6
timestamp 1731220469
transform 1 0 4712 0 1 5168
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5775_6
timestamp 1731220469
transform 1 0 4944 0 1 5168
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5774_6
timestamp 1731220469
transform 1 0 5184 0 1 5168
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5773_6
timestamp 1731220469
transform 1 0 5096 0 -1 5408
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5772_6
timestamp 1731220469
transform 1 0 4880 0 -1 5408
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5771_6
timestamp 1731220469
transform 1 0 4664 0 -1 5408
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5770_6
timestamp 1731220469
transform 1 0 4704 0 1 5428
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5769_6
timestamp 1731220469
transform 1 0 4856 0 1 5428
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5768_6
timestamp 1731220469
transform 1 0 5016 0 1 5428
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5767_6
timestamp 1731220469
transform 1 0 4984 0 -1 5652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5766_6
timestamp 1731220469
transform 1 0 4848 0 -1 5652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5765_6
timestamp 1731220469
transform 1 0 4712 0 -1 5652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5764_6
timestamp 1731220469
transform 1 0 4576 0 -1 5652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5763_6
timestamp 1731220469
transform 1 0 4440 0 -1 5652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5762_6
timestamp 1731220469
transform 1 0 4304 0 -1 5652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5761_6
timestamp 1731220469
transform 1 0 4248 0 1 5428
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5760_6
timestamp 1731220469
transform 1 0 4400 0 1 5428
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5759_6
timestamp 1731220469
transform 1 0 4552 0 1 5428
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5758_6
timestamp 1731220469
transform 1 0 4456 0 -1 5408
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5757_6
timestamp 1731220469
transform 1 0 4248 0 -1 5408
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5756_6
timestamp 1731220469
transform 1 0 4248 0 1 5168
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5755_6
timestamp 1731220469
transform 1 0 4480 0 1 5168
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5754_6
timestamp 1731220469
transform 1 0 4376 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5753_6
timestamp 1731220469
transform 1 0 4104 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5752_6
timestamp 1731220469
transform 1 0 4648 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5751_6
timestamp 1731220469
transform 1 0 4624 0 1 4904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5750_6
timestamp 1731220469
transform 1 0 4408 0 1 4904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5749_6
timestamp 1731220469
transform 1 0 4840 0 1 4904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5748_6
timestamp 1731220469
transform 1 0 4704 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5747_6
timestamp 1731220469
transform 1 0 4480 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5746_6
timestamp 1731220469
transform 1 0 4928 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5745_6
timestamp 1731220469
transform 1 0 5064 0 1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5744_6
timestamp 1731220469
transform 1 0 4760 0 1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5743_6
timestamp 1731220469
transform 1 0 4840 0 -1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5742_6
timestamp 1731220469
transform 1 0 5120 0 -1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5741_6
timestamp 1731220469
transform 1 0 5176 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5740_6
timestamp 1731220469
transform 1 0 4912 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5739_6
timestamp 1731220469
transform 1 0 4848 0 -1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5738_6
timestamp 1731220469
transform 1 0 5048 0 -1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5737_6
timestamp 1731220469
transform 1 0 5256 0 -1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5736_6
timestamp 1731220469
transform 1 0 5232 0 1 4200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5735_6
timestamp 1731220469
transform 1 0 4968 0 1 4200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5734_6
timestamp 1731220469
transform 1 0 4712 0 1 4200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5733_6
timestamp 1731220469
transform 1 0 4472 0 1 4200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5732_6
timestamp 1731220469
transform 1 0 4248 0 1 4200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5731_6
timestamp 1731220469
transform 1 0 4328 0 -1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5730_6
timestamp 1731220469
transform 1 0 4488 0 -1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5729_6
timestamp 1731220469
transform 1 0 4656 0 -1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5728_6
timestamp 1731220469
transform 1 0 4656 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5727_6
timestamp 1731220469
transform 1 0 4408 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5726_6
timestamp 1731220469
transform 1 0 4176 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5725_6
timestamp 1731220469
transform 1 0 4032 0 -1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5724_6
timestamp 1731220469
transform 1 0 4296 0 -1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5723_6
timestamp 1731220469
transform 1 0 4568 0 -1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5722_6
timestamp 1731220469
transform 1 0 4464 0 1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5721_6
timestamp 1731220469
transform 1 0 4184 0 1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5720_6
timestamp 1731220469
transform 1 0 3912 0 1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5719_6
timestamp 1731220469
transform 1 0 3856 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5718_6
timestamp 1731220469
transform 1 0 4040 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5717_6
timestamp 1731220469
transform 1 0 4256 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5716_6
timestamp 1731220469
transform 1 0 4208 0 1 4904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5715_6
timestamp 1731220469
transform 1 0 4016 0 1 4904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5714_6
timestamp 1731220469
transform 1 0 3856 0 1 4904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5713_6
timestamp 1731220469
transform 1 0 3856 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5712_6
timestamp 1731220469
transform 1 0 3648 0 1 4976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5711_6
timestamp 1731220469
transform 1 0 3648 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5710_6
timestamp 1731220469
transform 1 0 3464 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5709_6
timestamp 1731220469
transform 1 0 3256 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5708_6
timestamp 1731220469
transform 1 0 3376 0 1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5707_6
timestamp 1731220469
transform 1 0 3576 0 1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5706_6
timestamp 1731220469
transform 1 0 3576 0 -1 5424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5705_6
timestamp 1731220469
transform 1 0 3392 0 -1 5424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5704_6
timestamp 1731220469
transform 1 0 3216 0 -1 5424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5703_6
timestamp 1731220469
transform 1 0 3288 0 1 5432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5702_6
timestamp 1731220469
transform 1 0 3464 0 1 5432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5701_6
timestamp 1731220469
transform 1 0 3640 0 1 5432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5700_6
timestamp 1731220469
transform 1 0 3648 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5699_6
timestamp 1731220469
transform 1 0 3512 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5698_6
timestamp 1731220469
transform 1 0 3352 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5697_6
timestamp 1731220469
transform 1 0 3192 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5696_6
timestamp 1731220469
transform 1 0 3032 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5695_6
timestamp 1731220469
transform 1 0 2864 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5694_6
timestamp 1731220469
transform 1 0 2696 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5693_6
timestamp 1731220469
transform 1 0 2752 0 1 5432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5692_6
timestamp 1731220469
transform 1 0 2936 0 1 5432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5691_6
timestamp 1731220469
transform 1 0 3112 0 1 5432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5690_6
timestamp 1731220469
transform 1 0 3040 0 -1 5424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5689_6
timestamp 1731220469
transform 1 0 2856 0 -1 5424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5688_6
timestamp 1731220469
transform 1 0 3000 0 1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5687_6
timestamp 1731220469
transform 1 0 3184 0 1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5686_6
timestamp 1731220469
transform 1 0 3056 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5685_6
timestamp 1731220469
transform 1 0 2856 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5684_6
timestamp 1731220469
transform 1 0 2528 0 1 4976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5683_6
timestamp 1731220469
transform 1 0 3096 0 1 4976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5682_6
timestamp 1731220469
transform 1 0 2840 0 -1 4944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5681_6
timestamp 1731220469
transform 1 0 2976 0 -1 4944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5680_6
timestamp 1731220469
transform 1 0 3128 0 1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5679_6
timestamp 1731220469
transform 1 0 2928 0 1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5678_6
timestamp 1731220469
transform 1 0 2728 0 1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5677_6
timestamp 1731220469
transform 1 0 2664 0 -1 4692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5676_6
timestamp 1731220469
transform 1 0 2888 0 -1 4692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5675_6
timestamp 1731220469
transform 1 0 3336 0 -1 4692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5674_6
timestamp 1731220469
transform 1 0 3112 0 -1 4692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5673_6
timestamp 1731220469
transform 1 0 3000 0 1 4464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5672_6
timestamp 1731220469
transform 1 0 2792 0 1 4464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5671_6
timestamp 1731220469
transform 1 0 3200 0 1 4464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5670_6
timestamp 1731220469
transform 1 0 3400 0 1 4464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5669_6
timestamp 1731220469
transform 1 0 3608 0 1 4464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5668_6
timestamp 1731220469
transform 1 0 3648 0 -1 4456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5667_6
timestamp 1731220469
transform 1 0 3464 0 -1 4456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5666_6
timestamp 1731220469
transform 1 0 3256 0 -1 4456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5665_6
timestamp 1731220469
transform 1 0 3048 0 -1 4456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5664_6
timestamp 1731220469
transform 1 0 3448 0 1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5663_6
timestamp 1731220469
transform 1 0 3648 0 1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5662_6
timestamp 1731220469
transform 1 0 3856 0 1 4200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5661_6
timestamp 1731220469
transform 1 0 4040 0 1 4200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5660_6
timestamp 1731220469
transform 1 0 3856 0 -1 4164
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5659_6
timestamp 1731220469
transform 1 0 4944 0 -1 4164
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5658_6
timestamp 1731220469
transform 1 0 4384 0 -1 4164
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5657_6
timestamp 1731220469
transform 1 0 4168 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5656_6
timestamp 1731220469
transform 1 0 4000 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5655_6
timestamp 1731220469
transform 1 0 3856 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5654_6
timestamp 1731220469
transform 1 0 3648 0 -1 3968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5653_6
timestamp 1731220469
transform 1 0 3480 0 -1 3968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5652_6
timestamp 1731220469
transform 1 0 3288 0 -1 3968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5651_6
timestamp 1731220469
transform 1 0 3104 0 -1 3968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5650_6
timestamp 1731220469
transform 1 0 2912 0 -1 3968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5649_6
timestamp 1731220469
transform 1 0 3400 0 1 3732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5648_6
timestamp 1731220469
transform 1 0 3192 0 1 3732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5647_6
timestamp 1731220469
transform 1 0 2992 0 1 3732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5646_6
timestamp 1731220469
transform 1 0 2792 0 1 3732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5645_6
timestamp 1731220469
transform 1 0 2584 0 1 3732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5644_6
timestamp 1731220469
transform 1 0 2448 0 -1 3728
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5643_6
timestamp 1731220469
transform 1 0 2648 0 -1 3728
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5642_6
timestamp 1731220469
transform 1 0 2848 0 -1 3728
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5641_6
timestamp 1731220469
transform 1 0 3248 0 -1 3728
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5640_6
timestamp 1731220469
transform 1 0 3048 0 -1 3728
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5639_6
timestamp 1731220469
transform 1 0 2976 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5638_6
timestamp 1731220469
transform 1 0 2752 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5637_6
timestamp 1731220469
transform 1 0 3192 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5636_6
timestamp 1731220469
transform 1 0 3408 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5635_6
timestamp 1731220469
transform 1 0 3624 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5634_6
timestamp 1731220469
transform 1 0 3448 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5633_6
timestamp 1731220469
transform 1 0 3232 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5632_6
timestamp 1731220469
transform 1 0 3016 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5631_6
timestamp 1731220469
transform 1 0 3648 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5630_6
timestamp 1731220469
transform 1 0 3856 0 -1 3396
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5629_6
timestamp 1731220469
transform 1 0 4120 0 -1 3396
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5628_6
timestamp 1731220469
transform 1 0 3856 0 1 3172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5627_6
timestamp 1731220469
transform 1 0 3872 0 -1 3156
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5626_6
timestamp 1731220469
transform 1 0 3904 0 1 2932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5625_6
timestamp 1731220469
transform 1 0 3864 0 -1 2928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5624_6
timestamp 1731220469
transform 1 0 3856 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5623_6
timestamp 1731220469
transform 1 0 3992 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5622_6
timestamp 1731220469
transform 1 0 3928 0 -1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5621_6
timestamp 1731220469
transform 1 0 3856 0 1 2472
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5620_6
timestamp 1731220469
transform 1 0 4080 0 1 2472
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5619_6
timestamp 1731220469
transform 1 0 4056 0 -1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5618_6
timestamp 1731220469
transform 1 0 3856 0 -1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5617_6
timestamp 1731220469
transform 1 0 3648 0 -1 2476
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5616_6
timestamp 1731220469
transform 1 0 3648 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5615_6
timestamp 1731220469
transform 1 0 3480 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5614_6
timestamp 1731220469
transform 1 0 3408 0 -1 2476
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5613_6
timestamp 1731220469
transform 1 0 3152 0 -1 2476
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5612_6
timestamp 1731220469
transform 1 0 2896 0 -1 2476
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5611_6
timestamp 1731220469
transform 1 0 2824 0 1 2500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5610_6
timestamp 1731220469
transform 1 0 2960 0 1 2500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5609_6
timestamp 1731220469
transform 1 0 3096 0 1 2500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5608_6
timestamp 1731220469
transform 1 0 2984 0 -1 2736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5607_6
timestamp 1731220469
transform 1 0 2728 0 -1 2736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5606_6
timestamp 1731220469
transform 1 0 2472 0 -1 2736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5605_6
timestamp 1731220469
transform 1 0 2752 0 1 2740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5604_6
timestamp 1731220469
transform 1 0 3000 0 1 2740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5603_6
timestamp 1731220469
transform 1 0 2904 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5602_6
timestamp 1731220469
transform 1 0 3104 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5601_6
timestamp 1731220469
transform 1 0 3304 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5600_6
timestamp 1731220469
transform 1 0 3232 0 1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5599_6
timestamp 1731220469
transform 1 0 3464 0 1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5598_6
timestamp 1731220469
transform 1 0 3400 0 -1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5597_6
timestamp 1731220469
transform 1 0 3208 0 -1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5596_6
timestamp 1731220469
transform 1 0 3592 0 -1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5595_6
timestamp 1731220469
transform 1 0 3552 0 1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5594_6
timestamp 1731220469
transform 1 0 3368 0 1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5593_6
timestamp 1731220469
transform 1 0 3184 0 1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5592_6
timestamp 1731220469
transform 1 0 3000 0 1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5591_6
timestamp 1731220469
transform 1 0 2808 0 1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5590_6
timestamp 1731220469
transform 1 0 2832 0 -1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5589_6
timestamp 1731220469
transform 1 0 3024 0 -1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5588_6
timestamp 1731220469
transform 1 0 3000 0 1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5587_6
timestamp 1731220469
transform 1 0 2776 0 1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5586_6
timestamp 1731220469
transform 1 0 2712 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5585_6
timestamp 1731220469
transform 1 0 2504 0 1 2740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5584_6
timestamp 1731220469
transform 1 0 2216 0 -1 2736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5583_6
timestamp 1731220469
transform 1 0 2552 0 1 2500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5582_6
timestamp 1731220469
transform 1 0 2688 0 1 2500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5581_6
timestamp 1731220469
transform 1 0 2648 0 -1 2476
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5580_6
timestamp 1731220469
transform 1 0 2416 0 -1 2476
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5579_6
timestamp 1731220469
transform 1 0 2192 0 -1 2476
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5578_6
timestamp 1731220469
transform 1 0 2536 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5577_6
timestamp 1731220469
transform 1 0 2728 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5576_6
timestamp 1731220469
transform 1 0 2680 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5575_6
timestamp 1731220469
transform 1 0 2504 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5574_6
timestamp 1731220469
transform 1 0 2328 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5573_6
timestamp 1731220469
transform 1 0 2160 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5572_6
timestamp 1731220469
transform 1 0 1992 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5571_6
timestamp 1731220469
transform 1 0 2344 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5570_6
timestamp 1731220469
transform 1 0 2152 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5569_6
timestamp 1731220469
transform 1 0 1992 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5568_6
timestamp 1731220469
transform 1 0 1992 0 -1 2476
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5567_6
timestamp 1731220469
transform 1 0 1784 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5566_6
timestamp 1731220469
transform 1 0 1784 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5565_6
timestamp 1731220469
transform 1 0 1600 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5564_6
timestamp 1731220469
transform 1 0 1400 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5563_6
timestamp 1731220469
transform 1 0 1512 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5562_6
timestamp 1731220469
transform 1 0 1672 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5561_6
timestamp 1731220469
transform 1 0 1768 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5560_6
timestamp 1731220469
transform 1 0 1992 0 -1 2736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5559_6
timestamp 1731220469
transform 1 0 2008 0 1 2740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5558_6
timestamp 1731220469
transform 1 0 2256 0 1 2740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5557_6
timestamp 1731220469
transform 1 0 2112 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5556_6
timestamp 1731220469
transform 1 0 2312 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5555_6
timestamp 1731220469
transform 1 0 2512 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5554_6
timestamp 1731220469
transform 1 0 2552 0 1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5553_6
timestamp 1731220469
transform 1 0 2328 0 1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5552_6
timestamp 1731220469
transform 1 0 2432 0 -1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5551_6
timestamp 1731220469
transform 1 0 2632 0 -1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5550_6
timestamp 1731220469
transform 1 0 2616 0 1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5549_6
timestamp 1731220469
transform 1 0 2408 0 1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5548_6
timestamp 1731220469
transform 1 0 2800 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5547_6
timestamp 1731220469
transform 1 0 2584 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5546_6
timestamp 1731220469
transform 1 0 2512 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5545_6
timestamp 1731220469
transform 1 0 2248 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5544_6
timestamp 1731220469
transform 1 0 2248 0 -1 3728
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5543_6
timestamp 1731220469
transform 1 0 2368 0 1 3732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5542_6
timestamp 1731220469
transform 1 0 2136 0 1 3732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5541_6
timestamp 1731220469
transform 1 0 2088 0 -1 3968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5540_6
timestamp 1731220469
transform 1 0 2296 0 -1 3968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5539_6
timestamp 1731220469
transform 1 0 2712 0 -1 3968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5538_6
timestamp 1731220469
transform 1 0 2504 0 -1 3968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5537_6
timestamp 1731220469
transform 1 0 2424 0 1 3972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5536_6
timestamp 1731220469
transform 1 0 2288 0 1 3972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5535_6
timestamp 1731220469
transform 1 0 2832 0 1 3972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5534_6
timestamp 1731220469
transform 1 0 2696 0 1 3972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5533_6
timestamp 1731220469
transform 1 0 2560 0 1 3972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5532_6
timestamp 1731220469
transform 1 0 2536 0 -1 4216
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5531_6
timestamp 1731220469
transform 1 0 2672 0 -1 4216
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5530_6
timestamp 1731220469
transform 1 0 2808 0 -1 4216
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5529_6
timestamp 1731220469
transform 1 0 2944 0 -1 4216
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5528_6
timestamp 1731220469
transform 1 0 3224 0 1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5527_6
timestamp 1731220469
transform 1 0 3008 0 1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5526_6
timestamp 1731220469
transform 1 0 2808 0 1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5525_6
timestamp 1731220469
transform 1 0 2624 0 1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5524_6
timestamp 1731220469
transform 1 0 2456 0 1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5523_6
timestamp 1731220469
transform 1 0 2304 0 1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5522_6
timestamp 1731220469
transform 1 0 2840 0 -1 4456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5521_6
timestamp 1731220469
transform 1 0 2632 0 -1 4456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5520_6
timestamp 1731220469
transform 1 0 2416 0 -1 4456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5519_6
timestamp 1731220469
transform 1 0 2200 0 -1 4456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5518_6
timestamp 1731220469
transform 1 0 2096 0 1 4464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5517_6
timestamp 1731220469
transform 1 0 2344 0 1 4464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5516_6
timestamp 1731220469
transform 1 0 2576 0 1 4464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5515_6
timestamp 1731220469
transform 1 0 2440 0 -1 4692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5514_6
timestamp 1731220469
transform 1 0 2208 0 -1 4692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5513_6
timestamp 1731220469
transform 1 0 1992 0 -1 4692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5512_6
timestamp 1731220469
transform 1 0 2536 0 1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5511_6
timestamp 1731220469
transform 1 0 2344 0 1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5510_6
timestamp 1731220469
transform 1 0 2152 0 1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5509_6
timestamp 1731220469
transform 1 0 1992 0 1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5508_6
timestamp 1731220469
transform 1 0 1784 0 -1 4740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5507_6
timestamp 1731220469
transform 1 0 1544 0 -1 4740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5506_6
timestamp 1731220469
transform 1 0 1280 0 -1 4740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5505_6
timestamp 1731220469
transform 1 0 1488 0 1 4500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5504_6
timestamp 1731220469
transform 1 0 1784 0 1 4500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5503_6
timestamp 1731220469
transform 1 0 1648 0 -1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5502_6
timestamp 1731220469
transform 1 0 1648 0 1 4268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5501_6
timestamp 1731220469
transform 1 0 1464 0 1 4268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5500_6
timestamp 1731220469
transform 1 0 1464 0 -1 4252
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5499_6
timestamp 1731220469
transform 1 0 1736 0 -1 4252
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5498_6
timestamp 1731220469
transform 1 0 1600 0 -1 4252
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5497_6
timestamp 1731220469
transform 1 0 1544 0 1 4024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5496_6
timestamp 1731220469
transform 1 0 1408 0 1 4024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5495_6
timestamp 1731220469
transform 1 0 1272 0 1 4024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5494_6
timestamp 1731220469
transform 1 0 1288 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5493_6
timestamp 1731220469
transform 1 0 1120 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5492_6
timestamp 1731220469
transform 1 0 1160 0 1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5491_6
timestamp 1731220469
transform 1 0 936 0 1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5490_6
timestamp 1731220469
transform 1 0 1024 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5489_6
timestamp 1731220469
transform 1 0 1040 0 1 3512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5488_6
timestamp 1731220469
transform 1 0 1080 0 -1 3488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5487_6
timestamp 1731220469
transform 1 0 904 0 -1 3488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5486_6
timestamp 1731220469
transform 1 0 464 0 1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5485_6
timestamp 1731220469
transform 1 0 504 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5484_6
timestamp 1731220469
transform 1 0 424 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5483_6
timestamp 1731220469
transform 1 0 168 0 -1 2988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5482_6
timestamp 1731220469
transform 1 0 480 0 -1 2988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5481_6
timestamp 1731220469
transform 1 0 784 0 -1 2988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5480_6
timestamp 1731220469
transform 1 0 1008 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5479_6
timestamp 1731220469
transform 1 0 760 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5478_6
timestamp 1731220469
transform 1 0 520 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5477_6
timestamp 1731220469
transform 1 0 304 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5476_6
timestamp 1731220469
transform 1 0 128 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5475_6
timestamp 1731220469
transform 1 0 248 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5474_6
timestamp 1731220469
transform 1 0 424 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5473_6
timestamp 1731220469
transform 1 0 616 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5472_6
timestamp 1731220469
transform 1 0 824 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5471_6
timestamp 1731220469
transform 1 0 1048 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5470_6
timestamp 1731220469
transform 1 0 888 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5469_6
timestamp 1731220469
transform 1 0 728 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5468_6
timestamp 1731220469
transform 1 0 568 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5467_6
timestamp 1731220469
transform 1 0 784 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5466_6
timestamp 1731220469
transform 1 0 568 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5465_6
timestamp 1731220469
transform 1 0 352 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5464_6
timestamp 1731220469
transform 1 0 224 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5463_6
timestamp 1731220469
transform 1 0 520 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5462_6
timestamp 1731220469
transform 1 0 568 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5461_6
timestamp 1731220469
transform 1 0 336 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5460_6
timestamp 1731220469
transform 1 0 128 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5459_6
timestamp 1731220469
transform 1 0 128 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5458_6
timestamp 1731220469
transform 1 0 344 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5457_6
timestamp 1731220469
transform 1 0 592 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5456_6
timestamp 1731220469
transform 1 0 512 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5455_6
timestamp 1731220469
transform 1 0 376 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5454_6
timestamp 1731220469
transform 1 0 240 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5453_6
timestamp 1731220469
transform 1 0 184 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5452_6
timestamp 1731220469
transform 1 0 376 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5451_6
timestamp 1731220469
transform 1 0 344 0 -1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5450_6
timestamp 1731220469
transform 1 0 128 0 -1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5449_6
timestamp 1731220469
transform 1 0 128 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5448_6
timestamp 1731220469
transform 1 0 128 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5447_6
timestamp 1731220469
transform 1 0 344 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5446_6
timestamp 1731220469
transform 1 0 128 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5445_6
timestamp 1731220469
transform 1 0 128 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5444_6
timestamp 1731220469
transform 1 0 128 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5443_6
timestamp 1731220469
transform 1 0 144 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5442_6
timestamp 1731220469
transform 1 0 400 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5441_6
timestamp 1731220469
transform 1 0 232 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5440_6
timestamp 1731220469
transform 1 0 144 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5439_6
timestamp 1731220469
transform 1 0 128 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5438_6
timestamp 1731220469
transform 1 0 312 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5437_6
timestamp 1731220469
transform 1 0 344 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5436_6
timestamp 1731220469
transform 1 0 128 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5435_6
timestamp 1731220469
transform 1 0 152 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5434_6
timestamp 1731220469
transform 1 0 480 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5433_6
timestamp 1731220469
transform 1 0 456 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5432_6
timestamp 1731220469
transform 1 0 248 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5431_6
timestamp 1731220469
transform 1 0 264 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5430_6
timestamp 1731220469
transform 1 0 128 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5429_6
timestamp 1731220469
transform 1 0 400 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5428_6
timestamp 1731220469
transform 1 0 536 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5427_6
timestamp 1731220469
transform 1 0 672 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5426_6
timestamp 1731220469
transform 1 0 1080 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5425_6
timestamp 1731220469
transform 1 0 944 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5424_6
timestamp 1731220469
transform 1 0 808 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5423_6
timestamp 1731220469
transform 1 0 672 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5422_6
timestamp 1731220469
transform 1 0 1104 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5421_6
timestamp 1731220469
transform 1 0 888 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5420_6
timestamp 1731220469
transform 1 0 808 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5419_6
timestamp 1731220469
transform 1 0 1472 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5418_6
timestamp 1731220469
transform 1 0 1136 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5417_6
timestamp 1731220469
transform 1 0 968 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5416_6
timestamp 1731220469
transform 1 0 776 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5415_6
timestamp 1731220469
transform 1 0 568 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5414_6
timestamp 1731220469
transform 1 0 520 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5413_6
timestamp 1731220469
transform 1 0 904 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5412_6
timestamp 1731220469
transform 1 0 720 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5411_6
timestamp 1731220469
transform 1 0 640 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5410_6
timestamp 1731220469
transform 1 0 400 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5409_6
timestamp 1731220469
transform 1 0 456 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5408_6
timestamp 1731220469
transform 1 0 680 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5407_6
timestamp 1731220469
transform 1 0 656 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5406_6
timestamp 1731220469
transform 1 0 656 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5405_6
timestamp 1731220469
transform 1 0 472 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5404_6
timestamp 1731220469
transform 1 0 288 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5403_6
timestamp 1731220469
transform 1 0 328 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5402_6
timestamp 1731220469
transform 1 0 544 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5401_6
timestamp 1731220469
transform 1 0 408 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5400_6
timestamp 1731220469
transform 1 0 736 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5399_6
timestamp 1731220469
transform 1 0 576 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5398_6
timestamp 1731220469
transform 1 0 808 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5397_6
timestamp 1731220469
transform 1 0 976 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5396_6
timestamp 1731220469
transform 1 0 1272 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5395_6
timestamp 1731220469
transform 1 0 1160 0 -1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5394_6
timestamp 1731220469
transform 1 0 968 0 -1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5393_6
timestamp 1731220469
transform 1 0 1352 0 -1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5392_6
timestamp 1731220469
transform 1 0 1544 0 -1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5391_6
timestamp 1731220469
transform 1 0 1552 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5390_6
timestamp 1731220469
transform 1 0 1296 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5389_6
timestamp 1731220469
transform 1 0 1232 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5388_6
timestamp 1731220469
transform 1 0 1088 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5387_6
timestamp 1731220469
transform 1 0 1512 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5386_6
timestamp 1731220469
transform 1 0 1376 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5385_6
timestamp 1731220469
transform 1 0 1312 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5384_6
timestamp 1731220469
transform 1 0 1560 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5383_6
timestamp 1731220469
transform 1 0 1784 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5382_6
timestamp 1731220469
transform 1 0 1648 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5381_6
timestamp 1731220469
transform 1 0 1784 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5380_6
timestamp 1731220469
transform 1 0 1784 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5379_6
timestamp 1731220469
transform 1 0 1992 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5378_6
timestamp 1731220469
transform 1 0 2224 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5377_6
timestamp 1731220469
transform 1 0 2464 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5376_6
timestamp 1731220469
transform 1 0 2280 0 -1 1752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5375_6
timestamp 1731220469
transform 1 0 2128 0 -1 1752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5374_6
timestamp 1731220469
transform 1 0 1992 0 -1 1752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5373_6
timestamp 1731220469
transform 1 0 2440 0 -1 1752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5372_6
timestamp 1731220469
transform 1 0 2608 0 -1 1752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5371_6
timestamp 1731220469
transform 1 0 2768 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5370_6
timestamp 1731220469
transform 1 0 2632 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5369_6
timestamp 1731220469
transform 1 0 2496 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5368_6
timestamp 1731220469
transform 1 0 2360 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5367_6
timestamp 1731220469
transform 1 0 2224 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5366_6
timestamp 1731220469
transform 1 0 2088 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5365_6
timestamp 1731220469
transform 1 0 2536 0 -1 1500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5364_6
timestamp 1731220469
transform 1 0 2400 0 -1 1500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5363_6
timestamp 1731220469
transform 1 0 2264 0 -1 1500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5362_6
timestamp 1731220469
transform 1 0 2128 0 -1 1500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5361_6
timestamp 1731220469
transform 1 0 1992 0 -1 1500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5360_6
timestamp 1731220469
transform 1 0 2272 0 1 1268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5359_6
timestamp 1731220469
transform 1 0 1992 0 1 1268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5358_6
timestamp 1731220469
transform 1 0 1784 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5357_6
timestamp 1731220469
transform 1 0 1784 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5356_6
timestamp 1731220469
transform 1 0 1632 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5355_6
timestamp 1731220469
transform 1 0 1464 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5354_6
timestamp 1731220469
transform 1 0 1296 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5353_6
timestamp 1731220469
transform 1 0 1120 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5352_6
timestamp 1731220469
transform 1 0 1168 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5351_6
timestamp 1731220469
transform 1 0 1328 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5350_6
timestamp 1731220469
transform 1 0 1488 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5349_6
timestamp 1731220469
transform 1 0 1648 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5348_6
timestamp 1731220469
transform 1 0 1784 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5347_6
timestamp 1731220469
transform 1 0 1992 0 1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5346_6
timestamp 1731220469
transform 1 0 1992 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5345_6
timestamp 1731220469
transform 1 0 2160 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5344_6
timestamp 1731220469
transform 1 0 2344 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5343_6
timestamp 1731220469
transform 1 0 2176 0 1 776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5342_6
timestamp 1731220469
transform 1 0 1992 0 1 776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5341_6
timestamp 1731220469
transform 1 0 2400 0 1 776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5340_6
timestamp 1731220469
transform 1 0 2672 0 1 776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5339_6
timestamp 1731220469
transform 1 0 3320 0 1 776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5338_6
timestamp 1731220469
transform 1 0 2984 0 1 776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5337_6
timestamp 1731220469
transform 1 0 2728 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5336_6
timestamp 1731220469
transform 1 0 2536 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5335_6
timestamp 1731220469
transform 1 0 2360 0 1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5334_6
timestamp 1731220469
transform 1 0 2168 0 1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5333_6
timestamp 1731220469
transform 1 0 2800 0 -1 1244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5332_6
timestamp 1731220469
transform 1 0 2624 0 -1 1244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5331_6
timestamp 1731220469
transform 1 0 2560 0 1 1268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5330_6
timestamp 1731220469
transform 1 0 2840 0 1 1268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5329_6
timestamp 1731220469
transform 1 0 2808 0 -1 1500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5328_6
timestamp 1731220469
transform 1 0 2672 0 -1 1500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5327_6
timestamp 1731220469
transform 1 0 2944 0 -1 1500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5326_6
timestamp 1731220469
transform 1 0 3176 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5325_6
timestamp 1731220469
transform 1 0 3040 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5324_6
timestamp 1731220469
transform 1 0 2904 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5323_6
timestamp 1731220469
transform 1 0 2776 0 -1 1752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5322_6
timestamp 1731220469
transform 1 0 3120 0 -1 1752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5321_6
timestamp 1731220469
transform 1 0 2944 0 -1 1752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5320_6
timestamp 1731220469
transform 1 0 2904 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5319_6
timestamp 1731220469
transform 1 0 2688 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5318_6
timestamp 1731220469
transform 1 0 3104 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5317_6
timestamp 1731220469
transform 1 0 3096 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5316_6
timestamp 1731220469
transform 1 0 3232 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5315_6
timestamp 1731220469
transform 1 0 3368 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5314_6
timestamp 1731220469
transform 1 0 3376 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5313_6
timestamp 1731220469
transform 1 0 3240 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5312_6
timestamp 1731220469
transform 1 0 3104 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5311_6
timestamp 1731220469
transform 1 0 3016 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5310_6
timestamp 1731220469
transform 1 0 2848 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5309_6
timestamp 1731220469
transform 1 0 3176 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5308_6
timestamp 1731220469
transform 1 0 3112 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5307_6
timestamp 1731220469
transform 1 0 2920 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5306_6
timestamp 1731220469
transform 1 0 3296 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5305_6
timestamp 1731220469
transform 1 0 3336 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5304_6
timestamp 1731220469
transform 1 0 3504 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5303_6
timestamp 1731220469
transform 1 0 3648 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5302_6
timestamp 1731220469
transform 1 0 3648 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5301_6
timestamp 1731220469
transform 1 0 3512 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5300_6
timestamp 1731220469
transform 1 0 3640 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5299_6
timestamp 1731220469
transform 1 0 3504 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5298_6
timestamp 1731220469
transform 1 0 3480 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5297_6
timestamp 1731220469
transform 1 0 3296 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5296_6
timestamp 1731220469
transform 1 0 3648 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5295_6
timestamp 1731220469
transform 1 0 3856 0 -1 1744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5294_6
timestamp 1731220469
transform 1 0 4048 0 -1 1744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5293_6
timestamp 1731220469
transform 1 0 4152 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5292_6
timestamp 1731220469
transform 1 0 4128 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5291_6
timestamp 1731220469
transform 1 0 3992 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5290_6
timestamp 1731220469
transform 1 0 3856 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5289_6
timestamp 1731220469
transform 1 0 3856 0 1 1292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5288_6
timestamp 1731220469
transform 1 0 3648 0 1 1268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5287_6
timestamp 1731220469
transform 1 0 3392 0 1 1268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5286_6
timestamp 1731220469
transform 1 0 3120 0 1 1268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5285_6
timestamp 1731220469
transform 1 0 3512 0 -1 1244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5284_6
timestamp 1731220469
transform 1 0 3328 0 -1 1244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5283_6
timestamp 1731220469
transform 1 0 3152 0 -1 1244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5282_6
timestamp 1731220469
transform 1 0 2976 0 -1 1244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5281_6
timestamp 1731220469
transform 1 0 3216 0 1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5280_6
timestamp 1731220469
transform 1 0 3056 0 1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5279_6
timestamp 1731220469
transform 1 0 2888 0 1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5278_6
timestamp 1731220469
transform 1 0 2720 0 1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5277_6
timestamp 1731220469
transform 1 0 2544 0 1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5276_6
timestamp 1731220469
transform 1 0 3384 0 1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5275_6
timestamp 1731220469
transform 1 0 3280 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5274_6
timestamp 1731220469
transform 1 0 3096 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5273_6
timestamp 1731220469
transform 1 0 2912 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5272_6
timestamp 1731220469
transform 1 0 3464 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5271_6
timestamp 1731220469
transform 1 0 3648 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5270_6
timestamp 1731220469
transform 1 0 3648 0 1 776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5269_6
timestamp 1731220469
transform 1 0 3856 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5268_6
timestamp 1731220469
transform 1 0 3856 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5267_6
timestamp 1731220469
transform 1 0 3856 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5266_6
timestamp 1731220469
transform 1 0 4400 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5265_6
timestamp 1731220469
transform 1 0 4264 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5264_6
timestamp 1731220469
transform 1 0 4128 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5263_6
timestamp 1731220469
transform 1 0 3992 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5262_6
timestamp 1731220469
transform 1 0 3856 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5261_6
timestamp 1731220469
transform 1 0 3648 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5260_6
timestamp 1731220469
transform 1 0 3512 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5259_6
timestamp 1731220469
transform 1 0 3376 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5258_6
timestamp 1731220469
transform 1 0 3240 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5257_6
timestamp 1731220469
transform 1 0 3104 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5256_6
timestamp 1731220469
transform 1 0 3648 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5255_6
timestamp 1731220469
transform 1 0 3464 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5254_6
timestamp 1731220469
transform 1 0 3264 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5253_6
timestamp 1731220469
transform 1 0 3064 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5252_6
timestamp 1731220469
transform 1 0 2856 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5251_6
timestamp 1731220469
transform 1 0 3624 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5250_6
timestamp 1731220469
transform 1 0 3488 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5249_6
timestamp 1731220469
transform 1 0 3352 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5248_6
timestamp 1731220469
transform 1 0 3216 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5247_6
timestamp 1731220469
transform 1 0 3080 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5246_6
timestamp 1731220469
transform 1 0 2944 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5245_6
timestamp 1731220469
transform 1 0 3624 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5244_6
timestamp 1731220469
transform 1 0 3488 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5243_6
timestamp 1731220469
transform 1 0 3352 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5242_6
timestamp 1731220469
transform 1 0 3216 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5241_6
timestamp 1731220469
transform 1 0 3080 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5240_6
timestamp 1731220469
transform 1 0 2944 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5239_6
timestamp 1731220469
transform 1 0 2808 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5238_6
timestamp 1731220469
transform 1 0 2672 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5237_6
timestamp 1731220469
transform 1 0 2536 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5236_6
timestamp 1731220469
transform 1 0 2400 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5235_6
timestamp 1731220469
transform 1 0 2264 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5234_6
timestamp 1731220469
transform 1 0 2128 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5233_6
timestamp 1731220469
transform 1 0 1992 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5232_6
timestamp 1731220469
transform 1 0 2808 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5231_6
timestamp 1731220469
transform 1 0 2672 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5230_6
timestamp 1731220469
transform 1 0 2536 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5229_6
timestamp 1731220469
transform 1 0 2400 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5228_6
timestamp 1731220469
transform 1 0 2264 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5227_6
timestamp 1731220469
transform 1 0 2128 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5226_6
timestamp 1731220469
transform 1 0 1992 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5225_6
timestamp 1731220469
transform 1 0 2648 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5224_6
timestamp 1731220469
transform 1 0 2424 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5223_6
timestamp 1731220469
transform 1 0 2200 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5222_6
timestamp 1731220469
transform 1 0 1992 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5221_6
timestamp 1731220469
transform 1 0 1784 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5220_6
timestamp 1731220469
transform 1 0 1784 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5219_6
timestamp 1731220469
transform 1 0 1640 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5218_6
timestamp 1731220469
transform 1 0 1480 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5217_6
timestamp 1731220469
transform 1 0 1312 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5216_6
timestamp 1731220469
transform 1 0 1144 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5215_6
timestamp 1731220469
transform 1 0 1768 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5214_6
timestamp 1731220469
transform 1 0 1592 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5213_6
timestamp 1731220469
transform 1 0 1424 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5212_6
timestamp 1731220469
transform 1 0 1256 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5211_6
timestamp 1731220469
transform 1 0 1080 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5210_6
timestamp 1731220469
transform 1 0 872 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5209_6
timestamp 1731220469
transform 1 0 1096 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5208_6
timestamp 1731220469
transform 1 0 1320 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5207_6
timestamp 1731220469
transform 1 0 1544 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5206_6
timestamp 1731220469
transform 1 0 1360 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5205_6
timestamp 1731220469
transform 1 0 1128 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5204_6
timestamp 1731220469
transform 1 0 904 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5203_6
timestamp 1731220469
transform 1 0 920 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5202_6
timestamp 1731220469
transform 1 0 1184 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5201_6
timestamp 1731220469
transform 1 0 1000 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5200_6
timestamp 1731220469
transform 1 0 832 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5199_6
timestamp 1731220469
transform 1 0 744 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5198_6
timestamp 1731220469
transform 1 0 936 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5197_6
timestamp 1731220469
transform 1 0 1088 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5196_6
timestamp 1731220469
transform 1 0 1448 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5195_6
timestamp 1731220469
transform 1 0 1272 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5194_6
timestamp 1731220469
transform 1 0 1040 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5193_6
timestamp 1731220469
transform 1 0 680 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5192_6
timestamp 1731220469
transform 1 0 392 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5191_6
timestamp 1731220469
transform 1 0 560 0 -1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5190_6
timestamp 1731220469
transform 1 0 768 0 -1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5189_6
timestamp 1731220469
transform 1 0 1048 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5188_6
timestamp 1731220469
transform 1 0 808 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5187_6
timestamp 1731220469
transform 1 0 584 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5186_6
timestamp 1731220469
transform 1 0 656 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5185_6
timestamp 1731220469
transform 1 0 800 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5184_6
timestamp 1731220469
transform 1 0 944 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5183_6
timestamp 1731220469
transform 1 0 832 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5182_6
timestamp 1731220469
transform 1 0 1072 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5181_6
timestamp 1731220469
transform 1 0 1032 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5180_6
timestamp 1731220469
transform 1 0 800 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5179_6
timestamp 1731220469
transform 1 0 832 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5178_6
timestamp 1731220469
transform 1 0 1152 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5177_6
timestamp 1731220469
transform 1 0 1480 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5176_6
timestamp 1731220469
transform 1 0 1200 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5175_6
timestamp 1731220469
transform 1 0 992 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5174_6
timestamp 1731220469
transform 1 0 1040 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5173_6
timestamp 1731220469
transform 1 0 1192 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5172_6
timestamp 1731220469
transform 1 0 1352 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5171_6
timestamp 1731220469
transform 1 0 1280 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5170_6
timestamp 1731220469
transform 1 0 1520 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5169_6
timestamp 1731220469
transform 1 0 1536 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5168_6
timestamp 1731220469
transform 1 0 1272 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5167_6
timestamp 1731220469
transform 1 0 1080 0 -1 2988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5166_6
timestamp 1731220469
transform 1 0 1384 0 -1 2988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5165_6
timestamp 1731220469
transform 1 0 1688 0 -1 2988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5164_6
timestamp 1731220469
transform 1 0 1784 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5163_6
timestamp 1731220469
transform 1 0 1648 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5162_6
timestamp 1731220469
transform 1 0 1512 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5161_6
timestamp 1731220469
transform 1 0 1440 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5160_6
timestamp 1731220469
transform 1 0 1624 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5159_6
timestamp 1731220469
transform 1 0 1784 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5158_6
timestamp 1731220469
transform 1 0 1992 0 1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5157_6
timestamp 1731220469
transform 1 0 2192 0 1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5156_6
timestamp 1731220469
transform 1 0 2368 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5155_6
timestamp 1731220469
transform 1 0 2160 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5154_6
timestamp 1731220469
transform 1 0 1992 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5153_6
timestamp 1731220469
transform 1 0 1992 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5152_6
timestamp 1731220469
transform 1 0 1784 0 1 3512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5151_6
timestamp 1731220469
transform 1 0 1784 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5150_6
timestamp 1731220469
transform 1 0 1648 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5149_6
timestamp 1731220469
transform 1 0 1488 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5148_6
timestamp 1731220469
transform 1 0 1336 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5147_6
timestamp 1731220469
transform 1 0 1184 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5146_6
timestamp 1731220469
transform 1 0 856 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5145_6
timestamp 1731220469
transform 1 0 680 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5144_6
timestamp 1731220469
transform 1 0 1288 0 1 3512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5143_6
timestamp 1731220469
transform 1 0 1544 0 1 3512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5142_6
timestamp 1731220469
transform 1 0 1456 0 -1 3488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5141_6
timestamp 1731220469
transform 1 0 1264 0 -1 3488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5140_6
timestamp 1731220469
transform 1 0 1312 0 1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5139_6
timestamp 1731220469
transform 1 0 1264 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5138_6
timestamp 1731220469
transform 1 0 1080 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5137_6
timestamp 1731220469
transform 1 0 1376 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5136_6
timestamp 1731220469
transform 1 0 1240 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5135_6
timestamp 1731220469
transform 1 0 1104 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5134_6
timestamp 1731220469
transform 1 0 968 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5133_6
timestamp 1731220469
transform 1 0 832 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5132_6
timestamp 1731220469
transform 1 0 696 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5131_6
timestamp 1731220469
transform 1 0 560 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5130_6
timestamp 1731220469
transform 1 0 696 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5129_6
timestamp 1731220469
transform 1 0 888 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5128_6
timestamp 1731220469
transform 1 0 1088 0 1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5127_6
timestamp 1731220469
transform 1 0 872 0 1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5126_6
timestamp 1731220469
transform 1 0 664 0 1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5125_6
timestamp 1731220469
transform 1 0 728 0 -1 3488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5124_6
timestamp 1731220469
transform 1 0 568 0 -1 3488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5123_6
timestamp 1731220469
transform 1 0 416 0 -1 3488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5122_6
timestamp 1731220469
transform 1 0 272 0 -1 3488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5121_6
timestamp 1731220469
transform 1 0 800 0 1 3512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5120_6
timestamp 1731220469
transform 1 0 568 0 1 3512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5119_6
timestamp 1731220469
transform 1 0 352 0 1 3512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5118_6
timestamp 1731220469
transform 1 0 144 0 1 3512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5117_6
timestamp 1731220469
transform 1 0 128 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5116_6
timestamp 1731220469
transform 1 0 496 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5115_6
timestamp 1731220469
transform 1 0 304 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5114_6
timestamp 1731220469
transform 1 0 304 0 1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5113_6
timestamp 1731220469
transform 1 0 128 0 1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5112_6
timestamp 1731220469
transform 1 0 512 0 1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5111_6
timestamp 1731220469
transform 1 0 720 0 1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5110_6
timestamp 1731220469
transform 1 0 632 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5109_6
timestamp 1731220469
transform 1 0 480 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5108_6
timestamp 1731220469
transform 1 0 952 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5107_6
timestamp 1731220469
transform 1 0 792 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5106_6
timestamp 1731220469
transform 1 0 728 0 1 4024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5105_6
timestamp 1731220469
transform 1 0 864 0 1 4024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5104_6
timestamp 1731220469
transform 1 0 1000 0 1 4024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5103_6
timestamp 1731220469
transform 1 0 1136 0 1 4024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5102_6
timestamp 1731220469
transform 1 0 1328 0 -1 4252
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5101_6
timestamp 1731220469
transform 1 0 1192 0 -1 4252
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5100_6
timestamp 1731220469
transform 1 0 1056 0 -1 4252
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_599_6
timestamp 1731220469
transform 1 0 920 0 -1 4252
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_598_6
timestamp 1731220469
transform 1 0 784 0 -1 4252
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_597_6
timestamp 1731220469
transform 1 0 1288 0 1 4268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_596_6
timestamp 1731220469
transform 1 0 1120 0 1 4268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_595_6
timestamp 1731220469
transform 1 0 960 0 1 4268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_594_6
timestamp 1731220469
transform 1 0 808 0 1 4268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_593_6
timestamp 1731220469
transform 1 0 664 0 1 4268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_592_6
timestamp 1731220469
transform 1 0 1376 0 -1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_591_6
timestamp 1731220469
transform 1 0 1112 0 -1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_590_6
timestamp 1731220469
transform 1 0 856 0 -1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_589_6
timestamp 1731220469
transform 1 0 624 0 -1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_588_6
timestamp 1731220469
transform 1 0 416 0 -1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_587_6
timestamp 1731220469
transform 1 0 1192 0 1 4500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_586_6
timestamp 1731220469
transform 1 0 904 0 1 4500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_585_6
timestamp 1731220469
transform 1 0 640 0 1 4500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_584_6
timestamp 1731220469
transform 1 0 392 0 1 4500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_583_6
timestamp 1731220469
transform 1 0 168 0 1 4500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_582_6
timestamp 1731220469
transform 1 0 1024 0 -1 4740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_581_6
timestamp 1731220469
transform 1 0 776 0 -1 4740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_580_6
timestamp 1731220469
transform 1 0 536 0 -1 4740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_579_6
timestamp 1731220469
transform 1 0 312 0 -1 4740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_578_6
timestamp 1731220469
transform 1 0 128 0 -1 4740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_577_6
timestamp 1731220469
transform 1 0 672 0 1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_576_6
timestamp 1731220469
transform 1 0 536 0 1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_575_6
timestamp 1731220469
transform 1 0 400 0 1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_574_6
timestamp 1731220469
transform 1 0 264 0 1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_573_6
timestamp 1731220469
transform 1 0 128 0 1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_572_6
timestamp 1731220469
transform 1 0 128 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_571_6
timestamp 1731220469
transform 1 0 312 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_570_6
timestamp 1731220469
transform 1 0 720 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_569_6
timestamp 1731220469
transform 1 0 520 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_568_6
timestamp 1731220469
transform 1 0 480 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_567_6
timestamp 1731220469
transform 1 0 344 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_566_6
timestamp 1731220469
transform 1 0 616 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_565_6
timestamp 1731220469
transform 1 0 752 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_564_6
timestamp 1731220469
transform 1 0 888 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_563_6
timestamp 1731220469
transform 1 0 1032 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_562_6
timestamp 1731220469
transform 1 0 1336 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_561_6
timestamp 1731220469
transform 1 0 1184 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_560_6
timestamp 1731220469
transform 1 0 1096 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_559_6
timestamp 1731220469
transform 1 0 912 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_558_6
timestamp 1731220469
transform 1 0 1280 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_557_6
timestamp 1731220469
transform 1 0 1456 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_556_6
timestamp 1731220469
transform 1 0 1632 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_555_6
timestamp 1731220469
transform 1 0 1784 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_554_6
timestamp 1731220469
transform 1 0 1648 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_553_6
timestamp 1731220469
transform 1 0 1488 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_552_6
timestamp 1731220469
transform 1 0 1784 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_551_6
timestamp 1731220469
transform 1 0 1992 0 1 4976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_550_6
timestamp 1731220469
transform 1 0 1992 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_549_6
timestamp 1731220469
transform 1 0 2128 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_548_6
timestamp 1731220469
transform 1 0 2664 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_547_6
timestamp 1731220469
transform 1 0 2480 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_546_6
timestamp 1731220469
transform 1 0 2296 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_545_6
timestamp 1731220469
transform 1 0 2192 0 1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_544_6
timestamp 1731220469
transform 1 0 2336 0 1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_543_6
timestamp 1731220469
transform 1 0 2488 0 1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_542_6
timestamp 1731220469
transform 1 0 2648 0 1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_541_6
timestamp 1731220469
transform 1 0 2816 0 1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_540_6
timestamp 1731220469
transform 1 0 2672 0 -1 5424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_539_6
timestamp 1731220469
transform 1 0 2480 0 -1 5424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_538_6
timestamp 1731220469
transform 1 0 2280 0 -1 5424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_537_6
timestamp 1731220469
transform 1 0 2136 0 1 5432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_536_6
timestamp 1731220469
transform 1 0 2352 0 1 5432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_535_6
timestamp 1731220469
transform 1 0 2560 0 1 5432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_534_6
timestamp 1731220469
transform 1 0 2520 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_533_6
timestamp 1731220469
transform 1 0 2336 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_532_6
timestamp 1731220469
transform 1 0 2152 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_531_6
timestamp 1731220469
transform 1 0 1992 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_530_6
timestamp 1731220469
transform 1 0 1784 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_529_6
timestamp 1731220469
transform 1 0 1512 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_528_6
timestamp 1731220469
transform 1 0 1736 0 -1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_527_6
timestamp 1731220469
transform 1 0 1480 0 -1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_526_6
timestamp 1731220469
transform 1 0 1232 0 -1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_525_6
timestamp 1731220469
transform 1 0 1256 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_524_6
timestamp 1731220469
transform 1 0 1488 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_523_6
timestamp 1731220469
transform 1 0 1512 0 -1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_522_6
timestamp 1731220469
transform 1 0 1376 0 -1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_521_6
timestamp 1731220469
transform 1 0 1240 0 -1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_520_6
timestamp 1731220469
transform 1 0 1104 0 -1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_519_6
timestamp 1731220469
transform 1 0 968 0 -1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_518_6
timestamp 1731220469
transform 1 0 832 0 -1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_517_6
timestamp 1731220469
transform 1 0 696 0 -1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_516_6
timestamp 1731220469
transform 1 0 560 0 -1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_515_6
timestamp 1731220469
transform 1 0 1032 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_514_6
timestamp 1731220469
transform 1 0 816 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_513_6
timestamp 1731220469
transform 1 0 608 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_512_6
timestamp 1731220469
transform 1 0 408 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_511_6
timestamp 1731220469
transform 1 0 984 0 -1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_510_6
timestamp 1731220469
transform 1 0 736 0 -1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_59_6
timestamp 1731220469
transform 1 0 488 0 -1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_58_6
timestamp 1731220469
transform 1 0 248 0 -1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_57_6
timestamp 1731220469
transform 1 0 1224 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_56_6
timestamp 1731220469
transform 1 0 952 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_55_6
timestamp 1731220469
transform 1 0 696 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_54_6
timestamp 1731220469
transform 1 0 472 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_53_6
timestamp 1731220469
transform 1 0 272 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_52_6
timestamp 1731220469
transform 1 0 128 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_51_6
timestamp 1731220469
transform 1 0 264 0 -1 5756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_50_6
timestamp 1731220469
transform 1 0 128 0 -1 5756
box 3 5 132 108
<< end >>
